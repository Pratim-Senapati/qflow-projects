magic
tech scmos
magscale 1 2
timestamp 1740717622
<< nwell >>
rect -10 96 106 210
rect 12 88 66 96
<< ntransistor >>
rect 14 20 18 40
rect 30 20 34 60
rect 40 20 44 60
rect 56 20 60 60
rect 66 20 70 60
<< ptransistor >>
rect 14 140 18 180
rect 30 100 34 180
rect 40 100 44 180
rect 56 108 60 188
rect 66 108 70 188
<< ndiffusion >>
rect 24 56 30 60
rect 20 52 30 56
rect 4 39 14 40
rect 12 21 14 39
rect 4 20 14 21
rect 18 24 20 40
rect 28 24 30 52
rect 18 20 30 24
rect 34 20 40 60
rect 44 52 56 60
rect 44 24 46 52
rect 54 24 56 52
rect 44 20 56 24
rect 60 20 66 60
rect 70 59 80 60
rect 70 21 72 59
rect 70 20 80 21
<< pdiffusion >>
rect 46 184 56 188
rect 4 179 14 180
rect 12 141 14 179
rect 4 140 14 141
rect 18 140 20 180
rect 28 112 30 180
rect 24 100 30 112
rect 34 100 40 180
rect 44 116 46 180
rect 54 116 56 184
rect 44 108 56 116
rect 60 108 66 188
rect 70 187 80 188
rect 70 109 72 187
rect 70 108 80 109
rect 44 100 50 108
<< ndcontact >>
rect 4 21 12 39
rect 20 24 28 52
rect 46 24 54 52
rect 72 21 80 59
<< pdcontact >>
rect 4 141 12 179
rect 20 112 28 180
rect 46 116 54 184
rect 72 109 80 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
<< polysilicon >>
rect 14 190 44 194
rect 14 180 18 190
rect 30 180 34 184
rect 40 180 44 190
rect 56 188 60 192
rect 66 188 70 192
rect 14 138 18 140
rect 8 134 18 138
rect 8 86 12 134
rect 30 98 34 100
rect 24 94 34 98
rect 40 96 44 100
rect 24 86 28 94
rect 56 80 60 108
rect 66 106 70 108
rect 66 102 72 106
rect 8 46 12 78
rect 22 66 26 78
rect 50 76 60 80
rect 40 68 48 72
rect 22 62 34 66
rect 30 60 34 62
rect 40 60 44 68
rect 68 66 72 94
rect 56 60 60 64
rect 66 62 72 66
rect 66 60 70 62
rect 8 42 18 46
rect 14 40 18 42
rect 14 10 18 20
rect 30 16 34 20
rect 40 16 44 20
rect 56 10 60 20
rect 66 16 70 20
rect 14 6 60 10
<< polycontact >>
rect 4 78 12 86
rect 20 78 28 86
rect 42 72 50 80
rect 68 94 76 102
<< metal1 >>
rect -4 204 100 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 100 204
rect -4 194 100 196
rect 20 180 28 194
rect 4 179 12 180
rect 4 140 12 141
rect 4 106 10 140
rect 46 184 54 188
rect 72 187 80 194
rect 54 116 62 118
rect 46 112 62 116
rect 4 100 42 106
rect 4 86 12 94
rect 20 86 28 94
rect 36 72 42 100
rect 56 74 62 112
rect 72 108 80 109
rect 68 86 76 94
rect 36 68 46 72
rect 4 62 46 68
rect 56 66 76 74
rect 4 40 10 62
rect 56 60 62 66
rect 54 56 62 60
rect 20 52 28 56
rect 4 39 12 40
rect 4 20 12 21
rect 20 6 28 24
rect 46 52 62 56
rect 54 50 62 52
rect 72 59 80 60
rect 46 20 54 24
rect 72 6 80 21
rect -4 4 100 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 100 4
rect -4 -6 100 -4
<< m1p >>
rect 4 86 12 94
rect 20 86 28 94
rect 68 86 76 94
rect 68 66 76 74
<< labels >>
rlabel metal1 8 90 8 90 4 S
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 72 70 72 70 4 Y
rlabel metal1 72 90 72 90 4 A
rlabel metal1 24 90 24 90 4 B
<< end >>

magic
tech scmos
magscale 1 2
timestamp 1740717622
<< nwell >>
rect -14 96 136 210
<< ntransistor >>
rect 30 12 34 32
rect 46 12 50 32
rect 62 12 66 32
<< ptransistor >>
rect 14 128 18 188
rect 30 128 34 188
rect 46 128 50 188
rect 62 128 66 188
rect 94 120 98 180
rect 110 120 114 180
<< ndiffusion >>
rect 20 31 30 32
rect 28 13 30 31
rect 20 12 30 13
rect 34 31 46 32
rect 34 13 36 31
rect 44 13 46 31
rect 34 12 46 13
rect 50 24 62 32
rect 50 16 52 24
rect 60 16 62 24
rect 50 12 62 16
rect 66 31 76 32
rect 66 13 68 31
rect 66 12 76 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 129 14 187
rect 4 128 14 129
rect 18 187 30 188
rect 18 129 20 187
rect 28 129 30 187
rect 18 128 30 129
rect 34 187 46 188
rect 34 129 36 187
rect 44 129 46 187
rect 34 128 46 129
rect 50 176 62 188
rect 50 128 52 176
rect 60 128 62 176
rect 66 130 68 188
rect 84 179 94 180
rect 66 128 72 130
rect 92 121 94 179
rect 84 120 94 121
rect 98 172 110 180
rect 98 124 100 172
rect 108 124 110 172
rect 98 120 110 124
rect 114 179 124 180
rect 114 121 116 179
rect 114 120 124 121
<< ndcontact >>
rect 20 13 28 31
rect 36 13 44 31
rect 52 16 60 24
rect 68 13 76 31
<< pdcontact >>
rect 4 129 12 187
rect 20 129 28 187
rect 36 129 44 187
rect 52 128 60 176
rect 68 130 76 188
rect 84 121 92 179
rect 100 124 108 172
rect 116 121 124 179
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
rect 92 -4 100 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
rect 92 196 100 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 46 188 50 192
rect 62 188 66 192
rect 94 180 98 184
rect 110 180 114 184
rect 14 126 18 128
rect 30 126 34 128
rect 46 126 50 128
rect 62 126 66 128
rect 14 122 34 126
rect 30 54 34 122
rect 44 122 66 126
rect 44 74 48 122
rect 94 118 98 120
rect 110 118 114 120
rect 94 114 114 118
rect 94 112 98 114
rect 62 108 98 112
rect 62 94 66 108
rect 30 32 34 46
rect 46 32 50 66
rect 62 32 66 86
rect 30 8 34 12
rect 46 8 50 12
rect 62 8 66 12
<< polycontact >>
rect 60 86 68 94
rect 44 66 52 74
rect 30 46 38 54
<< metal1 >>
rect -4 204 132 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 92 204
rect 100 196 132 204
rect -4 194 132 196
rect 4 187 12 188
rect 4 128 12 129
rect 20 187 28 194
rect 20 128 28 129
rect 36 187 68 188
rect 44 182 68 187
rect 36 128 44 129
rect 86 182 122 188
rect 86 180 92 182
rect 84 179 92 180
rect 6 122 12 128
rect 36 122 42 128
rect 6 116 42 122
rect 54 124 60 128
rect 54 121 84 124
rect 116 180 122 182
rect 116 179 124 180
rect 54 120 92 121
rect 100 172 108 176
rect 100 120 108 124
rect 116 120 124 121
rect 54 118 90 120
rect 100 114 106 120
rect 100 112 108 114
rect 74 106 108 112
rect 52 86 60 94
rect 36 66 44 74
rect 20 46 30 54
rect 74 40 80 106
rect 40 34 80 40
rect 40 32 46 34
rect 20 31 28 32
rect 20 6 28 13
rect 36 31 46 32
rect 44 26 46 31
rect 68 32 80 34
rect 68 31 76 32
rect 36 12 44 13
rect 52 24 60 28
rect 52 6 60 16
rect 68 12 76 13
rect -4 4 132 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 92 4
rect 100 -4 132 4
rect -4 -6 132 -4
<< m1p >>
rect 100 106 108 114
rect 52 86 60 94
rect 36 66 44 74
rect 20 46 28 54
<< labels >>
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 40 70 40 70 4 B
rlabel metal1 56 90 56 90 4 C
rlabel metal1 24 50 24 50 4 A
rlabel metal1 104 110 104 110 4 Y
<< end >>

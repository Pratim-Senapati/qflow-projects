magic
tech scmos
magscale 1 2
timestamp 1743590271
<< metal1 >>
rect 552 606 558 614
rect 566 606 572 614
rect 580 606 586 614
rect 594 606 600 614
rect 669 577 691 583
rect 462 537 492 543
rect 77 517 124 523
rect 132 457 147 463
rect 45 437 67 443
rect 264 406 270 414
rect 278 406 284 414
rect 292 406 298 414
rect 306 406 312 414
rect 716 303 724 308
rect 541 297 563 303
rect 701 297 724 303
rect 404 277 419 283
rect 509 277 531 283
rect 525 257 531 277
rect 564 277 579 283
rect 621 277 675 283
rect 685 277 700 283
rect 621 263 627 277
rect 813 277 844 283
rect 589 257 627 263
rect 452 236 456 244
rect 552 206 558 214
rect 566 206 572 214
rect 580 206 586 214
rect 594 206 600 214
rect 333 157 396 163
rect 264 6 270 14
rect 278 6 284 14
rect 292 6 298 14
rect 306 6 312 14
<< m2contact >>
rect 558 606 566 614
rect 572 606 580 614
rect 586 606 594 614
rect 540 576 548 584
rect 732 576 740 584
rect 780 576 788 584
rect 300 556 308 564
rect 668 558 676 566
rect 812 556 820 564
rect 12 536 20 544
rect 268 536 276 544
rect 492 536 500 544
rect 588 536 596 544
rect 124 516 132 524
rect 172 516 180 524
rect 652 516 660 524
rect 700 516 708 524
rect 748 516 756 524
rect 12 496 20 504
rect 204 500 212 508
rect 124 456 132 464
rect 204 454 212 462
rect 28 436 36 444
rect 796 436 804 444
rect 270 406 278 414
rect 284 406 292 414
rect 298 406 306 414
rect 44 376 52 384
rect 332 336 340 344
rect 748 336 756 344
rect 44 316 52 324
rect 716 316 724 324
rect 44 296 52 304
rect 732 296 740 304
rect 780 296 788 304
rect 140 276 148 284
rect 396 276 404 284
rect 172 256 180 264
rect 556 276 564 284
rect 700 276 708 284
rect 844 276 852 284
rect 652 256 660 264
rect 748 256 756 264
rect 444 236 452 244
rect 558 206 566 214
rect 572 206 580 214
rect 586 206 594 214
rect 828 176 836 184
rect 172 156 180 164
rect 396 156 404 164
rect 668 156 676 164
rect 140 136 148 144
rect 636 136 644 144
rect 44 116 52 124
rect 252 116 260 124
rect 444 116 452 124
rect 540 116 548 124
rect 44 96 52 104
rect 572 100 580 108
rect 572 54 580 62
rect 44 36 52 44
rect 412 36 420 44
rect 270 6 278 14
rect 284 6 292 14
rect 298 6 306 14
<< metal2 >>
rect 301 637 323 643
rect 605 637 627 643
rect 717 637 739 643
rect 765 637 787 643
rect 269 544 275 576
rect 301 564 307 637
rect 552 606 558 614
rect 566 606 572 614
rect 580 606 586 614
rect 594 606 600 614
rect 621 564 627 637
rect 733 584 739 637
rect 781 584 787 637
rect 660 558 668 563
rect 660 557 675 558
rect 13 504 19 516
rect 29 444 35 516
rect 125 464 131 516
rect 301 504 307 556
rect 589 524 595 536
rect 653 524 659 556
rect 701 524 707 536
rect 813 524 819 556
rect 820 517 835 523
rect 29 303 35 436
rect 45 324 51 376
rect 29 297 44 303
rect 45 124 51 296
rect 173 264 179 496
rect 205 462 211 500
rect 264 406 270 414
rect 278 406 284 414
rect 292 406 298 414
rect 306 406 312 414
rect 141 144 147 176
rect 173 164 179 256
rect 397 164 403 276
rect 653 264 659 336
rect 701 304 707 516
rect 717 324 723 516
rect 781 304 787 336
rect 701 284 707 296
rect 445 184 451 236
rect 552 206 558 214
rect 566 206 572 214
rect 580 206 586 214
rect 594 206 600 214
rect 253 124 259 136
rect 397 124 403 156
rect 797 144 803 436
rect 829 184 835 517
rect 845 284 851 296
rect 541 124 547 136
rect 45 44 51 96
rect 573 62 579 100
rect 264 6 270 14
rect 278 6 284 14
rect 292 6 298 14
rect 306 6 312 14
rect 413 -17 419 36
rect 413 -23 435 -17
<< m3contact >>
rect 268 576 276 584
rect 558 606 566 614
rect 572 606 580 614
rect 586 606 594 614
rect 540 576 548 584
rect 620 556 628 564
rect 652 556 660 564
rect 12 536 20 544
rect 12 516 20 524
rect 28 516 36 524
rect 172 516 180 524
rect 172 496 180 504
rect 492 536 500 544
rect 700 536 708 544
rect 588 516 596 524
rect 716 516 724 524
rect 748 516 756 524
rect 812 516 820 524
rect 140 276 148 284
rect 300 496 308 504
rect 270 406 278 414
rect 284 406 292 414
rect 298 406 306 414
rect 332 336 340 344
rect 652 336 660 344
rect 556 276 564 284
rect 140 176 148 184
rect 748 336 756 344
rect 780 336 788 344
rect 700 296 708 304
rect 732 296 740 304
rect 476 256 484 264
rect 748 256 756 264
rect 558 206 566 214
rect 572 206 580 214
rect 586 206 594 214
rect 444 176 452 184
rect 172 156 180 164
rect 668 156 676 164
rect 252 136 260 144
rect 844 296 852 304
rect 540 136 548 144
rect 636 136 644 144
rect 796 136 804 144
rect 396 116 404 124
rect 444 116 452 124
rect 270 6 278 14
rect 284 6 292 14
rect 298 6 306 14
<< metal3 >>
rect 552 614 600 616
rect 552 606 556 614
rect 566 606 572 614
rect 580 606 586 614
rect 596 606 600 614
rect 552 604 600 606
rect 276 577 540 583
rect 628 557 652 563
rect 500 537 700 543
rect -19 517 12 523
rect 36 517 172 523
rect 596 517 716 523
rect 724 517 748 523
rect 756 517 812 523
rect -19 497 12 503
rect 180 497 300 503
rect 264 414 312 416
rect 264 406 268 414
rect 278 406 284 414
rect 292 406 298 414
rect 308 406 312 414
rect 264 404 312 406
rect 340 337 652 343
rect 660 337 748 343
rect 756 337 780 343
rect 708 297 732 303
rect 852 297 883 303
rect 148 277 556 283
rect 484 257 748 263
rect 552 214 600 216
rect 552 206 556 214
rect 566 206 572 214
rect 580 206 586 214
rect 596 206 600 214
rect 552 204 600 206
rect 148 177 444 183
rect 180 157 668 163
rect 260 137 540 143
rect 644 137 796 143
rect 404 117 444 123
rect 264 14 312 16
rect 264 6 268 14
rect 278 6 284 14
rect 292 6 298 14
rect 308 6 312 14
rect 264 4 312 6
<< m4contact >>
rect 556 606 558 614
rect 558 606 564 614
rect 572 606 580 614
rect 588 606 594 614
rect 594 606 596 614
rect 12 536 20 544
rect 12 496 20 504
rect 268 406 270 414
rect 270 406 276 414
rect 284 406 292 414
rect 300 406 306 414
rect 306 406 308 414
rect 556 206 558 214
rect 558 206 564 214
rect 572 206 580 214
rect 588 206 594 214
rect 594 206 596 214
rect 268 6 270 14
rect 270 6 276 14
rect 284 6 292 14
rect 300 6 306 14
rect 306 6 308 14
<< metal4 >>
rect 10 544 22 546
rect 10 536 12 544
rect 20 536 22 544
rect 10 504 22 536
rect 10 496 12 504
rect 20 496 22 504
rect 10 494 22 496
rect 264 414 312 640
rect 264 406 268 414
rect 276 406 284 414
rect 292 406 300 414
rect 308 406 312 414
rect 264 14 312 406
rect 264 6 268 14
rect 276 6 284 14
rect 292 6 300 14
rect 308 6 312 14
rect 264 -40 312 6
rect 552 614 600 640
rect 552 606 556 614
rect 564 606 572 614
rect 580 606 588 614
rect 596 606 600 614
rect 552 214 600 606
rect 552 206 556 214
rect 564 206 572 214
rect 580 206 588 214
rect 596 206 600 214
rect 552 -40 600 206
use DFFSR  DFFSR_4
timestamp 1743590271
transform 1 0 8 0 -1 210
box -4 -6 356 206
use FILL  FILL_0_0_0
timestamp 1743590271
transform -1 0 376 0 -1 210
box -4 -6 20 206
use DFFSR  DFFSR_3
timestamp 1743590271
transform 1 0 8 0 1 210
box -4 -6 356 206
use FILL  FILL_1_0_0
timestamp 1743590271
transform -1 0 376 0 1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1743590271
transform -1 0 392 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1743590271
transform -1 0 408 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_4
timestamp 1743590271
transform -1 0 456 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_1_0
timestamp 1743590271
transform 1 0 456 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1743590271
transform -1 0 392 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_2
timestamp 1743590271
transform -1 0 408 0 1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1743590271
transform 1 0 472 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_2
timestamp 1743590271
transform 1 0 488 0 -1 210
box -4 -6 20 206
use INVX1  INVX1_2
timestamp 1743590271
transform 1 0 520 0 1 210
box -4 -6 36 206
use XNOR2X1  XNOR2X1_1
timestamp 1743590271
transform -1 0 520 0 1 210
box -4 -6 116 206
use NAND3X1  NAND3X1_1
timestamp 1743590271
transform 1 0 712 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_1
timestamp 1743590271
transform -1 0 712 0 1 210
box -4 -6 68 206
use FILL  FILL_1_1_2
timestamp 1743590271
transform -1 0 648 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_1
timestamp 1743590271
transform -1 0 632 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_0
timestamp 1743590271
transform -1 0 616 0 1 210
box -4 -6 20 206
use NOR2X1  NOR2X1_1
timestamp 1743590271
transform -1 0 600 0 1 210
box -4 -6 52 206
use DFFSR  DFFSR_1
timestamp 1743590271
transform 1 0 504 0 -1 210
box -4 -6 356 206
use BUFX2  BUFX2_3
timestamp 1743590271
transform 1 0 776 0 1 210
box -4 -6 52 206
use FILL  FILL_2_1
timestamp 1743590271
transform 1 0 824 0 1 210
box -4 -6 20 206
use FILL  FILL_2_2
timestamp 1743590271
transform 1 0 840 0 1 210
box -4 -6 20 206
use INVX2  INVX2_1
timestamp 1743590271
transform 1 0 8 0 -1 610
box -4 -6 36 206
use BUFX2  BUFX2_6
timestamp 1743590271
transform -1 0 88 0 -1 610
box -4 -6 52 206
use FILL  FILL_2_0_0
timestamp 1743590271
transform 1 0 88 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1743590271
transform 1 0 104 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1743590271
transform 1 0 120 0 -1 610
box -4 -6 20 206
use DFFSR  DFFSR_2
timestamp 1743590271
transform 1 0 136 0 -1 610
box -4 -6 356 206
use XOR2X1  XOR2X1_1
timestamp 1743590271
transform -1 0 600 0 -1 610
box -4 -6 116 206
use FILL  FILL_2_1_0
timestamp 1743590271
transform 1 0 600 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1743590271
transform 1 0 616 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1743590271
transform 1 0 632 0 -1 610
box -4 -6 20 206
use BUFX2  BUFX2_5
timestamp 1743590271
transform 1 0 648 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_2
timestamp 1743590271
transform 1 0 696 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_1
timestamp 1743590271
transform 1 0 744 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_1
timestamp 1743590271
transform -1 0 824 0 -1 610
box -4 -6 36 206
use FILL  FILL_3_1
timestamp 1743590271
transform -1 0 840 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_2
timestamp 1743590271
transform -1 0 856 0 -1 610
box -4 -6 20 206
<< labels >>
flabel metal3 s -16 520 -16 520 7 FreeSans 24 0 0 0 vdd
port 0 nsew
flabel metal2 s 608 640 608 640 3 FreeSans 24 90 0 0 gnd
port 1 nsew
flabel metal2 s 317 637 323 643 3 FreeSans 24 90 0 0 clk
port 2 nsew
flabel metal3 s -19 497 -13 503 7 FreeSans 24 0 0 0 rst
port 3 nsew
flabel metal2 s 765 637 771 643 3 FreeSans 24 90 0 0 count[0]
port 4 nsew
flabel metal2 s 717 637 723 643 3 FreeSans 24 90 0 0 count[1]
port 5 nsew
flabel metal3 s 877 297 883 303 3 FreeSans 24 0 0 0 count[2]
port 6 nsew
flabel metal2 s 429 -23 435 -17 7 FreeSans 24 270 0 0 count[3]
port 7 nsew
<< end >>

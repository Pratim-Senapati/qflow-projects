magic
tech scmos
magscale 1 2
timestamp 1740717622
<< nwell >>
rect -14 96 70 210
<< ntransistor >>
rect 14 12 18 32
rect 30 12 34 32
rect 46 12 50 52
<< ptransistor >>
rect 14 108 18 188
rect 24 108 28 188
rect 40 108 44 188
<< ndiffusion >>
rect 40 48 46 52
rect 36 44 46 48
rect 4 31 14 32
rect 12 13 14 31
rect 4 12 14 13
rect 18 31 30 32
rect 18 13 20 31
rect 28 13 30 31
rect 18 12 30 13
rect 34 16 36 32
rect 44 16 46 44
rect 34 12 46 16
rect 50 51 60 52
rect 50 13 52 51
rect 50 12 60 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 109 14 187
rect 4 108 14 109
rect 18 108 24 188
rect 28 187 40 188
rect 28 109 30 187
rect 38 109 40 187
rect 28 108 40 109
rect 44 187 54 188
rect 44 109 46 187
rect 44 108 54 109
<< ndcontact >>
rect 4 13 12 31
rect 20 13 28 31
rect 36 16 44 44
rect 52 13 60 51
<< pdcontact >>
rect 4 109 12 187
rect 30 109 38 187
rect 46 109 54 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
<< polysilicon >>
rect 14 188 18 192
rect 24 188 28 192
rect 40 188 44 192
rect 14 106 18 108
rect 12 102 18 106
rect 12 38 16 102
rect 24 82 28 108
rect 40 102 44 108
rect 40 98 50 102
rect 32 74 34 78
rect 12 34 18 38
rect 14 32 18 34
rect 30 32 34 74
rect 46 52 50 98
rect 14 8 18 12
rect 30 8 34 12
rect 46 8 50 12
<< polycontact >>
rect 4 38 12 46
rect 38 90 46 98
rect 24 74 32 82
<< metal1 >>
rect -4 204 68 206
rect 4 196 28 204
rect 36 196 68 204
rect -4 194 68 196
rect 4 187 12 188
rect 4 102 12 109
rect 30 187 38 194
rect 30 108 38 109
rect 46 187 54 188
rect 54 109 60 114
rect 46 108 60 109
rect 4 98 44 102
rect 4 96 38 98
rect 54 94 60 108
rect 20 66 30 74
rect 40 60 46 90
rect 52 86 60 94
rect 22 54 46 60
rect 4 46 12 54
rect 22 32 28 54
rect 54 52 60 86
rect 52 51 60 52
rect 4 31 12 32
rect 4 6 12 13
rect 20 31 28 32
rect 20 12 28 13
rect 36 44 44 48
rect 36 6 44 16
rect 52 12 60 13
rect -4 4 68 6
rect 4 -4 28 4
rect 36 -4 68 4
rect -4 -6 68 -4
<< m1p >>
rect 52 86 60 94
rect 20 66 28 74
rect 4 46 12 54
<< labels >>
rlabel metal1 56 90 56 90 4 Y
rlabel metal1 24 70 24 70 4 B
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 50 8 50 4 A
<< end >>

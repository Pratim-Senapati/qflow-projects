magic
tech scmos
magscale 1 2
timestamp 1739819275
<< checkpaint >>
rect -79 -100 2351 2103
<< metal1 >>
rect 408 2006 412 2014
rect 420 2006 424 2014
rect 1336 2006 1340 2014
rect 1348 2006 1352 2014
rect 90 1936 92 1944
rect 381 1937 403 1943
rect 317 1917 332 1923
rect 381 1923 387 1937
rect 372 1917 387 1923
rect 61 1903 67 1916
rect 61 1897 83 1903
rect 477 1897 547 1903
rect 845 1903 851 1923
rect 845 1897 899 1903
rect 909 1897 947 1903
rect 1021 1903 1027 1923
rect 1012 1897 1027 1903
rect 1133 1897 1170 1903
rect 1934 1897 1987 1903
rect 61 1877 76 1883
rect 260 1877 280 1883
rect 637 1877 659 1883
rect 669 1877 707 1883
rect 653 1864 659 1877
rect 964 1877 995 1883
rect 1060 1877 1075 1883
rect 2093 1883 2099 1903
rect 2132 1897 2147 1903
rect 2164 1897 2179 1903
rect 2068 1877 2099 1883
rect 2205 1877 2252 1883
rect 189 1857 211 1863
rect 612 1856 620 1864
rect 1156 1857 1171 1863
rect 2100 1857 2115 1863
rect 138 1836 140 1844
rect 365 1837 380 1843
rect 872 1806 876 1814
rect 884 1806 888 1814
rect 1864 1806 1868 1814
rect 1876 1806 1880 1814
rect 1764 1776 1766 1784
rect 884 1757 899 1763
rect 1885 1757 1900 1763
rect 125 1737 140 1743
rect 756 1737 771 1743
rect 1149 1737 1171 1743
rect 1165 1724 1171 1737
rect 1661 1737 1708 1743
rect 45 1717 99 1723
rect 605 1717 643 1723
rect 637 1697 643 1717
rect 692 1717 723 1723
rect 733 1717 764 1723
rect 804 1717 819 1723
rect 909 1717 947 1723
rect 973 1717 1011 1723
rect 973 1697 979 1717
rect 1092 1717 1107 1723
rect 148 1677 163 1683
rect 948 1636 950 1644
rect 1066 1636 1068 1644
rect 408 1606 412 1614
rect 420 1606 424 1614
rect 1336 1606 1340 1614
rect 1348 1606 1352 1614
rect 132 1576 134 1584
rect 573 1497 611 1503
rect 701 1497 716 1503
rect 1773 1497 1811 1503
rect 2174 1497 2211 1503
rect 77 1477 108 1483
rect 653 1477 668 1483
rect 1566 1477 1603 1483
rect 1773 1477 1788 1483
rect 2237 1477 2252 1483
rect 1196 1464 1204 1468
rect 1565 1457 1580 1463
rect 1821 1457 1836 1463
rect 1636 1436 1640 1444
rect 872 1406 876 1414
rect 884 1406 888 1414
rect 1864 1406 1868 1414
rect 1876 1406 1880 1414
rect 260 1357 275 1363
rect 413 1357 435 1363
rect 1796 1357 1820 1363
rect 1828 1357 1843 1363
rect 93 1337 124 1343
rect 141 1337 195 1343
rect 1188 1337 1203 1343
rect 1476 1337 1491 1343
rect 1508 1337 1523 1343
rect 1748 1337 1779 1343
rect 413 1317 428 1323
rect 676 1317 706 1323
rect 1556 1317 1603 1323
rect 1629 1297 1644 1303
rect 564 1277 579 1283
rect 2205 1277 2252 1283
rect 408 1206 412 1214
rect 420 1206 424 1214
rect 1336 1206 1340 1214
rect 1348 1206 1352 1214
rect 676 1137 732 1143
rect 45 1097 82 1103
rect 573 1097 611 1103
rect 772 1097 787 1103
rect 1284 1097 1299 1103
rect 509 1077 563 1083
rect 1101 1077 1132 1083
rect 2221 1077 2252 1083
rect 557 1057 572 1063
rect 1178 1036 1180 1044
rect 872 1006 876 1014
rect 884 1006 888 1014
rect 1864 1006 1868 1014
rect 1876 1006 1880 1014
rect 285 944 291 963
rect 349 957 387 963
rect 2212 956 2214 964
rect 292 937 307 943
rect 1437 937 1452 943
rect 1661 937 1676 943
rect 260 917 275 923
rect 445 917 483 923
rect 29 897 51 903
rect 477 897 483 917
rect 589 917 604 923
rect 1005 917 1042 923
rect 1421 917 1436 923
rect 1668 917 1699 923
rect 1604 896 1608 904
rect 189 877 252 883
rect 408 806 412 814
rect 420 806 424 814
rect 1336 806 1340 814
rect 1348 806 1352 814
rect 541 743 547 763
rect 541 737 611 743
rect 666 736 668 744
rect 2205 737 2252 743
rect 604 724 612 728
rect 765 703 771 723
rect 676 697 723 703
rect 733 697 771 703
rect 781 697 812 703
rect 1997 697 2019 703
rect 2061 677 2099 683
rect 1933 657 1980 663
rect 2061 657 2067 677
rect 872 606 876 614
rect 884 606 888 614
rect 1864 606 1868 614
rect 1876 606 1880 614
rect 420 557 435 563
rect 1709 557 1731 563
rect 2212 557 2227 563
rect 445 537 460 543
rect 1645 537 1683 543
rect 45 517 82 523
rect 1764 517 1811 523
rect 548 497 563 503
rect 1236 497 1299 503
rect 1213 477 1244 483
rect 1812 436 1814 444
rect 408 406 412 414
rect 420 406 424 414
rect 1336 406 1340 414
rect 1348 406 1352 414
rect 1620 337 1635 343
rect 372 297 387 303
rect 964 297 979 303
rect 1501 297 1539 303
rect 2141 297 2179 303
rect 2196 297 2211 303
rect 461 277 483 283
rect 900 277 931 283
rect 1028 277 1043 283
rect 1524 277 1539 283
rect 1972 277 2003 283
rect 2013 277 2060 283
rect 2237 277 2252 283
rect 1437 257 1484 263
rect 872 206 876 214
rect 884 206 888 214
rect 1864 206 1868 214
rect 1876 206 1880 214
rect 372 157 387 163
rect 397 157 412 163
rect 452 157 483 163
rect 1428 137 1443 143
rect 413 117 435 123
rect 1294 117 1324 123
rect 1405 117 1443 123
rect 1588 117 1603 123
rect 2158 117 2195 123
rect 2221 77 2252 83
rect 1357 37 1372 43
rect 408 6 412 14
rect 420 6 424 14
rect 1336 6 1340 14
rect 1348 6 1352 14
<< m2contact >>
rect 412 2006 420 2014
rect 1340 2006 1348 2014
rect 764 1976 772 1984
rect 1100 1976 1108 1984
rect 1452 1976 1460 1984
rect 1548 1976 1556 1984
rect 1564 1976 1572 1984
rect 2012 1976 2020 1984
rect 1676 1958 1684 1966
rect 92 1936 100 1944
rect 284 1936 292 1944
rect 60 1916 68 1924
rect 124 1916 132 1924
rect 332 1916 340 1924
rect 364 1916 372 1924
rect 444 1936 452 1944
rect 604 1916 612 1924
rect 748 1916 756 1924
rect 28 1896 36 1904
rect 252 1896 260 1904
rect 300 1896 308 1904
rect 396 1896 404 1904
rect 684 1896 692 1904
rect 716 1896 724 1904
rect 796 1896 804 1904
rect 828 1896 836 1904
rect 876 1916 884 1924
rect 1004 1896 1012 1904
rect 1452 1916 1460 1924
rect 1676 1912 1684 1920
rect 1452 1896 1460 1904
rect 1516 1896 1524 1904
rect 1596 1896 1604 1904
rect 1628 1896 1636 1904
rect 1852 1896 1860 1904
rect 2076 1896 2084 1904
rect 12 1876 20 1884
rect 76 1876 84 1884
rect 156 1876 164 1884
rect 236 1876 244 1884
rect 252 1876 260 1884
rect 332 1876 340 1884
rect 492 1876 500 1884
rect 508 1876 516 1884
rect 556 1876 564 1884
rect 748 1876 756 1884
rect 812 1876 820 1884
rect 924 1876 932 1884
rect 956 1876 964 1884
rect 1052 1876 1060 1884
rect 1356 1876 1364 1884
rect 1740 1876 1748 1884
rect 2060 1876 2068 1884
rect 2124 1896 2132 1904
rect 2156 1896 2164 1904
rect 2252 1876 2260 1884
rect 108 1856 116 1864
rect 172 1856 180 1864
rect 428 1856 436 1864
rect 588 1856 596 1864
rect 604 1856 612 1864
rect 652 1856 660 1864
rect 956 1856 964 1864
rect 972 1856 980 1864
rect 1084 1856 1092 1864
rect 1148 1856 1156 1864
rect 1324 1856 1332 1864
rect 1772 1856 1780 1864
rect 2028 1856 2036 1864
rect 2092 1856 2100 1864
rect 2124 1856 2132 1864
rect 2156 1856 2164 1864
rect 140 1836 148 1844
rect 220 1836 228 1844
rect 380 1836 388 1844
rect 444 1836 452 1844
rect 524 1836 532 1844
rect 572 1836 580 1844
rect 1020 1836 1028 1844
rect 1932 1836 1940 1844
rect 2044 1836 2052 1844
rect 876 1806 884 1814
rect 1868 1806 1876 1814
rect 1244 1776 1252 1784
rect 1644 1776 1652 1784
rect 1756 1776 1764 1784
rect 1852 1776 1860 1784
rect 2236 1776 2244 1784
rect 316 1756 324 1764
rect 876 1756 884 1764
rect 1084 1756 1092 1764
rect 1196 1756 1204 1764
rect 1436 1756 1444 1764
rect 1628 1756 1636 1764
rect 1692 1756 1700 1764
rect 1900 1756 1908 1764
rect 2076 1756 2084 1764
rect 12 1736 20 1744
rect 76 1736 84 1744
rect 140 1736 148 1744
rect 348 1736 356 1744
rect 572 1736 580 1744
rect 636 1736 644 1744
rect 684 1736 692 1744
rect 748 1736 756 1744
rect 860 1736 868 1744
rect 924 1736 932 1744
rect 1036 1736 1044 1744
rect 1180 1736 1188 1744
rect 1404 1736 1412 1744
rect 1598 1736 1606 1744
rect 1708 1736 1716 1744
rect 2044 1736 2052 1744
rect 28 1716 36 1724
rect 236 1716 244 1724
rect 540 1716 548 1724
rect 588 1716 596 1724
rect 60 1696 68 1704
rect 124 1696 132 1704
rect 444 1696 452 1704
rect 556 1696 564 1704
rect 620 1696 628 1704
rect 668 1716 676 1724
rect 684 1716 692 1724
rect 764 1716 772 1724
rect 796 1716 804 1724
rect 700 1696 708 1704
rect 1020 1716 1028 1724
rect 1052 1716 1060 1724
rect 1084 1716 1092 1724
rect 1132 1716 1140 1724
rect 1164 1716 1172 1724
rect 1212 1716 1220 1724
rect 1308 1716 1316 1724
rect 1676 1716 1684 1724
rect 1724 1716 1732 1724
rect 1740 1716 1748 1724
rect 1788 1716 1796 1724
rect 1820 1716 1828 1724
rect 1868 1716 1876 1724
rect 1980 1716 1988 1724
rect 988 1696 996 1704
rect 1308 1696 1316 1704
rect 1948 1696 1956 1704
rect 140 1676 148 1684
rect 524 1676 532 1684
rect 444 1636 452 1644
rect 540 1636 548 1644
rect 940 1636 948 1644
rect 1068 1636 1076 1644
rect 1308 1636 1316 1644
rect 1948 1636 1956 1644
rect 412 1606 420 1614
rect 1340 1606 1348 1614
rect 124 1576 132 1584
rect 204 1576 212 1584
rect 1052 1576 1060 1584
rect 1276 1576 1284 1584
rect 492 1556 500 1564
rect 796 1558 804 1566
rect 1916 1558 1924 1566
rect 156 1516 164 1524
rect 204 1516 212 1524
rect 540 1516 548 1524
rect 796 1512 804 1520
rect 1276 1516 1284 1524
rect 1916 1512 1924 1520
rect 44 1496 52 1504
rect 60 1496 68 1504
rect 124 1496 132 1504
rect 236 1496 244 1504
rect 412 1496 420 1504
rect 716 1496 724 1504
rect 780 1496 788 1504
rect 972 1496 980 1504
rect 1276 1496 1284 1504
rect 1292 1496 1300 1504
rect 1708 1496 1716 1504
rect 1724 1496 1732 1504
rect 1980 1496 1988 1504
rect 2092 1496 2100 1504
rect 12 1476 20 1484
rect 108 1476 116 1484
rect 300 1476 308 1484
rect 588 1476 596 1484
rect 636 1480 644 1488
rect 668 1476 676 1484
rect 860 1476 868 1484
rect 1084 1476 1092 1484
rect 1372 1476 1380 1484
rect 1692 1476 1700 1484
rect 1788 1476 1796 1484
rect 1980 1476 1988 1484
rect 2252 1476 2260 1484
rect 92 1456 100 1464
rect 332 1456 340 1464
rect 668 1456 676 1464
rect 892 1456 900 1464
rect 1196 1456 1204 1464
rect 1404 1456 1412 1464
rect 1580 1456 1588 1464
rect 1836 1456 1844 1464
rect 2012 1456 2020 1464
rect 2172 1456 2180 1464
rect 540 1436 548 1444
rect 684 1436 692 1444
rect 1628 1436 1636 1444
rect 876 1406 884 1414
rect 1868 1406 1876 1414
rect 444 1376 452 1384
rect 636 1376 644 1384
rect 700 1376 708 1384
rect 1372 1376 1380 1384
rect 1452 1376 1460 1384
rect 1644 1376 1652 1384
rect 76 1356 84 1364
rect 156 1356 164 1364
rect 252 1356 260 1364
rect 396 1356 404 1364
rect 620 1356 628 1364
rect 860 1356 868 1364
rect 1468 1356 1476 1364
rect 1500 1356 1508 1364
rect 1628 1356 1636 1364
rect 1708 1356 1716 1364
rect 1724 1356 1732 1364
rect 1788 1356 1796 1364
rect 1820 1356 1828 1364
rect 1996 1356 2004 1364
rect 60 1336 68 1344
rect 124 1336 132 1344
rect 220 1336 228 1344
rect 300 1336 308 1344
rect 892 1336 900 1344
rect 1052 1336 1060 1344
rect 1180 1336 1188 1344
rect 1436 1336 1444 1344
rect 1468 1336 1476 1344
rect 1500 1336 1508 1344
rect 1564 1336 1572 1344
rect 1580 1336 1588 1344
rect 1692 1336 1700 1344
rect 1740 1336 1748 1344
rect 2028 1336 2036 1344
rect 28 1316 36 1324
rect 44 1316 52 1324
rect 108 1316 116 1324
rect 172 1316 180 1324
rect 236 1316 244 1324
rect 300 1316 308 1324
rect 428 1316 436 1324
rect 460 1316 468 1324
rect 492 1316 500 1324
rect 556 1316 564 1324
rect 668 1316 676 1324
rect 780 1316 788 1324
rect 1340 1316 1348 1324
rect 1420 1316 1428 1324
rect 1548 1316 1556 1324
rect 1676 1316 1684 1324
rect 1756 1316 1764 1324
rect 2028 1316 2036 1324
rect 2092 1316 2100 1324
rect 2172 1316 2180 1324
rect 12 1296 20 1304
rect 476 1296 484 1304
rect 540 1296 548 1304
rect 988 1296 996 1304
rect 1516 1296 1524 1304
rect 1644 1296 1652 1304
rect 2124 1296 2132 1304
rect 508 1276 516 1284
rect 556 1276 564 1284
rect 604 1276 612 1284
rect 2252 1276 2260 1284
rect 188 1236 196 1244
rect 348 1236 356 1244
rect 492 1236 500 1244
rect 556 1236 564 1244
rect 988 1236 996 1244
rect 1308 1236 1316 1244
rect 2124 1236 2132 1244
rect 412 1206 420 1214
rect 1340 1206 1348 1214
rect 76 1176 84 1184
rect 364 1176 372 1184
rect 444 1176 452 1184
rect 716 1176 724 1184
rect 828 1176 836 1184
rect 1260 1176 1268 1184
rect 1836 1176 1844 1184
rect 1436 1158 1444 1166
rect 652 1136 660 1144
rect 668 1136 676 1144
rect 732 1136 740 1144
rect 940 1136 948 1144
rect 364 1116 372 1124
rect 588 1116 596 1124
rect 684 1116 692 1124
rect 700 1116 708 1124
rect 1436 1112 1444 1120
rect 1836 1116 1844 1124
rect 364 1096 372 1104
rect 460 1096 468 1104
rect 524 1096 532 1104
rect 668 1096 676 1104
rect 716 1096 724 1104
rect 764 1096 772 1104
rect 860 1096 868 1104
rect 1020 1096 1028 1104
rect 1068 1096 1076 1104
rect 1148 1096 1156 1104
rect 1196 1096 1204 1104
rect 1212 1096 1220 1104
rect 1228 1096 1236 1104
rect 1276 1096 1284 1104
rect 1404 1096 1412 1104
rect 1612 1096 1620 1104
rect 1772 1096 1780 1104
rect 1836 1096 1844 1104
rect 2044 1096 2052 1104
rect 2188 1096 2196 1104
rect 12 1076 20 1084
rect 268 1076 276 1084
rect 476 1076 484 1084
rect 620 1076 628 1084
rect 764 1076 772 1084
rect 956 1076 964 1084
rect 1052 1076 1060 1084
rect 1132 1076 1140 1084
rect 1500 1076 1508 1084
rect 1756 1076 1764 1084
rect 1932 1076 1940 1084
rect 2252 1076 2260 1084
rect 236 1056 244 1064
rect 428 1056 436 1064
rect 540 1056 548 1064
rect 572 1056 580 1064
rect 1036 1056 1044 1064
rect 1532 1056 1540 1064
rect 1724 1056 1732 1064
rect 1740 1056 1748 1064
rect 1964 1056 1972 1064
rect 2124 1056 2132 1064
rect 2172 1056 2180 1064
rect 492 1036 500 1044
rect 652 1036 660 1044
rect 780 1036 788 1044
rect 988 1036 996 1044
rect 1180 1036 1188 1044
rect 1324 1036 1332 1044
rect 1692 1036 1700 1044
rect 2156 1036 2164 1044
rect 876 1006 884 1014
rect 1868 1006 1876 1014
rect 1036 976 1044 984
rect 1532 976 1540 984
rect 1724 976 1732 984
rect 1788 976 1796 984
rect 12 956 20 964
rect 252 956 260 964
rect 780 956 788 964
rect 1196 956 1204 964
rect 1452 956 1460 964
rect 1548 956 1556 964
rect 1980 956 1988 964
rect 2204 956 2212 964
rect 92 936 100 944
rect 284 936 292 944
rect 412 936 420 944
rect 476 936 484 944
rect 524 936 532 944
rect 540 936 548 944
rect 812 936 820 944
rect 1228 936 1236 944
rect 1404 936 1412 944
rect 1452 936 1460 944
rect 1484 936 1492 944
rect 1564 936 1572 944
rect 1676 936 1684 944
rect 1740 936 1748 944
rect 1948 936 1956 944
rect 60 916 68 924
rect 76 916 84 924
rect 124 916 132 924
rect 204 916 212 924
rect 252 916 260 924
rect 316 916 324 924
rect 428 916 436 924
rect 108 896 116 904
rect 220 896 228 904
rect 348 896 356 904
rect 396 896 404 904
rect 460 896 468 904
rect 508 916 516 924
rect 556 916 564 924
rect 604 916 612 924
rect 892 916 900 924
rect 1116 916 1124 924
rect 1308 916 1316 924
rect 1436 916 1444 924
rect 1500 916 1508 924
rect 1516 916 1524 924
rect 1660 916 1668 924
rect 1756 916 1764 924
rect 1852 916 1860 924
rect 2172 916 2180 924
rect 2188 916 2196 924
rect 2236 916 2244 924
rect 908 896 916 904
rect 1292 900 1300 908
rect 1388 896 1396 904
rect 1596 896 1604 904
rect 1724 896 1732 904
rect 1788 896 1796 904
rect 1884 900 1892 908
rect 140 876 148 884
rect 172 876 180 884
rect 252 876 260 884
rect 1452 876 1460 884
rect 156 856 164 864
rect 1292 854 1300 862
rect 1884 854 1892 862
rect 620 836 628 844
rect 908 836 916 844
rect 972 836 980 844
rect 2140 836 2148 844
rect 412 806 420 814
rect 1340 806 1348 814
rect 124 776 132 784
rect 412 776 420 784
rect 588 776 596 784
rect 1292 776 1300 784
rect 60 736 68 744
rect 524 736 532 744
rect 956 758 964 766
rect 1676 758 1684 766
rect 668 736 676 744
rect 1212 736 1220 744
rect 2252 736 2260 744
rect 412 716 420 724
rect 556 716 564 724
rect 572 716 580 724
rect 604 716 612 724
rect 636 716 644 724
rect 748 716 756 724
rect 44 696 52 704
rect 92 696 100 704
rect 380 696 388 704
rect 492 696 500 704
rect 540 696 548 704
rect 588 696 596 704
rect 668 696 676 704
rect 828 716 836 724
rect 956 712 964 720
rect 1292 716 1300 724
rect 1676 712 1684 720
rect 812 696 820 704
rect 860 696 868 704
rect 924 696 932 704
rect 940 696 948 704
rect 1308 696 1316 704
rect 1500 696 1508 704
rect 1644 696 1652 704
rect 1852 696 1860 704
rect 2108 696 2116 704
rect 2124 696 2132 704
rect 2172 696 2180 704
rect 12 676 20 684
rect 316 676 324 684
rect 684 676 692 684
rect 700 676 708 684
rect 796 676 804 684
rect 1020 676 1028 684
rect 1388 676 1396 684
rect 1740 676 1748 684
rect 2028 676 2036 684
rect 284 656 292 664
rect 476 656 484 664
rect 1052 656 1060 664
rect 1420 656 1428 664
rect 1772 656 1780 664
rect 1980 656 1988 664
rect 2044 656 2052 664
rect 2156 676 2164 684
rect 2076 656 2084 664
rect 1580 636 1588 644
rect 876 606 884 614
rect 1868 606 1876 614
rect 1212 576 1220 584
rect 1692 576 1700 584
rect 2236 576 2244 584
rect 76 556 84 564
rect 236 556 244 564
rect 412 556 420 564
rect 460 556 468 564
rect 540 556 548 564
rect 636 556 644 564
rect 828 556 836 564
rect 1020 556 1028 564
rect 1036 556 1044 564
rect 1452 556 1460 564
rect 1628 556 1636 564
rect 2028 556 2036 564
rect 2204 556 2212 564
rect 268 536 276 544
rect 460 536 468 544
rect 492 536 500 544
rect 860 536 868 544
rect 1052 536 1060 544
rect 1484 536 1492 544
rect 1772 536 1780 544
rect 1788 536 1796 544
rect 1996 536 2004 544
rect 348 516 356 524
rect 380 516 388 524
rect 460 516 468 524
rect 508 516 516 524
rect 572 516 580 524
rect 666 516 674 524
rect 940 516 948 524
rect 1228 516 1236 524
rect 1372 516 1380 524
rect 1596 516 1604 524
rect 1660 516 1668 524
rect 1756 516 1764 524
rect 1932 516 1940 524
rect 332 500 340 508
rect 540 496 548 504
rect 924 500 932 508
rect 1228 496 1236 504
rect 1548 500 1556 508
rect 1724 496 1732 504
rect 1836 496 1844 504
rect 1900 496 1908 504
rect 12 476 20 484
rect 588 476 596 484
rect 620 476 628 484
rect 1244 476 1252 484
rect 572 456 580 464
rect 1548 454 1556 462
rect 332 436 340 444
rect 524 436 532 444
rect 924 436 932 444
rect 1164 436 1172 444
rect 1228 436 1236 444
rect 1644 436 1652 444
rect 1804 436 1812 444
rect 1900 436 1908 444
rect 2188 436 2196 444
rect 412 406 420 414
rect 1340 406 1348 414
rect 28 376 36 384
rect 1148 376 1156 384
rect 1916 376 1924 384
rect 2124 376 2132 384
rect 220 356 228 364
rect 812 358 820 366
rect 1052 336 1060 344
rect 1612 336 1620 344
rect 316 316 324 324
rect 524 316 532 324
rect 812 312 820 320
rect 1148 316 1156 324
rect 1916 316 1924 324
rect 220 296 228 304
rect 364 296 372 304
rect 412 296 420 304
rect 492 296 500 304
rect 554 296 562 304
rect 844 296 852 304
rect 956 296 964 304
rect 1148 296 1156 304
rect 1356 296 1364 304
rect 1580 296 1588 304
rect 1596 296 1604 304
rect 1708 296 1716 304
rect 1900 296 1908 304
rect 1932 296 1940 304
rect 2028 296 2036 304
rect 2076 296 2084 304
rect 2092 296 2100 304
rect 2188 296 2196 304
rect 220 276 228 284
rect 428 276 436 284
rect 524 276 532 284
rect 748 276 756 284
rect 892 276 900 284
rect 1020 276 1028 284
rect 1244 276 1252 284
rect 1516 276 1524 284
rect 1820 276 1828 284
rect 1964 276 1972 284
rect 2060 276 2068 284
rect 2252 276 2260 284
rect 188 256 196 264
rect 444 256 452 264
rect 716 256 724 264
rect 1276 256 1284 264
rect 1484 256 1492 264
rect 1788 256 1796 264
rect 1980 256 1988 264
rect 2060 256 2068 264
rect 2188 256 2196 264
rect 1004 236 1012 244
rect 1628 236 1636 244
rect 876 206 884 214
rect 1868 206 1876 214
rect 1676 176 1684 184
rect 2156 176 2164 184
rect 28 156 36 164
rect 188 156 196 164
rect 364 156 372 164
rect 412 156 420 164
rect 444 156 452 164
rect 636 156 644 164
rect 1132 156 1140 164
rect 1388 156 1396 164
rect 1580 156 1588 164
rect 1692 156 1700 164
rect 1756 156 1764 164
rect 1996 156 2004 164
rect 220 136 228 144
rect 668 136 676 144
rect 828 136 836 144
rect 956 136 964 144
rect 1100 136 1108 144
rect 1420 136 1428 144
rect 1660 136 1668 144
rect 1804 136 1812 144
rect 1964 136 1972 144
rect 316 116 324 124
rect 556 116 564 124
rect 764 116 772 124
rect 1004 116 1012 124
rect 1324 116 1332 124
rect 1484 116 1492 124
rect 1500 116 1508 124
rect 1516 116 1524 124
rect 1564 116 1572 124
rect 1580 116 1588 124
rect 1644 116 1652 124
rect 1708 116 1716 124
rect 1788 116 1796 124
rect 1900 116 1908 124
rect 284 100 292 108
rect 732 100 740 108
rect 1036 100 1044 108
rect 1756 96 1764 104
rect 1868 96 1876 104
rect 2252 76 2260 84
rect 732 54 740 62
rect 1036 54 1044 62
rect 284 36 292 44
rect 1372 36 1380 44
rect 1548 36 1556 44
rect 1628 36 1636 44
rect 1740 36 1748 44
rect 1868 36 1876 44
rect 412 6 420 14
rect 1340 6 1348 14
<< metal2 >>
rect 408 2006 412 2014
rect 420 2006 424 2014
rect 445 1944 451 2043
rect 125 1904 131 1916
rect 13 1744 19 1876
rect 29 1804 35 1896
rect 77 1884 83 1896
rect 333 1884 339 1916
rect 365 1904 371 1916
rect 445 1904 451 1936
rect 557 1884 563 2043
rect 605 1903 611 1916
rect 621 1904 627 2043
rect 605 1897 620 1903
rect 237 1864 243 1876
rect 333 1864 339 1876
rect 429 1864 435 1876
rect 509 1864 515 1876
rect 29 1724 35 1796
rect 77 1744 83 1776
rect 141 1764 147 1836
rect 221 1784 227 1836
rect 381 1804 387 1836
rect 125 1584 131 1696
rect 13 1484 19 1496
rect 45 1363 51 1496
rect 125 1484 131 1496
rect 93 1364 99 1456
rect 45 1357 60 1363
rect 61 1344 67 1356
rect 45 1324 51 1336
rect 13 1184 19 1296
rect 77 1184 83 1356
rect 109 1324 115 1476
rect 141 1364 147 1676
rect 205 1524 211 1576
rect 125 1304 131 1336
rect 157 1284 163 1356
rect 221 1344 227 1756
rect 237 1504 243 1716
rect 317 1643 323 1756
rect 445 1724 451 1836
rect 525 1764 531 1836
rect 541 1724 547 1796
rect 557 1763 563 1876
rect 653 1864 659 2043
rect 765 2037 787 2043
rect 1101 2037 1123 2043
rect 1229 2037 1251 2043
rect 1533 2037 1555 2043
rect 765 1984 771 2037
rect 1101 1984 1107 2037
rect 733 1917 748 1923
rect 589 1844 595 1856
rect 573 1784 579 1836
rect 589 1764 595 1796
rect 557 1757 579 1763
rect 573 1744 579 1757
rect 445 1644 451 1696
rect 525 1684 531 1716
rect 557 1704 563 1736
rect 589 1724 595 1756
rect 621 1704 627 1776
rect 653 1764 659 1856
rect 717 1804 723 1896
rect 733 1744 739 1917
rect 797 1864 803 1896
rect 877 1864 883 1916
rect 749 1744 755 1856
rect 872 1806 876 1814
rect 884 1806 888 1814
rect 925 1744 931 1856
rect 957 1844 963 1856
rect 957 1744 963 1836
rect 1005 1744 1011 1896
rect 1053 1864 1059 1876
rect 1085 1764 1091 1856
rect 1245 1784 1251 2037
rect 1336 2006 1340 2014
rect 1348 2006 1352 2014
rect 1549 1984 1555 2037
rect 1565 2037 1587 2043
rect 1565 1984 1571 2037
rect 1837 2004 1843 2043
rect 1997 2037 2019 2043
rect 2013 1984 2019 2037
rect 1453 1924 1459 1976
rect 1677 1920 1683 1958
rect 1357 1884 1363 1896
rect 317 1637 339 1643
rect 301 1484 307 1536
rect 333 1464 339 1637
rect 408 1606 412 1614
rect 420 1606 424 1614
rect 541 1524 547 1636
rect 589 1484 595 1696
rect 637 1544 643 1736
rect 621 1480 636 1483
rect 621 1477 643 1480
rect 237 1284 243 1316
rect 13 1084 19 1096
rect 13 944 19 956
rect 77 924 83 956
rect 93 904 99 936
rect 109 904 115 996
rect 141 903 147 1056
rect 157 1004 163 1276
rect 189 1204 195 1236
rect 253 1184 259 1356
rect 301 1344 307 1356
rect 301 1244 307 1316
rect 269 1084 275 1196
rect 333 1084 339 1456
rect 445 1384 451 1476
rect 541 1384 547 1436
rect 461 1284 467 1316
rect 557 1264 563 1276
rect 589 1263 595 1476
rect 621 1364 627 1477
rect 685 1483 691 1716
rect 676 1477 691 1483
rect 637 1384 643 1396
rect 621 1344 627 1356
rect 621 1304 627 1336
rect 669 1324 675 1456
rect 589 1257 611 1263
rect 349 1164 355 1236
rect 408 1206 412 1214
rect 420 1206 424 1214
rect 445 1184 451 1256
rect 365 1124 371 1176
rect 461 1104 467 1236
rect 237 1064 243 1076
rect 461 1064 467 1096
rect 493 1083 499 1236
rect 525 1084 531 1096
rect 484 1077 499 1083
rect 557 1063 563 1236
rect 589 1124 595 1136
rect 548 1057 563 1063
rect 205 924 211 936
rect 221 904 227 916
rect 285 904 291 936
rect 317 924 323 936
rect 349 904 355 996
rect 413 924 419 936
rect 125 897 147 903
rect 13 684 19 696
rect 93 664 99 696
rect 13 484 19 496
rect 109 384 115 896
rect 125 784 131 897
rect 429 884 435 916
rect 408 806 412 814
rect 420 806 424 814
rect 125 704 131 776
rect 413 724 419 776
rect 317 684 323 716
rect 285 624 291 656
rect 237 564 243 616
rect 237 424 243 556
rect 269 524 275 536
rect 381 524 387 696
rect 461 564 467 756
rect 477 724 483 936
rect 493 923 499 1036
rect 525 944 531 996
rect 493 917 508 923
rect 525 764 531 936
rect 557 864 563 916
rect 573 744 579 1056
rect 605 1004 611 1257
rect 653 1144 659 1156
rect 669 1104 675 1136
rect 685 1124 691 1436
rect 701 1384 707 1696
rect 749 1684 755 1736
rect 765 1724 771 1736
rect 925 1704 931 1736
rect 1197 1723 1203 1756
rect 1325 1724 1331 1856
rect 1405 1744 1411 1776
rect 1437 1724 1443 1756
rect 1197 1717 1212 1723
rect 1293 1717 1308 1723
rect 1053 1704 1059 1716
rect 1133 1704 1139 1716
rect 717 1564 723 1676
rect 717 1504 723 1556
rect 765 1524 771 1696
rect 941 1604 947 1636
rect 797 1520 803 1558
rect 717 1184 723 1296
rect 685 1104 691 1116
rect 621 1084 627 1096
rect 701 1084 707 1116
rect 765 1104 771 1516
rect 781 1324 787 1496
rect 861 1484 867 1596
rect 1053 1584 1059 1696
rect 973 1484 979 1496
rect 872 1406 876 1414
rect 884 1406 888 1414
rect 893 1344 899 1376
rect 1053 1344 1059 1356
rect 781 1224 787 1316
rect 989 1244 995 1296
rect 829 1184 835 1216
rect 1069 1144 1075 1636
rect 1085 1444 1091 1476
rect 1165 1384 1171 1716
rect 1213 1704 1219 1716
rect 1277 1524 1283 1576
rect 1293 1504 1299 1717
rect 1309 1644 1315 1696
rect 1336 1606 1340 1614
rect 1348 1606 1352 1614
rect 1181 1344 1187 1436
rect 941 1124 947 1136
rect 1021 1104 1027 1116
rect 1133 1084 1139 1096
rect 1149 1084 1155 1096
rect 589 784 595 936
rect 605 924 611 936
rect 573 684 579 716
rect 589 704 595 736
rect 605 564 611 716
rect 621 703 627 836
rect 637 704 643 716
rect 621 697 636 703
rect 621 664 627 697
rect 653 703 659 1036
rect 653 697 668 703
rect 685 684 691 796
rect 701 724 707 1076
rect 765 1004 771 1076
rect 1181 1064 1187 1336
rect 1197 1104 1203 1336
rect 1213 1104 1219 1496
rect 1277 1484 1283 1496
rect 1373 1424 1379 1476
rect 1405 1464 1411 1716
rect 1453 1384 1459 1416
rect 1517 1364 1523 1896
rect 1597 1744 1603 1896
rect 1741 1823 1747 1876
rect 1853 1864 1859 1896
rect 2109 1883 2115 2043
rect 2109 1877 2131 1883
rect 1741 1817 1763 1823
rect 1693 1744 1699 1756
rect 1677 1584 1683 1716
rect 1693 1484 1699 1736
rect 1725 1724 1731 1816
rect 1757 1784 1763 1817
rect 1773 1764 1779 1856
rect 1933 1824 1939 1836
rect 1864 1806 1868 1814
rect 1876 1806 1880 1814
rect 1901 1764 1907 1816
rect 1741 1724 1747 1736
rect 1773 1724 1779 1756
rect 1981 1724 1987 1856
rect 2061 1844 2067 1876
rect 2125 1864 2131 1877
rect 2157 1864 2163 1896
rect 2253 1884 2259 1896
rect 2045 1744 2051 1836
rect 2157 1784 2163 1856
rect 1709 1717 1724 1723
rect 1709 1504 1715 1717
rect 1732 1497 1747 1503
rect 1581 1364 1587 1456
rect 1645 1384 1651 1416
rect 1476 1357 1491 1363
rect 1485 1343 1491 1357
rect 1581 1344 1587 1356
rect 1485 1337 1500 1343
rect 1565 1324 1571 1336
rect 1677 1324 1683 1376
rect 1741 1344 1747 1497
rect 1821 1364 1827 1716
rect 1949 1644 1955 1696
rect 1917 1520 1923 1558
rect 1981 1504 1987 1716
rect 2077 1604 2083 1756
rect 2013 1464 2019 1596
rect 1864 1406 1868 1414
rect 1876 1406 1880 1414
rect 2013 1403 2019 1456
rect 1997 1397 2019 1403
rect 1997 1364 2003 1397
rect 1789 1344 1795 1356
rect 2029 1344 2035 1356
rect 2093 1324 2099 1496
rect 2253 1484 2259 1496
rect 1261 1184 1267 1276
rect 1277 1124 1283 1316
rect 1421 1284 1427 1316
rect 1549 1284 1555 1316
rect 1229 1104 1235 1116
rect 1277 1104 1283 1116
rect 781 984 787 1036
rect 872 1006 876 1014
rect 884 1006 888 1014
rect 701 684 707 696
rect 797 684 803 816
rect 893 724 899 916
rect 909 844 915 896
rect 973 824 979 836
rect 989 804 995 1036
rect 1037 984 1043 1056
rect 1213 1044 1219 1096
rect 1309 1064 1315 1236
rect 1336 1206 1340 1214
rect 1348 1206 1352 1214
rect 1437 1120 1443 1158
rect 1181 1004 1187 1036
rect 957 720 963 758
rect 925 704 931 716
rect 813 684 819 696
rect 541 524 547 556
rect 573 524 579 536
rect 333 444 339 500
rect 349 424 355 516
rect 509 484 515 516
rect 541 504 547 516
rect 637 504 643 556
rect 685 544 691 676
rect 797 644 803 676
rect 872 606 876 614
rect 884 606 888 614
rect 573 464 579 476
rect 189 264 195 416
rect 221 304 227 356
rect 317 324 323 416
rect 408 406 412 414
rect 420 406 424 414
rect 525 324 531 436
rect 813 320 819 358
rect 189 164 195 256
rect 317 124 323 316
rect 365 284 371 296
rect 413 277 428 283
rect 413 164 419 277
rect 445 264 451 296
rect 493 284 499 296
rect 829 264 835 556
rect 861 504 867 536
rect 941 524 947 696
rect 1053 664 1059 956
rect 1229 944 1235 996
rect 1309 964 1315 1056
rect 1293 862 1299 900
rect 1053 544 1059 616
rect 1213 584 1219 676
rect 1229 584 1235 636
rect 1037 537 1052 543
rect 925 444 931 500
rect 637 164 643 256
rect 445 144 451 156
rect 829 144 835 256
rect 285 44 291 100
rect 669 24 675 136
rect 845 124 851 296
rect 893 284 899 296
rect 1005 244 1011 276
rect 872 206 876 214
rect 884 206 888 214
rect 957 144 963 156
rect 733 62 739 100
rect 408 6 412 14
rect 420 6 424 14
rect 621 -23 627 16
rect 957 -17 963 136
rect 1005 124 1011 236
rect 941 -23 963 -17
rect 989 -23 995 36
rect 1021 24 1027 276
rect 1037 164 1043 537
rect 1229 524 1235 576
rect 1245 504 1251 796
rect 1293 724 1299 776
rect 1309 704 1315 916
rect 1325 844 1331 1036
rect 1405 944 1411 956
rect 1389 904 1395 936
rect 1336 806 1340 814
rect 1348 806 1352 814
rect 1389 744 1395 896
rect 1421 684 1427 1056
rect 1501 1044 1507 1076
rect 1533 984 1539 1036
rect 1645 1004 1651 1296
rect 1757 1284 1763 1316
rect 1764 1277 1779 1283
rect 1773 1104 1779 1277
rect 2029 1243 2035 1316
rect 2125 1244 2131 1296
rect 2029 1237 2051 1243
rect 1837 1124 1843 1176
rect 2045 1104 2051 1237
rect 1933 1064 1939 1076
rect 1549 964 1555 976
rect 1565 944 1571 956
rect 1453 924 1459 936
rect 1437 904 1443 916
rect 1485 904 1491 936
rect 1677 924 1683 936
rect 1517 884 1523 916
rect 1389 624 1395 676
rect 1421 664 1427 676
rect 1245 484 1251 496
rect 1053 304 1059 336
rect 1149 324 1155 376
rect 1149 284 1155 296
rect 1165 264 1171 436
rect 1229 384 1235 436
rect 1336 406 1340 414
rect 1348 406 1352 414
rect 1373 383 1379 516
rect 1357 377 1379 383
rect 1357 304 1363 377
rect 1453 264 1459 556
rect 1485 544 1491 556
rect 1549 462 1555 500
rect 1597 404 1603 516
rect 1133 164 1139 256
rect 1389 124 1395 156
rect 1485 144 1491 256
rect 1501 124 1507 376
rect 1581 304 1587 316
rect 1597 304 1603 376
rect 1613 344 1619 916
rect 1629 564 1635 636
rect 1629 544 1635 556
rect 1661 524 1667 916
rect 1693 844 1699 1036
rect 1725 984 1731 1056
rect 1965 1023 1971 1056
rect 1965 1017 1987 1023
rect 1864 1006 1868 1014
rect 1876 1006 1880 1014
rect 1981 964 1987 1017
rect 1725 864 1731 896
rect 1757 844 1763 916
rect 1677 720 1683 758
rect 1773 684 1779 876
rect 1789 864 1795 896
rect 1853 704 1859 916
rect 1885 862 1891 900
rect 1981 884 1987 956
rect 1741 664 1747 676
rect 1773 664 1779 676
rect 1981 664 1987 696
rect 2077 664 2083 1096
rect 2157 1044 2163 1076
rect 2173 1064 2179 1316
rect 2253 1284 2259 1296
rect 2253 1084 2259 1096
rect 2157 924 2163 1036
rect 2205 944 2211 956
rect 2173 844 2179 916
rect 2109 704 2115 836
rect 2109 684 2115 696
rect 2141 684 2147 836
rect 2157 684 2163 696
rect 2173 684 2179 696
rect 2077 644 2083 656
rect 1693 584 1699 616
rect 1629 263 1635 516
rect 1661 504 1667 516
rect 1645 324 1651 436
rect 1629 257 1651 263
rect 1581 164 1587 236
rect 1517 124 1523 136
rect 1581 124 1587 156
rect 1645 124 1651 257
rect 1677 184 1683 276
rect 1693 203 1699 536
rect 1725 504 1731 576
rect 1773 544 1779 636
rect 1864 606 1868 614
rect 1876 606 1880 614
rect 1837 504 1843 576
rect 1901 444 1907 496
rect 1709 304 1715 396
rect 1805 384 1811 436
rect 1917 324 1923 376
rect 1933 304 1939 516
rect 2029 404 2035 556
rect 1693 197 1715 203
rect 1709 124 1715 197
rect 1757 104 1763 136
rect 1789 124 1795 236
rect 1864 206 1868 214
rect 1876 206 1880 214
rect 1805 144 1811 176
rect 1901 124 1907 296
rect 1965 144 1971 276
rect 1981 264 1987 376
rect 1997 264 2003 396
rect 2109 304 2115 676
rect 2205 564 2211 676
rect 2237 584 2243 916
rect 2125 384 2131 536
rect 2189 304 2195 436
rect 1997 164 2003 256
rect 2029 244 2035 296
rect 2093 284 2099 296
rect 2189 264 2195 296
rect 2253 284 2259 296
rect 2061 204 2067 256
rect 2157 184 2163 196
rect 1037 62 1043 100
rect 1869 44 1875 96
rect 2253 84 2259 96
rect 1069 -23 1075 16
rect 1336 6 1340 14
rect 1348 6 1352 14
rect 1373 -17 1379 36
rect 1549 -17 1555 36
rect 1629 -17 1635 36
rect 1741 -17 1747 36
rect 1357 -23 1379 -17
rect 1533 -23 1555 -17
rect 1613 -23 1635 -17
rect 1725 -23 1747 -17
<< m3contact >>
rect 412 2006 420 2014
rect 92 1936 100 1944
rect 284 1936 292 1944
rect 60 1916 68 1924
rect 76 1896 84 1904
rect 124 1896 132 1904
rect 252 1896 260 1904
rect 300 1896 308 1904
rect 12 1876 20 1884
rect 364 1896 372 1904
rect 396 1896 404 1904
rect 444 1896 452 1904
rect 620 1896 628 1904
rect 156 1876 164 1884
rect 252 1876 260 1884
rect 428 1876 436 1884
rect 492 1876 500 1884
rect 556 1876 564 1884
rect 108 1856 116 1864
rect 172 1856 180 1864
rect 236 1856 244 1864
rect 332 1856 340 1864
rect 508 1856 516 1864
rect 28 1796 36 1804
rect 76 1776 84 1784
rect 380 1796 388 1804
rect 220 1776 228 1784
rect 140 1756 148 1764
rect 220 1756 228 1764
rect 140 1736 148 1744
rect 60 1696 68 1704
rect 12 1496 20 1504
rect 60 1496 68 1504
rect 124 1476 132 1484
rect 60 1356 68 1364
rect 92 1356 100 1364
rect 44 1336 52 1344
rect 28 1316 36 1324
rect 156 1516 164 1524
rect 140 1356 148 1364
rect 124 1296 132 1304
rect 348 1736 356 1744
rect 540 1796 548 1804
rect 524 1756 532 1764
rect 684 1896 692 1904
rect 604 1856 612 1864
rect 588 1836 596 1844
rect 588 1796 596 1804
rect 572 1776 580 1784
rect 620 1776 628 1784
rect 588 1756 596 1764
rect 556 1736 564 1744
rect 444 1716 452 1724
rect 524 1716 532 1724
rect 716 1796 724 1804
rect 652 1756 660 1764
rect 828 1896 836 1904
rect 748 1876 756 1884
rect 812 1876 820 1884
rect 924 1876 932 1884
rect 956 1876 964 1884
rect 748 1856 756 1864
rect 796 1856 804 1864
rect 876 1856 884 1864
rect 924 1856 932 1864
rect 972 1856 980 1864
rect 876 1806 884 1814
rect 876 1756 884 1764
rect 956 1836 964 1844
rect 1052 1856 1060 1864
rect 1084 1856 1092 1864
rect 1148 1856 1156 1864
rect 1020 1836 1028 1844
rect 1340 2006 1348 2014
rect 1836 1996 1844 2004
rect 1356 1896 1364 1904
rect 1452 1896 1460 1904
rect 1628 1896 1636 1904
rect 2076 1896 2084 1904
rect 684 1736 692 1744
rect 732 1736 740 1744
rect 764 1736 772 1744
rect 860 1736 868 1744
rect 956 1736 964 1744
rect 1004 1736 1012 1744
rect 1036 1736 1044 1744
rect 1180 1736 1188 1744
rect 556 1696 564 1704
rect 588 1696 596 1704
rect 300 1536 308 1544
rect 412 1606 420 1614
rect 492 1556 500 1564
rect 412 1496 420 1504
rect 668 1716 676 1724
rect 636 1536 644 1544
rect 444 1476 452 1484
rect 332 1456 340 1464
rect 300 1356 308 1364
rect 172 1316 180 1324
rect 156 1276 164 1284
rect 236 1276 244 1284
rect 12 1176 20 1184
rect 76 1176 84 1184
rect 12 1096 20 1104
rect 140 1056 148 1064
rect 108 996 116 1004
rect 76 956 84 964
rect 12 936 20 944
rect 60 916 68 924
rect 124 916 132 924
rect 92 896 100 904
rect 188 1196 196 1204
rect 300 1236 308 1244
rect 268 1196 276 1204
rect 252 1176 260 1184
rect 540 1376 548 1384
rect 396 1356 404 1364
rect 428 1316 436 1324
rect 492 1316 500 1324
rect 556 1316 564 1324
rect 476 1296 484 1304
rect 540 1296 548 1304
rect 460 1276 468 1284
rect 508 1276 516 1284
rect 444 1256 452 1264
rect 556 1256 564 1264
rect 636 1396 644 1404
rect 620 1336 628 1344
rect 620 1296 628 1304
rect 604 1276 612 1284
rect 412 1206 420 1214
rect 460 1236 468 1244
rect 348 1156 356 1164
rect 364 1096 372 1104
rect 236 1076 244 1084
rect 332 1076 340 1084
rect 524 1076 532 1084
rect 428 1056 436 1064
rect 460 1056 468 1064
rect 588 1136 596 1144
rect 156 996 164 1004
rect 348 996 356 1004
rect 252 956 260 964
rect 204 936 212 944
rect 316 936 324 944
rect 220 916 228 924
rect 252 916 260 924
rect 412 916 420 924
rect 60 736 68 744
rect 12 696 20 704
rect 44 696 52 704
rect 92 656 100 664
rect 76 556 84 564
rect 12 496 20 504
rect 284 896 292 904
rect 396 896 404 904
rect 460 896 468 904
rect 140 876 148 884
rect 172 876 180 884
rect 252 876 260 884
rect 428 876 436 884
rect 156 856 164 864
rect 412 806 420 814
rect 460 756 468 764
rect 316 716 324 724
rect 124 696 132 704
rect 236 616 244 624
rect 284 616 292 624
rect 524 996 532 1004
rect 540 936 548 944
rect 556 856 564 864
rect 524 756 532 764
rect 652 1156 660 1164
rect 796 1716 804 1724
rect 1020 1716 1028 1724
rect 1084 1716 1092 1724
rect 1404 1776 1412 1784
rect 764 1696 772 1704
rect 924 1696 932 1704
rect 988 1696 996 1704
rect 1052 1696 1060 1704
rect 1132 1696 1140 1704
rect 716 1676 724 1684
rect 748 1676 756 1684
rect 716 1556 724 1564
rect 860 1596 868 1604
rect 940 1596 948 1604
rect 764 1516 772 1524
rect 716 1296 724 1304
rect 732 1136 740 1144
rect 620 1096 628 1104
rect 684 1096 692 1104
rect 780 1496 788 1504
rect 972 1476 980 1484
rect 892 1456 900 1464
rect 876 1406 884 1414
rect 892 1376 900 1384
rect 860 1356 868 1364
rect 1052 1356 1060 1364
rect 780 1216 788 1224
rect 828 1216 836 1224
rect 1084 1436 1092 1444
rect 1212 1696 1220 1704
rect 1324 1716 1332 1724
rect 1404 1716 1412 1724
rect 1436 1716 1444 1724
rect 1340 1606 1348 1614
rect 1212 1496 1220 1504
rect 1196 1456 1204 1464
rect 1180 1436 1188 1444
rect 1164 1376 1172 1384
rect 1196 1336 1204 1344
rect 1068 1136 1076 1144
rect 940 1116 948 1124
rect 1020 1116 1028 1124
rect 716 1096 724 1104
rect 860 1096 868 1104
rect 1068 1096 1076 1104
rect 1132 1096 1140 1104
rect 700 1076 708 1084
rect 956 1076 964 1084
rect 1052 1076 1060 1084
rect 1148 1076 1156 1084
rect 604 996 612 1004
rect 588 936 596 944
rect 604 936 612 944
rect 524 736 532 744
rect 572 736 580 744
rect 588 736 596 744
rect 476 716 484 724
rect 556 716 564 724
rect 492 696 500 704
rect 540 696 548 704
rect 572 676 580 684
rect 476 656 484 664
rect 636 696 644 704
rect 684 796 692 804
rect 668 736 676 744
rect 1276 1476 1284 1484
rect 1404 1456 1412 1464
rect 1372 1416 1380 1424
rect 1452 1416 1460 1424
rect 1372 1376 1380 1384
rect 1724 1816 1732 1824
rect 2124 1896 2132 1904
rect 2252 1896 2260 1904
rect 1852 1856 1860 1864
rect 1980 1856 1988 1864
rect 2028 1856 2036 1864
rect 1644 1776 1652 1784
rect 1628 1756 1636 1764
rect 1596 1736 1598 1744
rect 1598 1736 1604 1744
rect 1692 1736 1700 1744
rect 1708 1736 1716 1744
rect 1676 1576 1684 1584
rect 1900 1816 1908 1824
rect 1932 1816 1940 1824
rect 1868 1806 1876 1814
rect 1852 1776 1860 1784
rect 1772 1756 1780 1764
rect 1740 1736 1748 1744
rect 2092 1856 2100 1864
rect 2060 1836 2068 1844
rect 2156 1776 2164 1784
rect 2236 1776 2244 1784
rect 2076 1756 2084 1764
rect 1772 1716 1780 1724
rect 1788 1716 1796 1724
rect 1868 1716 1876 1724
rect 1708 1496 1716 1504
rect 1628 1436 1636 1444
rect 1644 1416 1652 1424
rect 1676 1376 1684 1384
rect 1436 1336 1444 1344
rect 1468 1336 1476 1344
rect 1500 1356 1508 1364
rect 1516 1356 1524 1364
rect 1580 1356 1588 1364
rect 1628 1356 1636 1364
rect 1708 1356 1716 1364
rect 1724 1356 1732 1364
rect 1788 1476 1796 1484
rect 2012 1596 2020 1604
rect 2076 1596 2084 1604
rect 1980 1476 1988 1484
rect 2252 1496 2260 1504
rect 1836 1456 1844 1464
rect 1868 1406 1876 1414
rect 2028 1356 2036 1364
rect 1692 1336 1700 1344
rect 1788 1336 1796 1344
rect 2172 1456 2180 1464
rect 1276 1316 1284 1324
rect 1340 1316 1348 1324
rect 1564 1316 1572 1324
rect 2172 1316 2180 1324
rect 1260 1276 1268 1284
rect 1516 1296 1524 1304
rect 1644 1296 1652 1304
rect 1420 1276 1428 1284
rect 1548 1276 1556 1284
rect 1228 1116 1236 1124
rect 1276 1116 1284 1124
rect 1180 1056 1188 1064
rect 764 996 772 1004
rect 876 1006 884 1014
rect 780 976 788 984
rect 780 956 788 964
rect 812 936 820 944
rect 892 916 900 924
rect 796 816 804 824
rect 700 716 708 724
rect 748 716 756 724
rect 700 696 708 704
rect 972 816 980 824
rect 1340 1206 1348 1214
rect 1404 1096 1412 1104
rect 1612 1096 1620 1104
rect 1308 1056 1316 1064
rect 1420 1056 1428 1064
rect 1212 1036 1220 1044
rect 1180 996 1188 1004
rect 1228 996 1236 1004
rect 1052 956 1060 964
rect 1196 956 1204 964
rect 988 796 996 804
rect 828 716 836 724
rect 892 716 900 724
rect 924 716 932 724
rect 860 696 868 704
rect 796 676 804 684
rect 812 676 820 684
rect 620 656 628 664
rect 412 556 420 564
rect 604 556 612 564
rect 460 536 468 544
rect 492 536 500 544
rect 572 536 580 544
rect 268 516 276 524
rect 460 516 468 524
rect 540 516 548 524
rect 796 636 804 644
rect 876 606 884 614
rect 684 536 692 544
rect 668 516 674 524
rect 674 516 676 524
rect 636 496 644 504
rect 508 476 516 484
rect 572 476 580 484
rect 588 476 596 484
rect 620 476 628 484
rect 188 416 196 424
rect 236 416 244 424
rect 316 416 324 424
rect 348 416 356 424
rect 28 376 36 384
rect 108 376 116 384
rect 412 406 420 414
rect 220 276 228 284
rect 188 256 196 264
rect 28 156 36 164
rect 220 136 228 144
rect 412 296 420 304
rect 444 296 452 304
rect 556 296 562 304
rect 562 296 564 304
rect 364 276 372 284
rect 428 276 436 284
rect 492 276 500 284
rect 524 276 532 284
rect 748 276 756 284
rect 1020 676 1028 684
rect 1308 956 1316 964
rect 1116 916 1124 924
rect 1244 796 1252 804
rect 1212 736 1220 744
rect 1212 676 1220 684
rect 1052 616 1060 624
rect 1020 556 1028 564
rect 1036 556 1044 564
rect 1228 636 1236 644
rect 1228 576 1236 584
rect 860 496 868 504
rect 844 296 852 304
rect 892 296 900 304
rect 956 296 964 304
rect 636 256 644 264
rect 716 256 724 264
rect 828 256 836 264
rect 364 156 372 164
rect 444 136 452 144
rect 316 116 324 124
rect 556 116 564 124
rect 1004 276 1012 284
rect 876 206 884 214
rect 956 156 964 164
rect 764 116 772 124
rect 844 116 852 124
rect 620 16 628 24
rect 668 16 676 24
rect 412 6 420 14
rect 988 36 996 44
rect 1404 956 1412 964
rect 1388 936 1396 944
rect 1324 836 1332 844
rect 1340 806 1348 814
rect 1388 736 1396 744
rect 1532 1056 1540 1064
rect 1500 1036 1508 1044
rect 1532 1036 1540 1044
rect 1756 1276 1764 1284
rect 1836 1096 1844 1104
rect 2076 1096 2084 1104
rect 1756 1076 1764 1084
rect 1740 1056 1748 1064
rect 1932 1056 1940 1064
rect 1644 996 1652 1004
rect 1548 976 1556 984
rect 1452 956 1460 964
rect 1564 956 1572 964
rect 1452 916 1460 924
rect 1500 916 1508 924
rect 1612 916 1620 924
rect 1676 916 1684 924
rect 1436 896 1444 904
rect 1484 896 1492 904
rect 1596 896 1604 904
rect 1452 876 1460 884
rect 1516 876 1524 884
rect 1500 696 1508 704
rect 1420 676 1428 684
rect 1580 636 1588 644
rect 1388 616 1396 624
rect 1484 556 1492 564
rect 1228 496 1236 504
rect 1244 496 1252 504
rect 1052 296 1060 304
rect 1148 276 1156 284
rect 1340 406 1348 414
rect 1228 376 1236 384
rect 1244 276 1252 284
rect 1596 396 1604 404
rect 1500 376 1508 384
rect 1596 376 1604 384
rect 1132 256 1140 264
rect 1164 256 1172 264
rect 1276 256 1284 264
rect 1452 256 1460 264
rect 1036 156 1044 164
rect 1100 136 1108 144
rect 1420 136 1428 144
rect 1484 136 1492 144
rect 1580 316 1588 324
rect 1644 696 1652 704
rect 1628 636 1636 644
rect 1628 536 1636 544
rect 1868 1006 1876 1014
rect 1788 976 1796 984
rect 1740 936 1748 944
rect 1948 936 1956 944
rect 1724 856 1732 864
rect 1772 876 1780 884
rect 1692 836 1700 844
rect 1756 836 1764 844
rect 1788 856 1796 864
rect 1980 876 1988 884
rect 1980 696 1988 704
rect 1772 676 1780 684
rect 2028 676 2036 684
rect 2156 1076 2164 1084
rect 2124 1056 2132 1064
rect 2252 1296 2260 1304
rect 2188 1096 2196 1104
rect 2252 1096 2260 1104
rect 2172 1056 2180 1064
rect 2204 936 2212 944
rect 2156 916 2164 924
rect 2188 916 2196 924
rect 2108 836 2116 844
rect 2172 836 2180 844
rect 2124 696 2132 704
rect 2156 696 2164 704
rect 2108 676 2116 684
rect 2140 676 2148 684
rect 2172 676 2180 684
rect 2204 676 2212 684
rect 1740 656 1748 664
rect 2044 656 2052 664
rect 1772 636 1780 644
rect 2076 636 2084 644
rect 1692 616 1700 624
rect 1724 576 1732 584
rect 1692 536 1700 544
rect 1628 516 1636 524
rect 1596 296 1604 304
rect 1516 276 1524 284
rect 1660 496 1668 504
rect 1644 316 1652 324
rect 1676 276 1684 284
rect 1580 236 1588 244
rect 1628 236 1636 244
rect 1516 136 1524 144
rect 1868 606 1876 614
rect 1836 576 1844 584
rect 1788 536 1796 544
rect 1756 516 1764 524
rect 1996 536 2004 544
rect 1708 396 1716 404
rect 1804 376 1812 384
rect 1996 396 2004 404
rect 2028 396 2036 404
rect 1980 376 1988 384
rect 1820 276 1828 284
rect 1788 256 1796 264
rect 1788 236 1796 244
rect 1692 156 1700 164
rect 1660 136 1668 144
rect 1756 156 1764 164
rect 1756 136 1764 144
rect 1324 116 1332 124
rect 1388 116 1396 124
rect 1484 116 1492 124
rect 1564 116 1572 124
rect 1644 116 1652 124
rect 1868 206 1876 214
rect 1804 176 1812 184
rect 2252 736 2260 744
rect 2124 536 2132 544
rect 2076 296 2084 304
rect 2108 296 2116 304
rect 2252 296 2260 304
rect 1996 256 2004 264
rect 2060 276 2068 284
rect 2092 276 2100 284
rect 2028 236 2036 244
rect 2060 196 2068 204
rect 2156 196 2164 204
rect 1788 116 1796 124
rect 2252 96 2260 104
rect 1020 16 1028 24
rect 1068 16 1076 24
rect 1340 6 1348 14
<< metal3 >>
rect 408 2014 424 2016
rect 408 2006 412 2014
rect 420 2006 424 2014
rect 408 2004 424 2006
rect 1336 2014 1352 2016
rect 1336 2006 1340 2014
rect 1348 2006 1352 2014
rect 1336 2004 1352 2006
rect 100 1937 284 1943
rect -19 1917 60 1923
rect 84 1897 124 1903
rect 260 1897 300 1903
rect 308 1897 364 1903
rect 404 1897 444 1903
rect 628 1897 684 1903
rect 836 1897 1356 1903
rect 1460 1897 1628 1903
rect 2084 1897 2124 1903
rect 2260 1897 2291 1903
rect -19 1877 12 1883
rect 20 1877 115 1883
rect 109 1864 115 1877
rect 164 1877 204 1883
rect 212 1877 252 1883
rect 436 1877 492 1883
rect 500 1877 556 1883
rect 756 1877 812 1883
rect 932 1877 956 1883
rect 116 1857 172 1863
rect 244 1857 332 1863
rect 340 1857 508 1863
rect 516 1857 604 1863
rect 756 1857 796 1863
rect 884 1857 924 1863
rect 980 1857 1052 1863
rect 1092 1857 1148 1863
rect 1860 1857 1980 1863
rect 2036 1857 2092 1863
rect 877 1843 883 1856
rect 596 1837 883 1843
rect 964 1837 1020 1843
rect 1773 1837 2060 1843
rect 1773 1823 1779 1837
rect 1732 1817 1779 1823
rect 1908 1817 1932 1823
rect 872 1814 888 1816
rect 872 1806 876 1814
rect 884 1806 888 1814
rect 872 1804 888 1806
rect 1864 1814 1880 1816
rect 1864 1806 1868 1814
rect 1876 1806 1880 1814
rect 1864 1804 1880 1806
rect 36 1797 380 1803
rect 388 1797 540 1803
rect 596 1797 716 1803
rect 84 1777 220 1783
rect 580 1777 620 1783
rect 1412 1777 1644 1783
rect 1844 1777 1852 1783
rect 2164 1777 2236 1783
rect 148 1757 220 1763
rect 532 1757 588 1763
rect 660 1757 876 1763
rect 1620 1757 1628 1763
rect 1780 1757 2076 1763
rect 148 1737 348 1743
rect 564 1737 684 1743
rect 692 1737 732 1743
rect 772 1737 860 1743
rect 868 1737 956 1743
rect 1012 1737 1036 1743
rect 1044 1737 1180 1743
rect 1604 1737 1692 1743
rect 1716 1737 1740 1743
rect 452 1717 524 1723
rect 676 1717 796 1723
rect 1028 1717 1084 1723
rect 1332 1717 1404 1723
rect 1412 1717 1436 1723
rect 1444 1717 1772 1723
rect 1796 1717 1868 1723
rect 68 1697 556 1703
rect 564 1697 588 1703
rect 772 1697 924 1703
rect 932 1697 988 1703
rect 1060 1697 1132 1703
rect 1140 1697 1212 1703
rect 724 1677 748 1683
rect 408 1614 424 1616
rect 408 1606 412 1614
rect 420 1606 424 1614
rect 408 1604 424 1606
rect 1336 1614 1352 1616
rect 1336 1606 1340 1614
rect 1348 1606 1352 1614
rect 1336 1604 1352 1606
rect 868 1597 940 1603
rect 2020 1597 2076 1603
rect 500 1557 716 1563
rect 308 1537 636 1543
rect 164 1517 764 1523
rect -19 1497 12 1503
rect 68 1497 76 1503
rect 372 1497 412 1503
rect 420 1497 780 1503
rect 1220 1497 1708 1503
rect 2260 1497 2291 1503
rect 132 1477 444 1483
rect 980 1477 1276 1483
rect 1796 1477 1980 1483
rect 340 1457 716 1463
rect 724 1457 892 1463
rect 900 1457 908 1463
rect 1204 1457 1404 1463
rect 1844 1457 2172 1463
rect 1092 1437 1180 1443
rect 1556 1437 1628 1443
rect 1380 1417 1452 1423
rect 1620 1417 1644 1423
rect 872 1414 888 1416
rect 872 1406 876 1414
rect 884 1406 888 1414
rect 872 1404 888 1406
rect 1864 1414 1880 1416
rect 1864 1406 1868 1414
rect 1876 1406 1880 1414
rect 1864 1404 1880 1406
rect 20 1397 636 1403
rect 548 1377 892 1383
rect 1172 1377 1372 1383
rect 1380 1377 1676 1383
rect 68 1357 92 1363
rect 100 1357 140 1363
rect 148 1357 300 1363
rect 308 1357 396 1363
rect 868 1357 908 1363
rect 916 1357 1052 1363
rect 1508 1357 1516 1363
rect 1524 1357 1580 1363
rect 1636 1357 1708 1363
rect 1732 1357 2028 1363
rect 52 1337 76 1343
rect 84 1337 620 1343
rect 1204 1337 1436 1343
rect 1444 1337 1468 1343
rect 1700 1337 1788 1343
rect 36 1317 172 1323
rect 436 1317 492 1323
rect 500 1317 556 1323
rect 1284 1317 1340 1323
rect 1572 1317 1580 1323
rect 1588 1317 2172 1323
rect -19 1297 12 1303
rect 132 1297 476 1303
rect 484 1297 540 1303
rect 628 1297 716 1303
rect 1524 1297 1644 1303
rect 2260 1297 2291 1303
rect 164 1277 236 1283
rect 468 1277 508 1283
rect 516 1277 604 1283
rect 1268 1277 1420 1283
rect 1428 1277 1548 1283
rect 1556 1277 1756 1283
rect 452 1257 556 1263
rect 308 1237 460 1243
rect 788 1217 828 1223
rect 408 1214 424 1216
rect 408 1206 412 1214
rect 420 1206 424 1214
rect 408 1204 424 1206
rect 1336 1214 1352 1216
rect 1336 1206 1340 1214
rect 1348 1206 1352 1214
rect 1336 1204 1352 1206
rect 196 1197 268 1203
rect 20 1177 76 1183
rect 84 1177 252 1183
rect 356 1157 652 1163
rect 596 1137 732 1143
rect 740 1137 1068 1143
rect 948 1117 1020 1123
rect 1028 1117 1228 1123
rect 1236 1117 1276 1123
rect -19 1097 12 1103
rect 628 1097 684 1103
rect 692 1097 716 1103
rect 868 1097 908 1103
rect 916 1097 1068 1103
rect 1140 1097 1404 1103
rect 1620 1097 1836 1103
rect 2084 1097 2188 1103
rect 2260 1097 2291 1103
rect 244 1077 332 1083
rect 532 1077 700 1083
rect 708 1077 956 1083
rect 1060 1077 1148 1083
rect 1764 1077 2156 1083
rect 148 1057 428 1063
rect 436 1057 460 1063
rect 1140 1057 1180 1063
rect 1316 1057 1420 1063
rect 1428 1057 1532 1063
rect 1748 1057 1932 1063
rect 2132 1057 2172 1063
rect 1220 1037 1228 1043
rect 1508 1037 1532 1043
rect 872 1014 888 1016
rect 872 1006 876 1014
rect 884 1006 888 1014
rect 872 1004 888 1006
rect 1864 1014 1880 1016
rect 1864 1006 1868 1014
rect 1876 1006 1880 1014
rect 1864 1004 1880 1006
rect 116 997 156 1003
rect 164 997 348 1003
rect 356 997 524 1003
rect 532 997 604 1003
rect 612 997 764 1003
rect 1188 997 1228 1003
rect 1652 997 1708 1003
rect 1556 977 1788 983
rect 84 957 204 963
rect 212 957 252 963
rect 724 957 780 963
rect 1060 957 1196 963
rect 1204 957 1308 963
rect 1412 957 1452 963
rect 1572 957 1580 963
rect -19 937 12 943
rect 20 937 204 943
rect 253 943 259 956
rect 253 937 316 943
rect 548 937 588 943
rect 612 937 812 943
rect 1396 937 1740 943
rect 1956 937 2204 943
rect 68 917 124 923
rect 228 917 252 923
rect 260 917 412 923
rect 900 917 1116 923
rect 1460 917 1500 923
rect 1508 917 1548 923
rect 1620 917 1676 923
rect 2164 917 2188 923
rect -19 897 92 903
rect 100 897 284 903
rect 404 897 460 903
rect 1444 897 1484 903
rect 1492 897 1596 903
rect 148 877 172 883
rect 260 877 428 883
rect 1460 877 1516 883
rect 1780 877 1980 883
rect 164 857 556 863
rect 1716 857 1724 863
rect 1732 857 1788 863
rect 1332 837 1388 843
rect 1700 837 1756 843
rect 1764 837 1772 843
rect 2116 837 2172 843
rect 788 817 796 823
rect 980 817 1004 823
rect 408 814 424 816
rect 408 806 412 814
rect 420 806 424 814
rect 408 804 424 806
rect 1336 814 1352 816
rect 1336 806 1340 814
rect 1348 806 1352 814
rect 1336 804 1352 806
rect 692 797 988 803
rect 996 797 1244 803
rect 468 757 524 763
rect -19 737 60 743
rect 532 737 572 743
rect 596 737 668 743
rect 749 737 1212 743
rect 749 724 755 737
rect 1220 737 1388 743
rect 2260 737 2291 743
rect 324 717 476 723
rect 564 717 700 723
rect 708 717 748 723
rect 836 717 892 723
rect 900 717 924 723
rect -19 697 12 703
rect 52 697 124 703
rect 500 697 540 703
rect 621 697 636 703
rect 644 697 700 703
rect 868 697 908 703
rect 1508 697 1644 703
rect 1988 697 2124 703
rect 2164 697 2291 703
rect 580 677 796 683
rect 820 677 1020 683
rect 1220 677 1228 683
rect 1428 677 1772 683
rect 2036 677 2108 683
rect 2148 677 2172 683
rect 2180 677 2204 683
rect 100 657 476 663
rect 484 657 620 663
rect 1748 657 2044 663
rect 804 637 1228 643
rect 1588 637 1628 643
rect 1780 637 2076 643
rect 244 617 284 623
rect 1060 617 1132 623
rect 1396 617 1692 623
rect 872 614 888 616
rect 872 606 876 614
rect 884 606 888 614
rect 872 604 888 606
rect 1864 614 1880 616
rect 1864 606 1868 614
rect 1876 606 1880 614
rect 1864 604 1880 606
rect 1236 577 1708 583
rect 1716 577 1724 583
rect 1732 577 1836 583
rect 84 557 412 563
rect 612 557 1020 563
rect 1044 557 1484 563
rect 468 537 492 543
rect 580 537 684 543
rect 1636 537 1692 543
rect 1700 537 1788 543
rect 2004 537 2124 543
rect 276 517 460 523
rect 548 517 668 523
rect 1396 517 1628 523
rect 1636 517 1756 523
rect -19 497 12 503
rect 644 497 860 503
rect 868 497 1228 503
rect 1252 497 1660 503
rect 516 477 572 483
rect 596 477 620 483
rect 196 417 236 423
rect 324 417 348 423
rect 408 414 424 416
rect 408 406 412 414
rect 420 406 424 414
rect 408 404 424 406
rect 1336 414 1352 416
rect 1336 406 1340 414
rect 1348 406 1352 414
rect 1336 404 1352 406
rect 1604 397 1708 403
rect 2004 397 2028 403
rect 36 377 108 383
rect 1236 377 1500 383
rect 1508 377 1596 383
rect 1812 377 1980 383
rect 1588 317 1644 323
rect 420 297 444 303
rect 452 297 556 303
rect 852 297 892 303
rect 916 297 956 303
rect 964 297 1052 303
rect 1604 297 2076 303
rect 2084 297 2108 303
rect 2260 297 2291 303
rect 228 277 364 283
rect 436 277 492 283
rect 532 277 748 283
rect 1012 277 1148 283
rect 1252 277 1516 283
rect 1684 277 1820 283
rect 2068 277 2092 283
rect 196 257 636 263
rect 644 257 716 263
rect 724 257 828 263
rect 1140 257 1164 263
rect 1172 257 1276 263
rect 1284 257 1452 263
rect 1460 257 1788 263
rect 1796 257 1996 263
rect 1588 237 1628 243
rect 1796 237 2028 243
rect 872 214 888 216
rect 872 206 876 214
rect 884 206 888 214
rect 872 204 888 206
rect 1864 214 1880 216
rect 1864 206 1868 214
rect 1876 206 1880 214
rect 1864 204 1880 206
rect 1901 197 2060 203
rect 1901 183 1907 197
rect 2068 197 2156 203
rect 1812 177 1907 183
rect 36 157 364 163
rect 964 157 1036 163
rect 1700 157 1756 163
rect 228 137 444 143
rect 1108 137 1420 143
rect 1492 137 1516 143
rect 1565 137 1660 143
rect 1565 124 1571 137
rect 1716 137 1756 143
rect 324 117 556 123
rect 772 117 844 123
rect 1332 117 1388 123
rect 1492 117 1564 123
rect 1652 117 1788 123
rect 2260 97 2291 103
rect 996 37 1004 43
rect 628 17 668 23
rect 1028 17 1068 23
rect 408 14 424 16
rect 408 6 412 14
rect 420 6 424 14
rect 408 4 424 6
rect 1336 14 1352 16
rect 1336 6 1340 14
rect 1348 6 1352 14
rect 1336 4 1352 6
<< m4contact >>
rect 412 2006 420 2014
rect 1340 2006 1348 2014
rect 1836 1996 1844 2004
rect 204 1876 212 1884
rect 876 1806 884 1814
rect 1868 1806 1876 1814
rect 1836 1776 1844 1784
rect 1612 1756 1620 1764
rect 412 1606 420 1614
rect 1340 1606 1348 1614
rect 1676 1576 1684 1584
rect 76 1496 84 1504
rect 364 1496 372 1504
rect 716 1456 724 1464
rect 908 1456 916 1464
rect 1548 1436 1556 1444
rect 1612 1416 1620 1424
rect 876 1406 884 1414
rect 1868 1406 1876 1414
rect 12 1396 20 1404
rect 1676 1376 1684 1384
rect 908 1356 916 1364
rect 76 1336 84 1344
rect 1580 1316 1588 1324
rect 12 1296 20 1304
rect 412 1206 420 1214
rect 1340 1206 1348 1214
rect 364 1096 372 1104
rect 908 1096 916 1104
rect 1132 1056 1140 1064
rect 1228 1036 1236 1044
rect 876 1006 884 1014
rect 1868 1006 1876 1014
rect 1708 996 1716 1004
rect 780 976 788 984
rect 204 956 212 964
rect 716 956 724 964
rect 1580 956 1588 964
rect 1548 916 1556 924
rect 1708 856 1716 864
rect 1388 836 1396 844
rect 1772 836 1780 844
rect 780 816 788 824
rect 1004 816 1012 824
rect 412 806 420 814
rect 1340 806 1348 814
rect 908 696 916 704
rect 1228 676 1236 684
rect 1772 636 1780 644
rect 1132 616 1140 624
rect 876 606 884 614
rect 1868 606 1876 614
rect 1708 576 1716 584
rect 1388 516 1396 524
rect 412 406 420 414
rect 1340 406 1348 414
rect 908 296 916 304
rect 876 206 884 214
rect 1868 206 1876 214
rect 1708 136 1716 144
rect 1004 36 1012 44
rect 412 6 420 14
rect 1340 6 1348 14
<< metal4 >>
rect 408 2014 424 2040
rect 408 2006 412 2014
rect 420 2006 424 2014
rect 202 1884 214 1886
rect 202 1876 204 1884
rect 212 1876 214 1884
rect 74 1504 86 1506
rect 74 1496 76 1504
rect 84 1496 86 1504
rect 10 1404 22 1406
rect 10 1396 12 1404
rect 20 1396 22 1404
rect 10 1304 22 1396
rect 74 1344 86 1496
rect 74 1336 76 1344
rect 84 1336 86 1344
rect 74 1334 86 1336
rect 10 1296 12 1304
rect 20 1296 22 1304
rect 10 1294 22 1296
rect 202 964 214 1876
rect 408 1614 424 2006
rect 408 1606 412 1614
rect 420 1606 424 1614
rect 362 1504 374 1506
rect 362 1496 364 1504
rect 372 1496 374 1504
rect 362 1104 374 1496
rect 362 1096 364 1104
rect 372 1096 374 1104
rect 362 1094 374 1096
rect 408 1214 424 1606
rect 872 1814 888 2040
rect 872 1806 876 1814
rect 884 1806 888 1814
rect 408 1206 412 1214
rect 420 1206 424 1214
rect 202 956 204 964
rect 212 956 214 964
rect 202 954 214 956
rect 408 814 424 1206
rect 714 1464 726 1466
rect 714 1456 716 1464
rect 724 1456 726 1464
rect 714 964 726 1456
rect 872 1414 888 1806
rect 1336 2014 1352 2040
rect 1336 2006 1340 2014
rect 1348 2006 1352 2014
rect 1336 1614 1352 2006
rect 1834 2004 1846 2006
rect 1834 1996 1836 2004
rect 1844 1996 1846 2004
rect 1834 1784 1846 1996
rect 1834 1776 1836 1784
rect 1844 1776 1846 1784
rect 1834 1774 1846 1776
rect 1864 1814 1880 2040
rect 1864 1806 1868 1814
rect 1876 1806 1880 1814
rect 1336 1606 1340 1614
rect 1348 1606 1352 1614
rect 872 1406 876 1414
rect 884 1406 888 1414
rect 872 1014 888 1406
rect 906 1464 918 1466
rect 906 1456 908 1464
rect 916 1456 918 1464
rect 906 1364 918 1456
rect 906 1356 908 1364
rect 916 1356 918 1364
rect 906 1354 918 1356
rect 1336 1214 1352 1606
rect 1610 1764 1622 1766
rect 1610 1756 1612 1764
rect 1620 1756 1622 1764
rect 1336 1206 1340 1214
rect 1348 1206 1352 1214
rect 872 1006 876 1014
rect 884 1006 888 1014
rect 714 956 716 964
rect 724 956 726 964
rect 714 954 726 956
rect 778 984 790 986
rect 778 976 780 984
rect 788 976 790 984
rect 778 824 790 976
rect 778 816 780 824
rect 788 816 790 824
rect 778 814 790 816
rect 408 806 412 814
rect 420 806 424 814
rect 408 414 424 806
rect 408 406 412 414
rect 420 406 424 414
rect 408 14 424 406
rect 408 6 412 14
rect 420 6 424 14
rect 408 -40 424 6
rect 872 614 888 1006
rect 872 606 876 614
rect 884 606 888 614
rect 872 214 888 606
rect 906 1104 918 1106
rect 906 1096 908 1104
rect 916 1096 918 1104
rect 906 704 918 1096
rect 1130 1064 1142 1066
rect 1130 1056 1132 1064
rect 1140 1056 1142 1064
rect 906 696 908 704
rect 916 696 918 704
rect 906 304 918 696
rect 906 296 908 304
rect 916 296 918 304
rect 906 294 918 296
rect 1002 824 1014 826
rect 1002 816 1004 824
rect 1012 816 1014 824
rect 872 206 876 214
rect 884 206 888 214
rect 872 -40 888 206
rect 1002 44 1014 816
rect 1130 624 1142 1056
rect 1226 1044 1238 1046
rect 1226 1036 1228 1044
rect 1236 1036 1238 1044
rect 1226 684 1238 1036
rect 1226 676 1228 684
rect 1236 676 1238 684
rect 1226 674 1238 676
rect 1336 814 1352 1206
rect 1546 1444 1558 1446
rect 1546 1436 1548 1444
rect 1556 1436 1558 1444
rect 1546 924 1558 1436
rect 1610 1424 1622 1756
rect 1610 1416 1612 1424
rect 1620 1416 1622 1424
rect 1610 1414 1622 1416
rect 1674 1584 1686 1586
rect 1674 1576 1676 1584
rect 1684 1576 1686 1584
rect 1674 1384 1686 1576
rect 1674 1376 1676 1384
rect 1684 1376 1686 1384
rect 1674 1374 1686 1376
rect 1864 1414 1880 1806
rect 1864 1406 1868 1414
rect 1876 1406 1880 1414
rect 1578 1324 1590 1326
rect 1578 1316 1580 1324
rect 1588 1316 1590 1324
rect 1578 964 1590 1316
rect 1864 1014 1880 1406
rect 1864 1006 1868 1014
rect 1876 1006 1880 1014
rect 1578 956 1580 964
rect 1588 956 1590 964
rect 1578 954 1590 956
rect 1706 1004 1718 1006
rect 1706 996 1708 1004
rect 1716 996 1718 1004
rect 1546 916 1548 924
rect 1556 916 1558 924
rect 1546 914 1558 916
rect 1706 864 1718 996
rect 1706 856 1708 864
rect 1716 856 1718 864
rect 1336 806 1340 814
rect 1348 806 1352 814
rect 1130 616 1132 624
rect 1140 616 1142 624
rect 1130 614 1142 616
rect 1002 36 1004 44
rect 1012 36 1014 44
rect 1002 34 1014 36
rect 1336 414 1352 806
rect 1386 844 1398 846
rect 1386 836 1388 844
rect 1396 836 1398 844
rect 1386 524 1398 836
rect 1386 516 1388 524
rect 1396 516 1398 524
rect 1386 514 1398 516
rect 1706 584 1718 856
rect 1770 844 1782 846
rect 1770 836 1772 844
rect 1780 836 1782 844
rect 1770 644 1782 836
rect 1770 636 1772 644
rect 1780 636 1782 644
rect 1770 634 1782 636
rect 1706 576 1708 584
rect 1716 576 1718 584
rect 1336 406 1340 414
rect 1348 406 1352 414
rect 1336 14 1352 406
rect 1706 144 1718 576
rect 1706 136 1708 144
rect 1716 136 1718 144
rect 1706 134 1718 136
rect 1864 614 1880 1006
rect 1864 606 1868 614
rect 1876 606 1880 614
rect 1864 214 1880 606
rect 1864 206 1868 214
rect 1876 206 1880 214
rect 1336 6 1340 14
rect 1348 6 1352 14
rect 1336 -40 1352 6
rect 1864 -40 1880 206
use FILL  FILL_55
timestamp 1739819275
transform -1 0 376 0 1 210
box -16 -6 32 210
use FILL  FILL_54
timestamp 1739819275
transform 1 0 360 0 -1 210
box -16 -6 32 210
use NOR2X1  NOR2X1_13
timestamp 1739819275
transform 1 0 376 0 -1 210
box -16 -6 64 210
use DFFSR  DFFSR_32
timestamp 1739819275
transform -1 0 360 0 1 210
box -16 -6 368 210
use DFFSR  DFFSR_31
timestamp 1739819275
transform -1 0 360 0 -1 210
box -16 -6 368 210
use AND2X2  AND2X2_3
timestamp 1739819275
transform -1 0 440 0 1 210
box -16 -6 80 210
use INVX1  INVX1_34
timestamp 1739819275
transform 1 0 440 0 1 210
box -18 -6 52 210
use INVX1  INVX1_33
timestamp 1739819275
transform -1 0 456 0 -1 210
box -18 -6 52 210
use DFFSR  DFFSR_30
timestamp 1739819275
transform -1 0 888 0 1 210
box -16 -6 368 210
use DFFSR  DFFSR_29
timestamp 1739819275
transform -1 0 808 0 -1 210
box -16 -6 368 210
use OAI21X1  OAI21X1_29
timestamp 1739819275
transform 1 0 472 0 1 210
box -16 -6 68 210
use FILL  FILL_53
timestamp 1739819275
transform -1 0 904 0 1 210
box -16 -6 32 210
use FILL  FILL_52
timestamp 1739819275
transform -1 0 824 0 -1 210
box -16 -6 32 210
use DFFSR  DFFSR_28
timestamp 1739819275
transform 1 0 1112 0 1 210
box -16 -6 368 210
use DFFSR  DFFSR_27
timestamp 1739819275
transform 1 0 968 0 -1 210
box -16 -6 368 210
use CLKBUF1  CLKBUF1_4
timestamp 1739819275
transform -1 0 968 0 -1 210
box -16 -6 160 210
use BUFX4  BUFX4_8
timestamp 1739819275
transform 1 0 968 0 1 210
box -18 -6 74 210
use BUFX4  BUFX4_7
timestamp 1739819275
transform -1 0 968 0 1 210
box -18 -6 74 210
use INVX8  INVX8_1
timestamp 1739819275
transform 1 0 1032 0 1 210
box -18 -6 90 210
use FILL  FILL_51
timestamp 1739819275
transform 1 0 1464 0 1 210
box -16 -6 32 210
use FILL  FILL_50
timestamp 1739819275
transform 1 0 1368 0 -1 210
box -16 -6 32 210
use BUFX2  BUFX2_25
timestamp 1739819275
transform 1 0 1512 0 -1 210
box -10 -6 56 210
use BUFX2  BUFX2_24
timestamp 1739819275
transform 1 0 1320 0 -1 210
box -10 -6 56 210
use INVX1  INVX1_32
timestamp 1739819275
transform 1 0 1480 0 1 210
box -18 -6 52 210
use INVX1  INVX1_31
timestamp 1739819275
transform 1 0 1384 0 -1 210
box -18 -6 52 210
use MUX2X1  MUX2X1_6
timestamp 1739819275
transform -1 0 1608 0 1 210
box -10 -6 106 210
use MUX2X1  MUX2X1_5
timestamp 1739819275
transform -1 0 1512 0 -1 210
box -10 -6 106 210
use FILL  FILL_49
timestamp 1739819275
transform 1 0 1816 0 -1 210
box -16 -6 32 210
use BUFX2  BUFX2_23
timestamp 1739819275
transform 1 0 1704 0 -1 210
box -10 -6 56 210
use BUFX2  BUFX2_22
timestamp 1739819275
transform 1 0 1592 0 -1 210
box -10 -6 56 210
use INVX1  INVX1_30
timestamp 1739819275
transform -1 0 1592 0 -1 210
box -18 -6 52 210
use AOI21X1  AOI21X1_13
timestamp 1739819275
transform 1 0 1640 0 -1 210
box -14 -6 78 210
use DFFSR  DFFSR_26
timestamp 1739819275
transform 1 0 1832 0 -1 210
box -16 -6 368 210
use DFFSR  DFFSR_25
timestamp 1739819275
transform -1 0 1960 0 1 210
box -16 -6 368 210
use OAI21X1  OAI21X1_28
timestamp 1739819275
transform -1 0 1816 0 -1 210
box -16 -6 68 210
use FILL  FILL_48
timestamp 1739819275
transform -1 0 1976 0 1 210
box -16 -6 32 210
use INVX1  INVX1_29
timestamp 1739819275
transform -1 0 2072 0 1 210
box -18 -6 52 210
use AOI21X1  AOI21X1_12
timestamp 1739819275
transform -1 0 2040 0 1 210
box -14 -6 78 210
use MUX2X1  MUX2X1_4
timestamp 1739819275
transform 1 0 2072 0 1 210
box -10 -6 106 210
use FILL  FILL_45
timestamp 1739819275
transform 1 0 2248 0 1 210
box -16 -6 32 210
use FILL  FILL_46
timestamp 1739819275
transform -1 0 2264 0 -1 210
box -16 -6 32 210
use FILL  FILL_47
timestamp 1739819275
transform -1 0 2248 0 -1 210
box -16 -6 32 210
use BUFX2  BUFX2_20
timestamp 1739819275
transform 1 0 2200 0 1 210
box -10 -6 56 210
use BUFX2  BUFX2_21
timestamp 1739819275
transform 1 0 2184 0 -1 210
box -10 -6 56 210
use INVX1  INVX1_28
timestamp 1739819275
transform -1 0 2200 0 1 210
box -18 -6 52 210
use BUFX2  BUFX2_19
timestamp 1739819275
transform -1 0 56 0 -1 610
box -10 -6 56 210
use DFFSR  DFFSR_24
timestamp 1739819275
transform -1 0 408 0 -1 610
box -16 -6 368 210
use FILL  FILL_44
timestamp 1739819275
transform 1 0 408 0 -1 610
box -16 -6 32 210
use INVX1  INVX1_27
timestamp 1739819275
transform -1 0 648 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_26
timestamp 1739819275
transform -1 0 552 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_25
timestamp 1739819275
transform 1 0 424 0 -1 610
box -18 -6 52 210
use AOI21X1  AOI21X1_11
timestamp 1739819275
transform -1 0 520 0 -1 610
box -14 -6 78 210
use DFFSR  DFFSR_23
timestamp 1739819275
transform -1 0 1000 0 -1 610
box -16 -6 368 210
use NAND3X1  NAND3X1_11
timestamp 1739819275
transform 1 0 552 0 -1 610
box -16 -6 80 210
use FILL  FILL_43
timestamp 1739819275
transform 1 0 1000 0 -1 610
box -16 -6 32 210
use INVX1  INVX1_24
timestamp 1739819275
transform 1 0 1016 0 -1 610
box -18 -6 52 210
use CLKBUF1  CLKBUF1_3
timestamp 1739819275
transform 1 0 1048 0 -1 610
box -16 -6 160 210
use FILL  FILL_42
timestamp 1739819275
transform -1 0 1272 0 -1 610
box -16 -6 32 210
use DFFSR  DFFSR_22
timestamp 1739819275
transform -1 0 1624 0 -1 610
box -16 -6 368 210
use NAND3X1  NAND3X1_10
timestamp 1739819275
transform -1 0 1256 0 -1 610
box -16 -6 80 210
use FILL  FILL_41
timestamp 1739819275
transform 1 0 1848 0 -1 610
box -16 -6 32 210
use INVX1  INVX1_23
timestamp 1739819275
transform 1 0 1624 0 -1 610
box -18 -6 52 210
use AOI21X1  AOI21X1_10
timestamp 1739819275
transform 1 0 1656 0 -1 610
box -14 -6 78 210
use DFFSR  DFFSR_21
timestamp 1739819275
transform 1 0 1864 0 -1 610
box -16 -6 368 210
use OAI21X1  OAI21X1_27
timestamp 1739819275
transform 1 0 1784 0 -1 610
box -16 -6 68 210
use OAI21X1  OAI21X1_26
timestamp 1739819275
transform -1 0 1784 0 -1 610
box -16 -6 68 210
use FILL  FILL_40
timestamp 1739819275
transform -1 0 2264 0 -1 610
box -16 -6 32 210
use INVX1  INVX1_22
timestamp 1739819275
transform 1 0 2216 0 -1 610
box -18 -6 52 210
use BUFX2  BUFX2_18
timestamp 1739819275
transform -1 0 104 0 1 610
box -10 -6 56 210
use BUFX2  BUFX2_17
timestamp 1739819275
transform -1 0 56 0 1 610
box -10 -6 56 210
use DFFSR  DFFSR_20
timestamp 1739819275
transform -1 0 456 0 1 610
box -16 -6 368 210
use FILL  FILL_39
timestamp 1739819275
transform 1 0 456 0 1 610
box -16 -6 32 210
use INVX1  INVX1_21
timestamp 1739819275
transform 1 0 472 0 1 610
box -18 -6 52 210
use NAND2X1  NAND2X1_6
timestamp 1739819275
transform -1 0 808 0 1 610
box -16 -6 64 210
use OAI21X1  OAI21X1_25
timestamp 1739819275
transform 1 0 696 0 1 610
box -16 -6 68 210
use OAI21X1  OAI21X1_24
timestamp 1739819275
transform -1 0 696 0 1 610
box -16 -6 68 210
use NAND3X1  NAND3X1_9
timestamp 1739819275
transform 1 0 568 0 1 610
box -16 -6 80 210
use NAND3X1  NAND3X1_8
timestamp 1739819275
transform -1 0 568 0 1 610
box -16 -6 80 210
use FILL  FILL_38
timestamp 1739819275
transform 1 0 872 0 1 610
box -16 -6 32 210
use DFFSR  DFFSR_19
timestamp 1739819275
transform 1 0 888 0 1 610
box -16 -6 368 210
use BUFX4  BUFX4_6
timestamp 1739819275
transform -1 0 872 0 1 610
box -18 -6 74 210
use FILL  FILL_37
timestamp 1739819275
transform 1 0 1240 0 1 610
box -16 -6 32 210
use DFFSR  DFFSR_18
timestamp 1739819275
transform 1 0 1256 0 1 610
box -16 -6 368 210
use DFFSR  DFFSR_17
timestamp 1739819275
transform 1 0 1608 0 1 610
box -16 -6 368 210
use FILL  FILL_36
timestamp 1739819275
transform 1 0 2248 0 1 610
box -16 -6 32 210
use FILL  FILL_35
timestamp 1739819275
transform 1 0 2232 0 1 610
box -16 -6 32 210
use FILL  FILL_34
timestamp 1739819275
transform 1 0 2216 0 1 610
box -16 -6 32 210
use FILL  FILL_33
timestamp 1739819275
transform 1 0 1960 0 1 610
box -16 -6 32 210
use BUFX2  BUFX2_16
timestamp 1739819275
transform 1 0 2168 0 1 610
box -10 -6 56 210
use BUFX2  BUFX2_15
timestamp 1739819275
transform 1 0 2120 0 1 610
box -10 -6 56 210
use INVX1  INVX1_20
timestamp 1739819275
transform 1 0 1976 0 1 610
box -18 -6 52 210
use NOR2X1  NOR2X1_12
timestamp 1739819275
transform 1 0 2072 0 1 610
box -16 -6 64 210
use AOI21X1  AOI21X1_9
timestamp 1739819275
transform 1 0 2008 0 1 610
box -14 -6 78 210
use FILL  FILL_32
timestamp 1739819275
transform 1 0 360 0 -1 1010
box -16 -6 32 210
use INVX1  INVX1_19
timestamp 1739819275
transform 1 0 376 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_18
timestamp 1739819275
transform -1 0 296 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_17
timestamp 1739819275
transform -1 0 264 0 -1 1010
box -18 -6 52 210
use INVX1  INVX1_16
timestamp 1739819275
transform 1 0 8 0 -1 1010
box -18 -6 52 210
use OAI21X1  OAI21X1_23
timestamp 1739819275
transform 1 0 296 0 -1 1010
box -16 -6 68 210
use OAI21X1  OAI21X1_22
timestamp 1739819275
transform -1 0 104 0 -1 1010
box -16 -6 68 210
use NAND3X1  NAND3X1_7
timestamp 1739819275
transform -1 0 232 0 -1 1010
box -16 -6 80 210
use NAND3X1  NAND3X1_6
timestamp 1739819275
transform 1 0 104 0 -1 1010
box -16 -6 80 210
use DFFSR  DFFSR_16
timestamp 1739819275
transform -1 0 952 0 -1 1010
box -16 -6 368 210
use OAI21X1  OAI21X1_21
timestamp 1739819275
transform -1 0 536 0 -1 1010
box -16 -6 68 210
use OAI21X1  OAI21X1_20
timestamp 1739819275
transform 1 0 408 0 -1 1010
box -16 -6 68 210
use AND2X2  AND2X2_2
timestamp 1739819275
transform 1 0 536 0 -1 1010
box -16 -6 80 210
use FILL  FILL_31
timestamp 1739819275
transform -1 0 968 0 -1 1010
box -16 -6 32 210
use BUFX2  BUFX2_14
timestamp 1739819275
transform -1 0 1016 0 -1 1010
box -10 -6 56 210
use DFFSR  DFFSR_15
timestamp 1739819275
transform -1 0 1368 0 -1 1010
box -16 -6 368 210
use FILL  FILL_30
timestamp 1739819275
transform -1 0 1384 0 -1 1010
box -16 -6 32 210
use NOR2X1  NOR2X1_11
timestamp 1739819275
transform -1 0 1560 0 -1 1010
box -16 -6 64 210
use AOI21X1  AOI21X1_8
timestamp 1739819275
transform -1 0 1512 0 -1 1010
box -14 -6 78 210
use OAI21X1  OAI21X1_19
timestamp 1739819275
transform -1 0 1448 0 -1 1010
box -16 -6 68 210
use FILL  FILL_29
timestamp 1739819275
transform 1 0 1800 0 -1 1010
box -16 -6 32 210
use DFFSR  DFFSR_14
timestamp 1739819275
transform 1 0 1816 0 -1 1010
box -16 -6 368 210
use OAI21X1  OAI21X1_18
timestamp 1739819275
transform 1 0 1736 0 -1 1010
box -16 -6 68 210
use OAI21X1  OAI21X1_17
timestamp 1739819275
transform 1 0 1672 0 -1 1010
box -16 -6 68 210
use XNOR2X1  XNOR2X1_1
timestamp 1739819275
transform -1 0 1672 0 -1 1010
box -16 -6 128 210
use MUX2X1  MUX2X1_3
timestamp 1739819275
transform 1 0 2168 0 -1 1010
box -10 -6 106 210
use BUFX2  BUFX2_13
timestamp 1739819275
transform -1 0 56 0 1 1010
box -10 -6 56 210
use DFFSR  DFFSR_13
timestamp 1739819275
transform -1 0 408 0 1 1010
box -16 -6 368 210
use FILL  FILL_28
timestamp 1739819275
transform 1 0 408 0 1 1010
box -16 -6 32 210
use INVX1  INVX1_15
timestamp 1739819275
transform 1 0 424 0 1 1010
box -18 -6 52 210
use NOR2X1  NOR2X1_10
timestamp 1739819275
transform 1 0 536 0 1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_5
timestamp 1739819275
transform -1 0 632 0 1 1010
box -16 -6 64 210
use NAND3X1  NAND3X1_5
timestamp 1739819275
transform 1 0 696 0 1 1010
box -16 -6 80 210
use NAND3X1  NAND3X1_4
timestamp 1739819275
transform -1 0 696 0 1 1010
box -16 -6 80 210
use AOI22X1  AOI22X1_1
timestamp 1739819275
transform -1 0 536 0 1 1010
box -16 -6 92 210
use INVX4  INVX4_0
timestamp 1739819275
transform 1 0 760 0 1 1010
box -18 -6 56 210
use FILL  FILL_27
timestamp 1739819275
transform -1 0 888 0 1 1010
box -16 -6 32 210
use INVX1  INVX1_14
timestamp 1739819275
transform 1 0 1032 0 1 1010
box -18 -6 52 210
use MUX2X1  MUX2X1_2
timestamp 1739819275
transform -1 0 1224 0 1 1010
box -10 -6 106 210
use BUFX4  BUFX4_5
timestamp 1739819275
transform 1 0 1064 0 1 1010
box -18 -6 74 210
use BUFX4  BUFX4_4
timestamp 1739819275
transform -1 0 1032 0 1 1010
box -18 -6 74 210
use BUFX4  BUFX4_3
timestamp 1739819275
transform -1 0 872 0 1 1010
box -18 -6 74 210
use INVX8  INVX8_0
timestamp 1739819275
transform -1 0 968 0 1 1010
box -18 -6 90 210
use FILL  FILL_26
timestamp 1739819275
transform 1 0 1352 0 1 1010
box -16 -6 32 210
use DFFSR  DFFSR_12
timestamp 1739819275
transform 1 0 1368 0 1 1010
box -16 -6 368 210
use BUFX4  BUFX4_2
timestamp 1739819275
transform 1 0 1288 0 1 1010
box -18 -6 74 210
use BUFX4  BUFX4_1
timestamp 1739819275
transform 1 0 1224 0 1 1010
box -18 -6 74 210
use FILL  FILL_25
timestamp 1739819275
transform 1 0 1784 0 1 1010
box -16 -6 32 210
use AOI21X1  AOI21X1_7
timestamp 1739819275
transform -1 0 1784 0 1 1010
box -14 -6 78 210
use DFFSR  DFFSR_11
timestamp 1739819275
transform 1 0 1800 0 1 1010
box -16 -6 368 210
use FILL  FILL_24
timestamp 1739819275
transform 1 0 2248 0 1 1010
box -16 -6 32 210
use FILL  FILL_23
timestamp 1739819275
transform 1 0 2232 0 1 1010
box -16 -6 32 210
use BUFX2  BUFX2_12
timestamp 1739819275
transform 1 0 2184 0 1 1010
box -10 -6 56 210
use INVX1  INVX1_13
timestamp 1739819275
transform -1 0 2184 0 1 1010
box -18 -6 52 210
use FILL  FILL_22
timestamp 1739819275
transform 1 0 376 0 -1 1410
box -16 -6 32 210
use INVX1  INVX1_12
timestamp 1739819275
transform 1 0 392 0 -1 1410
box -18 -6 52 210
use INVX1  INVX1_11
timestamp 1739819275
transform 1 0 72 0 -1 1410
box -18 -6 52 210
use AOI21X1  AOI21X1_6
timestamp 1739819275
transform 1 0 104 0 -1 1410
box -14 -6 78 210
use OAI21X1  OAI21X1_16
timestamp 1739819275
transform -1 0 72 0 -1 1410
box -16 -6 68 210
use NOR3X1  NOR3X1_0
timestamp 1739819275
transform 1 0 248 0 -1 1410
box -14 -6 136 210
use AOI22X1  AOI22X1_0
timestamp 1739819275
transform -1 0 248 0 -1 1410
box -16 -6 92 210
use BUFX2  BUFX2_11
timestamp 1739819275
transform -1 0 680 0 -1 1410
box -10 -6 56 210
use INVX1  INVX1_10
timestamp 1739819275
transform -1 0 632 0 -1 1410
box -18 -6 52 210
use NOR2X1  NOR2X1_9
timestamp 1739819275
transform 1 0 424 0 -1 1410
box -16 -6 64 210
use DFFSR  DFFSR_10
timestamp 1739819275
transform -1 0 1032 0 -1 1410
box -16 -6 368 210
use NAND3X1  NAND3X1_3
timestamp 1739819275
transform 1 0 536 0 -1 1410
box -16 -6 80 210
use NAND3X1  NAND3X1_2
timestamp 1739819275
transform 1 0 472 0 -1 1410
box -16 -6 80 210
use FILL  FILL_21
timestamp 1739819275
transform -1 0 1048 0 -1 1410
box -16 -6 32 210
use CLKBUF1  CLKBUF1_2
timestamp 1739819275
transform -1 0 1192 0 -1 1410
box -16 -6 160 210
use FILL  FILL_20
timestamp 1739819275
transform 1 0 1400 0 -1 1410
box -16 -6 32 210
use INVX1  INVX1_9
timestamp 1739819275
transform -1 0 1512 0 -1 1410
box -18 -6 52 210
use AOI21X1  AOI21X1_5
timestamp 1739819275
transform 1 0 1416 0 -1 1410
box -14 -6 78 210
use OAI21X1  OAI21X1_15
timestamp 1739819275
transform -1 0 1576 0 -1 1410
box -16 -6 68 210
use CLKBUF1  CLKBUF1_1
timestamp 1739819275
transform 1 0 1192 0 -1 1410
box -16 -6 160 210
use BUFX4  BUFX4_0
timestamp 1739819275
transform 1 0 1336 0 -1 1410
box -18 -6 74 210
use FILL  FILL_19
timestamp 1739819275
transform -1 0 1816 0 -1 1410
box -16 -6 32 210
use INVX1  INVX1_8
timestamp 1739819275
transform -1 0 1800 0 -1 1410
box -18 -6 52 210
use AOI21X1  AOI21X1_4
timestamp 1739819275
transform -1 0 1768 0 -1 1410
box -14 -6 78 210
use DFFSR  DFFSR_9
timestamp 1739819275
transform -1 0 2168 0 -1 1410
box -16 -6 368 210
use OAI21X1  OAI21X1_14
timestamp 1739819275
transform -1 0 1704 0 -1 1410
box -16 -6 68 210
use OAI21X1  OAI21X1_13
timestamp 1739819275
transform 1 0 1576 0 -1 1410
box -16 -6 68 210
use FILL  FILL_18
timestamp 1739819275
transform -1 0 2264 0 -1 1410
box -16 -6 32 210
use FILL  FILL_17
timestamp 1739819275
transform -1 0 2248 0 -1 1410
box -16 -6 32 210
use FILL  FILL_16
timestamp 1739819275
transform -1 0 2232 0 -1 1410
box -16 -6 32 210
use BUFX2  BUFX2_10
timestamp 1739819275
transform 1 0 2168 0 -1 1410
box -10 -6 56 210
use BUFX2  BUFX2_9
timestamp 1739819275
transform -1 0 56 0 1 1410
box -10 -6 56 210
use NOR2X1  NOR2X1_8
timestamp 1739819275
transform -1 0 104 0 1 1410
box -16 -6 64 210
use DFFSR  DFFSR_8
timestamp 1739819275
transform 1 0 168 0 1 1410
box -16 -6 368 210
use OAI21X1  OAI21X1_12
timestamp 1739819275
transform 1 0 104 0 1 1410
box -16 -6 68 210
use FILL  FILL_15
timestamp 1739819275
transform 1 0 712 0 1 1410
box -16 -6 32 210
use FILL  FILL_14
timestamp 1739819275
transform -1 0 536 0 1 1410
box -16 -6 32 210
use NOR2X1  NOR2X1_7
timestamp 1739819275
transform 1 0 664 0 1 1410
box -16 -6 64 210
use DFFSR  DFFSR_7
timestamp 1739819275
transform 1 0 728 0 1 1410
box -16 -6 368 210
use OAI21X1  OAI21X1_11
timestamp 1739819275
transform -1 0 600 0 1 1410
box -16 -6 68 210
use AND2X2  AND2X2_1
timestamp 1739819275
transform -1 0 664 0 1 1410
box -16 -6 80 210
use CLKBUF1  CLKBUF1_0
timestamp 1739819275
transform 1 0 1080 0 1 1410
box -16 -6 160 210
use FILL  FILL_13
timestamp 1739819275
transform 1 0 1224 0 1 1410
box -16 -6 32 210
use DFFSR  DFFSR_6
timestamp 1739819275
transform 1 0 1240 0 1 1410
box -16 -6 368 210
use FILL  FILL_12
timestamp 1739819275
transform 1 0 1832 0 1 1410
box -16 -6 32 210
use INVX1  INVX1_7
timestamp 1739819275
transform -1 0 1832 0 1 1410
box -18 -6 52 210
use DFFSR  DFFSR_5
timestamp 1739819275
transform 1 0 1848 0 1 1410
box -16 -6 368 210
use MUX2X1  MUX2X1_1
timestamp 1739819275
transform 1 0 1704 0 1 1410
box -10 -6 106 210
use XNOR2X1  XNOR2X1_0
timestamp 1739819275
transform 1 0 1592 0 1 1410
box -16 -6 128 210
use FILL  FILL_11
timestamp 1739819275
transform 1 0 2248 0 1 1410
box -16 -6 32 210
use BUFX2  BUFX2_8
timestamp 1739819275
transform 1 0 2200 0 1 1410
box -10 -6 56 210
use DFFSR  DFFSR_4
timestamp 1739819275
transform -1 0 488 0 -1 1810
box -16 -6 368 210
use OAI21X1  OAI21X1_10
timestamp 1739819275
transform 1 0 72 0 -1 1810
box -16 -6 68 210
use OAI21X1  OAI21X1_9
timestamp 1739819275
transform 1 0 8 0 -1 1810
box -16 -6 68 210
use FILL  FILL_10
timestamp 1739819275
transform -1 0 504 0 -1 1810
box -16 -6 32 210
use OAI21X1  OAI21X1_8
timestamp 1739819275
transform -1 0 760 0 -1 1810
box -16 -6 68 210
use OAI21X1  OAI21X1_7
timestamp 1739819275
transform -1 0 696 0 -1 1810
box -16 -6 68 210
use OAI21X1  OAI21X1_6
timestamp 1739819275
transform 1 0 568 0 -1 1810
box -16 -6 68 210
use NAND3X1  NAND3X1_1
timestamp 1739819275
transform -1 0 568 0 -1 1810
box -16 -6 80 210
use XOR2X1  XOR2X1_0
timestamp 1739819275
transform -1 0 872 0 -1 1810
box -16 -6 128 210
use FILL  FILL_9
timestamp 1739819275
transform 1 0 872 0 -1 1810
box -16 -6 32 210
use INVX1  INVX1_6
timestamp 1739819275
transform 1 0 888 0 -1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_6
timestamp 1739819275
transform -1 0 1096 0 -1 1810
box -16 -6 64 210
use OAI21X1  OAI21X1_5
timestamp 1739819275
transform -1 0 1048 0 -1 1810
box -16 -6 68 210
use OAI21X1  OAI21X1_4
timestamp 1739819275
transform 1 0 920 0 -1 1810
box -16 -6 68 210
use AND2X2  AND2X2_0
timestamp 1739819275
transform -1 0 1160 0 -1 1810
box -16 -6 80 210
use FILL  FILL_8
timestamp 1739819275
transform 1 0 1256 0 -1 1810
box -16 -6 32 210
use BUFX2  BUFX2_7
timestamp 1739819275
transform 1 0 1208 0 -1 1810
box -10 -6 56 210
use NOR2X1  NOR2X1_5
timestamp 1739819275
transform -1 0 1208 0 -1 1810
box -16 -6 64 210
use DFFSR  DFFSR_3
timestamp 1739819275
transform 1 0 1272 0 -1 1810
box -16 -6 368 210
use FILL  FILL_7
timestamp 1739819275
transform 1 0 1896 0 -1 1810
box -16 -6 32 210
use BUFX2  BUFX2_6
timestamp 1739819275
transform 1 0 1816 0 -1 1810
box -10 -6 56 210
use INVX1  INVX1_5
timestamp 1739819275
transform -1 0 1896 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_4
timestamp 1739819275
transform 1 0 1688 0 -1 1810
box -18 -6 52 210
use AOI21X1  AOI21X1_3
timestamp 1739819275
transform -1 0 1688 0 -1 1810
box -14 -6 78 210
use DFFSR  DFFSR_2
timestamp 1739819275
transform 1 0 1912 0 -1 1810
box -16 -6 368 210
use MUX2X1  MUX2X1_0
timestamp 1739819275
transform 1 0 1720 0 -1 1810
box -10 -6 106 210
use FILL  FILL_6
timestamp 1739819275
transform -1 0 392 0 1 1810
box -16 -6 32 210
use INVX1  INVX1_3
timestamp 1739819275
transform 1 0 168 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_4
timestamp 1739819275
transform -1 0 120 0 1 1810
box -16 -6 64 210
use AOI21X1  AOI21X1_2
timestamp 1739819275
transform -1 0 264 0 1 1810
box -14 -6 78 210
use NAND2X1  NAND2X1_4
timestamp 1739819275
transform 1 0 328 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_3
timestamp 1739819275
transform -1 0 168 0 1 1810
box -16 -6 64 210
use OAI21X1  OAI21X1_3
timestamp 1739819275
transform 1 0 8 0 1 1810
box -16 -6 68 210
use NAND3X1  NAND3X1_0
timestamp 1739819275
transform -1 0 328 0 1 1810
box -16 -6 80 210
use BUFX2  BUFX2_5
timestamp 1739819275
transform -1 0 808 0 1 1810
box -10 -6 56 210
use NOR2X1  NOR2X1_3
timestamp 1739819275
transform 1 0 648 0 1 1810
box -16 -6 64 210
use NOR2X1  NOR2X1_2
timestamp 1739819275
transform -1 0 440 0 1 1810
box -16 -6 64 210
use AOI21X1  AOI21X1_1
timestamp 1739819275
transform 1 0 536 0 1 1810
box -14 -6 78 210
use NAND2X1  NAND2X1_2
timestamp 1739819275
transform -1 0 648 0 1 1810
box -16 -6 64 210
use OAI21X1  OAI21X1_2
timestamp 1739819275
transform 1 0 696 0 1 1810
box -16 -6 68 210
use OAI21X1  OAI21X1_1
timestamp 1739819275
transform -1 0 504 0 1 1810
box -16 -6 68 210
use INVX2  INVX2_0
timestamp 1739819275
transform 1 0 504 0 1 1810
box -18 -6 52 210
use FILL  FILL_5
timestamp 1739819275
transform -1 0 872 0 1 1810
box -16 -6 32 210
use BUFX2  BUFX2_4
timestamp 1739819275
transform -1 0 1144 0 1 1810
box -10 -6 56 210
use INVX1  INVX1_2
timestamp 1739819275
transform -1 0 1096 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_1
timestamp 1739819275
transform -1 0 968 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_1
timestamp 1739819275
transform 1 0 968 0 1 1810
box -16 -6 64 210
use DFFSR  DFFSR_1
timestamp 1739819275
transform -1 0 1496 0 1 1810
box -16 -6 368 210
use NAND2X1  NAND2X1_1
timestamp 1739819275
transform -1 0 1064 0 1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_0
timestamp 1739819275
transform 1 0 808 0 1 1810
box -16 -6 64 210
use OAI21X1  OAI21X1_0
timestamp 1739819275
transform -1 0 936 0 1 1810
box -16 -6 68 210
use FILL  FILL_4
timestamp 1739819275
transform 1 0 1496 0 1 1810
box -16 -6 32 210
use BUFX2  BUFX2_3
timestamp 1739819275
transform 1 0 1512 0 1 1810
box -10 -6 56 210
use BUFX2  BUFX2_2
timestamp 1739819275
transform -1 0 1608 0 1 1810
box -10 -6 56 210
use DFFSR  DFFSR_0
timestamp 1739819275
transform 1 0 1608 0 1 1810
box -16 -6 368 210
use FILL  FILL_3
timestamp 1739819275
transform 1 0 2248 0 1 1810
box -16 -6 32 210
use FILL  FILL_2
timestamp 1739819275
transform 1 0 2232 0 1 1810
box -16 -6 32 210
use FILL  FILL_1
timestamp 1739819275
transform 1 0 2216 0 1 1810
box -16 -6 32 210
use FILL  FILL_0
timestamp 1739819275
transform 1 0 1960 0 1 1810
box -16 -6 32 210
use BUFX2  BUFX2_1
timestamp 1739819275
transform 1 0 2168 0 1 1810
box -10 -6 56 210
use BUFX2  BUFX2_0
timestamp 1739819275
transform 1 0 1976 0 1 1810
box -10 -6 56 210
use INVX1  INVX1_0
timestamp 1739819275
transform -1 0 2168 0 1 1810
box -18 -6 52 210
use NOR2X1  NOR2X1_0
timestamp 1739819275
transform -1 0 2136 0 1 1810
box -16 -6 64 210
use AOI21X1  AOI21X1_0
timestamp 1739819275
transform -1 0 2088 0 1 1810
box -14 -6 78 210
<< labels >>
flabel metal4 416 -36 416 -36 7 FreeSans 30 270 0 0 vdd
flabel metal4 880 -36 880 -36 7 FreeSans 30 270 0 0 gnd
flabel metal2 944 -20 944 -20 7 FreeSans 30 270 0 0 clock
flabel metal2 1072 -20 1072 -20 7 FreeSans 30 270 0 0 reset
flabel metal2 624 -20 624 -20 7 FreeSans 30 270 0 0 start
flabel metal2 2112 2040 2112 2040 3 FreeSans 30 90 0 0 N[0]
flabel metal2 656 2040 656 2040 3 FreeSans 30 90 0 0 N[1]
flabel metal2 624 2040 624 2040 3 FreeSans 30 90 0 0 N[2]
flabel metal2 560 2040 560 2040 3 FreeSans 30 90 0 0 N[3]
flabel metal2 448 2040 448 2040 3 FreeSans 30 90 0 0 N[4]
flabel metal3 -16 1880 -16 1880 7 FreeSans 30 0 0 0 N[5]
flabel metal3 -16 1920 -16 1920 7 FreeSans 30 0 0 0 N[6]
flabel metal3 -16 900 -16 900 7 FreeSans 30 0 0 0 N[7]
flabel metal3 -16 940 -16 940 7 FreeSans 30 0 0 0 N[8]
flabel metal3 2288 1900 2288 1900 3 FreeSans 30 0 0 0 dp[0]
flabel metal3 2288 700 2288 700 3 FreeSans 30 0 0 0 dp[1]
flabel metal2 1536 -20 1536 -20 7 FreeSans 30 270 0 0 dp[2]
flabel metal3 2288 300 2288 300 3 FreeSans 30 0 0 0 dp[3]
flabel metal2 1360 -20 1360 -20 7 FreeSans 30 270 0 0 dp[4]
flabel metal3 2288 740 2288 740 3 FreeSans 30 0 0 0 dp[5]
flabel metal2 992 -20 992 -20 7 FreeSans 30 270 0 0 dp[6]
flabel metal3 2288 1500 2288 1500 3 FreeSans 30 0 0 0 dp[7]
flabel metal2 2000 2040 2000 2040 3 FreeSans 30 90 0 0 dp[8]
flabel metal3 -16 500 -16 500 7 FreeSans 30 0 0 0 done
flabel metal2 1232 2040 1232 2040 3 FreeSans 30 90 0 0 counter[0]
flabel metal2 1120 2040 1120 2040 3 FreeSans 30 90 0 0 counter[1]
flabel metal2 784 2040 784 2040 3 FreeSans 30 90 0 0 counter[2]
flabel metal3 -16 1300 -16 1300 7 FreeSans 30 0 0 0 counter[3]
flabel metal3 -16 1500 -16 1500 7 FreeSans 30 0 0 0 counter[4]
flabel metal3 -16 1100 -16 1100 7 FreeSans 30 0 0 0 counter[5]
flabel metal3 -16 700 -16 700 7 FreeSans 30 0 0 0 counter[6]
flabel metal3 -16 740 -16 740 7 FreeSans 30 0 0 0 counter[7]
flabel metal3 2288 1100 2288 1100 3 FreeSans 30 0 0 0 sr[0]
flabel metal2 1728 -20 1728 -20 7 FreeSans 30 270 0 0 sr[1]
flabel metal3 2288 100 2288 100 3 FreeSans 30 0 0 0 sr[2]
flabel metal2 1616 -20 1616 -20 7 FreeSans 30 270 0 0 sr[3]
flabel metal3 2288 1300 2288 1300 3 FreeSans 30 0 0 0 sr[4]
flabel metal2 1536 2040 1536 2040 3 FreeSans 30 90 0 0 sr[5]
flabel metal2 1840 2040 1840 2040 3 FreeSans 30 90 0 0 sr[6]
flabel metal2 1584 2040 1584 2040 3 FreeSans 30 90 0 0 sr[7]
<< end >>

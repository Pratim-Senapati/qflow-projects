magic
tech scmos
magscale 1 2
timestamp 1744230924
<< metal1 >>
rect 2904 4206 2910 4214
rect 2918 4206 2924 4214
rect 2932 4206 2938 4214
rect 2946 4206 2952 4214
rect 93 4157 108 4163
rect 1460 4156 1468 4164
rect 61 4137 83 4143
rect 100 4137 131 4143
rect 301 4137 339 4143
rect 1348 4137 1395 4143
rect 189 4117 227 4123
rect 221 4097 227 4117
rect 253 4117 307 4123
rect 1693 4123 1699 4143
rect 1837 4143 1843 4163
rect 1853 4157 1891 4163
rect 2116 4157 2131 4163
rect 3997 4157 4012 4163
rect 1828 4137 1843 4143
rect 1940 4137 1971 4143
rect 2132 4137 2147 4143
rect 2685 4137 2700 4143
rect 3908 4137 3923 4143
rect 4372 4137 4387 4143
rect 4980 4137 4995 4143
rect 1693 4117 1724 4123
rect 2173 4123 2179 4136
rect 2157 4117 2179 4123
rect 2269 4117 2284 4123
rect 2701 4117 2732 4123
rect 356 4096 364 4104
rect 1036 4103 1044 4108
rect 1021 4097 1044 4103
rect 2701 4097 2707 4117
rect 3437 4117 3452 4123
rect 3533 4117 3548 4123
rect 3940 4117 3955 4123
rect 4420 4117 4467 4123
rect 3853 4097 3868 4103
rect 4317 4097 4332 4103
rect 4925 4097 4940 4103
rect 1268 4076 1272 4084
rect 1540 4076 1544 4084
rect 1352 4006 1358 4014
rect 1366 4006 1372 4014
rect 1380 4006 1386 4014
rect 1394 4006 1400 4014
rect 4440 4006 4446 4014
rect 4454 4006 4460 4014
rect 4468 4006 4474 4014
rect 4482 4006 4488 4014
rect 3012 3976 3014 3984
rect 1796 3956 1798 3964
rect 2356 3956 2358 3964
rect 1412 3936 1416 3944
rect 3284 3937 3299 3943
rect 61 3917 99 3923
rect 141 3917 179 3923
rect 189 3917 220 3923
rect 404 3916 412 3924
rect 253 3903 259 3916
rect 253 3897 275 3903
rect 285 3897 323 3903
rect 845 3903 851 3923
rect 1037 3917 1059 3923
rect 1092 3917 1107 3923
rect 781 3897 819 3903
rect 845 3897 883 3903
rect 1060 3897 1075 3903
rect 1732 3897 1747 3903
rect 1821 3903 1827 3923
rect 1933 3917 1948 3923
rect 2221 3917 2252 3923
rect 2381 3904 2387 3923
rect 3069 3917 3084 3923
rect 4365 3917 4380 3923
rect 4733 3917 4748 3923
rect 1821 3897 1859 3903
rect 2340 3897 2355 3903
rect 2388 3897 2419 3903
rect 2756 3897 2787 3903
rect 3124 3897 3155 3903
rect 3597 3897 3619 3903
rect 4125 3897 4140 3903
rect 4820 3897 4835 3903
rect 509 3877 540 3883
rect 557 3877 595 3883
rect 589 3857 595 3877
rect 644 3877 659 3883
rect 909 3877 924 3883
rect 957 3877 995 3883
rect 1012 3877 1027 3883
rect 1021 3857 1027 3877
rect 2061 3877 2115 3883
rect 2317 3877 2339 3883
rect 2484 3877 2515 3883
rect 2141 3857 2179 3863
rect 2509 3857 2515 3877
rect 2653 3877 2691 3883
rect 3188 3877 3203 3883
rect 3492 3877 3507 3883
rect 4788 3877 4803 3883
rect 3597 3857 3612 3863
rect 244 3836 246 3844
rect 938 3836 940 3844
rect 1524 3836 1528 3844
rect 1924 3836 1926 3844
rect 2596 3836 2600 3844
rect 2730 3836 2732 3844
rect 3098 3836 3100 3844
rect 4356 3836 4358 3844
rect 4906 3836 4908 3844
rect 2904 3806 2910 3814
rect 2918 3806 2924 3814
rect 2932 3806 2938 3814
rect 2946 3806 2952 3814
rect 1988 3776 1990 3784
rect 2340 3776 2344 3784
rect 1901 3743 1907 3763
rect 1924 3756 1932 3764
rect 1693 3737 1731 3743
rect 1821 3737 1875 3743
rect 1901 3737 1916 3743
rect 45 3717 83 3723
rect 45 3697 51 3717
rect 109 3723 115 3736
rect 109 3717 131 3723
rect 237 3717 252 3723
rect 413 3717 451 3723
rect 413 3697 419 3717
rect 1965 3723 1971 3743
rect 2004 3737 2019 3743
rect 2029 3737 2067 3743
rect 2260 3737 2275 3743
rect 2580 3737 2595 3743
rect 2989 3737 3020 3743
rect 3709 3743 3715 3763
rect 3709 3737 3747 3743
rect 4093 3737 4108 3743
rect 5332 3737 5347 3743
rect 5453 3737 5468 3743
rect 1933 3717 1971 3723
rect 2116 3717 2147 3723
rect 2157 3717 2195 3723
rect 2413 3717 2444 3723
rect 1636 3696 1640 3704
rect 2109 3697 2124 3703
rect 2157 3697 2163 3717
rect 2772 3717 2819 3723
rect 2845 3717 2883 3723
rect 2845 3697 2851 3717
rect 2900 3717 2963 3723
rect 3037 3717 3075 3723
rect 3181 3717 3196 3723
rect 3373 3717 3388 3723
rect 3597 3717 3628 3723
rect 3812 3717 3843 3723
rect 4068 3717 4083 3723
rect 4468 3717 4515 3723
rect 4877 3697 4892 3703
rect 20 3677 35 3683
rect 138 3676 140 3684
rect 1012 3676 1018 3684
rect 2084 3676 2086 3684
rect 2554 3676 2556 3684
rect 3802 3676 3804 3684
rect 2666 3636 2668 3644
rect 3076 3636 3078 3644
rect 3690 3636 3692 3644
rect 1352 3606 1358 3614
rect 1366 3606 1372 3614
rect 1380 3606 1386 3614
rect 1394 3606 1400 3614
rect 4440 3606 4446 3614
rect 4454 3606 4460 3614
rect 4468 3606 4474 3614
rect 4482 3606 4488 3614
rect 2692 3556 2696 3564
rect 3258 3556 3260 3564
rect 3316 3537 3331 3543
rect 4852 3536 4858 3544
rect 36 3516 44 3524
rect 280 3516 284 3524
rect 2004 3516 2014 3524
rect 2788 3516 2796 3524
rect 68 3497 83 3503
rect 77 3477 83 3497
rect 1933 3497 1964 3503
rect 2125 3497 2163 3503
rect 2205 3497 2227 3503
rect 2221 3484 2227 3497
rect 2292 3497 2355 3503
rect 2484 3497 2515 3503
rect 2813 3503 2819 3523
rect 4301 3504 4307 3523
rect 2772 3497 2787 3503
rect 2813 3497 2851 3503
rect 3156 3497 3187 3503
rect 3268 3497 3299 3503
rect 3652 3497 3667 3503
rect 4132 3497 4147 3503
rect 4180 3497 4211 3503
rect 4221 3497 4268 3503
rect 4308 3497 4339 3503
rect 317 3477 332 3483
rect 605 3477 620 3483
rect 772 3477 803 3483
rect 829 3477 867 3483
rect 925 3477 948 3483
rect 669 3457 707 3463
rect 717 3457 732 3463
rect 829 3457 835 3477
rect 940 3472 948 3477
rect 3069 3477 3123 3483
rect 3885 3477 3907 3483
rect 4365 3477 4380 3483
rect 4621 3477 4636 3483
rect 4644 3477 4659 3483
rect 4692 3477 4707 3483
rect 2973 3457 3011 3463
rect 3140 3457 3155 3463
rect 260 3436 264 3444
rect 1272 3436 1276 3444
rect 1357 3437 1404 3443
rect 1480 3436 1484 3444
rect 2260 3436 2264 3444
rect 2410 3436 2412 3444
rect 4564 3436 4566 3444
rect 4740 3436 4744 3444
rect 2904 3406 2910 3414
rect 2918 3406 2924 3414
rect 2932 3406 2938 3414
rect 2946 3406 2952 3414
rect 836 3376 838 3384
rect 2340 3376 2344 3384
rect 2717 3357 2732 3363
rect 2893 3357 2979 3363
rect 621 3337 643 3343
rect 1053 3337 1068 3343
rect 1245 3337 1260 3343
rect 1533 3337 1548 3343
rect 1604 3337 1619 3343
rect 2829 3337 2867 3343
rect 4429 3337 4476 3343
rect 4685 3337 4700 3343
rect 5821 3337 5852 3343
rect 429 3317 444 3323
rect 845 3317 883 3323
rect 557 3297 579 3303
rect 845 3297 851 3317
rect 916 3317 931 3323
rect 941 3317 956 3323
rect 1005 3317 1020 3323
rect 1069 3317 1100 3323
rect 1140 3317 1155 3323
rect 1236 3317 1283 3323
rect 1293 3317 1331 3323
rect 1357 3317 1388 3323
rect 900 3297 915 3303
rect 1204 3296 1214 3304
rect 1325 3297 1331 3317
rect 1684 3317 1699 3323
rect 1709 3317 1784 3323
rect 2196 3317 2227 3323
rect 2740 3317 2771 3323
rect 3165 3317 3203 3323
rect 3876 3317 3923 3323
rect 4013 3317 4028 3323
rect 4621 3317 4659 3323
rect 1661 3297 1683 3303
rect 2516 3297 2531 3303
rect 2573 3297 2595 3303
rect 3053 3297 3091 3303
rect 3108 3297 3123 3303
rect 4653 3297 4659 3317
rect 4692 3317 4723 3323
rect 4829 3317 4860 3323
rect 4669 3297 4684 3303
rect 474 3276 476 3284
rect 2493 3277 2540 3283
rect 3028 3276 3030 3284
rect 4372 3276 4376 3284
rect 2772 3256 2774 3264
rect 778 3236 780 3244
rect 1002 3236 1004 3244
rect 1476 3236 1480 3244
rect 2442 3236 2444 3244
rect 3268 3236 3272 3244
rect 3780 3236 3782 3244
rect 4564 3236 4566 3244
rect 1352 3206 1358 3214
rect 1366 3206 1372 3214
rect 1380 3206 1386 3214
rect 1394 3206 1400 3214
rect 4440 3206 4446 3214
rect 4454 3206 4460 3214
rect 4468 3206 4474 3214
rect 4482 3206 4488 3214
rect 4692 3176 4696 3184
rect 1204 3136 1206 3144
rect 189 3097 204 3103
rect 461 3103 467 3123
rect 484 3116 492 3124
rect 893 3117 915 3123
rect 1380 3117 1411 3123
rect 429 3097 467 3103
rect 516 3097 531 3103
rect 61 3077 76 3083
rect 525 3077 531 3097
rect 772 3097 787 3103
rect 1037 3097 1068 3103
rect 1165 3097 1203 3103
rect 1517 3103 1523 3123
rect 2308 3116 2316 3124
rect 3805 3104 3811 3123
rect 4333 3117 4355 3123
rect 1485 3097 1523 3103
rect 1549 3097 1564 3103
rect 2269 3097 2284 3103
rect 2381 3097 2396 3103
rect 2461 3097 2483 3103
rect 2541 3097 2595 3103
rect 2653 3097 2668 3103
rect 669 3077 684 3083
rect 932 3077 947 3083
rect 1565 3077 1580 3083
rect 1620 3077 1635 3083
rect 1661 3077 1715 3083
rect 1725 3077 1747 3083
rect 77 3057 83 3076
rect 1725 3064 1731 3077
rect 2333 3077 2355 3083
rect 2669 3083 2675 3096
rect 3316 3097 3347 3103
rect 3364 3097 3411 3103
rect 3444 3097 3475 3103
rect 3540 3097 3587 3103
rect 3764 3097 3779 3103
rect 3773 3084 3779 3097
rect 3812 3097 3843 3103
rect 3972 3097 3987 3103
rect 4356 3097 4371 3103
rect 4557 3103 4563 3123
rect 4404 3097 4435 3103
rect 4525 3097 4563 3103
rect 5380 3097 5395 3103
rect 2580 3077 2595 3083
rect 2669 3077 2691 3083
rect 2908 3077 2924 3083
rect 3197 3077 3212 3083
rect 3261 3077 3299 3083
rect 3501 3077 3523 3083
rect 3533 3077 3548 3083
rect 93 3057 131 3063
rect 212 3057 227 3063
rect 1677 3057 1692 3063
rect 3533 3057 3539 3077
rect 3933 3077 3955 3083
rect 4292 3077 4323 3083
rect 4397 3077 4412 3083
rect 4317 3057 4323 3077
rect 4644 3077 4659 3083
rect 4637 3057 4643 3076
rect 330 3036 332 3044
rect 564 3036 568 3044
rect 650 3036 652 3044
rect 1290 3036 1292 3044
rect 3700 3036 3704 3044
rect 4260 3036 4262 3044
rect 4445 3037 4492 3043
rect 2904 3006 2910 3014
rect 2918 3006 2924 3014
rect 2932 3006 2938 3014
rect 2946 3006 2952 3014
rect 4884 2976 4888 2984
rect 1149 2957 1171 2963
rect 1684 2957 1699 2963
rect 804 2937 819 2943
rect 1309 2937 1347 2943
rect 1540 2937 1555 2943
rect 1725 2937 1756 2943
rect 1789 2943 1795 2956
rect 1789 2937 1811 2943
rect 1980 2943 1988 2948
rect 109 2917 124 2923
rect 292 2917 323 2923
rect 420 2917 435 2923
rect 541 2917 579 2923
rect 605 2917 652 2923
rect 253 2897 275 2903
rect 573 2897 579 2917
rect 685 2917 723 2923
rect 685 2897 691 2917
rect 765 2917 803 2923
rect 916 2917 963 2923
rect 1037 2917 1068 2923
rect 1380 2917 1459 2923
rect 1869 2923 1875 2943
rect 1965 2937 1988 2943
rect 3149 2937 3171 2943
rect 3292 2943 3300 2948
rect 3261 2937 3300 2943
rect 3965 2937 3987 2943
rect 5773 2937 5788 2943
rect 1860 2917 1875 2923
rect 2468 2917 2515 2923
rect 3044 2917 3091 2923
rect 3197 2917 3235 2923
rect 4084 2917 4099 2923
rect 4509 2917 4547 2923
rect 5325 2917 5362 2923
rect 1117 2897 1132 2903
rect 1373 2897 1379 2916
rect 1620 2896 1628 2904
rect 1645 2897 1667 2903
rect 4061 2897 4083 2903
rect 5700 2897 5715 2903
rect 1908 2876 1912 2884
rect 3908 2876 3912 2884
rect 4612 2876 4614 2884
rect 5238 2876 5244 2884
rect 5837 2877 5852 2883
rect 602 2856 604 2864
rect 1092 2856 1094 2864
rect 4372 2856 4376 2864
rect 106 2836 108 2844
rect 660 2836 662 2844
rect 1352 2806 1358 2814
rect 1366 2806 1372 2814
rect 1380 2806 1386 2814
rect 1394 2806 1400 2814
rect 4440 2806 4446 2814
rect 4454 2806 4460 2814
rect 4468 2806 4474 2814
rect 4482 2806 4488 2814
rect 4552 2776 4556 2784
rect 196 2737 211 2743
rect 2212 2736 2216 2744
rect 2605 2737 2620 2743
rect 3652 2736 3656 2744
rect 4132 2737 4147 2743
rect 1524 2716 1532 2724
rect 253 2697 268 2703
rect 541 2697 556 2703
rect 692 2697 707 2703
rect 1236 2697 1267 2703
rect 1533 2697 1580 2703
rect 1645 2697 1683 2703
rect 1677 2684 1683 2697
rect 1741 2703 1747 2723
rect 1709 2697 1747 2703
rect 1853 2697 1868 2703
rect 2045 2697 2060 2703
rect 2461 2703 2467 2723
rect 2445 2697 2467 2703
rect 269 2677 291 2683
rect 285 2664 291 2677
rect 420 2677 451 2683
rect 468 2677 499 2683
rect 1028 2677 1043 2683
rect 1053 2677 1091 2683
rect 1149 2677 1164 2683
rect 1053 2664 1059 2677
rect 1229 2677 1244 2683
rect 1357 2677 1443 2683
rect 2285 2683 2291 2696
rect 2445 2684 2451 2697
rect 2516 2697 2531 2703
rect 3044 2697 3075 2703
rect 3124 2697 3155 2703
rect 3348 2697 3363 2703
rect 3716 2697 3747 2703
rect 3757 2697 3795 2703
rect 4413 2697 4444 2703
rect 5524 2697 5539 2703
rect 2269 2677 2291 2683
rect 2333 2677 2371 2683
rect 2333 2657 2339 2677
rect 2628 2677 2643 2683
rect 2685 2677 2707 2683
rect 2964 2677 3027 2683
rect 3037 2677 3052 2683
rect 3037 2657 3043 2677
rect 3092 2677 3107 2683
rect 3268 2677 3283 2683
rect 4013 2677 4028 2683
rect 5837 2677 5852 2683
rect 4068 2657 4083 2663
rect 628 2636 632 2644
rect 740 2636 742 2644
rect 920 2636 924 2644
rect 2740 2636 2744 2644
rect 2884 2636 2888 2644
rect 3322 2636 3324 2644
rect 2904 2606 2910 2614
rect 2918 2606 2924 2614
rect 2932 2606 2938 2614
rect 2946 2606 2952 2614
rect 2900 2577 2915 2583
rect 3300 2576 3302 2584
rect 4906 2576 4908 2584
rect 5096 2576 5100 2584
rect 5208 2576 5212 2584
rect 5320 2576 5324 2584
rect 173 2537 204 2543
rect 445 2537 460 2543
rect 493 2543 499 2556
rect 493 2537 515 2543
rect 717 2537 748 2543
rect 813 2543 819 2563
rect 1236 2557 1251 2563
rect 3540 2557 3555 2563
rect 4957 2557 4988 2563
rect 788 2537 803 2543
rect 813 2537 828 2543
rect 1428 2537 1443 2543
rect 1876 2537 1891 2543
rect 3261 2537 3276 2543
rect 3316 2537 3331 2543
rect 3389 2537 3427 2543
rect 3508 2537 3523 2543
rect 4765 2537 4803 2543
rect 4941 2543 4947 2556
rect 4925 2537 4947 2543
rect 5005 2537 5020 2543
rect 45 2517 83 2523
rect 77 2497 83 2517
rect 317 2517 332 2523
rect 724 2517 739 2523
rect 820 2517 851 2523
rect 1213 2523 1219 2536
rect 1213 2517 1235 2523
rect 1581 2517 1612 2523
rect 141 2497 156 2503
rect 877 2497 899 2503
rect 948 2497 963 2503
rect 1069 2497 1091 2503
rect 1581 2497 1587 2517
rect 1741 2517 1756 2523
rect 1853 2517 1868 2523
rect 1908 2517 1923 2523
rect 1940 2517 1955 2523
rect 2845 2517 2892 2523
rect 3309 2517 3324 2523
rect 1652 2497 1667 2503
rect 1677 2497 1715 2503
rect 3309 2497 3315 2517
rect 3572 2517 3603 2523
rect 4100 2517 4115 2523
rect 4724 2517 4739 2523
rect 5037 2523 5043 2543
rect 5252 2537 5267 2543
rect 5837 2537 5852 2543
rect 5028 2517 5043 2523
rect 3348 2496 3356 2504
rect 4692 2497 4723 2503
rect 4852 2496 4860 2504
rect 916 2477 931 2483
rect 1044 2476 1046 2484
rect 1940 2477 1955 2483
rect 3140 2476 3144 2484
rect 378 2436 380 2444
rect 548 2436 552 2444
rect 1316 2436 1320 2444
rect 1476 2436 1480 2444
rect 1850 2436 1852 2444
rect 1352 2406 1358 2414
rect 1366 2406 1372 2414
rect 1380 2406 1386 2414
rect 1394 2406 1400 2414
rect 4440 2406 4446 2414
rect 4454 2406 4460 2414
rect 4468 2406 4474 2414
rect 4482 2406 4488 2414
rect 4330 2376 4332 2384
rect 5805 2377 5852 2383
rect 852 2336 856 2344
rect 2582 2336 2588 2344
rect 2970 2336 2972 2344
rect 4205 2337 4220 2343
rect 4436 2337 4515 2343
rect 4554 2336 4556 2344
rect 4856 2336 4860 2344
rect 1540 2316 1548 2324
rect 1565 2303 1571 2323
rect 1565 2297 1596 2303
rect 2948 2297 2963 2303
rect 2845 2277 2867 2283
rect 2877 2277 2956 2283
rect 3309 2277 3331 2283
rect 3341 2277 3363 2283
rect 3325 2264 3331 2277
rect 3820 2277 3844 2283
rect 4317 2283 4323 2303
rect 4532 2297 4547 2303
rect 5444 2297 5459 2303
rect 4204 2277 4227 2283
rect 4285 2277 4323 2283
rect 4621 2277 4636 2283
rect 4204 2272 4212 2277
rect 4676 2277 4691 2283
rect 2989 2257 3011 2263
rect 3028 2257 3043 2263
rect 4244 2257 4275 2263
rect 4525 2257 4540 2263
rect 356 2236 360 2244
rect 1444 2236 1448 2244
rect 3290 2236 3292 2244
rect 4602 2236 4604 2244
rect 2904 2206 2910 2214
rect 2918 2206 2924 2214
rect 2932 2206 2938 2214
rect 2946 2206 2952 2214
rect 3880 2176 3884 2184
rect 5096 2176 5100 2184
rect 5208 2176 5212 2184
rect 1757 2157 1779 2163
rect 1924 2157 1939 2163
rect 2260 2157 2275 2163
rect 2285 2157 2307 2163
rect 2749 2157 2771 2163
rect 2877 2157 2924 2163
rect 4660 2156 4668 2164
rect 1332 2137 1364 2143
rect 1757 2137 1772 2143
rect 1940 2137 1955 2143
rect 2285 2137 2300 2143
rect 2884 2137 2963 2143
rect 3677 2137 3699 2143
rect 3917 2137 3932 2143
rect 4637 2137 4652 2143
rect 4692 2137 4707 2143
rect 5028 2137 5043 2143
rect 5309 2137 5324 2143
rect 1421 2117 1436 2123
rect 1613 2117 1628 2123
rect 1805 2117 1836 2123
rect 1853 2117 1884 2123
rect 2237 2117 2268 2123
rect 2333 2117 2364 2123
rect 2381 2117 2428 2123
rect 2852 2117 2867 2123
rect 2973 2117 2996 2123
rect 2988 2114 2996 2117
rect 3949 2117 3964 2123
rect 4509 2117 4547 2123
rect 4708 2117 4723 2123
rect 4733 2117 4764 2123
rect 4797 2117 4828 2123
rect 5252 2117 5267 2123
rect 5325 2117 5363 2123
rect 5389 2123 5395 2143
rect 5380 2117 5395 2123
rect 3988 2096 3996 2104
rect 5357 2097 5388 2103
rect 1917 2077 1932 2083
rect 2166 2076 2172 2084
rect 2500 2076 2502 2084
rect 2797 2077 2812 2083
rect 3716 2076 3718 2084
rect 1988 2036 1990 2044
rect 1352 2006 1358 2014
rect 1366 2006 1372 2014
rect 1380 2006 1386 2014
rect 1394 2006 1400 2014
rect 4440 2006 4446 2014
rect 4454 2006 4460 2014
rect 4468 2006 4474 2014
rect 4482 2006 4488 2014
rect 2648 1976 2652 1984
rect 3268 1976 3272 1984
rect 3512 1976 3516 1984
rect 3940 1976 3942 1984
rect 4461 1977 4508 1983
rect 4712 1976 4716 1984
rect 5048 1976 5052 1984
rect 2026 1936 2028 1944
rect 3053 1937 3068 1943
rect 5293 1937 5324 1943
rect 788 1917 819 1923
rect 884 1917 899 1923
rect 77 1897 92 1903
rect 644 1897 675 1903
rect 909 1897 940 1903
rect 1021 1903 1027 1923
rect 1165 1917 1187 1923
rect 1908 1916 1916 1924
rect 1101 1903 1107 1916
rect 957 1897 995 1903
rect 1021 1897 1059 1903
rect 1069 1897 1107 1903
rect 1572 1897 1587 1903
rect 1725 1897 1756 1903
rect 1949 1903 1955 1923
rect 3028 1917 3043 1923
rect 1924 1897 1955 1903
rect 2180 1896 2184 1904
rect 2484 1897 2508 1903
rect 2525 1897 2547 1903
rect 3005 1897 3036 1903
rect 3740 1903 3748 1906
rect 3740 1897 3763 1903
rect 3853 1903 3859 1923
rect 4573 1917 4595 1923
rect 4813 1917 4835 1923
rect 3844 1897 3859 1903
rect 589 1877 627 1883
rect 845 1877 867 1883
rect 1140 1877 1155 1883
rect 1149 1857 1155 1877
rect 2093 1877 2115 1883
rect 2125 1877 2147 1883
rect 2125 1864 2131 1877
rect 2356 1876 2358 1884
rect 2692 1877 2707 1883
rect 3069 1877 3084 1883
rect 3165 1877 3180 1883
rect 3332 1877 3347 1883
rect 3389 1877 3411 1883
rect 3949 1883 3955 1903
rect 5277 1903 5283 1923
rect 5245 1897 5283 1903
rect 5588 1896 5592 1904
rect 3949 1877 3987 1883
rect 4909 1877 4947 1883
rect 5261 1877 5276 1883
rect 5428 1877 5443 1883
rect 5517 1877 5555 1883
rect 4061 1857 4076 1863
rect 570 1836 572 1844
rect 618 1836 620 1844
rect 1114 1836 1116 1844
rect 1194 1836 1196 1844
rect 1405 1837 1452 1843
rect 1962 1836 1964 1844
rect 2074 1836 2076 1844
rect 2904 1806 2910 1814
rect 2918 1806 2924 1814
rect 2932 1806 2938 1814
rect 2946 1806 2952 1814
rect 3844 1776 3846 1784
rect 4856 1776 4860 1784
rect 5092 1776 5094 1784
rect 701 1757 716 1763
rect 2492 1744 2500 1748
rect 253 1723 259 1743
rect 685 1737 700 1743
rect 733 1737 771 1743
rect 1940 1737 1955 1743
rect 2253 1737 2291 1743
rect 2772 1736 2774 1744
rect 253 1717 307 1723
rect 484 1717 515 1723
rect 708 1717 739 1723
rect 772 1717 787 1723
rect 1261 1717 1324 1723
rect 1933 1717 1964 1723
rect 1885 1697 1923 1703
rect 1933 1697 1939 1717
rect 2061 1717 2083 1723
rect 2141 1717 2156 1723
rect 3149 1723 3155 1743
rect 3197 1737 3212 1743
rect 3229 1737 3244 1743
rect 3581 1743 3587 1763
rect 3549 1737 3587 1743
rect 3709 1743 3715 1763
rect 5540 1757 5555 1763
rect 3668 1737 3715 1743
rect 4781 1737 4796 1743
rect 3117 1717 3155 1723
rect 3245 1717 3283 1723
rect 3293 1717 3347 1723
rect 3357 1717 3395 1723
rect 3245 1697 3251 1717
rect 3453 1717 3484 1723
rect 3629 1717 3667 1723
rect 4045 1717 4083 1723
rect 4157 1717 4195 1723
rect 3348 1696 3356 1704
rect 3949 1697 3964 1703
rect 4157 1697 4163 1717
rect 4324 1717 4339 1723
rect 4925 1717 4963 1723
rect 4973 1717 5011 1723
rect 5005 1697 5011 1717
rect 5236 1717 5267 1723
rect 5300 1717 5331 1723
rect 5404 1717 5420 1723
rect 5404 1712 5412 1717
rect 5645 1717 5660 1723
rect 328 1676 332 1684
rect 788 1676 790 1684
rect 2202 1676 2204 1684
rect 3046 1676 3052 1684
rect 5805 1677 5852 1683
rect 440 1656 444 1664
rect 1784 1656 1788 1664
rect 5274 1656 5276 1664
rect 1000 1636 1004 1644
rect 4042 1636 4044 1644
rect 1352 1606 1358 1614
rect 1366 1606 1372 1614
rect 1380 1606 1386 1614
rect 1394 1606 1400 1614
rect 4440 1606 4446 1614
rect 4454 1606 4460 1614
rect 4468 1606 4474 1614
rect 4482 1606 4488 1614
rect 420 1576 422 1584
rect 3562 1576 3564 1584
rect 5592 1576 5596 1584
rect 744 1536 748 1544
rect 1076 1537 1091 1543
rect 2392 1536 2396 1544
rect 3078 1536 3084 1544
rect 445 1517 483 1523
rect 2493 1517 2515 1523
rect 564 1497 579 1503
rect 589 1497 643 1503
rect 941 1497 963 1503
rect 1037 1503 1043 1516
rect 980 1497 1011 1503
rect 1021 1497 1043 1503
rect 2093 1503 2099 1516
rect 2029 1497 2099 1503
rect 2820 1496 2824 1504
rect 3533 1503 3539 1523
rect 3844 1516 3852 1524
rect 4349 1517 4371 1523
rect 3501 1497 3539 1503
rect 3661 1497 3676 1503
rect 3764 1497 3779 1503
rect 4212 1497 4243 1503
rect 4637 1503 4643 1523
rect 5197 1517 5212 1523
rect 4605 1497 4643 1503
rect 4653 1497 4668 1503
rect 4788 1497 4803 1503
rect 5037 1497 5068 1503
rect 1220 1477 1251 1483
rect 1261 1477 1315 1483
rect 2324 1477 2339 1483
rect 2541 1477 2572 1483
rect 2596 1477 2611 1483
rect 1332 1456 1340 1464
rect 2605 1457 2611 1477
rect 3581 1477 3603 1483
rect 3965 1477 4003 1483
rect 4036 1477 4083 1483
rect 4292 1477 4307 1483
rect 4413 1477 4444 1483
rect 4477 1477 4531 1483
rect 4541 1477 4579 1483
rect 5197 1477 5219 1483
rect 5384 1477 5404 1483
rect 5524 1477 5539 1483
rect 2621 1457 2636 1463
rect 4100 1456 4108 1464
rect 1480 1436 1484 1444
rect 1928 1436 1932 1444
rect 2200 1436 2204 1444
rect 4004 1436 4006 1444
rect 5460 1436 5462 1444
rect 5821 1437 5836 1443
rect 2904 1406 2910 1414
rect 2918 1406 2924 1414
rect 2932 1406 2938 1414
rect 2946 1406 2952 1414
rect 442 1376 444 1384
rect 500 1376 502 1384
rect 612 1376 614 1384
rect 1290 1376 1292 1384
rect 3866 1376 3868 1384
rect 4020 1376 4022 1384
rect 4264 1376 4268 1384
rect 4756 1377 4771 1383
rect 5156 1376 5158 1384
rect 5348 1376 5350 1384
rect 5716 1376 5720 1384
rect 173 1357 211 1363
rect 308 1357 323 1363
rect 61 1337 92 1343
rect 189 1317 204 1323
rect 461 1323 467 1343
rect 1316 1337 1379 1343
rect 1805 1337 1843 1343
rect 397 1317 435 1323
rect 461 1317 499 1323
rect 509 1317 547 1323
rect 365 1297 380 1303
rect 429 1297 435 1317
rect 509 1304 515 1317
rect 797 1317 835 1323
rect 861 1317 899 1323
rect 829 1297 835 1317
rect 957 1317 995 1323
rect 1021 1317 1059 1323
rect 1133 1317 1148 1323
rect 989 1297 995 1317
rect 1053 1304 1059 1317
rect 1181 1317 1219 1323
rect 1245 1317 1260 1323
rect 1069 1297 1107 1303
rect 1213 1297 1219 1317
rect 1901 1317 1916 1323
rect 2013 1317 2035 1323
rect 2013 1304 2019 1317
rect 2125 1323 2131 1343
rect 2541 1343 2547 1363
rect 2596 1357 2611 1363
rect 4381 1344 4387 1363
rect 4397 1357 4483 1363
rect 4621 1357 4643 1363
rect 2541 1337 2579 1343
rect 2621 1337 2643 1343
rect 2797 1337 2812 1343
rect 2893 1337 2940 1343
rect 3469 1337 3484 1343
rect 2125 1317 2140 1323
rect 2173 1317 2211 1323
rect 1869 1297 1884 1303
rect 2205 1297 2211 1317
rect 2365 1317 2419 1323
rect 2589 1317 2627 1323
rect 2692 1317 2723 1323
rect 2829 1317 2867 1323
rect 3597 1323 3603 1343
rect 3613 1337 3651 1343
rect 3732 1337 3747 1343
rect 3837 1337 3852 1343
rect 3965 1337 4019 1343
rect 4052 1337 4099 1343
rect 4125 1337 4179 1343
rect 4365 1337 4380 1343
rect 5149 1337 5187 1343
rect 3588 1317 3603 1323
rect 3933 1317 3955 1323
rect 3933 1304 3939 1317
rect 4509 1317 4547 1323
rect 4557 1317 4588 1323
rect 4701 1317 4716 1323
rect 2724 1296 2732 1304
rect 3426 1296 3436 1304
rect 3629 1297 3644 1303
rect 3709 1297 3731 1303
rect 3844 1297 3859 1303
rect 4621 1297 4636 1303
rect 5213 1297 5251 1303
rect 5364 1297 5379 1303
rect 5444 1297 5459 1303
rect 20 1277 35 1283
rect 1734 1276 1740 1284
rect 2106 1276 2108 1284
rect 3320 1256 3324 1264
rect 116 1236 118 1244
rect 228 1236 230 1244
rect 714 1236 716 1244
rect 1018 1236 1020 1244
rect 1524 1236 1528 1244
rect 1940 1236 1942 1244
rect 2042 1236 2044 1244
rect 2234 1236 2236 1244
rect 2660 1236 2662 1244
rect 3016 1236 3020 1244
rect 5604 1236 5608 1244
rect 1352 1206 1358 1214
rect 1366 1206 1372 1214
rect 1380 1206 1386 1214
rect 1394 1206 1400 1214
rect 4440 1206 4446 1214
rect 4454 1206 4460 1214
rect 4468 1206 4474 1214
rect 4482 1206 4488 1214
rect 1188 1176 1190 1184
rect 2520 1176 2524 1184
rect 4170 1176 4172 1184
rect 1380 1157 1427 1163
rect 776 1136 780 1144
rect 1892 1137 1907 1143
rect 2888 1136 2892 1144
rect 5174 1136 5180 1144
rect 525 1117 563 1123
rect 2324 1116 2332 1124
rect 2621 1117 2659 1123
rect 3908 1116 3916 1124
rect 205 1097 220 1103
rect 285 1097 316 1103
rect 397 1097 428 1103
rect 589 1097 604 1103
rect 877 1097 892 1103
rect 1172 1097 1187 1103
rect 1261 1097 1276 1103
rect 1572 1097 1619 1103
rect 1748 1097 1763 1103
rect 1997 1097 2012 1103
rect 2356 1097 2387 1103
rect 3005 1097 3043 1103
rect 3524 1097 3539 1103
rect 3693 1097 3747 1103
rect 3853 1097 3868 1103
rect 3876 1097 3907 1103
rect 4029 1097 4051 1103
rect 4068 1097 4099 1103
rect 4109 1097 4124 1103
rect 4596 1097 4611 1103
rect 5556 1097 5571 1103
rect 317 1077 332 1083
rect 612 1077 627 1083
rect 637 1077 652 1083
rect 621 1057 627 1077
rect 692 1077 723 1083
rect 1149 1077 1171 1083
rect 1293 1077 1331 1083
rect 1437 1077 1475 1083
rect 1437 1064 1443 1077
rect 1853 1077 1884 1083
rect 2100 1077 2131 1083
rect 2701 1077 2716 1083
rect 4045 1077 4083 1083
rect 957 1057 988 1063
rect 1908 1057 1939 1063
rect 122 1036 124 1044
rect 916 1036 918 1044
rect 1540 1036 1544 1044
rect 5288 1036 5292 1044
rect 5400 1036 5404 1044
rect 2904 1006 2910 1014
rect 2918 1006 2924 1014
rect 2932 1006 2938 1014
rect 2946 1006 2952 1014
rect 874 976 876 984
rect 2708 976 2710 984
rect 2884 977 2931 983
rect 3736 976 3740 984
rect 4106 976 4108 984
rect 4493 977 4508 983
rect 4616 976 4620 984
rect 397 957 419 963
rect 397 937 412 943
rect 509 943 515 963
rect 584 956 588 964
rect 932 956 940 964
rect 1133 957 1148 963
rect 500 937 515 943
rect 989 937 1043 943
rect 1277 937 1331 943
rect 1517 937 1555 943
rect 1821 943 1827 963
rect 1837 957 1868 963
rect 1917 943 1923 963
rect 1789 937 1827 943
rect 1885 937 1923 943
rect 1933 937 1948 943
rect 2093 943 2099 963
rect 2084 937 2099 943
rect 2109 937 2147 943
rect 2397 937 2412 943
rect 2541 937 2556 943
rect 2772 937 2787 943
rect 2980 937 2995 943
rect 3005 937 3020 943
rect 3533 937 3580 943
rect 148 917 163 923
rect 173 917 204 923
rect 477 917 508 923
rect 701 917 732 923
rect 797 917 812 923
rect 941 917 956 923
rect 61 897 83 903
rect 429 897 451 903
rect 813 897 835 903
rect 852 897 867 903
rect 941 897 947 917
rect 1437 917 1452 923
rect 1997 917 2028 923
rect 2285 917 2323 923
rect 2420 917 2451 923
rect 2813 917 2828 923
rect 3677 924 3683 943
rect 3885 937 3900 943
rect 4125 937 4140 943
rect 4532 937 4563 943
rect 4856 937 4883 943
rect 5292 937 5316 943
rect 5805 937 5852 943
rect 3645 917 3676 923
rect 4013 917 4051 923
rect 4728 917 4780 923
rect 1165 897 1187 903
rect 2612 896 2616 904
rect 2717 897 2739 903
rect 3028 897 3059 903
rect 3613 897 3635 903
rect 4212 896 4220 904
rect 4797 897 4819 903
rect 1133 877 1148 883
rect 2845 877 2908 883
rect 3446 876 3452 884
rect 5670 876 5676 884
rect 474 856 476 864
rect 1434 836 1436 844
rect 2058 836 2060 844
rect 1352 806 1358 814
rect 1366 806 1372 814
rect 1380 806 1386 814
rect 1394 806 1400 814
rect 4440 806 4446 814
rect 4454 806 4460 814
rect 4468 806 4474 814
rect 4482 806 4488 814
rect 1764 776 1766 784
rect 1850 776 1852 784
rect 1946 776 1948 784
rect 2004 776 2006 784
rect 2762 776 2764 784
rect 3924 776 3926 784
rect 4680 776 4684 784
rect 5290 776 5292 784
rect 2292 736 2294 744
rect 308 716 316 724
rect 477 717 499 723
rect 644 716 652 724
rect 893 717 915 723
rect 1060 716 1068 724
rect 516 697 531 703
rect 564 697 579 703
rect 628 697 643 703
rect 1277 703 1283 723
rect 1293 717 1331 723
rect 1789 717 1804 723
rect 2045 717 2083 723
rect 2100 716 2108 724
rect 2317 717 2339 723
rect 2973 717 2995 723
rect 3133 717 3155 723
rect 1245 697 1283 703
rect 1357 697 1436 703
rect 2109 697 2124 703
rect 2276 697 2291 703
rect 2653 697 2684 703
rect 2996 697 3011 703
rect 3949 703 3955 723
rect 4861 717 4883 723
rect 5021 717 5043 723
rect 3885 697 3923 703
rect 3949 697 3987 703
rect 4093 697 4124 703
rect 4173 697 4195 703
rect 4388 697 4435 703
rect 4829 697 4844 703
rect 4884 697 4899 703
rect 4932 697 4963 703
rect 5044 697 5059 703
rect 5261 703 5267 723
rect 5204 697 5219 703
rect 5229 697 5267 703
rect 5364 697 5379 703
rect 109 677 124 683
rect 221 677 243 683
rect 397 677 428 683
rect 541 677 572 683
rect 605 677 620 683
rect 557 657 595 663
rect 605 657 611 677
rect 1117 677 1155 683
rect 1149 657 1155 677
rect 2173 677 2227 683
rect 2781 677 2796 683
rect 2813 677 2828 683
rect 2916 677 2956 683
rect 3309 677 3324 683
rect 2349 657 2364 663
rect 2445 657 2460 663
rect 3172 657 3187 663
rect 3284 657 3299 663
rect 3309 657 3315 677
rect 3540 676 3542 684
rect 3732 676 3734 684
rect 3804 677 3827 683
rect 3804 672 3812 677
rect 4020 677 4035 683
rect 4045 677 4083 683
rect 4285 677 4339 683
rect 4516 677 4547 683
rect 4813 677 4844 683
rect 5117 677 5148 683
rect 5837 677 5852 683
rect 3844 657 3875 663
rect 4260 656 4268 664
rect 52 636 56 644
rect 1012 636 1014 644
rect 1476 636 1480 644
rect 3384 636 3388 644
rect 2904 606 2910 614
rect 2918 606 2924 614
rect 2932 606 2938 614
rect 2946 606 2952 614
rect 2056 576 2060 584
rect 2472 576 2476 584
rect 3946 576 3948 584
rect 5192 576 5196 584
rect 1476 557 1491 563
rect 45 543 51 556
rect 45 537 67 543
rect 244 537 275 543
rect 372 537 387 543
rect 573 543 579 556
rect 557 537 579 543
rect 941 537 979 543
rect 996 537 1011 543
rect 1085 537 1100 543
rect 1325 543 1331 556
rect 1325 537 1395 543
rect 1540 537 1555 543
rect 2285 543 2291 563
rect 2813 557 2828 563
rect 2973 557 2995 563
rect 4797 557 4835 563
rect 4845 557 4860 563
rect 2285 537 2323 543
rect 2765 537 2780 543
rect 3021 537 3036 543
rect 3069 537 3084 543
rect 4205 537 4220 543
rect 4228 537 4243 543
rect 4621 537 4636 543
rect 4708 537 4739 543
rect 4957 537 4972 543
rect 5117 543 5123 556
rect 5069 537 5107 543
rect 5117 537 5139 543
rect 212 517 227 523
rect 349 517 371 523
rect 692 517 723 523
rect 1197 517 1219 523
rect 1533 517 1603 523
rect 2141 517 2211 523
rect 2221 517 2259 523
rect 2340 517 2371 523
rect 2749 517 2764 523
rect 3037 517 3052 523
rect 3309 517 3324 523
rect 3421 517 3459 523
rect 100 497 131 503
rect 1437 497 1459 503
rect 2372 496 2380 504
rect 3085 497 3107 503
rect 3453 497 3459 517
rect 4301 517 4371 523
rect 4509 517 4547 523
rect 3917 497 3939 503
rect 4397 497 4435 503
rect 4541 497 4547 517
rect 5309 517 5324 523
rect 3084 484 3092 488
rect 1720 476 1724 484
rect 3846 476 3852 484
rect 180 436 182 444
rect 820 436 822 444
rect 1028 436 1030 444
rect 1588 436 1592 444
rect 4372 436 4374 444
rect 1352 406 1358 414
rect 1366 406 1372 414
rect 1380 406 1386 414
rect 1394 406 1400 414
rect 4440 406 4446 414
rect 4454 406 4460 414
rect 4468 406 4474 414
rect 4482 406 4488 414
rect 1928 376 1932 384
rect 2692 376 2694 384
rect 2884 376 2886 384
rect 3002 376 3004 384
rect 3178 376 3180 384
rect 4196 376 4198 384
rect 4884 376 4886 384
rect 4954 376 4956 384
rect 5332 376 5336 384
rect 5700 376 5704 384
rect 349 303 355 323
rect 1700 316 1708 324
rect 349 297 387 303
rect 804 297 819 303
rect 957 297 1004 303
rect 1709 297 1756 303
rect 1805 303 1811 323
rect 2264 316 2268 324
rect 1773 297 1811 303
rect 2125 297 2163 303
rect 29 277 51 283
rect 260 277 275 283
rect 1725 277 1740 283
rect 2157 277 2163 297
rect 2413 283 2419 303
rect 2573 303 2579 316
rect 2557 297 2579 303
rect 2717 303 2723 323
rect 2964 317 2979 323
rect 2717 297 2755 303
rect 2772 297 2819 303
rect 2829 297 2860 303
rect 3069 297 3084 303
rect 3149 303 3155 323
rect 3117 297 3155 303
rect 3364 297 3395 303
rect 3501 303 3507 323
rect 3517 317 3532 323
rect 4269 317 4307 323
rect 4612 316 4620 324
rect 5533 317 5548 323
rect 3492 297 3507 303
rect 3860 297 3875 303
rect 4072 297 4124 303
rect 4228 297 4243 303
rect 4365 297 4387 303
rect 2356 277 2371 283
rect 2381 277 2419 283
rect 477 257 492 263
rect 1556 257 1587 263
rect 2365 257 2371 277
rect 2468 277 2515 283
rect 2605 277 2643 283
rect 2788 277 2803 283
rect 3405 277 3436 283
rect 3533 277 3548 283
rect 3597 277 3612 283
rect 3629 277 3651 283
rect 3981 277 4019 283
rect 4237 277 4243 297
rect 4381 284 4387 297
rect 4413 297 4492 303
rect 4868 297 4883 303
rect 5117 297 5139 303
rect 5156 297 5171 303
rect 5396 297 5411 303
rect 4301 277 4332 283
rect 4452 277 4499 283
rect 4509 277 4547 283
rect 4637 277 4675 283
rect 5213 277 5267 283
rect 5389 277 5404 283
rect 5421 277 5459 283
rect 3428 257 3443 263
rect 5453 257 5459 277
rect 68 236 70 244
rect 648 236 652 244
rect 1300 236 1304 244
rect 1480 236 1484 244
rect 1556 236 1558 244
rect 2180 236 2182 244
rect 4260 236 4262 244
rect 2904 206 2910 214
rect 2918 206 2924 214
rect 2932 206 2938 214
rect 2946 206 2952 214
rect 1880 176 1884 184
rect 2458 176 2460 184
rect 2888 176 2892 184
rect 3146 176 3148 184
rect 4088 176 4092 184
rect 4554 176 4556 184
rect 1652 157 1667 163
rect 1693 143 1699 163
rect 3226 156 3228 164
rect 5108 157 5123 163
rect 5341 144 5347 163
rect 1661 137 1699 143
rect 1789 137 1820 143
rect 2109 137 2147 143
rect 1469 117 1539 123
rect 1629 117 1651 123
rect 1965 117 2019 123
rect 2045 117 2083 123
rect 1565 97 1587 103
rect 2045 97 2051 117
rect 2157 117 2179 123
rect 2253 123 2259 143
rect 2301 137 2316 143
rect 2925 137 2972 143
rect 3997 137 4012 143
rect 4429 137 4460 143
rect 4484 137 4499 143
rect 2244 117 2259 123
rect 2484 117 2515 123
rect 3005 117 3043 123
rect 2173 97 2204 103
rect 2285 97 2307 103
rect 2589 97 2627 103
rect 3037 97 3043 117
rect 3341 117 3372 123
rect 4205 117 4243 123
rect 3117 97 3139 103
rect 4237 97 4243 117
rect 4573 123 4579 136
rect 4797 124 4803 143
rect 5085 137 5116 143
rect 5348 137 5379 143
rect 4573 117 4595 123
rect 4804 117 4835 123
rect 4845 117 4883 123
rect 4532 97 4547 103
rect 4760 96 4764 104
rect 4877 97 4883 117
rect 5229 117 5244 123
rect 5284 117 5315 123
rect 5325 117 5356 123
rect 4964 96 4972 104
rect 5229 97 5251 103
rect 232 76 236 84
rect 344 76 348 84
rect 2564 76 2566 84
rect 2712 76 2716 84
rect 4308 77 4323 83
rect 5821 77 5852 83
rect 2020 56 2022 64
rect 2392 56 2396 64
rect 1352 6 1358 14
rect 1366 6 1372 14
rect 1380 6 1386 14
rect 1394 6 1400 14
rect 4440 6 4446 14
rect 4454 6 4460 14
rect 4468 6 4474 14
rect 4482 6 4488 14
<< m2contact >>
rect 2910 4206 2918 4214
rect 2924 4206 2932 4214
rect 2938 4206 2946 4214
rect 396 4176 404 4184
rect 460 4176 468 4184
rect 2204 4176 2212 4184
rect 4604 4176 4612 4184
rect 108 4156 116 4164
rect 284 4156 292 4164
rect 1452 4156 1460 4164
rect 92 4136 100 4144
rect 172 4136 180 4144
rect 268 4136 276 4144
rect 444 4136 452 4144
rect 620 4136 628 4144
rect 812 4136 820 4144
rect 844 4136 852 4144
rect 972 4136 980 4144
rect 988 4136 996 4144
rect 1196 4136 1204 4144
rect 1228 4136 1236 4144
rect 1324 4136 1332 4144
rect 1340 4136 1348 4144
rect 1436 4136 1444 4144
rect 1484 4136 1492 4144
rect 1500 4136 1508 4144
rect 1596 4136 1604 4144
rect 1612 4136 1620 4144
rect 28 4116 36 4124
rect 44 4116 52 4124
rect 12 4096 20 4104
rect 204 4096 212 4104
rect 236 4116 244 4124
rect 316 4116 324 4124
rect 348 4116 356 4124
rect 428 4116 436 4124
rect 588 4118 596 4126
rect 780 4118 788 4126
rect 1100 4116 1108 4124
rect 1164 4118 1172 4126
rect 1420 4116 1428 4124
rect 1676 4116 1684 4124
rect 1708 4136 1716 4144
rect 1740 4136 1748 4144
rect 1820 4136 1828 4144
rect 1980 4156 1988 4164
rect 2028 4156 2036 4164
rect 2092 4156 2100 4164
rect 2108 4156 2116 4164
rect 2412 4156 2420 4164
rect 3724 4156 3732 4164
rect 4012 4156 4020 4164
rect 4188 4156 4196 4164
rect 4508 4156 4516 4164
rect 4796 4156 4804 4164
rect 5068 4156 5076 4164
rect 5292 4156 5300 4164
rect 5660 4156 5668 4164
rect 1916 4136 1924 4144
rect 1932 4136 1940 4144
rect 2124 4136 2132 4144
rect 2172 4136 2180 4144
rect 2668 4136 2676 4144
rect 2700 4136 2708 4144
rect 2716 4136 2724 4144
rect 2940 4136 2948 4144
rect 3020 4136 3028 4144
rect 3148 4136 3156 4144
rect 3404 4136 3412 4144
rect 3756 4136 3764 4144
rect 3900 4136 3908 4144
rect 3932 4136 3940 4144
rect 3980 4136 3988 4144
rect 4220 4136 4228 4144
rect 4364 4136 4372 4144
rect 4396 4136 4404 4144
rect 4492 4136 4500 4144
rect 4828 4136 4836 4144
rect 4972 4136 4980 4144
rect 5004 4136 5012 4144
rect 5052 4136 5060 4144
rect 5260 4136 5268 4144
rect 5692 4136 5700 4144
rect 1724 4116 1732 4124
rect 1788 4116 1796 4124
rect 1804 4116 1812 4124
rect 1868 4116 1876 4124
rect 1932 4116 1940 4124
rect 1948 4116 1956 4124
rect 1996 4116 2004 4124
rect 2012 4116 2020 4124
rect 2076 4116 2084 4124
rect 2284 4116 2292 4124
rect 2332 4118 2340 4126
rect 2396 4116 2404 4124
rect 2492 4116 2500 4124
rect 2556 4118 2564 4126
rect 2652 4116 2660 4124
rect 348 4096 356 4104
rect 380 4096 388 4104
rect 1388 4096 1396 4104
rect 1452 4096 1460 4104
rect 1644 4096 1652 4104
rect 1660 4096 1668 4104
rect 1756 4096 1764 4104
rect 1772 4096 1780 4104
rect 2732 4116 2740 4124
rect 2748 4116 2756 4124
rect 2908 4118 2916 4126
rect 3228 4116 3236 4124
rect 3292 4118 3300 4126
rect 3388 4116 3396 4124
rect 3452 4116 3460 4124
rect 3548 4116 3556 4124
rect 3852 4116 3860 4124
rect 3932 4116 3940 4124
rect 4316 4116 4324 4124
rect 4412 4116 4420 4124
rect 4556 4116 4564 4124
rect 4572 4116 4580 4124
rect 4924 4116 4932 4124
rect 5020 4116 5028 4124
rect 5084 4116 5092 4124
rect 5148 4116 5156 4124
rect 5372 4116 5380 4124
rect 5580 4116 5588 4124
rect 2764 4096 2772 4104
rect 3868 4096 3876 4104
rect 3900 4096 3908 4104
rect 4332 4096 4340 4104
rect 4364 4096 4372 4104
rect 4940 4096 4948 4104
rect 4972 4096 4980 4104
rect 5196 4100 5204 4108
rect 5788 4096 5796 4104
rect 220 4076 228 4084
rect 652 4076 660 4084
rect 1260 4076 1268 4084
rect 1532 4076 1540 4084
rect 4540 4076 4548 4084
rect 2780 4056 2788 4064
rect 76 4036 84 4044
rect 156 4036 164 4044
rect 1004 4036 1012 4044
rect 1036 4036 1044 4044
rect 1628 4036 1636 4044
rect 1884 4036 1892 4044
rect 2092 4036 2100 4044
rect 2188 4036 2196 4044
rect 2204 4036 2212 4044
rect 2428 4036 2436 4044
rect 3164 4036 3172 4044
rect 3564 4036 3572 4044
rect 4028 4036 4036 4044
rect 4636 4036 4644 4044
rect 5196 4036 5204 4044
rect 5452 4036 5460 4044
rect 5500 4036 5508 4044
rect 5788 4036 5796 4044
rect 1358 4006 1366 4014
rect 1372 4006 1380 4014
rect 1386 4006 1394 4014
rect 4446 4006 4454 4014
rect 4460 4006 4468 4014
rect 4474 4006 4482 4014
rect 2908 3996 2916 4004
rect 5084 3996 5092 4004
rect 2268 3976 2276 3984
rect 3004 3976 3012 3984
rect 3052 3976 3060 3984
rect 5068 3976 5076 3984
rect 5436 3976 5444 3984
rect 1788 3956 1796 3964
rect 2348 3956 2356 3964
rect 5116 3958 5124 3966
rect 5180 3958 5188 3966
rect 5532 3958 5540 3966
rect 1404 3936 1412 3944
rect 3276 3936 3284 3944
rect 108 3916 116 3924
rect 124 3916 132 3924
rect 220 3916 228 3924
rect 252 3916 260 3924
rect 380 3916 388 3924
rect 412 3916 420 3924
rect 444 3916 452 3924
rect 524 3916 532 3924
rect 28 3896 36 3904
rect 412 3896 420 3904
rect 540 3896 548 3904
rect 636 3896 644 3904
rect 860 3916 868 3924
rect 924 3916 932 3924
rect 972 3916 980 3924
rect 1084 3916 1092 3924
rect 1644 3916 1652 3924
rect 1660 3916 1668 3924
rect 1724 3916 1732 3924
rect 892 3896 900 3904
rect 1052 3896 1060 3904
rect 1196 3896 1204 3904
rect 1260 3894 1268 3902
rect 1612 3896 1620 3904
rect 1692 3896 1700 3904
rect 1724 3896 1732 3904
rect 1788 3896 1796 3904
rect 1836 3916 1844 3924
rect 1948 3916 1956 3924
rect 2028 3916 2036 3924
rect 2204 3916 2212 3924
rect 2252 3916 2260 3924
rect 2396 3916 2404 3924
rect 2668 3916 2676 3924
rect 2716 3916 2724 3924
rect 2812 3916 2820 3924
rect 3084 3916 3092 3924
rect 3132 3916 3140 3924
rect 3244 3916 3252 3924
rect 3260 3916 3268 3924
rect 4380 3916 4388 3924
rect 4748 3916 4756 3924
rect 4780 3916 4788 3924
rect 4892 3916 4900 3924
rect 5180 3912 5188 3920
rect 5532 3912 5540 3920
rect 1868 3896 1876 3904
rect 1996 3896 2004 3904
rect 2076 3896 2084 3904
rect 2092 3896 2100 3904
rect 2156 3896 2164 3904
rect 2332 3896 2340 3904
rect 2380 3896 2388 3904
rect 2492 3896 2500 3904
rect 2540 3896 2548 3904
rect 2748 3896 2756 3904
rect 3020 3896 3028 3904
rect 3116 3896 3124 3904
rect 3164 3896 3172 3904
rect 3212 3896 3220 3904
rect 3420 3894 3428 3902
rect 3484 3896 3492 3904
rect 3532 3896 3540 3904
rect 3692 3896 3700 3904
rect 3740 3896 3748 3904
rect 3772 3896 3780 3904
rect 3964 3896 3972 3904
rect 4028 3894 4036 3902
rect 4140 3896 4148 3904
rect 4188 3896 4196 3904
rect 4236 3896 4244 3904
rect 4284 3896 4292 3904
rect 4732 3896 4740 3904
rect 4812 3896 4820 3904
rect 4988 3896 4996 3904
rect 5052 3896 5060 3904
rect 5100 3896 5108 3904
rect 5148 3896 5156 3904
rect 5516 3896 5524 3904
rect 12 3876 20 3884
rect 76 3876 84 3884
rect 156 3876 164 3884
rect 204 3876 212 3884
rect 220 3876 228 3884
rect 332 3876 340 3884
rect 428 3876 436 3884
rect 476 3876 484 3884
rect 492 3876 500 3884
rect 540 3876 548 3884
rect 300 3856 308 3864
rect 364 3856 372 3864
rect 572 3856 580 3864
rect 620 3876 628 3884
rect 636 3876 644 3884
rect 748 3876 756 3884
rect 796 3876 804 3884
rect 828 3876 836 3884
rect 924 3876 932 3884
rect 1004 3876 1012 3884
rect 764 3856 772 3864
rect 1084 3876 1092 3884
rect 1292 3876 1300 3884
rect 1372 3876 1380 3884
rect 1468 3876 1476 3884
rect 1484 3876 1492 3884
rect 1580 3876 1588 3884
rect 1596 3876 1604 3884
rect 1628 3876 1636 3884
rect 1660 3876 1668 3884
rect 1708 3876 1716 3884
rect 1756 3876 1764 3884
rect 1772 3876 1780 3884
rect 1884 3876 1892 3884
rect 1900 3876 1908 3884
rect 1964 3876 1972 3884
rect 1980 3876 1988 3884
rect 2012 3876 2020 3884
rect 2124 3876 2132 3884
rect 2236 3876 2244 3884
rect 2284 3876 2292 3884
rect 2428 3876 2436 3884
rect 2476 3876 2484 3884
rect 1116 3856 1124 3864
rect 2044 3856 2052 3864
rect 2188 3856 2196 3864
rect 2300 3856 2308 3864
rect 2444 3856 2452 3864
rect 2556 3876 2564 3884
rect 2700 3876 2708 3884
rect 2748 3876 2756 3884
rect 2764 3876 2772 3884
rect 2828 3876 2836 3884
rect 2924 3876 2932 3884
rect 3036 3876 3044 3884
rect 3116 3876 3124 3884
rect 3180 3876 3188 3884
rect 3228 3876 3236 3884
rect 3388 3876 3396 3884
rect 3484 3876 3492 3884
rect 3580 3876 3588 3884
rect 3884 3876 3892 3884
rect 4220 3876 4228 3884
rect 4332 3876 4340 3884
rect 4636 3876 4644 3884
rect 4780 3876 4788 3884
rect 4812 3876 4820 3884
rect 4860 3876 4868 3884
rect 4924 3876 4932 3884
rect 5244 3876 5252 3884
rect 5596 3876 5604 3884
rect 2988 3856 2996 3864
rect 3276 3856 3284 3864
rect 3516 3856 3524 3864
rect 3612 3856 3620 3864
rect 3644 3856 3652 3864
rect 4028 3856 4036 3864
rect 4604 3856 4612 3864
rect 4876 3856 4884 3864
rect 4956 3856 4964 3864
rect 5276 3856 5284 3864
rect 5628 3856 5636 3864
rect 60 3836 68 3844
rect 236 3836 244 3844
rect 348 3836 356 3844
rect 444 3836 452 3844
rect 604 3836 612 3844
rect 700 3836 708 3844
rect 940 3836 948 3844
rect 1132 3836 1140 3844
rect 1516 3836 1524 3844
rect 1916 3836 1924 3844
rect 2460 3836 2468 3844
rect 2524 3836 2532 3844
rect 2588 3836 2596 3844
rect 2732 3836 2740 3844
rect 2812 3836 2820 3844
rect 2876 3836 2884 3844
rect 3100 3836 3108 3844
rect 3628 3836 3636 3844
rect 3900 3836 3908 3844
rect 4348 3836 4356 3844
rect 4444 3836 4452 3844
rect 4908 3836 4916 3844
rect 5020 3836 5028 3844
rect 5788 3836 5796 3844
rect 2910 3806 2918 3814
rect 2924 3806 2932 3814
rect 2938 3806 2946 3814
rect 332 3776 340 3784
rect 412 3776 420 3784
rect 1980 3776 1988 3784
rect 2332 3776 2340 3784
rect 2460 3776 2468 3784
rect 2620 3776 2628 3784
rect 2716 3776 2724 3784
rect 3116 3776 3124 3784
rect 3308 3776 3316 3784
rect 3692 3776 3700 3784
rect 3868 3776 3876 3784
rect 5308 3776 5316 3784
rect 5804 3776 5812 3784
rect 156 3756 164 3764
rect 188 3756 196 3764
rect 316 3756 324 3764
rect 1100 3756 1108 3764
rect 1292 3756 1300 3764
rect 1804 3756 1812 3764
rect 12 3736 20 3744
rect 108 3736 116 3744
rect 172 3736 180 3744
rect 252 3736 260 3744
rect 300 3736 308 3744
rect 364 3736 372 3744
rect 476 3736 484 3744
rect 652 3736 660 3744
rect 732 3736 740 3744
rect 764 3736 772 3744
rect 1500 3736 1508 3744
rect 1596 3736 1604 3744
rect 1916 3756 1924 3764
rect 2028 3756 2036 3764
rect 2428 3756 2436 3764
rect 2700 3756 2708 3764
rect 2780 3756 2788 3764
rect 2876 3756 2884 3764
rect 3020 3756 3028 3764
rect 1916 3736 1924 3744
rect 1948 3736 1956 3744
rect 92 3716 100 3724
rect 220 3716 228 3724
rect 252 3716 260 3724
rect 348 3716 356 3724
rect 380 3716 388 3724
rect 60 3696 68 3704
rect 204 3696 212 3704
rect 268 3696 276 3704
rect 284 3696 292 3704
rect 460 3716 468 3724
rect 620 3718 628 3726
rect 716 3716 724 3724
rect 844 3716 852 3724
rect 908 3718 916 3726
rect 1100 3718 1108 3726
rect 1276 3716 1284 3724
rect 1532 3718 1540 3726
rect 1724 3716 1732 3724
rect 1772 3716 1780 3724
rect 1788 3716 1796 3724
rect 1836 3716 1844 3724
rect 1852 3716 1860 3724
rect 1996 3736 2004 3744
rect 2124 3736 2132 3744
rect 2204 3736 2212 3744
rect 2236 3736 2244 3744
rect 2252 3736 2260 3744
rect 2284 3736 2292 3744
rect 2300 3736 2308 3744
rect 2396 3736 2404 3744
rect 2508 3736 2516 3744
rect 2572 3736 2580 3744
rect 2684 3736 2692 3744
rect 2732 3736 2740 3744
rect 2796 3736 2804 3744
rect 2828 3736 2836 3744
rect 2892 3736 2900 3744
rect 3020 3736 3028 3744
rect 3052 3736 3060 3744
rect 3500 3736 3508 3744
rect 3612 3736 3620 3744
rect 3724 3756 3732 3764
rect 3852 3756 3860 3764
rect 4284 3756 4292 3764
rect 4556 3756 4564 3764
rect 4748 3756 4756 3764
rect 4972 3756 4980 3764
rect 5148 3756 5156 3764
rect 5644 3756 5652 3764
rect 3820 3736 3828 3744
rect 4108 3736 4116 3744
rect 4316 3736 4324 3744
rect 4540 3736 4548 3744
rect 4780 3736 4788 3744
rect 4956 3736 4964 3744
rect 5116 3736 5124 3744
rect 5324 3736 5332 3744
rect 5468 3736 5476 3744
rect 5612 3736 5620 3744
rect 2076 3716 2084 3724
rect 2108 3716 2116 3724
rect 428 3696 436 3704
rect 684 3696 692 3704
rect 1628 3696 1636 3704
rect 1916 3696 1924 3704
rect 1996 3696 2004 3704
rect 2044 3696 2052 3704
rect 2124 3696 2132 3704
rect 2444 3716 2452 3724
rect 2492 3716 2500 3724
rect 2524 3716 2532 3724
rect 2556 3716 2564 3724
rect 2668 3716 2676 3724
rect 2748 3716 2756 3724
rect 2764 3716 2772 3724
rect 2172 3696 2180 3704
rect 2220 3696 2228 3704
rect 2252 3696 2260 3704
rect 2620 3696 2628 3704
rect 2636 3696 2644 3704
rect 2892 3716 2900 3724
rect 3196 3716 3204 3724
rect 3244 3718 3252 3726
rect 3388 3716 3396 3724
rect 3436 3718 3444 3726
rect 3516 3716 3524 3724
rect 3532 3716 3540 3724
rect 3628 3716 3636 3724
rect 3644 3716 3652 3724
rect 3676 3716 3684 3724
rect 3756 3716 3764 3724
rect 3804 3716 3812 3724
rect 3932 3716 3940 3724
rect 3996 3718 4004 3726
rect 4060 3716 4068 3724
rect 4412 3716 4420 3724
rect 4460 3716 4468 3724
rect 4876 3716 4884 3724
rect 4924 3716 4932 3724
rect 5020 3716 5028 3724
rect 5420 3716 5428 3724
rect 5516 3716 5524 3724
rect 2860 3696 2868 3704
rect 3100 3696 3108 3704
rect 3548 3696 3556 3704
rect 3660 3696 3668 3704
rect 3772 3696 3780 3704
rect 4380 3700 4388 3708
rect 4892 3696 4900 3704
rect 5020 3696 5028 3704
rect 5548 3700 5556 3708
rect 12 3676 20 3684
rect 140 3676 148 3684
rect 972 3676 980 3684
rect 1004 3676 1012 3684
rect 2076 3676 2084 3684
rect 2556 3676 2564 3684
rect 3804 3676 3812 3684
rect 1164 3656 1172 3664
rect 492 3636 500 3644
rect 748 3636 756 3644
rect 780 3636 788 3644
rect 1404 3636 1412 3644
rect 1900 3636 1908 3644
rect 2668 3636 2676 3644
rect 3068 3636 3076 3644
rect 3692 3636 3700 3644
rect 4124 3636 4132 3644
rect 4588 3636 4596 3644
rect 5020 3636 5028 3644
rect 5356 3636 5364 3644
rect 5452 3636 5460 3644
rect 5548 3636 5556 3644
rect 1358 3606 1366 3614
rect 1372 3606 1380 3614
rect 1386 3606 1394 3614
rect 4446 3606 4454 3614
rect 4460 3606 4468 3614
rect 4474 3606 4482 3614
rect 204 3576 212 3584
rect 348 3576 356 3584
rect 2508 3576 2516 3584
rect 2620 3576 2628 3584
rect 4812 3576 4820 3584
rect 5116 3576 5124 3584
rect 5532 3576 5540 3584
rect 2684 3556 2692 3564
rect 3260 3556 3268 3564
rect 5148 3558 5156 3566
rect 5212 3558 5220 3566
rect 3308 3536 3316 3544
rect 4844 3536 4852 3544
rect 12 3516 20 3524
rect 44 3516 52 3524
rect 284 3516 292 3524
rect 492 3516 500 3524
rect 604 3516 612 3524
rect 892 3516 900 3524
rect 1132 3516 1140 3524
rect 1356 3516 1364 3524
rect 1996 3516 2004 3524
rect 2332 3516 2340 3524
rect 2396 3516 2404 3524
rect 2476 3516 2484 3524
rect 2556 3516 2564 3524
rect 2780 3516 2788 3524
rect 44 3496 52 3504
rect 60 3496 68 3504
rect 60 3476 68 3484
rect 412 3496 420 3504
rect 476 3496 484 3504
rect 524 3496 532 3504
rect 572 3496 580 3504
rect 620 3496 628 3504
rect 652 3496 660 3504
rect 684 3496 692 3504
rect 764 3496 772 3504
rect 780 3496 788 3504
rect 876 3496 884 3504
rect 1004 3496 1012 3504
rect 1068 3494 1076 3502
rect 1596 3496 1604 3504
rect 1660 3494 1668 3502
rect 1788 3496 1796 3504
rect 1852 3494 1860 3502
rect 1916 3496 1924 3504
rect 1964 3496 1972 3504
rect 2092 3496 2100 3504
rect 2284 3496 2292 3504
rect 2364 3496 2372 3504
rect 2476 3496 2484 3504
rect 2764 3496 2772 3504
rect 2828 3516 2836 3524
rect 3036 3516 3044 3524
rect 3228 3516 3236 3524
rect 4124 3516 4132 3524
rect 4188 3516 4196 3524
rect 4316 3516 4324 3524
rect 4412 3516 4420 3524
rect 4508 3516 4516 3524
rect 4572 3516 4580 3524
rect 4684 3516 4692 3524
rect 5212 3512 5220 3520
rect 5532 3516 5540 3524
rect 2924 3496 2932 3504
rect 2988 3496 2996 3504
rect 3132 3496 3140 3504
rect 3148 3496 3156 3504
rect 3260 3496 3268 3504
rect 3388 3496 3396 3504
rect 3452 3494 3460 3502
rect 3516 3496 3524 3504
rect 3644 3496 3652 3504
rect 3740 3496 3748 3504
rect 4060 3494 4068 3502
rect 4124 3496 4132 3504
rect 4156 3496 4164 3504
rect 4172 3496 4180 3504
rect 4268 3496 4276 3504
rect 4300 3496 4308 3504
rect 4348 3496 4356 3504
rect 4524 3496 4532 3504
rect 4636 3496 4644 3504
rect 4940 3494 4948 3502
rect 5180 3496 5188 3504
rect 5516 3496 5524 3504
rect 5532 3496 5540 3504
rect 172 3476 180 3484
rect 220 3476 228 3484
rect 332 3476 340 3484
rect 380 3476 388 3484
rect 460 3476 468 3484
rect 508 3476 516 3484
rect 540 3476 548 3484
rect 556 3476 564 3484
rect 620 3476 628 3484
rect 636 3476 644 3484
rect 764 3476 772 3484
rect 188 3456 196 3464
rect 332 3456 340 3464
rect 364 3456 372 3464
rect 428 3456 436 3464
rect 732 3456 740 3464
rect 1164 3476 1172 3484
rect 1196 3476 1204 3484
rect 1212 3476 1220 3484
rect 1308 3476 1316 3484
rect 1324 3476 1332 3484
rect 1420 3476 1428 3484
rect 1516 3476 1524 3484
rect 1964 3476 1972 3484
rect 2060 3476 2068 3484
rect 2076 3476 2084 3484
rect 2140 3476 2148 3484
rect 2188 3476 2196 3484
rect 2220 3476 2228 3484
rect 2316 3476 2324 3484
rect 2380 3476 2388 3484
rect 2428 3476 2436 3484
rect 2444 3476 2452 3484
rect 2492 3476 2500 3484
rect 2540 3476 2548 3484
rect 2636 3476 2644 3484
rect 2652 3476 2660 3484
rect 2748 3476 2756 3484
rect 2764 3476 2772 3484
rect 2860 3476 2868 3484
rect 2940 3476 2948 3484
rect 3276 3476 3284 3484
rect 3484 3476 3492 3484
rect 3708 3476 3716 3484
rect 3788 3476 3796 3484
rect 3916 3476 3924 3484
rect 4028 3476 4036 3484
rect 4172 3476 4180 3484
rect 4236 3476 4244 3484
rect 4252 3476 4260 3484
rect 4380 3476 4388 3484
rect 4540 3476 4548 3484
rect 4636 3476 4644 3484
rect 4684 3476 4692 3484
rect 4876 3476 4884 3484
rect 4972 3476 4980 3484
rect 5004 3476 5012 3484
rect 5276 3476 5284 3484
rect 5470 3476 5478 3484
rect 5628 3476 5636 3484
rect 844 3456 852 3464
rect 1948 3456 1956 3464
rect 2092 3456 2100 3464
rect 2156 3456 2164 3464
rect 2956 3456 2964 3464
rect 3020 3456 3028 3464
rect 3084 3456 3092 3464
rect 3100 3456 3108 3464
rect 3132 3456 3140 3464
rect 3212 3456 3220 3464
rect 3308 3456 3316 3464
rect 3452 3456 3460 3464
rect 3532 3456 3540 3464
rect 3676 3456 3684 3464
rect 4396 3456 4404 3464
rect 4428 3456 4436 3464
rect 4492 3456 4500 3464
rect 4588 3456 4596 3464
rect 5308 3456 5316 3464
rect 5660 3456 5668 3464
rect 124 3436 132 3444
rect 204 3436 212 3444
rect 252 3436 260 3444
rect 348 3436 356 3444
rect 444 3436 452 3444
rect 748 3436 756 3444
rect 812 3436 820 3444
rect 892 3436 900 3444
rect 940 3436 948 3444
rect 1132 3436 1140 3444
rect 1180 3436 1188 3444
rect 1276 3436 1284 3444
rect 1404 3436 1412 3444
rect 1484 3436 1492 3444
rect 1532 3436 1540 3444
rect 1724 3436 1732 3444
rect 2252 3436 2260 3444
rect 2412 3436 2420 3444
rect 2476 3436 2484 3444
rect 2620 3436 2628 3444
rect 3116 3436 3124 3444
rect 3196 3436 3204 3444
rect 3548 3436 3556 3444
rect 3836 3436 3844 3444
rect 3900 3436 3908 3444
rect 3932 3436 3940 3444
rect 4300 3436 4308 3444
rect 4556 3436 4564 3444
rect 4604 3436 4612 3444
rect 4684 3436 4692 3444
rect 4732 3436 4740 3444
rect 5116 3436 5124 3444
rect 5820 3436 5828 3444
rect 2910 3406 2918 3414
rect 2924 3406 2932 3414
rect 2938 3406 2946 3414
rect 220 3376 228 3384
rect 828 3376 836 3384
rect 1132 3376 1140 3384
rect 2332 3376 2340 3384
rect 2668 3376 2676 3384
rect 3340 3376 3348 3384
rect 3564 3376 3572 3384
rect 4748 3376 4756 3384
rect 4940 3376 4948 3384
rect 5132 3376 5140 3384
rect 5212 3376 5220 3384
rect 268 3356 276 3364
rect 588 3356 596 3364
rect 604 3356 612 3364
rect 1036 3356 1044 3364
rect 1164 3356 1172 3364
rect 1596 3356 1604 3364
rect 1628 3356 1636 3364
rect 1644 3356 1652 3364
rect 2684 3356 2692 3364
rect 2700 3356 2708 3364
rect 2732 3356 2740 3364
rect 2812 3356 2820 3364
rect 2988 3356 2996 3364
rect 3116 3356 3124 3364
rect 3180 3356 3188 3364
rect 3548 3356 3556 3364
rect 4636 3356 4644 3364
rect 5372 3356 5380 3364
rect 12 3336 20 3344
rect 108 3336 116 3344
rect 188 3336 196 3344
rect 380 3336 388 3344
rect 412 3336 420 3344
rect 492 3336 500 3344
rect 796 3336 804 3344
rect 812 3336 820 3344
rect 892 3336 900 3344
rect 956 3336 964 3344
rect 1020 3336 1028 3344
rect 1068 3336 1076 3344
rect 1084 3336 1092 3344
rect 1180 3336 1188 3344
rect 1260 3336 1268 3344
rect 1340 3336 1348 3344
rect 1372 3336 1380 3344
rect 1436 3336 1444 3344
rect 1548 3336 1556 3344
rect 1564 3336 1572 3344
rect 1596 3336 1604 3344
rect 1724 3336 1732 3344
rect 1740 3336 1748 3344
rect 1836 3336 1844 3344
rect 1980 3336 1988 3344
rect 2108 3336 2116 3344
rect 2188 3336 2196 3344
rect 2284 3336 2292 3344
rect 2300 3336 2308 3344
rect 2396 3336 2404 3344
rect 2460 3336 2468 3344
rect 2508 3336 2516 3344
rect 2620 3336 2628 3344
rect 2652 3336 2660 3344
rect 2748 3336 2756 3344
rect 3004 3336 3012 3344
rect 3068 3336 3076 3344
rect 3148 3336 3156 3344
rect 3228 3336 3236 3344
rect 3324 3336 3332 3344
rect 3452 3336 3460 3344
rect 3676 3336 3684 3344
rect 3756 3336 3764 3344
rect 3820 3336 3828 3344
rect 3884 3336 3892 3344
rect 3900 3336 3908 3344
rect 4108 3336 4116 3344
rect 4236 3336 4244 3344
rect 4332 3336 4340 3344
rect 4476 3336 4484 3344
rect 4540 3336 4548 3344
rect 4700 3336 4708 3344
rect 4972 3336 4980 3344
rect 5404 3336 5412 3344
rect 5852 3336 5860 3344
rect 140 3316 148 3324
rect 252 3316 260 3324
rect 300 3316 308 3324
rect 364 3316 372 3324
rect 444 3316 452 3324
rect 476 3316 484 3324
rect 540 3316 548 3324
rect 716 3316 724 3324
rect 780 3316 788 3324
rect 444 3296 452 3304
rect 668 3296 676 3304
rect 732 3296 740 3304
rect 748 3296 756 3304
rect 908 3316 916 3324
rect 956 3316 964 3324
rect 1020 3316 1028 3324
rect 1100 3316 1108 3324
rect 1132 3316 1140 3324
rect 1196 3316 1204 3324
rect 1228 3316 1236 3324
rect 860 3296 868 3304
rect 892 3296 900 3304
rect 972 3296 980 3304
rect 1132 3296 1140 3304
rect 1196 3296 1204 3304
rect 1308 3296 1316 3304
rect 1388 3316 1396 3324
rect 1548 3316 1556 3324
rect 1580 3316 1588 3324
rect 1676 3316 1684 3324
rect 2124 3318 2132 3326
rect 2188 3316 2196 3324
rect 2348 3316 2356 3324
rect 2444 3316 2452 3324
rect 2540 3316 2548 3324
rect 2636 3316 2644 3324
rect 2732 3316 2740 3324
rect 2844 3316 2852 3324
rect 2956 3316 2964 3324
rect 3020 3316 3028 3324
rect 3212 3316 3220 3324
rect 3404 3316 3412 3324
rect 3468 3318 3476 3326
rect 3532 3316 3540 3324
rect 3692 3318 3700 3326
rect 3772 3316 3780 3324
rect 3804 3316 3812 3324
rect 3852 3316 3860 3324
rect 3868 3316 3876 3324
rect 4028 3316 4036 3324
rect 4076 3318 4084 3326
rect 4268 3318 4276 3326
rect 4492 3316 4500 3324
rect 4556 3316 4564 3324
rect 4604 3316 4612 3324
rect 2412 3296 2420 3304
rect 2476 3296 2484 3304
rect 2508 3296 2516 3304
rect 2796 3296 2804 3304
rect 3100 3296 3108 3304
rect 3836 3296 3844 3304
rect 3932 3296 3940 3304
rect 4588 3296 4596 3304
rect 4684 3316 4692 3324
rect 4860 3316 4868 3324
rect 4876 3316 4884 3324
rect 5004 3318 5012 3326
rect 5068 3316 5076 3324
rect 5148 3316 5156 3324
rect 5468 3316 5476 3324
rect 5612 3316 5620 3324
rect 5660 3316 5668 3324
rect 5740 3316 5748 3324
rect 5788 3316 5796 3324
rect 4684 3296 4692 3304
rect 4748 3296 4756 3304
rect 5500 3296 5508 3304
rect 476 3276 484 3284
rect 524 3276 532 3284
rect 652 3276 660 3284
rect 700 3276 708 3284
rect 2540 3276 2548 3284
rect 2556 3276 2564 3284
rect 3020 3276 3028 3284
rect 4364 3276 4372 3284
rect 5772 3276 5780 3284
rect 716 3256 724 3264
rect 2764 3256 2772 3264
rect 60 3236 68 3244
rect 220 3236 228 3244
rect 284 3236 292 3244
rect 332 3236 340 3244
rect 412 3236 420 3244
rect 540 3236 548 3244
rect 780 3236 788 3244
rect 1004 3236 1012 3244
rect 1468 3236 1476 3244
rect 1868 3236 1876 3244
rect 1996 3236 2004 3244
rect 2444 3236 2452 3244
rect 2604 3236 2612 3244
rect 2892 3236 2900 3244
rect 3260 3236 3268 3244
rect 3772 3236 3780 3244
rect 3948 3236 3956 3244
rect 4140 3236 4148 3244
rect 4556 3236 4564 3244
rect 5500 3236 5508 3244
rect 5548 3236 5556 3244
rect 1358 3206 1366 3214
rect 1372 3206 1380 3214
rect 1386 3206 1394 3214
rect 4446 3206 4454 3214
rect 4460 3206 4468 3214
rect 4474 3206 4482 3214
rect 748 3176 756 3184
rect 2732 3176 2740 3184
rect 3516 3176 3524 3184
rect 3788 3176 3796 3184
rect 4684 3176 4692 3184
rect 4764 3176 4772 3184
rect 4972 3176 4980 3184
rect 1196 3136 1204 3144
rect 1996 3136 2004 3144
rect 4044 3136 4052 3144
rect 5628 3136 5636 3144
rect 12 3116 20 3124
rect 252 3116 260 3124
rect 316 3116 324 3124
rect 444 3116 452 3124
rect 44 3096 52 3104
rect 108 3096 116 3104
rect 156 3096 164 3104
rect 204 3096 212 3104
rect 284 3096 292 3104
rect 364 3096 372 3104
rect 492 3116 500 3124
rect 636 3116 644 3124
rect 988 3116 996 3124
rect 1100 3116 1108 3124
rect 1228 3116 1236 3124
rect 1276 3116 1284 3124
rect 1372 3116 1380 3124
rect 1500 3116 1508 3124
rect 492 3096 500 3104
rect 508 3096 516 3104
rect 76 3076 84 3084
rect 172 3076 180 3084
rect 268 3076 276 3084
rect 300 3076 308 3084
rect 348 3076 356 3084
rect 412 3076 420 3084
rect 508 3076 516 3084
rect 716 3096 724 3104
rect 764 3096 772 3104
rect 844 3096 852 3104
rect 956 3096 964 3104
rect 1068 3096 1076 3104
rect 1116 3096 1124 3104
rect 1324 3096 1332 3104
rect 1436 3096 1444 3104
rect 2284 3116 2292 3124
rect 2316 3116 2324 3124
rect 2348 3116 2356 3124
rect 2556 3116 2564 3124
rect 3228 3116 3236 3124
rect 3276 3116 3284 3124
rect 3324 3116 3332 3124
rect 3388 3116 3396 3124
rect 3452 3116 3460 3124
rect 4444 3116 4452 3124
rect 4540 3116 4548 3124
rect 1564 3096 1572 3104
rect 1580 3096 1588 3104
rect 1692 3096 1700 3104
rect 1756 3096 1764 3104
rect 1868 3096 1876 3104
rect 1932 3094 1940 3102
rect 2124 3094 2132 3102
rect 2220 3096 2228 3104
rect 2284 3096 2292 3104
rect 2316 3096 2324 3104
rect 2396 3096 2404 3104
rect 2428 3096 2436 3104
rect 2524 3096 2532 3104
rect 2636 3096 2644 3104
rect 2668 3096 2676 3104
rect 2716 3096 2724 3104
rect 620 3076 628 3084
rect 684 3076 692 3084
rect 700 3076 708 3084
rect 796 3076 804 3084
rect 828 3076 836 3084
rect 860 3076 868 3084
rect 924 3076 932 3084
rect 1052 3076 1060 3084
rect 1084 3076 1092 3084
rect 1132 3076 1140 3084
rect 1180 3076 1188 3084
rect 1308 3076 1316 3084
rect 1420 3076 1428 3084
rect 1452 3076 1460 3084
rect 1468 3076 1476 3084
rect 1516 3076 1524 3084
rect 1580 3076 1588 3084
rect 1612 3076 1620 3084
rect 2108 3076 2116 3084
rect 2396 3076 2404 3084
rect 2444 3076 2452 3084
rect 2508 3076 2516 3084
rect 2572 3076 2580 3084
rect 2860 3094 2868 3102
rect 3036 3096 3044 3104
rect 3100 3094 3108 3102
rect 3164 3096 3172 3104
rect 3308 3096 3316 3104
rect 3356 3096 3364 3104
rect 3420 3096 3428 3104
rect 3436 3096 3444 3104
rect 3484 3096 3492 3104
rect 3532 3096 3540 3104
rect 3756 3096 3764 3104
rect 3804 3096 3812 3104
rect 3852 3096 3860 3104
rect 3884 3096 3892 3104
rect 3916 3096 3924 3104
rect 3964 3096 3972 3104
rect 4108 3096 4116 3104
rect 4172 3094 4180 3102
rect 4236 3096 4244 3104
rect 4300 3096 4308 3104
rect 4348 3096 4356 3104
rect 4380 3096 4388 3104
rect 4396 3096 4404 3104
rect 5292 3116 5300 3124
rect 5340 3116 5348 3124
rect 5356 3116 5364 3124
rect 4572 3096 4580 3104
rect 4588 3096 4596 3104
rect 4844 3094 4852 3102
rect 5292 3096 5300 3104
rect 5372 3096 5380 3104
rect 5500 3094 5508 3102
rect 5692 3094 5700 3102
rect 2828 3076 2836 3084
rect 2924 3076 2932 3084
rect 3212 3076 3220 3084
rect 3308 3076 3316 3084
rect 3372 3076 3380 3084
rect 3436 3076 3444 3084
rect 204 3056 212 3064
rect 236 3056 244 3064
rect 396 3056 404 3064
rect 684 3056 692 3064
rect 876 3056 884 3064
rect 924 3056 932 3064
rect 1004 3056 1012 3064
rect 1164 3056 1172 3064
rect 1244 3056 1252 3064
rect 1340 3056 1348 3064
rect 1612 3056 1620 3064
rect 1692 3056 1700 3064
rect 1724 3056 1732 3064
rect 2204 3054 2212 3062
rect 2412 3056 2420 3064
rect 2492 3056 2500 3064
rect 3548 3076 3556 3084
rect 3644 3076 3652 3084
rect 3660 3076 3668 3084
rect 3756 3076 3764 3084
rect 3772 3076 3780 3084
rect 3868 3076 3876 3084
rect 4012 3076 4020 3084
rect 4252 3076 4260 3084
rect 4284 3076 4292 3084
rect 3820 3056 3828 3064
rect 3884 3056 3892 3064
rect 3964 3056 3972 3064
rect 4028 3056 4036 3064
rect 4412 3076 4420 3084
rect 4508 3076 4516 3084
rect 4604 3076 4612 3084
rect 4636 3076 4644 3084
rect 4748 3076 4756 3084
rect 4876 3076 4884 3084
rect 5196 3076 5204 3084
rect 5372 3076 5380 3084
rect 5420 3076 5428 3084
rect 5516 3076 5524 3084
rect 5660 3076 5668 3084
rect 4780 3056 4788 3064
rect 5004 3056 5012 3064
rect 5164 3056 5172 3064
rect 5436 3056 5444 3064
rect 12 3036 20 3044
rect 140 3036 148 3044
rect 332 3036 340 3044
rect 380 3036 388 3044
rect 556 3036 564 3044
rect 652 3036 660 3044
rect 812 3036 820 3044
rect 988 3036 996 3044
rect 1020 3036 1028 3044
rect 1148 3036 1156 3044
rect 1260 3036 1268 3044
rect 1292 3036 1300 3044
rect 1500 3036 1508 3044
rect 1596 3036 1604 3044
rect 1708 3036 1716 3044
rect 1788 3036 1796 3044
rect 1804 3036 1812 3044
rect 2972 3036 2980 3044
rect 3228 3036 3236 3044
rect 3692 3036 3700 3044
rect 3948 3036 3956 3044
rect 4252 3036 4260 3044
rect 4332 3036 4340 3044
rect 4492 3036 4500 3044
rect 4620 3036 4628 3044
rect 5820 3036 5828 3044
rect 2316 3016 2324 3024
rect 2910 3006 2918 3014
rect 2924 3006 2932 3014
rect 2938 3006 2946 3014
rect 460 2976 468 2984
rect 764 2976 772 2984
rect 908 2976 916 2984
rect 1036 2976 1044 2984
rect 1500 2976 1508 2984
rect 1564 2976 1572 2984
rect 2444 2976 2452 2984
rect 3676 2976 3684 2984
rect 4140 2976 4148 2984
rect 4876 2976 4884 2984
rect 12 2956 20 2964
rect 60 2956 68 2964
rect 284 2956 292 2964
rect 364 2956 372 2964
rect 780 2956 788 2964
rect 1132 2956 1140 2964
rect 1308 2956 1316 2964
rect 1516 2956 1524 2964
rect 1580 2956 1588 2964
rect 1676 2956 1684 2964
rect 1788 2956 1796 2964
rect 2108 2956 2116 2964
rect 2236 2958 2244 2966
rect 3276 2956 3284 2964
rect 4044 2956 4052 2964
rect 4492 2956 4500 2964
rect 5516 2956 5524 2964
rect 5788 2956 5796 2964
rect 124 2936 132 2944
rect 204 2936 212 2944
rect 348 2936 356 2944
rect 396 2936 404 2944
rect 444 2936 452 2944
rect 476 2936 484 2944
rect 508 2936 516 2944
rect 620 2936 628 2944
rect 636 2936 644 2944
rect 732 2936 740 2944
rect 796 2936 804 2944
rect 844 2936 852 2944
rect 876 2936 884 2944
rect 924 2936 932 2944
rect 1020 2936 1028 2944
rect 1052 2936 1060 2944
rect 1068 2936 1076 2944
rect 1196 2936 1204 2944
rect 1228 2936 1236 2944
rect 1276 2936 1284 2944
rect 1292 2936 1300 2944
rect 1468 2936 1476 2944
rect 1532 2936 1540 2944
rect 1596 2936 1604 2944
rect 1756 2936 1764 2944
rect 1836 2936 1844 2944
rect 124 2916 132 2924
rect 172 2916 180 2924
rect 220 2916 228 2924
rect 236 2916 244 2924
rect 284 2916 292 2924
rect 332 2916 340 2924
rect 412 2916 420 2924
rect 492 2916 500 2924
rect 524 2916 532 2924
rect 28 2896 36 2904
rect 76 2896 84 2904
rect 188 2896 196 2904
rect 300 2896 308 2904
rect 556 2896 564 2904
rect 652 2916 660 2924
rect 748 2916 756 2924
rect 860 2916 868 2924
rect 908 2916 916 2924
rect 1068 2916 1076 2924
rect 1084 2916 1092 2924
rect 1212 2916 1220 2924
rect 1260 2916 1268 2924
rect 1372 2916 1380 2924
rect 1484 2916 1492 2924
rect 1532 2916 1540 2924
rect 1612 2916 1620 2924
rect 1740 2916 1748 2924
rect 1756 2916 1764 2924
rect 1820 2916 1828 2924
rect 1852 2916 1860 2924
rect 2316 2936 2324 2944
rect 2460 2936 2468 2944
rect 2556 2936 2564 2944
rect 3004 2936 3012 2944
rect 3052 2936 3060 2944
rect 3212 2936 3220 2944
rect 3404 2936 3412 2944
rect 3868 2936 3876 2944
rect 4028 2936 4036 2944
rect 4124 2936 4132 2944
rect 4332 2936 4340 2944
rect 4428 2936 4436 2944
rect 4524 2936 4532 2944
rect 4572 2936 4580 2944
rect 4588 2936 4596 2944
rect 4668 2936 4676 2944
rect 4844 2936 4852 2944
rect 4940 2936 4948 2944
rect 4956 2936 4964 2944
rect 5084 2936 5092 2944
rect 5116 2936 5124 2944
rect 5164 2936 5172 2944
rect 5548 2936 5556 2944
rect 5692 2936 5700 2944
rect 5788 2936 5796 2944
rect 2044 2916 2052 2924
rect 2108 2918 2116 2926
rect 2204 2916 2212 2924
rect 2220 2916 2228 2924
rect 2332 2916 2340 2924
rect 2460 2916 2468 2924
rect 2636 2916 2644 2924
rect 2700 2918 2708 2926
rect 2828 2916 2836 2924
rect 2892 2918 2900 2926
rect 3036 2916 3044 2924
rect 3420 2918 3428 2926
rect 3548 2916 3556 2924
rect 3612 2918 3620 2926
rect 3740 2916 3748 2924
rect 3804 2918 3812 2926
rect 4012 2916 4020 2924
rect 4076 2916 4084 2924
rect 4108 2916 4116 2924
rect 4204 2916 4212 2924
rect 4252 2916 4260 2924
rect 4604 2916 4612 2924
rect 4700 2918 4708 2926
rect 5148 2918 5156 2926
rect 5644 2916 5652 2924
rect 5740 2916 5748 2924
rect 5804 2916 5812 2924
rect 700 2896 708 2904
rect 908 2896 916 2904
rect 1132 2896 1140 2904
rect 1228 2896 1236 2904
rect 1324 2896 1332 2904
rect 1436 2896 1444 2904
rect 1612 2896 1620 2904
rect 1852 2896 1860 2904
rect 3020 2896 3028 2904
rect 3036 2896 3044 2904
rect 3164 2896 3172 2904
rect 3980 2896 3988 2904
rect 4572 2896 4580 2904
rect 4636 2896 4644 2904
rect 5644 2896 5652 2904
rect 5692 2896 5700 2904
rect 5724 2896 5732 2904
rect 156 2876 164 2884
rect 1900 2876 1908 2884
rect 3900 2876 3908 2884
rect 4604 2876 4612 2884
rect 4828 2876 4836 2884
rect 5244 2876 5252 2884
rect 5276 2876 5284 2884
rect 5852 2876 5860 2884
rect 604 2856 612 2864
rect 1084 2856 1092 2864
rect 1980 2856 1988 2864
rect 4364 2856 4372 2864
rect 44 2836 52 2844
rect 108 2836 116 2844
rect 172 2836 180 2844
rect 364 2836 372 2844
rect 652 2836 660 2844
rect 812 2836 820 2844
rect 1164 2836 1172 2844
rect 1356 2836 1364 2844
rect 1692 2836 1700 2844
rect 1756 2836 1764 2844
rect 2572 2836 2580 2844
rect 2764 2836 2772 2844
rect 3292 2836 3300 2844
rect 3484 2836 3492 2844
rect 5292 2836 5300 2844
rect 1358 2806 1366 2814
rect 1372 2806 1380 2814
rect 1386 2806 1394 2814
rect 4446 2806 4454 2814
rect 4460 2806 4468 2814
rect 4474 2806 4482 2814
rect 300 2776 308 2784
rect 572 2776 580 2784
rect 1260 2776 1268 2784
rect 3868 2776 3876 2784
rect 4092 2776 4100 2784
rect 4108 2776 4116 2784
rect 4556 2776 4564 2784
rect 4620 2776 4628 2784
rect 188 2736 196 2744
rect 1788 2736 1796 2744
rect 2204 2736 2212 2744
rect 2620 2736 2628 2744
rect 3644 2736 3652 2744
rect 3852 2736 3860 2744
rect 4124 2736 4132 2744
rect 4828 2736 4836 2744
rect 5212 2736 5220 2744
rect 5596 2736 5604 2744
rect 5788 2736 5796 2744
rect 220 2716 228 2724
rect 316 2716 324 2724
rect 796 2716 804 2724
rect 1180 2716 1188 2724
rect 1276 2716 1284 2724
rect 1372 2716 1380 2724
rect 1484 2716 1492 2724
rect 1500 2716 1508 2724
rect 1532 2716 1540 2724
rect 1724 2716 1732 2724
rect 60 2696 68 2704
rect 268 2696 276 2704
rect 348 2696 356 2704
rect 428 2696 436 2704
rect 476 2696 484 2704
rect 556 2696 564 2704
rect 684 2696 692 2704
rect 716 2696 724 2704
rect 764 2696 772 2704
rect 828 2696 836 2704
rect 972 2696 980 2704
rect 1100 2696 1108 2704
rect 1116 2696 1124 2704
rect 1212 2696 1220 2704
rect 1228 2696 1236 2704
rect 1308 2696 1316 2704
rect 1452 2696 1460 2704
rect 1468 2696 1476 2704
rect 1580 2696 1588 2704
rect 1612 2696 1620 2704
rect 1628 2696 1636 2704
rect 1692 2696 1700 2704
rect 2396 2716 2404 2724
rect 1868 2696 1876 2704
rect 1916 2694 1924 2702
rect 2060 2696 2068 2704
rect 2108 2694 2116 2702
rect 2284 2696 2292 2704
rect 2332 2696 2340 2704
rect 2380 2696 2388 2704
rect 2412 2696 2420 2704
rect 2428 2696 2436 2704
rect 2588 2716 2596 2724
rect 2684 2716 2692 2724
rect 3132 2716 3140 2724
rect 3308 2716 3316 2724
rect 3724 2716 3732 2724
rect 3820 2716 3828 2724
rect 3948 2716 3956 2724
rect 3980 2716 3988 2724
rect 4044 2716 4052 2724
rect 4380 2716 4388 2724
rect 4636 2716 4644 2724
rect 44 2676 52 2684
rect 76 2676 84 2684
rect 172 2676 180 2684
rect 364 2676 372 2684
rect 412 2676 420 2684
rect 460 2676 468 2684
rect 524 2676 532 2684
rect 588 2676 596 2684
rect 684 2676 692 2684
rect 844 2676 852 2684
rect 860 2676 868 2684
rect 956 2676 964 2684
rect 988 2676 996 2684
rect 1020 2676 1028 2684
rect 1164 2676 1172 2684
rect 1244 2676 1252 2684
rect 1324 2676 1332 2684
rect 1340 2676 1348 2684
rect 1548 2676 1556 2684
rect 1596 2676 1604 2684
rect 1660 2676 1668 2684
rect 1676 2676 1684 2684
rect 1772 2676 1780 2684
rect 1852 2676 1860 2684
rect 2172 2676 2180 2684
rect 2492 2696 2500 2704
rect 2508 2696 2516 2704
rect 2652 2696 2660 2704
rect 3004 2696 3012 2704
rect 3036 2696 3044 2704
rect 3084 2696 3092 2704
rect 3116 2696 3124 2704
rect 3164 2696 3172 2704
rect 3212 2696 3220 2704
rect 3244 2696 3252 2704
rect 3340 2696 3348 2704
rect 3548 2694 3556 2702
rect 3708 2696 3716 2704
rect 3836 2696 3844 2704
rect 3884 2696 3892 2704
rect 4060 2696 4068 2704
rect 4204 2696 4212 2704
rect 4268 2694 4276 2702
rect 4332 2696 4340 2704
rect 4396 2696 4404 2704
rect 4444 2696 4452 2704
rect 4700 2694 4708 2702
rect 4892 2694 4900 2702
rect 4956 2696 4964 2704
rect 5100 2696 5108 2704
rect 5276 2694 5284 2702
rect 5468 2694 5476 2702
rect 5516 2696 5524 2704
rect 5660 2694 5668 2702
rect 5804 2696 5812 2704
rect 2300 2676 2308 2684
rect 12 2656 20 2664
rect 188 2656 196 2664
rect 284 2656 292 2664
rect 380 2656 388 2664
rect 460 2656 468 2664
rect 556 2656 564 2664
rect 1004 2656 1012 2664
rect 1020 2656 1028 2664
rect 1052 2656 1060 2664
rect 1068 2656 1076 2664
rect 1580 2656 1588 2664
rect 2444 2676 2452 2684
rect 2460 2676 2468 2684
rect 2508 2676 2516 2684
rect 2556 2680 2564 2688
rect 2572 2676 2580 2684
rect 2620 2676 2628 2684
rect 2796 2676 2804 2684
rect 2812 2676 2820 2684
rect 2844 2676 2852 2684
rect 2940 2676 2948 2684
rect 2956 2676 2964 2684
rect 2348 2656 2356 2664
rect 2828 2656 2836 2664
rect 3052 2676 3060 2684
rect 3084 2676 3092 2684
rect 3180 2676 3188 2684
rect 3196 2676 3204 2684
rect 3260 2676 3268 2684
rect 3340 2676 3348 2684
rect 3388 2676 3396 2684
rect 3516 2676 3524 2684
rect 3580 2676 3588 2684
rect 3612 2676 3620 2684
rect 3708 2676 3716 2684
rect 3772 2676 3780 2684
rect 3900 2676 3908 2684
rect 4028 2676 4036 2684
rect 4300 2676 4308 2684
rect 4428 2676 4436 2684
rect 4492 2676 4500 2684
rect 4588 2676 4596 2684
rect 4604 2676 4612 2684
rect 4668 2676 4676 2684
rect 4924 2676 4932 2684
rect 5116 2676 5124 2684
rect 5244 2676 5252 2684
rect 5340 2676 5348 2684
rect 5436 2676 5444 2684
rect 5628 2676 5636 2684
rect 5852 2676 5860 2684
rect 3052 2656 3060 2664
rect 3116 2656 3124 2664
rect 3212 2656 3220 2664
rect 3292 2656 3300 2664
rect 3404 2656 3412 2664
rect 3804 2656 3812 2664
rect 3932 2656 3940 2664
rect 3964 2656 3972 2664
rect 4028 2656 4036 2664
rect 4060 2656 4068 2664
rect 4124 2656 4132 2664
rect 4364 2656 4372 2664
rect 28 2636 36 2644
rect 124 2636 132 2644
rect 220 2636 228 2644
rect 316 2636 324 2644
rect 396 2636 404 2644
rect 508 2636 516 2644
rect 620 2636 628 2644
rect 732 2636 740 2644
rect 796 2636 804 2644
rect 924 2636 932 2644
rect 1180 2636 1188 2644
rect 1276 2636 1284 2644
rect 1740 2636 1748 2644
rect 1980 2636 1988 2644
rect 2732 2636 2740 2644
rect 2876 2636 2884 2644
rect 3324 2636 3332 2644
rect 3420 2636 3428 2644
rect 3916 2636 3924 2644
rect 3980 2636 3988 2644
rect 4092 2636 4100 2644
rect 4108 2636 4116 2644
rect 4348 2636 4356 2644
rect 5020 2636 5028 2644
rect 5404 2636 5412 2644
rect 2910 2606 2918 2614
rect 2924 2606 2932 2614
rect 2938 2606 2946 2614
rect 412 2576 420 2584
rect 476 2576 484 2584
rect 764 2576 772 2584
rect 1580 2576 1588 2584
rect 1708 2576 1716 2584
rect 1996 2576 2004 2584
rect 2188 2576 2196 2584
rect 2620 2576 2628 2584
rect 2892 2576 2900 2584
rect 3292 2576 3300 2584
rect 3452 2576 3460 2584
rect 3676 2576 3684 2584
rect 3964 2576 3972 2584
rect 3996 2576 4004 2584
rect 4188 2576 4196 2584
rect 4412 2576 4420 2584
rect 4572 2576 4580 2584
rect 4636 2576 4644 2584
rect 4908 2576 4916 2584
rect 5100 2576 5108 2584
rect 5212 2576 5220 2584
rect 5324 2576 5332 2584
rect 156 2556 164 2564
rect 236 2556 244 2564
rect 492 2556 500 2564
rect 780 2556 788 2564
rect 12 2536 20 2544
rect 108 2536 116 2544
rect 124 2536 132 2544
rect 204 2536 212 2544
rect 220 2536 228 2544
rect 396 2536 404 2544
rect 460 2536 468 2544
rect 604 2536 612 2544
rect 620 2536 628 2544
rect 748 2536 756 2544
rect 780 2536 788 2544
rect 908 2556 916 2564
rect 940 2556 948 2564
rect 1100 2556 1108 2564
rect 1148 2556 1156 2564
rect 1228 2556 1236 2564
rect 1260 2556 1268 2564
rect 1804 2556 1812 2564
rect 1900 2556 1908 2564
rect 1932 2556 1940 2564
rect 1980 2556 1988 2564
rect 2316 2556 2324 2564
rect 3404 2556 3412 2564
rect 3500 2556 3508 2564
rect 3532 2556 3540 2564
rect 3564 2556 3572 2564
rect 3660 2556 3668 2564
rect 3948 2556 3956 2564
rect 4428 2556 4436 2564
rect 4588 2556 4596 2564
rect 4684 2556 4692 2564
rect 4940 2556 4948 2564
rect 4988 2556 4996 2564
rect 5020 2556 5028 2564
rect 828 2536 836 2544
rect 876 2536 884 2544
rect 1020 2536 1028 2544
rect 1180 2536 1188 2544
rect 1212 2536 1220 2544
rect 1276 2536 1284 2544
rect 1372 2536 1380 2544
rect 1420 2536 1428 2544
rect 1532 2536 1540 2544
rect 1548 2536 1556 2544
rect 1596 2536 1604 2544
rect 1692 2536 1700 2544
rect 1756 2536 1764 2544
rect 1868 2536 1876 2544
rect 2588 2536 2596 2544
rect 2812 2536 2820 2544
rect 3100 2536 3108 2544
rect 3196 2536 3204 2544
rect 3212 2536 3220 2544
rect 3276 2536 3284 2544
rect 3308 2536 3316 2544
rect 3484 2536 3492 2544
rect 3500 2536 3508 2544
rect 3628 2536 3636 2544
rect 3740 2536 3748 2544
rect 3836 2536 3844 2544
rect 3884 2536 3892 2544
rect 3916 2536 3924 2544
rect 4156 2536 4164 2544
rect 4300 2536 4308 2544
rect 4396 2536 4404 2544
rect 4620 2536 4628 2544
rect 4652 2536 4660 2544
rect 4812 2536 4820 2544
rect 4876 2536 4884 2544
rect 5020 2536 5028 2544
rect 28 2516 36 2524
rect 60 2496 68 2504
rect 188 2516 196 2524
rect 252 2516 260 2524
rect 268 2516 276 2524
rect 332 2516 340 2524
rect 380 2516 388 2524
rect 460 2516 468 2524
rect 716 2516 724 2524
rect 812 2516 820 2524
rect 972 2516 980 2524
rect 1036 2516 1044 2524
rect 1116 2516 1124 2524
rect 1132 2516 1140 2524
rect 1196 2516 1204 2524
rect 156 2496 164 2504
rect 348 2496 356 2504
rect 412 2496 420 2504
rect 940 2496 948 2504
rect 1164 2496 1172 2504
rect 1612 2516 1620 2524
rect 1628 2516 1636 2524
rect 1756 2516 1764 2524
rect 1772 2516 1780 2524
rect 1868 2516 1876 2524
rect 1900 2516 1908 2524
rect 1932 2516 1940 2524
rect 2060 2516 2068 2524
rect 2124 2518 2132 2526
rect 2252 2516 2260 2524
rect 2300 2516 2308 2524
rect 2412 2516 2420 2524
rect 2556 2518 2564 2526
rect 2684 2516 2692 2524
rect 2748 2518 2756 2526
rect 2892 2516 2900 2524
rect 2972 2516 2980 2524
rect 3036 2518 3044 2526
rect 3244 2516 3252 2524
rect 1644 2496 1652 2504
rect 1820 2496 1828 2504
rect 3212 2496 3220 2504
rect 3324 2516 3332 2524
rect 3340 2516 3348 2524
rect 3372 2516 3380 2524
rect 3436 2516 3444 2524
rect 3532 2516 3540 2524
rect 3564 2516 3572 2524
rect 3612 2516 3620 2524
rect 3804 2518 3812 2526
rect 3868 2516 3876 2524
rect 3900 2516 3908 2524
rect 3932 2516 3940 2524
rect 3980 2516 3988 2524
rect 4092 2516 4100 2524
rect 4316 2518 4324 2526
rect 4380 2516 4388 2524
rect 4524 2516 4532 2524
rect 4556 2516 4564 2524
rect 4604 2516 4612 2524
rect 4668 2516 4676 2524
rect 4716 2516 4724 2524
rect 4748 2516 4756 2524
rect 4860 2516 4868 2524
rect 4972 2516 4980 2524
rect 4988 2516 4996 2524
rect 5020 2516 5028 2524
rect 5132 2536 5140 2544
rect 5148 2536 5156 2544
rect 5244 2536 5252 2544
rect 5356 2536 5364 2544
rect 5436 2536 5444 2544
rect 5628 2536 5636 2544
rect 5852 2536 5860 2544
rect 5420 2518 5428 2526
rect 5564 2516 5572 2524
rect 5660 2518 5668 2526
rect 5804 2516 5812 2524
rect 3340 2496 3348 2504
rect 3452 2496 3460 2504
rect 3580 2496 3588 2504
rect 3644 2496 3652 2504
rect 4540 2496 4548 2504
rect 4684 2496 4692 2504
rect 4780 2496 4788 2504
rect 4828 2496 4836 2504
rect 4860 2496 4868 2504
rect 4892 2496 4900 2504
rect 908 2476 916 2484
rect 988 2476 996 2484
rect 1036 2476 1044 2484
rect 1772 2476 1780 2484
rect 1932 2476 1940 2484
rect 3132 2476 3140 2484
rect 4508 2476 4516 2484
rect 5548 2476 5556 2484
rect 5596 2476 5604 2484
rect 5788 2476 5796 2484
rect 4524 2456 4532 2464
rect 92 2436 100 2444
rect 300 2436 308 2444
rect 380 2436 388 2444
rect 540 2436 548 2444
rect 668 2436 676 2444
rect 972 2436 980 2444
rect 1308 2436 1316 2444
rect 1468 2436 1476 2444
rect 1852 2436 1860 2444
rect 2380 2436 2388 2444
rect 2428 2436 2436 2444
rect 1358 2406 1366 2414
rect 1372 2406 1380 2414
rect 1386 2406 1394 2414
rect 4446 2406 4454 2414
rect 4460 2406 4468 2414
rect 4474 2406 4482 2414
rect 4332 2376 4340 2384
rect 4396 2376 4404 2384
rect 4508 2376 4516 2384
rect 5852 2376 5860 2384
rect 4012 2356 4020 2364
rect 844 2336 852 2344
rect 2396 2336 2404 2344
rect 2588 2336 2596 2344
rect 2972 2336 2980 2344
rect 3580 2336 3588 2344
rect 4220 2336 4228 2344
rect 4412 2336 4420 2344
rect 4428 2336 4436 2344
rect 4556 2336 4564 2344
rect 4860 2336 4868 2344
rect 5084 2336 5092 2344
rect 5276 2336 5284 2344
rect 5324 2336 5332 2344
rect 5516 2336 5524 2344
rect 5708 2336 5716 2344
rect 924 2316 932 2324
rect 1532 2316 1540 2324
rect 140 2294 148 2302
rect 556 2294 564 2302
rect 668 2294 676 2302
rect 1100 2294 1108 2302
rect 1292 2294 1300 2302
rect 1532 2296 1540 2304
rect 1628 2316 1636 2324
rect 2892 2316 2900 2324
rect 3052 2316 3060 2324
rect 3276 2316 3284 2324
rect 3388 2316 3396 2324
rect 4252 2316 4260 2324
rect 4380 2316 4388 2324
rect 4444 2316 4452 2324
rect 4588 2316 4596 2324
rect 4652 2316 4660 2324
rect 4668 2316 4676 2324
rect 1596 2296 1604 2304
rect 1772 2294 1780 2302
rect 1964 2296 1972 2304
rect 2044 2296 2052 2304
rect 2108 2294 2116 2302
rect 2236 2296 2244 2304
rect 2300 2294 2308 2302
rect 2428 2296 2436 2304
rect 2492 2294 2500 2302
rect 2700 2296 2708 2304
rect 2940 2296 2948 2304
rect 3068 2296 3076 2304
rect 3148 2296 3156 2304
rect 3452 2294 3460 2302
rect 3516 2296 3524 2304
rect 3596 2296 3604 2304
rect 3756 2296 3764 2304
rect 3884 2294 3892 2302
rect 3948 2296 3956 2304
rect 4076 2294 4084 2302
rect 4140 2296 4148 2304
rect 4300 2296 4308 2304
rect 124 2276 132 2284
rect 204 2276 212 2284
rect 300 2276 308 2284
rect 316 2276 324 2284
rect 412 2276 420 2284
rect 700 2276 708 2284
rect 812 2276 820 2284
rect 908 2276 916 2284
rect 956 2276 964 2284
rect 1068 2276 1076 2284
rect 1324 2276 1332 2284
rect 1404 2276 1412 2284
rect 1500 2276 1508 2284
rect 1516 2276 1524 2284
rect 1580 2276 1588 2284
rect 1708 2276 1716 2284
rect 1804 2276 1812 2284
rect 1836 2276 1844 2284
rect 2460 2276 2468 2284
rect 2652 2276 2660 2284
rect 2956 2276 2964 2284
rect 3100 2276 3108 2284
rect 3628 2276 3636 2284
rect 4044 2276 4052 2284
rect 4428 2296 4436 2304
rect 4524 2296 4532 2304
rect 4700 2296 4708 2304
rect 4732 2296 4740 2304
rect 4956 2294 4964 2302
rect 5148 2294 5156 2302
rect 5292 2296 5300 2304
rect 5388 2294 5396 2302
rect 5436 2296 5444 2304
rect 5580 2294 5588 2302
rect 5724 2296 5732 2304
rect 5772 2296 5780 2304
rect 4636 2276 4644 2284
rect 4668 2276 4676 2284
rect 4748 2276 4756 2284
rect 4796 2276 4804 2284
rect 4892 2276 4900 2284
rect 4924 2276 4932 2284
rect 5116 2276 5124 2284
rect 5548 2276 5556 2284
rect 5644 2276 5652 2284
rect 5756 2276 5764 2284
rect 556 2256 564 2264
rect 2364 2256 2372 2264
rect 2828 2256 2836 2264
rect 3020 2256 3028 2264
rect 3324 2256 3332 2264
rect 4348 2256 4356 2264
rect 4364 2256 4372 2264
rect 4540 2256 4548 2264
rect 4572 2256 4580 2264
rect 4764 2256 4772 2264
rect 12 2236 20 2244
rect 252 2236 260 2244
rect 348 2236 356 2244
rect 428 2236 436 2244
rect 796 2236 804 2244
rect 924 2236 932 2244
rect 972 2236 980 2244
rect 1164 2236 1172 2244
rect 1436 2236 1444 2244
rect 1628 2236 1636 2244
rect 1644 2236 1652 2244
rect 1980 2236 1988 2244
rect 2172 2236 2180 2244
rect 2380 2236 2388 2244
rect 2620 2236 2628 2244
rect 2812 2236 2820 2244
rect 3260 2236 3268 2244
rect 3292 2236 3300 2244
rect 3388 2236 3396 2244
rect 3644 2236 3652 2244
rect 4284 2236 4292 2244
rect 4604 2236 4612 2244
rect 4700 2236 4708 2244
rect 4780 2236 4788 2244
rect 2910 2206 2918 2214
rect 2924 2206 2932 2214
rect 2938 2206 2946 2214
rect 2204 2176 2212 2184
rect 2716 2176 2724 2184
rect 2844 2176 2852 2184
rect 2988 2176 2996 2184
rect 3644 2176 3652 2184
rect 3884 2176 3892 2184
rect 4076 2176 4084 2184
rect 4412 2176 4420 2184
rect 4556 2176 4564 2184
rect 4860 2176 4868 2184
rect 4956 2176 4964 2184
rect 5100 2176 5108 2184
rect 5212 2176 5220 2184
rect 5420 2176 5428 2184
rect 1740 2156 1748 2164
rect 1884 2156 1892 2164
rect 1916 2156 1924 2164
rect 2252 2156 2260 2164
rect 2732 2156 2740 2164
rect 2924 2156 2932 2164
rect 2940 2156 2948 2164
rect 3420 2156 3428 2164
rect 3660 2156 3668 2164
rect 3804 2156 3812 2164
rect 3932 2156 3940 2164
rect 4380 2156 4388 2164
rect 4428 2156 4436 2164
rect 4572 2156 4580 2164
rect 4652 2156 4660 2164
rect 4876 2156 4884 2164
rect 5292 2156 5300 2164
rect 556 2136 564 2144
rect 940 2136 948 2144
rect 972 2136 980 2144
rect 1100 2136 1108 2144
rect 1276 2136 1284 2144
rect 1324 2136 1332 2144
rect 1772 2136 1780 2144
rect 1820 2136 1828 2144
rect 1932 2136 1940 2144
rect 1964 2136 1972 2144
rect 2044 2136 2052 2144
rect 2300 2136 2308 2144
rect 2348 2136 2356 2144
rect 2412 2136 2420 2144
rect 2460 2136 2468 2144
rect 2476 2136 2484 2144
rect 2812 2136 2820 2144
rect 2876 2136 2884 2144
rect 3100 2136 3108 2144
rect 3180 2136 3188 2144
rect 3484 2136 3492 2144
rect 3756 2136 3764 2144
rect 3820 2136 3828 2144
rect 3932 2136 3940 2144
rect 4012 2136 4020 2144
rect 4028 2136 4036 2144
rect 4124 2136 4132 2144
rect 4156 2136 4164 2144
rect 4364 2136 4372 2144
rect 4492 2136 4500 2144
rect 4588 2136 4596 2144
rect 4652 2136 4660 2144
rect 4684 2136 4692 2144
rect 4764 2136 4772 2144
rect 4828 2136 4836 2144
rect 4892 2136 4900 2144
rect 4908 2136 4916 2144
rect 4972 2136 4980 2144
rect 4988 2136 4996 2144
rect 5004 2136 5012 2144
rect 5020 2136 5028 2144
rect 5132 2136 5140 2144
rect 5148 2136 5156 2144
rect 5244 2136 5252 2144
rect 5276 2136 5284 2144
rect 5324 2136 5332 2144
rect 5372 2136 5380 2144
rect 60 2118 68 2126
rect 124 2116 132 2124
rect 268 2116 276 2124
rect 316 2116 324 2124
rect 524 2118 532 2126
rect 652 2116 660 2124
rect 700 2116 708 2124
rect 908 2118 916 2126
rect 1180 2116 1188 2124
rect 1244 2118 1252 2126
rect 1436 2116 1444 2124
rect 1468 2116 1476 2124
rect 1628 2116 1636 2124
rect 1660 2116 1668 2124
rect 1836 2116 1844 2124
rect 1884 2116 1892 2124
rect 1916 2116 1924 2124
rect 1980 2116 1988 2124
rect 2076 2118 2084 2126
rect 2220 2116 2228 2124
rect 2268 2116 2276 2124
rect 2364 2116 2372 2124
rect 2428 2116 2436 2124
rect 2492 2116 2500 2124
rect 2588 2118 2596 2126
rect 2652 2116 2660 2124
rect 2796 2116 2804 2124
rect 2844 2116 2852 2124
rect 3052 2116 3060 2124
rect 3116 2118 3124 2126
rect 3212 2116 3220 2124
rect 3292 2116 3300 2124
rect 3356 2118 3364 2126
rect 3452 2116 3460 2124
rect 3516 2118 3524 2126
rect 3580 2116 3588 2124
rect 3708 2116 3716 2124
rect 3772 2116 3780 2124
rect 3964 2116 3972 2124
rect 3996 2116 4004 2124
rect 4188 2118 4196 2126
rect 4252 2116 4260 2124
rect 4332 2116 4340 2124
rect 4396 2116 4404 2124
rect 4604 2116 4612 2124
rect 4700 2116 4708 2124
rect 4764 2116 4772 2124
rect 4780 2116 4788 2124
rect 4828 2116 4836 2124
rect 4924 2116 4932 2124
rect 4956 2116 4964 2124
rect 5244 2116 5252 2124
rect 5372 2116 5380 2124
rect 5644 2136 5652 2144
rect 5676 2136 5684 2144
rect 5484 2118 5492 2126
rect 5548 2116 5556 2124
rect 5692 2116 5700 2124
rect 5820 2116 5828 2124
rect 1868 2096 1876 2104
rect 2012 2096 2020 2104
rect 2396 2096 2404 2104
rect 2460 2096 2468 2104
rect 2524 2096 2532 2104
rect 2844 2096 2852 2104
rect 3740 2096 3748 2104
rect 3804 2096 3812 2104
rect 3964 2096 3972 2104
rect 3996 2096 4004 2104
rect 4524 2096 4532 2104
rect 4636 2096 4644 2104
rect 4652 2096 4660 2104
rect 4748 2096 4756 2104
rect 4812 2096 4820 2104
rect 4860 2096 4868 2104
rect 5020 2096 5028 2104
rect 5340 2096 5348 2104
rect 5388 2096 5396 2104
rect 5420 2096 5428 2104
rect 1932 2076 1940 2084
rect 2172 2076 2180 2084
rect 2332 2076 2340 2084
rect 2492 2076 2500 2084
rect 2812 2076 2820 2084
rect 3228 2076 3236 2084
rect 3708 2076 3716 2084
rect 4316 2076 4324 2084
rect 5612 2076 5620 2084
rect 5804 2076 5812 2084
rect 5852 2076 5860 2084
rect 188 2036 196 2044
rect 380 2036 388 2044
rect 396 2036 404 2044
rect 764 2036 772 2044
rect 780 2036 788 2044
rect 1116 2036 1124 2044
rect 1532 2036 1540 2044
rect 1724 2036 1732 2044
rect 1804 2036 1812 2044
rect 1980 2036 1988 2044
rect 1358 2006 1366 2014
rect 1372 2006 1380 2014
rect 1386 2006 1394 2014
rect 4446 2006 4454 2014
rect 4460 2006 4468 2014
rect 4474 2006 4482 2014
rect 2652 1976 2660 1984
rect 3260 1976 3268 1984
rect 3516 1976 3524 1984
rect 3740 1976 3748 1984
rect 3804 1976 3812 1984
rect 3932 1976 3940 1984
rect 4028 1976 4036 1984
rect 4092 1976 4100 1984
rect 4508 1976 4516 1984
rect 4716 1976 4724 1984
rect 4972 1976 4980 1984
rect 5052 1976 5060 1984
rect 5244 1976 5252 1984
rect 5340 1976 5348 1984
rect 5372 1976 5380 1984
rect 2028 1936 2036 1944
rect 3068 1936 3076 1944
rect 5324 1936 5332 1944
rect 396 1916 404 1924
rect 492 1916 500 1924
rect 556 1916 564 1924
rect 604 1916 612 1924
rect 652 1916 660 1924
rect 780 1916 788 1924
rect 860 1916 868 1924
rect 876 1916 884 1924
rect 92 1896 100 1904
rect 124 1896 132 1904
rect 252 1894 260 1902
rect 316 1896 324 1904
rect 540 1896 548 1904
rect 636 1896 644 1904
rect 684 1896 692 1904
rect 940 1896 948 1904
rect 1036 1916 1044 1924
rect 1100 1916 1108 1924
rect 1884 1916 1892 1924
rect 1916 1916 1924 1924
rect 1292 1896 1300 1904
rect 1516 1894 1524 1902
rect 1564 1896 1572 1904
rect 1756 1896 1764 1904
rect 1916 1896 1924 1904
rect 1996 1916 2004 1924
rect 2060 1916 2068 1924
rect 2444 1916 2452 1924
rect 2556 1916 2564 1924
rect 2732 1916 2740 1924
rect 3020 1916 3028 1924
rect 3116 1916 3124 1924
rect 3212 1916 3220 1924
rect 3388 1916 3396 1924
rect 3436 1916 3444 1924
rect 2028 1896 2036 1904
rect 2172 1896 2180 1904
rect 2300 1894 2308 1902
rect 2476 1896 2484 1904
rect 2508 1896 2516 1904
rect 2796 1894 2804 1902
rect 3036 1896 3044 1904
rect 3148 1896 3156 1904
rect 3356 1896 3364 1904
rect 3612 1894 3620 1902
rect 3772 1896 3780 1904
rect 3820 1896 3828 1904
rect 3836 1896 3844 1904
rect 4908 1916 4916 1924
rect 5116 1916 5124 1924
rect 5180 1916 5188 1924
rect 3884 1896 3892 1904
rect 428 1876 436 1884
rect 460 1876 468 1884
rect 636 1876 644 1884
rect 700 1876 708 1884
rect 716 1876 724 1884
rect 732 1880 740 1888
rect 924 1876 932 1884
rect 972 1876 980 1884
rect 1084 1876 1092 1884
rect 1132 1876 1140 1884
rect 444 1856 452 1864
rect 508 1856 516 1864
rect 780 1856 788 1864
rect 876 1856 884 1864
rect 940 1856 948 1864
rect 1212 1876 1220 1884
rect 1276 1876 1284 1884
rect 1708 1876 1716 1884
rect 1932 1876 1940 1884
rect 1980 1876 1988 1884
rect 2044 1876 2052 1884
rect 2236 1876 2244 1884
rect 2268 1876 2276 1884
rect 2348 1876 2356 1884
rect 2460 1876 2468 1884
rect 2492 1876 2500 1884
rect 2588 1876 2596 1884
rect 2684 1876 2692 1884
rect 2764 1876 2772 1884
rect 2988 1876 2996 1884
rect 3084 1876 3092 1884
rect 3100 1876 3108 1884
rect 3132 1876 3140 1884
rect 3180 1876 3188 1884
rect 3228 1876 3236 1884
rect 3324 1876 3332 1884
rect 3420 1876 3428 1884
rect 3452 1876 3460 1884
rect 3548 1876 3556 1884
rect 3580 1876 3588 1884
rect 3852 1876 3860 1884
rect 3900 1876 3908 1884
rect 3964 1896 3972 1904
rect 4076 1896 4084 1904
rect 4204 1896 4212 1904
rect 4332 1894 4340 1902
rect 4524 1896 4532 1904
rect 4620 1896 4628 1904
rect 4780 1896 4788 1904
rect 4876 1896 4884 1904
rect 4924 1896 4932 1904
rect 5164 1896 5172 1904
rect 5388 1916 5396 1924
rect 5484 1916 5492 1924
rect 5452 1896 5460 1904
rect 5500 1896 5508 1904
rect 5580 1896 5588 1904
rect 5708 1894 5716 1902
rect 4252 1876 4260 1884
rect 4540 1876 4548 1884
rect 4604 1876 4612 1884
rect 4636 1876 4644 1884
rect 4652 1876 4660 1884
rect 4748 1876 4756 1884
rect 4764 1876 4772 1884
rect 4812 1876 4820 1884
rect 4860 1876 4868 1884
rect 4988 1876 4996 1884
rect 5084 1876 5092 1884
rect 5212 1876 5220 1884
rect 5276 1876 5284 1884
rect 5308 1876 5316 1884
rect 5356 1876 5364 1884
rect 5420 1876 5428 1884
rect 5484 1876 5492 1884
rect 5644 1876 5652 1884
rect 5676 1876 5684 1884
rect 1852 1856 1860 1864
rect 2124 1856 2132 1864
rect 2508 1856 2516 1864
rect 2572 1856 2580 1864
rect 3916 1856 3924 1864
rect 3996 1856 4004 1864
rect 4012 1856 4020 1864
rect 4044 1856 4052 1864
rect 4076 1856 4084 1864
rect 4332 1856 4340 1864
rect 4572 1856 4580 1864
rect 4844 1856 4852 1864
rect 4972 1856 4980 1864
rect 5100 1856 5108 1864
rect 5132 1856 5140 1864
rect 5244 1856 5252 1864
rect 5324 1856 5332 1864
rect 5532 1856 5540 1864
rect 188 1836 196 1844
rect 380 1836 388 1844
rect 396 1836 404 1844
rect 524 1836 532 1844
rect 572 1836 580 1844
rect 620 1836 628 1844
rect 764 1836 772 1844
rect 812 1836 820 1844
rect 1020 1836 1028 1844
rect 1116 1836 1124 1844
rect 1196 1836 1204 1844
rect 1452 1836 1460 1844
rect 1644 1836 1652 1844
rect 1836 1836 1844 1844
rect 1868 1836 1876 1844
rect 1964 1836 1972 1844
rect 2076 1836 2084 1844
rect 2428 1836 2436 1844
rect 2732 1836 2740 1844
rect 2924 1836 2932 1844
rect 3212 1836 3220 1844
rect 3740 1836 3748 1844
rect 5148 1836 5156 1844
rect 5180 1836 5188 1844
rect 5404 1836 5412 1844
rect 5836 1836 5844 1844
rect 2910 1806 2918 1814
rect 2924 1806 2932 1814
rect 2938 1806 2946 1814
rect 3084 1776 3092 1784
rect 3260 1776 3268 1784
rect 3516 1776 3524 1784
rect 3724 1776 3732 1784
rect 3788 1776 3796 1784
rect 3836 1776 3844 1784
rect 3948 1776 3956 1784
rect 4156 1776 4164 1784
rect 4396 1776 4404 1784
rect 4748 1776 4756 1784
rect 4764 1776 4772 1784
rect 4860 1776 4868 1784
rect 4924 1776 4932 1784
rect 5004 1776 5012 1784
rect 5084 1776 5092 1784
rect 5196 1776 5204 1784
rect 556 1756 564 1764
rect 716 1756 724 1764
rect 2012 1756 2020 1764
rect 2076 1756 2084 1764
rect 2092 1756 2100 1764
rect 3404 1756 3412 1764
rect 3564 1756 3572 1764
rect 124 1736 132 1744
rect 140 1718 148 1726
rect 220 1716 228 1724
rect 236 1716 244 1724
rect 268 1736 276 1744
rect 380 1736 388 1744
rect 476 1736 484 1744
rect 540 1736 548 1744
rect 588 1736 596 1744
rect 668 1736 676 1744
rect 700 1736 708 1744
rect 828 1736 836 1744
rect 924 1736 932 1744
rect 940 1736 948 1744
rect 1036 1736 1044 1744
rect 1068 1736 1076 1744
rect 1244 1736 1252 1744
rect 1548 1736 1556 1744
rect 1724 1736 1732 1744
rect 1820 1736 1828 1744
rect 1836 1736 1844 1744
rect 1900 1736 1908 1744
rect 1932 1736 1940 1744
rect 2044 1736 2052 1744
rect 2108 1736 2116 1744
rect 2220 1736 2228 1744
rect 2236 1736 2244 1744
rect 2348 1736 2356 1744
rect 2492 1736 2500 1744
rect 2524 1736 2532 1744
rect 2652 1736 2660 1744
rect 2684 1736 2692 1744
rect 2764 1736 2772 1744
rect 2924 1736 2932 1744
rect 3132 1736 3140 1744
rect 476 1716 484 1724
rect 524 1716 532 1724
rect 604 1716 612 1724
rect 636 1716 644 1724
rect 652 1716 660 1724
rect 700 1716 708 1724
rect 748 1716 756 1724
rect 764 1716 772 1724
rect 876 1716 884 1724
rect 1100 1718 1108 1726
rect 1324 1716 1332 1724
rect 1388 1718 1396 1726
rect 1452 1716 1460 1724
rect 1580 1718 1588 1726
rect 1644 1716 1652 1724
rect 1852 1716 1860 1724
rect 1868 1716 1876 1724
rect 204 1696 212 1704
rect 492 1696 500 1704
rect 620 1696 628 1704
rect 812 1696 820 1704
rect 1276 1696 1284 1704
rect 1964 1716 1972 1724
rect 1980 1716 1988 1724
rect 2028 1716 2036 1724
rect 2124 1716 2132 1724
rect 2156 1716 2164 1724
rect 2204 1716 2212 1724
rect 2380 1718 2388 1726
rect 2716 1718 2724 1726
rect 2956 1718 2964 1726
rect 3212 1736 3220 1744
rect 3244 1736 3252 1744
rect 3308 1736 3316 1744
rect 3372 1736 3380 1744
rect 3420 1736 3428 1744
rect 3484 1736 3492 1744
rect 3628 1756 3636 1764
rect 3644 1756 3652 1764
rect 3692 1756 3700 1764
rect 3660 1736 3668 1744
rect 3772 1756 3780 1764
rect 3932 1756 3940 1764
rect 4092 1756 4100 1764
rect 5292 1756 5300 1764
rect 5420 1756 5428 1764
rect 5436 1756 5444 1764
rect 5532 1756 5540 1764
rect 5564 1756 5572 1764
rect 3740 1736 3748 1744
rect 3820 1736 3828 1744
rect 3868 1736 3876 1744
rect 3964 1736 3972 1744
rect 4060 1736 4068 1744
rect 4108 1736 4116 1744
rect 4204 1736 4212 1744
rect 4332 1736 4340 1744
rect 4460 1736 4468 1744
rect 4556 1736 4564 1744
rect 4588 1736 4596 1744
rect 4796 1736 4804 1744
rect 4892 1736 4900 1744
rect 4908 1736 4916 1744
rect 4940 1736 4948 1744
rect 5052 1736 5060 1744
rect 5068 1736 5076 1744
rect 5132 1736 5140 1744
rect 5164 1736 5172 1744
rect 5244 1736 5252 1744
rect 5340 1736 5348 1744
rect 3164 1716 3172 1724
rect 1996 1696 2004 1704
rect 2156 1696 2164 1704
rect 2172 1696 2180 1704
rect 2268 1696 2276 1704
rect 2300 1696 2308 1704
rect 2316 1696 2324 1704
rect 3100 1696 3108 1704
rect 3196 1696 3204 1704
rect 3436 1716 3444 1724
rect 3484 1716 3492 1724
rect 3532 1716 3540 1724
rect 3612 1716 3620 1724
rect 3756 1716 3764 1724
rect 3804 1716 3812 1724
rect 3884 1716 3892 1724
rect 3900 1716 3908 1724
rect 4124 1716 4132 1724
rect 4268 1718 4276 1726
rect 3260 1696 3268 1704
rect 3324 1696 3332 1704
rect 3356 1696 3364 1704
rect 3468 1696 3476 1704
rect 3516 1696 3524 1704
rect 3852 1696 3860 1704
rect 3916 1696 3924 1704
rect 3964 1696 3972 1704
rect 3996 1696 4004 1704
rect 4012 1696 4020 1704
rect 4316 1716 4324 1724
rect 4524 1716 4532 1724
rect 4620 1718 4628 1726
rect 4684 1716 4692 1724
rect 4172 1696 4180 1704
rect 4988 1696 4996 1704
rect 5036 1716 5044 1724
rect 5116 1716 5124 1724
rect 5180 1716 5188 1724
rect 5228 1716 5236 1724
rect 5292 1716 5300 1724
rect 5388 1716 5396 1724
rect 5420 1716 5428 1724
rect 5452 1716 5460 1724
rect 5484 1716 5492 1724
rect 5500 1716 5508 1724
rect 5532 1716 5540 1724
rect 5660 1716 5668 1724
rect 5692 1716 5700 1724
rect 5772 1716 5780 1724
rect 5100 1696 5108 1704
rect 5196 1696 5204 1704
rect 5308 1696 5316 1704
rect 5404 1696 5412 1704
rect 5468 1696 5476 1704
rect 332 1676 340 1684
rect 780 1676 788 1684
rect 2204 1676 2212 1684
rect 2844 1676 2852 1684
rect 3052 1676 3060 1684
rect 3612 1676 3620 1684
rect 5132 1676 5140 1684
rect 5372 1676 5380 1684
rect 5500 1676 5508 1684
rect 5756 1676 5764 1684
rect 5852 1676 5860 1684
rect 444 1656 452 1664
rect 1788 1656 1796 1664
rect 5276 1656 5284 1664
rect 12 1636 20 1644
rect 556 1636 564 1644
rect 1004 1636 1012 1644
rect 1228 1636 1236 1644
rect 1516 1636 1524 1644
rect 1708 1636 1716 1644
rect 2508 1636 2516 1644
rect 3980 1636 3988 1644
rect 4044 1636 4052 1644
rect 5356 1636 5364 1644
rect 5516 1636 5524 1644
rect 1358 1606 1366 1614
rect 1372 1606 1380 1614
rect 1386 1606 1394 1614
rect 4446 1606 4454 1614
rect 4460 1606 4468 1614
rect 4474 1606 4482 1614
rect 204 1576 212 1584
rect 412 1576 420 1584
rect 3564 1576 3572 1584
rect 4188 1576 4196 1584
rect 4476 1576 4484 1584
rect 4860 1576 4868 1584
rect 5484 1576 5492 1584
rect 5596 1576 5604 1584
rect 748 1536 756 1544
rect 1068 1536 1076 1544
rect 2396 1536 2404 1544
rect 3084 1536 3092 1544
rect 5388 1536 5396 1544
rect 124 1516 132 1524
rect 188 1516 196 1524
rect 332 1516 340 1524
rect 492 1516 500 1524
rect 540 1516 548 1524
rect 604 1516 612 1524
rect 668 1516 676 1524
rect 1036 1516 1044 1524
rect 2092 1516 2100 1524
rect 2556 1516 2564 1524
rect 2716 1516 2724 1524
rect 3516 1516 3524 1524
rect 28 1496 36 1504
rect 156 1496 164 1504
rect 252 1496 260 1504
rect 284 1496 292 1504
rect 316 1496 324 1504
rect 364 1496 372 1504
rect 412 1496 420 1504
rect 556 1496 564 1504
rect 796 1496 804 1504
rect 860 1496 868 1504
rect 876 1496 884 1504
rect 972 1496 980 1504
rect 1148 1496 1156 1504
rect 1228 1496 1236 1504
rect 1292 1496 1300 1504
rect 1356 1496 1364 1504
rect 1580 1494 1588 1502
rect 1644 1496 1652 1504
rect 1724 1496 1732 1504
rect 2252 1496 2260 1504
rect 2636 1496 2644 1504
rect 2668 1496 2676 1504
rect 2700 1496 2708 1504
rect 2748 1496 2756 1504
rect 2812 1496 2820 1504
rect 2988 1494 2996 1502
rect 3052 1496 3060 1504
rect 3180 1494 3188 1502
rect 3484 1496 3492 1504
rect 3676 1516 3684 1524
rect 3740 1516 3748 1524
rect 3804 1516 3812 1524
rect 3820 1516 3828 1524
rect 3852 1516 3860 1524
rect 3884 1516 3892 1524
rect 4620 1516 4628 1524
rect 3564 1496 3572 1504
rect 3644 1496 3652 1504
rect 3676 1496 3684 1504
rect 3708 1496 3716 1504
rect 3756 1496 3764 1504
rect 3852 1496 3860 1504
rect 3916 1496 3924 1504
rect 3980 1496 3988 1504
rect 4044 1496 4052 1504
rect 4060 1496 4068 1504
rect 4124 1496 4132 1504
rect 4140 1496 4148 1504
rect 4156 1496 4164 1504
rect 4204 1496 4212 1504
rect 4284 1496 4292 1504
rect 4396 1496 4404 1504
rect 4508 1496 4516 1504
rect 4588 1496 4596 1504
rect 5020 1516 5028 1524
rect 5212 1516 5220 1524
rect 5244 1516 5252 1524
rect 5308 1516 5316 1524
rect 5420 1516 5428 1524
rect 5468 1516 5476 1524
rect 4668 1496 4676 1504
rect 4732 1494 4740 1502
rect 4780 1496 4788 1504
rect 4876 1496 4884 1504
rect 5068 1496 5076 1504
rect 5132 1496 5140 1504
rect 5164 1496 5172 1504
rect 5276 1496 5284 1504
rect 5292 1496 5300 1504
rect 5340 1496 5348 1504
rect 5356 1496 5364 1504
rect 5404 1496 5412 1504
rect 5484 1496 5492 1504
rect 5708 1496 5716 1504
rect 12 1476 20 1484
rect 92 1476 100 1484
rect 140 1476 148 1484
rect 236 1476 244 1484
rect 300 1476 308 1484
rect 380 1476 388 1484
rect 396 1476 404 1484
rect 460 1476 468 1484
rect 508 1476 516 1484
rect 556 1476 564 1484
rect 620 1476 628 1484
rect 684 1476 692 1484
rect 780 1476 788 1484
rect 812 1476 820 1484
rect 844 1476 852 1484
rect 892 1476 900 1484
rect 924 1476 932 1484
rect 1068 1476 1076 1484
rect 1116 1476 1124 1484
rect 1212 1476 1220 1484
rect 1340 1476 1348 1484
rect 1420 1476 1428 1484
rect 1852 1476 1860 1484
rect 1964 1476 1972 1484
rect 1980 1476 1988 1484
rect 2076 1476 2084 1484
rect 2124 1476 2132 1484
rect 2140 1476 2148 1484
rect 2236 1476 2244 1484
rect 2316 1476 2324 1484
rect 2428 1476 2436 1484
rect 2460 1476 2468 1484
rect 2572 1476 2580 1484
rect 2588 1476 2596 1484
rect 76 1456 84 1464
rect 188 1456 196 1464
rect 204 1456 212 1464
rect 268 1456 276 1464
rect 668 1456 676 1464
rect 972 1456 980 1464
rect 988 1456 996 1464
rect 1100 1456 1108 1464
rect 1276 1456 1284 1464
rect 1340 1456 1348 1464
rect 2284 1456 2292 1464
rect 2316 1456 2324 1464
rect 2444 1456 2452 1464
rect 2652 1476 2660 1484
rect 2732 1476 2740 1484
rect 2764 1476 2772 1484
rect 2780 1476 2788 1484
rect 2876 1476 2884 1484
rect 3148 1476 3156 1484
rect 3324 1476 3332 1484
rect 3468 1476 3476 1484
rect 3628 1476 3636 1484
rect 3692 1476 3700 1484
rect 3756 1476 3764 1484
rect 3804 1476 3812 1484
rect 3868 1476 3876 1484
rect 3900 1476 3908 1484
rect 3932 1476 3940 1484
rect 4028 1476 4036 1484
rect 4108 1476 4116 1484
rect 4252 1476 4260 1484
rect 4284 1476 4292 1484
rect 4444 1476 4452 1484
rect 4668 1476 4676 1484
rect 4700 1476 4708 1484
rect 5004 1476 5012 1484
rect 5052 1476 5060 1484
rect 5084 1476 5092 1484
rect 5116 1476 5124 1484
rect 5148 1476 5156 1484
rect 5260 1476 5268 1484
rect 5404 1476 5412 1484
rect 5436 1476 5444 1484
rect 5516 1476 5524 1484
rect 5628 1476 5636 1484
rect 5692 1476 5700 1484
rect 2636 1456 2644 1464
rect 3612 1456 3620 1464
rect 3740 1456 3748 1464
rect 3948 1456 3956 1464
rect 4108 1456 4116 1464
rect 4284 1456 4292 1464
rect 4316 1456 4324 1464
rect 4332 1456 4340 1464
rect 4492 1456 4500 1464
rect 4556 1456 4564 1464
rect 5324 1456 5332 1464
rect 5516 1456 5524 1464
rect 60 1436 68 1444
rect 220 1436 228 1444
rect 332 1436 340 1444
rect 540 1436 548 1444
rect 828 1436 836 1444
rect 908 1436 916 1444
rect 1036 1436 1044 1444
rect 1484 1436 1492 1444
rect 1708 1436 1716 1444
rect 1932 1436 1940 1444
rect 2092 1436 2100 1444
rect 2204 1436 2212 1444
rect 2268 1436 2276 1444
rect 2300 1436 2308 1444
rect 2508 1436 2516 1444
rect 3116 1436 3124 1444
rect 3308 1436 3316 1444
rect 3436 1436 3444 1444
rect 3996 1436 4004 1444
rect 4364 1436 4372 1444
rect 5100 1436 5108 1444
rect 5244 1436 5252 1444
rect 5452 1436 5460 1444
rect 5836 1436 5844 1444
rect 2910 1406 2918 1414
rect 2924 1406 2932 1414
rect 2938 1406 2946 1414
rect 268 1376 276 1384
rect 444 1376 452 1384
rect 492 1376 500 1384
rect 604 1376 612 1384
rect 1212 1376 1220 1384
rect 1292 1376 1300 1384
rect 2012 1376 2020 1384
rect 2428 1376 2436 1384
rect 2764 1376 2772 1384
rect 3244 1376 3252 1384
rect 3708 1376 3716 1384
rect 3804 1376 3812 1384
rect 3868 1376 3876 1384
rect 3932 1376 3940 1384
rect 4012 1376 4020 1384
rect 4108 1376 4116 1384
rect 4268 1376 4276 1384
rect 4492 1376 4500 1384
rect 4540 1376 4548 1384
rect 4620 1376 4628 1384
rect 4748 1376 4756 1384
rect 4796 1376 4804 1384
rect 5148 1376 5156 1384
rect 5212 1376 5220 1384
rect 5340 1376 5348 1384
rect 5404 1376 5412 1384
rect 5708 1376 5716 1384
rect 12 1356 20 1364
rect 76 1356 84 1364
rect 156 1356 164 1364
rect 284 1356 292 1364
rect 300 1356 308 1364
rect 332 1356 340 1364
rect 348 1356 356 1364
rect 908 1356 916 1364
rect 1100 1356 1108 1364
rect 1644 1356 1652 1364
rect 1884 1356 1892 1364
rect 2060 1356 2068 1364
rect 92 1336 100 1344
rect 380 1336 388 1344
rect 44 1316 52 1324
rect 108 1316 116 1324
rect 204 1316 212 1324
rect 236 1316 244 1324
rect 252 1316 260 1324
rect 300 1316 308 1324
rect 476 1336 484 1344
rect 524 1336 532 1344
rect 572 1336 580 1344
rect 588 1336 596 1344
rect 652 1336 660 1344
rect 764 1336 772 1344
rect 828 1336 836 1344
rect 876 1336 884 1344
rect 924 1336 932 1344
rect 1036 1336 1044 1344
rect 1084 1336 1092 1344
rect 1148 1336 1156 1344
rect 1164 1336 1172 1344
rect 1260 1336 1268 1344
rect 1308 1336 1316 1344
rect 1468 1336 1476 1344
rect 1484 1336 1492 1344
rect 1580 1336 1588 1344
rect 1788 1336 1796 1344
rect 1916 1336 1924 1344
rect 1980 1336 1988 1344
rect 140 1296 148 1304
rect 380 1296 388 1304
rect 412 1296 420 1304
rect 684 1316 692 1324
rect 732 1316 740 1324
rect 748 1316 756 1324
rect 780 1316 788 1324
rect 508 1296 516 1304
rect 572 1296 580 1304
rect 620 1296 628 1304
rect 812 1296 820 1304
rect 940 1316 948 1324
rect 972 1296 980 1304
rect 1148 1316 1156 1324
rect 1052 1296 1060 1304
rect 1196 1296 1204 1304
rect 1260 1316 1268 1324
rect 1644 1318 1652 1326
rect 1916 1316 1924 1324
rect 1932 1316 1940 1324
rect 2108 1316 2116 1324
rect 2140 1336 2148 1344
rect 2252 1336 2260 1344
rect 2268 1336 2276 1344
rect 2316 1336 2324 1344
rect 2332 1336 2340 1344
rect 2508 1336 2516 1344
rect 2556 1356 2564 1364
rect 2588 1356 2596 1364
rect 2812 1356 2820 1364
rect 3692 1356 3700 1364
rect 3772 1356 3780 1364
rect 3788 1356 3796 1364
rect 3980 1356 3988 1364
rect 4188 1356 4196 1364
rect 4524 1356 4532 1364
rect 5388 1356 5396 1364
rect 5500 1356 5508 1364
rect 2700 1336 2708 1344
rect 2812 1336 2820 1344
rect 2844 1336 2852 1344
rect 2940 1336 2948 1344
rect 2956 1336 2964 1344
rect 3052 1336 3060 1344
rect 3084 1336 3092 1344
rect 3148 1336 3156 1344
rect 3260 1336 3268 1344
rect 3356 1336 3364 1344
rect 3372 1336 3380 1344
rect 3484 1336 3492 1344
rect 3580 1336 3588 1344
rect 2140 1316 2148 1324
rect 2156 1316 2164 1324
rect 1276 1296 1284 1304
rect 1820 1296 1828 1304
rect 1852 1296 1860 1304
rect 1884 1296 1892 1304
rect 1964 1296 1972 1304
rect 2012 1296 2020 1304
rect 2076 1296 2084 1304
rect 2188 1296 2196 1304
rect 2236 1316 2244 1324
rect 2284 1316 2292 1324
rect 2348 1316 2356 1324
rect 2460 1316 2468 1324
rect 2476 1316 2484 1324
rect 2492 1316 2500 1324
rect 2524 1316 2532 1324
rect 2652 1316 2660 1324
rect 2684 1316 2692 1324
rect 3116 1318 3124 1326
rect 3548 1316 3556 1324
rect 3580 1316 3588 1324
rect 3724 1336 3732 1344
rect 3756 1336 3764 1344
rect 3852 1336 3860 1344
rect 3884 1336 3892 1344
rect 3900 1336 3908 1344
rect 4044 1336 4052 1344
rect 4204 1336 4212 1344
rect 4300 1336 4308 1344
rect 4332 1336 4340 1344
rect 4380 1336 4388 1344
rect 4572 1336 4580 1344
rect 4668 1336 4676 1344
rect 4956 1336 4964 1344
rect 4988 1336 4996 1344
rect 5132 1336 5140 1344
rect 5228 1336 5236 1344
rect 5276 1336 5284 1344
rect 5324 1336 5332 1344
rect 5436 1336 5444 1344
rect 5484 1336 5492 1344
rect 5564 1336 5572 1344
rect 5660 1336 5668 1344
rect 5676 1336 5684 1344
rect 5772 1336 5780 1344
rect 3996 1316 4004 1324
rect 4060 1316 4068 1324
rect 4076 1316 4084 1324
rect 4140 1316 4148 1324
rect 4156 1316 4164 1324
rect 4348 1316 4356 1324
rect 4412 1316 4420 1324
rect 4588 1316 4596 1324
rect 4684 1316 4692 1324
rect 4716 1316 4724 1324
rect 4748 1316 4756 1324
rect 4908 1316 4916 1324
rect 5548 1316 5556 1324
rect 5788 1316 5796 1324
rect 2316 1296 2324 1304
rect 2380 1296 2388 1304
rect 2684 1296 2692 1304
rect 2716 1296 2724 1304
rect 2748 1296 2756 1304
rect 2764 1296 2772 1304
rect 2892 1296 2900 1304
rect 3436 1296 3444 1304
rect 3644 1296 3652 1304
rect 3676 1296 3684 1304
rect 3804 1296 3812 1304
rect 3836 1296 3844 1304
rect 3932 1296 3940 1304
rect 4316 1296 4324 1304
rect 4636 1296 4644 1304
rect 4652 1296 4660 1304
rect 4716 1296 4724 1304
rect 4732 1296 4740 1304
rect 5164 1296 5172 1304
rect 5260 1296 5268 1304
rect 5356 1296 5364 1304
rect 5404 1296 5412 1304
rect 5436 1296 5444 1304
rect 12 1276 20 1284
rect 1740 1276 1748 1284
rect 2108 1276 2116 1284
rect 3660 1276 3668 1284
rect 4764 1276 4772 1284
rect 5532 1276 5540 1284
rect 5804 1276 5812 1284
rect 3324 1256 3332 1264
rect 44 1236 52 1244
rect 108 1236 116 1244
rect 220 1236 228 1244
rect 636 1236 644 1244
rect 716 1236 724 1244
rect 1020 1236 1028 1244
rect 1420 1236 1428 1244
rect 1516 1236 1524 1244
rect 1772 1236 1780 1244
rect 1932 1236 1940 1244
rect 2044 1236 2052 1244
rect 2236 1236 2244 1244
rect 2652 1236 2660 1244
rect 3020 1236 3028 1244
rect 3820 1236 3828 1244
rect 5100 1236 5108 1244
rect 5292 1236 5300 1244
rect 5596 1236 5604 1244
rect 1358 1206 1366 1214
rect 1372 1206 1380 1214
rect 1386 1206 1394 1214
rect 4446 1206 4454 1214
rect 4460 1206 4468 1214
rect 4474 1206 4482 1214
rect 1180 1176 1188 1184
rect 2524 1176 2532 1184
rect 3068 1176 3076 1184
rect 3452 1176 3460 1184
rect 3484 1176 3492 1184
rect 3564 1176 3572 1184
rect 4172 1176 4180 1184
rect 4492 1176 4500 1184
rect 4572 1176 4580 1184
rect 4636 1176 4644 1184
rect 5020 1176 5028 1184
rect 5212 1176 5220 1184
rect 5820 1176 5828 1184
rect 1372 1156 1380 1164
rect 780 1136 788 1144
rect 1820 1136 1828 1144
rect 1884 1136 1892 1144
rect 2892 1136 2900 1144
rect 3628 1136 3636 1144
rect 5180 1136 5188 1144
rect 5628 1136 5636 1144
rect 60 1116 68 1124
rect 460 1116 468 1124
rect 924 1116 932 1124
rect 1084 1116 1092 1124
rect 1148 1116 1156 1124
rect 1212 1116 1220 1124
rect 1916 1116 1924 1124
rect 1964 1116 1972 1124
rect 2108 1116 2116 1124
rect 2300 1116 2308 1124
rect 2332 1116 2340 1124
rect 2604 1116 2612 1124
rect 2748 1116 2756 1124
rect 2812 1116 2820 1124
rect 3708 1116 3716 1124
rect 3820 1116 3828 1124
rect 3900 1116 3908 1124
rect 3932 1116 3940 1124
rect 3948 1116 3956 1124
rect 4124 1116 4132 1124
rect 4140 1116 4148 1124
rect 28 1096 36 1104
rect 76 1096 84 1104
rect 140 1096 148 1104
rect 220 1096 228 1104
rect 316 1096 324 1104
rect 364 1096 372 1104
rect 428 1096 436 1104
rect 444 1096 452 1104
rect 508 1096 516 1104
rect 604 1096 612 1104
rect 700 1096 708 1104
rect 844 1096 852 1104
rect 892 1096 900 1104
rect 972 1096 980 1104
rect 988 1096 996 1104
rect 1052 1096 1060 1104
rect 1116 1096 1124 1104
rect 1164 1096 1172 1104
rect 1276 1096 1284 1104
rect 1308 1096 1316 1104
rect 1340 1096 1348 1104
rect 1484 1096 1492 1104
rect 1564 1096 1572 1104
rect 1692 1094 1700 1102
rect 1740 1096 1748 1104
rect 2012 1096 2020 1104
rect 2028 1096 2036 1104
rect 2092 1096 2100 1104
rect 2172 1096 2180 1104
rect 2204 1096 2212 1104
rect 2220 1096 2228 1104
rect 2284 1096 2292 1104
rect 2332 1096 2340 1104
rect 2348 1096 2356 1104
rect 2428 1096 2436 1104
rect 2444 1096 2452 1104
rect 2684 1096 2692 1104
rect 2780 1096 2788 1104
rect 2796 1096 2804 1104
rect 3132 1094 3140 1102
rect 3324 1094 3332 1102
rect 3516 1096 3524 1104
rect 3596 1096 3604 1104
rect 3676 1096 3684 1104
rect 3756 1096 3764 1104
rect 3788 1096 3796 1104
rect 3804 1096 3812 1104
rect 3868 1096 3876 1104
rect 4060 1096 4068 1104
rect 4124 1096 4132 1104
rect 4172 1096 4180 1104
rect 4236 1096 4244 1104
rect 4364 1094 4372 1102
rect 4588 1096 4596 1104
rect 4668 1096 4676 1104
rect 4732 1096 4740 1104
rect 4892 1094 4900 1102
rect 4956 1096 4964 1104
rect 5084 1094 5092 1102
rect 5516 1096 5524 1104
rect 5548 1096 5556 1104
rect 5692 1094 5700 1102
rect 12 1076 20 1084
rect 92 1076 100 1084
rect 124 1076 132 1084
rect 188 1076 196 1084
rect 220 1076 228 1084
rect 332 1076 340 1084
rect 380 1076 388 1084
rect 412 1076 420 1084
rect 604 1076 612 1084
rect 60 1056 68 1064
rect 156 1056 164 1064
rect 332 1056 340 1064
rect 348 1056 356 1064
rect 476 1056 484 1064
rect 540 1056 548 1064
rect 652 1076 660 1084
rect 684 1076 692 1084
rect 812 1076 820 1084
rect 828 1076 836 1084
rect 892 1076 900 1084
rect 1036 1076 1044 1084
rect 1068 1076 1076 1084
rect 1100 1076 1108 1084
rect 1500 1076 1508 1084
rect 1596 1076 1604 1084
rect 1836 1076 1844 1084
rect 1884 1076 1892 1084
rect 1948 1076 1956 1084
rect 2012 1076 2020 1084
rect 2044 1076 2052 1084
rect 2076 1076 2084 1084
rect 2092 1076 2100 1084
rect 2140 1076 2148 1084
rect 2188 1076 2196 1084
rect 2236 1076 2244 1084
rect 2252 1076 2260 1084
rect 2268 1076 2276 1084
rect 2348 1076 2356 1084
rect 2460 1076 2468 1084
rect 2556 1076 2564 1084
rect 2636 1076 2644 1084
rect 2716 1076 2724 1084
rect 2764 1076 2772 1084
rect 2828 1076 2836 1084
rect 2924 1076 2932 1084
rect 2988 1076 2996 1084
rect 3148 1076 3156 1084
rect 3292 1076 3300 1084
rect 3660 1076 3668 1084
rect 3868 1076 3876 1084
rect 3884 1076 3892 1084
rect 3980 1076 3988 1084
rect 4188 1076 4196 1084
rect 4204 1076 4212 1084
rect 4300 1076 4308 1084
rect 4332 1076 4340 1084
rect 4588 1076 4596 1084
rect 4620 1076 4628 1084
rect 4684 1076 4692 1084
rect 4780 1076 4788 1084
rect 4796 1076 4804 1084
rect 5100 1076 5108 1084
rect 5228 1076 5236 1084
rect 5324 1076 5332 1084
rect 5340 1076 5348 1084
rect 5436 1076 5444 1084
rect 5660 1076 5668 1084
rect 652 1056 660 1064
rect 940 1056 948 1064
rect 988 1056 996 1064
rect 1020 1056 1028 1064
rect 1228 1056 1236 1064
rect 1276 1056 1284 1064
rect 1356 1056 1364 1064
rect 1436 1056 1444 1064
rect 1452 1056 1460 1064
rect 1628 1056 1636 1064
rect 1692 1056 1700 1064
rect 2156 1056 2164 1064
rect 2396 1056 2404 1064
rect 2572 1056 2580 1064
rect 2732 1056 2740 1064
rect 3820 1056 3828 1064
rect 3996 1056 4004 1064
rect 4060 1056 4068 1064
rect 124 1036 132 1044
rect 172 1036 180 1044
rect 492 1036 500 1044
rect 556 1036 564 1044
rect 668 1036 676 1044
rect 908 1036 916 1044
rect 1004 1036 1012 1044
rect 1244 1036 1252 1044
rect 1532 1036 1540 1044
rect 1964 1036 1972 1044
rect 2060 1036 2068 1044
rect 2588 1036 2596 1044
rect 2652 1036 2660 1044
rect 3004 1036 3012 1044
rect 3260 1036 3268 1044
rect 3564 1036 3572 1044
rect 3948 1036 3956 1044
rect 4012 1036 4020 1044
rect 4812 1036 4820 1044
rect 5292 1036 5300 1044
rect 5404 1036 5412 1044
rect 2910 1006 2918 1014
rect 2924 1006 2932 1014
rect 2938 1006 2946 1014
rect 28 976 36 984
rect 220 976 228 984
rect 284 976 292 984
rect 876 976 884 984
rect 1052 976 1060 984
rect 1260 976 1268 984
rect 1468 976 1476 984
rect 1756 976 1764 984
rect 2236 976 2244 984
rect 2700 976 2708 984
rect 2876 976 2884 984
rect 3740 976 3748 984
rect 3932 976 3940 984
rect 4076 976 4084 984
rect 4108 976 4116 984
rect 4508 976 4516 984
rect 4620 976 4628 984
rect 4908 976 4916 984
rect 5100 976 5108 984
rect 5116 976 5124 984
rect 5500 976 5508 984
rect 44 956 52 964
rect 268 956 276 964
rect 316 956 324 964
rect 12 936 20 944
rect 140 936 148 944
rect 348 936 356 944
rect 412 936 420 944
rect 492 936 500 944
rect 524 956 532 964
rect 588 956 596 964
rect 604 956 612 964
rect 844 956 852 964
rect 940 956 948 964
rect 1004 956 1012 964
rect 1068 956 1076 964
rect 1148 956 1156 964
rect 1244 956 1252 964
rect 1308 956 1316 964
rect 1804 956 1812 964
rect 636 936 644 944
rect 668 936 676 944
rect 732 936 740 944
rect 780 936 788 944
rect 892 936 900 944
rect 908 936 916 944
rect 972 936 980 944
rect 1100 936 1108 944
rect 1196 936 1204 944
rect 1228 936 1236 944
rect 1452 936 1460 944
rect 1564 936 1572 944
rect 1660 936 1668 944
rect 1868 956 1876 964
rect 1900 956 1908 964
rect 1948 936 1956 944
rect 1964 936 1972 944
rect 2076 936 2084 944
rect 2332 956 2340 964
rect 2428 956 2436 964
rect 2748 956 2756 964
rect 3036 956 3044 964
rect 3564 956 3572 964
rect 3788 956 3796 964
rect 3948 956 3956 964
rect 4780 956 4788 964
rect 4796 956 4804 964
rect 2172 936 2180 944
rect 2204 936 2212 944
rect 2300 936 2308 944
rect 2364 936 2372 944
rect 2412 936 2420 944
rect 2556 936 2564 944
rect 2572 936 2580 944
rect 2668 936 2676 944
rect 2684 936 2692 944
rect 2764 936 2772 944
rect 2860 936 2868 944
rect 2972 936 2980 944
rect 3020 936 3028 944
rect 3068 936 3076 944
rect 3580 936 3588 944
rect 3660 936 3668 944
rect 92 916 100 924
rect 140 916 148 924
rect 204 916 212 924
rect 252 916 260 924
rect 300 916 308 924
rect 364 916 372 924
rect 508 916 516 924
rect 556 916 564 924
rect 620 916 628 924
rect 652 916 660 924
rect 684 916 692 924
rect 732 916 740 924
rect 812 916 820 924
rect 188 896 196 904
rect 396 896 404 904
rect 540 896 548 904
rect 716 896 724 904
rect 764 896 772 904
rect 844 896 852 904
rect 956 916 964 924
rect 1020 916 1028 924
rect 1084 916 1092 924
rect 1212 916 1220 924
rect 1292 916 1300 924
rect 1340 916 1348 924
rect 1452 916 1460 924
rect 1500 916 1508 924
rect 1628 918 1636 926
rect 1692 916 1700 924
rect 1772 916 1780 924
rect 1852 916 1860 924
rect 1868 916 1876 924
rect 1948 916 1956 924
rect 1980 916 1988 924
rect 2028 916 2036 924
rect 2060 916 2068 924
rect 2124 916 2132 924
rect 2188 916 2196 924
rect 2268 916 2276 924
rect 2348 916 2356 924
rect 2412 916 2420 924
rect 2460 916 2468 924
rect 2476 916 2484 924
rect 2492 916 2500 924
rect 2540 916 2548 924
rect 2828 916 2836 924
rect 2956 916 2964 924
rect 3164 918 3172 926
rect 3228 916 3236 924
rect 3356 918 3364 926
rect 3772 936 3780 944
rect 3836 936 3844 944
rect 3900 936 3908 944
rect 3916 936 3924 944
rect 3964 936 3972 944
rect 4028 936 4036 944
rect 4140 936 4148 944
rect 4236 936 4244 944
rect 4268 936 4276 944
rect 4300 936 4308 944
rect 4332 936 4340 944
rect 4524 936 4532 944
rect 4652 936 4660 944
rect 4668 936 4676 944
rect 4764 936 4772 944
rect 4940 936 4948 944
rect 5420 936 5428 944
rect 5516 936 5524 944
rect 5548 936 5556 944
rect 5852 936 5860 944
rect 3420 916 3428 924
rect 3500 916 3508 924
rect 3676 916 3684 924
rect 3820 916 3828 924
rect 3852 916 3860 924
rect 3900 916 3908 924
rect 3980 916 3988 924
rect 4172 916 4180 924
rect 4220 916 4228 924
rect 4284 916 4292 924
rect 4364 918 4372 926
rect 4780 916 4788 924
rect 4828 916 4836 924
rect 4972 918 4980 926
rect 5036 916 5044 924
rect 5180 916 5188 924
rect 5244 918 5252 926
rect 5372 916 5380 924
rect 5580 918 5588 926
rect 5724 916 5732 924
rect 5772 916 5780 924
rect 1404 896 1412 904
rect 1468 896 1476 904
rect 1532 896 1540 904
rect 2012 896 2020 904
rect 2028 896 2036 904
rect 2236 896 2244 904
rect 2252 896 2260 904
rect 2604 896 2612 904
rect 2828 896 2836 904
rect 2924 896 2932 904
rect 3020 896 3028 904
rect 3100 896 3108 904
rect 3884 896 3892 904
rect 4076 896 4084 904
rect 4092 896 4100 904
rect 4188 896 4196 904
rect 4220 896 4228 904
rect 4252 896 4260 904
rect 4908 896 4916 904
rect 108 876 116 884
rect 332 876 340 884
rect 572 876 580 884
rect 748 876 756 884
rect 1148 876 1156 884
rect 2908 876 2916 884
rect 3452 876 3460 884
rect 3484 876 3492 884
rect 3820 876 3828 884
rect 4844 876 4852 884
rect 5484 876 5492 884
rect 5676 876 5684 884
rect 5708 876 5716 884
rect 5756 876 5764 884
rect 476 856 484 864
rect 92 836 100 844
rect 1436 836 1444 844
rect 2060 836 2068 844
rect 2140 836 2148 844
rect 2396 836 2404 844
rect 3084 836 3092 844
rect 3292 836 3300 844
rect 1358 806 1366 814
rect 1372 806 1380 814
rect 1386 806 1394 814
rect 4446 806 4454 814
rect 4460 806 4468 814
rect 4474 806 4482 814
rect 780 776 788 784
rect 1756 776 1764 784
rect 1852 776 1860 784
rect 1900 776 1908 784
rect 1948 776 1956 784
rect 1996 776 2004 784
rect 2220 776 2228 784
rect 2764 776 2772 784
rect 2860 776 2868 784
rect 3612 776 3620 784
rect 3836 776 3844 784
rect 3916 776 3924 784
rect 4284 776 4292 784
rect 4684 776 4692 784
rect 5292 776 5300 784
rect 732 736 740 744
rect 828 736 836 744
rect 2284 736 2292 744
rect 2444 736 2452 744
rect 2876 736 2884 744
rect 5180 736 5188 744
rect 5324 736 5332 744
rect 5596 736 5604 744
rect 5788 736 5796 744
rect 124 716 132 724
rect 220 716 228 724
rect 268 716 276 724
rect 284 716 292 724
rect 316 716 324 724
rect 636 716 644 724
rect 668 716 676 724
rect 972 716 980 724
rect 1020 716 1028 724
rect 1052 716 1060 724
rect 1084 716 1092 724
rect 1260 716 1268 724
rect 188 696 196 704
rect 316 696 324 704
rect 412 696 420 704
rect 444 696 452 704
rect 508 696 516 704
rect 556 696 564 704
rect 620 696 628 704
rect 796 696 804 704
rect 1052 696 1060 704
rect 1100 696 1108 704
rect 1164 696 1172 704
rect 1196 696 1204 704
rect 1228 696 1236 704
rect 1804 716 1812 724
rect 1916 716 1924 724
rect 2028 716 2036 724
rect 2108 716 2116 724
rect 2476 716 2484 724
rect 2540 716 2548 724
rect 2588 716 2596 724
rect 2604 716 2612 724
rect 2716 716 2724 724
rect 2732 716 2740 724
rect 2844 716 2852 724
rect 3852 716 3860 724
rect 1436 696 1444 704
rect 1596 694 1604 702
rect 1660 696 1668 704
rect 1756 696 1764 704
rect 1820 696 1828 704
rect 1836 696 1844 704
rect 1932 696 1940 704
rect 1996 696 2004 704
rect 2124 696 2132 704
rect 2188 696 2196 704
rect 2268 696 2276 704
rect 2412 696 2420 704
rect 2460 696 2468 704
rect 2508 696 2516 704
rect 2684 696 2692 704
rect 2700 696 2708 704
rect 2764 696 2772 704
rect 2828 696 2836 704
rect 2860 696 2868 704
rect 2988 696 2996 704
rect 3020 696 3028 704
rect 3100 696 3108 704
rect 3116 696 3124 704
rect 3228 696 3236 704
rect 3244 696 3252 704
rect 3964 716 3972 724
rect 4060 716 4068 724
rect 4108 716 4116 724
rect 4140 716 4148 724
rect 4268 716 4276 724
rect 4780 716 4788 724
rect 4940 716 4948 724
rect 5244 716 5252 724
rect 3484 694 3492 702
rect 3676 694 3684 702
rect 3996 696 4004 704
rect 4124 696 4132 704
rect 4316 696 4324 704
rect 4380 696 4388 704
rect 4556 696 4564 704
rect 4588 696 4596 704
rect 4748 696 4756 704
rect 4844 696 4852 704
rect 4876 696 4884 704
rect 4908 696 4916 704
rect 4924 696 4932 704
rect 4972 696 4980 704
rect 5036 696 5044 704
rect 5068 696 5076 704
rect 5100 696 5108 704
rect 5180 696 5188 704
rect 5196 696 5204 704
rect 5292 696 5300 704
rect 5356 696 5364 704
rect 5468 694 5476 702
rect 5660 694 5668 702
rect 5804 696 5812 704
rect 12 676 20 684
rect 124 676 132 684
rect 156 676 164 684
rect 172 676 180 684
rect 332 676 340 684
rect 364 676 372 684
rect 428 676 436 684
rect 460 676 468 684
rect 572 676 580 684
rect 380 656 388 664
rect 508 656 516 664
rect 620 676 628 684
rect 748 676 756 684
rect 860 676 868 684
rect 940 676 948 684
rect 988 676 996 684
rect 1036 676 1044 684
rect 764 656 772 664
rect 924 656 932 664
rect 1132 656 1140 664
rect 1180 676 1188 684
rect 1212 676 1220 684
rect 1308 676 1316 684
rect 1340 676 1348 684
rect 1372 676 1380 684
rect 1436 676 1444 684
rect 1532 676 1540 684
rect 1740 676 1748 684
rect 1884 676 1892 684
rect 1980 676 1988 684
rect 2124 676 2132 684
rect 2268 676 2276 684
rect 2396 676 2404 684
rect 2492 676 2500 684
rect 2540 676 2548 684
rect 2556 676 2564 684
rect 2668 676 2676 684
rect 2796 676 2804 684
rect 2828 676 2836 684
rect 2908 676 2916 684
rect 2956 676 2964 684
rect 3036 676 3044 684
rect 3084 676 3092 684
rect 3212 676 3220 684
rect 1804 656 1812 664
rect 1868 656 1876 664
rect 1964 656 1972 664
rect 2060 656 2068 664
rect 2140 656 2148 664
rect 2156 656 2164 664
rect 2204 656 2212 664
rect 2236 656 2244 664
rect 2252 656 2260 664
rect 2364 656 2372 664
rect 2460 656 2468 664
rect 2620 656 2628 664
rect 2636 656 2644 664
rect 2796 656 2804 664
rect 2956 656 2964 664
rect 3068 656 3076 664
rect 3164 656 3172 664
rect 3196 656 3204 664
rect 3276 656 3284 664
rect 3324 676 3332 684
rect 3420 676 3428 684
rect 3452 676 3460 684
rect 3532 676 3540 684
rect 3644 676 3652 684
rect 3724 676 3732 684
rect 3900 676 3908 684
rect 4012 676 4020 684
rect 4124 676 4132 684
rect 4236 676 4244 684
rect 4380 676 4388 684
rect 4476 676 4484 684
rect 4508 676 4516 684
rect 4572 676 4580 684
rect 4604 676 4612 684
rect 4620 676 4628 684
rect 4716 676 4724 684
rect 4732 676 4740 684
rect 4844 676 4852 684
rect 4924 676 4932 684
rect 4988 676 4996 684
rect 5084 676 5092 684
rect 5148 676 5156 684
rect 5196 676 5204 684
rect 5308 676 5316 684
rect 5404 676 5412 684
rect 5500 676 5508 684
rect 5676 676 5684 684
rect 5724 676 5732 684
rect 5852 676 5860 684
rect 4156 656 4164 664
rect 4220 656 4228 664
rect 4268 656 4276 664
rect 4300 656 4308 664
rect 4364 656 4372 664
rect 4780 656 4788 664
rect 4796 656 4804 664
rect 4844 656 4852 664
rect 5004 656 5012 664
rect 5132 656 5140 664
rect 5148 656 5156 664
rect 44 636 52 644
rect 124 636 132 644
rect 268 636 276 644
rect 348 636 356 644
rect 700 636 708 644
rect 780 636 788 644
rect 892 636 900 644
rect 972 636 980 644
rect 1004 636 1012 644
rect 1468 636 1476 644
rect 1724 636 1732 644
rect 2380 636 2388 644
rect 2588 636 2596 644
rect 3052 636 3060 644
rect 3260 636 3268 644
rect 3388 636 3396 644
rect 3804 636 3812 644
rect 4204 636 4212 644
rect 4348 636 4356 644
rect 2910 606 2918 614
rect 2924 606 2932 614
rect 2938 606 2946 614
rect 28 576 36 584
rect 92 576 100 584
rect 860 576 868 584
rect 1212 576 1220 584
rect 1436 576 1444 584
rect 1500 576 1508 584
rect 1964 576 1972 584
rect 2060 576 2068 584
rect 2220 576 2228 584
rect 2268 576 2276 584
rect 2476 576 2484 584
rect 2668 576 2676 584
rect 2796 576 2804 584
rect 2844 576 2852 584
rect 2972 576 2980 584
rect 3244 576 3252 584
rect 3692 576 3700 584
rect 3948 576 3956 584
rect 4156 576 4164 584
rect 4540 576 4548 584
rect 4924 576 4932 584
rect 4988 576 4996 584
rect 5052 576 5060 584
rect 5100 576 5108 584
rect 5196 576 5204 584
rect 5420 576 5428 584
rect 5628 576 5636 584
rect 44 556 52 564
rect 156 556 164 564
rect 332 556 340 564
rect 572 556 580 564
rect 604 556 612 564
rect 620 556 628 564
rect 636 556 644 564
rect 1068 556 1076 564
rect 1164 556 1172 564
rect 1228 556 1236 564
rect 1308 556 1316 564
rect 1324 556 1332 564
rect 1468 556 1476 564
rect 2236 556 2244 564
rect 108 536 116 544
rect 204 536 212 544
rect 236 536 244 544
rect 300 536 308 544
rect 364 536 372 544
rect 412 536 420 544
rect 508 536 516 544
rect 668 536 676 544
rect 796 536 804 544
rect 892 536 900 544
rect 988 536 996 544
rect 1100 536 1108 544
rect 1132 536 1140 544
rect 1260 536 1268 544
rect 1292 536 1300 544
rect 1516 536 1524 544
rect 1532 536 1540 544
rect 1644 536 1652 544
rect 1660 536 1668 544
rect 1756 536 1764 544
rect 1788 536 1796 544
rect 1980 536 1988 544
rect 1996 536 2004 544
rect 2092 536 2100 544
rect 2124 536 2132 544
rect 2156 536 2164 544
rect 2172 536 2180 544
rect 2300 556 2308 564
rect 2828 556 2836 564
rect 2860 556 2868 564
rect 3004 556 3012 564
rect 3116 556 3124 564
rect 3164 556 3172 564
rect 3324 556 3332 564
rect 3900 556 3908 564
rect 4412 556 4420 564
rect 4764 556 4772 564
rect 4780 556 4788 564
rect 4860 556 4868 564
rect 4940 556 4948 564
rect 4972 556 4980 564
rect 5036 556 5044 564
rect 5116 556 5124 564
rect 2348 536 2356 544
rect 2412 536 2420 544
rect 2508 536 2516 544
rect 2556 536 2564 544
rect 2780 536 2788 544
rect 2924 536 2932 544
rect 3036 536 3044 544
rect 3052 536 3060 544
rect 3084 536 3092 544
rect 3148 536 3156 544
rect 3180 536 3188 544
rect 3228 536 3236 544
rect 3260 536 3268 544
rect 3388 536 3396 544
rect 3500 536 3508 544
rect 3532 536 3540 544
rect 3724 536 3732 544
rect 3964 536 3972 544
rect 3996 536 4004 544
rect 4092 536 4100 544
rect 4220 536 4228 544
rect 4332 536 4340 544
rect 4348 536 4356 544
rect 4492 536 4500 544
rect 4588 536 4596 544
rect 4604 536 4612 544
rect 4636 536 4644 544
rect 4700 536 4708 544
rect 4876 536 4884 544
rect 4972 536 4980 544
rect 5004 536 5012 544
rect 5228 536 5236 544
rect 5500 536 5508 544
rect 5596 536 5604 544
rect 5724 536 5732 544
rect 12 516 20 524
rect 188 516 196 524
rect 204 516 212 524
rect 252 516 260 524
rect 284 516 292 524
rect 316 516 324 524
rect 396 516 404 524
rect 428 516 436 524
rect 476 516 484 524
rect 540 516 548 524
rect 684 516 692 524
rect 764 516 772 524
rect 780 516 788 524
rect 812 516 820 524
rect 1020 516 1028 524
rect 1116 516 1124 524
rect 1180 516 1188 524
rect 1276 516 1284 524
rect 1404 516 1412 524
rect 1820 518 1828 526
rect 2332 516 2340 524
rect 2524 516 2532 524
rect 2588 516 2596 524
rect 2636 516 2644 524
rect 2732 516 2740 524
rect 2764 516 2772 524
rect 2780 516 2788 524
rect 2828 516 2836 524
rect 2940 516 2948 524
rect 3052 516 3060 524
rect 3132 516 3140 524
rect 3196 516 3204 524
rect 3212 516 3220 524
rect 3276 516 3284 524
rect 3292 516 3300 524
rect 3324 516 3332 524
rect 3340 516 3348 524
rect 3404 516 3412 524
rect 92 496 100 504
rect 140 496 148 504
rect 236 496 244 504
rect 492 496 500 504
rect 508 496 516 504
rect 844 496 852 504
rect 860 496 868 504
rect 908 496 916 504
rect 956 496 964 504
rect 1052 496 1060 504
rect 1148 496 1156 504
rect 1244 496 1252 504
rect 2108 496 2116 504
rect 2364 496 2372 504
rect 2396 496 2404 504
rect 2972 496 2980 504
rect 3436 496 3444 504
rect 3468 516 3476 524
rect 3484 516 3492 524
rect 3564 518 3572 526
rect 3756 518 3764 526
rect 4028 518 4036 526
rect 4172 516 4180 524
rect 4524 496 4532 504
rect 4572 516 4580 524
rect 4684 516 4692 524
rect 4716 516 4724 524
rect 4812 516 4820 524
rect 4860 516 4868 524
rect 4892 516 4900 524
rect 5020 516 5028 524
rect 5084 516 5092 524
rect 5324 516 5332 524
rect 5356 516 5364 524
rect 5564 518 5572 526
rect 5756 518 5764 526
rect 4636 496 4644 504
rect 4652 496 4660 504
rect 4924 496 4932 504
rect 460 476 468 484
rect 1724 476 1732 484
rect 3084 476 3092 484
rect 3372 476 3380 484
rect 3852 476 3860 484
rect 3884 476 3892 484
rect 2700 456 2708 464
rect 172 436 180 444
rect 444 436 452 444
rect 588 436 596 444
rect 636 436 644 444
rect 732 436 740 444
rect 812 436 820 444
rect 924 436 932 444
rect 1020 436 1028 444
rect 1308 436 1316 444
rect 1580 436 1588 444
rect 1948 436 1956 444
rect 2188 436 2196 444
rect 2620 436 2628 444
rect 2668 436 2676 444
rect 2748 436 2756 444
rect 4364 436 4372 444
rect 4764 436 4772 444
rect 5436 436 5444 444
rect 1358 406 1366 414
rect 1372 406 1380 414
rect 1386 406 1394 414
rect 4446 406 4454 414
rect 4460 406 4468 414
rect 4474 406 4482 414
rect 508 376 516 384
rect 556 376 564 384
rect 876 376 884 384
rect 1932 376 1940 384
rect 2540 376 2548 384
rect 2684 376 2692 384
rect 2876 376 2884 384
rect 3004 376 3012 384
rect 3180 376 3188 384
rect 3212 376 3220 384
rect 3260 376 3268 384
rect 4188 376 4196 384
rect 4716 376 4724 384
rect 4876 376 4884 384
rect 4956 376 4964 384
rect 5100 376 5108 384
rect 5324 376 5332 384
rect 5564 376 5572 384
rect 5692 376 5700 384
rect 2332 356 2340 364
rect 4364 356 4372 364
rect 108 336 116 344
rect 4556 336 4564 344
rect 76 316 84 324
rect 124 316 132 324
rect 204 316 212 324
rect 188 296 196 304
rect 236 296 244 304
rect 300 296 308 304
rect 364 316 372 324
rect 1004 316 1012 324
rect 1564 316 1572 324
rect 1644 316 1652 324
rect 1708 316 1716 324
rect 1788 316 1796 324
rect 396 296 404 304
rect 428 296 436 304
rect 524 296 532 304
rect 764 296 772 304
rect 796 296 804 304
rect 1004 296 1012 304
rect 1036 296 1044 304
rect 1116 294 1124 302
rect 1180 296 1188 304
rect 1676 296 1684 304
rect 1756 296 1764 304
rect 2108 316 2116 324
rect 2188 316 2196 324
rect 2268 316 2276 324
rect 2316 316 2324 324
rect 2572 316 2580 324
rect 2620 316 2628 324
rect 1836 296 1844 304
rect 1980 296 1988 304
rect 2060 296 2068 304
rect 92 276 100 284
rect 172 276 180 284
rect 252 276 260 284
rect 316 276 324 284
rect 412 276 420 284
rect 444 276 452 284
rect 588 276 596 284
rect 684 276 692 284
rect 892 276 900 284
rect 988 276 996 284
rect 1004 276 1012 284
rect 1052 276 1060 284
rect 1084 276 1092 284
rect 1260 276 1268 284
rect 1356 276 1364 284
rect 1420 276 1428 284
rect 1516 276 1524 284
rect 1532 276 1540 284
rect 1612 276 1620 284
rect 1628 276 1636 284
rect 1660 276 1668 284
rect 1740 276 1748 284
rect 1820 276 1828 284
rect 1852 276 1860 284
rect 1868 276 1876 284
rect 1964 276 1972 284
rect 1996 276 2004 284
rect 2044 276 2052 284
rect 2140 276 2148 284
rect 2396 296 2404 304
rect 2204 276 2212 284
rect 2300 276 2308 284
rect 2348 276 2356 284
rect 2476 296 2484 304
rect 2492 296 2500 304
rect 2684 296 2692 304
rect 2732 316 2740 324
rect 2844 316 2852 324
rect 2908 316 2916 324
rect 2956 316 2964 324
rect 3132 316 3140 324
rect 2764 296 2772 304
rect 2860 296 2868 304
rect 2876 296 2884 304
rect 3004 296 3012 304
rect 3084 296 3092 304
rect 3100 296 3108 304
rect 3324 316 3332 324
rect 3180 296 3188 304
rect 3292 296 3300 304
rect 3308 296 3316 304
rect 3340 296 3348 304
rect 3356 296 3364 304
rect 3484 296 3492 304
rect 3532 316 3540 324
rect 3596 316 3604 324
rect 4156 316 4164 324
rect 4220 316 4228 324
rect 4316 316 4324 324
rect 4428 316 4436 324
rect 4524 316 4532 324
rect 4572 316 4580 324
rect 4588 316 4596 324
rect 4620 316 4628 324
rect 4652 316 4660 324
rect 4908 316 4916 324
rect 4924 316 4932 324
rect 4988 316 4996 324
rect 5516 316 5524 324
rect 5548 316 5556 324
rect 5596 316 5604 324
rect 5820 316 5828 324
rect 3564 296 3572 304
rect 3676 296 3684 304
rect 3804 294 3812 302
rect 3852 296 3860 304
rect 3948 296 3956 304
rect 4124 296 4132 304
rect 4188 296 4196 304
rect 4220 296 4228 304
rect 12 256 20 264
rect 140 256 148 264
rect 460 256 468 264
rect 492 256 500 264
rect 2028 256 2036 264
rect 2428 276 2436 284
rect 2460 276 2468 284
rect 2540 276 2548 284
rect 2652 276 2660 284
rect 2668 276 2676 284
rect 2780 276 2788 284
rect 2860 276 2868 284
rect 3020 276 3028 284
rect 3084 276 3092 284
rect 3196 276 3204 284
rect 3372 276 3380 284
rect 3436 276 3444 284
rect 3468 276 3476 284
rect 3548 276 3556 284
rect 3612 276 3620 284
rect 3740 276 3748 284
rect 4108 276 4116 284
rect 4124 276 4132 284
rect 4140 276 4148 284
rect 4172 276 4180 284
rect 4396 296 4404 304
rect 4492 296 4500 304
rect 4620 296 4628 304
rect 4700 296 4708 304
rect 4764 296 4772 304
rect 4780 296 4788 304
rect 4844 296 4852 304
rect 4860 296 4868 304
rect 4956 296 4964 304
rect 5020 296 5028 304
rect 5052 296 5060 304
rect 5148 296 5156 304
rect 5196 296 5204 304
rect 5228 296 5236 304
rect 5276 296 5284 304
rect 5388 296 5396 304
rect 5500 296 5508 304
rect 5628 296 5636 304
rect 5788 296 5796 304
rect 4284 276 4292 284
rect 4332 276 4340 284
rect 4380 276 4388 284
rect 4444 276 4452 284
rect 4684 276 4692 284
rect 4716 276 4724 284
rect 4748 276 4756 284
rect 4796 276 4804 284
rect 4828 276 4836 284
rect 4860 276 4868 284
rect 4972 276 4980 284
rect 5004 276 5012 284
rect 5036 276 5044 284
rect 5068 276 5076 284
rect 5100 276 5108 284
rect 5180 276 5188 284
rect 5292 276 5300 284
rect 5404 276 5412 284
rect 3036 256 3044 264
rect 3228 256 3236 264
rect 3244 256 3252 264
rect 3276 256 3284 264
rect 3420 256 3428 264
rect 3612 256 3620 264
rect 4332 256 4340 264
rect 5148 256 5156 264
rect 5244 256 5252 264
rect 5436 256 5444 264
rect 5484 276 5492 284
rect 5548 276 5556 284
rect 5612 276 5620 284
rect 5644 276 5652 284
rect 5660 276 5668 284
rect 5756 276 5764 284
rect 5772 276 5780 284
rect 5804 276 5812 284
rect 5580 256 5588 264
rect 60 236 68 244
rect 156 236 164 244
rect 204 236 212 244
rect 348 236 356 244
rect 652 236 660 244
rect 1244 236 1252 244
rect 1292 236 1300 244
rect 1484 236 1492 244
rect 1548 236 1556 244
rect 1596 236 1604 244
rect 2012 236 2020 244
rect 2092 236 2100 244
rect 2108 236 2116 244
rect 2172 236 2180 244
rect 2444 236 2452 244
rect 2572 236 2580 244
rect 3052 236 3060 244
rect 3452 236 3460 244
rect 3932 236 3940 244
rect 4252 236 4260 244
rect 4812 236 4820 244
rect 5468 236 5476 244
rect 2910 206 2918 214
rect 2924 206 2932 214
rect 2938 206 2946 214
rect 572 176 580 184
rect 764 176 772 184
rect 956 176 964 184
rect 1148 176 1156 184
rect 1340 176 1348 184
rect 1564 176 1572 184
rect 1884 176 1892 184
rect 2204 176 2212 184
rect 2460 176 2468 184
rect 2812 176 2820 184
rect 2892 176 2900 184
rect 3148 176 3156 184
rect 3564 176 3572 184
rect 3756 176 3764 184
rect 4092 176 4100 184
rect 4236 176 4244 184
rect 4380 176 4388 184
rect 4524 176 4532 184
rect 4556 176 4564 184
rect 4604 176 4612 184
rect 5052 176 5060 184
rect 5132 176 5140 184
rect 5164 176 5172 184
rect 5420 176 5428 184
rect 5516 176 5524 184
rect 5596 176 5604 184
rect 5772 176 5780 184
rect 12 156 20 164
rect 1596 156 1604 164
rect 1612 156 1620 164
rect 1644 156 1652 164
rect 1676 156 1684 164
rect 28 136 36 144
rect 156 136 164 144
rect 172 136 180 144
rect 268 136 276 144
rect 284 136 292 144
rect 380 136 388 144
rect 604 136 612 144
rect 796 136 804 144
rect 988 136 996 144
rect 1180 136 1188 144
rect 1404 136 1412 144
rect 1500 136 1508 144
rect 1516 136 1524 144
rect 1708 156 1716 164
rect 2124 156 2132 164
rect 2188 156 2196 164
rect 2316 156 2324 164
rect 3100 156 3108 164
rect 3228 156 3236 164
rect 4140 156 4148 164
rect 4156 156 4164 164
rect 4412 156 4420 164
rect 4620 156 4628 164
rect 4684 156 4692 164
rect 5004 156 5012 164
rect 5068 156 5076 164
rect 5100 156 5108 164
rect 5212 156 5220 164
rect 5356 156 5364 164
rect 5436 156 5444 164
rect 5532 156 5540 164
rect 1724 136 1732 144
rect 1820 136 1828 144
rect 1916 136 1924 144
rect 1932 136 1940 144
rect 1996 136 2004 144
rect 2236 136 2244 144
rect 76 116 84 124
rect 124 116 132 124
rect 140 116 148 124
rect 444 118 452 126
rect 508 116 516 124
rect 636 118 644 126
rect 700 116 708 124
rect 828 118 836 126
rect 892 116 900 124
rect 1020 118 1028 126
rect 1084 116 1092 124
rect 1228 116 1236 124
rect 1740 116 1748 124
rect 1756 116 1764 124
rect 1948 116 1956 124
rect 92 96 100 104
rect 108 96 116 104
rect 1980 96 1988 104
rect 2092 116 2100 124
rect 2236 116 2244 124
rect 2316 136 2324 144
rect 2332 136 2340 144
rect 2428 136 2436 144
rect 2476 136 2484 144
rect 2492 136 2500 144
rect 2540 136 2548 144
rect 2604 136 2612 144
rect 2652 136 2660 144
rect 2748 136 2756 144
rect 2764 136 2772 144
rect 2828 136 2836 144
rect 2972 136 2980 144
rect 2988 136 2996 144
rect 3084 136 3092 144
rect 3164 136 3172 144
rect 3276 136 3284 144
rect 3372 136 3380 144
rect 3852 136 3860 144
rect 4012 136 4020 144
rect 4028 136 4036 144
rect 4124 136 4132 144
rect 4172 136 4180 144
rect 4284 136 4292 144
rect 4300 136 4308 144
rect 4460 136 4468 144
rect 4476 136 4484 144
rect 4572 136 4580 144
rect 4636 136 4644 144
rect 4700 136 4708 144
rect 2476 116 2484 124
rect 2556 116 2564 124
rect 2780 116 2788 124
rect 2060 96 2068 104
rect 2204 96 2212 104
rect 2444 96 2452 104
rect 2524 96 2532 104
rect 2636 96 2644 104
rect 2812 96 2820 104
rect 3020 96 3028 104
rect 3052 116 3060 124
rect 3068 116 3076 124
rect 3196 116 3204 124
rect 3244 116 3252 124
rect 3260 116 3268 124
rect 3372 116 3380 124
rect 3436 118 3444 126
rect 3500 116 3508 124
rect 3628 118 3636 126
rect 3692 116 3700 124
rect 3820 118 3828 126
rect 3964 116 3972 124
rect 4188 116 4196 124
rect 4220 96 4228 104
rect 4268 116 4276 124
rect 4348 116 4356 124
rect 4812 136 4820 144
rect 4892 136 4900 144
rect 4924 136 4932 144
rect 4940 136 4948 144
rect 5020 136 5028 144
rect 5116 136 5124 144
rect 5260 136 5268 144
rect 5292 136 5300 144
rect 5340 136 5348 144
rect 5404 136 5412 144
rect 5452 136 5460 144
rect 5468 136 5476 144
rect 5548 136 5556 144
rect 5612 136 5620 144
rect 5708 136 5716 144
rect 5724 136 5732 144
rect 4652 116 4660 124
rect 4796 116 4804 124
rect 4332 96 4340 104
rect 4524 96 4532 104
rect 4684 96 4692 104
rect 4764 96 4772 104
rect 4860 96 4868 104
rect 4908 116 4916 124
rect 4956 116 4964 124
rect 5100 116 5108 124
rect 5196 116 5204 124
rect 5244 116 5252 124
rect 5276 116 5284 124
rect 5356 116 5364 124
rect 5388 116 5396 124
rect 5484 116 5492 124
rect 5500 116 5508 124
rect 5564 116 5572 124
rect 5644 116 5652 124
rect 5740 116 5748 124
rect 5788 116 5796 124
rect 4956 96 4964 104
rect 4988 96 4996 104
rect 5772 96 5780 104
rect 60 76 68 84
rect 236 76 244 84
rect 348 76 356 84
rect 2268 76 2276 84
rect 2556 76 2564 84
rect 2716 76 2724 84
rect 3948 76 3956 84
rect 4300 76 4308 84
rect 5852 76 5860 84
rect 76 56 84 64
rect 2012 56 2020 64
rect 2396 56 2404 64
rect 1358 6 1366 14
rect 1372 6 1380 14
rect 1386 6 1394 14
rect 4446 6 4454 14
rect 4460 6 4468 14
rect 4474 6 4482 14
<< metal2 >>
rect 973 4204 979 4243
rect 2904 4206 2910 4214
rect 2918 4206 2924 4214
rect 2932 4206 2938 4214
rect 2946 4206 2952 4214
rect 397 4164 403 4176
rect 109 4144 115 4156
rect 285 4144 291 4156
rect 93 4124 99 4136
rect 29 3944 35 4116
rect 205 4104 211 4116
rect 77 3964 83 4036
rect 29 3904 35 3936
rect 109 3884 115 3916
rect 13 3744 19 3876
rect 61 3744 67 3836
rect 13 3524 19 3676
rect 29 3383 35 3736
rect 61 3704 67 3716
rect 52 3517 67 3523
rect 61 3504 67 3517
rect 61 3464 67 3476
rect 77 3464 83 3876
rect 125 3744 131 3916
rect 157 3904 163 4036
rect 221 3984 227 4076
rect 237 3883 243 4116
rect 269 4044 275 4136
rect 349 4124 355 4156
rect 461 4143 467 4176
rect 973 4144 979 4196
rect 2205 4164 2211 4176
rect 452 4137 467 4143
rect 381 4064 387 4096
rect 429 4084 435 4116
rect 781 4104 787 4118
rect 381 3944 387 4036
rect 228 3877 243 3883
rect 157 3844 163 3876
rect 157 3764 163 3836
rect 93 3624 99 3716
rect 157 3544 163 3756
rect 189 3644 195 3756
rect 205 3704 211 3876
rect 237 3724 243 3836
rect 253 3744 259 3916
rect 333 3884 339 3936
rect 381 3924 387 3936
rect 397 3897 412 3903
rect 333 3784 339 3856
rect 349 3784 355 3836
rect 317 3744 323 3756
rect 365 3744 371 3756
rect 221 3664 227 3716
rect 205 3584 211 3616
rect 173 3484 179 3496
rect 189 3484 195 3536
rect 221 3484 227 3636
rect 253 3604 259 3716
rect 269 3624 275 3696
rect 301 3644 307 3736
rect 189 3464 195 3476
rect 13 3377 35 3383
rect 13 3344 19 3377
rect 109 3344 115 3356
rect 13 3124 19 3136
rect 45 3084 51 3096
rect 13 2964 19 3036
rect 61 2984 67 3236
rect 77 3084 83 3236
rect 125 3104 131 3436
rect 189 3344 195 3416
rect 189 3144 195 3336
rect 205 3144 211 3436
rect 221 3384 227 3456
rect 253 3364 259 3436
rect 269 3244 275 3356
rect 317 3344 323 3716
rect 349 3704 355 3716
rect 349 3584 355 3616
rect 365 3464 371 3696
rect 381 3664 387 3716
rect 381 3503 387 3656
rect 397 3624 403 3897
rect 429 3884 435 3956
rect 477 3884 483 3896
rect 493 3884 499 3976
rect 525 3904 531 3916
rect 541 3904 547 3956
rect 573 3864 579 4076
rect 621 3904 627 4056
rect 621 3884 627 3896
rect 637 3884 643 3896
rect 765 3864 771 3936
rect 797 3884 803 3916
rect 413 3784 419 3856
rect 429 3684 435 3696
rect 429 3544 435 3676
rect 381 3497 403 3503
rect 365 3444 371 3456
rect 285 3244 291 3296
rect 221 3124 227 3236
rect 285 3104 291 3236
rect 301 3124 307 3316
rect 317 3124 323 3136
rect 109 3084 115 3096
rect 13 2664 19 2956
rect 109 2864 115 3076
rect 157 3064 163 3096
rect 125 2964 131 3056
rect 141 2964 147 3036
rect 125 2944 131 2956
rect 125 2864 131 2916
rect 45 2684 51 2836
rect 61 2644 67 2696
rect 77 2684 83 2856
rect 141 2724 147 2956
rect 205 2944 211 2956
rect 221 2924 227 2996
rect 269 2963 275 3076
rect 285 3064 291 3096
rect 333 3084 339 3236
rect 349 3084 355 3436
rect 381 3404 387 3476
rect 397 3343 403 3497
rect 445 3464 451 3836
rect 461 3704 467 3716
rect 477 3624 483 3736
rect 493 3543 499 3636
rect 477 3537 499 3543
rect 477 3504 483 3537
rect 429 3444 435 3456
rect 388 3337 403 3343
rect 445 3324 451 3436
rect 477 3324 483 3456
rect 493 3344 499 3516
rect 525 3444 531 3496
rect 541 3484 547 3616
rect 605 3604 611 3836
rect 573 3504 579 3596
rect 637 3484 643 3536
rect 653 3504 659 3516
rect 541 3404 547 3476
rect 589 3364 595 3396
rect 605 3364 611 3456
rect 685 3444 691 3496
rect 365 3304 371 3316
rect 445 3304 451 3316
rect 541 3304 547 3316
rect 413 3244 419 3256
rect 413 3144 419 3236
rect 445 3124 451 3136
rect 500 3117 515 3123
rect 509 3104 515 3117
rect 269 2957 284 2963
rect 157 2844 163 2876
rect 173 2704 179 2836
rect 189 2784 195 2896
rect 189 2744 195 2776
rect 221 2724 227 2736
rect 29 2524 35 2636
rect 61 2504 67 2616
rect 109 2544 115 2576
rect 125 2544 131 2636
rect 189 2624 195 2656
rect 93 1904 99 2436
rect 141 2302 147 2596
rect 205 2584 211 2696
rect 221 2564 227 2636
rect 237 2564 243 2716
rect 189 2524 195 2556
rect 205 2284 211 2536
rect 253 2524 259 2936
rect 269 2724 275 2957
rect 301 2924 307 3076
rect 349 3064 355 3076
rect 333 3024 339 3036
rect 365 2984 371 3096
rect 285 2744 291 2916
rect 317 2903 323 2976
rect 349 2944 355 2956
rect 365 2944 371 2956
rect 333 2904 339 2916
rect 308 2897 323 2903
rect 301 2784 307 2876
rect 333 2684 339 2896
rect 349 2704 355 2796
rect 365 2724 371 2836
rect 381 2664 387 3036
rect 397 2944 403 2956
rect 413 2924 419 2976
rect 445 2944 451 3016
rect 461 2984 467 2996
rect 477 2944 483 2996
rect 509 2984 515 3076
rect 509 2944 515 2956
rect 429 2704 435 2736
rect 445 2683 451 2936
rect 525 2924 531 3176
rect 541 3144 547 3236
rect 605 3143 611 3356
rect 701 3324 707 3836
rect 733 3744 739 3756
rect 733 3684 739 3736
rect 765 3724 771 3736
rect 733 3464 739 3676
rect 765 3664 771 3716
rect 749 3644 755 3656
rect 749 3504 755 3636
rect 765 3504 771 3656
rect 781 3484 787 3496
rect 765 3464 771 3476
rect 749 3404 755 3436
rect 797 3424 803 3876
rect 845 3744 851 4136
rect 989 4064 995 4136
rect 1101 4124 1107 4136
rect 893 3904 899 3916
rect 925 3904 931 3916
rect 989 3884 995 4056
rect 1005 3944 1011 4036
rect 1037 3884 1043 4036
rect 845 3724 851 3736
rect 941 3724 947 3836
rect 1101 3764 1107 4116
rect 1165 4084 1171 4118
rect 1197 3904 1203 4136
rect 1261 4084 1267 4096
rect 1325 3984 1331 4136
rect 1389 4104 1395 4156
rect 1501 4144 1507 4156
rect 1741 4144 1747 4156
rect 1981 4144 1987 4156
rect 1421 4104 1427 4116
rect 1352 4006 1358 4014
rect 1366 4006 1372 4014
rect 1380 4006 1386 4014
rect 1394 4006 1400 4014
rect 1453 3964 1459 4096
rect 1485 3944 1491 4136
rect 1597 4044 1603 4136
rect 1613 3984 1619 4136
rect 1661 4044 1667 4096
rect 1405 3904 1411 3936
rect 1581 3884 1587 3916
rect 1597 3884 1603 3936
rect 1629 3904 1635 4036
rect 1709 3944 1715 4136
rect 1725 4084 1731 4116
rect 1773 4104 1779 4116
rect 1789 4104 1795 4116
rect 1821 4104 1827 4136
rect 1757 4004 1763 4096
rect 1869 4024 1875 4116
rect 1917 4084 1923 4136
rect 2109 4124 2115 4156
rect 2173 4144 2179 4156
rect 1933 4044 1939 4116
rect 1997 4104 2003 4116
rect 1885 3984 1891 4036
rect 2093 4024 2099 4036
rect 1741 3957 1788 3963
rect 1645 3937 1683 3943
rect 1645 3924 1651 3937
rect 1661 3904 1667 3916
rect 1677 3904 1683 3937
rect 1741 3923 1747 3957
rect 1732 3917 1747 3923
rect 1613 3884 1619 3896
rect 1117 3864 1123 3876
rect 1277 3724 1283 3816
rect 1293 3764 1299 3876
rect 1373 3864 1379 3876
rect 1293 3744 1299 3756
rect 1469 3724 1475 3876
rect 1485 3844 1491 3876
rect 1629 3864 1635 3876
rect 1693 3864 1699 3896
rect 1709 3884 1715 3916
rect 1757 3884 1763 3936
rect 1773 3884 1779 3916
rect 1789 3884 1795 3896
rect 1517 3804 1523 3836
rect 1101 3704 1107 3718
rect 861 3517 876 3523
rect 813 3384 819 3436
rect 829 3384 835 3456
rect 717 3324 723 3356
rect 781 3324 787 3376
rect 813 3344 819 3356
rect 669 3264 675 3296
rect 717 3264 723 3296
rect 605 3137 627 3143
rect 621 3084 627 3137
rect 637 3124 643 3136
rect 557 2943 563 3036
rect 621 2964 627 3076
rect 669 2984 675 3136
rect 685 3084 691 3156
rect 733 3144 739 3296
rect 749 3184 755 3196
rect 717 3104 723 3116
rect 733 3097 764 3103
rect 733 3083 739 3097
rect 708 3077 739 3083
rect 685 3024 691 3056
rect 637 2944 643 2976
rect 541 2937 563 2943
rect 493 2884 499 2916
rect 525 2904 531 2916
rect 477 2704 483 2756
rect 525 2684 531 2736
rect 445 2677 460 2683
rect 269 2524 275 2556
rect 317 2524 323 2636
rect 333 2564 339 2636
rect 397 2563 403 2636
rect 413 2584 419 2656
rect 461 2644 467 2656
rect 381 2557 403 2563
rect 333 2524 339 2556
rect 381 2524 387 2557
rect 461 2544 467 2636
rect 477 2584 483 2656
rect 493 2564 499 2636
rect 509 2564 515 2636
rect 541 2604 547 2937
rect 621 2924 627 2936
rect 557 2904 563 2916
rect 557 2764 563 2896
rect 573 2784 579 2916
rect 557 2664 563 2696
rect 589 2684 595 2756
rect 653 2704 659 2836
rect 685 2724 691 2936
rect 701 2864 707 2896
rect 701 2804 707 2856
rect 685 2704 691 2716
rect 717 2704 723 3036
rect 765 2984 771 3076
rect 781 2984 787 3236
rect 797 3204 803 3336
rect 845 3324 851 3456
rect 861 3304 867 3517
rect 877 3504 883 3516
rect 893 3484 899 3516
rect 1005 3504 1011 3676
rect 1165 3504 1171 3656
rect 1309 3524 1315 3636
rect 1352 3606 1358 3614
rect 1366 3606 1372 3614
rect 1380 3606 1386 3614
rect 1394 3606 1400 3614
rect 1501 3544 1507 3736
rect 1533 3726 1539 3776
rect 1757 3764 1763 3876
rect 1805 3764 1811 3976
rect 1837 3924 1843 3956
rect 1597 3604 1603 3736
rect 1789 3724 1795 3756
rect 1853 3724 1859 3956
rect 1997 3904 2003 3976
rect 1869 3864 1875 3896
rect 1885 3884 1891 3896
rect 1965 3884 1971 3896
rect 2029 3884 2035 3916
rect 1901 3864 1907 3876
rect 1965 3864 1971 3876
rect 1725 3684 1731 3716
rect 1773 3644 1779 3716
rect 1869 3704 1875 3856
rect 1917 3783 1923 3836
rect 1901 3777 1923 3783
rect 1901 3703 1907 3777
rect 1949 3744 1955 3756
rect 1965 3744 1971 3856
rect 1981 3784 1987 3876
rect 1924 3737 1939 3743
rect 1901 3697 1916 3703
rect 1933 3684 1939 3737
rect 1997 3704 2003 3716
rect 1901 3644 1907 3676
rect 2013 3644 2019 3876
rect 2045 3864 2051 3916
rect 2077 3764 2083 3896
rect 2045 3704 2051 3756
rect 2093 3724 2099 3896
rect 2109 3764 2115 4116
rect 2285 4104 2291 4116
rect 2189 4044 2195 4096
rect 2141 3824 2147 3936
rect 2157 3904 2163 3976
rect 2189 3923 2195 4036
rect 2205 3944 2211 4036
rect 2269 3984 2275 4036
rect 2189 3917 2204 3923
rect 2125 3704 2131 3736
rect 2157 3684 2163 3896
rect 2189 3724 2195 3856
rect 2205 3744 2211 3876
rect 2253 3863 2259 3916
rect 2285 3904 2291 4096
rect 2333 3904 2339 3996
rect 2404 3917 2419 3923
rect 2381 3884 2387 3896
rect 2253 3857 2300 3863
rect 2301 3744 2307 3756
rect 2397 3744 2403 3756
rect 2173 3704 2179 3716
rect 893 3364 899 3436
rect 941 3324 947 3436
rect 1021 3384 1027 3476
rect 1069 3464 1075 3494
rect 1133 3403 1139 3436
rect 1165 3424 1171 3476
rect 1181 3444 1187 3516
rect 1213 3484 1219 3496
rect 1309 3484 1315 3516
rect 1325 3484 1331 3496
rect 1117 3397 1139 3403
rect 1021 3364 1027 3376
rect 957 3344 963 3356
rect 1021 3344 1027 3356
rect 1085 3344 1091 3376
rect 893 3304 899 3316
rect 813 3063 819 3256
rect 845 3084 851 3096
rect 861 3084 867 3296
rect 829 3064 835 3076
rect 797 3057 819 3063
rect 733 2944 739 2976
rect 749 2924 755 2956
rect 765 2924 771 2956
rect 781 2924 787 2956
rect 797 2944 803 3057
rect 749 2904 755 2916
rect 813 2884 819 3036
rect 829 2884 835 2996
rect 845 2944 851 3056
rect 893 2944 899 3296
rect 909 3164 915 3316
rect 973 3304 979 3336
rect 973 3084 979 3296
rect 1005 3123 1011 3236
rect 996 3117 1011 3123
rect 909 3077 924 3083
rect 909 3024 915 3077
rect 1021 3064 1027 3316
rect 909 2984 915 3016
rect 925 2944 931 3056
rect 989 2984 995 3036
rect 1037 2984 1043 3076
rect 1053 3064 1059 3076
rect 1021 2963 1027 2976
rect 1085 2963 1091 3076
rect 1101 2984 1107 3116
rect 1117 3104 1123 3397
rect 1165 3364 1171 3416
rect 1181 3364 1187 3436
rect 1181 3344 1187 3356
rect 1197 3324 1203 3416
rect 1229 3324 1235 3436
rect 1133 3084 1139 3296
rect 1229 3124 1235 3196
rect 1245 3124 1251 3376
rect 1277 3164 1283 3436
rect 1309 3344 1315 3476
rect 1373 3464 1379 3516
rect 1597 3504 1603 3536
rect 1661 3502 1667 3576
rect 1789 3504 1795 3536
rect 1853 3502 1859 3556
rect 1901 3543 1907 3636
rect 1901 3537 1923 3543
rect 1917 3504 1923 3537
rect 1517 3443 1523 3476
rect 1725 3444 1731 3476
rect 1517 3437 1532 3443
rect 1405 3384 1411 3436
rect 1517 3424 1523 3437
rect 1533 3404 1539 3436
rect 1549 3344 1555 3436
rect 1629 3364 1635 3376
rect 1725 3344 1731 3376
rect 1741 3344 1747 3396
rect 1837 3344 1843 3476
rect 1949 3464 1955 3596
rect 2013 3544 2019 3636
rect 2077 3484 2083 3516
rect 2141 3484 2147 3496
rect 1949 3444 1955 3456
rect 2061 3384 2067 3476
rect 2093 3464 2099 3476
rect 2157 3464 2163 3536
rect 2205 3483 2211 3736
rect 2237 3664 2243 3736
rect 2253 3684 2259 3696
rect 2237 3584 2243 3656
rect 2397 3524 2403 3696
rect 2413 3684 2419 3917
rect 2429 3884 2435 3936
rect 2445 3864 2451 4136
rect 2557 4126 2563 4156
rect 3149 4144 3155 4176
rect 3725 4144 3731 4156
rect 3757 4144 3763 4243
rect 3933 4184 3939 4243
rect 2493 4104 2499 4116
rect 2557 4024 2563 4118
rect 2669 4044 2675 4136
rect 2676 4037 2691 4043
rect 2477 3884 2483 3936
rect 2541 3924 2547 4016
rect 2493 3844 2499 3896
rect 2541 3864 2547 3896
rect 2557 3864 2563 3876
rect 2461 3784 2467 3816
rect 2525 3784 2531 3836
rect 2541 3824 2547 3856
rect 2589 3804 2595 3836
rect 2621 3784 2627 3796
rect 2429 3764 2435 3776
rect 2525 3724 2531 3776
rect 2557 3724 2563 3756
rect 2573 3724 2579 3736
rect 2445 3584 2451 3616
rect 2493 3584 2499 3716
rect 2557 3704 2563 3716
rect 2621 3704 2627 3716
rect 2637 3684 2643 3696
rect 2509 3584 2515 3676
rect 2653 3663 2659 3876
rect 2669 3804 2675 3916
rect 2685 3744 2691 4037
rect 2701 3904 2707 4136
rect 3229 4124 3235 4136
rect 2733 3984 2739 4116
rect 2749 3904 2755 4116
rect 2765 3924 2771 4096
rect 2909 4004 2915 4118
rect 3405 4123 3411 4136
rect 3396 4117 3411 4123
rect 3005 3984 3011 4076
rect 3172 4037 3187 4043
rect 3053 3984 3059 3996
rect 2701 3884 2707 3896
rect 2717 3784 2723 3856
rect 2701 3764 2707 3776
rect 2733 3744 2739 3836
rect 2765 3784 2771 3876
rect 2781 3764 2787 3976
rect 2749 3724 2755 3756
rect 2781 3704 2787 3756
rect 2797 3744 2803 3916
rect 2813 3904 2819 3916
rect 3117 3904 3123 3916
rect 3165 3904 3171 3976
rect 2925 3884 2931 3896
rect 2637 3657 2659 3663
rect 2317 3484 2323 3496
rect 2445 3484 2451 3576
rect 2196 3477 2211 3483
rect 2189 3464 2195 3476
rect 2317 3464 2323 3476
rect 2317 3443 2323 3456
rect 2301 3437 2323 3443
rect 2189 3344 2195 3376
rect 2301 3344 2307 3437
rect 2413 3384 2419 3436
rect 2397 3344 2403 3356
rect 1373 3324 1379 3336
rect 1549 3324 1555 3336
rect 1981 3324 1987 3336
rect 1309 3304 1315 3316
rect 1309 3204 1315 3296
rect 1352 3206 1358 3214
rect 1366 3206 1372 3214
rect 1380 3206 1386 3214
rect 1394 3206 1400 3214
rect 1149 3004 1155 3036
rect 1133 2964 1139 2976
rect 1021 2957 1043 2963
rect 861 2924 867 2936
rect 877 2924 883 2936
rect 765 2704 771 2876
rect 797 2724 803 2776
rect 717 2524 723 2696
rect 733 2544 739 2636
rect 765 2584 771 2676
rect 781 2564 787 2576
rect 349 2504 355 2516
rect 461 2504 467 2516
rect 301 2284 307 2436
rect 317 2284 323 2496
rect 381 2304 387 2436
rect 413 2284 419 2296
rect 125 2144 131 2276
rect 125 2124 131 2136
rect 125 1904 131 2116
rect 13 1484 19 1636
rect 29 1504 35 1836
rect 125 1744 131 1896
rect 189 1864 195 2036
rect 253 1902 259 2236
rect 349 2164 355 2236
rect 269 2124 275 2156
rect 317 2124 323 2136
rect 317 1904 323 2116
rect 381 1864 387 2036
rect 429 1944 435 2236
rect 541 2224 547 2436
rect 557 2302 563 2336
rect 669 2302 675 2436
rect 797 2324 803 2636
rect 813 2524 819 2836
rect 829 2664 835 2696
rect 861 2684 867 2916
rect 957 2764 963 2916
rect 957 2684 963 2756
rect 925 2624 931 2636
rect 909 2564 915 2576
rect 829 2524 835 2536
rect 925 2503 931 2616
rect 1021 2604 1027 2656
rect 973 2524 979 2536
rect 1037 2524 1043 2957
rect 1069 2957 1091 2963
rect 1069 2944 1075 2957
rect 1053 2683 1059 2936
rect 1085 2924 1091 2936
rect 1069 2704 1075 2916
rect 1133 2904 1139 2936
rect 1165 2884 1171 3056
rect 1181 3044 1187 3076
rect 1245 3064 1251 3116
rect 1309 3084 1315 3196
rect 1373 3124 1379 3136
rect 1581 3123 1587 3316
rect 1677 3124 1683 3316
rect 1565 3117 1587 3123
rect 1437 3104 1443 3116
rect 1501 3104 1507 3116
rect 1341 3064 1347 3096
rect 1517 3084 1523 3116
rect 1197 2944 1203 2956
rect 1213 2924 1219 3036
rect 1261 2924 1267 3036
rect 1277 2944 1283 3036
rect 1293 3024 1299 3036
rect 1229 2844 1235 2896
rect 1293 2864 1299 2936
rect 1325 2904 1331 2956
rect 1373 2924 1379 2976
rect 1053 2677 1075 2683
rect 1069 2664 1075 2677
rect 1053 2544 1059 2656
rect 925 2497 940 2503
rect 909 2284 915 2476
rect 973 2283 979 2436
rect 964 2277 979 2283
rect 525 2126 531 2196
rect 557 2144 563 2256
rect 653 2124 659 2216
rect 701 2144 707 2276
rect 925 2203 931 2236
rect 973 2224 979 2236
rect 909 2197 931 2203
rect 701 2124 707 2136
rect 909 2126 915 2197
rect 788 2037 803 2043
rect 397 1904 403 1916
rect 429 1884 435 1916
rect 445 1884 451 2036
rect 765 1964 771 2036
rect 445 1864 451 1876
rect 461 1864 467 1876
rect 141 1726 147 1756
rect 237 1724 243 1776
rect 253 1764 259 1856
rect 205 1584 211 1696
rect 189 1524 195 1576
rect 221 1544 227 1716
rect 13 1364 19 1476
rect 29 1463 35 1496
rect 77 1464 83 1496
rect 29 1457 51 1463
rect 13 1104 19 1276
rect 29 1104 35 1457
rect 45 1344 51 1457
rect 61 1457 76 1463
rect 61 1444 67 1457
rect 93 1344 99 1476
rect 45 1324 51 1336
rect 109 1324 115 1496
rect 148 1477 163 1483
rect 141 1304 147 1376
rect 157 1364 163 1477
rect 205 1464 211 1496
rect 237 1484 243 1556
rect 253 1504 259 1756
rect 269 1744 275 1836
rect 397 1784 403 1836
rect 300 1750 308 1756
rect 269 1564 275 1736
rect 381 1724 387 1736
rect 509 1723 515 1856
rect 525 1764 531 1836
rect 541 1744 547 1896
rect 605 1864 611 1916
rect 653 1904 659 1916
rect 685 1904 691 1916
rect 573 1724 579 1836
rect 509 1717 524 1723
rect 333 1684 339 1716
rect 333 1584 339 1676
rect 413 1584 419 1716
rect 317 1504 323 1516
rect 333 1504 339 1516
rect 365 1504 371 1516
rect 477 1504 483 1716
rect 589 1704 595 1736
rect 605 1724 611 1756
rect 621 1704 627 1836
rect 669 1744 675 1896
rect 701 1744 707 1876
rect 717 1764 723 1876
rect 733 1864 739 1880
rect 749 1744 755 1856
rect 749 1724 755 1736
rect 765 1724 771 1836
rect 493 1684 499 1696
rect 493 1524 499 1536
rect 557 1524 563 1636
rect 637 1544 643 1716
rect 749 1524 755 1536
rect 500 1517 515 1523
rect 13 1084 19 1096
rect 29 1084 35 1096
rect 29 1043 35 1076
rect 13 1037 35 1043
rect 13 944 19 1037
rect 29 984 35 1016
rect 45 964 51 1236
rect 109 1124 115 1236
rect 125 1084 131 1156
rect 141 1104 147 1256
rect 189 1084 195 1436
rect 205 1324 211 1456
rect 221 1264 227 1436
rect 237 1364 243 1476
rect 253 1424 259 1496
rect 317 1484 323 1496
rect 269 1384 275 1456
rect 301 1384 307 1476
rect 381 1464 387 1476
rect 397 1464 403 1476
rect 413 1444 419 1496
rect 461 1464 467 1476
rect 333 1404 339 1436
rect 301 1364 307 1376
rect 349 1364 355 1416
rect 445 1384 451 1436
rect 285 1344 291 1356
rect 253 1284 259 1316
rect 301 1304 307 1316
rect 221 1104 227 1236
rect 333 1104 339 1356
rect 381 1344 387 1356
rect 445 1324 451 1376
rect 365 1104 371 1116
rect 93 1024 99 1076
rect 13 684 19 936
rect 93 863 99 916
rect 109 884 115 916
rect 93 857 115 863
rect 93 764 99 836
rect 76 664 84 670
rect 45 564 51 636
rect 93 584 99 596
rect 109 584 115 857
rect 125 744 131 1036
rect 141 944 147 996
rect 148 937 163 943
rect 141 804 147 916
rect 141 704 147 796
rect 157 724 163 937
rect 173 824 179 1036
rect 189 904 195 1016
rect 221 984 227 1016
rect 285 984 291 1036
rect 317 964 323 1096
rect 381 1084 387 1096
rect 413 1084 419 1136
rect 461 1124 467 1456
rect 477 1344 483 1416
rect 493 1384 499 1496
rect 509 1484 515 1517
rect 653 1517 668 1523
rect 541 1483 547 1516
rect 557 1504 563 1516
rect 605 1504 611 1516
rect 541 1477 556 1483
rect 557 1444 563 1476
rect 621 1464 627 1476
rect 525 1304 531 1336
rect 541 1304 547 1436
rect 589 1344 595 1456
rect 653 1444 659 1517
rect 797 1504 803 2037
rect 877 1924 883 1956
rect 1037 1924 1043 2216
rect 1069 2144 1075 2276
rect 877 1864 883 1916
rect 925 1864 931 1876
rect 941 1864 947 1896
rect 1037 1884 1043 1916
rect 813 1723 819 1836
rect 1021 1784 1027 1836
rect 829 1744 835 1756
rect 925 1744 931 1776
rect 1069 1744 1075 2136
rect 1085 1884 1091 2796
rect 1117 2704 1123 2836
rect 1245 2704 1251 2736
rect 1277 2724 1283 2756
rect 1101 2684 1107 2696
rect 1165 2664 1171 2676
rect 1101 2564 1107 2596
rect 1117 2524 1123 2536
rect 1165 2504 1171 2656
rect 1181 2604 1187 2636
rect 1181 2544 1187 2576
rect 1197 2524 1203 2676
rect 1213 2544 1219 2696
rect 1229 2684 1235 2696
rect 1293 2684 1299 2856
rect 1325 2783 1331 2876
rect 1352 2806 1358 2814
rect 1366 2806 1372 2814
rect 1380 2806 1386 2814
rect 1394 2806 1400 2814
rect 1325 2777 1347 2783
rect 1309 2684 1315 2696
rect 1341 2684 1347 2777
rect 1373 2724 1379 2736
rect 1252 2677 1260 2683
rect 1261 2564 1267 2676
rect 1325 2664 1331 2676
rect 1341 2644 1347 2676
rect 1277 2544 1283 2636
rect 1373 2544 1379 2636
rect 1421 2544 1427 3076
rect 1469 3064 1475 3076
rect 1501 3024 1507 3036
rect 1437 2784 1443 2896
rect 1453 2764 1459 3016
rect 1533 2944 1539 3116
rect 1565 3104 1571 3117
rect 1565 3084 1571 3096
rect 1581 3084 1587 3096
rect 1725 3064 1731 3236
rect 1869 3104 1875 3236
rect 1933 3102 1939 3116
rect 1997 3104 2003 3136
rect 1597 3024 1603 3036
rect 1549 2964 1555 3016
rect 1565 2984 1571 2996
rect 1517 2937 1532 2943
rect 1485 2904 1491 2916
rect 1469 2723 1475 2876
rect 1485 2724 1491 2736
rect 1453 2717 1475 2723
rect 1453 2704 1459 2717
rect 1517 2684 1523 2937
rect 1533 2904 1539 2916
rect 1581 2904 1587 2956
rect 1597 2944 1603 2956
rect 1613 2924 1619 3056
rect 1693 2984 1699 3056
rect 1677 2964 1683 2976
rect 1709 2964 1715 3036
rect 1789 2984 1795 3036
rect 1757 2944 1763 2976
rect 1757 2924 1763 2936
rect 1805 2924 1811 3036
rect 1821 2924 1827 2976
rect 1837 2944 1843 3036
rect 1853 2924 1859 2936
rect 1869 2924 1875 3096
rect 2109 3084 2115 3336
rect 2285 3284 2291 3336
rect 2125 3102 2131 3196
rect 2285 3124 2291 3156
rect 2301 3103 2307 3336
rect 2413 3304 2419 3376
rect 2429 3364 2435 3476
rect 2477 3464 2483 3496
rect 2493 3484 2499 3496
rect 2445 3344 2451 3456
rect 2493 3444 2499 3476
rect 2461 3344 2467 3356
rect 2445 3324 2451 3336
rect 2349 3124 2355 3176
rect 2292 3097 2307 3103
rect 2109 2964 2115 3076
rect 2221 3063 2227 3096
rect 2301 3084 2307 3097
rect 2205 3062 2227 3063
rect 2212 3057 2227 3062
rect 2205 2924 2211 3054
rect 2324 3017 2339 3023
rect 2221 2958 2236 2963
rect 2221 2957 2243 2958
rect 2221 2924 2227 2957
rect 1620 2917 1635 2923
rect 1629 2884 1635 2917
rect 1741 2844 1747 2916
rect 1853 2884 1859 2896
rect 1533 2684 1539 2716
rect 1549 2664 1555 2676
rect 1565 2544 1571 2836
rect 1693 2744 1699 2836
rect 1661 2684 1667 2716
rect 1597 2664 1603 2676
rect 1581 2584 1587 2656
rect 1549 2524 1555 2536
rect 1309 2384 1315 2436
rect 1352 2406 1358 2414
rect 1366 2406 1372 2414
rect 1380 2406 1386 2414
rect 1394 2406 1400 2414
rect 1101 2302 1107 2376
rect 1293 2302 1299 2336
rect 1405 2284 1411 2316
rect 1501 2284 1507 2516
rect 1597 2484 1603 2536
rect 1613 2504 1619 2516
rect 1581 2477 1596 2483
rect 1517 2284 1523 2416
rect 1581 2304 1587 2477
rect 1629 2324 1635 2516
rect 1645 2504 1651 2656
rect 1677 2604 1683 2676
rect 1757 2644 1763 2836
rect 1789 2724 1795 2736
rect 1869 2704 1875 2916
rect 1917 2702 1923 2736
rect 1709 2584 1715 2596
rect 1693 2544 1699 2576
rect 1693 2524 1699 2536
rect 1581 2284 1587 2296
rect 1101 2144 1107 2256
rect 1165 2224 1171 2236
rect 1325 2144 1331 2276
rect 1181 2124 1187 2136
rect 1213 1884 1219 1956
rect 1277 1884 1283 2136
rect 1437 2124 1443 2236
rect 1629 2124 1635 2236
rect 1645 2164 1651 2236
rect 1709 2124 1715 2276
rect 1741 2183 1747 2636
rect 1821 2544 1827 2636
rect 1757 2484 1763 2516
rect 1773 2484 1779 2496
rect 1789 2383 1795 2516
rect 1821 2504 1827 2536
rect 1773 2377 1795 2383
rect 1773 2302 1779 2377
rect 1805 2284 1811 2456
rect 1821 2424 1827 2496
rect 1853 2464 1859 2676
rect 1901 2564 1907 2596
rect 1981 2564 1987 2596
rect 1997 2564 2003 2576
rect 1869 2544 1875 2556
rect 1933 2524 1939 2556
rect 2061 2524 2067 2696
rect 2173 2684 2179 2716
rect 2285 2704 2291 2836
rect 2157 2524 2163 2636
rect 2317 2564 2323 2936
rect 2333 2924 2339 3017
rect 2349 2664 2355 3116
rect 2397 3104 2403 3296
rect 2445 3144 2451 3236
rect 2413 3064 2419 3136
rect 2445 3084 2451 3116
rect 2461 3104 2467 3336
rect 2477 3304 2483 3436
rect 2541 3384 2547 3476
rect 2557 3464 2563 3516
rect 2637 3484 2643 3657
rect 2669 3544 2675 3636
rect 2765 3504 2771 3536
rect 2813 3523 2819 3836
rect 2829 3744 2835 3876
rect 2989 3864 2995 3876
rect 3021 3864 3027 3896
rect 3181 3884 3187 4037
rect 2861 3704 2867 3836
rect 2877 3784 2883 3816
rect 2904 3806 2910 3814
rect 2918 3806 2924 3814
rect 2932 3806 2938 3814
rect 2946 3806 2952 3814
rect 2813 3517 2828 3523
rect 2653 3484 2659 3496
rect 2749 3484 2755 3496
rect 2516 3377 2531 3383
rect 2509 3344 2515 3376
rect 2525 3324 2531 3377
rect 2541 3364 2547 3376
rect 2509 3304 2515 3316
rect 2477 3124 2483 3296
rect 2541 3284 2547 3316
rect 2557 3304 2563 3456
rect 2621 3424 2627 3436
rect 2621 3344 2627 3396
rect 2637 3364 2643 3476
rect 2669 3384 2675 3396
rect 2701 3364 2707 3376
rect 2461 2983 2467 3096
rect 2493 3064 2499 3136
rect 2509 3084 2515 3096
rect 2525 3084 2531 3096
rect 2541 2984 2547 3276
rect 2557 3264 2563 3276
rect 2557 3124 2563 3256
rect 2605 3164 2611 3236
rect 2637 3104 2643 3136
rect 2669 3104 2675 3296
rect 2685 3184 2691 3356
rect 2717 3124 2723 3416
rect 2749 3344 2755 3456
rect 2765 3344 2771 3476
rect 2829 3384 2835 3516
rect 2861 3484 2867 3696
rect 2893 3584 2899 3716
rect 2925 3504 2931 3536
rect 2941 3504 2947 3516
rect 2989 3504 2995 3856
rect 3021 3764 3027 3856
rect 3053 3744 3059 3796
rect 3021 3704 3027 3736
rect 3101 3704 3107 3836
rect 3117 3804 3123 3876
rect 3181 3764 3187 3876
rect 3197 3724 3203 4096
rect 3245 3924 3251 3976
rect 3277 3904 3283 3936
rect 3229 3864 3235 3876
rect 3277 3864 3283 3896
rect 2941 3484 2947 3496
rect 2845 3364 2851 3456
rect 2904 3406 2910 3414
rect 2918 3406 2924 3414
rect 2932 3406 2938 3414
rect 2946 3406 2952 3414
rect 2989 3364 2995 3436
rect 3069 3364 3075 3636
rect 3229 3524 3235 3796
rect 3309 3784 3315 3976
rect 3421 3884 3427 3894
rect 3549 3884 3555 4116
rect 3389 3724 3395 3876
rect 3613 3864 3619 3896
rect 3501 3857 3516 3863
rect 3501 3744 3507 3857
rect 3677 3863 3683 4016
rect 3693 3884 3699 3896
rect 3677 3857 3699 3863
rect 3437 3726 3443 3736
rect 3245 3704 3251 3718
rect 3501 3724 3507 3736
rect 3517 3724 3523 3756
rect 3613 3744 3619 3856
rect 3629 3764 3635 3836
rect 3645 3744 3651 3856
rect 3693 3784 3699 3857
rect 3725 3784 3731 4136
rect 3757 4104 3763 4136
rect 3869 4104 3875 4136
rect 3741 3884 3747 3896
rect 3885 3884 3891 4176
rect 3933 4144 3939 4176
rect 3981 4104 3987 4136
rect 4013 4084 4019 4156
rect 4221 4144 4227 4243
rect 4221 4104 4227 4136
rect 4333 4104 4339 4136
rect 4029 4004 4035 4036
rect 4109 3884 4115 4036
rect 4381 3924 4387 4243
rect 4589 4237 4611 4243
rect 4605 4184 4611 4237
rect 4781 4204 4787 4243
rect 4397 4144 4403 4176
rect 4221 3897 4236 3903
rect 4189 3884 4195 3896
rect 4221 3884 4227 3897
rect 3741 3764 3747 3876
rect 3853 3777 3868 3783
rect 3853 3764 3859 3777
rect 3732 3757 3740 3763
rect 3629 3724 3635 3736
rect 3677 3724 3683 3756
rect 3821 3744 3827 3756
rect 3853 3744 3859 3756
rect 3133 3464 3139 3496
rect 3261 3484 3267 3496
rect 3213 3464 3219 3476
rect 3085 3404 3091 3456
rect 3117 3424 3123 3436
rect 3133 3404 3139 3456
rect 3277 3444 3283 3476
rect 3309 3464 3315 3536
rect 3117 3364 3123 3396
rect 2733 3324 2739 3336
rect 2749 3324 2755 3336
rect 2765 3304 2771 3336
rect 2845 3324 2851 3356
rect 2893 3144 2899 3236
rect 2717 3104 2723 3116
rect 2452 2977 2467 2983
rect 2461 2944 2467 2956
rect 2573 2943 2579 3076
rect 2564 2937 2579 2943
rect 2701 2926 2707 2936
rect 2829 2924 2835 3076
rect 2904 3006 2910 3014
rect 2918 3006 2924 3014
rect 2932 3006 2938 3014
rect 2946 3006 2952 3014
rect 2397 2684 2403 2716
rect 2413 2704 2419 2716
rect 2493 2704 2499 2716
rect 2573 2684 2579 2696
rect 2445 2664 2451 2676
rect 2605 2604 2611 2836
rect 2621 2664 2627 2676
rect 2301 2524 2307 2556
rect 2413 2524 2419 2576
rect 2557 2526 2563 2536
rect 2589 2524 2595 2536
rect 2637 2524 2643 2916
rect 2973 2904 2979 3036
rect 3005 2944 3011 3336
rect 3021 3324 3027 3356
rect 3149 3344 3155 3376
rect 3181 3364 3187 3416
rect 3197 3364 3203 3436
rect 3197 3323 3203 3356
rect 3325 3344 3331 3396
rect 3341 3384 3347 3616
rect 3389 3504 3395 3716
rect 3533 3704 3539 3716
rect 3533 3464 3539 3696
rect 3549 3684 3555 3696
rect 3645 3504 3651 3716
rect 3757 3704 3763 3716
rect 3773 3704 3779 3716
rect 3805 3704 3811 3716
rect 3661 3684 3667 3696
rect 3773 3683 3779 3696
rect 3757 3677 3779 3683
rect 3693 3584 3699 3636
rect 3453 3344 3459 3456
rect 3565 3384 3571 3396
rect 3549 3324 3555 3356
rect 3677 3344 3683 3456
rect 3757 3404 3763 3677
rect 3789 3484 3795 3576
rect 3885 3564 3891 3876
rect 3901 3764 3907 3836
rect 3933 3724 3939 3776
rect 4029 3484 4035 3856
rect 4109 3744 4115 3876
rect 4333 3824 4339 3876
rect 4349 3804 4355 3836
rect 4109 3544 4115 3736
rect 4189 3524 4195 3716
rect 4173 3504 4179 3516
rect 3757 3344 3763 3396
rect 3197 3317 3212 3323
rect 3261 3204 3267 3236
rect 3101 3102 3107 3136
rect 3165 3104 3171 3116
rect 3277 3104 3283 3116
rect 3309 3104 3315 3116
rect 3037 3084 3043 3096
rect 3213 2944 3219 3076
rect 3325 3064 3331 3116
rect 3373 3084 3379 3156
rect 3389 3084 3395 3116
rect 3229 2944 3235 3036
rect 2685 2724 2691 2736
rect 2797 2664 2803 2676
rect 2829 2664 2835 2896
rect 3037 2704 3043 2896
rect 3053 2744 3059 2936
rect 2957 2684 2963 2696
rect 3053 2684 3059 2736
rect 3133 2724 3139 2736
rect 3117 2704 3123 2716
rect 3092 2697 3107 2703
rect 2845 2664 2851 2676
rect 3101 2644 3107 2697
rect 3181 2684 3187 2836
rect 3213 2723 3219 2936
rect 3197 2717 3219 2723
rect 3197 2684 3203 2717
rect 3277 2704 3283 2956
rect 3405 2944 3411 3316
rect 3517 3184 3523 3276
rect 3421 3104 3427 3156
rect 3437 3104 3443 3116
rect 3533 3104 3539 3136
rect 3549 3084 3555 3136
rect 3645 3084 3651 3176
rect 3757 3124 3763 3336
rect 3837 3324 3843 3436
rect 3901 3364 3907 3436
rect 3917 3404 3923 3476
rect 3933 3404 3939 3436
rect 3869 3324 3875 3336
rect 3773 3284 3779 3316
rect 3773 3164 3779 3236
rect 3789 3184 3795 3296
rect 3805 3244 3811 3316
rect 3757 3104 3763 3116
rect 3437 3064 3443 3076
rect 3757 3064 3763 3076
rect 3437 3004 3443 3056
rect 3677 2984 3683 2996
rect 3693 2944 3699 3036
rect 3773 3024 3779 3076
rect 3821 3064 3827 3216
rect 3853 3184 3859 3316
rect 3885 3244 3891 3336
rect 3901 3224 3907 3336
rect 4029 3324 4035 3476
rect 4189 3404 4195 3516
rect 4077 3326 4083 3376
rect 3917 3104 3923 3236
rect 3917 3044 3923 3096
rect 3933 3084 3939 3296
rect 3949 3224 3955 3236
rect 4109 3104 4115 3336
rect 4141 3084 4147 3236
rect 4173 3102 4179 3176
rect 3965 3064 3971 3076
rect 4013 3057 4028 3063
rect 3405 2924 3411 2936
rect 3613 2926 3619 2936
rect 3421 2884 3427 2918
rect 3485 2744 3491 2836
rect 3645 2724 3651 2736
rect 3117 2664 3123 2676
rect 2733 2564 2739 2636
rect 2904 2606 2910 2614
rect 2918 2606 2924 2614
rect 2932 2606 2938 2614
rect 2946 2606 2952 2614
rect 3197 2584 3203 2676
rect 3245 2624 3251 2696
rect 2893 2524 2899 2576
rect 3197 2544 3203 2556
rect 3245 2544 3251 2616
rect 3261 2564 3267 2676
rect 3293 2664 3299 2676
rect 3309 2623 3315 2716
rect 3549 2702 3555 2716
rect 3613 2684 3619 2696
rect 3309 2617 3331 2623
rect 3293 2584 3299 2616
rect 3277 2544 3283 2576
rect 3309 2544 3315 2576
rect 3325 2544 3331 2617
rect 3325 2524 3331 2536
rect 3341 2524 3347 2656
rect 3421 2644 3427 2676
rect 3453 2584 3459 2656
rect 3405 2564 3411 2576
rect 3485 2557 3500 2563
rect 3485 2544 3491 2557
rect 3437 2524 3443 2536
rect 1853 2304 1859 2436
rect 2061 2303 2067 2516
rect 2052 2297 2067 2303
rect 2109 2302 2115 2336
rect 2253 2303 2259 2516
rect 2381 2344 2387 2436
rect 2397 2324 2403 2336
rect 2244 2297 2259 2303
rect 2301 2302 2307 2316
rect 2429 2304 2435 2436
rect 2589 2344 2595 2516
rect 2749 2504 2755 2518
rect 3229 2503 3235 2516
rect 3229 2497 3244 2503
rect 3133 2484 3139 2496
rect 3277 2324 3283 2336
rect 2877 2317 2892 2323
rect 2461 2284 2467 2296
rect 2493 2284 2499 2294
rect 1805 2184 1811 2276
rect 1837 2264 1843 2276
rect 2365 2244 2371 2256
rect 2381 2244 2387 2276
rect 1741 2177 1763 2183
rect 1352 2006 1358 2014
rect 1366 2006 1372 2014
rect 1380 2006 1386 2014
rect 1394 2006 1400 2014
rect 1117 1744 1123 1836
rect 813 1717 835 1723
rect 781 1464 787 1476
rect 605 1384 611 1436
rect 621 1343 627 1396
rect 605 1337 627 1343
rect 573 1324 579 1336
rect 509 1184 515 1296
rect 429 1084 435 1096
rect 333 1044 339 1056
rect 269 944 275 956
rect 189 723 195 896
rect 205 784 211 916
rect 253 744 259 916
rect 317 904 323 956
rect 365 924 371 1076
rect 381 944 387 1076
rect 461 1024 467 1116
rect 477 1084 483 1176
rect 477 1064 483 1076
rect 493 1044 499 1116
rect 493 944 499 1036
rect 525 983 531 1176
rect 541 1164 547 1296
rect 605 1104 611 1337
rect 621 1304 627 1316
rect 653 1304 659 1336
rect 685 1324 691 1356
rect 749 1324 755 1416
rect 637 1244 643 1276
rect 637 1104 643 1236
rect 653 1144 659 1296
rect 701 1104 707 1196
rect 717 1084 723 1236
rect 733 1204 739 1316
rect 749 1124 755 1316
rect 797 1304 803 1496
rect 829 1484 835 1717
rect 820 1477 828 1483
rect 829 1364 835 1436
rect 845 1363 851 1476
rect 861 1384 867 1496
rect 877 1463 883 1496
rect 877 1457 899 1463
rect 893 1444 899 1457
rect 845 1357 867 1363
rect 829 1184 835 1336
rect 845 1104 851 1116
rect 541 1064 547 1076
rect 605 1064 611 1076
rect 829 1064 835 1076
rect 509 977 531 983
rect 509 924 515 977
rect 557 924 563 1036
rect 605 944 611 956
rect 669 944 675 1036
rect 733 944 739 956
rect 653 924 659 936
rect 733 904 739 916
rect 781 904 787 936
rect 189 717 211 723
rect 125 684 131 696
rect 173 684 179 716
rect 157 664 163 676
rect 125 563 131 636
rect 157 564 163 656
rect 205 624 211 717
rect 221 664 227 716
rect 109 557 131 563
rect 13 264 19 516
rect 45 204 51 556
rect 109 544 115 557
rect 205 544 211 616
rect 237 544 243 736
rect 269 724 275 756
rect 285 724 291 776
rect 301 703 307 816
rect 397 764 403 896
rect 541 884 547 896
rect 573 864 579 876
rect 781 784 787 896
rect 413 704 419 776
rect 829 764 835 1056
rect 845 964 851 1096
rect 861 1024 867 1357
rect 877 1244 883 1336
rect 893 1284 899 1436
rect 909 1404 915 1436
rect 925 1384 931 1476
rect 909 1364 915 1376
rect 941 1324 947 1736
rect 1037 1624 1043 1736
rect 1197 1704 1203 1836
rect 1037 1524 1043 1536
rect 989 1464 995 1496
rect 1069 1484 1075 1496
rect 1037 1444 1043 1456
rect 1037 1344 1043 1436
rect 1085 1344 1091 1556
rect 1101 1544 1107 1636
rect 1101 1464 1107 1536
rect 1117 1484 1123 1616
rect 1213 1484 1219 1876
rect 1533 1824 1539 2036
rect 1565 1904 1571 2116
rect 1709 1884 1715 2116
rect 1725 1864 1731 2036
rect 1757 1904 1763 2177
rect 1917 2164 1923 2236
rect 1837 2124 1843 2136
rect 1917 2124 1923 2156
rect 2045 2144 2051 2176
rect 1805 1904 1811 2036
rect 1869 1964 1875 2096
rect 1885 2084 1891 2116
rect 1933 2084 1939 2116
rect 1965 2104 1971 2136
rect 2077 2126 2083 2136
rect 2173 2124 2179 2236
rect 2253 2164 2259 2176
rect 2381 2123 2387 2236
rect 2413 2124 2419 2136
rect 2477 2124 2483 2136
rect 2589 2126 2595 2136
rect 2372 2117 2387 2123
rect 2653 2124 2659 2276
rect 2013 2084 2019 2096
rect 2333 2084 2339 2096
rect 1629 1837 1644 1843
rect 1453 1724 1459 1736
rect 1389 1664 1395 1718
rect 1229 1584 1235 1636
rect 1352 1606 1358 1614
rect 1366 1606 1372 1614
rect 1380 1606 1386 1614
rect 1394 1606 1400 1614
rect 1085 1324 1091 1336
rect 1117 1304 1123 1476
rect 1165 1344 1171 1464
rect 1213 1384 1219 1456
rect 1229 1444 1235 1496
rect 1133 1337 1148 1343
rect 1133 1324 1139 1337
rect 973 1284 979 1296
rect 1021 1204 1027 1236
rect 1053 1224 1059 1296
rect 1085 1124 1091 1156
rect 973 1104 979 1116
rect 1117 1104 1123 1116
rect 877 984 883 1076
rect 893 1064 899 1076
rect 845 944 851 956
rect 909 944 915 1036
rect 1005 984 1011 1036
rect 1053 984 1059 1036
rect 1069 964 1075 1076
rect 1085 964 1091 1096
rect 1101 1064 1107 1076
rect 989 924 995 956
rect 1085 924 1091 956
rect 1117 943 1123 1096
rect 1108 937 1123 943
rect 669 724 675 756
rect 445 704 451 716
rect 301 697 316 703
rect 429 684 435 696
rect 317 644 323 656
rect 93 504 99 516
rect 109 363 115 536
rect 93 357 115 363
rect 93 303 99 357
rect 125 324 131 536
rect 253 524 259 576
rect 141 504 147 516
rect 189 504 195 516
rect 173 304 179 436
rect 269 344 275 636
rect 301 544 307 576
rect 317 524 323 636
rect 333 604 339 676
rect 381 644 387 656
rect 333 564 339 596
rect 349 544 355 636
rect 365 544 371 556
rect 349 504 355 536
rect 381 524 387 556
rect 413 544 419 576
rect 429 524 435 616
rect 461 484 467 676
rect 509 644 515 656
rect 557 624 563 696
rect 573 564 579 676
rect 605 564 611 676
rect 637 644 643 716
rect 749 684 755 716
rect 765 684 771 756
rect 797 704 803 736
rect 1021 724 1027 916
rect 973 684 979 716
rect 1037 684 1043 796
rect 1133 744 1139 1316
rect 1149 1244 1155 1316
rect 1181 1284 1187 1376
rect 1181 1184 1187 1276
rect 1149 1124 1155 1176
rect 1149 964 1155 996
rect 637 564 643 636
rect 477 537 508 543
rect 477 524 483 537
rect 541 524 547 556
rect 669 544 675 556
rect 205 324 211 336
rect 301 304 307 356
rect 429 344 435 476
rect 397 304 403 316
rect 429 304 435 336
rect 445 304 451 436
rect 509 384 515 496
rect 557 384 563 496
rect 525 304 531 336
rect 77 297 99 303
rect 13 164 19 196
rect 61 84 67 236
rect 77 124 83 297
rect 93 104 99 276
rect 141 264 147 296
rect 317 284 323 296
rect 173 264 179 276
rect 413 264 419 276
rect 493 264 499 296
rect 589 284 595 436
rect 637 324 643 436
rect 685 284 691 376
rect 701 344 707 636
rect 749 524 755 676
rect 765 664 771 676
rect 861 664 867 676
rect 925 664 931 676
rect 941 664 947 676
rect 973 663 979 676
rect 1037 664 1043 676
rect 973 657 995 663
rect 781 564 787 636
rect 797 544 803 616
rect 893 563 899 636
rect 973 584 979 636
rect 893 557 915 563
rect 813 524 819 556
rect 765 484 771 516
rect 861 504 867 556
rect 909 524 915 557
rect 989 544 995 657
rect 1053 644 1059 696
rect 909 504 915 516
rect 957 504 963 536
rect 1005 484 1011 636
rect 1069 564 1075 656
rect 1085 624 1091 716
rect 1165 704 1171 1096
rect 1229 1064 1235 1436
rect 1261 1344 1267 1496
rect 1277 1424 1283 1456
rect 1293 1384 1299 1496
rect 1357 1424 1363 1496
rect 1421 1484 1427 1536
rect 1517 1464 1523 1636
rect 1581 1502 1587 1516
rect 1629 1444 1635 1837
rect 1853 1824 1859 1856
rect 1725 1744 1731 1816
rect 1869 1784 1875 1836
rect 1821 1724 1827 1736
rect 1645 1504 1651 1716
rect 1709 1624 1715 1636
rect 1485 1364 1491 1436
rect 1469 1344 1475 1356
rect 1581 1344 1587 1436
rect 1645 1364 1651 1496
rect 1245 1004 1251 1036
rect 1261 984 1267 1316
rect 1485 1304 1491 1336
rect 1277 1284 1283 1296
rect 1352 1206 1358 1214
rect 1366 1206 1372 1214
rect 1380 1206 1386 1214
rect 1394 1206 1400 1214
rect 1309 1104 1315 1176
rect 1341 1104 1347 1116
rect 1277 1064 1283 1076
rect 1197 977 1235 983
rect 1197 944 1203 977
rect 1229 963 1235 977
rect 1229 957 1244 963
rect 1213 924 1219 956
rect 1213 824 1219 856
rect 1101 644 1107 696
rect 1181 624 1187 676
rect 1197 624 1203 696
rect 1213 684 1219 816
rect 1101 544 1107 556
rect 1133 544 1139 616
rect 1021 524 1027 536
rect 1117 524 1123 536
rect 1149 524 1155 616
rect 1213 584 1219 636
rect 1229 564 1235 636
rect 1229 544 1235 556
rect 1245 523 1251 916
rect 1277 723 1283 1056
rect 1309 964 1315 1096
rect 1341 924 1347 976
rect 1268 717 1283 723
rect 1293 604 1299 916
rect 1405 904 1411 936
rect 1352 806 1358 814
rect 1366 806 1372 814
rect 1380 806 1386 814
rect 1394 806 1400 814
rect 1309 684 1315 736
rect 1373 684 1379 736
rect 1421 704 1427 1236
rect 1485 1123 1491 1296
rect 1581 1283 1587 1336
rect 1709 1324 1715 1436
rect 1837 1424 1843 1736
rect 1853 1724 1859 1756
rect 1853 1484 1859 1696
rect 1885 1564 1891 1916
rect 1901 1744 1907 1956
rect 1933 1884 1939 2076
rect 1981 1964 1987 2036
rect 2013 1903 2019 2076
rect 2173 1924 2179 2076
rect 2397 2064 2403 2096
rect 2013 1897 2028 1903
rect 2061 1883 2067 1916
rect 2237 1884 2243 1956
rect 2269 1884 2275 1916
rect 2301 1902 2307 1936
rect 2429 1923 2435 2116
rect 2461 2084 2467 2096
rect 2429 1917 2444 1923
rect 2477 1904 2483 2116
rect 2493 2104 2499 2116
rect 2493 1884 2499 2056
rect 2525 2044 2531 2096
rect 2701 2084 2707 2296
rect 2813 2244 2819 2256
rect 2733 2164 2739 2236
rect 2829 2184 2835 2256
rect 2845 2184 2851 2296
rect 2829 2143 2835 2176
rect 2877 2144 2883 2317
rect 3453 2302 3459 2496
rect 3517 2304 3523 2676
rect 3709 2644 3715 2676
rect 3565 2544 3571 2556
rect 3533 2504 3539 2516
rect 3581 2504 3587 2616
rect 3725 2604 3731 2716
rect 3773 2704 3779 3016
rect 3949 2984 3955 3036
rect 3869 2944 3875 2976
rect 3805 2864 3811 2918
rect 3981 2904 3987 3036
rect 4013 2924 4019 3057
rect 4141 2984 4147 3016
rect 3821 2724 3827 2736
rect 3821 2684 3827 2716
rect 3837 2704 3843 2896
rect 3981 2784 3987 2896
rect 4029 2744 4035 2936
rect 4045 2904 4051 2956
rect 4093 2917 4108 2923
rect 4093 2784 4099 2917
rect 4125 2903 4131 2936
rect 4205 2924 4211 3776
rect 4285 3764 4291 3776
rect 4381 3744 4387 3916
rect 4397 3824 4403 4136
rect 4493 4104 4499 4136
rect 4509 4084 4515 4156
rect 4557 4083 4563 4116
rect 4548 4077 4563 4083
rect 4440 4006 4446 4014
rect 4454 4006 4460 4014
rect 4468 4006 4474 4014
rect 4482 4006 4488 4014
rect 4445 3804 4451 3836
rect 4381 3708 4387 3716
rect 4253 3484 4259 3536
rect 4317 3524 4323 3536
rect 4269 3504 4275 3516
rect 4269 3484 4275 3496
rect 4237 3464 4243 3476
rect 4397 3464 4403 3796
rect 4509 3764 4515 4076
rect 4573 4004 4579 4116
rect 4637 3884 4643 3916
rect 4749 3884 4755 3916
rect 4797 3864 4803 4156
rect 4829 4144 4835 4243
rect 4829 4104 4835 4136
rect 4893 3924 4899 4243
rect 5085 4143 5091 4243
rect 5069 4137 5091 4143
rect 4941 4104 4947 4136
rect 4861 3884 4867 3916
rect 4605 3784 4611 3856
rect 4749 3764 4755 3856
rect 4813 3824 4819 3876
rect 4877 3764 4883 3856
rect 4440 3606 4446 3614
rect 4454 3606 4460 3614
rect 4468 3606 4474 3614
rect 4482 3606 4488 3614
rect 4493 3464 4499 3476
rect 4509 3464 4515 3516
rect 4573 3504 4579 3516
rect 4429 3444 4435 3456
rect 4301 3344 4307 3436
rect 4493 3324 4499 3396
rect 4365 3284 4371 3316
rect 4237 3084 4243 3096
rect 4253 3084 4259 3116
rect 4253 2924 4259 3036
rect 4109 2897 4131 2903
rect 4109 2784 4115 2897
rect 3853 2724 3859 2736
rect 3965 2717 3980 2723
rect 3885 2704 3891 2716
rect 3661 2564 3667 2576
rect 3661 2524 3667 2556
rect 3677 2544 3683 2576
rect 3741 2544 3747 2676
rect 3837 2644 3843 2696
rect 3869 2524 3875 2696
rect 3901 2684 3907 2696
rect 3965 2664 3971 2717
rect 4029 2684 4035 2736
rect 4061 2664 4067 2696
rect 4125 2664 4131 2736
rect 4205 2704 4211 2916
rect 3933 2644 3939 2656
rect 3885 2544 3891 2636
rect 3917 2544 3923 2636
rect 3933 2524 3939 2596
rect 3965 2584 3971 2636
rect 3981 2604 3987 2636
rect 4061 2584 4067 2656
rect 4093 2524 4099 2636
rect 4109 2564 4115 2636
rect 4221 2344 4227 2736
rect 4269 2702 4275 3256
rect 4440 3206 4446 3214
rect 4454 3206 4460 3214
rect 4468 3206 4474 3214
rect 4482 3206 4488 3214
rect 4285 3084 4291 3156
rect 4445 3124 4451 3136
rect 4349 3104 4355 3116
rect 4381 3104 4387 3116
rect 4509 3084 4515 3396
rect 4557 3324 4563 3436
rect 4573 3264 4579 3496
rect 4589 3484 4595 3636
rect 4749 3544 4755 3756
rect 4893 3744 4899 3916
rect 4909 3703 4915 3836
rect 4925 3824 4931 3876
rect 4900 3697 4915 3703
rect 4989 3644 4995 3896
rect 5005 3824 5011 4136
rect 5053 4104 5059 4136
rect 5069 3984 5075 4137
rect 5149 4124 5155 4156
rect 5085 4004 5091 4116
rect 5197 4044 5203 4100
rect 5293 4043 5299 4156
rect 5277 4037 5299 4043
rect 5021 3764 5027 3836
rect 5101 3804 5107 3896
rect 5021 3724 5027 3756
rect 5117 3744 5123 3958
rect 5181 3920 5187 3958
rect 5149 3844 5155 3896
rect 5245 3804 5251 3876
rect 5277 3864 5283 4037
rect 5373 4024 5379 4116
rect 5437 3984 5443 4136
rect 5453 3884 5459 4036
rect 5149 3724 5155 3756
rect 5277 3724 5283 3856
rect 5309 3784 5315 3796
rect 5325 3744 5331 3816
rect 5469 3744 5475 4116
rect 5021 3644 5027 3696
rect 5117 3584 5123 3716
rect 5421 3644 5427 3716
rect 4637 3504 4643 3516
rect 4941 3502 4947 3503
rect 4589 3464 4595 3476
rect 4589 3304 4595 3456
rect 4605 3344 4611 3436
rect 4637 3364 4643 3476
rect 4685 3324 4691 3436
rect 4701 3344 4707 3396
rect 4733 3384 4739 3436
rect 4749 3384 4755 3464
rect 4877 3324 4883 3476
rect 4941 3384 4947 3494
rect 5005 3484 5011 3556
rect 4973 3344 4979 3476
rect 5117 3444 5123 3456
rect 5117 3324 5123 3436
rect 5149 3324 5155 3558
rect 5213 3520 5219 3558
rect 5213 3384 5219 3476
rect 5309 3404 5315 3456
rect 5453 3403 5459 3636
rect 5453 3397 5475 3403
rect 5373 3364 5379 3396
rect 5405 3344 5411 3356
rect 5469 3324 5475 3397
rect 5501 3364 5507 4036
rect 5661 4024 5667 4156
rect 5789 4044 5795 4096
rect 5517 3904 5523 4016
rect 5533 3920 5539 3958
rect 5517 3724 5523 3896
rect 5629 3864 5635 4016
rect 5629 3823 5635 3856
rect 5629 3817 5651 3823
rect 5645 3764 5651 3817
rect 5517 3504 5523 3716
rect 5549 3644 5555 3700
rect 5645 3643 5651 3756
rect 5789 3744 5795 3836
rect 5805 3784 5811 4136
rect 5645 3637 5667 3643
rect 5533 3524 5539 3576
rect 5533 3344 5539 3496
rect 5661 3464 5667 3637
rect 5661 3404 5667 3456
rect 5789 3324 5795 3436
rect 4557 3123 4563 3236
rect 4548 3117 4563 3123
rect 4413 3064 4419 3076
rect 4333 2944 4339 3036
rect 4493 2964 4499 3036
rect 4525 2944 4531 3076
rect 4525 2904 4531 2936
rect 4541 2924 4547 3116
rect 4589 3104 4595 3136
rect 4637 3084 4643 3276
rect 4765 3184 4771 3256
rect 4749 3084 4755 3096
rect 4621 3044 4627 3056
rect 4813 3044 4819 3096
rect 4861 3063 4867 3316
rect 5005 3184 5011 3318
rect 5341 3084 5347 3116
rect 5165 3064 5171 3076
rect 5373 3064 5379 3076
rect 5469 3064 5475 3316
rect 5501 3244 5507 3296
rect 4861 3057 4883 3063
rect 4440 2806 4446 2814
rect 4454 2806 4460 2814
rect 4468 2806 4474 2814
rect 4482 2806 4488 2814
rect 4557 2784 4563 3036
rect 4621 2944 4627 3036
rect 4877 2984 4883 3057
rect 5165 2944 5171 3056
rect 4573 2884 4579 2896
rect 4621 2784 4627 2916
rect 4333 2704 4339 2736
rect 4413 2677 4428 2683
rect 4301 2544 4307 2676
rect 4349 2604 4355 2636
rect 4365 2583 4371 2656
rect 4349 2577 4371 2583
rect 4317 2526 4323 2576
rect 3588 2337 3603 2343
rect 3597 2304 3603 2337
rect 4253 2324 4259 2356
rect 4301 2304 4307 2336
rect 2957 2284 2963 2296
rect 2904 2206 2910 2214
rect 2918 2206 2924 2214
rect 2932 2206 2938 2214
rect 2946 2206 2952 2214
rect 2941 2164 2947 2176
rect 2989 2164 2995 2176
rect 3101 2144 3107 2276
rect 3149 2224 3155 2296
rect 3629 2284 3635 2296
rect 3325 2244 3331 2256
rect 2820 2137 2835 2143
rect 3181 2124 3187 2136
rect 2653 1984 2659 2076
rect 2733 1924 2739 2096
rect 2052 1877 2067 1883
rect 1981 1864 1987 1876
rect 1933 1744 1939 1776
rect 1965 1724 1971 1836
rect 2077 1783 2083 1836
rect 2077 1777 2099 1783
rect 2013 1744 2019 1756
rect 2045 1744 2051 1776
rect 2093 1764 2099 1777
rect 2109 1764 2115 1836
rect 2109 1744 2115 1756
rect 1981 1704 1987 1716
rect 1997 1704 2003 1736
rect 2173 1704 2179 1756
rect 2349 1744 2355 1876
rect 2429 1844 2435 1856
rect 2493 1744 2499 1876
rect 2509 1864 2515 1896
rect 2765 1884 2771 2116
rect 2813 2084 2819 2096
rect 2989 1884 2995 2036
rect 3037 1904 3043 1916
rect 2685 1864 2691 1876
rect 2525 1744 2531 1796
rect 2765 1744 2771 1876
rect 2925 1844 2931 1856
rect 2904 1806 2910 1814
rect 2918 1806 2924 1814
rect 2932 1806 2938 1814
rect 2946 1806 2952 1814
rect 2237 1704 2243 1736
rect 2269 1704 2275 1716
rect 2317 1684 2323 1696
rect 2253 1504 2259 1516
rect 2141 1484 2147 1496
rect 1932 1464 1940 1470
rect 1821 1304 1827 1316
rect 1581 1277 1603 1283
rect 1517 1184 1523 1236
rect 1485 1117 1507 1123
rect 1501 1084 1507 1117
rect 1597 1084 1603 1277
rect 1693 1102 1699 1136
rect 1741 1104 1747 1276
rect 1773 1204 1779 1236
rect 1837 1084 1843 1336
rect 1885 1324 1891 1356
rect 1917 1344 1923 1464
rect 1933 1364 1939 1436
rect 1965 1344 1971 1476
rect 1981 1464 1987 1476
rect 2061 1364 2067 1416
rect 1981 1344 1987 1356
rect 1885 1144 1891 1296
rect 1917 1124 1923 1316
rect 1965 1304 1971 1336
rect 2093 1303 2099 1436
rect 2109 1304 2115 1316
rect 2084 1297 2099 1303
rect 1933 1124 1939 1236
rect 1917 1104 1923 1116
rect 2013 1104 2019 1176
rect 2045 1124 2051 1236
rect 2077 1184 2083 1296
rect 2125 1164 2131 1476
rect 2141 1344 2147 1456
rect 2237 1344 2243 1476
rect 2285 1464 2291 1476
rect 2324 1457 2339 1463
rect 2285 1444 2291 1456
rect 2269 1404 2275 1436
rect 2253 1344 2259 1376
rect 2301 1364 2307 1436
rect 2269 1344 2275 1356
rect 2333 1344 2339 1457
rect 2429 1384 2435 1476
rect 2445 1464 2451 1576
rect 2461 1484 2467 1496
rect 2157 1324 2163 1336
rect 2141 1224 2147 1316
rect 2237 1304 2243 1316
rect 1501 1064 1507 1076
rect 1597 1064 1603 1076
rect 1469 984 1475 1016
rect 1453 944 1459 976
rect 1533 924 1539 1036
rect 1453 904 1459 916
rect 1501 904 1507 916
rect 1533 904 1539 916
rect 1469 884 1475 896
rect 1565 864 1571 936
rect 1629 926 1635 936
rect 1437 704 1443 836
rect 1277 524 1283 596
rect 1325 564 1331 576
rect 1245 517 1267 523
rect 1149 504 1155 516
rect 733 384 739 436
rect 765 304 771 316
rect 813 304 819 436
rect 877 384 883 456
rect 925 324 931 436
rect 157 163 163 236
rect 205 184 211 236
rect 141 157 163 163
rect 141 124 147 157
rect 285 144 291 256
rect 349 204 355 236
rect 573 184 579 256
rect 765 184 771 196
rect 381 144 387 176
rect 797 144 803 296
rect 989 284 995 376
rect 1021 323 1027 436
rect 1012 317 1027 323
rect 1037 304 1043 336
rect 1053 284 1059 496
rect 1245 484 1251 496
rect 1181 304 1187 316
rect 157 104 163 136
rect 269 124 275 136
rect 605 124 611 136
rect 109 84 115 96
rect 349 84 355 96
rect 445 84 451 118
rect 989 124 995 136
rect 1021 126 1027 236
rect 829 104 835 118
rect 1085 124 1091 276
rect 1181 144 1187 296
rect 1261 284 1267 517
rect 1293 504 1299 536
rect 1341 443 1347 676
rect 1437 644 1443 676
rect 1533 664 1539 676
rect 1469 624 1475 636
rect 1405 524 1411 616
rect 1469 524 1475 556
rect 1325 437 1347 443
rect 1309 344 1315 436
rect 1325 304 1331 437
rect 1352 406 1358 414
rect 1366 406 1372 414
rect 1380 406 1386 414
rect 1394 406 1400 414
rect 1357 284 1363 296
rect 1229 124 1235 236
rect 1245 224 1251 236
rect 1341 184 1347 236
rect 1405 184 1411 356
rect 1485 324 1491 616
rect 1501 584 1507 596
rect 1517 544 1523 556
rect 1533 544 1539 636
rect 1565 604 1571 856
rect 1661 704 1667 936
rect 1693 924 1699 1056
rect 1837 984 1843 1076
rect 1757 964 1763 976
rect 1837 964 1843 976
rect 1757 784 1763 876
rect 1645 544 1651 656
rect 1661 624 1667 696
rect 1741 684 1747 736
rect 1773 703 1779 916
rect 1805 724 1811 956
rect 1853 784 1859 916
rect 1869 744 1875 916
rect 1885 723 1891 1076
rect 1965 1004 1971 1036
rect 1901 964 1907 976
rect 1965 944 1971 976
rect 2013 944 2019 1036
rect 2029 984 2035 1096
rect 2077 1084 2083 1116
rect 2093 1104 2099 1156
rect 2109 1104 2115 1116
rect 2141 1084 2147 1216
rect 2173 1104 2179 1116
rect 2221 1104 2227 1296
rect 2237 1104 2243 1236
rect 2269 1224 2275 1336
rect 2285 1324 2291 1336
rect 2381 1304 2387 1336
rect 2477 1324 2483 1636
rect 2525 1524 2531 1736
rect 2717 1704 2723 1718
rect 2957 1664 2963 1718
rect 2989 1704 2995 1876
rect 3053 1684 3059 2116
rect 3213 2083 3219 2116
rect 3213 2077 3228 2083
rect 3261 1984 3267 2216
rect 3293 2184 3299 2236
rect 3293 2124 3299 2136
rect 3357 2126 3363 2156
rect 3389 2124 3395 2236
rect 3453 2124 3459 2236
rect 3885 2184 3891 2294
rect 4045 2284 4051 2296
rect 4349 2303 4355 2577
rect 4397 2544 4403 2596
rect 4413 2584 4419 2677
rect 4445 2644 4451 2696
rect 4605 2684 4611 2696
rect 4397 2384 4403 2436
rect 4413 2344 4419 2516
rect 4429 2504 4435 2556
rect 4493 2464 4499 2676
rect 4525 2524 4531 2596
rect 4573 2584 4579 2636
rect 4589 2604 4595 2676
rect 4637 2584 4643 2716
rect 4669 2684 4675 2936
rect 4845 2744 4851 2936
rect 4941 2924 4947 2936
rect 4589 2523 4595 2556
rect 4685 2544 4691 2556
rect 4589 2517 4604 2523
rect 4509 2484 4515 2516
rect 4557 2484 4563 2516
rect 4605 2484 4611 2516
rect 4525 2464 4531 2476
rect 4440 2406 4446 2414
rect 4454 2406 4460 2414
rect 4468 2406 4474 2414
rect 4482 2406 4488 2414
rect 4509 2384 4515 2416
rect 4557 2404 4563 2476
rect 4621 2364 4627 2536
rect 4653 2384 4659 2536
rect 4701 2503 4707 2694
rect 4701 2497 4723 2503
rect 4349 2297 4364 2303
rect 4077 2184 4083 2294
rect 4141 2223 4147 2296
rect 4365 2264 4371 2296
rect 4141 2217 4163 2223
rect 3652 2177 3667 2183
rect 3661 2164 3667 2177
rect 3661 2144 3667 2156
rect 3709 2124 3715 2176
rect 4157 2144 4163 2217
rect 4413 2184 4419 2336
rect 4669 2324 4675 2396
rect 4429 2304 4435 2316
rect 4445 2264 4451 2316
rect 4525 2304 4531 2316
rect 4429 2164 4435 2196
rect 3517 1984 3523 2118
rect 3213 1924 3219 1936
rect 3101 1864 3107 1876
rect 3133 1864 3139 1876
rect 3101 1704 3107 1856
rect 3149 1844 3155 1896
rect 3156 1837 3171 1843
rect 3133 1744 3139 1776
rect 3165 1724 3171 1837
rect 3181 1704 3187 1876
rect 3229 1864 3235 1876
rect 3213 1764 3219 1836
rect 3261 1784 3267 1796
rect 3325 1764 3331 1856
rect 3357 1844 3363 1896
rect 3197 1704 3203 1716
rect 3213 1704 3219 1736
rect 2557 1504 2563 1516
rect 2509 1364 2515 1436
rect 2557 1364 2563 1496
rect 2701 1483 2707 1496
rect 2717 1484 2723 1516
rect 2989 1502 2995 1536
rect 3053 1504 3059 1676
rect 2685 1477 2707 1483
rect 2589 1464 2595 1476
rect 2589 1444 2595 1456
rect 2653 1444 2659 1476
rect 2589 1364 2595 1436
rect 2493 1357 2508 1363
rect 2493 1324 2499 1357
rect 2557 1344 2563 1356
rect 1949 904 1955 916
rect 1901 784 1907 816
rect 1949 784 1955 896
rect 1869 717 1891 723
rect 1764 697 1779 703
rect 1837 644 1843 696
rect 1869 684 1875 717
rect 1885 684 1891 696
rect 1869 664 1875 676
rect 1917 644 1923 716
rect 1981 703 1987 916
rect 2013 904 2019 936
rect 2029 924 2035 936
rect 2061 924 2067 1036
rect 2125 924 2131 996
rect 2157 904 2163 1056
rect 2189 1044 2195 1076
rect 2205 1024 2211 1096
rect 2205 1004 2211 1016
rect 2029 884 2035 896
rect 1997 784 2003 836
rect 1981 697 1996 703
rect 1965 664 1971 676
rect 1981 664 1987 676
rect 1661 544 1667 596
rect 1789 544 1795 616
rect 1725 484 1731 516
rect 1517 284 1523 356
rect 1533 284 1539 416
rect 1565 324 1571 456
rect 1581 384 1587 436
rect 1581 303 1587 336
rect 1645 324 1651 376
rect 1565 297 1587 303
rect 1421 224 1427 276
rect 1533 264 1539 276
rect 1485 184 1491 236
rect 1405 144 1411 176
rect 1549 164 1555 236
rect 1565 184 1571 297
rect 1645 283 1651 316
rect 1645 277 1660 283
rect 1597 224 1603 236
rect 1613 164 1619 276
rect 1661 163 1667 276
rect 1725 224 1731 296
rect 1741 284 1747 456
rect 1757 304 1763 396
rect 1661 157 1676 163
rect 1517 144 1523 156
rect 1613 144 1619 156
rect 1725 144 1731 216
rect 1773 204 1779 436
rect 1837 404 1843 636
rect 1965 584 1971 636
rect 1997 563 2003 696
rect 2029 684 2035 716
rect 2061 704 2067 836
rect 2141 703 2147 836
rect 2173 824 2179 936
rect 2189 924 2195 976
rect 2189 704 2195 856
rect 2205 744 2211 936
rect 2221 903 2227 1096
rect 2269 1084 2275 1176
rect 2285 1104 2291 1176
rect 2340 1117 2355 1123
rect 2301 1064 2307 1116
rect 2349 1104 2355 1117
rect 2429 1104 2435 1116
rect 2445 1104 2451 1316
rect 2461 1284 2467 1316
rect 2509 1224 2515 1336
rect 2653 1324 2659 1336
rect 2685 1324 2691 1477
rect 2701 1344 2707 1456
rect 2525 1304 2531 1316
rect 2525 1184 2531 1276
rect 2653 1184 2659 1236
rect 2653 1124 2659 1176
rect 2333 1084 2339 1096
rect 2237 984 2243 1056
rect 2333 984 2339 1076
rect 2349 1044 2355 1076
rect 2397 1064 2403 1076
rect 2301 944 2307 976
rect 2333 924 2339 956
rect 2413 944 2419 1096
rect 2429 964 2435 1036
rect 2445 924 2451 1096
rect 2461 964 2467 1076
rect 2573 1044 2579 1056
rect 2605 1024 2611 1116
rect 2653 1024 2659 1036
rect 2701 984 2707 1216
rect 2733 1164 2739 1476
rect 2749 1464 2755 1496
rect 2765 1384 2771 1476
rect 2781 1424 2787 1476
rect 2877 1444 2883 1476
rect 2749 1224 2755 1296
rect 2765 1204 2771 1296
rect 2733 1123 2739 1156
rect 2733 1117 2748 1123
rect 2781 1104 2787 1116
rect 2797 1104 2803 1436
rect 2904 1406 2910 1414
rect 2918 1406 2924 1414
rect 2932 1406 2938 1414
rect 2946 1406 2952 1414
rect 2813 1364 2819 1376
rect 2957 1344 2963 1356
rect 3085 1344 3091 1536
rect 3117 1424 3123 1436
rect 3149 1344 3155 1476
rect 3197 1463 3203 1696
rect 3309 1684 3315 1736
rect 3325 1704 3331 1756
rect 3373 1724 3379 1736
rect 3389 1723 3395 1916
rect 3437 1864 3443 1916
rect 3581 1884 3587 2116
rect 3741 1984 3747 2096
rect 3821 2083 3827 2136
rect 3805 2077 3827 2083
rect 3805 1984 3811 2077
rect 3933 1984 3939 2136
rect 3965 2084 3971 2096
rect 4013 1984 4019 2136
rect 4029 1984 4035 2136
rect 4125 2124 4131 2136
rect 3933 1904 3939 1976
rect 3949 1897 3964 1903
rect 3380 1717 3395 1723
rect 3421 1704 3427 1736
rect 3437 1724 3443 1796
rect 3453 1764 3459 1876
rect 3517 1784 3523 1836
rect 3613 1804 3619 1894
rect 3725 1784 3731 1896
rect 3741 1804 3747 1836
rect 3789 1784 3795 1856
rect 3837 1784 3843 1896
rect 3853 1884 3859 1896
rect 3885 1884 3891 1896
rect 3901 1784 3907 1876
rect 3565 1744 3571 1756
rect 3613 1724 3619 1736
rect 3645 1724 3651 1756
rect 3485 1704 3491 1716
rect 3469 1684 3475 1696
rect 3613 1684 3619 1696
rect 3565 1584 3571 1656
rect 3181 1457 3203 1463
rect 2820 1337 2835 1343
rect 2461 924 2467 956
rect 2685 944 2691 976
rect 2429 917 2444 923
rect 2221 897 2236 903
rect 2221 784 2227 876
rect 2253 844 2259 896
rect 2269 704 2275 916
rect 2349 904 2355 916
rect 2132 697 2147 703
rect 2029 584 2035 676
rect 2125 644 2131 676
rect 2237 664 2243 676
rect 2221 657 2236 663
rect 2141 623 2147 656
rect 2205 644 2211 656
rect 2125 617 2147 623
rect 2061 584 2067 616
rect 1981 557 2003 563
rect 1981 544 1987 557
rect 2125 544 2131 617
rect 2221 584 2227 657
rect 2285 663 2291 676
rect 2260 657 2291 663
rect 2269 584 2275 636
rect 2349 583 2355 896
rect 2397 844 2403 896
rect 2397 703 2403 836
rect 2397 697 2412 703
rect 2340 577 2355 583
rect 2157 544 2163 576
rect 1933 384 1939 476
rect 1956 437 1971 443
rect 1789 224 1795 316
rect 1965 304 1971 437
rect 1981 424 1987 536
rect 1997 464 2003 536
rect 2173 524 2179 536
rect 2109 464 2115 496
rect 1981 284 1987 296
rect 1997 284 2003 316
rect 2045 284 2051 316
rect 2061 284 2067 296
rect 1821 264 1827 276
rect 1853 224 1859 276
rect 1741 124 1747 176
rect 1773 123 1779 196
rect 1789 124 1795 216
rect 1869 184 1875 276
rect 1965 264 1971 276
rect 1885 184 1891 196
rect 1917 144 1923 176
rect 1933 144 1939 216
rect 1997 163 2003 176
rect 1981 157 2003 163
rect 1949 124 1955 156
rect 1764 117 1779 123
rect 1981 104 1987 157
rect 1997 124 2003 136
rect 2013 84 2019 236
rect 2029 204 2035 256
rect 2061 104 2067 116
rect 2077 103 2083 456
rect 2173 364 2179 516
rect 2189 384 2195 436
rect 2189 343 2195 356
rect 2173 337 2195 343
rect 2109 304 2115 316
rect 2093 244 2099 256
rect 2109 184 2115 236
rect 2157 184 2163 316
rect 2173 264 2179 337
rect 2189 264 2195 296
rect 2205 284 2211 536
rect 2301 524 2307 556
rect 2333 524 2339 576
rect 2349 524 2355 536
rect 2365 504 2371 656
rect 2429 584 2435 917
rect 2493 864 2499 916
rect 2541 904 2547 916
rect 2573 884 2579 936
rect 2445 644 2451 716
rect 2477 644 2483 716
rect 2509 704 2515 716
rect 2589 704 2595 716
rect 2701 704 2707 736
rect 2717 724 2723 1076
rect 2749 964 2755 1096
rect 2765 944 2771 1076
rect 2813 1064 2819 1116
rect 2829 1104 2835 1337
rect 2845 1324 2851 1336
rect 2829 1044 2835 1076
rect 2925 1044 2931 1076
rect 2877 984 2883 1016
rect 2904 1006 2910 1014
rect 2918 1006 2924 1014
rect 2932 1006 2938 1014
rect 2946 1006 2952 1014
rect 2829 924 2835 956
rect 2973 944 2979 1096
rect 2989 1084 2995 1316
rect 3117 1284 3123 1318
rect 3069 1184 3075 1256
rect 2989 944 2995 1076
rect 3005 964 3011 1036
rect 3037 964 3043 976
rect 2829 884 2835 896
rect 2765 784 2771 876
rect 2861 784 2867 936
rect 2925 904 2931 936
rect 3021 904 3027 916
rect 2541 684 2547 696
rect 2685 684 2691 696
rect 2557 664 2563 676
rect 2621 644 2627 656
rect 2477 584 2483 636
rect 2397 504 2403 576
rect 2413 544 2419 556
rect 2589 544 2595 636
rect 2669 584 2675 676
rect 2733 644 2739 716
rect 2861 704 2867 716
rect 2877 704 2883 736
rect 3037 704 3043 956
rect 3101 904 3107 1216
rect 3133 1102 3139 1236
rect 3149 1084 3155 1336
rect 3181 1324 3187 1457
rect 3245 1384 3251 1556
rect 3645 1544 3651 1716
rect 3693 1684 3699 1756
rect 3741 1744 3747 1776
rect 3773 1744 3779 1756
rect 3677 1677 3692 1683
rect 3677 1524 3683 1677
rect 3325 1484 3331 1516
rect 3469 1464 3475 1476
rect 3309 1444 3315 1456
rect 3261 1344 3267 1416
rect 3373 1344 3379 1456
rect 3437 1384 3443 1436
rect 3485 1424 3491 1496
rect 3517 1424 3523 1516
rect 3549 1350 3555 1476
rect 3565 1444 3571 1496
rect 3629 1464 3635 1476
rect 3581 1364 3587 1456
rect 3581 1344 3587 1356
rect 3613 1344 3619 1456
rect 3453 1184 3459 1276
rect 3485 1184 3491 1336
rect 3565 1184 3571 1276
rect 3325 1102 3331 1136
rect 3501 1097 3516 1103
rect 3261 1024 3267 1036
rect 3165 904 3171 918
rect 3501 924 3507 1097
rect 3565 964 3571 1016
rect 3581 944 3587 1316
rect 3629 1144 3635 1416
rect 3645 1384 3651 1496
rect 3693 1484 3699 1536
rect 3709 1504 3715 1556
rect 3725 1484 3731 1736
rect 3741 1704 3747 1736
rect 3821 1724 3827 1736
rect 3869 1724 3875 1736
rect 3741 1544 3747 1696
rect 3757 1664 3763 1716
rect 3805 1704 3811 1716
rect 3885 1704 3891 1716
rect 3917 1704 3923 1816
rect 3949 1784 3955 1897
rect 3997 1824 4003 1856
rect 4013 1784 4019 1856
rect 4045 1784 4051 1856
rect 3933 1704 3939 1756
rect 3965 1744 3971 1756
rect 4061 1744 4067 1876
rect 4077 1763 4083 1856
rect 4077 1757 4092 1763
rect 4061 1724 4067 1736
rect 4013 1704 4019 1716
rect 3757 1584 3763 1656
rect 3757 1504 3763 1556
rect 3773 1443 3779 1676
rect 3805 1564 3811 1696
rect 3853 1684 3859 1696
rect 3917 1684 3923 1696
rect 3981 1604 3987 1636
rect 3805 1524 3811 1536
rect 3821 1464 3827 1516
rect 3885 1504 3891 1516
rect 3981 1504 3987 1576
rect 3853 1444 3859 1496
rect 3757 1437 3779 1443
rect 3645 1304 3651 1376
rect 3693 1364 3699 1376
rect 3677 1304 3683 1336
rect 3677 1104 3683 1116
rect 3741 984 3747 1396
rect 3757 1344 3763 1437
rect 3805 1384 3811 1436
rect 3837 1304 3843 1376
rect 3853 1324 3859 1336
rect 3805 1104 3811 1176
rect 3821 1124 3827 1236
rect 3789 1064 3795 1096
rect 3661 944 3667 976
rect 3789 964 3795 1016
rect 3357 884 3363 918
rect 3501 883 3507 916
rect 3773 884 3779 936
rect 3492 877 3507 883
rect 3085 724 3091 836
rect 3293 744 3299 836
rect 2836 697 2851 703
rect 2525 444 2531 516
rect 2557 504 2563 536
rect 2541 384 2547 396
rect 2324 317 2339 323
rect 2173 224 2179 236
rect 2189 164 2195 256
rect 2301 244 2307 276
rect 2125 144 2131 156
rect 2205 117 2236 123
rect 2068 97 2083 103
rect 2093 84 2099 116
rect 2205 104 2211 117
rect 2253 84 2259 176
rect 2317 164 2323 236
rect 2333 224 2339 317
rect 2349 284 2355 316
rect 2397 224 2403 296
rect 2429 284 2435 336
rect 2461 284 2467 316
rect 2477 304 2483 376
rect 2509 337 2595 343
rect 2509 324 2515 337
rect 2589 324 2595 337
rect 2452 237 2467 243
rect 2461 223 2467 237
rect 2541 224 2547 276
rect 2461 217 2515 223
rect 2445 184 2451 216
rect 2493 144 2499 196
rect 2509 183 2515 217
rect 2509 177 2540 183
rect 77 64 83 76
rect 2333 64 2339 136
rect 2429 84 2435 136
rect 2445 104 2451 136
rect 2461 123 2467 136
rect 2557 124 2563 276
rect 2461 117 2476 123
rect 2573 103 2579 236
rect 2605 144 2611 576
rect 2733 524 2739 596
rect 2765 564 2771 696
rect 2804 677 2819 683
rect 2797 584 2803 656
rect 2813 604 2819 677
rect 2845 664 2851 697
rect 3069 703 3075 716
rect 3069 697 3084 703
rect 2964 677 3011 683
rect 2781 544 2787 576
rect 2829 564 2835 656
rect 2845 584 2851 656
rect 2909 643 2915 676
rect 2964 657 2979 663
rect 2877 637 2915 643
rect 2861 564 2867 636
rect 2877 604 2883 637
rect 2904 606 2910 614
rect 2918 606 2924 614
rect 2932 606 2938 614
rect 2946 606 2952 614
rect 2973 584 2979 657
rect 3005 623 3011 677
rect 3021 644 3027 696
rect 3037 664 3043 676
rect 3101 644 3107 696
rect 3165 664 3171 736
rect 3213 664 3219 676
rect 3245 644 3251 696
rect 3037 623 3043 636
rect 3005 617 3043 623
rect 3053 563 3059 636
rect 3245 584 3251 636
rect 3261 564 3267 636
rect 3037 557 3059 563
rect 2829 544 2835 556
rect 3037 544 3043 557
rect 2781 504 2787 516
rect 2653 444 2659 476
rect 2621 344 2627 436
rect 2669 384 2675 436
rect 2685 384 2691 476
rect 2781 464 2787 496
rect 2621 304 2627 316
rect 2685 304 2691 356
rect 2749 323 2755 436
rect 2877 384 2883 416
rect 2941 344 2947 516
rect 3005 384 3011 536
rect 3069 523 3075 556
rect 3060 517 3075 523
rect 2845 324 2851 336
rect 2740 317 2755 323
rect 2733 304 2739 316
rect 2861 304 2867 316
rect 2957 304 2963 316
rect 2653 244 2659 276
rect 2765 244 2771 296
rect 2781 264 2787 276
rect 2637 104 2643 156
rect 2653 144 2659 196
rect 2813 184 2819 296
rect 2877 184 2883 296
rect 2904 206 2910 214
rect 2918 206 2924 214
rect 2932 206 2938 214
rect 2946 206 2952 214
rect 2973 164 2979 276
rect 2749 144 2755 156
rect 2765 144 2771 156
rect 2973 144 2979 156
rect 2989 144 2995 336
rect 3005 244 3011 296
rect 3021 284 3027 316
rect 3037 264 3043 376
rect 3085 304 3091 476
rect 3117 304 3123 556
rect 3133 464 3139 516
rect 3181 424 3187 536
rect 3197 503 3203 516
rect 3197 497 3219 503
rect 3133 324 3139 336
rect 3108 297 3116 303
rect 3165 303 3171 396
rect 3181 384 3187 396
rect 3213 384 3219 497
rect 3261 384 3267 536
rect 3293 524 3299 696
rect 3453 684 3459 876
rect 3677 702 3683 716
rect 3325 564 3331 676
rect 3341 524 3347 636
rect 3389 564 3395 636
rect 3421 604 3427 676
rect 3485 624 3491 694
rect 3805 684 3811 1096
rect 3821 1004 3827 1036
rect 3821 924 3827 996
rect 3853 964 3859 1316
rect 3869 1104 3875 1356
rect 3885 1344 3891 1356
rect 3917 1263 3923 1496
rect 4029 1484 4035 1596
rect 4045 1544 4051 1636
rect 4061 1504 4067 1676
rect 4093 1504 4099 1756
rect 4109 1744 4115 2076
rect 4109 1724 4115 1736
rect 4125 1703 4131 1716
rect 4109 1697 4131 1703
rect 4068 1497 4083 1503
rect 4045 1483 4051 1496
rect 4045 1477 4067 1483
rect 3933 1384 3939 1476
rect 3997 1364 4003 1436
rect 4013 1384 4019 1436
rect 3981 1344 3987 1356
rect 4045 1344 4051 1376
rect 4061 1324 4067 1477
rect 4077 1324 4083 1497
rect 4109 1484 4115 1697
rect 4141 1504 4147 1796
rect 4157 1784 4163 2116
rect 4189 2104 4195 2118
rect 4205 1844 4211 1896
rect 4253 1884 4259 2116
rect 4365 2044 4371 2136
rect 4381 1904 4387 2156
rect 4445 2104 4451 2256
rect 4493 2144 4499 2296
rect 4548 2257 4563 2263
rect 4493 2043 4499 2136
rect 4525 2104 4531 2196
rect 4557 2184 4563 2257
rect 4589 2204 4595 2256
rect 4493 2037 4515 2043
rect 4253 1824 4259 1876
rect 4173 1584 4179 1696
rect 4189 1584 4195 1736
rect 4205 1724 4211 1736
rect 4205 1564 4211 1716
rect 4157 1504 4163 1516
rect 4109 1384 4115 1436
rect 4141 1424 4147 1496
rect 4205 1464 4211 1496
rect 4269 1404 4275 1718
rect 4285 1444 4291 1456
rect 4301 1384 4307 1896
rect 4333 1744 4339 1856
rect 4317 1704 4323 1716
rect 4333 1444 4339 1456
rect 3933 1284 3939 1296
rect 3917 1257 3939 1263
rect 3885 1084 3891 1136
rect 3933 1124 3939 1257
rect 3949 1124 3955 1136
rect 3933 984 3939 1116
rect 3965 1084 3971 1276
rect 4061 1204 4067 1316
rect 4077 1284 4083 1316
rect 3949 984 3955 1036
rect 3981 1024 3987 1076
rect 3997 1064 4003 1196
rect 4141 1164 4147 1316
rect 4157 1304 4163 1316
rect 4173 1184 4179 1316
rect 4189 1264 4195 1356
rect 4301 1324 4307 1336
rect 4317 1304 4323 1416
rect 4333 1344 4339 1436
rect 4196 1257 4211 1263
rect 4061 1104 4067 1136
rect 3821 884 3827 896
rect 3837 784 3843 936
rect 3853 904 3859 916
rect 3885 904 3891 976
rect 3901 944 3907 956
rect 3917 924 3923 936
rect 3949 884 3955 956
rect 3965 944 3971 1016
rect 3997 943 4003 1056
rect 3988 937 4003 943
rect 3981 924 3987 936
rect 4013 884 4019 1036
rect 4061 1024 4067 1056
rect 4077 984 4083 1116
rect 4141 1084 4147 1116
rect 4173 1104 4179 1156
rect 4205 1084 4211 1257
rect 4317 1184 4323 1296
rect 4349 1284 4355 1316
rect 4365 1284 4371 1436
rect 4381 1404 4387 1896
rect 4397 1784 4403 2036
rect 4440 2006 4446 2014
rect 4454 2006 4460 2014
rect 4468 2006 4474 2014
rect 4482 2006 4488 2014
rect 4509 1984 4515 2037
rect 4525 1924 4531 2096
rect 4525 1884 4531 1896
rect 4541 1884 4547 1896
rect 4573 1864 4579 2136
rect 4589 2124 4595 2136
rect 4605 2124 4611 2236
rect 4621 1904 4627 1996
rect 4637 1884 4643 2096
rect 4653 2044 4659 2096
rect 4669 2084 4675 2276
rect 4685 2144 4691 2456
rect 4701 2304 4707 2316
rect 4701 2204 4707 2236
rect 4669 2064 4675 2076
rect 4685 2004 4691 2136
rect 4701 2044 4707 2116
rect 4717 1984 4723 2497
rect 4749 2424 4755 2516
rect 4797 2503 4803 2736
rect 4829 2724 4835 2736
rect 4893 2702 4899 2716
rect 4813 2544 4819 2596
rect 4877 2544 4883 2616
rect 4909 2584 4915 2916
rect 4957 2724 4963 2936
rect 5117 2704 5123 2936
rect 5149 2884 5155 2918
rect 5213 2724 5219 2736
rect 4788 2497 4803 2503
rect 4829 2444 4835 2496
rect 4733 2244 4739 2296
rect 4749 2224 4755 2276
rect 4765 2264 4771 2336
rect 4861 2324 4867 2336
rect 4925 2284 4931 2676
rect 5021 2624 5027 2636
rect 4941 2564 4947 2596
rect 5101 2584 5107 2696
rect 5117 2684 5123 2696
rect 5213 2584 5219 2696
rect 5245 2684 5251 2876
rect 5277 2702 5283 2716
rect 5293 2584 5299 2836
rect 5325 2584 5331 3036
rect 5373 2964 5379 3056
rect 5501 3044 5507 3094
rect 5517 2964 5523 3076
rect 5517 2704 5523 2956
rect 5613 2784 5619 3316
rect 5629 3124 5635 3136
rect 5693 3102 5699 3116
rect 5741 2964 5747 3316
rect 5773 3284 5779 3296
rect 5789 2964 5795 3056
rect 5693 2944 5699 2956
rect 5725 2904 5731 2936
rect 5805 2884 5811 2916
rect 5853 2884 5859 2896
rect 5796 2737 5811 2743
rect 5597 2724 5603 2736
rect 5661 2702 5667 2716
rect 5805 2704 5811 2737
rect 5853 2684 5859 2696
rect 5437 2544 5443 2676
rect 5149 2524 5155 2536
rect 4957 2302 4963 2316
rect 4973 2304 4979 2516
rect 4989 2344 4995 2516
rect 4797 2264 4803 2276
rect 4893 2244 4899 2276
rect 5021 2264 5027 2516
rect 5085 2324 5091 2336
rect 5149 2302 5155 2316
rect 4765 2144 4771 2156
rect 4781 2124 4787 2236
rect 4861 2184 4867 2236
rect 4909 2144 4915 2156
rect 4749 2104 4755 2116
rect 4829 2104 4835 2116
rect 4749 2084 4755 2096
rect 4749 1884 4755 2036
rect 4605 1864 4611 1876
rect 4653 1864 4659 1876
rect 4765 1864 4771 1876
rect 4573 1804 4579 1856
rect 4781 1843 4787 1896
rect 4765 1837 4787 1843
rect 4589 1744 4595 1816
rect 4749 1784 4755 1836
rect 4765 1804 4771 1837
rect 4765 1784 4771 1796
rect 4797 1744 4803 2076
rect 4813 2064 4819 2096
rect 4813 2004 4819 2056
rect 4861 1884 4867 1996
rect 4893 1917 4908 1923
rect 4845 1844 4851 1856
rect 4893 1844 4899 1917
rect 4925 1884 4931 1896
rect 4941 1884 4947 2196
rect 4957 2184 4963 2256
rect 4973 2144 4979 2216
rect 5101 2184 5107 2236
rect 5213 2184 5219 2296
rect 5245 2244 5251 2536
rect 5284 2337 5299 2343
rect 5293 2304 5299 2337
rect 4989 2144 4995 2156
rect 5245 2144 5251 2156
rect 4957 2124 4963 2136
rect 4973 1984 4979 2116
rect 4989 2004 4995 2136
rect 5021 2104 5027 2136
rect 5021 2084 5027 2096
rect 5053 1984 5059 2076
rect 5149 1924 5155 2136
rect 5277 2124 5283 2136
rect 4973 1864 4979 1876
rect 4861 1784 4867 1816
rect 4893 1744 4899 1836
rect 4925 1784 4931 1836
rect 4941 1744 4947 1856
rect 4989 1824 4995 1876
rect 4440 1606 4446 1614
rect 4454 1606 4460 1614
rect 4468 1606 4474 1614
rect 4482 1606 4488 1614
rect 4557 1584 4563 1736
rect 4685 1643 4691 1716
rect 4685 1637 4707 1643
rect 4397 1504 4403 1536
rect 4509 1504 4515 1516
rect 4445 1464 4451 1476
rect 4445 1384 4451 1456
rect 4493 1384 4499 1456
rect 4557 1424 4563 1456
rect 4493 1364 4499 1376
rect 4317 1164 4323 1176
rect 4333 1084 4339 1196
rect 4381 1104 4387 1336
rect 4440 1206 4446 1214
rect 4454 1206 4460 1214
rect 4468 1206 4474 1214
rect 4482 1206 4488 1214
rect 4109 984 4115 1076
rect 4029 904 4035 936
rect 4077 904 4083 916
rect 4093 904 4099 956
rect 4141 904 4147 936
rect 4173 924 4179 1036
rect 4189 944 4195 1076
rect 4301 1064 4307 1076
rect 4237 944 4243 976
rect 4269 944 4275 956
rect 4333 944 4339 1076
rect 4189 904 4195 936
rect 3917 784 3923 876
rect 3389 524 3395 536
rect 3405 524 3411 536
rect 3485 524 3491 556
rect 3533 544 3539 676
rect 3693 564 3699 576
rect 3725 544 3731 676
rect 3805 604 3811 636
rect 3277 484 3283 516
rect 3293 404 3299 516
rect 3309 344 3315 516
rect 3501 504 3507 536
rect 3757 526 3763 576
rect 3853 564 3859 716
rect 3901 564 3907 596
rect 3949 584 3955 696
rect 3965 684 3971 716
rect 3997 704 4003 716
rect 4077 704 4083 896
rect 4013 604 4019 676
rect 3965 544 3971 556
rect 4093 544 4099 816
rect 4109 704 4115 716
rect 4125 704 4131 876
rect 4237 784 4243 936
rect 4285 784 4291 916
rect 4333 824 4339 936
rect 4365 884 4371 918
rect 4141 724 4147 756
rect 4237 684 4243 736
rect 4269 724 4275 776
rect 4381 744 4387 1096
rect 4509 984 4515 1396
rect 4621 1384 4627 1416
rect 4525 1004 4531 1356
rect 4573 1324 4579 1336
rect 4573 1184 4579 1316
rect 4589 1124 4595 1316
rect 4637 1304 4643 1556
rect 4701 1484 4707 1637
rect 4749 1384 4755 1476
rect 4797 1384 4803 1736
rect 4909 1584 4915 1736
rect 4669 1344 4675 1356
rect 4909 1344 4915 1576
rect 5021 1524 5027 1756
rect 5037 1724 5043 1796
rect 5085 1784 5091 1816
rect 5069 1744 5075 1776
rect 5101 1764 5107 1856
rect 5165 1844 5171 1896
rect 5149 1764 5155 1836
rect 5181 1764 5187 1836
rect 5197 1784 5203 1916
rect 5213 1884 5219 2116
rect 5245 1984 5251 2116
rect 5277 1884 5283 1996
rect 5309 1884 5315 2136
rect 5325 1944 5331 2136
rect 5341 2104 5347 2116
rect 5341 1984 5347 2096
rect 5357 1963 5363 2536
rect 5421 2184 5427 2518
rect 5437 2304 5443 2536
rect 5565 2524 5571 2616
rect 5629 2544 5635 2676
rect 5597 2484 5603 2496
rect 5661 2484 5667 2518
rect 5716 2337 5731 2343
rect 5517 2324 5523 2336
rect 5581 2302 5587 2316
rect 5725 2304 5731 2337
rect 5773 2304 5779 2636
rect 5805 2483 5811 2516
rect 5796 2477 5811 2483
rect 5757 2284 5763 2296
rect 5549 2124 5555 2276
rect 5645 2144 5651 2276
rect 5373 1984 5379 2116
rect 5485 2084 5491 2118
rect 5341 1957 5363 1963
rect 5325 1884 5331 1936
rect 5053 1704 5059 1736
rect 5117 1724 5123 1756
rect 5140 1737 5155 1743
rect 4989 1344 4995 1476
rect 4685 1324 4691 1336
rect 4637 1184 4643 1296
rect 4733 1144 4739 1296
rect 4589 1104 4595 1116
rect 4621 1084 4627 1096
rect 4589 1004 4595 1076
rect 4621 1064 4627 1076
rect 4669 1044 4675 1096
rect 4797 1084 4803 1156
rect 4621 984 4627 1016
rect 4653 944 4659 956
rect 4669 944 4675 996
rect 4685 984 4691 1076
rect 4781 1064 4787 1076
rect 4797 1004 4803 1076
rect 4781 964 4787 976
rect 4440 806 4446 814
rect 4454 806 4460 814
rect 4468 806 4474 814
rect 4482 806 4488 814
rect 4125 624 4131 676
rect 4125 564 4131 616
rect 4157 584 4163 656
rect 4221 604 4227 656
rect 4157 564 4163 576
rect 3373 484 3379 496
rect 3165 297 3180 303
rect 3005 164 3011 236
rect 3101 204 3107 296
rect 2829 123 2835 136
rect 2820 117 2835 123
rect 2781 104 2787 116
rect 2813 104 2819 116
rect 3021 104 3027 196
rect 3149 184 3155 276
rect 3229 264 3235 316
rect 3309 304 3315 336
rect 3245 264 3251 276
rect 3277 264 3283 296
rect 3101 164 3107 176
rect 3165 164 3171 256
rect 3069 124 3075 156
rect 3085 144 3091 156
rect 3165 144 3171 156
rect 3245 124 3251 196
rect 3325 184 3331 316
rect 3341 304 3347 316
rect 3485 304 3491 476
rect 3501 384 3507 496
rect 3853 484 3859 536
rect 3549 284 3555 376
rect 3565 304 3571 416
rect 3853 304 3859 476
rect 3949 304 3955 476
rect 4029 444 4035 518
rect 4173 484 4179 516
rect 4173 344 4179 476
rect 4189 384 4195 396
rect 4221 324 4227 536
rect 3373 244 3379 276
rect 3469 257 3475 276
rect 3421 244 3427 256
rect 3453 204 3459 236
rect 3565 184 3571 216
rect 3277 144 3283 156
rect 3373 144 3379 176
rect 3757 164 3763 176
rect 3853 144 3859 296
rect 3949 143 3955 296
rect 4157 283 4163 316
rect 4157 277 4172 283
rect 4076 264 4084 270
rect 4109 224 4115 276
rect 4125 264 4131 276
rect 4093 184 4099 196
rect 4029 144 4035 156
rect 4173 144 4179 276
rect 4189 224 4195 296
rect 3949 137 3971 143
rect 3261 124 3267 136
rect 3501 124 3507 136
rect 2532 97 2579 103
rect 2525 84 2531 96
rect 3437 64 3443 118
rect 3693 124 3699 136
rect 3965 124 3971 137
rect 3629 84 3635 118
rect 3949 84 3955 116
rect 4125 104 4131 136
rect 4189 124 4195 216
rect 4237 203 4243 596
rect 4285 556 4291 716
rect 4525 704 4531 936
rect 4685 784 4691 876
rect 4557 684 4563 696
rect 4605 684 4611 736
rect 4765 723 4771 936
rect 4781 924 4787 956
rect 4781 744 4787 916
rect 4829 844 4835 916
rect 4845 864 4851 876
rect 4756 717 4771 723
rect 4749 704 4755 716
rect 4781 684 4787 716
rect 4365 644 4371 656
rect 4349 584 4355 636
rect 4381 564 4387 676
rect 4333 544 4339 556
rect 4253 304 4259 356
rect 4221 197 4243 203
rect 4221 144 4227 197
rect 4221 104 4227 136
rect 4253 123 4259 236
rect 4269 204 4275 296
rect 4301 163 4307 496
rect 4317 324 4323 376
rect 4397 304 4403 576
rect 4413 564 4419 636
rect 4477 464 4483 676
rect 4509 604 4515 676
rect 4509 483 4515 596
rect 4541 584 4547 656
rect 4557 584 4563 676
rect 4525 504 4531 576
rect 4573 564 4579 676
rect 4589 544 4595 676
rect 4621 664 4627 676
rect 4717 664 4723 676
rect 4733 624 4739 676
rect 4797 664 4803 756
rect 4861 703 4867 1116
rect 4893 1024 4899 1094
rect 4909 984 4915 1316
rect 4957 1104 4963 1336
rect 5021 1184 5027 1516
rect 5053 1484 5059 1556
rect 5085 1484 5091 1716
rect 5117 1704 5123 1716
rect 5101 1684 5107 1696
rect 5117 1484 5123 1696
rect 5133 1604 5139 1676
rect 5149 1644 5155 1737
rect 5165 1684 5171 1736
rect 5133 1504 5139 1516
rect 5101 1404 5107 1436
rect 5149 1384 5155 1476
rect 5165 1464 5171 1496
rect 5165 1284 5171 1296
rect 4941 1097 4956 1103
rect 4941 944 4947 1097
rect 5101 1084 5107 1236
rect 5117 1003 5123 1276
rect 5197 1183 5203 1556
rect 5213 1524 5219 1856
rect 5229 1724 5235 1756
rect 5245 1744 5251 1756
rect 5229 1524 5235 1716
rect 5245 1624 5251 1736
rect 5261 1564 5267 1856
rect 5277 1704 5283 1876
rect 5309 1784 5315 1876
rect 5341 1824 5347 1957
rect 5389 1904 5395 1916
rect 5357 1864 5363 1876
rect 5309 1744 5315 1776
rect 5293 1684 5299 1716
rect 5309 1704 5315 1716
rect 5309 1584 5315 1696
rect 5325 1544 5331 1796
rect 5341 1744 5347 1756
rect 5389 1744 5395 1896
rect 5405 1804 5411 1836
rect 5421 1724 5427 1756
rect 5453 1744 5459 1896
rect 5373 1664 5379 1676
rect 5389 1664 5395 1716
rect 5405 1624 5411 1696
rect 5245 1504 5251 1516
rect 5277 1504 5283 1516
rect 5341 1504 5347 1576
rect 5229 1344 5235 1416
rect 5197 1177 5212 1183
rect 5101 997 5123 1003
rect 5101 984 5107 997
rect 5133 983 5139 1176
rect 5245 1143 5251 1436
rect 5341 1384 5347 1476
rect 5357 1464 5363 1496
rect 5229 1137 5251 1143
rect 5124 977 5139 983
rect 5181 924 5187 1136
rect 5229 1084 5235 1137
rect 5277 1104 5283 1336
rect 5373 1304 5379 1616
rect 5421 1464 5427 1516
rect 5437 1504 5443 1736
rect 5501 1724 5507 1896
rect 5677 1884 5683 2136
rect 5693 2084 5699 2116
rect 5821 2083 5827 2116
rect 5853 2084 5859 2096
rect 5812 2077 5827 2083
rect 5533 1764 5539 1856
rect 5565 1764 5571 1776
rect 5453 1664 5459 1716
rect 5453 1503 5459 1656
rect 5469 1524 5475 1636
rect 5485 1584 5491 1716
rect 5533 1624 5539 1716
rect 5453 1497 5475 1503
rect 5405 1384 5411 1456
rect 5389 1344 5395 1356
rect 5389 1284 5395 1336
rect 5405 1244 5411 1296
rect 5293 1124 5299 1236
rect 5325 1084 5331 1236
rect 5453 1144 5459 1436
rect 5341 1084 5347 1136
rect 5469 1084 5475 1497
rect 5485 1424 5491 1496
rect 5517 1484 5523 1596
rect 5533 1424 5539 1616
rect 5597 1584 5603 1836
rect 5661 1724 5667 1816
rect 5677 1723 5683 1876
rect 5837 1824 5843 1836
rect 5677 1717 5692 1723
rect 5693 1484 5699 1716
rect 5773 1683 5779 1716
rect 5853 1684 5859 1696
rect 5764 1677 5779 1683
rect 5709 1504 5715 1636
rect 5501 1344 5507 1356
rect 5565 1344 5571 1376
rect 5661 1344 5667 1396
rect 5709 1384 5715 1476
rect 5773 1344 5779 1356
rect 5485 1244 5491 1336
rect 5549 1283 5555 1316
rect 5540 1277 5555 1283
rect 5597 1104 5603 1236
rect 5677 1184 5683 1336
rect 5789 1283 5795 1316
rect 5789 1277 5804 1283
rect 5629 1124 5635 1136
rect 5693 1102 5699 1116
rect 5549 1084 5555 1096
rect 5293 1024 5299 1036
rect 4909 883 4915 896
rect 4973 884 4979 918
rect 5245 884 5251 918
rect 4909 877 4931 883
rect 4877 704 4883 856
rect 4925 704 4931 877
rect 4941 724 4947 736
rect 5037 704 5043 836
rect 5293 784 5299 876
rect 5181 723 5187 736
rect 5325 724 5331 736
rect 5181 717 5203 723
rect 5197 704 5203 717
rect 5357 704 5363 1036
rect 5373 924 5379 1016
rect 4852 697 4867 703
rect 4605 544 4611 576
rect 4765 564 4771 656
rect 4781 564 4787 616
rect 4797 584 4803 656
rect 4861 583 4867 697
rect 5469 702 5475 1036
rect 5501 984 5507 1076
rect 5549 944 5555 1076
rect 5837 1024 5843 1436
rect 4909 584 4915 696
rect 4932 677 4947 683
rect 4925 584 4931 636
rect 4845 577 4867 583
rect 4701 544 4707 556
rect 4685 524 4691 536
rect 4717 524 4723 536
rect 4573 504 4579 516
rect 4765 504 4771 556
rect 4637 484 4643 496
rect 4509 477 4524 483
rect 4440 406 4446 414
rect 4454 406 4460 414
rect 4468 406 4474 414
rect 4482 406 4488 414
rect 4525 324 4531 476
rect 4589 324 4595 376
rect 4413 317 4428 323
rect 4317 297 4355 303
rect 4317 284 4323 297
rect 4349 263 4355 297
rect 4397 284 4403 296
rect 4413 263 4419 317
rect 4349 257 4419 263
rect 4333 204 4339 256
rect 4445 204 4451 276
rect 4285 157 4307 163
rect 4285 144 4291 157
rect 4253 117 4268 123
rect 4333 104 4339 156
rect 4349 124 4355 196
rect 4381 184 4387 196
rect 4413 164 4419 196
rect 4477 144 4483 316
rect 4493 304 4499 316
rect 4573 224 4579 316
rect 4580 217 4595 223
rect 4525 184 4531 216
rect 4557 184 4563 196
rect 4589 164 4595 217
rect 4605 184 4611 356
rect 4653 324 4659 336
rect 4628 317 4643 323
rect 4621 284 4627 296
rect 4637 284 4643 317
rect 4685 304 4691 496
rect 4845 484 4851 577
rect 4861 524 4867 536
rect 4877 524 4883 536
rect 4893 524 4899 576
rect 4941 564 4947 677
rect 4941 544 4947 556
rect 4909 497 4924 503
rect 4701 323 4707 436
rect 4717 384 4723 396
rect 4765 384 4771 436
rect 4701 317 4723 323
rect 4685 284 4691 296
rect 4717 284 4723 317
rect 4573 144 4579 156
rect 4525 104 4531 136
rect 4621 104 4627 156
rect 4637 144 4643 216
rect 4669 164 4675 236
rect 4749 204 4755 276
rect 4765 264 4771 296
rect 4781 244 4787 296
rect 4797 284 4803 376
rect 4845 304 4851 476
rect 4861 304 4867 376
rect 4813 144 4819 216
rect 4829 204 4835 276
rect 4701 103 4707 136
rect 4692 97 4707 103
rect 4845 103 4851 296
rect 4877 283 4883 356
rect 4868 277 4883 283
rect 4893 144 4899 356
rect 4909 324 4915 497
rect 4909 124 4915 236
rect 4925 164 4931 316
rect 4941 303 4947 396
rect 4957 384 4963 576
rect 4973 564 4979 656
rect 4989 584 4995 656
rect 5005 644 5011 656
rect 5037 564 5043 636
rect 5053 584 5059 676
rect 5021 484 5027 516
rect 4989 324 4995 376
rect 5021 304 5027 316
rect 4941 297 4956 303
rect 5037 284 5043 496
rect 5069 404 5075 696
rect 5101 684 5107 696
rect 5085 564 5091 676
rect 5293 664 5299 696
rect 5101 584 5107 656
rect 5133 563 5139 656
rect 5197 584 5203 656
rect 5421 584 5427 636
rect 5124 557 5139 563
rect 5229 544 5235 576
rect 5501 544 5507 676
rect 5517 584 5523 936
rect 5773 924 5779 1016
rect 5581 884 5587 918
rect 5725 883 5731 916
rect 5757 884 5763 896
rect 5716 877 5731 883
rect 5597 724 5603 736
rect 5661 702 5667 716
rect 5677 684 5683 876
rect 5796 737 5811 743
rect 5805 704 5811 737
rect 5853 684 5859 696
rect 5085 524 5091 536
rect 5501 524 5507 536
rect 5085 364 5091 516
rect 5101 384 5107 476
rect 4973 244 4979 276
rect 5005 243 5011 276
rect 5053 264 5059 296
rect 5069 264 5075 276
rect 5085 243 5091 316
rect 5005 237 5091 243
rect 5005 164 5011 196
rect 5053 184 5059 216
rect 5069 164 5075 196
rect 5117 164 5123 516
rect 5149 244 5155 256
rect 5133 184 5139 196
rect 5165 184 5171 496
rect 5197 304 5203 396
rect 5325 384 5331 516
rect 5181 264 5187 276
rect 5124 137 5164 143
rect 4861 104 4867 116
rect 4845 97 4860 103
rect 4925 103 4931 136
rect 4941 124 4947 136
rect 4957 124 4963 136
rect 5197 124 5203 216
rect 5229 184 5235 296
rect 4989 104 4995 116
rect 5213 104 5219 156
rect 5245 124 5251 256
rect 5261 144 5267 236
rect 5277 224 5283 296
rect 5293 284 5299 336
rect 5389 204 5395 296
rect 5405 284 5411 316
rect 5437 264 5443 296
rect 5501 284 5507 296
rect 5277 124 5283 136
rect 5389 124 5395 196
rect 5421 184 5427 216
rect 5469 164 5475 236
rect 5485 224 5491 276
rect 5517 263 5523 316
rect 5533 283 5539 676
rect 5725 544 5731 676
rect 5565 384 5571 496
rect 5533 277 5548 283
rect 5581 264 5587 436
rect 5693 384 5699 516
rect 5613 264 5619 276
rect 5501 257 5523 263
rect 5501 183 5507 257
rect 5517 184 5523 236
rect 5597 184 5603 196
rect 5645 184 5651 276
rect 5661 224 5667 276
rect 5757 264 5763 276
rect 5773 244 5779 276
rect 5773 184 5779 216
rect 5492 177 5507 183
rect 5437 144 5443 156
rect 5405 124 5411 136
rect 5469 124 5475 136
rect 5485 124 5491 176
rect 5501 124 5507 136
rect 5533 104 5539 156
rect 5709 144 5715 156
rect 5725 144 5731 176
rect 5565 104 5571 116
rect 5613 104 5619 136
rect 5789 124 5795 276
rect 5805 104 5811 276
rect 5821 184 5827 316
rect 4925 97 4956 103
rect 5853 84 5859 96
rect 1352 6 1358 14
rect 1366 6 1372 14
rect 1380 6 1386 14
rect 1394 6 1400 14
rect 4440 6 4446 14
rect 4454 6 4460 14
rect 4468 6 4474 14
rect 4482 6 4488 14
<< m3contact >>
rect 2910 4206 2918 4214
rect 2924 4206 2932 4214
rect 2938 4206 2946 4214
rect 972 4196 980 4204
rect 348 4156 356 4164
rect 396 4156 404 4164
rect 108 4136 116 4144
rect 172 4136 180 4144
rect 284 4136 292 4144
rect 44 4116 52 4124
rect 92 4116 100 4124
rect 204 4116 212 4124
rect 12 4096 20 4104
rect 76 3956 84 3964
rect 28 3936 36 3944
rect 12 3876 20 3884
rect 76 3876 84 3884
rect 108 3876 116 3884
rect 28 3736 36 3744
rect 60 3736 68 3744
rect 60 3716 68 3724
rect 44 3496 52 3504
rect 220 3976 228 3984
rect 220 3916 228 3924
rect 156 3896 164 3904
rect 220 3876 228 3884
rect 444 4136 452 4144
rect 3148 4176 3156 4184
rect 1388 4156 1396 4164
rect 1452 4156 1460 4164
rect 1500 4156 1508 4164
rect 1740 4156 1748 4164
rect 2028 4156 2036 4164
rect 2092 4156 2100 4164
rect 2172 4156 2180 4164
rect 2204 4156 2212 4164
rect 2412 4156 2420 4164
rect 2556 4156 2564 4164
rect 620 4136 628 4144
rect 812 4136 820 4144
rect 844 4136 852 4144
rect 1100 4136 1108 4144
rect 1228 4136 1236 4144
rect 1340 4136 1348 4144
rect 316 4116 324 4124
rect 428 4116 436 4124
rect 588 4118 596 4124
rect 588 4116 596 4118
rect 348 4096 356 4104
rect 780 4096 788 4104
rect 428 4076 436 4084
rect 572 4076 580 4084
rect 652 4076 660 4084
rect 380 4056 388 4064
rect 268 4036 276 4044
rect 380 4036 388 4044
rect 492 3976 500 3984
rect 428 3956 436 3964
rect 332 3936 340 3944
rect 380 3936 388 3944
rect 252 3916 260 3924
rect 156 3836 164 3844
rect 108 3736 116 3744
rect 124 3736 132 3744
rect 140 3676 148 3684
rect 92 3616 100 3624
rect 172 3736 180 3744
rect 412 3916 420 3924
rect 300 3856 308 3864
rect 332 3856 340 3864
rect 364 3856 372 3864
rect 348 3776 356 3784
rect 364 3756 372 3764
rect 316 3736 324 3744
rect 236 3716 244 3724
rect 204 3696 212 3704
rect 220 3656 228 3664
rect 188 3636 196 3644
rect 220 3636 228 3644
rect 204 3616 212 3624
rect 156 3536 164 3544
rect 188 3536 196 3544
rect 172 3496 180 3504
rect 284 3696 292 3704
rect 316 3716 324 3724
rect 300 3636 308 3644
rect 268 3616 276 3624
rect 252 3596 260 3604
rect 284 3516 292 3524
rect 188 3476 196 3484
rect 60 3456 68 3464
rect 76 3456 84 3464
rect 220 3456 228 3464
rect 108 3356 116 3364
rect 76 3236 84 3244
rect 12 3136 20 3144
rect 44 3076 52 3084
rect 188 3416 196 3424
rect 140 3316 148 3324
rect 252 3356 260 3364
rect 268 3356 276 3364
rect 252 3316 260 3324
rect 348 3696 356 3704
rect 364 3696 372 3704
rect 348 3616 356 3624
rect 332 3476 340 3484
rect 380 3656 388 3664
rect 444 3916 452 3924
rect 476 3896 484 3904
rect 540 3956 548 3964
rect 524 3896 532 3904
rect 540 3876 548 3884
rect 620 4056 628 4064
rect 764 3936 772 3944
rect 620 3896 628 3904
rect 636 3876 644 3884
rect 748 3876 756 3884
rect 796 3916 804 3924
rect 828 3876 836 3884
rect 412 3856 420 3864
rect 428 3676 436 3684
rect 396 3616 404 3624
rect 428 3536 436 3544
rect 332 3456 340 3464
rect 364 3436 372 3444
rect 316 3336 324 3344
rect 300 3316 308 3324
rect 284 3296 292 3304
rect 268 3236 276 3244
rect 188 3136 196 3144
rect 204 3136 212 3144
rect 220 3116 228 3124
rect 252 3116 260 3124
rect 316 3136 324 3144
rect 300 3116 308 3124
rect 124 3096 132 3104
rect 204 3096 212 3104
rect 108 3076 116 3084
rect 60 2976 68 2984
rect 60 2956 68 2964
rect 28 2896 36 2904
rect 76 2896 84 2904
rect 172 3076 180 3084
rect 124 3056 132 3064
rect 156 3056 164 3064
rect 204 3056 212 3064
rect 236 3056 244 3064
rect 220 2996 228 3004
rect 124 2956 132 2964
rect 140 2956 148 2964
rect 204 2956 212 2964
rect 76 2856 84 2864
rect 108 2856 116 2864
rect 124 2856 132 2864
rect 108 2836 116 2844
rect 380 3396 388 3404
rect 412 3496 420 3504
rect 476 3736 484 3744
rect 460 3696 468 3704
rect 492 3636 500 3644
rect 476 3616 484 3624
rect 540 3616 548 3624
rect 492 3516 500 3524
rect 460 3476 468 3484
rect 444 3456 452 3464
rect 476 3456 484 3464
rect 428 3436 436 3444
rect 412 3336 420 3344
rect 508 3476 516 3484
rect 652 3736 660 3744
rect 620 3718 628 3724
rect 620 3716 628 3718
rect 684 3696 692 3704
rect 572 3596 580 3604
rect 604 3596 612 3604
rect 636 3536 644 3544
rect 604 3516 612 3524
rect 620 3496 628 3504
rect 652 3516 660 3524
rect 684 3496 692 3504
rect 556 3476 564 3484
rect 620 3476 628 3484
rect 524 3436 532 3444
rect 604 3456 612 3464
rect 540 3396 548 3404
rect 588 3396 596 3404
rect 684 3436 692 3444
rect 364 3296 372 3304
rect 540 3296 548 3304
rect 476 3276 484 3284
rect 524 3276 532 3284
rect 412 3256 420 3264
rect 524 3176 532 3184
rect 412 3136 420 3144
rect 444 3136 452 3144
rect 364 3096 372 3104
rect 492 3096 500 3104
rect 300 3076 308 3084
rect 332 3076 340 3084
rect 284 3056 292 3064
rect 252 2936 260 2944
rect 172 2916 180 2924
rect 236 2916 244 2924
rect 156 2836 164 2844
rect 140 2716 148 2724
rect 188 2776 196 2784
rect 220 2736 228 2744
rect 236 2716 244 2724
rect 172 2696 180 2704
rect 204 2696 212 2704
rect 172 2676 180 2684
rect 60 2636 68 2644
rect 12 2536 20 2544
rect 60 2616 68 2624
rect 108 2576 116 2584
rect 188 2616 196 2624
rect 140 2596 148 2604
rect 12 2236 20 2244
rect 60 2118 68 2124
rect 60 2116 68 2118
rect 204 2576 212 2584
rect 156 2556 164 2564
rect 188 2556 196 2564
rect 220 2556 228 2564
rect 220 2536 228 2544
rect 156 2496 164 2504
rect 348 3056 356 3064
rect 332 3016 340 3024
rect 412 3076 420 3084
rect 508 3076 516 3084
rect 396 3056 404 3064
rect 316 2976 324 2984
rect 364 2976 372 2984
rect 300 2916 308 2924
rect 348 2956 356 2964
rect 364 2936 372 2944
rect 332 2896 340 2904
rect 300 2876 308 2884
rect 284 2736 292 2744
rect 268 2716 276 2724
rect 316 2716 324 2724
rect 268 2696 276 2704
rect 348 2796 356 2804
rect 364 2716 372 2724
rect 348 2696 356 2704
rect 332 2676 340 2684
rect 364 2676 372 2684
rect 444 3016 452 3024
rect 412 2976 420 2984
rect 396 2956 404 2964
rect 460 2996 468 3004
rect 476 2996 484 3004
rect 508 2976 516 2984
rect 508 2956 516 2964
rect 428 2736 436 2744
rect 412 2676 420 2684
rect 540 3136 548 3144
rect 732 3756 740 3764
rect 716 3716 724 3724
rect 764 3716 772 3724
rect 732 3676 740 3684
rect 748 3656 756 3664
rect 764 3656 772 3664
rect 780 3636 788 3644
rect 748 3496 756 3504
rect 780 3476 788 3484
rect 764 3456 772 3464
rect 988 4056 996 4064
rect 860 3916 868 3924
rect 892 3916 900 3924
rect 972 3916 980 3924
rect 924 3896 932 3904
rect 1004 3936 1012 3944
rect 1084 3916 1092 3924
rect 1052 3896 1060 3904
rect 924 3876 932 3884
rect 988 3876 996 3884
rect 1004 3876 1012 3884
rect 1036 3876 1044 3884
rect 1084 3876 1092 3884
rect 844 3736 852 3744
rect 1164 4076 1172 4084
rect 1260 4096 1268 4104
rect 1436 4136 1444 4144
rect 1484 4136 1492 4144
rect 1932 4136 1940 4144
rect 1980 4136 1988 4144
rect 1420 4096 1428 4104
rect 1358 4006 1366 4014
rect 1372 4006 1380 4014
rect 1386 4006 1394 4014
rect 1324 3976 1332 3984
rect 1452 3956 1460 3964
rect 1532 4076 1540 4084
rect 1596 4036 1604 4044
rect 1676 4116 1684 4124
rect 1644 4096 1652 4104
rect 1660 4036 1668 4044
rect 1612 3976 1620 3984
rect 1484 3936 1492 3944
rect 1596 3936 1604 3944
rect 1580 3916 1588 3924
rect 1260 3902 1268 3904
rect 1260 3896 1268 3902
rect 1404 3896 1412 3904
rect 1772 4116 1780 4124
rect 1804 4116 1812 4124
rect 1868 4116 1876 4124
rect 1788 4096 1796 4104
rect 1820 4096 1828 4104
rect 1724 4076 1732 4084
rect 2124 4136 2132 4144
rect 2444 4136 2452 4144
rect 1948 4116 1956 4124
rect 2012 4116 2020 4124
rect 2076 4116 2084 4124
rect 2108 4116 2116 4124
rect 2332 4118 2340 4124
rect 2332 4116 2340 4118
rect 2396 4116 2404 4124
rect 1916 4076 1924 4084
rect 1996 4096 2004 4104
rect 1932 4036 1940 4044
rect 1868 4016 1876 4024
rect 1756 3996 1764 4004
rect 2092 4016 2100 4024
rect 1804 3976 1812 3984
rect 1884 3976 1892 3984
rect 1996 3976 2004 3984
rect 1708 3936 1716 3944
rect 1708 3916 1716 3924
rect 1756 3936 1764 3944
rect 1628 3896 1636 3904
rect 1660 3896 1668 3904
rect 1676 3896 1684 3904
rect 1116 3876 1124 3884
rect 1612 3876 1620 3884
rect 1660 3876 1668 3884
rect 1132 3836 1140 3844
rect 1276 3816 1284 3824
rect 908 3718 916 3724
rect 908 3716 916 3718
rect 940 3716 948 3724
rect 1372 3856 1380 3864
rect 1292 3736 1300 3744
rect 1724 3896 1732 3904
rect 1772 3916 1780 3924
rect 1788 3876 1796 3884
rect 1628 3856 1636 3864
rect 1692 3856 1700 3864
rect 1484 3836 1492 3844
rect 1516 3796 1524 3804
rect 1532 3776 1540 3784
rect 1500 3736 1508 3744
rect 1468 3716 1476 3724
rect 1100 3696 1108 3704
rect 972 3676 980 3684
rect 828 3456 836 3464
rect 796 3416 804 3424
rect 748 3396 756 3404
rect 780 3376 788 3384
rect 812 3376 820 3384
rect 716 3356 724 3364
rect 812 3356 820 3364
rect 700 3316 708 3324
rect 716 3296 724 3304
rect 748 3296 756 3304
rect 652 3276 660 3284
rect 700 3276 708 3284
rect 668 3256 676 3264
rect 684 3156 692 3164
rect 636 3136 644 3144
rect 668 3136 676 3144
rect 652 3036 660 3044
rect 748 3196 756 3204
rect 732 3136 740 3144
rect 716 3116 724 3124
rect 764 3076 772 3084
rect 716 3036 724 3044
rect 684 3016 692 3024
rect 636 2976 644 2984
rect 668 2976 676 2984
rect 620 2956 628 2964
rect 524 2896 532 2904
rect 492 2876 500 2884
rect 476 2756 484 2764
rect 524 2736 532 2744
rect 284 2656 292 2664
rect 412 2656 420 2664
rect 476 2656 484 2664
rect 332 2636 340 2644
rect 268 2556 276 2564
rect 332 2556 340 2564
rect 460 2636 468 2644
rect 492 2636 500 2644
rect 684 2936 692 2944
rect 556 2916 564 2924
rect 572 2916 580 2924
rect 620 2916 628 2924
rect 652 2916 660 2924
rect 604 2856 612 2864
rect 556 2756 564 2764
rect 588 2756 596 2764
rect 700 2856 708 2864
rect 700 2796 708 2804
rect 684 2716 692 2724
rect 844 3316 852 3324
rect 876 3516 884 3524
rect 1164 3656 1172 3664
rect 1132 3516 1140 3524
rect 1308 3636 1316 3644
rect 1404 3636 1412 3644
rect 1358 3606 1366 3614
rect 1372 3606 1380 3614
rect 1386 3606 1394 3614
rect 1836 3956 1844 3964
rect 1852 3956 1860 3964
rect 1756 3756 1764 3764
rect 1788 3756 1796 3764
rect 1804 3756 1812 3764
rect 1948 3916 1956 3924
rect 2044 3916 2052 3924
rect 1884 3896 1892 3904
rect 1964 3896 1972 3904
rect 1900 3876 1908 3884
rect 2028 3876 2036 3884
rect 1868 3856 1876 3864
rect 1900 3856 1908 3864
rect 1964 3856 1972 3864
rect 1836 3716 1844 3724
rect 1628 3696 1636 3704
rect 1724 3676 1732 3684
rect 1868 3696 1876 3704
rect 1916 3756 1924 3764
rect 1948 3756 1956 3764
rect 1964 3736 1972 3744
rect 1996 3736 2004 3744
rect 1996 3716 2004 3724
rect 1900 3676 1908 3684
rect 1932 3676 1940 3684
rect 2028 3756 2036 3764
rect 2044 3756 2052 3764
rect 2076 3756 2084 3764
rect 2188 4096 2196 4104
rect 2284 4096 2292 4104
rect 2268 4036 2276 4044
rect 2156 3976 2164 3984
rect 2140 3936 2148 3944
rect 2124 3876 2132 3884
rect 2204 3936 2212 3944
rect 2140 3816 2148 3824
rect 2108 3756 2116 3764
rect 2124 3736 2132 3744
rect 2076 3716 2084 3724
rect 2092 3716 2100 3724
rect 2108 3716 2116 3724
rect 2044 3696 2052 3704
rect 2204 3876 2212 3884
rect 2236 3876 2244 3884
rect 2428 4036 2436 4044
rect 2332 3996 2340 4004
rect 2348 3956 2356 3964
rect 2428 3936 2436 3944
rect 2284 3896 2292 3904
rect 2284 3876 2292 3884
rect 2380 3876 2388 3884
rect 2332 3776 2340 3784
rect 2300 3756 2308 3764
rect 2396 3756 2404 3764
rect 2252 3736 2260 3744
rect 2284 3736 2292 3744
rect 2300 3736 2308 3744
rect 2172 3716 2180 3724
rect 2188 3716 2196 3724
rect 2076 3676 2084 3684
rect 2156 3676 2164 3684
rect 1772 3636 1780 3644
rect 2012 3636 2020 3644
rect 1596 3596 1604 3604
rect 1660 3576 1668 3584
rect 1500 3536 1508 3544
rect 1596 3536 1604 3544
rect 1180 3516 1188 3524
rect 1308 3516 1316 3524
rect 1356 3516 1364 3524
rect 1372 3516 1380 3524
rect 1164 3496 1172 3504
rect 892 3476 900 3484
rect 1020 3476 1028 3484
rect 892 3356 900 3364
rect 892 3336 900 3344
rect 1068 3456 1076 3464
rect 1212 3496 1220 3504
rect 1324 3496 1332 3504
rect 1196 3476 1204 3484
rect 1228 3436 1236 3444
rect 1164 3416 1172 3424
rect 1020 3376 1028 3384
rect 1084 3376 1092 3384
rect 956 3356 964 3364
rect 1020 3356 1028 3364
rect 1036 3356 1044 3364
rect 972 3336 980 3344
rect 1068 3336 1076 3344
rect 892 3316 900 3324
rect 940 3316 948 3324
rect 956 3316 964 3324
rect 812 3256 820 3264
rect 796 3196 804 3204
rect 796 3076 804 3084
rect 844 3076 852 3084
rect 732 2976 740 2984
rect 780 2976 788 2984
rect 748 2956 756 2964
rect 764 2956 772 2964
rect 828 3056 836 3064
rect 844 3056 852 3064
rect 876 3056 884 3064
rect 764 2916 772 2924
rect 780 2916 788 2924
rect 748 2896 756 2904
rect 828 2996 836 3004
rect 1020 3316 1028 3324
rect 1100 3316 1108 3324
rect 908 3156 916 3164
rect 956 3096 964 3104
rect 972 3076 980 3084
rect 1068 3096 1076 3104
rect 1036 3076 1044 3084
rect 924 3056 932 3064
rect 1004 3056 1012 3064
rect 1020 3056 1028 3064
rect 908 3016 916 3024
rect 1020 3036 1028 3044
rect 1052 3056 1060 3064
rect 988 2976 996 2984
rect 1020 2976 1028 2984
rect 1132 3376 1140 3384
rect 1196 3416 1204 3424
rect 1180 3356 1188 3364
rect 1244 3376 1252 3384
rect 1132 3316 1140 3324
rect 1132 3296 1140 3304
rect 1196 3296 1204 3304
rect 1228 3196 1236 3204
rect 1196 3136 1204 3144
rect 1260 3336 1268 3344
rect 1852 3556 1860 3564
rect 1788 3536 1796 3544
rect 1948 3596 1956 3604
rect 1420 3476 1428 3484
rect 1724 3476 1732 3484
rect 1836 3476 1844 3484
rect 1372 3456 1380 3464
rect 1484 3436 1492 3444
rect 1548 3436 1556 3444
rect 1516 3416 1524 3424
rect 1532 3396 1540 3404
rect 1404 3376 1412 3384
rect 1740 3396 1748 3404
rect 1628 3376 1636 3384
rect 1724 3376 1732 3384
rect 1596 3356 1604 3364
rect 1644 3356 1652 3364
rect 2012 3536 2020 3544
rect 2156 3536 2164 3544
rect 1996 3516 2004 3524
rect 2076 3516 2084 3524
rect 1964 3496 1972 3504
rect 2092 3496 2100 3504
rect 2140 3496 2148 3504
rect 1964 3476 1972 3484
rect 2092 3476 2100 3484
rect 1948 3436 1956 3444
rect 2220 3696 2228 3704
rect 2396 3696 2404 3704
rect 2252 3676 2260 3684
rect 2236 3656 2244 3664
rect 2236 3576 2244 3584
rect 3884 4176 3892 4184
rect 3932 4176 3940 4184
rect 2668 4136 2676 4144
rect 2716 4136 2724 4144
rect 2940 4136 2948 4144
rect 3020 4136 3028 4144
rect 3228 4136 3236 4144
rect 3724 4136 3732 4144
rect 3868 4136 3876 4144
rect 2492 4096 2500 4104
rect 2652 4116 2660 4124
rect 2668 4036 2676 4044
rect 2540 4016 2548 4024
rect 2556 4016 2564 4024
rect 2476 3936 2484 3944
rect 2540 3916 2548 3924
rect 2652 3876 2660 3884
rect 2540 3856 2548 3864
rect 2556 3856 2564 3864
rect 2460 3836 2468 3844
rect 2492 3836 2500 3844
rect 2460 3816 2468 3824
rect 2540 3816 2548 3824
rect 2588 3796 2596 3804
rect 2620 3796 2628 3804
rect 2428 3776 2436 3784
rect 2524 3776 2532 3784
rect 2508 3736 2516 3744
rect 2556 3756 2564 3764
rect 2444 3716 2452 3724
rect 2572 3716 2580 3724
rect 2620 3716 2628 3724
rect 2412 3676 2420 3684
rect 2444 3616 2452 3624
rect 2556 3696 2564 3704
rect 2508 3676 2516 3684
rect 2556 3676 2564 3684
rect 2636 3676 2644 3684
rect 2668 3796 2676 3804
rect 2732 4116 2740 4124
rect 2732 3976 2740 3984
rect 2716 3916 2724 3924
rect 2780 4056 2788 4064
rect 3292 4118 3300 4124
rect 3292 4116 3300 4118
rect 3388 4116 3396 4124
rect 3452 4116 3460 4124
rect 3548 4116 3556 4124
rect 3196 4096 3204 4104
rect 3004 4076 3012 4084
rect 3052 3996 3060 4004
rect 2780 3976 2788 3984
rect 3164 3976 3172 3984
rect 2764 3916 2772 3924
rect 2700 3896 2708 3904
rect 2748 3876 2756 3884
rect 2716 3856 2724 3864
rect 2700 3776 2708 3784
rect 2764 3776 2772 3784
rect 2796 3916 2804 3924
rect 3084 3916 3092 3924
rect 3116 3916 3124 3924
rect 3132 3916 3140 3924
rect 2748 3756 2756 3764
rect 2668 3716 2676 3724
rect 2764 3716 2772 3724
rect 2812 3896 2820 3904
rect 2924 3896 2932 3904
rect 2988 3876 2996 3884
rect 2796 3736 2804 3744
rect 2780 3696 2788 3704
rect 2444 3576 2452 3584
rect 2492 3576 2500 3584
rect 2620 3576 2628 3584
rect 2332 3516 2340 3524
rect 2284 3496 2292 3504
rect 2316 3496 2324 3504
rect 2364 3496 2372 3504
rect 2476 3516 2484 3524
rect 2556 3516 2564 3524
rect 2492 3496 2500 3504
rect 2220 3476 2228 3484
rect 2380 3476 2388 3484
rect 2188 3456 2196 3464
rect 2316 3456 2324 3464
rect 2252 3436 2260 3444
rect 2060 3376 2068 3384
rect 2188 3376 2196 3384
rect 2332 3376 2340 3384
rect 2412 3376 2420 3384
rect 2396 3356 2404 3364
rect 1308 3336 1316 3344
rect 1340 3336 1348 3344
rect 1436 3336 1444 3344
rect 1564 3336 1572 3344
rect 1596 3336 1604 3344
rect 1308 3316 1316 3324
rect 1372 3316 1380 3324
rect 1388 3316 1396 3324
rect 1980 3316 1988 3324
rect 1468 3236 1476 3244
rect 1358 3206 1366 3214
rect 1372 3206 1380 3214
rect 1386 3206 1394 3214
rect 1308 3196 1316 3204
rect 1276 3156 1284 3164
rect 1244 3116 1252 3124
rect 1276 3116 1284 3124
rect 1148 2996 1156 3004
rect 1100 2976 1108 2984
rect 1132 2976 1140 2984
rect 860 2936 868 2944
rect 892 2936 900 2944
rect 1020 2936 1028 2944
rect 876 2916 884 2924
rect 908 2916 916 2924
rect 956 2916 964 2924
rect 764 2876 772 2884
rect 812 2876 820 2884
rect 828 2876 836 2884
rect 796 2776 804 2784
rect 652 2696 660 2704
rect 764 2696 772 2704
rect 684 2676 692 2684
rect 556 2656 564 2664
rect 620 2636 628 2644
rect 540 2596 548 2604
rect 508 2556 516 2564
rect 396 2536 404 2544
rect 604 2536 612 2544
rect 620 2536 628 2544
rect 764 2676 772 2684
rect 780 2576 788 2584
rect 732 2536 740 2544
rect 748 2536 756 2544
rect 780 2536 788 2544
rect 316 2516 324 2524
rect 348 2516 356 2524
rect 316 2496 324 2504
rect 412 2496 420 2504
rect 460 2496 468 2504
rect 380 2296 388 2304
rect 412 2296 420 2304
rect 124 2136 132 2144
rect 28 1836 36 1844
rect 268 2156 276 2164
rect 348 2156 356 2164
rect 316 2136 324 2144
rect 396 2036 404 2044
rect 556 2336 564 2344
rect 908 2896 916 2904
rect 956 2756 964 2764
rect 972 2696 980 2704
rect 844 2676 852 2684
rect 988 2676 996 2684
rect 1020 2676 1028 2684
rect 828 2656 836 2664
rect 1004 2656 1012 2664
rect 924 2616 932 2624
rect 908 2576 916 2584
rect 876 2536 884 2544
rect 828 2516 836 2524
rect 1020 2596 1028 2604
rect 940 2556 948 2564
rect 972 2536 980 2544
rect 1020 2536 1028 2544
rect 1052 2936 1060 2944
rect 1084 2936 1092 2944
rect 1132 2936 1140 2944
rect 1372 3136 1380 3144
rect 1436 3116 1444 3124
rect 1516 3116 1524 3124
rect 1532 3116 1540 3124
rect 1724 3236 1732 3244
rect 1996 3236 2004 3244
rect 1324 3096 1332 3104
rect 1340 3096 1348 3104
rect 1500 3096 1508 3104
rect 1308 3076 1316 3084
rect 1452 3076 1460 3084
rect 1180 3036 1188 3044
rect 1212 3036 1220 3044
rect 1276 3036 1284 3044
rect 1196 2956 1204 2964
rect 1196 2936 1204 2944
rect 1228 2936 1236 2944
rect 1292 3016 1300 3024
rect 1372 2976 1380 2984
rect 1308 2956 1316 2964
rect 1324 2956 1332 2964
rect 1164 2876 1172 2884
rect 1084 2856 1092 2864
rect 1324 2896 1332 2904
rect 1324 2876 1332 2884
rect 1292 2856 1300 2864
rect 1116 2836 1124 2844
rect 1164 2836 1172 2844
rect 1228 2836 1236 2844
rect 1084 2796 1092 2804
rect 1068 2696 1076 2704
rect 1052 2536 1060 2544
rect 988 2476 996 2484
rect 1036 2476 1044 2484
rect 844 2336 852 2344
rect 796 2316 804 2324
rect 924 2316 932 2324
rect 812 2276 820 2284
rect 540 2216 548 2224
rect 524 2196 532 2204
rect 652 2216 660 2224
rect 556 2136 564 2144
rect 796 2236 804 2244
rect 972 2216 980 2224
rect 1036 2216 1044 2224
rect 700 2136 708 2144
rect 940 2136 948 2144
rect 972 2136 980 2144
rect 444 2036 452 2044
rect 428 1936 436 1944
rect 428 1916 436 1924
rect 396 1896 404 1904
rect 764 1956 772 1964
rect 492 1916 500 1924
rect 556 1916 564 1924
rect 684 1916 692 1924
rect 780 1916 788 1924
rect 444 1876 452 1884
rect 188 1856 196 1864
rect 252 1856 260 1864
rect 380 1856 388 1864
rect 460 1856 468 1864
rect 508 1856 516 1864
rect 188 1836 196 1844
rect 236 1776 244 1784
rect 140 1756 148 1764
rect 268 1836 276 1844
rect 380 1836 388 1844
rect 252 1756 260 1764
rect 188 1576 196 1584
rect 236 1556 244 1564
rect 220 1536 228 1544
rect 124 1516 132 1524
rect 76 1496 84 1504
rect 108 1496 116 1504
rect 156 1496 164 1504
rect 204 1496 212 1504
rect 92 1476 100 1484
rect 12 1356 20 1364
rect 12 1276 20 1284
rect 76 1356 84 1364
rect 44 1336 52 1344
rect 140 1476 148 1484
rect 140 1376 148 1384
rect 396 1776 404 1784
rect 300 1756 308 1764
rect 476 1736 484 1744
rect 332 1716 340 1724
rect 380 1716 388 1724
rect 412 1716 420 1724
rect 524 1756 532 1764
rect 636 1896 644 1904
rect 652 1896 660 1904
rect 668 1896 676 1904
rect 636 1876 644 1884
rect 604 1856 612 1864
rect 556 1756 564 1764
rect 540 1736 548 1744
rect 604 1756 612 1764
rect 572 1716 580 1724
rect 444 1656 452 1664
rect 332 1576 340 1584
rect 268 1556 276 1564
rect 316 1516 324 1524
rect 364 1516 372 1524
rect 604 1716 612 1724
rect 716 1876 724 1884
rect 732 1856 740 1864
rect 748 1856 756 1864
rect 780 1856 788 1864
rect 700 1736 708 1744
rect 748 1736 756 1744
rect 652 1716 660 1724
rect 700 1716 708 1724
rect 588 1696 596 1704
rect 492 1676 500 1684
rect 492 1536 500 1544
rect 780 1676 788 1684
rect 636 1536 644 1544
rect 284 1496 292 1504
rect 332 1496 340 1504
rect 412 1496 420 1504
rect 476 1496 484 1504
rect 492 1496 500 1504
rect 188 1456 196 1464
rect 188 1436 196 1444
rect 140 1256 148 1264
rect 12 1096 20 1104
rect 28 1076 36 1084
rect 28 1016 36 1024
rect 124 1156 132 1164
rect 60 1116 68 1124
rect 108 1116 116 1124
rect 76 1096 84 1104
rect 316 1476 324 1484
rect 252 1416 260 1424
rect 380 1456 388 1464
rect 396 1456 404 1464
rect 460 1456 468 1464
rect 412 1436 420 1444
rect 444 1436 452 1444
rect 348 1416 356 1424
rect 332 1396 340 1404
rect 300 1376 308 1384
rect 236 1356 244 1364
rect 332 1356 340 1364
rect 380 1356 388 1364
rect 284 1336 292 1344
rect 236 1316 244 1324
rect 300 1296 308 1304
rect 252 1276 260 1284
rect 220 1256 228 1264
rect 444 1316 452 1324
rect 380 1296 388 1304
rect 412 1296 420 1304
rect 412 1136 420 1144
rect 364 1116 372 1124
rect 332 1096 340 1104
rect 380 1096 388 1104
rect 220 1076 228 1084
rect 60 1056 68 1064
rect 156 1056 164 1064
rect 284 1036 292 1044
rect 92 1016 100 1024
rect 108 916 116 924
rect 92 756 100 764
rect 76 656 84 664
rect 28 576 36 584
rect 92 596 100 604
rect 140 996 148 1004
rect 140 796 148 804
rect 124 736 132 744
rect 124 716 132 724
rect 188 1016 196 1024
rect 220 1016 228 1024
rect 476 1416 484 1424
rect 556 1516 564 1524
rect 604 1496 612 1504
rect 588 1456 596 1464
rect 620 1456 628 1464
rect 556 1436 564 1444
rect 748 1516 756 1524
rect 876 1956 884 1964
rect 1068 2136 1076 2144
rect 860 1916 868 1924
rect 940 1896 948 1904
rect 972 1876 980 1884
rect 1036 1876 1044 1884
rect 924 1856 932 1864
rect 924 1776 932 1784
rect 1020 1776 1028 1784
rect 828 1756 836 1764
rect 1260 2776 1268 2784
rect 1276 2756 1284 2764
rect 1244 2736 1252 2744
rect 1180 2716 1188 2724
rect 1212 2696 1220 2704
rect 1244 2696 1252 2704
rect 1100 2676 1108 2684
rect 1196 2676 1204 2684
rect 1164 2656 1172 2664
rect 1100 2596 1108 2604
rect 1148 2556 1156 2564
rect 1116 2536 1124 2544
rect 1132 2516 1140 2524
rect 1180 2596 1188 2604
rect 1180 2576 1188 2584
rect 1356 2836 1364 2844
rect 1358 2806 1366 2814
rect 1372 2806 1380 2814
rect 1386 2806 1394 2814
rect 1372 2736 1380 2744
rect 1228 2676 1236 2684
rect 1260 2676 1268 2684
rect 1292 2676 1300 2684
rect 1308 2676 1316 2684
rect 1324 2656 1332 2664
rect 1340 2636 1348 2644
rect 1372 2636 1380 2644
rect 1228 2556 1236 2564
rect 1468 3056 1476 3064
rect 1452 3016 1460 3024
rect 1500 3016 1508 3024
rect 1436 2896 1444 2904
rect 1436 2776 1444 2784
rect 1500 2976 1508 2984
rect 1516 2956 1524 2964
rect 1676 3116 1684 3124
rect 1692 3096 1700 3104
rect 1564 3076 1572 3084
rect 1580 3076 1588 3084
rect 1612 3076 1620 3084
rect 1932 3116 1940 3124
rect 1756 3096 1764 3104
rect 1724 3056 1732 3064
rect 1548 3016 1556 3024
rect 1596 3016 1604 3024
rect 1564 2996 1572 3004
rect 1548 2956 1556 2964
rect 1596 2956 1604 2964
rect 1468 2936 1476 2944
rect 1484 2896 1492 2904
rect 1468 2876 1476 2884
rect 1452 2756 1460 2764
rect 1484 2736 1492 2744
rect 1500 2716 1508 2724
rect 1468 2696 1476 2704
rect 1836 3036 1844 3044
rect 1676 2976 1684 2984
rect 1692 2976 1700 2984
rect 1756 2976 1764 2984
rect 1788 2976 1796 2984
rect 1708 2956 1716 2964
rect 1788 2956 1796 2964
rect 1820 2976 1828 2984
rect 1852 2936 1860 2944
rect 1996 3096 2004 3104
rect 2124 3318 2132 3324
rect 2124 3316 2132 3318
rect 2188 3316 2196 3324
rect 2284 3276 2292 3284
rect 2124 3196 2132 3204
rect 2284 3156 2292 3164
rect 2348 3316 2356 3324
rect 2444 3456 2452 3464
rect 2476 3456 2484 3464
rect 2428 3356 2436 3364
rect 2492 3436 2500 3444
rect 2460 3356 2468 3364
rect 2444 3336 2452 3344
rect 2396 3296 2404 3304
rect 2348 3176 2356 3184
rect 2316 3116 2324 3124
rect 2316 3096 2324 3104
rect 2300 3076 2308 3084
rect 1532 2896 1540 2904
rect 1580 2896 1588 2904
rect 1612 2896 1620 2904
rect 1804 2916 1812 2924
rect 1868 2916 1876 2924
rect 2044 2916 2052 2924
rect 2108 2918 2116 2924
rect 2108 2916 2116 2918
rect 1628 2876 1636 2884
rect 1852 2876 1860 2884
rect 1564 2836 1572 2844
rect 1740 2836 1748 2844
rect 1516 2676 1524 2684
rect 1532 2676 1540 2684
rect 1548 2656 1556 2664
rect 1692 2736 1700 2744
rect 1660 2716 1668 2724
rect 1724 2716 1732 2724
rect 1580 2696 1588 2704
rect 1612 2696 1620 2704
rect 1628 2696 1636 2704
rect 1692 2696 1700 2704
rect 1596 2656 1604 2664
rect 1644 2656 1652 2664
rect 1532 2536 1540 2544
rect 1564 2536 1572 2544
rect 1500 2516 1508 2524
rect 1548 2516 1556 2524
rect 1468 2436 1476 2444
rect 1358 2406 1366 2414
rect 1372 2406 1380 2414
rect 1386 2406 1394 2414
rect 1100 2376 1108 2384
rect 1308 2376 1316 2384
rect 1292 2336 1300 2344
rect 1404 2316 1412 2324
rect 1612 2496 1620 2504
rect 1516 2416 1524 2424
rect 1532 2316 1540 2324
rect 1596 2476 1604 2484
rect 1788 2716 1796 2724
rect 1900 2876 1908 2884
rect 1980 2856 1988 2864
rect 2284 2836 2292 2844
rect 1916 2736 1924 2744
rect 2204 2736 2212 2744
rect 2172 2716 2180 2724
rect 2108 2702 2116 2704
rect 2108 2696 2116 2702
rect 1772 2676 1780 2684
rect 1756 2636 1764 2644
rect 1820 2636 1828 2644
rect 1676 2596 1684 2604
rect 1708 2596 1716 2604
rect 1692 2576 1700 2584
rect 1692 2516 1700 2524
rect 1532 2296 1540 2304
rect 1580 2296 1588 2304
rect 1596 2296 1604 2304
rect 1516 2276 1524 2284
rect 1100 2256 1108 2264
rect 1164 2216 1172 2224
rect 1180 2136 1188 2144
rect 1244 2118 1252 2124
rect 1244 2116 1252 2118
rect 1116 2036 1124 2044
rect 1212 1956 1220 1964
rect 1100 1916 1108 1924
rect 1644 2156 1652 2164
rect 1804 2556 1812 2564
rect 1756 2536 1764 2544
rect 1820 2536 1828 2544
rect 1772 2516 1780 2524
rect 1788 2516 1796 2524
rect 1772 2496 1780 2504
rect 1756 2476 1764 2484
rect 1804 2456 1812 2464
rect 1980 2636 1988 2644
rect 1900 2596 1908 2604
rect 1980 2596 1988 2604
rect 1868 2556 1876 2564
rect 1932 2556 1940 2564
rect 1996 2556 2004 2564
rect 2300 2676 2308 2684
rect 2156 2636 2164 2644
rect 2188 2576 2196 2584
rect 2332 2696 2340 2704
rect 2412 3136 2420 3144
rect 2444 3136 2452 3144
rect 2396 3076 2404 3084
rect 2444 3116 2452 3124
rect 2428 3096 2436 3104
rect 2684 3556 2692 3564
rect 2668 3536 2676 3544
rect 2764 3536 2772 3544
rect 2780 3516 2788 3524
rect 3036 3876 3044 3884
rect 3020 3856 3028 3864
rect 2860 3836 2868 3844
rect 2876 3836 2884 3844
rect 2876 3816 2884 3824
rect 2910 3806 2918 3814
rect 2924 3806 2932 3814
rect 2938 3806 2946 3814
rect 2876 3776 2884 3784
rect 2876 3756 2884 3764
rect 2892 3736 2900 3744
rect 2860 3696 2868 3704
rect 2652 3496 2660 3504
rect 2748 3496 2756 3504
rect 2556 3456 2564 3464
rect 2508 3376 2516 3384
rect 2540 3376 2548 3384
rect 2540 3356 2548 3364
rect 2508 3316 2516 3324
rect 2524 3316 2532 3324
rect 2620 3416 2628 3424
rect 2620 3396 2628 3404
rect 2748 3456 2756 3464
rect 2716 3416 2724 3424
rect 2668 3396 2676 3404
rect 2700 3376 2708 3384
rect 2636 3356 2644 3364
rect 2684 3356 2692 3364
rect 2652 3336 2660 3344
rect 2636 3316 2644 3324
rect 2556 3296 2564 3304
rect 2668 3296 2676 3304
rect 2492 3136 2500 3144
rect 2476 3116 2484 3124
rect 2460 3096 2468 3104
rect 2508 3096 2516 3104
rect 2524 3076 2532 3084
rect 2556 3256 2564 3264
rect 2604 3156 2612 3164
rect 2636 3136 2644 3144
rect 2684 3176 2692 3184
rect 2732 3356 2740 3364
rect 2892 3576 2900 3584
rect 2924 3536 2932 3544
rect 2940 3516 2948 3524
rect 3052 3796 3060 3804
rect 3020 3736 3028 3744
rect 3052 3736 3060 3744
rect 3116 3796 3124 3804
rect 3116 3776 3124 3784
rect 3180 3756 3188 3764
rect 3244 3976 3252 3984
rect 3308 3976 3316 3984
rect 3260 3916 3268 3924
rect 3212 3896 3220 3904
rect 3276 3896 3284 3904
rect 3228 3856 3236 3864
rect 3228 3796 3236 3804
rect 3020 3696 3028 3704
rect 3036 3516 3044 3524
rect 2940 3496 2948 3504
rect 2988 3496 2996 3504
rect 2844 3456 2852 3464
rect 2956 3456 2964 3464
rect 3020 3456 3028 3464
rect 2828 3376 2836 3384
rect 2988 3436 2996 3444
rect 2910 3406 2918 3414
rect 2924 3406 2932 3414
rect 2938 3406 2946 3414
rect 3484 3896 3492 3904
rect 3532 3896 3540 3904
rect 3564 4036 3572 4044
rect 3676 4016 3684 4024
rect 3612 3896 3620 3904
rect 3420 3876 3428 3884
rect 3484 3876 3492 3884
rect 3548 3876 3556 3884
rect 3580 3876 3588 3884
rect 3692 3876 3700 3884
rect 3516 3756 3524 3764
rect 3436 3736 3444 3744
rect 3628 3756 3636 3764
rect 3852 4116 3860 4124
rect 3756 4096 3764 4104
rect 3772 3896 3780 3904
rect 4188 4156 4196 4164
rect 3900 4136 3908 4144
rect 3932 4116 3940 4124
rect 3900 4096 3908 4104
rect 3980 4096 3988 4104
rect 4332 4136 4340 4144
rect 4364 4136 4372 4144
rect 4316 4116 4324 4124
rect 4220 4096 4228 4104
rect 4364 4096 4372 4104
rect 4012 4076 4020 4084
rect 4108 4036 4116 4044
rect 4028 3996 4036 4004
rect 3964 3896 3972 3904
rect 4028 3902 4036 3904
rect 4028 3896 4036 3902
rect 4780 4196 4788 4204
rect 4396 4176 4404 4184
rect 4796 4156 4804 4164
rect 4140 3896 4148 3904
rect 4236 3896 4244 3904
rect 4284 3896 4292 3904
rect 3740 3876 3748 3884
rect 4108 3876 4116 3884
rect 4188 3876 4196 3884
rect 3724 3776 3732 3784
rect 3676 3756 3684 3764
rect 3740 3756 3748 3764
rect 3820 3756 3828 3764
rect 3612 3736 3620 3744
rect 3628 3736 3636 3744
rect 3644 3736 3652 3744
rect 3852 3736 3860 3744
rect 3500 3716 3508 3724
rect 3772 3716 3780 3724
rect 3244 3696 3252 3704
rect 3340 3616 3348 3624
rect 3260 3556 3268 3564
rect 3148 3496 3156 3504
rect 3212 3476 3220 3484
rect 3260 3476 3268 3484
rect 3100 3456 3108 3464
rect 3116 3416 3124 3424
rect 3308 3456 3316 3464
rect 3276 3436 3284 3444
rect 3180 3416 3188 3424
rect 3084 3396 3092 3404
rect 3116 3396 3124 3404
rect 3132 3396 3140 3404
rect 3148 3376 3156 3384
rect 2812 3356 2820 3364
rect 2844 3356 2852 3364
rect 3020 3356 3028 3364
rect 3068 3356 3076 3364
rect 3116 3356 3124 3364
rect 2732 3336 2740 3344
rect 2764 3336 2772 3344
rect 2748 3316 2756 3324
rect 3004 3336 3012 3344
rect 2956 3316 2964 3324
rect 2764 3296 2772 3304
rect 2796 3296 2804 3304
rect 2764 3256 2772 3264
rect 2732 3176 2740 3184
rect 2892 3136 2900 3144
rect 2716 3116 2724 3124
rect 2860 3102 2868 3104
rect 2860 3096 2868 3102
rect 2924 3076 2932 3084
rect 2540 2976 2548 2984
rect 2460 2956 2468 2964
rect 2700 2936 2708 2944
rect 2460 2916 2468 2924
rect 2636 2916 2644 2924
rect 2910 3006 2918 3014
rect 2924 3006 2932 3014
rect 2938 3006 2946 3014
rect 2828 2916 2836 2924
rect 2892 2918 2900 2924
rect 2892 2916 2900 2918
rect 2572 2836 2580 2844
rect 2604 2836 2612 2844
rect 2412 2716 2420 2724
rect 2492 2716 2500 2724
rect 2588 2716 2596 2724
rect 2380 2696 2388 2704
rect 2428 2696 2436 2704
rect 2508 2696 2516 2704
rect 2572 2696 2580 2704
rect 2396 2676 2404 2684
rect 2460 2676 2468 2684
rect 2508 2676 2516 2684
rect 2556 2680 2564 2684
rect 2556 2676 2564 2680
rect 2348 2656 2356 2664
rect 2444 2656 2452 2664
rect 2620 2736 2628 2744
rect 2620 2656 2628 2664
rect 2604 2596 2612 2604
rect 2412 2576 2420 2584
rect 2620 2576 2628 2584
rect 2300 2556 2308 2564
rect 2556 2536 2564 2544
rect 1868 2516 1876 2524
rect 1900 2516 1908 2524
rect 2124 2518 2132 2524
rect 2124 2516 2132 2518
rect 2156 2516 2164 2524
rect 3324 3396 3332 3404
rect 3196 3356 3204 3364
rect 3068 3336 3076 3344
rect 3532 3696 3540 3704
rect 3452 3502 3460 3504
rect 3452 3496 3460 3502
rect 3516 3496 3524 3504
rect 3484 3476 3492 3484
rect 3548 3676 3556 3684
rect 3756 3696 3764 3704
rect 3804 3696 3812 3704
rect 3660 3676 3668 3684
rect 3692 3576 3700 3584
rect 3644 3496 3652 3504
rect 3740 3496 3748 3504
rect 3708 3476 3716 3484
rect 3548 3436 3556 3444
rect 3564 3396 3572 3404
rect 3228 3336 3236 3344
rect 3804 3676 3812 3684
rect 3788 3576 3796 3584
rect 3932 3776 3940 3784
rect 3900 3756 3908 3764
rect 3996 3718 4004 3724
rect 3996 3716 4004 3718
rect 3884 3556 3892 3564
rect 4332 3816 4340 3824
rect 4348 3796 4356 3804
rect 4204 3776 4212 3784
rect 4284 3776 4292 3784
rect 4060 3716 4068 3724
rect 4188 3716 4196 3724
rect 4124 3636 4132 3644
rect 4108 3536 4116 3544
rect 4124 3516 4132 3524
rect 4172 3516 4180 3524
rect 4060 3502 4068 3504
rect 4060 3496 4068 3502
rect 4124 3496 4132 3504
rect 4156 3496 4164 3504
rect 4028 3476 4036 3484
rect 4172 3476 4180 3484
rect 3756 3396 3764 3404
rect 3820 3336 3828 3344
rect 3468 3318 3476 3324
rect 3468 3316 3476 3318
rect 3532 3316 3540 3324
rect 3548 3316 3556 3324
rect 3692 3318 3700 3324
rect 3692 3316 3700 3318
rect 3100 3296 3108 3304
rect 3020 3276 3028 3284
rect 3260 3196 3268 3204
rect 3372 3156 3380 3164
rect 3100 3136 3108 3144
rect 3164 3116 3172 3124
rect 3228 3116 3236 3124
rect 3308 3116 3316 3124
rect 3276 3096 3284 3104
rect 3036 3076 3044 3084
rect 3308 3076 3316 3084
rect 3356 3096 3364 3104
rect 3388 3116 3396 3124
rect 3388 3076 3396 3084
rect 3324 3056 3332 3064
rect 3228 2936 3236 2944
rect 3036 2916 3044 2924
rect 2828 2896 2836 2904
rect 2972 2896 2980 2904
rect 3020 2896 3028 2904
rect 2764 2836 2772 2844
rect 2684 2736 2692 2744
rect 2652 2696 2660 2704
rect 2812 2676 2820 2684
rect 3164 2896 3172 2904
rect 3180 2836 3188 2844
rect 3052 2736 3060 2744
rect 3132 2736 3140 2744
rect 2956 2696 2964 2704
rect 3004 2696 3012 2704
rect 3036 2696 3044 2704
rect 3116 2716 3124 2724
rect 2940 2676 2948 2684
rect 3084 2676 3092 2684
rect 2796 2656 2804 2664
rect 2828 2656 2836 2664
rect 2844 2656 2852 2664
rect 3052 2656 3060 2664
rect 3164 2696 3172 2704
rect 3516 3276 3524 3284
rect 3644 3176 3652 3184
rect 3420 3156 3428 3164
rect 3532 3136 3540 3144
rect 3548 3136 3556 3144
rect 3436 3116 3444 3124
rect 3452 3116 3460 3124
rect 3484 3096 3492 3104
rect 3916 3396 3924 3404
rect 3932 3396 3940 3404
rect 3900 3356 3908 3364
rect 3868 3336 3876 3344
rect 3836 3316 3844 3324
rect 3788 3296 3796 3304
rect 3772 3276 3780 3284
rect 3836 3296 3844 3304
rect 3804 3236 3812 3244
rect 3820 3216 3828 3224
rect 3772 3156 3780 3164
rect 3756 3116 3764 3124
rect 3804 3096 3812 3104
rect 3660 3076 3668 3084
rect 3436 3056 3444 3064
rect 3756 3056 3764 3064
rect 3436 2996 3444 3004
rect 3676 2996 3684 3004
rect 3884 3236 3892 3244
rect 4188 3396 4196 3404
rect 4076 3376 4084 3384
rect 4108 3336 4116 3344
rect 3916 3236 3924 3244
rect 3900 3216 3908 3224
rect 3852 3176 3860 3184
rect 3852 3096 3860 3104
rect 3884 3096 3892 3104
rect 3868 3076 3876 3084
rect 3820 3056 3828 3064
rect 3884 3056 3892 3064
rect 3948 3216 3956 3224
rect 4044 3136 4052 3144
rect 3964 3096 3972 3104
rect 4172 3176 4180 3184
rect 3932 3076 3940 3084
rect 3964 3076 3972 3084
rect 4012 3076 4020 3084
rect 4140 3076 4148 3084
rect 3916 3036 3924 3044
rect 3980 3036 3988 3044
rect 3772 3016 3780 3024
rect 3612 2936 3620 2944
rect 3692 2936 3700 2944
rect 3404 2916 3412 2924
rect 3548 2916 3556 2924
rect 3740 2916 3748 2924
rect 3420 2876 3428 2884
rect 3292 2836 3300 2844
rect 3484 2736 3492 2744
rect 3548 2716 3556 2724
rect 3644 2716 3652 2724
rect 3212 2696 3220 2704
rect 3276 2696 3284 2704
rect 3116 2676 3124 2684
rect 3180 2676 3188 2684
rect 2876 2636 2884 2644
rect 3100 2636 3108 2644
rect 2910 2606 2918 2614
rect 2924 2606 2932 2614
rect 2938 2606 2946 2614
rect 3212 2656 3220 2664
rect 3292 2676 3300 2684
rect 3244 2616 3252 2624
rect 3196 2576 3204 2584
rect 2732 2556 2740 2564
rect 2812 2536 2820 2544
rect 2588 2516 2596 2524
rect 2636 2516 2644 2524
rect 2684 2516 2692 2524
rect 3196 2556 3204 2564
rect 3292 2616 3300 2624
rect 3340 2696 3348 2704
rect 3612 2696 3620 2704
rect 3708 2696 3716 2704
rect 3340 2676 3348 2684
rect 3388 2676 3396 2684
rect 3420 2676 3428 2684
rect 3580 2676 3588 2684
rect 3340 2656 3348 2664
rect 3404 2656 3412 2664
rect 3324 2636 3332 2644
rect 3276 2576 3284 2584
rect 3308 2576 3316 2584
rect 3260 2556 3268 2564
rect 3100 2536 3108 2544
rect 3212 2536 3220 2544
rect 3244 2536 3252 2544
rect 3324 2536 3332 2544
rect 3452 2656 3460 2664
rect 3404 2576 3412 2584
rect 3500 2556 3508 2564
rect 3436 2536 3444 2544
rect 3500 2536 3508 2544
rect 1932 2476 1940 2484
rect 1852 2456 1860 2464
rect 1820 2416 1828 2424
rect 1852 2296 1860 2304
rect 1964 2296 1972 2304
rect 2044 2296 2052 2304
rect 2108 2336 2116 2344
rect 2236 2296 2244 2304
rect 2380 2336 2388 2344
rect 2300 2316 2308 2324
rect 2396 2316 2404 2324
rect 2972 2516 2980 2524
rect 3036 2518 3044 2524
rect 3036 2516 3044 2518
rect 3228 2516 3236 2524
rect 3244 2516 3252 2524
rect 3340 2516 3348 2524
rect 3372 2516 3380 2524
rect 2748 2496 2756 2504
rect 3132 2496 3140 2504
rect 3212 2496 3220 2504
rect 3244 2496 3252 2504
rect 3340 2496 3348 2504
rect 3452 2496 3460 2504
rect 2972 2336 2980 2344
rect 3276 2336 3284 2344
rect 2460 2296 2468 2304
rect 2844 2296 2852 2304
rect 2380 2276 2388 2284
rect 2492 2276 2500 2284
rect 1836 2256 1844 2264
rect 1916 2236 1924 2244
rect 1980 2236 1988 2244
rect 2172 2236 2180 2244
rect 2364 2236 2372 2244
rect 2620 2236 2628 2244
rect 1740 2156 1748 2164
rect 1468 2116 1476 2124
rect 1564 2116 1572 2124
rect 1660 2116 1668 2124
rect 1708 2116 1716 2124
rect 1358 2006 1366 2014
rect 1372 2006 1380 2014
rect 1386 2006 1394 2014
rect 1292 1896 1300 1904
rect 1516 1902 1524 1904
rect 1516 1896 1524 1902
rect 1084 1876 1092 1884
rect 1132 1876 1140 1884
rect 940 1736 948 1744
rect 1116 1736 1124 1744
rect 812 1696 820 1704
rect 684 1476 692 1484
rect 668 1456 676 1464
rect 780 1456 788 1464
rect 604 1436 612 1444
rect 652 1436 660 1444
rect 748 1416 756 1424
rect 620 1396 628 1404
rect 684 1356 692 1364
rect 572 1316 580 1324
rect 524 1296 532 1304
rect 540 1296 548 1304
rect 572 1296 580 1304
rect 476 1176 484 1184
rect 508 1176 516 1184
rect 524 1176 532 1184
rect 444 1096 452 1104
rect 332 1076 340 1084
rect 364 1076 372 1084
rect 412 1076 420 1084
rect 428 1076 436 1084
rect 348 1056 356 1064
rect 332 1036 340 1044
rect 268 936 276 944
rect 300 916 308 924
rect 172 816 180 824
rect 156 716 164 724
rect 172 716 180 724
rect 204 776 212 784
rect 348 936 356 944
rect 492 1116 500 1124
rect 476 1076 484 1084
rect 508 1096 516 1104
rect 460 1016 468 1024
rect 540 1156 548 1164
rect 620 1316 628 1324
rect 764 1336 772 1344
rect 780 1316 788 1324
rect 652 1296 660 1304
rect 636 1276 644 1284
rect 700 1196 708 1204
rect 652 1136 660 1144
rect 636 1096 644 1104
rect 732 1196 740 1204
rect 876 1716 884 1724
rect 860 1496 868 1504
rect 828 1476 836 1484
rect 828 1356 836 1364
rect 892 1476 900 1484
rect 892 1436 900 1444
rect 860 1376 868 1384
rect 796 1296 804 1304
rect 812 1296 820 1304
rect 828 1176 836 1184
rect 780 1136 788 1144
rect 748 1116 756 1124
rect 844 1116 852 1124
rect 540 1076 548 1084
rect 652 1076 660 1084
rect 684 1076 692 1084
rect 716 1076 724 1084
rect 812 1076 820 1084
rect 604 1056 612 1064
rect 652 1056 660 1064
rect 828 1056 836 1064
rect 380 936 388 944
rect 412 936 420 944
rect 524 956 532 964
rect 588 956 596 964
rect 732 956 740 964
rect 604 936 612 944
rect 636 936 644 944
rect 652 936 660 944
rect 364 916 372 924
rect 620 916 628 924
rect 684 916 692 924
rect 812 916 820 924
rect 316 896 324 904
rect 716 896 724 904
rect 732 896 740 904
rect 764 896 772 904
rect 780 896 788 904
rect 332 876 340 884
rect 300 816 308 824
rect 284 776 292 784
rect 268 756 276 764
rect 236 736 244 744
rect 252 736 260 744
rect 124 696 132 704
rect 140 696 148 704
rect 188 696 196 704
rect 172 676 180 684
rect 156 656 164 664
rect 108 576 116 584
rect 220 656 228 664
rect 204 616 212 624
rect 12 516 20 524
rect 12 256 20 264
rect 540 876 548 884
rect 748 876 756 884
rect 476 856 484 864
rect 572 856 580 864
rect 412 776 420 784
rect 780 776 788 784
rect 396 756 404 764
rect 316 716 324 724
rect 908 1396 916 1404
rect 908 1376 916 1384
rect 924 1376 932 1384
rect 924 1336 932 1344
rect 1004 1636 1012 1644
rect 1100 1718 1108 1724
rect 1100 1716 1108 1718
rect 1196 1696 1204 1704
rect 1100 1636 1108 1644
rect 1036 1616 1044 1624
rect 1084 1556 1092 1564
rect 1036 1536 1044 1544
rect 1068 1536 1076 1544
rect 972 1496 980 1504
rect 988 1496 996 1504
rect 1068 1496 1076 1504
rect 972 1456 980 1464
rect 1036 1456 1044 1464
rect 1116 1616 1124 1624
rect 1100 1536 1108 1544
rect 1148 1496 1156 1504
rect 1452 1836 1460 1844
rect 1804 2176 1812 2184
rect 2044 2176 2052 2184
rect 1884 2156 1892 2164
rect 1772 2136 1780 2144
rect 1820 2136 1828 2144
rect 1836 2136 1844 2144
rect 1932 2136 1940 2144
rect 2076 2136 2084 2144
rect 1932 2116 1940 2124
rect 1868 2096 1876 2104
rect 1980 2116 1988 2124
rect 2204 2176 2212 2184
rect 2252 2176 2260 2184
rect 2300 2136 2308 2144
rect 2348 2136 2356 2144
rect 2172 2116 2180 2124
rect 2220 2116 2228 2124
rect 2268 2116 2276 2124
rect 2460 2136 2468 2144
rect 2588 2136 2596 2144
rect 2412 2116 2420 2124
rect 2476 2116 2484 2124
rect 2652 2116 2660 2124
rect 1964 2096 1972 2104
rect 2332 2096 2340 2104
rect 1884 2076 1892 2084
rect 2012 2076 2020 2084
rect 1868 1956 1876 1964
rect 1900 1956 1908 1964
rect 1804 1896 1812 1904
rect 1724 1856 1732 1864
rect 1532 1816 1540 1824
rect 1244 1736 1252 1744
rect 1452 1736 1460 1744
rect 1548 1736 1556 1744
rect 1324 1716 1332 1724
rect 1276 1696 1284 1704
rect 1580 1718 1588 1724
rect 1580 1716 1588 1718
rect 1388 1656 1396 1664
rect 1358 1606 1366 1614
rect 1372 1606 1380 1614
rect 1386 1606 1394 1614
rect 1228 1576 1236 1584
rect 1420 1536 1428 1544
rect 1260 1496 1268 1504
rect 1100 1356 1108 1364
rect 940 1316 948 1324
rect 1084 1316 1092 1324
rect 1212 1456 1220 1464
rect 1228 1436 1236 1444
rect 1180 1376 1188 1384
rect 1164 1336 1172 1344
rect 1132 1316 1140 1324
rect 1148 1316 1156 1324
rect 1116 1296 1124 1304
rect 892 1276 900 1284
rect 972 1276 980 1284
rect 876 1236 884 1244
rect 1052 1216 1060 1224
rect 1020 1196 1028 1204
rect 1084 1156 1092 1164
rect 924 1116 932 1124
rect 972 1116 980 1124
rect 1116 1116 1124 1124
rect 892 1096 900 1104
rect 988 1096 996 1104
rect 1052 1096 1060 1104
rect 1084 1096 1092 1104
rect 876 1076 884 1084
rect 1036 1076 1044 1084
rect 860 1016 868 1024
rect 892 1056 900 1064
rect 940 1056 948 1064
rect 988 1056 996 1064
rect 1020 1056 1028 1064
rect 1052 1036 1060 1044
rect 1004 976 1012 984
rect 1100 1056 1108 1064
rect 940 956 948 964
rect 988 956 996 964
rect 1004 956 1012 964
rect 1084 956 1092 964
rect 844 936 852 944
rect 892 936 900 944
rect 908 936 916 944
rect 972 936 980 944
rect 956 916 964 924
rect 988 916 996 924
rect 1084 916 1092 924
rect 844 896 852 904
rect 668 756 676 764
rect 764 756 772 764
rect 828 756 836 764
rect 732 736 740 744
rect 444 716 452 724
rect 668 716 676 724
rect 748 716 756 724
rect 428 696 436 704
rect 508 696 516 704
rect 556 696 564 704
rect 620 696 628 704
rect 364 676 372 684
rect 316 656 324 664
rect 316 636 324 644
rect 252 576 260 584
rect 124 536 132 544
rect 236 536 244 544
rect 92 516 100 524
rect 76 316 84 324
rect 108 336 116 344
rect 140 516 148 524
rect 204 516 212 524
rect 188 496 196 504
rect 236 496 244 504
rect 124 316 132 324
rect 300 576 308 584
rect 380 636 388 644
rect 332 596 340 604
rect 428 616 436 624
rect 412 576 420 584
rect 364 556 372 564
rect 380 556 388 564
rect 348 536 356 544
rect 284 516 292 524
rect 380 516 388 524
rect 396 516 404 524
rect 348 496 356 504
rect 508 636 516 644
rect 604 676 612 684
rect 620 676 628 684
rect 556 616 564 624
rect 796 736 804 744
rect 828 736 836 744
rect 1036 796 1044 804
rect 1020 716 1028 724
rect 1196 1296 1204 1304
rect 1180 1276 1188 1284
rect 1148 1236 1156 1244
rect 1148 1176 1156 1184
rect 1212 1116 1220 1124
rect 1148 996 1156 1004
rect 1148 876 1156 884
rect 1132 736 1140 744
rect 1052 716 1060 724
rect 764 676 772 684
rect 924 676 932 684
rect 972 676 980 684
rect 988 676 996 684
rect 636 636 644 644
rect 540 556 548 564
rect 620 556 628 564
rect 668 556 676 564
rect 684 516 692 524
rect 492 496 500 504
rect 556 496 564 504
rect 428 476 436 484
rect 300 356 308 364
rect 204 336 212 344
rect 268 336 276 344
rect 428 336 436 344
rect 364 316 372 324
rect 396 316 404 324
rect 524 336 532 344
rect 12 196 20 204
rect 44 196 52 204
rect 28 136 36 144
rect 140 296 148 304
rect 172 296 180 304
rect 188 296 196 304
rect 236 296 244 304
rect 316 296 324 304
rect 444 296 452 304
rect 492 296 500 304
rect 92 276 100 284
rect 252 276 260 284
rect 444 276 452 284
rect 684 376 692 384
rect 636 316 644 324
rect 860 656 868 664
rect 940 656 948 664
rect 796 616 804 624
rect 780 556 788 564
rect 860 576 868 584
rect 812 556 820 564
rect 860 556 868 564
rect 972 576 980 584
rect 748 516 756 524
rect 780 516 788 524
rect 892 536 900 544
rect 1036 656 1044 664
rect 1068 656 1076 664
rect 1052 636 1060 644
rect 956 536 964 544
rect 908 516 916 524
rect 844 496 852 504
rect 1276 1416 1284 1424
rect 1340 1476 1348 1484
rect 1340 1456 1348 1464
rect 1580 1516 1588 1524
rect 1468 1456 1476 1464
rect 1516 1456 1524 1464
rect 1836 1836 1844 1844
rect 1724 1816 1732 1824
rect 1852 1816 1860 1824
rect 1868 1776 1876 1784
rect 1852 1756 1860 1764
rect 1836 1736 1844 1744
rect 1820 1716 1828 1724
rect 1788 1656 1796 1664
rect 1708 1616 1716 1624
rect 1644 1496 1652 1504
rect 1724 1496 1732 1504
rect 1580 1436 1588 1444
rect 1628 1436 1636 1444
rect 1356 1416 1364 1424
rect 1468 1356 1476 1364
rect 1484 1356 1492 1364
rect 1260 1336 1268 1344
rect 1308 1336 1316 1344
rect 1260 1316 1268 1324
rect 1244 996 1252 1004
rect 1484 1296 1492 1304
rect 1276 1276 1284 1284
rect 1358 1206 1366 1214
rect 1372 1206 1380 1214
rect 1386 1206 1394 1214
rect 1308 1176 1316 1184
rect 1372 1156 1380 1164
rect 1340 1116 1348 1124
rect 1276 1096 1284 1104
rect 1276 1076 1284 1084
rect 1212 956 1220 964
rect 1228 936 1236 944
rect 1244 916 1252 924
rect 1212 856 1220 864
rect 1212 816 1220 824
rect 1164 696 1172 704
rect 1132 656 1140 664
rect 1100 636 1108 644
rect 1228 696 1236 704
rect 1212 636 1220 644
rect 1228 636 1236 644
rect 1084 616 1092 624
rect 1132 616 1140 624
rect 1148 616 1156 624
rect 1180 616 1188 624
rect 1196 616 1204 624
rect 1100 556 1108 564
rect 1020 536 1028 544
rect 1116 536 1124 544
rect 1164 556 1172 564
rect 1228 536 1236 544
rect 1148 516 1156 524
rect 1180 516 1188 524
rect 1356 1056 1364 1064
rect 1340 976 1348 984
rect 1308 956 1316 964
rect 1404 936 1412 944
rect 1358 806 1366 814
rect 1372 806 1380 814
rect 1386 806 1394 814
rect 1308 736 1316 744
rect 1372 736 1380 744
rect 1868 1716 1876 1724
rect 1852 1696 1860 1704
rect 1916 1916 1924 1924
rect 1916 1896 1924 1904
rect 1980 1956 1988 1964
rect 1996 1916 2004 1924
rect 2028 1936 2036 1944
rect 2396 2056 2404 2064
rect 2236 1956 2244 1964
rect 2172 1916 2180 1924
rect 1932 1876 1940 1884
rect 2044 1876 2052 1884
rect 2172 1896 2180 1904
rect 2300 1936 2308 1944
rect 2268 1916 2276 1924
rect 2460 2076 2468 2084
rect 2492 2096 2500 2104
rect 2492 2076 2500 2084
rect 2492 2056 2500 2064
rect 2812 2256 2820 2264
rect 2732 2236 2740 2244
rect 2716 2176 2724 2184
rect 2828 2176 2836 2184
rect 3052 2316 3060 2324
rect 3388 2316 3396 2324
rect 2940 2296 2948 2304
rect 2956 2296 2964 2304
rect 3068 2296 3076 2304
rect 3708 2636 3716 2644
rect 3580 2616 3588 2624
rect 3532 2556 3540 2564
rect 3564 2536 3572 2544
rect 3564 2516 3572 2524
rect 3868 2976 3876 2984
rect 3948 2976 3956 2984
rect 4140 3016 4148 3024
rect 4028 2936 4036 2944
rect 4012 2916 4020 2924
rect 3836 2896 3844 2904
rect 3804 2856 3812 2864
rect 3820 2736 3828 2744
rect 3772 2696 3780 2704
rect 3900 2876 3908 2884
rect 3868 2776 3876 2784
rect 3980 2776 3988 2784
rect 4076 2916 4084 2924
rect 4044 2896 4052 2904
rect 4412 4116 4420 4124
rect 4492 4096 4500 4104
rect 4508 4076 4516 4084
rect 4446 4006 4454 4014
rect 4460 4006 4468 4014
rect 4474 4006 4482 4014
rect 4396 3816 4404 3824
rect 4396 3796 4404 3804
rect 4444 3796 4452 3804
rect 4316 3736 4324 3744
rect 4380 3736 4388 3744
rect 4380 3716 4388 3724
rect 4252 3536 4260 3544
rect 4316 3536 4324 3544
rect 4268 3516 4276 3524
rect 4300 3496 4308 3504
rect 4348 3496 4356 3504
rect 4268 3476 4276 3484
rect 4380 3476 4388 3484
rect 4636 4036 4644 4044
rect 4572 3996 4580 4004
rect 4636 3916 4644 3924
rect 4780 3916 4788 3924
rect 4732 3896 4740 3904
rect 4748 3876 4756 3884
rect 4780 3876 4788 3884
rect 4828 4096 4836 4104
rect 5068 4156 5076 4164
rect 4940 4136 4948 4144
rect 4972 4136 4980 4144
rect 5148 4156 5156 4164
rect 4924 4116 4932 4124
rect 4972 4096 4980 4104
rect 4860 3916 4868 3924
rect 4812 3896 4820 3904
rect 4748 3856 4756 3864
rect 4796 3856 4804 3864
rect 4604 3776 4612 3784
rect 4876 3856 4884 3864
rect 4812 3816 4820 3824
rect 4508 3756 4516 3764
rect 4556 3756 4564 3764
rect 4876 3756 4884 3764
rect 4540 3736 4548 3744
rect 4412 3716 4420 3724
rect 4460 3716 4468 3724
rect 4446 3606 4454 3614
rect 4460 3606 4468 3614
rect 4474 3606 4482 3614
rect 4412 3516 4420 3524
rect 4508 3516 4516 3524
rect 4492 3476 4500 3484
rect 4524 3496 4532 3504
rect 4572 3496 4580 3504
rect 4540 3476 4548 3484
rect 4236 3456 4244 3464
rect 4508 3456 4516 3464
rect 4428 3436 4436 3444
rect 4556 3436 4564 3444
rect 4492 3396 4500 3404
rect 4508 3396 4516 3404
rect 4236 3336 4244 3344
rect 4300 3336 4308 3344
rect 4332 3336 4340 3344
rect 4476 3336 4484 3344
rect 4268 3318 4276 3324
rect 4268 3316 4276 3318
rect 4364 3316 4372 3324
rect 4268 3256 4276 3264
rect 4252 3116 4260 3124
rect 4236 3076 4244 3084
rect 4028 2736 4036 2744
rect 3852 2716 3860 2724
rect 3884 2716 3892 2724
rect 3948 2716 3956 2724
rect 3868 2696 3876 2704
rect 3900 2696 3908 2704
rect 3740 2676 3748 2684
rect 3772 2676 3780 2684
rect 3820 2676 3828 2684
rect 3724 2596 3732 2604
rect 3660 2576 3668 2584
rect 3628 2536 3636 2544
rect 3804 2656 3812 2664
rect 3836 2636 3844 2644
rect 3676 2536 3684 2544
rect 3836 2536 3844 2544
rect 3980 2716 3988 2724
rect 4044 2716 4052 2724
rect 4220 2736 4228 2744
rect 4028 2656 4036 2664
rect 4124 2656 4132 2664
rect 3884 2636 3892 2644
rect 3932 2636 3940 2644
rect 3964 2636 3972 2644
rect 3932 2596 3940 2604
rect 3980 2596 3988 2604
rect 3996 2576 4004 2584
rect 4060 2576 4068 2584
rect 3948 2556 3956 2564
rect 4188 2576 4196 2584
rect 4108 2556 4116 2564
rect 4156 2536 4164 2544
rect 3612 2516 3620 2524
rect 3660 2516 3668 2524
rect 3804 2518 3812 2524
rect 3804 2516 3812 2518
rect 3900 2516 3908 2524
rect 3980 2516 3988 2524
rect 4092 2516 4100 2524
rect 3532 2496 3540 2504
rect 3644 2496 3652 2504
rect 4012 2356 4020 2364
rect 4446 3206 4454 3214
rect 4460 3206 4468 3214
rect 4474 3206 4482 3214
rect 4284 3156 4292 3164
rect 4444 3136 4452 3144
rect 4348 3116 4356 3124
rect 4380 3116 4388 3124
rect 4300 3096 4308 3104
rect 4396 3096 4404 3104
rect 4540 3336 4548 3344
rect 4556 3316 4564 3324
rect 4988 3896 4996 3904
rect 4780 3736 4788 3744
rect 4892 3736 4900 3744
rect 4876 3716 4884 3724
rect 4956 3856 4964 3864
rect 4924 3816 4932 3824
rect 4972 3756 4980 3764
rect 4956 3736 4964 3744
rect 4924 3716 4932 3724
rect 5020 4116 5028 4124
rect 5052 4096 5060 4104
rect 5260 4136 5268 4144
rect 5436 4136 5444 4144
rect 5052 3896 5060 3904
rect 5020 3836 5028 3844
rect 5004 3816 5012 3824
rect 5100 3796 5108 3804
rect 5020 3756 5028 3764
rect 5148 3836 5156 3844
rect 5372 4016 5380 4024
rect 5468 4116 5476 4124
rect 5580 4116 5588 4124
rect 5452 3876 5460 3884
rect 5244 3796 5252 3804
rect 5324 3816 5332 3824
rect 5308 3796 5316 3804
rect 5116 3716 5124 3724
rect 5148 3716 5156 3724
rect 5276 3716 5284 3724
rect 4988 3636 4996 3644
rect 5356 3636 5364 3644
rect 5420 3636 5428 3644
rect 4812 3576 4820 3584
rect 5004 3556 5012 3564
rect 4748 3536 4756 3544
rect 4844 3536 4852 3544
rect 4636 3516 4644 3524
rect 4684 3516 4692 3524
rect 4588 3476 4596 3484
rect 4684 3476 4692 3484
rect 4636 3356 4644 3364
rect 4604 3336 4612 3344
rect 4700 3396 4708 3404
rect 4732 3376 4740 3384
rect 5116 3456 5124 3464
rect 4604 3316 4612 3324
rect 5132 3376 5140 3384
rect 5180 3496 5188 3504
rect 5212 3476 5220 3484
rect 5276 3476 5284 3484
rect 5308 3456 5316 3464
rect 5308 3396 5316 3404
rect 5372 3396 5380 3404
rect 5468 3476 5470 3484
rect 5470 3476 5476 3484
rect 5404 3356 5412 3364
rect 5692 4136 5700 4144
rect 5804 4136 5812 4144
rect 5516 4016 5524 4024
rect 5628 4016 5636 4024
rect 5660 4016 5668 4024
rect 5596 3876 5604 3884
rect 5612 3736 5620 3744
rect 5788 3736 5796 3744
rect 5500 3356 5508 3364
rect 5628 3476 5636 3484
rect 5788 3436 5796 3444
rect 5820 3436 5828 3444
rect 5660 3396 5668 3404
rect 5532 3336 5540 3344
rect 5852 3336 5860 3344
rect 4684 3296 4692 3304
rect 4748 3296 4756 3304
rect 4636 3276 4644 3284
rect 4572 3256 4580 3264
rect 4540 3116 4548 3124
rect 4588 3136 4596 3144
rect 4508 3076 4516 3084
rect 4524 3076 4532 3084
rect 4412 3056 4420 3064
rect 4428 2936 4436 2944
rect 4572 3096 4580 3104
rect 4764 3256 4772 3264
rect 4684 3176 4692 3184
rect 4748 3096 4756 3104
rect 4812 3096 4820 3104
rect 4844 3102 4852 3104
rect 4844 3096 4852 3102
rect 4604 3076 4612 3084
rect 4620 3056 4628 3064
rect 4780 3056 4788 3064
rect 5068 3316 5076 3324
rect 5116 3316 5124 3324
rect 5660 3316 5668 3324
rect 4972 3176 4980 3184
rect 5004 3176 5012 3184
rect 5292 3116 5300 3124
rect 5356 3116 5364 3124
rect 5292 3096 5300 3104
rect 5372 3096 5380 3104
rect 4876 3076 4884 3084
rect 5164 3076 5172 3084
rect 5196 3076 5204 3084
rect 5340 3076 5348 3084
rect 5420 3076 5428 3084
rect 5548 3236 5556 3244
rect 4556 3036 4564 3044
rect 4812 3036 4820 3044
rect 4540 2916 4548 2924
rect 4524 2896 4532 2904
rect 4364 2856 4372 2864
rect 4446 2806 4454 2814
rect 4460 2806 4468 2814
rect 4474 2806 4482 2814
rect 5004 3056 5012 3064
rect 5372 3056 5380 3064
rect 5436 3056 5444 3064
rect 5468 3056 5476 3064
rect 5324 3036 5332 3044
rect 4572 2936 4580 2944
rect 4588 2936 4596 2944
rect 4620 2936 4628 2944
rect 4956 2936 4964 2944
rect 5084 2936 5092 2944
rect 5116 2936 5124 2944
rect 4604 2916 4612 2924
rect 4620 2916 4628 2924
rect 4572 2876 4580 2884
rect 4604 2876 4612 2884
rect 4636 2896 4644 2904
rect 4332 2736 4340 2744
rect 4380 2716 4388 2724
rect 4396 2696 4404 2704
rect 4604 2696 4612 2704
rect 4300 2676 4308 2684
rect 4348 2596 4356 2604
rect 4316 2576 4324 2584
rect 4396 2596 4404 2604
rect 4300 2536 4308 2544
rect 4332 2376 4340 2384
rect 4252 2356 4260 2364
rect 4300 2336 4308 2344
rect 3020 2256 3028 2264
rect 2910 2206 2918 2214
rect 2924 2206 2932 2214
rect 2938 2206 2946 2214
rect 2940 2176 2948 2184
rect 2924 2156 2932 2164
rect 2988 2156 2996 2164
rect 3628 2296 3636 2304
rect 3756 2296 3764 2304
rect 3948 2296 3956 2304
rect 4044 2296 4052 2304
rect 3260 2236 3268 2244
rect 3324 2236 3332 2244
rect 3452 2236 3460 2244
rect 3644 2236 3652 2244
rect 3148 2216 3156 2224
rect 3260 2216 3268 2224
rect 3100 2136 3108 2144
rect 2764 2116 2772 2124
rect 2796 2116 2804 2124
rect 2844 2116 2852 2124
rect 3116 2118 3124 2124
rect 3116 2116 3124 2118
rect 3180 2116 3188 2124
rect 2732 2096 2740 2104
rect 2652 2076 2660 2084
rect 2700 2076 2708 2084
rect 2524 2036 2532 2044
rect 2556 1916 2564 1924
rect 2460 1876 2468 1884
rect 1980 1856 1988 1864
rect 2124 1856 2132 1864
rect 2108 1836 2116 1844
rect 1932 1776 1940 1784
rect 1900 1736 1908 1744
rect 2044 1776 2052 1784
rect 2076 1756 2084 1764
rect 2108 1756 2116 1764
rect 2172 1756 2180 1764
rect 1996 1736 2004 1744
rect 2012 1736 2020 1744
rect 2028 1716 2036 1724
rect 2124 1716 2132 1724
rect 2156 1716 2164 1724
rect 2428 1856 2436 1864
rect 2812 2096 2820 2104
rect 2844 2096 2852 2104
rect 2988 2036 2996 2044
rect 2796 1902 2804 1904
rect 2796 1896 2804 1902
rect 3020 1916 3028 1924
rect 3036 1916 3044 1924
rect 2588 1876 2596 1884
rect 2572 1856 2580 1864
rect 2684 1856 2692 1864
rect 2732 1836 2740 1844
rect 2524 1796 2532 1804
rect 2924 1856 2932 1864
rect 2910 1806 2918 1814
rect 2924 1806 2932 1814
rect 2938 1806 2946 1814
rect 2220 1736 2228 1744
rect 2652 1736 2660 1744
rect 2684 1736 2692 1744
rect 2924 1736 2932 1744
rect 2204 1716 2212 1724
rect 2268 1716 2276 1724
rect 2380 1718 2388 1724
rect 2380 1716 2388 1718
rect 1980 1696 1988 1704
rect 2156 1696 2164 1704
rect 2236 1696 2244 1704
rect 2300 1696 2308 1704
rect 2204 1676 2212 1684
rect 2316 1676 2324 1684
rect 2476 1636 2484 1644
rect 2508 1636 2516 1644
rect 2444 1576 2452 1584
rect 1884 1556 1892 1564
rect 2396 1536 2404 1544
rect 2092 1516 2100 1524
rect 2252 1516 2260 1524
rect 2140 1496 2148 1504
rect 1964 1476 1972 1484
rect 2076 1476 2084 1484
rect 2236 1476 2244 1484
rect 2284 1476 2292 1484
rect 2316 1476 2324 1484
rect 1836 1416 1844 1424
rect 1788 1336 1796 1344
rect 1836 1336 1844 1344
rect 1644 1318 1652 1324
rect 1644 1316 1652 1318
rect 1708 1316 1716 1324
rect 1820 1316 1828 1324
rect 1516 1176 1524 1184
rect 1484 1096 1492 1104
rect 1564 1096 1572 1104
rect 1692 1136 1700 1144
rect 1772 1196 1780 1204
rect 1820 1136 1828 1144
rect 1932 1456 1940 1464
rect 1932 1356 1940 1364
rect 1980 1456 1988 1464
rect 2060 1416 2068 1424
rect 2012 1376 2020 1384
rect 1980 1356 1988 1364
rect 2060 1356 2068 1364
rect 1964 1336 1972 1344
rect 1884 1316 1892 1324
rect 1932 1316 1940 1324
rect 1852 1296 1860 1304
rect 2012 1296 2020 1304
rect 2108 1296 2116 1304
rect 2012 1176 2020 1184
rect 1932 1116 1940 1124
rect 1964 1116 1972 1124
rect 2108 1276 2116 1284
rect 2076 1176 2084 1184
rect 2140 1456 2148 1464
rect 2204 1436 2212 1444
rect 2316 1456 2324 1464
rect 2284 1436 2292 1444
rect 2268 1396 2276 1404
rect 2252 1376 2260 1384
rect 2268 1356 2276 1364
rect 2300 1356 2308 1364
rect 2460 1496 2468 1504
rect 2444 1456 2452 1464
rect 2156 1336 2164 1344
rect 2236 1336 2244 1344
rect 2284 1336 2292 1344
rect 2316 1336 2324 1344
rect 2380 1336 2388 1344
rect 2156 1316 2164 1324
rect 2188 1296 2196 1304
rect 2220 1296 2228 1304
rect 2236 1296 2244 1304
rect 2140 1216 2148 1224
rect 2092 1156 2100 1164
rect 2124 1156 2132 1164
rect 2044 1116 2052 1124
rect 2076 1116 2084 1124
rect 1916 1096 1924 1104
rect 1948 1076 1956 1084
rect 2012 1076 2020 1084
rect 1436 1056 1444 1064
rect 1452 1056 1460 1064
rect 1500 1056 1508 1064
rect 1596 1056 1604 1064
rect 1628 1056 1636 1064
rect 1468 1016 1476 1024
rect 1452 976 1460 984
rect 1628 936 1636 944
rect 1532 916 1540 924
rect 1452 896 1460 904
rect 1500 896 1508 904
rect 1468 876 1476 884
rect 1564 856 1572 864
rect 1420 696 1428 704
rect 1276 596 1284 604
rect 1292 596 1300 604
rect 1260 536 1268 544
rect 1324 576 1332 584
rect 1308 556 1316 564
rect 1052 496 1060 504
rect 764 476 772 484
rect 1004 476 1012 484
rect 876 456 884 464
rect 732 376 740 384
rect 700 336 708 344
rect 764 316 772 324
rect 988 376 996 384
rect 924 316 932 324
rect 812 296 820 304
rect 588 276 596 284
rect 172 256 180 264
rect 284 256 292 264
rect 412 256 420 264
rect 460 256 468 264
rect 572 256 580 264
rect 204 176 212 184
rect 348 196 356 204
rect 652 236 660 244
rect 764 196 772 204
rect 380 176 388 184
rect 1036 336 1044 344
rect 1004 296 1012 304
rect 1244 476 1252 484
rect 1180 316 1188 324
rect 1116 302 1124 304
rect 1116 296 1124 302
rect 892 276 900 284
rect 1004 276 1012 284
rect 1020 236 1028 244
rect 956 176 964 184
rect 172 136 180 144
rect 124 116 132 124
rect 268 116 276 124
rect 92 96 100 104
rect 156 96 164 104
rect 348 96 356 104
rect 508 116 516 124
rect 604 116 612 124
rect 636 118 644 124
rect 636 116 644 118
rect 700 116 708 124
rect 892 116 900 124
rect 988 116 996 124
rect 1148 176 1156 184
rect 1292 496 1300 504
rect 1532 656 1540 664
rect 1436 636 1444 644
rect 1532 636 1540 644
rect 1404 616 1412 624
rect 1468 616 1476 624
rect 1484 616 1492 624
rect 1436 576 1444 584
rect 1468 516 1476 524
rect 1308 336 1316 344
rect 1358 406 1366 414
rect 1372 406 1380 414
rect 1386 406 1394 414
rect 1404 356 1412 364
rect 1324 296 1332 304
rect 1356 296 1364 304
rect 1228 236 1236 244
rect 1292 236 1300 244
rect 1340 236 1348 244
rect 1244 216 1252 224
rect 1500 596 1508 604
rect 1516 556 1524 564
rect 1836 976 1844 984
rect 1756 956 1764 964
rect 1804 956 1812 964
rect 1836 956 1844 964
rect 1868 956 1876 964
rect 1772 916 1780 924
rect 1756 876 1764 884
rect 1740 736 1748 744
rect 1596 702 1604 704
rect 1596 696 1604 702
rect 1644 656 1652 664
rect 1564 596 1572 604
rect 1868 736 1876 744
rect 2012 1036 2020 1044
rect 1964 996 1972 1004
rect 1900 976 1908 984
rect 1964 976 1972 984
rect 2108 1096 2116 1104
rect 2172 1116 2180 1124
rect 2348 1316 2356 1324
rect 2716 1696 2724 1704
rect 2844 1676 2852 1684
rect 2988 1696 2996 1704
rect 3292 2176 3300 2184
rect 3356 2156 3364 2164
rect 3292 2136 3300 2144
rect 3420 2156 3428 2164
rect 4444 2636 4452 2644
rect 4380 2516 4388 2524
rect 4412 2516 4420 2524
rect 4396 2436 4404 2444
rect 4428 2496 4436 2504
rect 4572 2636 4580 2644
rect 4524 2596 4532 2604
rect 4588 2596 4596 2604
rect 4700 2918 4708 2924
rect 4700 2916 4708 2918
rect 4828 2876 4836 2884
rect 4908 2916 4916 2924
rect 4940 2916 4948 2924
rect 4796 2736 4804 2744
rect 4844 2736 4852 2744
rect 4668 2676 4676 2684
rect 4508 2516 4516 2524
rect 4620 2536 4628 2544
rect 4684 2536 4692 2544
rect 4540 2496 4548 2504
rect 4524 2476 4532 2484
rect 4556 2476 4564 2484
rect 4604 2476 4612 2484
rect 4492 2456 4500 2464
rect 4508 2416 4516 2424
rect 4446 2406 4454 2414
rect 4460 2406 4468 2414
rect 4474 2406 4482 2414
rect 4556 2396 4564 2404
rect 4668 2516 4676 2524
rect 4684 2496 4692 2504
rect 4716 2516 4724 2524
rect 4748 2516 4756 2524
rect 4684 2456 4692 2464
rect 4668 2396 4676 2404
rect 4652 2376 4660 2384
rect 4620 2356 4628 2364
rect 4428 2336 4436 2344
rect 4556 2336 4564 2344
rect 4380 2316 4388 2324
rect 4364 2296 4372 2304
rect 4348 2256 4356 2264
rect 4284 2236 4292 2244
rect 3708 2176 3716 2184
rect 3484 2136 3492 2144
rect 3660 2136 3668 2144
rect 3388 2116 3396 2124
rect 3804 2156 3812 2164
rect 3932 2156 3940 2164
rect 4428 2316 4436 2324
rect 4524 2316 4532 2324
rect 4588 2316 4596 2324
rect 4652 2316 4660 2324
rect 4492 2296 4500 2304
rect 4444 2256 4452 2264
rect 4428 2196 4436 2204
rect 3756 2136 3764 2144
rect 3772 2116 3780 2124
rect 3068 1936 3076 1944
rect 3212 1936 3220 1944
rect 3116 1916 3124 1924
rect 3084 1876 3092 1884
rect 3100 1856 3108 1864
rect 3132 1856 3140 1864
rect 3084 1776 3092 1784
rect 3324 1876 3332 1884
rect 3148 1836 3156 1844
rect 3132 1776 3140 1784
rect 3228 1856 3236 1864
rect 3324 1856 3332 1864
rect 3260 1796 3268 1804
rect 3356 1836 3364 1844
rect 3212 1756 3220 1764
rect 3324 1756 3332 1764
rect 3244 1736 3252 1744
rect 3196 1716 3204 1724
rect 3180 1696 3188 1704
rect 3212 1696 3220 1704
rect 3260 1696 3268 1704
rect 2956 1656 2964 1664
rect 2988 1536 2996 1544
rect 2524 1516 2532 1524
rect 2556 1496 2564 1504
rect 2636 1496 2644 1504
rect 2668 1496 2676 1504
rect 2572 1476 2580 1484
rect 2812 1496 2820 1504
rect 2588 1456 2596 1464
rect 2636 1456 2644 1464
rect 2588 1436 2596 1444
rect 2652 1436 2660 1444
rect 2508 1356 2516 1364
rect 2556 1336 2564 1344
rect 2652 1336 2660 1344
rect 2444 1316 2452 1324
rect 2476 1316 2484 1324
rect 2316 1296 2324 1304
rect 2268 1216 2276 1224
rect 2268 1176 2276 1184
rect 2284 1176 2292 1184
rect 2236 1096 2244 1104
rect 2044 1076 2052 1084
rect 2092 1076 2100 1084
rect 2028 976 2036 984
rect 1948 936 1956 944
rect 2012 936 2020 944
rect 2028 936 2036 944
rect 1980 916 1988 924
rect 1948 896 1956 904
rect 1900 816 1908 824
rect 1820 696 1828 704
rect 1740 676 1748 684
rect 1804 656 1812 664
rect 1884 696 1892 704
rect 1868 676 1876 684
rect 1932 696 1940 704
rect 2124 996 2132 1004
rect 2076 936 2084 944
rect 2188 1036 2196 1044
rect 2204 1016 2212 1024
rect 2204 996 2212 1004
rect 2188 976 2196 984
rect 2172 936 2180 944
rect 2156 896 2164 904
rect 2028 876 2036 884
rect 1996 836 2004 844
rect 1964 676 1972 684
rect 1980 656 1988 664
rect 1724 636 1732 644
rect 1836 636 1844 644
rect 1916 636 1924 644
rect 1964 636 1972 644
rect 1660 616 1668 624
rect 1788 616 1796 624
rect 1660 596 1668 604
rect 1756 536 1764 544
rect 1724 516 1732 524
rect 1820 518 1828 524
rect 1820 516 1828 518
rect 1564 456 1572 464
rect 1740 456 1748 464
rect 1532 416 1540 424
rect 1516 356 1524 364
rect 1484 316 1492 324
rect 1580 376 1588 384
rect 1644 376 1652 384
rect 1580 336 1588 344
rect 1708 316 1716 324
rect 1420 276 1428 284
rect 1532 256 1540 264
rect 1420 216 1428 224
rect 1404 176 1412 184
rect 1484 176 1492 184
rect 1612 276 1620 284
rect 1628 276 1636 284
rect 1676 296 1684 304
rect 1724 296 1732 304
rect 1596 216 1604 224
rect 1516 156 1524 164
rect 1548 156 1556 164
rect 1596 156 1604 164
rect 1644 156 1652 164
rect 1772 436 1780 444
rect 1756 396 1764 404
rect 1724 216 1732 224
rect 1708 156 1716 164
rect 2108 716 2116 724
rect 2060 696 2068 704
rect 2188 856 2196 864
rect 2172 816 2180 824
rect 2236 1076 2244 1084
rect 2252 1076 2260 1084
rect 2428 1116 2436 1124
rect 2460 1276 2468 1284
rect 2716 1476 2724 1484
rect 2700 1456 2708 1464
rect 2524 1296 2532 1304
rect 2684 1296 2692 1304
rect 2716 1296 2724 1304
rect 2524 1276 2532 1284
rect 2508 1216 2516 1224
rect 2700 1216 2708 1224
rect 2652 1176 2660 1184
rect 2652 1116 2660 1124
rect 2412 1096 2420 1104
rect 2332 1076 2340 1084
rect 2396 1076 2404 1084
rect 2236 1056 2244 1064
rect 2300 1056 2308 1064
rect 2348 1036 2356 1044
rect 2300 976 2308 984
rect 2332 976 2340 984
rect 2428 1036 2436 1044
rect 2364 936 2372 944
rect 2556 1076 2564 1084
rect 2572 1036 2580 1044
rect 2588 1036 2596 1044
rect 2684 1096 2692 1104
rect 2636 1076 2644 1084
rect 2604 1016 2612 1024
rect 2652 1016 2660 1024
rect 2748 1456 2756 1464
rect 2796 1436 2804 1444
rect 2876 1436 2884 1444
rect 2780 1416 2788 1424
rect 2764 1376 2772 1384
rect 2748 1216 2756 1224
rect 2764 1196 2772 1204
rect 2732 1156 2740 1164
rect 2780 1116 2788 1124
rect 2910 1406 2918 1414
rect 2924 1406 2932 1414
rect 2938 1406 2946 1414
rect 2812 1376 2820 1384
rect 2956 1356 2964 1364
rect 3180 1502 3188 1504
rect 3180 1496 3188 1502
rect 3116 1416 3124 1424
rect 3372 1716 3380 1724
rect 3420 1876 3428 1884
rect 3804 2096 3812 2104
rect 3708 2076 3716 2084
rect 3964 2116 3972 2124
rect 3996 2116 4004 2124
rect 3996 2096 4004 2104
rect 3964 2076 3972 2084
rect 4124 2116 4132 2124
rect 4156 2116 4164 2124
rect 4108 2076 4116 2084
rect 4012 1976 4020 1984
rect 4092 1976 4100 1984
rect 3724 1896 3732 1904
rect 3772 1896 3780 1904
rect 3820 1896 3828 1904
rect 3852 1896 3860 1904
rect 3932 1896 3940 1904
rect 3548 1876 3556 1884
rect 3436 1856 3444 1864
rect 3436 1796 3444 1804
rect 3404 1756 3412 1764
rect 3516 1836 3524 1844
rect 3612 1796 3620 1804
rect 3788 1856 3796 1864
rect 3740 1796 3748 1804
rect 3884 1876 3892 1884
rect 3916 1856 3924 1864
rect 3916 1816 3924 1824
rect 3740 1776 3748 1784
rect 3900 1776 3908 1784
rect 3452 1756 3460 1764
rect 3628 1756 3636 1764
rect 3484 1736 3492 1744
rect 3564 1736 3572 1744
rect 3612 1736 3620 1744
rect 3660 1736 3668 1744
rect 3532 1716 3540 1724
rect 3644 1716 3652 1724
rect 3356 1696 3364 1704
rect 3420 1696 3428 1704
rect 3484 1696 3492 1704
rect 3516 1696 3524 1704
rect 3612 1696 3620 1704
rect 3308 1676 3316 1684
rect 3468 1676 3476 1684
rect 3564 1656 3572 1664
rect 3244 1556 3252 1564
rect 2812 1336 2820 1344
rect 2748 1096 2756 1104
rect 2716 1076 2724 1084
rect 2684 976 2692 984
rect 2460 956 2468 964
rect 2556 936 2564 944
rect 2668 936 2676 944
rect 2332 916 2340 924
rect 2412 916 2420 924
rect 2236 896 2244 904
rect 2220 876 2228 884
rect 2252 836 2260 844
rect 2204 736 2212 744
rect 2348 896 2356 904
rect 2396 896 2404 904
rect 2284 736 2292 744
rect 2188 696 2196 704
rect 2028 676 2036 684
rect 2236 676 2244 684
rect 2268 676 2276 684
rect 2284 676 2292 684
rect 2060 656 2068 664
rect 2140 656 2148 664
rect 2156 656 2164 664
rect 2124 636 2132 644
rect 2060 616 2068 624
rect 2204 636 2212 644
rect 2028 576 2036 584
rect 2268 636 2276 644
rect 2156 576 2164 584
rect 2332 576 2340 584
rect 2396 676 2404 684
rect 2236 556 2244 564
rect 1980 536 1988 544
rect 2092 536 2100 544
rect 2204 536 2212 544
rect 1932 476 1940 484
rect 1836 396 1844 404
rect 2172 516 2180 524
rect 1996 456 2004 464
rect 2076 456 2084 464
rect 2108 456 2116 464
rect 1980 416 1988 424
rect 1996 316 2004 324
rect 2044 316 2052 324
rect 1836 296 1844 304
rect 1964 296 1972 304
rect 1980 276 1988 284
rect 2060 276 2068 284
rect 1820 256 1828 264
rect 1788 216 1796 224
rect 1852 216 1860 224
rect 1772 196 1780 204
rect 1740 176 1748 184
rect 1500 136 1508 144
rect 1612 136 1620 144
rect 1964 256 1972 264
rect 1932 216 1940 224
rect 1884 196 1892 204
rect 1868 176 1876 184
rect 1916 176 1924 184
rect 1996 176 2004 184
rect 1948 156 1956 164
rect 1820 136 1828 144
rect 1788 116 1796 124
rect 1996 116 2004 124
rect 828 96 836 104
rect 2028 196 2036 204
rect 2060 116 2068 124
rect 2188 376 2196 384
rect 2172 356 2180 364
rect 2188 356 2196 364
rect 2156 316 2164 324
rect 2108 296 2116 304
rect 2140 276 2148 284
rect 2092 256 2100 264
rect 2188 316 2196 324
rect 2188 296 2196 304
rect 2300 516 2308 524
rect 2348 516 2356 524
rect 2380 636 2388 644
rect 2444 916 2452 924
rect 2476 916 2484 924
rect 2540 896 2548 904
rect 2604 896 2612 904
rect 2572 876 2580 884
rect 2492 856 2500 864
rect 2444 736 2452 744
rect 2700 736 2708 744
rect 2444 716 2452 724
rect 2508 716 2516 724
rect 2540 716 2548 724
rect 2604 716 2612 724
rect 2460 696 2468 704
rect 2460 656 2468 664
rect 2732 1056 2740 1064
rect 2764 1076 2772 1084
rect 2940 1336 2948 1344
rect 3052 1336 3060 1344
rect 2844 1316 2852 1324
rect 2988 1316 2996 1324
rect 2892 1296 2900 1304
rect 2892 1136 2900 1144
rect 2828 1096 2836 1104
rect 2972 1096 2980 1104
rect 2812 1056 2820 1064
rect 2828 1036 2836 1044
rect 2924 1036 2932 1044
rect 2876 1016 2884 1024
rect 2910 1006 2918 1014
rect 2924 1006 2932 1014
rect 2938 1006 2946 1014
rect 2828 956 2836 964
rect 3116 1276 3124 1284
rect 3068 1256 3076 1264
rect 3020 1236 3028 1244
rect 3132 1236 3140 1244
rect 3100 1216 3108 1224
rect 3036 976 3044 984
rect 3004 956 3012 964
rect 2924 936 2932 944
rect 2988 936 2996 944
rect 3020 936 3028 944
rect 2764 876 2772 884
rect 2828 876 2836 884
rect 2956 916 2964 924
rect 3020 916 3028 924
rect 2908 876 2916 884
rect 2844 716 2852 724
rect 2860 716 2868 724
rect 2540 696 2548 704
rect 2588 696 2596 704
rect 2492 676 2500 684
rect 2684 676 2692 684
rect 2556 656 2564 664
rect 2636 656 2644 664
rect 2444 636 2452 644
rect 2476 636 2484 644
rect 2620 636 2628 644
rect 2396 576 2404 584
rect 2428 576 2436 584
rect 2412 556 2420 564
rect 3068 936 3076 944
rect 3724 1736 3732 1744
rect 3772 1736 3780 1744
rect 3644 1536 3652 1544
rect 3692 1676 3700 1684
rect 3708 1556 3716 1564
rect 3692 1536 3700 1544
rect 3324 1516 3332 1524
rect 3516 1516 3524 1524
rect 3484 1496 3492 1504
rect 3308 1456 3316 1464
rect 3372 1456 3380 1464
rect 3468 1456 3476 1464
rect 3260 1416 3268 1424
rect 3644 1496 3652 1504
rect 3676 1496 3684 1504
rect 3548 1476 3556 1484
rect 3484 1416 3492 1424
rect 3516 1416 3524 1424
rect 3436 1376 3444 1384
rect 3580 1456 3588 1464
rect 3628 1456 3636 1464
rect 3564 1436 3572 1444
rect 3580 1356 3588 1364
rect 3628 1416 3636 1424
rect 3356 1336 3364 1344
rect 3484 1336 3492 1344
rect 3612 1336 3620 1344
rect 3180 1316 3188 1324
rect 3436 1296 3444 1304
rect 3452 1276 3460 1284
rect 3324 1256 3332 1264
rect 3548 1316 3556 1324
rect 3564 1276 3572 1284
rect 3324 1136 3332 1144
rect 3148 1076 3156 1084
rect 3292 1076 3300 1084
rect 3260 1016 3268 1024
rect 3228 916 3236 924
rect 3516 1096 3524 1104
rect 3564 1036 3572 1044
rect 3564 1016 3572 1024
rect 3564 956 3572 964
rect 3820 1716 3828 1724
rect 3868 1716 3876 1724
rect 3900 1716 3908 1724
rect 3740 1696 3748 1704
rect 4076 1896 4084 1904
rect 4060 1876 4068 1884
rect 3996 1816 4004 1824
rect 4012 1776 4020 1784
rect 4044 1776 4052 1784
rect 3964 1756 3972 1764
rect 4012 1716 4020 1724
rect 4060 1716 4068 1724
rect 3804 1696 3812 1704
rect 3884 1696 3892 1704
rect 3932 1696 3940 1704
rect 3964 1696 3972 1704
rect 3996 1696 4004 1704
rect 3772 1676 3780 1684
rect 3756 1656 3764 1664
rect 3756 1576 3764 1584
rect 3756 1556 3764 1564
rect 3740 1536 3748 1544
rect 3740 1516 3748 1524
rect 3724 1476 3732 1484
rect 3756 1476 3764 1484
rect 3740 1456 3748 1464
rect 3852 1676 3860 1684
rect 3916 1676 3924 1684
rect 4060 1676 4068 1684
rect 3980 1596 3988 1604
rect 4028 1596 4036 1604
rect 3980 1576 3988 1584
rect 3804 1556 3812 1564
rect 3804 1536 3812 1544
rect 3852 1516 3860 1524
rect 3804 1476 3812 1484
rect 3884 1496 3892 1504
rect 3820 1456 3828 1464
rect 3868 1476 3876 1484
rect 3900 1476 3908 1484
rect 3740 1396 3748 1404
rect 3644 1376 3652 1384
rect 3692 1376 3700 1384
rect 3708 1376 3716 1384
rect 3676 1336 3684 1344
rect 3724 1336 3732 1344
rect 3660 1276 3668 1284
rect 3628 1136 3636 1144
rect 3676 1116 3684 1124
rect 3708 1116 3716 1124
rect 3596 1096 3604 1104
rect 3660 1076 3668 1084
rect 3804 1436 3812 1444
rect 3852 1436 3860 1444
rect 3836 1376 3844 1384
rect 3868 1376 3876 1384
rect 3772 1356 3780 1364
rect 3788 1356 3796 1364
rect 3868 1356 3876 1364
rect 3884 1356 3892 1364
rect 3852 1316 3860 1324
rect 3804 1296 3812 1304
rect 3804 1176 3812 1184
rect 3756 1096 3764 1104
rect 3788 1056 3796 1064
rect 3788 1016 3796 1024
rect 3660 976 3668 984
rect 3788 956 3796 964
rect 3580 936 3588 944
rect 3164 896 3172 904
rect 3420 916 3428 924
rect 3676 916 3684 924
rect 3356 876 3364 884
rect 3772 876 3780 884
rect 3164 736 3172 744
rect 3292 736 3300 744
rect 3068 716 3076 724
rect 3084 716 3092 724
rect 2732 636 2740 644
rect 2732 596 2740 604
rect 2604 576 2612 584
rect 2668 576 2676 584
rect 2508 536 2516 544
rect 2556 536 2564 544
rect 2588 536 2596 544
rect 2524 516 2532 524
rect 2588 516 2596 524
rect 2556 496 2564 504
rect 2524 436 2532 444
rect 2540 396 2548 404
rect 2476 376 2484 384
rect 2332 356 2340 364
rect 2428 336 2436 344
rect 2268 316 2276 324
rect 2204 276 2212 284
rect 2172 256 2180 264
rect 2188 256 2196 264
rect 2172 216 2180 224
rect 2108 176 2116 184
rect 2156 176 2164 184
rect 2300 236 2308 244
rect 2316 236 2324 244
rect 2204 176 2212 184
rect 2252 176 2260 184
rect 2124 136 2132 144
rect 2236 136 2244 144
rect 2348 316 2356 324
rect 2460 316 2468 324
rect 2508 316 2516 324
rect 2572 316 2580 324
rect 2588 316 2596 324
rect 2492 296 2500 304
rect 2556 276 2564 284
rect 2332 216 2340 224
rect 2396 216 2404 224
rect 2444 216 2452 224
rect 2492 196 2500 204
rect 2444 176 2452 184
rect 2460 176 2468 184
rect 2540 216 2548 224
rect 2540 176 2548 184
rect 2316 136 2324 144
rect 2444 136 2452 144
rect 2460 136 2468 144
rect 2476 136 2484 144
rect 2540 136 2548 144
rect 76 76 84 84
rect 108 76 116 84
rect 236 76 244 84
rect 444 76 452 84
rect 2012 76 2020 84
rect 2092 76 2100 84
rect 2252 76 2260 84
rect 2268 76 2276 84
rect 2828 676 2836 684
rect 2876 696 2884 704
rect 2988 696 2996 704
rect 3036 696 3044 704
rect 3084 696 3092 704
rect 3116 696 3124 704
rect 2828 656 2836 664
rect 2844 656 2852 664
rect 2812 596 2820 604
rect 2780 576 2788 584
rect 2764 556 2772 564
rect 2860 636 2868 644
rect 2910 606 2918 614
rect 2924 606 2932 614
rect 2938 606 2946 614
rect 2876 596 2884 604
rect 3084 676 3092 684
rect 3036 656 3044 664
rect 3068 656 3076 664
rect 3228 696 3236 704
rect 3292 696 3300 704
rect 3196 656 3204 664
rect 3212 656 3220 664
rect 3276 656 3284 664
rect 3020 636 3028 644
rect 3036 636 3044 644
rect 3100 636 3108 644
rect 3244 636 3252 644
rect 3004 556 3012 564
rect 3068 556 3076 564
rect 3164 556 3172 564
rect 3260 556 3268 564
rect 2828 536 2836 544
rect 2924 536 2932 544
rect 3004 536 3012 544
rect 3052 536 3060 544
rect 2636 516 2644 524
rect 2764 516 2772 524
rect 2828 516 2836 524
rect 2780 496 2788 504
rect 2652 476 2660 484
rect 2684 476 2692 484
rect 2652 436 2660 444
rect 2700 456 2708 464
rect 2780 456 2788 464
rect 2668 376 2676 384
rect 2684 356 2692 364
rect 2620 336 2628 344
rect 2876 416 2884 424
rect 2972 496 2980 504
rect 3084 536 3092 544
rect 3036 376 3044 384
rect 2844 336 2852 344
rect 2940 336 2948 344
rect 2988 336 2996 344
rect 2860 316 2868 324
rect 2908 316 2916 324
rect 2620 296 2628 304
rect 2732 296 2740 304
rect 2812 296 2820 304
rect 2956 296 2964 304
rect 2668 276 2676 284
rect 2780 256 2788 264
rect 2652 236 2660 244
rect 2764 236 2772 244
rect 2652 196 2660 204
rect 2636 156 2644 164
rect 2604 136 2612 144
rect 2860 276 2868 284
rect 2972 276 2980 284
rect 2910 206 2918 214
rect 2924 206 2932 214
rect 2938 206 2946 214
rect 2876 176 2884 184
rect 2892 176 2900 184
rect 2748 156 2756 164
rect 2764 156 2772 164
rect 2972 156 2980 164
rect 3020 316 3028 324
rect 3148 536 3156 544
rect 3228 536 3236 544
rect 3132 456 3140 464
rect 3212 516 3220 524
rect 3180 416 3188 424
rect 3164 396 3172 404
rect 3180 396 3188 404
rect 3132 336 3140 344
rect 3116 296 3124 304
rect 3612 776 3620 784
rect 3676 716 3684 724
rect 3324 676 3332 684
rect 3340 636 3348 644
rect 3820 1056 3828 1064
rect 3820 1036 3828 1044
rect 3820 996 3828 1004
rect 3900 1336 3908 1344
rect 4044 1536 4052 1544
rect 4140 1796 4148 1804
rect 4108 1716 4116 1724
rect 3948 1456 3956 1464
rect 4012 1436 4020 1444
rect 4044 1376 4052 1384
rect 3996 1356 4004 1364
rect 3980 1336 3988 1344
rect 4092 1496 4100 1504
rect 4332 2116 4340 2124
rect 4188 2096 4196 2104
rect 4316 2076 4324 2084
rect 4364 2036 4372 2044
rect 4396 2116 4404 2124
rect 4636 2276 4644 2284
rect 4524 2196 4532 2204
rect 4444 2096 4452 2104
rect 4396 2036 4404 2044
rect 4572 2256 4580 2264
rect 4588 2256 4596 2264
rect 4588 2196 4596 2204
rect 4572 2156 4580 2164
rect 4572 2136 4580 2144
rect 4300 1896 4308 1904
rect 4332 1902 4340 1904
rect 4332 1896 4340 1902
rect 4380 1896 4388 1904
rect 4204 1836 4212 1844
rect 4252 1816 4260 1824
rect 4188 1736 4196 1744
rect 4204 1716 4212 1724
rect 4172 1576 4180 1584
rect 4204 1556 4212 1564
rect 4156 1516 4164 1524
rect 4124 1496 4132 1504
rect 4108 1476 4116 1484
rect 4108 1456 4116 1464
rect 4108 1436 4116 1444
rect 4252 1476 4260 1484
rect 4204 1456 4212 1464
rect 4140 1416 4148 1424
rect 4284 1496 4292 1504
rect 4284 1476 4292 1484
rect 4284 1436 4292 1444
rect 4268 1396 4276 1404
rect 4316 1696 4324 1704
rect 4316 1456 4324 1464
rect 4332 1436 4340 1444
rect 4316 1416 4324 1424
rect 4268 1376 4276 1384
rect 4300 1376 4308 1384
rect 3996 1316 4004 1324
rect 4172 1316 4180 1324
rect 3932 1276 3940 1284
rect 3964 1276 3972 1284
rect 3884 1136 3892 1144
rect 3948 1136 3956 1144
rect 3900 1116 3908 1124
rect 3868 1076 3876 1084
rect 4076 1276 4084 1284
rect 3996 1196 4004 1204
rect 4060 1196 4068 1204
rect 3964 1076 3972 1084
rect 4156 1296 4164 1304
rect 4204 1336 4212 1344
rect 4300 1316 4308 1324
rect 4348 1316 4356 1324
rect 4188 1256 4196 1264
rect 4140 1156 4148 1164
rect 4172 1156 4180 1164
rect 4060 1136 4068 1144
rect 4076 1116 4084 1124
rect 4124 1116 4132 1124
rect 3964 1016 3972 1024
rect 3980 1016 3988 1024
rect 3884 976 3892 984
rect 3948 976 3956 984
rect 3852 956 3860 964
rect 3820 896 3828 904
rect 3900 956 3908 964
rect 3900 916 3908 924
rect 3916 916 3924 924
rect 3852 896 3860 904
rect 3980 936 3988 944
rect 4060 1016 4068 1024
rect 4124 1096 4132 1104
rect 4172 1096 4180 1104
rect 4446 2006 4454 2014
rect 4460 2006 4468 2014
rect 4474 2006 4482 2014
rect 4524 1916 4532 1924
rect 4540 1896 4548 1904
rect 4524 1876 4532 1884
rect 4652 2156 4660 2164
rect 4652 2136 4660 2144
rect 4588 2116 4596 2124
rect 4636 2096 4644 2104
rect 4620 1996 4628 2004
rect 4620 1896 4628 1904
rect 4700 2316 4708 2324
rect 4700 2196 4708 2204
rect 4668 2076 4676 2084
rect 4668 2056 4676 2064
rect 4652 2036 4660 2044
rect 4700 2036 4708 2044
rect 4684 1996 4692 2004
rect 4828 2716 4836 2724
rect 4892 2716 4900 2724
rect 4876 2616 4884 2624
rect 4812 2596 4820 2604
rect 4956 2716 4964 2724
rect 5148 2876 5156 2884
rect 5276 2876 5284 2884
rect 5212 2716 5220 2724
rect 4956 2696 4964 2704
rect 5116 2696 5124 2704
rect 5212 2696 5220 2704
rect 4860 2516 4868 2524
rect 4860 2496 4868 2504
rect 4892 2496 4900 2504
rect 4828 2436 4836 2444
rect 4748 2416 4756 2424
rect 4764 2336 4772 2344
rect 4732 2236 4740 2244
rect 4860 2316 4868 2324
rect 5020 2616 5028 2624
rect 4940 2596 4948 2604
rect 5276 2716 5284 2724
rect 5516 3076 5524 3084
rect 5500 3036 5508 3044
rect 5372 2956 5380 2964
rect 5548 2936 5556 2944
rect 5628 3116 5636 3124
rect 5692 3116 5700 3124
rect 5660 3076 5668 3084
rect 5772 3296 5780 3304
rect 5788 3056 5796 3064
rect 5820 3036 5828 3044
rect 5692 2956 5700 2964
rect 5740 2956 5748 2964
rect 5724 2936 5732 2944
rect 5788 2936 5796 2944
rect 5644 2916 5652 2924
rect 5740 2916 5748 2924
rect 5644 2896 5652 2904
rect 5692 2896 5700 2904
rect 5852 2896 5860 2904
rect 5804 2876 5812 2884
rect 5612 2776 5620 2784
rect 5596 2716 5604 2724
rect 5660 2716 5668 2724
rect 5468 2702 5476 2704
rect 5468 2696 5476 2702
rect 5852 2696 5860 2704
rect 5340 2676 5348 2684
rect 5436 2676 5444 2684
rect 5628 2676 5636 2684
rect 5404 2636 5412 2644
rect 5292 2576 5300 2584
rect 4988 2556 4996 2564
rect 5020 2556 5028 2564
rect 5564 2616 5572 2624
rect 5020 2536 5028 2544
rect 5132 2536 5140 2544
rect 5148 2516 5156 2524
rect 4956 2316 4964 2324
rect 4988 2336 4996 2344
rect 4972 2296 4980 2304
rect 4796 2256 4804 2264
rect 5084 2316 5092 2324
rect 5148 2316 5156 2324
rect 5212 2296 5220 2304
rect 5116 2276 5124 2284
rect 4956 2256 4964 2264
rect 5020 2256 5028 2264
rect 4860 2236 4868 2244
rect 4892 2236 4900 2244
rect 4748 2216 4756 2224
rect 4764 2156 4772 2164
rect 4940 2196 4948 2204
rect 4876 2156 4884 2164
rect 4908 2156 4916 2164
rect 4828 2136 4836 2144
rect 4892 2136 4900 2144
rect 4748 2116 4756 2124
rect 4764 2116 4772 2124
rect 4924 2116 4932 2124
rect 4828 2096 4836 2104
rect 4860 2096 4868 2104
rect 4748 2076 4756 2084
rect 4796 2076 4804 2084
rect 4748 2036 4756 2044
rect 4780 1896 4788 1904
rect 4636 1876 4644 1884
rect 4764 1876 4772 1884
rect 4604 1856 4612 1864
rect 4652 1856 4660 1864
rect 4764 1856 4772 1864
rect 4748 1836 4756 1844
rect 4588 1816 4596 1824
rect 4572 1796 4580 1804
rect 4764 1796 4772 1804
rect 4812 2056 4820 2064
rect 4812 1996 4820 2004
rect 4860 1996 4868 2004
rect 4876 1896 4884 1904
rect 4812 1876 4820 1884
rect 5100 2236 5108 2244
rect 4972 2216 4980 2224
rect 5324 2336 5332 2344
rect 5244 2236 5252 2244
rect 4988 2156 4996 2164
rect 5244 2156 5252 2164
rect 5292 2156 5300 2164
rect 4956 2136 4964 2144
rect 4972 2136 4980 2144
rect 5004 2136 5012 2144
rect 5132 2136 5140 2144
rect 5308 2136 5316 2144
rect 4972 2116 4980 2124
rect 5020 2076 5028 2084
rect 5052 2076 5060 2084
rect 4988 1996 4996 2004
rect 5212 2116 5220 2124
rect 5276 2116 5284 2124
rect 5116 1916 5124 1924
rect 5148 1916 5156 1924
rect 5180 1916 5188 1924
rect 5196 1916 5204 1924
rect 5164 1896 5172 1904
rect 4924 1876 4932 1884
rect 4940 1876 4948 1884
rect 4972 1876 4980 1884
rect 5084 1876 5092 1884
rect 4940 1856 4948 1864
rect 4844 1836 4852 1844
rect 4892 1836 4900 1844
rect 4924 1836 4932 1844
rect 4860 1816 4868 1824
rect 5132 1856 5140 1864
rect 4988 1816 4996 1824
rect 5084 1816 5092 1824
rect 5036 1796 5044 1804
rect 5004 1776 5012 1784
rect 5020 1756 5028 1764
rect 4460 1736 4468 1744
rect 4908 1736 4916 1744
rect 4524 1716 4532 1724
rect 4446 1606 4454 1614
rect 4460 1606 4468 1614
rect 4474 1606 4482 1614
rect 4620 1718 4628 1724
rect 4620 1716 4628 1718
rect 4476 1576 4484 1584
rect 4556 1576 4564 1584
rect 4636 1556 4644 1564
rect 4396 1536 4404 1544
rect 4508 1516 4516 1524
rect 4620 1516 4628 1524
rect 4588 1496 4596 1504
rect 4444 1456 4452 1464
rect 4380 1396 4388 1404
rect 4556 1416 4564 1424
rect 4620 1416 4628 1424
rect 4508 1396 4516 1404
rect 4444 1376 4452 1384
rect 4492 1356 4500 1364
rect 4348 1276 4356 1284
rect 4364 1276 4372 1284
rect 4332 1196 4340 1204
rect 4316 1176 4324 1184
rect 4316 1156 4324 1164
rect 4236 1096 4244 1104
rect 4412 1316 4420 1324
rect 4446 1206 4454 1214
rect 4460 1206 4468 1214
rect 4474 1206 4482 1214
rect 4492 1176 4500 1184
rect 4364 1102 4372 1104
rect 4364 1096 4372 1102
rect 4380 1096 4388 1104
rect 4108 1076 4116 1084
rect 4140 1076 4148 1084
rect 4172 1036 4180 1044
rect 4092 956 4100 964
rect 4076 916 4084 924
rect 4300 1056 4308 1064
rect 4236 976 4244 984
rect 4268 956 4276 964
rect 4188 936 4196 944
rect 4300 936 4308 944
rect 4220 916 4228 924
rect 4028 896 4036 904
rect 4140 896 4148 904
rect 4188 896 4196 904
rect 4220 896 4228 904
rect 3916 876 3924 884
rect 3948 876 3956 884
rect 4012 876 4020 884
rect 3996 716 4004 724
rect 4060 716 4068 724
rect 3532 676 3540 684
rect 3644 676 3652 684
rect 3804 676 3812 684
rect 3484 616 3492 624
rect 3420 596 3428 604
rect 3388 556 3396 564
rect 3484 556 3492 564
rect 3404 536 3412 544
rect 3692 556 3700 564
rect 3804 596 3812 604
rect 3756 576 3764 584
rect 3308 516 3316 524
rect 3324 516 3332 524
rect 3388 516 3396 524
rect 3468 516 3476 524
rect 3276 476 3284 484
rect 3292 396 3300 404
rect 3948 696 3956 704
rect 3900 676 3908 684
rect 3900 596 3908 604
rect 4124 876 4132 884
rect 4092 816 4100 824
rect 4076 696 4084 704
rect 3964 676 3972 684
rect 4012 596 4020 604
rect 3852 556 3860 564
rect 3964 556 3972 564
rect 4252 896 4260 904
rect 4364 876 4372 884
rect 4332 816 4340 824
rect 4236 776 4244 784
rect 4268 776 4276 784
rect 4140 756 4148 764
rect 4236 736 4244 744
rect 4140 716 4148 724
rect 4108 696 4116 704
rect 4540 1376 4548 1384
rect 4572 1316 4580 1324
rect 4668 1496 4676 1504
rect 4732 1502 4740 1504
rect 4732 1496 4740 1502
rect 4780 1496 4788 1504
rect 4668 1476 4676 1484
rect 4748 1476 4756 1484
rect 4988 1696 4996 1704
rect 4860 1576 4868 1584
rect 4908 1576 4916 1584
rect 4876 1496 4884 1504
rect 4668 1356 4676 1364
rect 5068 1776 5076 1784
rect 5164 1836 5172 1844
rect 5276 1996 5284 2004
rect 5340 2116 5348 2124
rect 5388 2302 5396 2304
rect 5388 2296 5396 2302
rect 5772 2636 5780 2644
rect 5596 2496 5604 2504
rect 5548 2476 5556 2484
rect 5660 2476 5668 2484
rect 5516 2316 5524 2324
rect 5580 2316 5588 2324
rect 5852 2536 5860 2544
rect 5852 2376 5860 2384
rect 5756 2296 5764 2304
rect 5548 2276 5556 2284
rect 5372 2136 5380 2144
rect 5388 2096 5396 2104
rect 5420 2096 5428 2104
rect 5484 2076 5492 2084
rect 5612 2076 5620 2084
rect 5324 1876 5332 1884
rect 5212 1856 5220 1864
rect 5244 1856 5252 1864
rect 5260 1856 5268 1864
rect 5100 1756 5108 1764
rect 5116 1756 5124 1764
rect 5148 1756 5156 1764
rect 5180 1756 5188 1764
rect 5036 1716 5044 1724
rect 5084 1716 5092 1724
rect 5052 1696 5060 1704
rect 5052 1556 5060 1564
rect 4988 1476 4996 1484
rect 5004 1476 5012 1484
rect 4684 1336 4692 1344
rect 4908 1336 4916 1344
rect 4716 1316 4724 1324
rect 4748 1316 4756 1324
rect 4652 1296 4660 1304
rect 4716 1296 4724 1304
rect 4764 1276 4772 1284
rect 4796 1156 4804 1164
rect 4732 1136 4740 1144
rect 4588 1116 4596 1124
rect 4620 1096 4628 1104
rect 4732 1096 4740 1104
rect 4620 1056 4628 1064
rect 4860 1116 4868 1124
rect 4668 1036 4676 1044
rect 4620 1016 4628 1024
rect 4524 996 4532 1004
rect 4588 996 4596 1004
rect 4668 996 4676 1004
rect 4652 956 4660 964
rect 4780 1056 4788 1064
rect 4812 1036 4820 1044
rect 4796 996 4804 1004
rect 4684 976 4692 984
rect 4780 976 4788 984
rect 4796 956 4804 964
rect 4446 806 4454 814
rect 4460 806 4468 814
rect 4474 806 4482 814
rect 4380 736 4388 744
rect 4284 716 4292 724
rect 4268 656 4276 664
rect 4124 616 4132 624
rect 4204 636 4212 644
rect 4220 596 4228 604
rect 4236 596 4244 604
rect 4124 556 4132 564
rect 4156 556 4164 564
rect 3852 536 3860 544
rect 3996 536 4004 544
rect 3564 518 3572 524
rect 3564 516 3572 518
rect 3372 496 3380 504
rect 3436 496 3444 504
rect 3500 496 3508 504
rect 3484 476 3492 484
rect 3308 336 3316 344
rect 3228 316 3236 324
rect 3084 276 3092 284
rect 3004 236 3012 244
rect 3052 236 3060 244
rect 3148 276 3156 284
rect 3196 276 3204 284
rect 3020 196 3028 204
rect 3100 196 3108 204
rect 3004 156 3012 164
rect 2812 116 2820 124
rect 3340 316 3348 324
rect 3276 296 3284 304
rect 3292 296 3300 304
rect 3244 276 3252 284
rect 3164 256 3172 264
rect 3100 176 3108 184
rect 3244 196 3252 204
rect 3068 156 3076 164
rect 3084 156 3092 164
rect 3164 156 3172 164
rect 3228 156 3236 164
rect 3884 476 3892 484
rect 3948 476 3956 484
rect 3564 416 3572 424
rect 3500 376 3508 384
rect 3548 376 3556 384
rect 3532 316 3540 324
rect 3356 296 3364 304
rect 3596 316 3604 324
rect 4172 476 4180 484
rect 4028 436 4036 444
rect 4188 396 4196 404
rect 4172 336 4180 344
rect 4220 316 4228 324
rect 3676 296 3684 304
rect 3804 302 3812 304
rect 3804 296 3812 302
rect 4124 296 4132 304
rect 3436 276 3444 284
rect 3468 276 3476 284
rect 3612 276 3620 284
rect 3740 276 3748 284
rect 3612 256 3620 264
rect 3372 236 3380 244
rect 3420 236 3428 244
rect 3564 216 3572 224
rect 3452 196 3460 204
rect 3324 176 3332 184
rect 3372 176 3380 184
rect 3276 156 3284 164
rect 3756 156 3764 164
rect 3932 236 3940 244
rect 3260 136 3268 144
rect 3500 136 3508 144
rect 3692 136 3700 144
rect 3852 136 3860 144
rect 4140 276 4148 284
rect 4220 296 4228 304
rect 4076 256 4084 264
rect 4124 256 4132 264
rect 4108 216 4116 224
rect 4092 196 4100 204
rect 4028 156 4036 164
rect 4140 156 4148 164
rect 4156 156 4164 164
rect 4188 216 4196 224
rect 3052 116 3060 124
rect 3196 116 3204 124
rect 3372 116 3380 124
rect 2780 96 2788 104
rect 3020 96 3028 104
rect 2428 76 2436 84
rect 2524 76 2532 84
rect 2556 76 2564 84
rect 2716 76 2724 84
rect 4012 136 4020 144
rect 4124 136 4132 144
rect 4172 136 4180 144
rect 3820 118 3828 124
rect 3820 116 3828 118
rect 3948 116 3956 124
rect 4684 876 4692 884
rect 4604 736 4612 744
rect 4316 696 4324 704
rect 4380 696 4388 704
rect 4524 696 4532 704
rect 4588 696 4596 704
rect 4748 716 4756 724
rect 4844 856 4852 864
rect 4828 836 4836 844
rect 4796 756 4804 764
rect 4780 736 4788 744
rect 4780 716 4788 724
rect 4380 676 4388 684
rect 4556 676 4564 684
rect 4588 676 4596 684
rect 4780 676 4788 684
rect 4300 656 4308 664
rect 4364 636 4372 644
rect 4348 576 4356 584
rect 4412 636 4420 644
rect 4396 576 4404 584
rect 4332 556 4340 564
rect 4380 556 4388 564
rect 4348 536 4356 544
rect 4300 496 4308 504
rect 4252 356 4260 364
rect 4252 296 4260 304
rect 4268 296 4276 304
rect 4236 176 4244 184
rect 4220 136 4228 144
rect 4284 276 4292 284
rect 4268 196 4276 204
rect 4364 436 4372 444
rect 4316 376 4324 384
rect 4364 356 4372 364
rect 4540 656 4548 664
rect 4508 596 4516 604
rect 4492 536 4500 544
rect 4524 576 4532 584
rect 4556 576 4564 584
rect 4572 556 4580 564
rect 4620 656 4628 664
rect 4716 656 4724 664
rect 4892 1016 4900 1024
rect 5068 1496 5076 1504
rect 5116 1696 5124 1704
rect 5100 1676 5108 1684
rect 5132 1676 5140 1684
rect 5180 1716 5188 1724
rect 5196 1696 5204 1704
rect 5164 1676 5172 1684
rect 5148 1636 5156 1644
rect 5132 1596 5140 1604
rect 5196 1556 5204 1564
rect 5132 1516 5140 1524
rect 5164 1496 5172 1504
rect 5100 1396 5108 1404
rect 5164 1456 5172 1464
rect 5132 1336 5140 1344
rect 5116 1276 5124 1284
rect 5164 1276 5172 1284
rect 5084 1102 5092 1104
rect 5084 1096 5092 1102
rect 5132 1176 5140 1184
rect 5228 1756 5236 1764
rect 5244 1756 5252 1764
rect 5244 1616 5252 1624
rect 5324 1856 5332 1864
rect 5484 1916 5492 1924
rect 5388 1896 5396 1904
rect 5580 1896 5588 1904
rect 5356 1856 5364 1864
rect 5340 1816 5348 1824
rect 5324 1796 5332 1804
rect 5308 1776 5316 1784
rect 5292 1756 5300 1764
rect 5308 1736 5316 1744
rect 5308 1716 5316 1724
rect 5276 1696 5284 1704
rect 5292 1676 5300 1684
rect 5276 1656 5284 1664
rect 5308 1576 5316 1584
rect 5260 1556 5268 1564
rect 5340 1756 5348 1764
rect 5420 1876 5428 1884
rect 5404 1796 5412 1804
rect 5436 1756 5444 1764
rect 5388 1736 5396 1744
rect 5484 1876 5492 1884
rect 5436 1736 5444 1744
rect 5452 1736 5460 1744
rect 5372 1676 5380 1684
rect 5372 1656 5380 1664
rect 5388 1656 5396 1664
rect 5356 1636 5364 1644
rect 5372 1616 5380 1624
rect 5404 1616 5412 1624
rect 5340 1576 5348 1584
rect 5324 1536 5332 1544
rect 5228 1516 5236 1524
rect 5276 1516 5284 1524
rect 5308 1516 5316 1524
rect 5244 1496 5252 1504
rect 5292 1496 5300 1504
rect 5340 1496 5348 1504
rect 5260 1476 5268 1484
rect 5340 1476 5348 1484
rect 5324 1456 5332 1464
rect 5228 1416 5236 1424
rect 5212 1376 5220 1384
rect 5356 1456 5364 1464
rect 5324 1336 5332 1344
rect 5260 1296 5268 1304
rect 5388 1536 5396 1544
rect 5404 1496 5412 1504
rect 5404 1476 5412 1484
rect 5692 2076 5700 2084
rect 5852 2096 5860 2104
rect 5708 1902 5716 1904
rect 5708 1896 5716 1902
rect 5644 1876 5652 1884
rect 5596 1836 5604 1844
rect 5564 1776 5572 1784
rect 5468 1696 5476 1704
rect 5452 1656 5460 1664
rect 5436 1496 5444 1504
rect 5468 1636 5476 1644
rect 5500 1676 5508 1684
rect 5516 1636 5524 1644
rect 5532 1616 5540 1624
rect 5516 1596 5524 1604
rect 5436 1476 5444 1484
rect 5404 1456 5412 1464
rect 5420 1456 5428 1464
rect 5388 1336 5396 1344
rect 5436 1336 5444 1344
rect 5356 1296 5364 1304
rect 5372 1296 5380 1304
rect 5436 1296 5444 1304
rect 5388 1276 5396 1284
rect 5324 1236 5332 1244
rect 5404 1236 5412 1244
rect 5292 1116 5300 1124
rect 5276 1096 5284 1104
rect 5340 1136 5348 1144
rect 5452 1136 5460 1144
rect 5484 1496 5492 1504
rect 5516 1456 5524 1464
rect 5660 1816 5668 1824
rect 5836 1816 5844 1824
rect 5852 1696 5860 1704
rect 5708 1636 5716 1644
rect 5628 1476 5636 1484
rect 5708 1476 5716 1484
rect 5484 1416 5492 1424
rect 5532 1416 5540 1424
rect 5660 1396 5668 1404
rect 5564 1376 5572 1384
rect 5772 1356 5780 1364
rect 5500 1336 5508 1344
rect 5484 1236 5492 1244
rect 5676 1176 5684 1184
rect 5820 1176 5828 1184
rect 5628 1116 5636 1124
rect 5692 1116 5700 1124
rect 5516 1096 5524 1104
rect 5596 1096 5604 1104
rect 5436 1076 5444 1084
rect 5468 1076 5476 1084
rect 5500 1076 5508 1084
rect 5548 1076 5556 1084
rect 5660 1076 5668 1084
rect 5356 1036 5364 1044
rect 5404 1036 5412 1044
rect 5468 1036 5476 1044
rect 5292 1016 5300 1024
rect 5036 916 5044 924
rect 5180 916 5188 924
rect 4876 856 4884 864
rect 4972 876 4980 884
rect 5244 876 5252 884
rect 5292 876 5300 884
rect 5036 836 5044 844
rect 4940 736 4948 744
rect 5244 716 5252 724
rect 5324 716 5332 724
rect 5372 1016 5380 1024
rect 5420 936 5428 944
rect 4844 676 4852 684
rect 4764 656 4772 664
rect 4780 656 4788 664
rect 4844 656 4852 664
rect 4732 616 4740 624
rect 4604 576 4612 584
rect 4780 616 4788 624
rect 4796 576 4804 584
rect 4972 696 4980 704
rect 5068 696 5076 704
rect 5180 696 5188 704
rect 5772 1016 5780 1024
rect 5836 1016 5844 1024
rect 5548 936 5556 944
rect 5484 876 5492 884
rect 4924 676 4932 684
rect 4924 636 4932 644
rect 4700 556 4708 564
rect 4588 536 4596 544
rect 4636 536 4644 544
rect 4684 536 4692 544
rect 4716 536 4724 544
rect 4812 516 4820 524
rect 4572 496 4580 504
rect 4652 496 4660 504
rect 4684 496 4692 504
rect 4764 496 4772 504
rect 4524 476 4532 484
rect 4636 476 4644 484
rect 4476 456 4484 464
rect 4446 406 4454 414
rect 4460 406 4468 414
rect 4474 406 4482 414
rect 4588 376 4596 384
rect 4556 336 4564 344
rect 4604 356 4612 364
rect 4316 276 4324 284
rect 4332 276 4340 284
rect 4380 276 4388 284
rect 4396 276 4404 284
rect 4476 316 4484 324
rect 4492 316 4500 324
rect 4332 196 4340 204
rect 4348 196 4356 204
rect 4380 196 4388 204
rect 4412 196 4420 204
rect 4444 196 4452 204
rect 4332 156 4340 164
rect 4300 136 4308 144
rect 4524 216 4532 224
rect 4572 216 4580 224
rect 4556 196 4564 204
rect 4652 336 4660 344
rect 4892 576 4900 584
rect 4908 576 4916 584
rect 4860 556 4868 564
rect 4860 536 4868 544
rect 4988 676 4996 684
rect 5052 676 5060 684
rect 4972 656 4980 664
rect 4988 656 4996 664
rect 4956 576 4964 584
rect 4940 536 4948 544
rect 4876 516 4884 524
rect 4844 476 4852 484
rect 4700 436 4708 444
rect 4716 396 4724 404
rect 4764 376 4772 384
rect 4796 376 4804 384
rect 4684 296 4692 304
rect 4700 296 4708 304
rect 4620 276 4628 284
rect 4636 276 4644 284
rect 4668 236 4676 244
rect 4636 216 4644 224
rect 4572 156 4580 164
rect 4588 156 4596 164
rect 4460 136 4468 144
rect 4524 136 4532 144
rect 4764 256 4772 264
rect 4860 376 4868 384
rect 4876 376 4884 384
rect 4876 356 4884 364
rect 4892 356 4900 364
rect 4844 296 4852 304
rect 4780 236 4788 244
rect 4812 236 4820 244
rect 4812 216 4820 224
rect 4748 196 4756 204
rect 4668 156 4676 164
rect 4684 156 4692 164
rect 4828 196 4836 204
rect 4652 116 4660 124
rect 4124 96 4132 104
rect 4620 96 4628 104
rect 4684 96 4692 104
rect 4796 116 4804 124
rect 4764 96 4772 104
rect 4924 496 4932 504
rect 4940 396 4948 404
rect 4908 236 4916 244
rect 5004 636 5012 644
rect 5036 636 5044 644
rect 4972 536 4980 544
rect 5004 536 5012 544
rect 5036 496 5044 504
rect 5020 476 5028 484
rect 4988 376 4996 384
rect 5020 316 5028 324
rect 5100 676 5108 684
rect 5148 676 5156 684
rect 5196 676 5204 684
rect 5308 676 5316 684
rect 5404 676 5412 684
rect 5100 656 5108 664
rect 5148 656 5156 664
rect 5196 656 5204 664
rect 5292 656 5300 664
rect 5084 556 5092 564
rect 5116 556 5124 564
rect 5420 636 5428 644
rect 5228 576 5236 584
rect 5852 936 5860 944
rect 5580 876 5588 884
rect 5756 896 5764 904
rect 5596 716 5604 724
rect 5660 716 5668 724
rect 5852 696 5860 704
rect 5532 676 5540 684
rect 5516 576 5524 584
rect 5084 536 5092 544
rect 5116 516 5124 524
rect 5356 516 5364 524
rect 5500 516 5508 524
rect 5068 396 5076 404
rect 5100 476 5108 484
rect 5084 356 5092 364
rect 5084 316 5092 324
rect 4972 236 4980 244
rect 5052 256 5060 264
rect 5068 256 5076 264
rect 5100 276 5108 284
rect 5052 216 5060 224
rect 5004 196 5012 204
rect 5068 196 5076 204
rect 5164 496 5172 504
rect 5148 296 5156 304
rect 5148 236 5156 244
rect 5132 196 5140 204
rect 5196 396 5204 404
rect 5436 436 5444 444
rect 5292 336 5300 344
rect 5180 256 5188 264
rect 5196 216 5204 224
rect 4924 156 4932 164
rect 5068 156 5076 164
rect 5100 156 5108 164
rect 5116 156 5124 164
rect 4956 136 4964 144
rect 5020 136 5028 144
rect 5164 136 5172 144
rect 4860 116 4868 124
rect 5228 176 5236 184
rect 4940 116 4948 124
rect 4988 116 4996 124
rect 5100 116 5108 124
rect 5260 236 5268 244
rect 5404 316 5412 324
rect 5276 216 5284 224
rect 5436 296 5444 304
rect 5500 296 5508 304
rect 5500 276 5508 284
rect 5420 216 5428 224
rect 5388 196 5396 204
rect 5356 156 5364 164
rect 5276 136 5284 144
rect 5292 136 5300 144
rect 5340 136 5348 144
rect 5628 576 5636 584
rect 5596 536 5604 544
rect 5724 536 5732 544
rect 5564 518 5572 524
rect 5564 516 5572 518
rect 5692 516 5700 524
rect 5756 518 5764 524
rect 5756 516 5764 518
rect 5564 496 5572 504
rect 5580 436 5588 444
rect 5548 316 5556 324
rect 5548 276 5556 284
rect 5596 316 5604 324
rect 5628 296 5636 304
rect 5788 296 5796 304
rect 5644 276 5652 284
rect 5788 276 5796 284
rect 5484 216 5492 224
rect 5484 176 5492 184
rect 5612 256 5620 264
rect 5516 236 5524 244
rect 5596 196 5604 204
rect 5756 256 5764 264
rect 5772 236 5780 244
rect 5660 216 5668 224
rect 5772 216 5780 224
rect 5644 176 5652 184
rect 5724 176 5732 184
rect 5468 156 5476 164
rect 5436 136 5444 144
rect 5452 136 5460 144
rect 5708 156 5716 164
rect 5500 136 5508 144
rect 5356 116 5364 124
rect 5404 116 5412 124
rect 5468 116 5476 124
rect 5548 136 5556 144
rect 5644 116 5652 124
rect 5740 116 5748 124
rect 5820 176 5828 184
rect 5212 96 5220 104
rect 5532 96 5540 104
rect 5564 96 5572 104
rect 5612 96 5620 104
rect 5772 96 5780 104
rect 5804 96 5812 104
rect 5852 96 5860 104
rect 3628 76 3636 84
rect 4300 76 4308 84
rect 2012 56 2020 64
rect 2332 56 2340 64
rect 2396 56 2404 64
rect 3436 56 3444 64
rect 1358 6 1366 14
rect 1372 6 1380 14
rect 1386 6 1394 14
rect 4446 6 4454 14
rect 4460 6 4468 14
rect 4474 6 4482 14
<< metal3 >>
rect 2904 4214 2952 4216
rect 2904 4206 2908 4214
rect 2918 4206 2924 4214
rect 2932 4206 2938 4214
rect 2948 4206 2952 4214
rect 2904 4204 2952 4206
rect 980 4197 1948 4203
rect 4772 4197 4780 4203
rect 1949 4183 1955 4196
rect 1949 4177 3148 4183
rect 3156 4177 3884 4183
rect 3940 4177 4396 4183
rect 356 4157 396 4163
rect 1396 4157 1452 4163
rect 1508 4157 1740 4163
rect 2036 4157 2092 4163
rect 2180 4157 2204 4163
rect 2420 4157 2556 4163
rect 4196 4157 4796 4163
rect 5076 4157 5148 4163
rect 116 4137 172 4143
rect 180 4137 284 4143
rect 292 4137 444 4143
rect 628 4137 812 4143
rect 820 4137 844 4143
rect 852 4137 1100 4143
rect 1236 4137 1340 4143
rect 1444 4137 1484 4143
rect 1501 4137 1932 4143
rect 52 4117 92 4123
rect 100 4117 204 4123
rect 212 4117 316 4123
rect 324 4117 380 4123
rect 388 4117 428 4123
rect 1501 4123 1507 4137
rect 1988 4137 2124 4143
rect 2132 4137 2444 4143
rect 2676 4137 2716 4143
rect 2948 4137 3020 4143
rect 3028 4137 3228 4143
rect 3236 4137 3724 4143
rect 3876 4137 3900 4143
rect 4340 4137 4364 4143
rect 4948 4137 4972 4143
rect 5268 4137 5436 4143
rect 5700 4137 5804 4143
rect 596 4117 1507 4123
rect 1684 4117 1772 4123
rect 1812 4117 1868 4123
rect 1956 4117 2012 4123
rect 2084 4117 2108 4123
rect 2340 4117 2396 4123
rect 2660 4117 2732 4123
rect 3300 4117 3388 4123
rect 3460 4117 3548 4123
rect 3860 4117 3932 4123
rect 4324 4117 4412 4123
rect 4932 4117 5020 4123
rect 5476 4117 5580 4123
rect 20 4097 348 4103
rect 788 4097 1260 4103
rect 1428 4097 1644 4103
rect 1652 4097 1788 4103
rect 1828 4097 1996 4103
rect 2004 4097 2188 4103
rect 2292 4097 2492 4103
rect 2500 4097 3196 4103
rect 3764 4097 3900 4103
rect 3908 4097 3980 4103
rect 4228 4097 4364 4103
rect 4372 4097 4492 4103
rect 4836 4097 4972 4103
rect 4980 4097 5052 4103
rect 436 4077 572 4083
rect 580 4077 652 4083
rect 1172 4077 1532 4083
rect 1732 4077 1916 4083
rect 1924 4077 3004 4083
rect 4020 4077 4508 4083
rect 388 4057 620 4063
rect 996 4057 2780 4063
rect 276 4037 380 4043
rect 1604 4037 1660 4043
rect 1668 4037 1932 4043
rect 1940 4037 2268 4043
rect 2436 4037 2668 4043
rect 3572 4037 4108 4043
rect 1876 4017 2012 4023
rect 2100 4017 2540 4023
rect 2564 4017 3676 4023
rect 5380 4017 5516 4023
rect 5636 4017 5660 4023
rect 1352 4014 1400 4016
rect 1352 4006 1356 4014
rect 1366 4006 1372 4014
rect 1380 4006 1386 4014
rect 1396 4006 1400 4014
rect 1352 4004 1400 4006
rect 4440 4014 4488 4016
rect 4440 4006 4444 4014
rect 4454 4006 4460 4014
rect 4468 4006 4474 4014
rect 4484 4006 4488 4014
rect 4440 4004 4488 4006
rect 1764 3997 2332 4003
rect 2340 3997 3052 4003
rect 4036 3997 4380 4003
rect 4580 3997 4732 4003
rect 228 3977 492 3983
rect 1332 3977 1612 3983
rect 1620 3977 1804 3983
rect 1892 3977 1996 3983
rect 2020 3977 2156 3983
rect 2740 3977 2780 3983
rect 2788 3977 3164 3983
rect 3172 3977 3244 3983
rect 3252 3977 3308 3983
rect 84 3957 428 3963
rect 436 3957 540 3963
rect 1460 3957 1836 3963
rect 1844 3957 1852 3963
rect 1860 3957 2348 3963
rect 36 3937 332 3943
rect 388 3937 764 3943
rect 772 3937 1004 3943
rect 1492 3937 1596 3943
rect 1604 3937 1708 3943
rect 1716 3937 1756 3943
rect 1764 3937 2140 3943
rect 2212 3937 2428 3943
rect 2436 3937 2476 3943
rect 228 3917 252 3923
rect 420 3917 444 3923
rect 804 3917 860 3923
rect 900 3917 972 3923
rect 980 3917 1084 3923
rect 1092 3917 1148 3923
rect 1588 3917 1708 3923
rect 1716 3917 1772 3923
rect 1780 3917 1948 3923
rect 1956 3917 2044 3923
rect 2276 3917 2428 3923
rect 2548 3917 2716 3923
rect 2772 3917 2796 3923
rect 3092 3917 3116 3923
rect 3140 3917 3260 3923
rect 4644 3917 4764 3923
rect 4772 3917 4780 3923
rect 4788 3917 4860 3923
rect 164 3897 476 3903
rect 484 3897 524 3903
rect 628 3897 924 3903
rect 932 3897 1052 3903
rect 1268 3897 1404 3903
rect 1636 3897 1660 3903
rect 1684 3897 1724 3903
rect 1892 3897 1964 3903
rect 1988 3897 2284 3903
rect 2708 3897 2812 3903
rect 3133 3903 3139 3916
rect 2932 3897 3139 3903
rect 3220 3897 3276 3903
rect 3492 3897 3532 3903
rect 3540 3897 3612 3903
rect 3780 3897 3964 3903
rect 4036 3897 4140 3903
rect 4148 3897 4236 3903
rect 4244 3897 4284 3903
rect 4740 3897 4812 3903
rect 4996 3897 5052 3903
rect 20 3877 76 3883
rect 116 3877 220 3883
rect 548 3877 636 3883
rect 756 3877 828 3883
rect 932 3877 988 3883
rect 996 3877 1004 3883
rect 1044 3877 1084 3883
rect 1092 3877 1116 3883
rect 1124 3877 1244 3883
rect 1620 3877 1660 3883
rect 1796 3877 1900 3883
rect 2036 3877 2124 3883
rect 2212 3877 2236 3883
rect 2292 3877 2380 3883
rect 2660 3877 2748 3883
rect 2996 3877 3036 3883
rect 3428 3877 3484 3883
rect 3556 3877 3580 3883
rect 3588 3877 3692 3883
rect 3700 3877 3740 3883
rect 4116 3877 4188 3883
rect 4756 3877 4780 3883
rect 5460 3877 5596 3883
rect 308 3857 332 3863
rect 372 3857 412 3863
rect 1380 3857 1628 3863
rect 1700 3857 1868 3863
rect 1908 3857 1916 3863
rect 1972 3857 2540 3863
rect 2564 3857 2716 3863
rect 3028 3857 3228 3863
rect 4756 3857 4796 3863
rect 4884 3857 4956 3863
rect 164 3837 1132 3843
rect 1492 3837 2460 3843
rect 2500 3837 2860 3843
rect 5028 3837 5148 3843
rect 1284 3817 1955 3823
rect 644 3797 1516 3803
rect 1949 3803 1955 3817
rect 2148 3817 2460 3823
rect 2548 3817 2876 3823
rect 4340 3817 4396 3823
rect 4404 3817 4812 3823
rect 4820 3817 4924 3823
rect 4932 3817 5004 3823
rect 5012 3817 5324 3823
rect 5332 3817 5340 3823
rect 2904 3814 2952 3816
rect 2904 3806 2908 3814
rect 2918 3806 2924 3814
rect 2932 3806 2938 3814
rect 2948 3806 2952 3814
rect 2904 3804 2952 3806
rect 1949 3797 2588 3803
rect 2628 3797 2668 3803
rect 3060 3797 3116 3803
rect 3124 3797 3228 3803
rect 4404 3797 4444 3803
rect 5108 3797 5116 3803
rect 5252 3797 5308 3803
rect 356 3777 892 3783
rect 1540 3777 2332 3783
rect 2532 3777 2700 3783
rect 2708 3777 2764 3783
rect 2884 3777 3116 3783
rect 3732 3777 3932 3783
rect 3940 3777 4204 3783
rect 4212 3777 4284 3783
rect 4292 3777 4604 3783
rect 324 3757 364 3763
rect 372 3757 732 3763
rect 1764 3757 1788 3763
rect 1812 3757 1916 3763
rect 1956 3757 2028 3763
rect 2052 3757 2076 3763
rect 2116 3757 2300 3763
rect 2404 3757 2556 3763
rect 2756 3757 2876 3763
rect 2893 3757 3180 3763
rect 2893 3744 2899 3757
rect 3524 3757 3628 3763
rect 3636 3757 3676 3763
rect 3748 3757 3820 3763
rect 3828 3757 3900 3763
rect 4516 3757 4556 3763
rect 4564 3757 4876 3763
rect 4980 3757 5020 3763
rect 36 3737 60 3743
rect 116 3737 124 3743
rect 132 3737 172 3743
rect 324 3737 476 3743
rect 660 3737 844 3743
rect 1300 3737 1500 3743
rect 1972 3737 1996 3743
rect 2132 3737 2252 3743
rect 2276 3737 2284 3743
rect 2308 3737 2508 3743
rect 2516 3737 2796 3743
rect 2804 3737 2892 3743
rect 3028 3737 3052 3743
rect 3444 3737 3612 3743
rect 3636 3737 3644 3743
rect 3652 3737 3852 3743
rect 4324 3737 4380 3743
rect 4388 3737 4540 3743
rect 4788 3737 4892 3743
rect 4900 3737 4956 3743
rect 5620 3737 5788 3743
rect 68 3717 236 3723
rect 244 3717 316 3723
rect 628 3717 636 3723
rect 724 3717 764 3723
rect 916 3717 940 3723
rect 1476 3717 1836 3723
rect 1844 3717 1996 3723
rect 2004 3717 2076 3723
rect 2084 3717 2092 3723
rect 2100 3717 2108 3723
rect 2180 3717 2188 3723
rect 2196 3717 2444 3723
rect 2452 3717 2572 3723
rect 2628 3717 2668 3723
rect 2676 3717 2764 3723
rect 3508 3717 3772 3723
rect 4004 3717 4060 3723
rect 4068 3717 4188 3723
rect 4356 3717 4380 3723
rect 4420 3717 4460 3723
rect 4884 3717 4924 3723
rect 5124 3717 5148 3723
rect 5156 3717 5276 3723
rect 212 3697 284 3703
rect 356 3697 364 3703
rect 372 3697 460 3703
rect 468 3697 684 3703
rect 1108 3697 1628 3703
rect 1876 3697 2044 3703
rect 2052 3697 2220 3703
rect 2228 3697 2396 3703
rect 2564 3697 2780 3703
rect 2868 3697 3020 3703
rect 3252 3697 3532 3703
rect 3764 3697 3804 3703
rect 148 3677 428 3683
rect 740 3677 972 3683
rect 1732 3677 1900 3683
rect 1940 3677 2076 3683
rect 2164 3677 2252 3683
rect 2260 3677 2412 3683
rect 2420 3677 2508 3683
rect 2564 3677 2636 3683
rect 3556 3677 3660 3683
rect 3668 3677 3804 3683
rect 68 3657 220 3663
rect 388 3657 748 3663
rect 772 3657 1164 3663
rect 1924 3657 2236 3663
rect 196 3637 220 3643
rect 228 3637 300 3643
rect 308 3637 492 3643
rect 788 3637 988 3643
rect 1316 3637 1404 3643
rect 1780 3637 2012 3643
rect 4996 3637 5180 3643
rect 5188 3637 5356 3643
rect 5364 3637 5420 3643
rect 100 3617 204 3623
rect 212 3617 268 3623
rect 356 3617 396 3623
rect 484 3617 540 3623
rect 2452 3617 3340 3623
rect 1352 3614 1400 3616
rect 1352 3606 1356 3614
rect 1366 3606 1372 3614
rect 1380 3606 1386 3614
rect 1396 3606 1400 3614
rect 1352 3604 1400 3606
rect 4440 3614 4488 3616
rect 4440 3606 4444 3614
rect 4454 3606 4460 3614
rect 4468 3606 4474 3614
rect 4484 3606 4488 3614
rect 4440 3604 4488 3606
rect 260 3597 572 3603
rect 580 3597 604 3603
rect 1604 3597 1948 3603
rect 1965 3597 2876 3603
rect 1965 3583 1971 3597
rect 1668 3577 1971 3583
rect 2244 3577 2444 3583
rect 2500 3577 2620 3583
rect 2628 3577 2892 3583
rect 3700 3577 3788 3583
rect 4740 3577 4812 3583
rect 1860 3557 2684 3563
rect 2708 3557 3260 3563
rect 3892 3557 4924 3563
rect 4932 3557 5004 3563
rect 164 3537 188 3543
rect 436 3537 636 3543
rect 1508 3537 1596 3543
rect 1604 3537 1788 3543
rect 1796 3537 1980 3543
rect 2020 3537 2156 3543
rect 2173 3537 2579 3543
rect 292 3517 492 3523
rect 612 3517 652 3523
rect 884 3517 1132 3523
rect 1140 3517 1180 3523
rect 1316 3517 1356 3523
rect 1380 3517 1996 3523
rect 2173 3523 2179 3537
rect 2084 3517 2179 3523
rect 2484 3517 2556 3523
rect 2573 3523 2579 3537
rect 2676 3537 2764 3543
rect 2772 3537 2924 3543
rect 4116 3537 4252 3543
rect 4260 3537 4316 3543
rect 4756 3537 4844 3543
rect 2573 3517 2684 3523
rect 2701 3517 2780 3523
rect 52 3497 60 3503
rect 180 3497 412 3503
rect 420 3497 620 3503
rect 692 3497 748 3503
rect 1172 3497 1212 3503
rect 1220 3497 1324 3503
rect 1972 3497 2092 3503
rect 2148 3497 2284 3503
rect 2324 3497 2364 3503
rect 2372 3497 2492 3503
rect 2701 3503 2707 3517
rect 2948 3517 3036 3523
rect 4132 3517 4172 3523
rect 4276 3517 4412 3523
rect 4516 3517 4636 3523
rect 4644 3517 4684 3523
rect 2660 3497 2707 3503
rect 2756 3497 2940 3503
rect 2996 3497 3148 3503
rect 3460 3497 3516 3503
rect 3652 3497 3740 3503
rect 4068 3497 4124 3503
rect 4164 3497 4300 3503
rect 4356 3497 4524 3503
rect 4532 3497 4572 3503
rect 5156 3497 5180 3503
rect 196 3477 332 3483
rect 340 3477 460 3483
rect 468 3477 476 3483
rect 516 3477 556 3483
rect 628 3477 780 3483
rect 788 3477 796 3483
rect 900 3477 1020 3483
rect 1028 3477 1196 3483
rect 1204 3477 1420 3483
rect 1428 3477 1724 3483
rect 1732 3477 1836 3483
rect 1972 3477 2092 3483
rect 2228 3477 2380 3483
rect 2388 3477 3027 3483
rect 3021 3464 3027 3477
rect 3220 3477 3260 3483
rect 3492 3477 3708 3483
rect 3716 3477 4028 3483
rect 4180 3477 4268 3483
rect 4388 3477 4492 3483
rect 4500 3477 4540 3483
rect 4596 3477 4684 3483
rect 5220 3477 5276 3483
rect 5476 3477 5628 3483
rect 68 3457 76 3463
rect 84 3457 220 3463
rect 340 3457 380 3463
rect 452 3457 476 3463
rect 612 3457 764 3463
rect 772 3457 828 3463
rect 1076 3457 1372 3463
rect 2196 3457 2316 3463
rect 2452 3457 2476 3463
rect 2564 3457 2748 3463
rect 2852 3457 2956 3463
rect 3028 3457 3100 3463
rect 3108 3457 3308 3463
rect 4244 3457 4508 3463
rect 5124 3457 5308 3463
rect 372 3437 428 3443
rect 436 3437 524 3443
rect 692 3437 1228 3443
rect 1492 3437 1548 3443
rect 1956 3437 2252 3443
rect 2500 3437 2988 3443
rect 2996 3437 3276 3443
rect 3284 3437 3548 3443
rect 4436 3437 4556 3443
rect 5796 3437 5820 3443
rect 196 3417 796 3423
rect 1172 3417 1196 3423
rect 1204 3417 1516 3423
rect 2628 3417 2716 3423
rect 3124 3417 3180 3423
rect 2904 3414 2952 3416
rect 2904 3406 2908 3414
rect 2918 3406 2924 3414
rect 2932 3406 2938 3414
rect 2948 3406 2952 3414
rect 2904 3404 2952 3406
rect 388 3397 540 3403
rect 548 3397 588 3403
rect 596 3397 748 3403
rect 1540 3397 1740 3403
rect 2628 3397 2668 3403
rect 3092 3397 3116 3403
rect 3140 3397 3324 3403
rect 3332 3397 3564 3403
rect 3764 3397 3916 3403
rect 3940 3397 3964 3403
rect 4196 3397 4492 3403
rect 4500 3397 4508 3403
rect 4516 3397 4700 3403
rect 5316 3397 5372 3403
rect 5380 3397 5660 3403
rect 788 3377 812 3383
rect 1028 3377 1084 3383
rect 1140 3377 1244 3383
rect 1412 3377 1628 3383
rect 1636 3377 1724 3383
rect 2068 3377 2188 3383
rect 2196 3377 2332 3383
rect 2420 3377 2508 3383
rect 2548 3377 2700 3383
rect 2836 3377 3148 3383
rect 4084 3377 4732 3383
rect 5124 3377 5132 3383
rect 116 3357 252 3363
rect 276 3357 316 3363
rect 724 3357 812 3363
rect 820 3357 892 3363
rect 964 3357 1020 3363
rect 1044 3357 1180 3363
rect 1245 3357 1596 3363
rect 324 3337 412 3343
rect 900 3337 972 3343
rect 1245 3343 1251 3357
rect 1604 3357 1644 3363
rect 2404 3357 2428 3363
rect 2436 3357 2460 3363
rect 2468 3357 2540 3363
rect 2644 3357 2684 3363
rect 2740 3357 2812 3363
rect 2852 3357 3020 3363
rect 3076 3357 3107 3363
rect 1076 3337 1251 3343
rect 1268 3337 1308 3343
rect 1348 3337 1436 3343
rect 1572 3337 1596 3343
rect 2452 3337 2652 3343
rect 2660 3337 2732 3343
rect 2772 3337 3004 3343
rect 3012 3337 3068 3343
rect 3101 3343 3107 3357
rect 3124 3357 3196 3363
rect 3876 3357 3900 3363
rect 4541 3357 4636 3363
rect 4541 3344 4547 3357
rect 5412 3357 5500 3363
rect 3101 3337 3228 3343
rect 3828 3337 3868 3343
rect 4116 3337 4236 3343
rect 4308 3337 4332 3343
rect 4388 3337 4476 3343
rect 4484 3337 4540 3343
rect 5380 3337 5532 3343
rect 5860 3337 5891 3343
rect 148 3317 252 3323
rect 260 3317 300 3323
rect 580 3317 700 3323
rect 852 3317 892 3323
rect 900 3317 940 3323
rect 964 3317 1020 3323
rect 1108 3317 1132 3323
rect 1316 3317 1372 3323
rect 1565 3323 1571 3336
rect 1396 3317 1571 3323
rect 1956 3317 1980 3323
rect 2132 3317 2188 3323
rect 2356 3317 2508 3323
rect 2532 3317 2636 3323
rect 2756 3317 2956 3323
rect 3476 3317 3532 3323
rect 3556 3317 3692 3323
rect 3700 3317 3836 3323
rect 4276 3317 4364 3323
rect 4564 3317 4604 3323
rect 5076 3317 5116 3323
rect 292 3297 364 3303
rect 548 3297 604 3303
rect 724 3297 748 3303
rect 1140 3297 1196 3303
rect 2404 3297 2556 3303
rect 2676 3297 2764 3303
rect 2804 3297 3100 3303
rect 3796 3297 3836 3303
rect 4692 3297 4748 3303
rect 5780 3297 5891 3303
rect 484 3277 524 3283
rect 660 3277 700 3283
rect 2292 3277 3020 3283
rect 3524 3277 3772 3283
rect 420 3257 668 3263
rect 676 3257 812 3263
rect 2564 3257 2764 3263
rect 4276 3257 4572 3263
rect 4580 3257 4764 3263
rect 84 3237 268 3243
rect 1732 3237 1996 3243
rect 3812 3237 3884 3243
rect 3892 3237 3916 3243
rect 5540 3237 5548 3243
rect 3828 3217 3900 3223
rect 3908 3217 3948 3223
rect 1352 3214 1400 3216
rect 1352 3206 1356 3214
rect 1366 3206 1372 3214
rect 1380 3206 1386 3214
rect 1396 3206 1400 3214
rect 1352 3204 1400 3206
rect 4440 3214 4488 3216
rect 4440 3206 4444 3214
rect 4454 3206 4460 3214
rect 4468 3206 4474 3214
rect 4484 3206 4488 3214
rect 4440 3204 4488 3206
rect 756 3197 796 3203
rect 804 3197 1228 3203
rect 1236 3197 1308 3203
rect 2132 3197 3260 3203
rect 484 3177 524 3183
rect 2340 3177 2348 3183
rect 2356 3177 2684 3183
rect 2692 3177 2732 3183
rect 3652 3177 3852 3183
rect 4180 3177 4684 3183
rect 4980 3177 5004 3183
rect 692 3157 908 3163
rect 2292 3157 2604 3163
rect 3380 3157 3420 3163
rect 3428 3157 3772 3163
rect 4132 3157 4284 3163
rect 20 3137 188 3143
rect 212 3137 316 3143
rect 420 3137 444 3143
rect 548 3137 636 3143
rect 676 3137 732 3143
rect 1204 3137 1372 3143
rect 2420 3137 2444 3143
rect 2500 3137 2636 3143
rect 2644 3137 2892 3143
rect 3108 3137 3532 3143
rect 3556 3137 4044 3143
rect 4452 3137 4588 3143
rect 4596 3137 4604 3143
rect 228 3117 252 3123
rect 308 3117 716 3123
rect 724 3117 924 3123
rect 1252 3117 1276 3123
rect 1444 3117 1516 3123
rect 1540 3117 1676 3123
rect 1940 3117 2316 3123
rect 2452 3117 2476 3123
rect 2724 3117 3164 3123
rect 3236 3117 3308 3123
rect 3396 3117 3436 3123
rect 3460 3117 3756 3123
rect 4260 3117 4348 3123
rect 4388 3117 4540 3123
rect 5300 3117 5356 3123
rect 5636 3117 5692 3123
rect 212 3097 364 3103
rect 500 3097 803 3103
rect 797 3084 803 3097
rect 900 3097 956 3103
rect 1076 3097 1324 3103
rect 1348 3097 1500 3103
rect 1508 3097 1692 3103
rect 1700 3097 1756 3103
rect 1764 3097 1996 3103
rect 2324 3097 2428 3103
rect 2468 3097 2508 3103
rect 2868 3097 3276 3103
rect 3284 3097 3356 3103
rect 3492 3097 3804 3103
rect 3860 3097 3884 3103
rect 3892 3097 3964 3103
rect 4308 3097 4396 3103
rect 4580 3097 4748 3103
rect 4820 3097 4844 3103
rect 5300 3097 5372 3103
rect 5421 3097 5891 3103
rect 5421 3084 5427 3097
rect 52 3077 108 3083
rect 116 3077 172 3083
rect 180 3077 300 3083
rect 340 3077 412 3083
rect 420 3077 508 3083
rect 612 3077 764 3083
rect 852 3077 972 3083
rect 980 3077 1036 3083
rect 1316 3077 1452 3083
rect 1540 3077 1564 3083
rect 1588 3077 1612 3083
rect 2308 3077 2396 3083
rect 2404 3077 2524 3083
rect 2932 3077 3036 3083
rect 3316 3077 3388 3083
rect 3668 3077 3843 3083
rect 132 3057 156 3063
rect 164 3057 204 3063
rect 244 3057 284 3063
rect 356 3057 396 3063
rect 836 3057 844 3063
rect 852 3057 876 3063
rect 932 3057 1004 3063
rect 1012 3057 1020 3063
rect 1028 3057 1052 3063
rect 1060 3057 1468 3063
rect 1476 3057 1724 3063
rect 3332 3057 3436 3063
rect 3764 3057 3820 3063
rect 3837 3063 3843 3077
rect 3940 3077 3964 3083
rect 3972 3077 4012 3083
rect 4020 3077 4140 3083
rect 4244 3077 4508 3083
rect 4516 3077 4524 3083
rect 4532 3077 4604 3083
rect 4884 3077 5164 3083
rect 5204 3077 5340 3083
rect 5348 3077 5420 3083
rect 5524 3077 5660 3083
rect 3837 3057 3884 3063
rect 4420 3057 4620 3063
rect 4788 3057 5004 3063
rect 5348 3057 5372 3063
rect 5444 3057 5468 3063
rect 5476 3057 5788 3063
rect 660 3037 716 3043
rect 1028 3037 1180 3043
rect 1188 3037 1212 3043
rect 1284 3037 1836 3043
rect 3924 3037 3980 3043
rect 4564 3037 4812 3043
rect 5332 3037 5500 3043
rect 340 3017 444 3023
rect 692 3017 908 3023
rect 1300 3017 1452 3023
rect 1508 3017 1548 3023
rect 1572 3017 1596 3023
rect 3780 3017 4140 3023
rect 2904 3014 2952 3016
rect 2904 3006 2908 3014
rect 2918 3006 2924 3014
rect 2932 3006 2938 3014
rect 2948 3006 2952 3014
rect 2904 3004 2952 3006
rect 228 2997 460 3003
rect 484 2997 828 3003
rect 1092 2997 1148 3003
rect 1188 2997 1564 3003
rect 3444 2997 3676 3003
rect 324 2977 364 2983
rect 372 2977 412 2983
rect 484 2977 508 2983
rect 516 2977 636 2983
rect 644 2977 668 2983
rect 676 2977 732 2983
rect 772 2977 780 2983
rect 996 2977 1020 2983
rect 1108 2977 1132 2983
rect 1140 2977 1372 2983
rect 1508 2977 1676 2983
rect 1700 2977 1756 2983
rect 1764 2977 1788 2983
rect 1796 2977 1820 2983
rect 2461 2977 2540 2983
rect 2461 2964 2467 2977
rect 3876 2977 3948 2983
rect 68 2957 124 2963
rect 148 2957 204 2963
rect 356 2957 380 2963
rect 388 2957 396 2963
rect 404 2957 508 2963
rect 516 2957 540 2963
rect 628 2957 748 2963
rect 772 2957 1180 2963
rect 1204 2957 1308 2963
rect 1332 2957 1516 2963
rect 1556 2957 1596 2963
rect 1716 2957 1788 2963
rect 5380 2957 5692 2963
rect 5748 2957 5788 2963
rect 196 2937 252 2943
rect 260 2937 364 2943
rect 372 2937 684 2943
rect 868 2937 892 2943
rect 900 2937 1020 2943
rect 1028 2937 1052 2943
rect 1140 2937 1196 2943
rect 1220 2937 1228 2943
rect 1252 2937 1468 2943
rect 1476 2937 1852 2943
rect 2708 2937 3228 2943
rect 3620 2937 3692 2943
rect 3876 2937 4028 2943
rect 4436 2937 4572 2943
rect 4596 2937 4620 2943
rect 4932 2937 4956 2943
rect 5092 2937 5116 2943
rect 5556 2937 5724 2943
rect 5732 2937 5788 2943
rect 5796 2937 5891 2943
rect 180 2917 236 2923
rect 308 2917 556 2923
rect 580 2917 620 2923
rect 660 2917 764 2923
rect 788 2917 876 2923
rect 884 2917 892 2923
rect 900 2917 908 2923
rect 964 2917 1804 2923
rect 1876 2917 2044 2923
rect 2116 2917 2460 2923
rect 2644 2917 2828 2923
rect 2900 2917 3036 2923
rect 3412 2917 3548 2923
rect 3556 2917 3740 2923
rect 4020 2917 4076 2923
rect 4548 2917 4604 2923
rect 4628 2917 4700 2923
rect 4916 2917 4940 2923
rect 5652 2917 5740 2923
rect 36 2897 76 2903
rect 340 2897 524 2903
rect 756 2897 908 2903
rect 1156 2897 1324 2903
rect 1444 2897 1484 2903
rect 1540 2897 1564 2903
rect 1588 2897 1612 2903
rect 2836 2897 2972 2903
rect 3028 2897 3164 2903
rect 3844 2897 3964 2903
rect 3972 2897 4044 2903
rect 4532 2897 4636 2903
rect 5652 2897 5692 2903
rect 5860 2897 5891 2903
rect 308 2877 492 2883
rect 772 2877 812 2883
rect 836 2877 1107 2883
rect 84 2857 108 2863
rect 132 2857 604 2863
rect 708 2857 1084 2863
rect 1101 2863 1107 2877
rect 1172 2877 1324 2883
rect 1476 2877 1532 2883
rect 1636 2877 1852 2883
rect 1860 2877 1900 2883
rect 3428 2877 3900 2883
rect 4580 2877 4604 2883
rect 4836 2877 5148 2883
rect 5284 2877 5804 2883
rect 1101 2857 1212 2863
rect 1300 2857 1980 2863
rect 3812 2857 4364 2863
rect 116 2837 156 2843
rect 932 2837 1116 2843
rect 1172 2837 1228 2843
rect 1316 2837 1356 2843
rect 1364 2837 1564 2843
rect 1572 2837 1740 2843
rect 2292 2837 2572 2843
rect 2612 2837 2764 2843
rect 3188 2837 3292 2843
rect 1352 2814 1400 2816
rect 1352 2806 1356 2814
rect 1366 2806 1372 2814
rect 1380 2806 1386 2814
rect 1396 2806 1400 2814
rect 1352 2804 1400 2806
rect 4440 2814 4488 2816
rect 4440 2806 4444 2814
rect 4454 2806 4460 2814
rect 4468 2806 4474 2814
rect 4484 2806 4488 2814
rect 4440 2804 4488 2806
rect 356 2797 700 2803
rect 996 2797 1084 2803
rect 196 2777 796 2783
rect 1268 2777 1436 2783
rect 3876 2777 3980 2783
rect 5620 2777 5628 2783
rect 484 2757 556 2763
rect 564 2757 588 2763
rect 596 2757 956 2763
rect 1284 2757 1452 2763
rect 228 2737 284 2743
rect 436 2737 524 2743
rect 532 2737 1244 2743
rect 1316 2737 1372 2743
rect 1492 2737 1692 2743
rect 1924 2737 2204 2743
rect 2628 2737 2684 2743
rect 3060 2737 3132 2743
rect 3140 2737 3484 2743
rect 3828 2737 4028 2743
rect 4228 2737 4332 2743
rect 4340 2737 4796 2743
rect 4804 2737 4844 2743
rect 148 2717 156 2723
rect 244 2717 268 2723
rect 324 2717 364 2723
rect 692 2717 1180 2723
rect 1188 2717 1212 2723
rect 1508 2717 1564 2723
rect 1572 2717 1635 2723
rect 1629 2704 1635 2717
rect 1668 2717 1724 2723
rect 1732 2717 1788 2723
rect 2180 2717 2412 2723
rect 2500 2717 2588 2723
rect 2596 2717 3116 2723
rect 3556 2717 3644 2723
rect 3860 2717 3884 2723
rect 3892 2717 3948 2723
rect 3988 2717 4044 2723
rect 4836 2717 4892 2723
rect 4964 2717 4988 2723
rect 5220 2717 5276 2723
rect 5604 2717 5660 2723
rect 180 2697 204 2703
rect 276 2697 348 2703
rect 612 2697 652 2703
rect 772 2697 972 2703
rect 1076 2697 1212 2703
rect 1252 2697 1468 2703
rect 1588 2697 1612 2703
rect 1636 2697 1692 2703
rect 2116 2697 2332 2703
rect 2388 2697 2428 2703
rect 2436 2697 2508 2703
rect 2580 2697 2652 2703
rect 2660 2697 2956 2703
rect 3012 2697 3036 2703
rect 3172 2697 3212 2703
rect 3220 2697 3276 2703
rect 3284 2697 3340 2703
rect 3620 2697 3708 2703
rect 3780 2697 3868 2703
rect 3876 2697 3900 2703
rect 4404 2697 4604 2703
rect 4964 2697 5116 2703
rect 5220 2697 5468 2703
rect 5860 2697 5891 2703
rect 180 2677 332 2683
rect 372 2677 412 2683
rect 548 2677 684 2683
rect 772 2677 844 2683
rect 996 2677 1020 2683
rect 1108 2677 1196 2683
rect 1204 2677 1228 2683
rect 1268 2677 1292 2683
rect 1316 2677 1516 2683
rect 1540 2677 1772 2683
rect 2308 2677 2396 2683
rect 2404 2677 2460 2683
rect 2516 2677 2556 2683
rect 2564 2677 2812 2683
rect 2948 2677 3084 2683
rect 3053 2664 3059 2677
rect 3124 2677 3180 2683
rect 3300 2677 3340 2683
rect 3348 2677 3388 2683
rect 3396 2677 3420 2683
rect 3588 2677 3740 2683
rect 3780 2677 3820 2683
rect 4308 2677 4668 2683
rect 5348 2677 5436 2683
rect 5444 2677 5628 2683
rect 292 2657 412 2663
rect 484 2657 556 2663
rect 836 2657 1004 2663
rect 1172 2657 1324 2663
rect 1332 2657 1548 2663
rect 1556 2657 1596 2663
rect 1604 2657 1644 2663
rect 2356 2657 2444 2663
rect 2452 2657 2620 2663
rect 2804 2657 2828 2663
rect 2852 2657 3036 2663
rect 3076 2657 3212 2663
rect 3348 2657 3404 2663
rect 3412 2657 3452 2663
rect 3812 2657 3891 2663
rect 3885 2644 3891 2657
rect 4036 2657 4124 2663
rect 68 2637 332 2643
rect 468 2637 492 2643
rect 500 2637 620 2643
rect 1348 2637 1372 2643
rect 1380 2637 1756 2643
rect 1828 2637 1980 2643
rect 2164 2637 2876 2643
rect 3108 2637 3324 2643
rect 3716 2637 3836 2643
rect 3892 2637 3932 2643
rect 3940 2637 3964 2643
rect 4452 2637 4572 2643
rect 5412 2637 5772 2643
rect 68 2617 188 2623
rect 196 2617 924 2623
rect 3252 2617 3292 2623
rect 3300 2617 3580 2623
rect 4388 2617 4876 2623
rect 5028 2617 5564 2623
rect 2904 2614 2952 2616
rect 2904 2606 2908 2614
rect 2918 2606 2924 2614
rect 2932 2606 2938 2614
rect 2948 2606 2952 2614
rect 2904 2604 2952 2606
rect 148 2597 540 2603
rect 1028 2597 1100 2603
rect 1108 2597 1180 2603
rect 1684 2597 1708 2603
rect 1908 2597 1980 2603
rect 1988 2597 2604 2603
rect 3732 2597 3932 2603
rect 3940 2597 3980 2603
rect 4356 2597 4396 2603
rect 4404 2597 4524 2603
rect 4596 2597 4636 2603
rect 4644 2597 4812 2603
rect 4820 2597 4940 2603
rect 116 2577 204 2583
rect 788 2577 908 2583
rect 916 2577 1180 2583
rect 1700 2577 2188 2583
rect 2420 2577 2620 2583
rect 3204 2577 3276 2583
rect 3284 2577 3308 2583
rect 3316 2577 3404 2583
rect 3668 2577 3996 2583
rect 4068 2577 4188 2583
rect 4324 2577 5292 2583
rect 196 2557 220 2563
rect 228 2557 268 2563
rect 340 2557 508 2563
rect 900 2557 940 2563
rect 1156 2557 1228 2563
rect 1812 2557 1868 2563
rect 1940 2557 1996 2563
rect 2308 2557 2732 2563
rect 3204 2557 3260 2563
rect 3508 2557 3532 2563
rect 3956 2557 4108 2563
rect 4996 2557 5020 2563
rect 20 2537 220 2543
rect 404 2537 476 2543
rect 628 2537 732 2543
rect 756 2537 780 2543
rect 884 2537 972 2543
rect 1028 2537 1052 2543
rect 1060 2537 1116 2543
rect 1540 2537 1564 2543
rect 1764 2537 1820 2543
rect 2564 2537 2812 2543
rect 3108 2537 3212 2543
rect 3236 2537 3244 2543
rect 3332 2537 3436 2543
rect 3444 2537 3500 2543
rect 3572 2537 3628 2543
rect 3636 2537 3676 2543
rect 3844 2537 4156 2543
rect 4164 2537 4300 2543
rect 4628 2537 4684 2543
rect 5028 2537 5132 2543
rect 5860 2537 5891 2543
rect 324 2517 348 2523
rect 836 2517 1132 2523
rect 1508 2517 1548 2523
rect 1556 2517 1692 2523
rect 1780 2517 1788 2523
rect 1796 2517 1868 2523
rect 1876 2517 1900 2523
rect 2132 2517 2156 2523
rect 2596 2517 2636 2523
rect 2644 2517 2684 2523
rect 2692 2517 2972 2523
rect 3044 2517 3228 2523
rect 3252 2517 3340 2523
rect 3380 2517 3564 2523
rect 3620 2517 3660 2523
rect 3812 2517 3900 2523
rect 3988 2517 4092 2523
rect 4388 2517 4412 2523
rect 4420 2517 4508 2523
rect 4676 2517 4716 2523
rect 4756 2517 4860 2523
rect 5092 2517 5148 2523
rect 164 2497 316 2503
rect 324 2497 412 2503
rect 420 2497 460 2503
rect 1620 2497 1772 2503
rect 2756 2497 3132 2503
rect 3220 2497 3228 2503
rect 3252 2497 3340 2503
rect 3460 2497 3532 2503
rect 3540 2497 3644 2503
rect 4436 2497 4540 2503
rect 4548 2497 4684 2503
rect 4868 2497 4892 2503
rect 5604 2497 5891 2503
rect 996 2477 1036 2483
rect 1444 2477 1468 2483
rect 1604 2477 1756 2483
rect 1764 2477 1932 2483
rect 4532 2477 4556 2483
rect 4580 2477 4604 2483
rect 5556 2477 5660 2483
rect 1812 2457 1852 2463
rect 4500 2457 4684 2463
rect 4404 2437 4828 2443
rect 1524 2417 1820 2423
rect 4516 2417 4748 2423
rect 1352 2414 1400 2416
rect 1352 2406 1356 2414
rect 1366 2406 1372 2414
rect 1380 2406 1386 2414
rect 1396 2406 1400 2414
rect 1352 2404 1400 2406
rect 4440 2414 4488 2416
rect 4440 2406 4444 2414
rect 4454 2406 4460 2414
rect 4468 2406 4474 2414
rect 4484 2406 4488 2414
rect 4440 2404 4488 2406
rect 4564 2397 4668 2403
rect 1108 2377 1308 2383
rect 4340 2377 4652 2383
rect 5860 2377 5891 2383
rect 4020 2357 4252 2363
rect 4260 2357 4620 2363
rect 564 2337 844 2343
rect 1300 2337 1564 2343
rect 2116 2337 2380 2343
rect 2980 2337 3276 2343
rect 4308 2337 4428 2343
rect 4564 2337 4764 2343
rect 4772 2337 4988 2343
rect 5332 2337 5891 2343
rect 804 2317 924 2323
rect 1412 2317 1532 2323
rect 2308 2317 2396 2323
rect 3060 2317 3388 2323
rect 4388 2317 4428 2323
rect 4436 2317 4524 2323
rect 4532 2317 4588 2323
rect 4660 2317 4700 2323
rect 4868 2317 4956 2323
rect 5092 2317 5148 2323
rect 5524 2317 5580 2323
rect 388 2297 412 2303
rect 1540 2297 1580 2303
rect 1604 2297 1852 2303
rect 1972 2297 2044 2303
rect 2052 2297 2236 2303
rect 2244 2297 2460 2303
rect 2852 2297 2940 2303
rect 2964 2297 3068 2303
rect 3636 2297 3756 2303
rect 3956 2297 4044 2303
rect 4372 2297 4492 2303
rect 4500 2297 4972 2303
rect 5220 2297 5388 2303
rect 5764 2297 5891 2303
rect 772 2277 812 2283
rect 1220 2277 1516 2283
rect 2388 2277 2492 2283
rect 4932 2277 5116 2283
rect 5124 2277 5548 2283
rect 1108 2257 1820 2263
rect 1828 2257 1836 2263
rect 1844 2257 1948 2263
rect 2820 2257 3020 2263
rect 4356 2257 4380 2263
rect 4388 2257 4444 2263
rect 4596 2257 4796 2263
rect 4964 2257 5020 2263
rect 20 2237 28 2243
rect 804 2237 924 2243
rect 1924 2237 1980 2243
rect 2180 2237 2364 2243
rect 2628 2237 2732 2243
rect 2740 2237 2844 2243
rect 3268 2237 3324 2243
rect 3460 2237 3644 2243
rect 4292 2237 4732 2243
rect 4868 2237 4892 2243
rect 5108 2237 5244 2243
rect 548 2217 652 2223
rect 900 2217 972 2223
rect 1044 2217 1164 2223
rect 3156 2217 3260 2223
rect 4756 2217 4972 2223
rect 2904 2214 2952 2216
rect 2904 2206 2908 2214
rect 2918 2206 2924 2214
rect 2932 2206 2938 2214
rect 2948 2206 2952 2214
rect 2904 2204 2952 2206
rect 532 2197 572 2203
rect 4436 2197 4524 2203
rect 4532 2197 4588 2203
rect 4708 2197 4940 2203
rect 1812 2177 2044 2183
rect 2212 2177 2252 2183
rect 2724 2177 2828 2183
rect 2852 2177 2940 2183
rect 3300 2177 3708 2183
rect 276 2157 348 2163
rect 1652 2157 1740 2163
rect 1748 2157 1884 2163
rect 2932 2157 2988 2163
rect 3364 2157 3420 2163
rect 3812 2157 3932 2163
rect 4580 2157 4652 2163
rect 4660 2157 4764 2163
rect 4772 2157 4876 2163
rect 4916 2157 4988 2163
rect 5252 2157 5292 2163
rect 132 2137 316 2143
rect 324 2137 556 2143
rect 564 2137 700 2143
rect 708 2137 940 2143
rect 948 2137 972 2143
rect 980 2137 1068 2143
rect 1076 2137 1180 2143
rect 1780 2137 1820 2143
rect 1844 2137 1932 2143
rect 1940 2137 2076 2143
rect 2308 2137 2348 2143
rect 2468 2137 2588 2143
rect 3108 2137 3292 2143
rect 3300 2137 3484 2143
rect 3668 2137 3756 2143
rect 4660 2137 4828 2143
rect 4900 2137 4956 2143
rect 4980 2137 5004 2143
rect 5140 2137 5308 2143
rect 5316 2137 5372 2143
rect 1252 2117 1276 2123
rect 1476 2117 1564 2123
rect 1572 2117 1660 2123
rect 1668 2117 1708 2123
rect 1940 2117 1980 2123
rect 2180 2117 2220 2123
rect 2276 2117 2412 2123
rect 2420 2117 2476 2123
rect 2660 2117 2764 2123
rect 2804 2117 2844 2123
rect 3124 2117 3180 2123
rect 3396 2117 3772 2123
rect 3972 2117 3996 2123
rect 4132 2117 4156 2123
rect 4340 2117 4396 2123
rect 4404 2117 4588 2123
rect 4644 2117 4748 2123
rect 4772 2117 4924 2123
rect 4980 2117 5084 2123
rect 5220 2117 5276 2123
rect 5284 2117 5340 2123
rect 1876 2097 1964 2103
rect 2340 2097 2492 2103
rect 2500 2097 2732 2103
rect 2820 2097 2844 2103
rect 3812 2097 3987 2103
rect 1892 2077 2012 2083
rect 2468 2077 2492 2083
rect 2660 2077 2700 2083
rect 3716 2077 3964 2083
rect 3981 2083 3987 2097
rect 4004 2097 4188 2103
rect 4452 2097 4636 2103
rect 4836 2097 4860 2103
rect 5396 2097 5420 2103
rect 5860 2097 5891 2103
rect 3981 2077 4108 2083
rect 4324 2077 4668 2083
rect 4756 2077 4796 2083
rect 4804 2077 5020 2083
rect 5060 2077 5484 2083
rect 5620 2077 5692 2083
rect 2404 2057 2492 2063
rect 4676 2057 4812 2063
rect 404 2037 444 2043
rect 2532 2037 2988 2043
rect 4372 2037 4396 2043
rect 4404 2037 4652 2043
rect 4660 2037 4700 2043
rect 4708 2037 4748 2043
rect 1352 2014 1400 2016
rect 1352 2006 1356 2014
rect 1366 2006 1372 2014
rect 1380 2006 1386 2014
rect 1396 2006 1400 2014
rect 1352 2004 1400 2006
rect 4440 2014 4488 2016
rect 4440 2006 4444 2014
rect 4454 2006 4460 2014
rect 4468 2006 4474 2014
rect 4484 2006 4488 2014
rect 4440 2004 4488 2006
rect 4628 1997 4684 2003
rect 4820 1997 4860 2003
rect 4868 1997 4988 2003
rect 4996 1997 5276 2003
rect 4020 1977 4092 1983
rect 772 1957 876 1963
rect 884 1957 1212 1963
rect 1876 1957 1900 1963
rect 1988 1957 2236 1963
rect 356 1937 428 1943
rect 2036 1937 2300 1943
rect 3076 1937 3212 1943
rect 436 1917 492 1923
rect 500 1917 556 1923
rect 692 1917 780 1923
rect 868 1917 1100 1923
rect 1924 1917 1996 1923
rect 2180 1917 2268 1923
rect 2564 1917 3020 1923
rect 3044 1917 3116 1923
rect 4532 1917 4540 1923
rect 5124 1917 5148 1923
rect 5156 1917 5180 1923
rect 5204 1917 5484 1923
rect 404 1897 636 1903
rect 660 1897 668 1903
rect 676 1897 940 1903
rect 1300 1897 1436 1903
rect 1476 1897 1516 1903
rect 1812 1897 1916 1903
rect 2180 1897 2796 1903
rect 3732 1897 3772 1903
rect 3828 1897 3852 1903
rect 3940 1897 4076 1903
rect 4308 1897 4332 1903
rect 4388 1897 4540 1903
rect 4548 1897 4620 1903
rect 4788 1897 4876 1903
rect 5172 1897 5388 1903
rect 5588 1897 5708 1903
rect 452 1877 636 1883
rect 644 1877 716 1883
rect 980 1877 988 1883
rect 996 1877 1036 1883
rect 1092 1877 1132 1883
rect 1940 1877 2044 1883
rect 2468 1877 2588 1883
rect 3092 1877 3324 1883
rect 3428 1877 3548 1883
rect 3892 1877 4060 1883
rect 4532 1877 4636 1883
rect 4644 1877 4764 1883
rect 4820 1877 4924 1883
rect 4948 1877 4972 1883
rect 4980 1877 5084 1883
rect 5332 1877 5420 1883
rect 5492 1877 5644 1883
rect 196 1857 252 1863
rect 388 1857 460 1863
rect 468 1857 508 1863
rect 516 1857 604 1863
rect 612 1857 732 1863
rect 740 1857 748 1863
rect 756 1857 780 1863
rect 1085 1863 1091 1876
rect 932 1857 1091 1863
rect 1732 1857 1980 1863
rect 1988 1857 2124 1863
rect 2436 1857 2572 1863
rect 2580 1857 2684 1863
rect 2932 1857 3100 1863
rect 3140 1857 3228 1863
rect 3332 1857 3436 1863
rect 3796 1857 3916 1863
rect 4612 1857 4652 1863
rect 4772 1857 4940 1863
rect 4948 1857 5132 1863
rect 5140 1857 5212 1863
rect 5220 1857 5244 1863
rect 5268 1857 5324 1863
rect 5332 1857 5356 1863
rect 36 1837 188 1843
rect 276 1837 380 1843
rect 1460 1837 1500 1843
rect 1844 1837 2108 1843
rect 2740 1837 3148 1843
rect 3156 1837 3356 1843
rect 3524 1837 4204 1843
rect 4756 1837 4844 1843
rect 4852 1837 4892 1843
rect 4932 1837 5164 1843
rect 5604 1837 5660 1843
rect 1540 1817 1724 1823
rect 1732 1817 1852 1823
rect 3924 1817 3996 1823
rect 4260 1817 4588 1823
rect 4868 1817 4988 1823
rect 5092 1817 5340 1823
rect 5668 1817 5836 1823
rect 2904 1814 2952 1816
rect 2904 1806 2908 1814
rect 2918 1806 2924 1814
rect 2932 1806 2938 1814
rect 2948 1806 2952 1814
rect 2904 1804 2952 1806
rect 1828 1797 2524 1803
rect 3268 1797 3436 1803
rect 3444 1797 3612 1803
rect 3748 1797 4140 1803
rect 4580 1797 4764 1803
rect 5044 1797 5324 1803
rect 5332 1797 5404 1803
rect 244 1777 396 1783
rect 932 1777 1020 1783
rect 1876 1777 1932 1783
rect 1940 1777 2044 1783
rect 3092 1777 3132 1783
rect 3140 1777 3411 1783
rect 3405 1764 3411 1777
rect 3748 1777 3900 1783
rect 3908 1777 4012 1783
rect 4020 1777 4044 1783
rect 5012 1777 5068 1783
rect 5316 1777 5564 1783
rect 132 1757 140 1763
rect 260 1757 300 1763
rect 532 1757 556 1763
rect 612 1757 828 1763
rect 1860 1757 2076 1763
rect 2116 1757 2172 1763
rect 3220 1757 3324 1763
rect 3412 1757 3452 1763
rect 3636 1757 3964 1763
rect 5028 1757 5100 1763
rect 5124 1757 5148 1763
rect 5188 1757 5228 1763
rect 5252 1757 5292 1763
rect 5348 1757 5436 1763
rect 548 1737 700 1743
rect 756 1737 940 1743
rect 1124 1737 1244 1743
rect 1460 1737 1548 1743
rect 1844 1737 1900 1743
rect 1908 1737 1996 1743
rect 2004 1737 2012 1743
rect 2125 1737 2220 1743
rect 340 1717 380 1723
rect 477 1723 483 1736
rect 2125 1724 2131 1737
rect 2660 1737 2684 1743
rect 2692 1737 2924 1743
rect 3252 1737 3484 1743
rect 3572 1737 3580 1743
rect 3620 1737 3660 1743
rect 3732 1737 3772 1743
rect 4196 1737 4460 1743
rect 4916 1737 5308 1743
rect 5396 1737 5436 1743
rect 420 1717 483 1723
rect 580 1717 604 1723
rect 660 1717 700 1723
rect 884 1717 1100 1723
rect 1332 1717 1580 1723
rect 1828 1717 1868 1723
rect 2036 1717 2124 1723
rect 2164 1717 2204 1723
rect 2212 1717 2268 1723
rect 2276 1717 2380 1723
rect 3204 1717 3372 1723
rect 3540 1717 3644 1723
rect 3652 1717 3820 1723
rect 3828 1717 3868 1723
rect 3908 1717 4012 1723
rect 4068 1717 4092 1723
rect 4116 1717 4204 1723
rect 4532 1717 4620 1723
rect 5044 1717 5084 1723
rect 5092 1717 5180 1723
rect 5453 1723 5459 1736
rect 5316 1717 5459 1723
rect 596 1697 812 1703
rect 820 1697 1196 1703
rect 1204 1697 1276 1703
rect 1828 1697 1852 1703
rect 1988 1697 2156 1703
rect 2164 1697 2236 1703
rect 2308 1697 2716 1703
rect 2996 1697 3068 1703
rect 3076 1697 3180 1703
rect 3220 1697 3260 1703
rect 3364 1697 3420 1703
rect 3492 1697 3516 1703
rect 3620 1697 3740 1703
rect 3812 1697 3884 1703
rect 3892 1697 3932 1703
rect 3972 1697 3996 1703
rect 4996 1697 5052 1703
rect 5060 1697 5084 1703
rect 5124 1697 5196 1703
rect 5284 1697 5308 1703
rect 5316 1697 5468 1703
rect 5860 1697 5891 1703
rect 500 1677 780 1683
rect 2212 1677 2316 1683
rect 2852 1677 3308 1683
rect 3316 1677 3468 1683
rect 3700 1677 3772 1683
rect 3780 1677 3852 1683
rect 3860 1677 3916 1683
rect 3924 1677 4060 1683
rect 5108 1677 5132 1683
rect 5172 1677 5292 1683
rect 5380 1677 5500 1683
rect 452 1657 1388 1663
rect 1796 1657 2956 1663
rect 3572 1657 3756 1663
rect 5284 1657 5372 1663
rect 5396 1657 5452 1663
rect 1012 1637 1100 1643
rect 2484 1637 2508 1643
rect 5156 1637 5356 1643
rect 5476 1637 5516 1643
rect 5540 1637 5708 1643
rect 1044 1617 1116 1623
rect 1716 1617 2684 1623
rect 5252 1617 5372 1623
rect 5412 1617 5532 1623
rect 1352 1614 1400 1616
rect 1352 1606 1356 1614
rect 1366 1606 1372 1614
rect 1380 1606 1386 1614
rect 1396 1606 1400 1614
rect 1352 1604 1400 1606
rect 4440 1614 4488 1616
rect 4440 1606 4444 1614
rect 4454 1606 4460 1614
rect 4468 1606 4474 1614
rect 4484 1606 4488 1614
rect 4440 1604 4488 1606
rect 3988 1597 4028 1603
rect 5140 1597 5516 1603
rect 196 1577 332 1583
rect 1236 1577 2444 1583
rect 3764 1577 3980 1583
rect 3988 1577 4172 1583
rect 4484 1577 4556 1583
rect 4868 1577 4908 1583
rect 5316 1577 5340 1583
rect 244 1557 268 1563
rect 1092 1557 1884 1563
rect 3252 1557 3708 1563
rect 3716 1557 3756 1563
rect 3764 1557 3804 1563
rect 4212 1557 4636 1563
rect 5060 1557 5196 1563
rect 5204 1557 5260 1563
rect 132 1537 220 1543
rect 500 1537 636 1543
rect 1044 1537 1068 1543
rect 1108 1537 1420 1543
rect 2404 1537 2988 1543
rect 3460 1537 3644 1543
rect 3652 1537 3692 1543
rect 3748 1537 3804 1543
rect 4052 1537 4396 1543
rect 5332 1537 5388 1543
rect 132 1517 316 1523
rect 372 1517 556 1523
rect 756 1517 1580 1523
rect 2100 1517 2252 1523
rect 2532 1517 3324 1523
rect 3524 1517 3740 1523
rect 3860 1517 4156 1523
rect 4164 1517 4508 1523
rect 4628 1517 4732 1523
rect 5140 1517 5228 1523
rect 5236 1517 5276 1523
rect 84 1497 108 1503
rect 116 1497 156 1503
rect 164 1497 204 1503
rect 292 1497 332 1503
rect 420 1497 476 1503
rect 500 1497 604 1503
rect 868 1497 972 1503
rect 996 1497 1068 1503
rect 1076 1497 1148 1503
rect 1156 1497 1260 1503
rect 1652 1497 1724 1503
rect 2468 1497 2556 1503
rect 2564 1497 2636 1503
rect 2644 1497 2668 1503
rect 2820 1497 3180 1503
rect 3492 1497 3644 1503
rect 3684 1497 3884 1503
rect 4100 1497 4124 1503
rect 4292 1497 4588 1503
rect 4676 1497 4732 1503
rect 4788 1497 4876 1503
rect 4884 1497 4924 1503
rect 5076 1497 5164 1503
rect 5252 1497 5292 1503
rect 5348 1497 5404 1503
rect 5444 1497 5484 1503
rect 100 1477 140 1483
rect 324 1477 684 1483
rect 836 1477 892 1483
rect 1325 1477 1340 1483
rect 196 1457 380 1463
rect 404 1457 460 1463
rect 468 1457 588 1463
rect 596 1457 620 1463
rect 676 1457 780 1463
rect 980 1457 1036 1463
rect 1325 1463 1331 1477
rect 1972 1477 2076 1483
rect 2084 1477 2236 1483
rect 2292 1477 2316 1483
rect 2580 1477 2716 1483
rect 3556 1477 3724 1483
rect 3732 1477 3756 1483
rect 3812 1477 3868 1483
rect 3908 1477 4108 1483
rect 4260 1477 4284 1483
rect 4676 1477 4748 1483
rect 4996 1477 5004 1483
rect 5268 1477 5340 1483
rect 5412 1477 5436 1483
rect 5636 1477 5708 1483
rect 1220 1457 1331 1463
rect 1348 1457 1468 1463
rect 1524 1457 1932 1463
rect 1940 1457 1980 1463
rect 1988 1457 2140 1463
rect 2148 1457 2316 1463
rect 2452 1457 2588 1463
rect 2644 1457 2700 1463
rect 2708 1457 2748 1463
rect 3316 1457 3372 1463
rect 3380 1457 3468 1463
rect 3476 1457 3580 1463
rect 3588 1457 3628 1463
rect 3748 1457 3820 1463
rect 3869 1463 3875 1476
rect 3869 1457 3948 1463
rect 4116 1457 4204 1463
rect 4324 1457 4444 1463
rect 5172 1457 5324 1463
rect 5364 1457 5404 1463
rect 5428 1457 5516 1463
rect 5524 1457 5532 1463
rect 196 1437 412 1443
rect 452 1437 556 1443
rect 612 1437 652 1443
rect 900 1437 1228 1443
rect 1588 1437 1628 1443
rect 2212 1437 2284 1443
rect 2596 1437 2652 1443
rect 2804 1437 2876 1443
rect 3572 1437 3804 1443
rect 3860 1437 4012 1443
rect 4100 1437 4108 1443
rect 4292 1437 4332 1443
rect 260 1417 348 1423
rect 356 1417 476 1423
rect 756 1417 988 1423
rect 996 1417 1276 1423
rect 1284 1417 1356 1423
rect 1364 1417 1836 1423
rect 2068 1417 2780 1423
rect 3124 1417 3260 1423
rect 3268 1417 3484 1423
rect 3524 1417 3628 1423
rect 4148 1417 4316 1423
rect 4564 1417 4620 1423
rect 5236 1417 5484 1423
rect 5508 1417 5532 1423
rect 2904 1414 2952 1416
rect 2904 1406 2908 1414
rect 2918 1406 2924 1414
rect 2932 1406 2938 1414
rect 2948 1406 2952 1414
rect 2904 1404 2952 1406
rect 292 1397 332 1403
rect 628 1397 908 1403
rect 2244 1397 2268 1403
rect 3748 1397 4268 1403
rect 4388 1397 4508 1403
rect 5108 1397 5660 1403
rect 148 1377 300 1383
rect 868 1377 908 1383
rect 932 1377 1180 1383
rect 2020 1377 2252 1383
rect 2772 1377 2812 1383
rect 3428 1377 3436 1383
rect 3652 1377 3692 1383
rect 3716 1377 3836 1383
rect 3876 1377 4044 1383
rect 4276 1377 4300 1383
rect 4452 1377 4540 1383
rect 5220 1377 5564 1383
rect 20 1357 76 1363
rect 244 1357 332 1363
rect 340 1357 380 1363
rect 692 1357 700 1363
rect 708 1357 828 1363
rect 1108 1357 1468 1363
rect 1492 1357 1564 1363
rect 1940 1357 1980 1363
rect 1988 1357 2060 1363
rect 2276 1357 2300 1363
rect 2516 1357 2956 1363
rect 3588 1357 3676 1363
rect 3684 1357 3772 1363
rect 3796 1357 3868 1363
rect 3876 1357 3884 1363
rect 4004 1357 4483 1363
rect 52 1337 284 1343
rect 772 1337 924 1343
rect 932 1337 1164 1343
rect 1268 1337 1308 1343
rect 1796 1337 1836 1343
rect 1844 1337 1964 1343
rect 2148 1337 2156 1343
rect 2244 1337 2284 1343
rect 2324 1337 2380 1343
rect 2564 1337 2620 1343
rect 2628 1337 2652 1343
rect 2692 1337 2812 1343
rect 2948 1337 3052 1343
rect 3364 1337 3484 1343
rect 3620 1337 3676 1343
rect 3684 1337 3724 1343
rect 3757 1337 3900 1343
rect 244 1317 444 1323
rect 580 1317 620 1323
rect 788 1317 940 1323
rect 1092 1317 1132 1323
rect 1156 1317 1260 1323
rect 1572 1317 1644 1323
rect 1716 1317 1820 1323
rect 1828 1317 1884 1323
rect 1892 1317 1932 1323
rect 1940 1317 2156 1323
rect 2221 1317 2348 1323
rect 2221 1304 2227 1317
rect 2452 1317 2476 1323
rect 2484 1317 2844 1323
rect 2852 1317 2988 1323
rect 2996 1317 3180 1323
rect 3757 1323 3763 1337
rect 3908 1337 3980 1343
rect 3988 1337 4204 1343
rect 4477 1343 4483 1357
rect 4500 1357 4668 1363
rect 5325 1357 5772 1363
rect 5325 1344 5331 1357
rect 4477 1337 4684 1343
rect 4916 1337 5132 1343
rect 5140 1337 5324 1343
rect 5396 1337 5436 1343
rect 5444 1337 5500 1343
rect 3556 1317 3763 1323
rect 3860 1317 3996 1323
rect 4180 1317 4300 1323
rect 4356 1317 4412 1323
rect 4420 1317 4572 1323
rect 4724 1317 4748 1323
rect 308 1297 380 1303
rect 388 1297 412 1303
rect 420 1297 524 1303
rect 548 1297 572 1303
rect 660 1297 796 1303
rect 804 1297 812 1303
rect 820 1297 1116 1303
rect 1124 1297 1196 1303
rect 1204 1297 1484 1303
rect 1860 1297 2012 1303
rect 2116 1297 2188 1303
rect 2196 1297 2220 1303
rect 2244 1297 2316 1303
rect 2324 1297 2524 1303
rect 2692 1297 2716 1303
rect 2884 1297 2892 1303
rect 3444 1297 3804 1303
rect 3812 1297 4156 1303
rect 4660 1297 4716 1303
rect 5268 1297 5356 1303
rect 5380 1297 5436 1303
rect 20 1277 252 1283
rect 644 1277 892 1283
rect 900 1277 972 1283
rect 1188 1277 1276 1283
rect 2116 1277 2460 1283
rect 2532 1277 3116 1283
rect 3572 1277 3580 1283
rect 3668 1277 3932 1283
rect 3972 1277 4076 1283
rect 4084 1277 4348 1283
rect 4372 1277 4764 1283
rect 5124 1277 5164 1283
rect 5172 1277 5388 1283
rect 148 1257 220 1263
rect 964 1257 1116 1263
rect 3332 1257 4188 1263
rect 884 1237 1148 1243
rect 3028 1237 3132 1243
rect 5332 1237 5404 1243
rect 5412 1237 5484 1243
rect 1028 1217 1052 1223
rect 2148 1217 2268 1223
rect 2516 1217 2700 1223
rect 2708 1217 2748 1223
rect 2756 1217 3100 1223
rect 1352 1214 1400 1216
rect 1352 1206 1356 1214
rect 1366 1206 1372 1214
rect 1380 1206 1386 1214
rect 1396 1206 1400 1214
rect 1352 1204 1400 1206
rect 4440 1214 4488 1216
rect 4440 1206 4444 1214
rect 4454 1206 4460 1214
rect 4468 1206 4474 1214
rect 4484 1206 4488 1214
rect 4440 1204 4488 1206
rect 708 1197 732 1203
rect 740 1197 1020 1203
rect 1780 1197 2748 1203
rect 2756 1197 2764 1203
rect 4004 1197 4060 1203
rect 4324 1197 4332 1203
rect 484 1177 508 1183
rect 532 1177 828 1183
rect 1156 1177 1308 1183
rect 1316 1177 1516 1183
rect 2020 1177 2076 1183
rect 2244 1177 2268 1183
rect 2292 1177 2652 1183
rect 3812 1177 4316 1183
rect 4500 1177 4540 1183
rect 5092 1177 5132 1183
rect 5140 1177 5676 1183
rect 5796 1177 5820 1183
rect 132 1157 540 1163
rect 1092 1157 1372 1163
rect 2100 1157 2124 1163
rect 2132 1157 2732 1163
rect 4148 1157 4172 1163
rect 4324 1157 4796 1163
rect 5284 1157 5372 1163
rect 420 1137 652 1143
rect 788 1137 1692 1143
rect 1828 1137 2620 1143
rect 2900 1137 3324 1143
rect 3636 1137 3884 1143
rect 3892 1137 3948 1143
rect 3956 1137 4060 1143
rect 4740 1137 4764 1143
rect 5348 1137 5452 1143
rect 68 1117 108 1123
rect 372 1117 492 1123
rect 756 1117 764 1123
rect 852 1117 892 1123
rect 900 1117 924 1123
rect 932 1117 972 1123
rect 989 1117 1116 1123
rect 989 1104 995 1117
rect 1220 1117 1340 1123
rect 1940 1117 1964 1123
rect 2052 1117 2076 1123
rect 2180 1117 2428 1123
rect 2660 1117 2780 1123
rect 3716 1117 3900 1123
rect 4084 1117 4124 1123
rect 4596 1117 4604 1123
rect 4868 1117 5292 1123
rect 5636 1117 5692 1123
rect 20 1097 76 1103
rect 340 1097 380 1103
rect 452 1097 499 1103
rect 36 1077 220 1083
rect 340 1077 364 1083
rect 372 1077 412 1083
rect 436 1077 476 1083
rect 493 1083 499 1097
rect 516 1097 636 1103
rect 900 1097 988 1103
rect 1060 1097 1084 1103
rect 1284 1097 1484 1103
rect 1492 1097 1564 1103
rect 1924 1097 2108 1103
rect 2244 1097 2412 1103
rect 2420 1097 2684 1103
rect 2756 1097 2828 1103
rect 2836 1097 2972 1103
rect 3524 1097 3596 1103
rect 3764 1097 4092 1103
rect 4132 1097 4172 1103
rect 4244 1097 4364 1103
rect 4388 1097 4620 1103
rect 4740 1097 5084 1103
rect 5220 1097 5276 1103
rect 5524 1097 5596 1103
rect 493 1077 540 1083
rect 548 1077 643 1083
rect 68 1057 156 1063
rect 356 1057 604 1063
rect 637 1063 643 1077
rect 660 1077 684 1083
rect 724 1077 812 1083
rect 884 1077 1036 1083
rect 1044 1077 1276 1083
rect 1956 1077 2012 1083
rect 2052 1077 2092 1083
rect 2100 1077 2236 1083
rect 2260 1077 2332 1083
rect 2404 1077 2556 1083
rect 2644 1077 2716 1083
rect 2724 1077 2764 1083
rect 3156 1077 3292 1083
rect 3668 1077 3868 1083
rect 3876 1077 3964 1083
rect 4116 1077 4140 1083
rect 5444 1077 5468 1083
rect 5476 1077 5500 1083
rect 5556 1077 5628 1083
rect 5636 1077 5660 1083
rect 637 1057 652 1063
rect 836 1057 892 1063
rect 900 1057 924 1063
rect 932 1057 940 1063
rect 996 1057 1020 1063
rect 1028 1057 1100 1063
rect 1364 1057 1436 1063
rect 1460 1057 1500 1063
rect 1604 1057 1628 1063
rect 2244 1057 2300 1063
rect 2740 1057 2812 1063
rect 3796 1057 3820 1063
rect 4100 1057 4300 1063
rect 4628 1057 4780 1063
rect 292 1037 332 1043
rect 1028 1037 1052 1043
rect 2020 1037 2188 1043
rect 2196 1037 2348 1043
rect 2356 1037 2428 1043
rect 2436 1037 2572 1043
rect 2596 1037 2828 1043
rect 2861 1037 2924 1043
rect 36 1017 92 1023
rect 100 1017 188 1023
rect 228 1017 460 1023
rect 868 1017 1468 1023
rect 2212 1017 2604 1023
rect 2861 1023 2867 1037
rect 3572 1037 3820 1043
rect 4180 1037 4668 1043
rect 4676 1037 4812 1043
rect 4820 1037 5356 1043
rect 5412 1037 5468 1043
rect 2660 1017 2867 1023
rect 3268 1017 3564 1023
rect 3796 1017 3964 1023
rect 3972 1017 3980 1023
rect 3988 1017 4060 1023
rect 4628 1017 4892 1023
rect 5300 1017 5372 1023
rect 5780 1017 5836 1023
rect 2904 1014 2952 1016
rect 2904 1006 2908 1014
rect 2918 1006 2924 1014
rect 2932 1006 2938 1014
rect 2948 1006 2952 1014
rect 2904 1004 2952 1006
rect 36 997 140 1003
rect 1156 997 1244 1003
rect 1972 997 2124 1003
rect 2132 997 2204 1003
rect 3828 997 4524 1003
rect 4532 997 4588 1003
rect 4596 997 4668 1003
rect 1012 977 1020 983
rect 1060 977 1340 983
rect 1348 977 1452 983
rect 1844 977 1900 983
rect 1908 977 1964 983
rect 1972 977 2028 983
rect 2036 977 2172 983
rect 2180 977 2188 983
rect 2308 977 2332 983
rect 2692 977 2748 983
rect 2756 977 3036 983
rect 3668 977 3884 983
rect 3892 977 3948 983
rect 4244 977 4636 983
rect 4644 977 4684 983
rect 4772 977 4780 983
rect 532 957 572 963
rect 596 957 732 963
rect 948 957 988 963
rect 1012 957 1084 963
rect 1220 957 1308 963
rect 1764 957 1804 963
rect 1812 957 1836 963
rect 1876 957 2460 963
rect 2788 957 2828 963
rect 2836 957 3004 963
rect 3012 957 3292 963
rect 3572 957 3788 963
rect 3860 957 3900 963
rect 3908 957 4092 963
rect 4276 957 4652 963
rect 4740 957 4796 963
rect 276 937 348 943
rect 356 937 380 943
rect 420 937 604 943
rect 660 937 700 943
rect 852 937 892 943
rect 916 937 972 943
rect 980 937 1228 943
rect 1236 937 1404 943
rect 1444 937 1628 943
rect 1956 937 2012 943
rect 2036 937 2076 943
rect 2180 937 2364 943
rect 2564 937 2668 943
rect 2932 937 2972 943
rect 2980 937 2988 943
rect 3028 937 3068 943
rect 3588 937 3980 943
rect 4196 937 4300 943
rect 5428 937 5548 943
rect 5860 937 5891 943
rect 116 917 124 923
rect 308 917 364 923
rect 628 917 684 923
rect 820 917 956 923
rect 996 917 1052 923
rect 1092 917 1244 923
rect 1252 917 1532 923
rect 1780 917 1980 923
rect 2340 917 2412 923
rect 2452 917 2476 923
rect 2964 917 3020 923
rect 3028 917 3036 923
rect 3236 917 3420 923
rect 3684 917 3900 923
rect 3924 917 4076 923
rect 4228 917 4604 923
rect 5044 917 5180 923
rect 324 897 508 903
rect 516 897 716 903
rect 740 897 764 903
rect 788 897 844 903
rect 1133 897 1436 903
rect 340 877 380 883
rect 388 877 540 883
rect 1133 883 1139 897
rect 1460 897 1468 903
rect 1476 897 1500 903
rect 1956 897 2156 903
rect 2244 897 2348 903
rect 2404 897 2540 903
rect 2612 897 3164 903
rect 3828 897 3852 903
rect 3860 897 4028 903
rect 4148 897 4188 903
rect 4228 897 4252 903
rect 5764 897 5891 903
rect 756 877 1139 883
rect 1156 877 1468 883
rect 1764 877 2028 883
rect 2228 877 2572 883
rect 2772 877 2828 883
rect 2916 877 3356 883
rect 3780 877 3916 883
rect 3956 877 4012 883
rect 4132 877 4364 883
rect 4692 877 4972 883
rect 5252 877 5292 883
rect 5492 877 5580 883
rect 484 857 572 863
rect 1220 857 1564 863
rect 2196 857 2492 863
rect 4852 857 4876 863
rect 2004 837 2252 843
rect 4836 837 5036 843
rect 180 817 300 823
rect 1028 817 1212 823
rect 1908 817 2172 823
rect 4100 817 4332 823
rect 1352 814 1400 816
rect 1352 806 1356 814
rect 1366 806 1372 814
rect 1380 806 1386 814
rect 1396 806 1400 814
rect 1352 804 1400 806
rect 4440 814 4488 816
rect 4440 806 4444 814
rect 4454 806 4460 814
rect 4468 806 4474 814
rect 4484 806 4488 814
rect 4440 804 4488 806
rect 148 797 348 803
rect 356 797 1036 803
rect 212 777 284 783
rect 420 777 780 783
rect 3620 777 4236 783
rect 4244 777 4268 783
rect 100 757 268 763
rect 404 757 668 763
rect 772 757 828 763
rect 4148 757 4796 763
rect 132 737 236 743
rect 260 737 732 743
rect 740 737 796 743
rect 836 737 1132 743
rect 1140 737 1308 743
rect 1316 737 1372 743
rect 1748 737 1868 743
rect 1876 737 2204 743
rect 2292 737 2444 743
rect 2708 737 3164 743
rect 3300 737 4236 743
rect 4244 737 4380 743
rect 4612 737 4636 743
rect 4788 737 4940 743
rect 132 717 156 723
rect 164 717 172 723
rect 324 717 444 723
rect 676 717 748 723
rect 756 717 764 723
rect 1028 717 1052 723
rect 2116 717 2435 723
rect 132 697 140 703
rect 148 697 188 703
rect 436 697 508 703
rect 564 697 620 703
rect 1172 697 1228 703
rect 1428 697 1596 703
rect 1828 697 1884 703
rect 1892 697 1932 703
rect 2068 697 2188 703
rect 2429 703 2435 717
rect 2452 717 2508 723
rect 2548 717 2604 723
rect 2612 717 2844 723
rect 2868 717 3068 723
rect 3092 717 3676 723
rect 4004 717 4060 723
rect 4068 717 4140 723
rect 4292 717 4748 723
rect 4788 717 4796 723
rect 4964 717 5244 723
rect 5252 717 5324 723
rect 5604 717 5660 723
rect 2429 697 2460 703
rect 2548 697 2588 703
rect 2884 697 2988 703
rect 3044 697 3068 703
rect 3092 697 3116 703
rect 3236 697 3292 703
rect 3956 697 4076 703
rect 4084 697 4108 703
rect 4324 697 4380 703
rect 4388 697 4524 703
rect 4596 697 4604 703
rect 4980 697 4988 703
rect 5076 697 5180 703
rect 5860 697 5891 703
rect 180 677 364 683
rect 509 683 515 696
rect 509 677 604 683
rect 628 677 764 683
rect 932 677 956 683
rect 964 677 972 683
rect 1028 677 1740 683
rect 1876 677 1964 683
rect 1972 677 2028 683
rect 2244 677 2268 683
rect 2292 677 2396 683
rect 2445 677 2492 683
rect 84 657 156 663
rect 164 657 220 663
rect 228 657 316 663
rect 365 663 371 676
rect 365 657 860 663
rect 868 657 940 663
rect 1044 657 1068 663
rect 1076 657 1132 663
rect 1140 657 1532 663
rect 1540 657 1644 663
rect 1741 663 1747 676
rect 1741 657 1804 663
rect 1812 657 1980 663
rect 2068 657 2140 663
rect 2445 663 2451 677
rect 2692 677 2812 683
rect 2836 677 3084 683
rect 3092 677 3324 683
rect 3540 677 3644 683
rect 3812 677 3900 683
rect 3908 677 3964 683
rect 4388 677 4556 683
rect 4596 677 4780 683
rect 4852 677 4924 683
rect 4996 677 5052 683
rect 5092 677 5100 683
rect 5156 677 5196 683
rect 5316 677 5404 683
rect 5412 677 5532 683
rect 2164 657 2451 663
rect 2468 657 2556 663
rect 2628 657 2636 663
rect 2644 657 2828 663
rect 2852 657 3036 663
rect 3044 657 3068 663
rect 3085 657 3196 663
rect 324 637 380 643
rect 516 637 636 643
rect 1060 637 1100 643
rect 1108 637 1212 643
rect 1236 637 1436 643
rect 1444 637 1500 643
rect 1508 637 1532 643
rect 1844 637 1916 643
rect 1924 637 1964 643
rect 2132 637 2204 643
rect 2212 637 2268 643
rect 2388 637 2444 643
rect 2484 637 2620 643
rect 2628 637 2732 643
rect 2820 637 2860 643
rect 2877 637 2995 643
rect 212 617 428 623
rect 436 617 556 623
rect 564 617 796 623
rect 1092 617 1132 623
rect 1156 617 1180 623
rect 1204 617 1404 623
rect 1412 617 1468 623
rect 1492 617 1660 623
rect 1668 617 1788 623
rect 2877 623 2883 637
rect 2068 617 2883 623
rect 2989 623 2995 637
rect 3012 637 3020 643
rect 3085 643 3091 657
rect 3220 657 3276 663
rect 4276 657 4300 663
rect 4308 657 4348 663
rect 4548 657 4620 663
rect 4724 657 4764 663
rect 4788 657 4844 663
rect 4852 657 4972 663
rect 5108 657 5148 663
rect 5204 657 5292 663
rect 3044 637 3091 643
rect 3108 637 3244 643
rect 3300 637 3340 643
rect 4212 637 4364 643
rect 4372 637 4412 643
rect 4932 637 5004 643
rect 5012 637 5036 643
rect 5412 637 5420 643
rect 2989 617 3484 623
rect 4132 617 4732 623
rect 4740 617 4780 623
rect 2904 614 2952 616
rect 2904 606 2908 614
rect 2918 606 2924 614
rect 2932 606 2938 614
rect 2948 606 2952 614
rect 2904 604 2952 606
rect 100 597 332 603
rect 1284 597 1292 603
rect 1300 597 1347 603
rect 36 577 108 583
rect 116 577 252 583
rect 308 577 412 583
rect 420 577 860 583
rect 980 577 1324 583
rect 1341 583 1347 597
rect 1476 597 1500 603
rect 1572 597 1660 603
rect 2740 597 2780 603
rect 2820 597 2876 603
rect 3012 597 3420 603
rect 3812 597 3900 603
rect 3908 597 4012 603
rect 4228 597 4236 603
rect 4244 597 4508 603
rect 1341 577 1436 583
rect 2036 577 2156 583
rect 2164 577 2332 583
rect 2404 577 2428 583
rect 2436 577 2604 583
rect 2676 577 2780 583
rect 2820 577 3756 583
rect 4356 577 4396 583
rect 4404 577 4524 583
rect 4564 577 4604 583
rect 4804 577 4892 583
rect 4916 577 4956 583
rect 4964 577 5228 583
rect 5524 577 5628 583
rect 292 557 364 563
rect 388 557 540 563
rect 628 557 668 563
rect 788 557 812 563
rect 868 557 1100 563
rect 1108 557 1164 563
rect 1316 557 1516 563
rect 2180 557 2236 563
rect 2244 557 2412 563
rect 2772 557 3004 563
rect 3076 557 3164 563
rect 3268 557 3379 563
rect 132 537 236 543
rect 356 537 892 543
rect 900 537 956 543
rect 964 537 1020 543
rect 1124 537 1228 543
rect 1268 537 1756 543
rect 1988 537 2092 543
rect 2212 537 2508 543
rect 2516 537 2556 543
rect 2596 537 2812 543
rect 2836 537 2924 543
rect 3044 537 3052 543
rect 3092 537 3148 543
rect 3156 537 3228 543
rect 3373 543 3379 557
rect 3396 557 3484 563
rect 3700 557 3852 563
rect 3860 557 3964 563
rect 3972 557 4124 563
rect 4164 557 4332 563
rect 4340 557 4380 563
rect 4580 557 4700 563
rect 4868 557 5084 563
rect 5092 557 5116 563
rect 3373 537 3404 543
rect 3860 537 3996 543
rect 4500 537 4588 543
rect 4644 537 4684 543
rect 4692 537 4716 543
rect 4868 537 4940 543
rect 4980 537 5004 543
rect 5604 537 5724 543
rect 20 517 92 523
rect 148 517 204 523
rect 292 517 380 523
rect 404 517 684 523
rect 756 517 780 523
rect 916 517 1148 523
rect 1188 517 1468 523
rect 1732 517 1820 523
rect 2180 517 2300 523
rect 2308 517 2348 523
rect 2532 517 2588 523
rect 2596 517 2636 523
rect 2772 517 2828 523
rect 2836 517 3212 523
rect 3220 517 3308 523
rect 3332 517 3388 523
rect 3476 517 3564 523
rect 4388 517 4812 523
rect 4820 517 4876 523
rect 4884 517 5116 523
rect 5124 517 5212 523
rect 5364 517 5500 523
rect 5572 517 5692 523
rect 196 497 236 503
rect 244 497 348 503
rect 500 497 508 503
rect 564 497 844 503
rect 852 497 988 503
rect 996 497 1052 503
rect 1060 497 1292 503
rect 2564 497 2780 503
rect 3380 497 3436 503
rect 3444 497 3500 503
rect 4308 497 4572 503
rect 4580 497 4652 503
rect 4692 497 4764 503
rect 4932 497 4956 503
rect 4964 497 5036 503
rect 5172 497 5276 503
rect 5508 497 5564 503
rect 436 477 764 483
rect 1012 477 1244 483
rect 1940 477 2652 483
rect 2692 477 3276 483
rect 3284 477 3484 483
rect 3892 477 3948 483
rect 3956 477 4172 483
rect 4532 477 4636 483
rect 4644 477 4844 483
rect 5028 477 5100 483
rect 884 457 1564 463
rect 1572 457 1740 463
rect 1748 457 1996 463
rect 2084 457 2108 463
rect 2116 457 2700 463
rect 2788 457 3132 463
rect 4484 457 4508 463
rect 1780 437 2524 443
rect 2660 437 4028 443
rect 4372 437 4700 443
rect 5444 437 5532 443
rect 5540 437 5580 443
rect 1540 417 1980 423
rect 2884 417 3180 423
rect 3188 417 3564 423
rect 1352 414 1400 416
rect 1352 406 1356 414
rect 1366 406 1372 414
rect 1380 406 1386 414
rect 1396 406 1400 414
rect 1352 404 1400 406
rect 4440 414 4488 416
rect 4440 406 4444 414
rect 4454 406 4460 414
rect 4468 406 4474 414
rect 4484 406 4488 414
rect 4440 404 4488 406
rect 1764 397 1836 403
rect 2548 397 3164 403
rect 3188 397 3292 403
rect 4196 397 4419 403
rect 692 377 732 383
rect 996 377 1580 383
rect 1652 377 2188 383
rect 2484 377 2668 383
rect 2676 377 3036 383
rect 3508 377 3548 383
rect 4260 377 4316 383
rect 4413 383 4419 397
rect 4724 397 4940 403
rect 5076 397 5196 403
rect 4413 377 4588 383
rect 4612 377 4732 383
rect 4772 377 4796 383
rect 4804 377 4860 383
rect 4884 377 4988 383
rect 308 357 531 363
rect 525 344 531 357
rect 1412 357 1516 363
rect 1524 357 2172 363
rect 2196 357 2268 363
rect 2340 357 2684 363
rect 4260 357 4284 363
rect 4372 357 4588 363
rect 4612 357 4876 363
rect 4900 357 5084 363
rect 116 337 204 343
rect 276 337 428 343
rect 532 337 700 343
rect 1044 337 1308 343
rect 1588 337 2428 343
rect 2468 337 2483 343
rect 84 317 124 323
rect 372 317 380 323
rect 404 317 636 323
rect 772 317 924 323
rect 1188 317 1484 323
rect 1716 317 1996 323
rect 2004 317 2044 323
rect 2164 317 2188 323
rect 2276 317 2348 323
rect 2404 317 2460 323
rect 2477 323 2483 337
rect 2500 337 2620 343
rect 2628 337 2844 343
rect 2852 337 2940 343
rect 2948 337 2988 343
rect 3140 337 3308 343
rect 4180 337 4348 343
rect 4564 337 4652 343
rect 4660 337 5292 343
rect 2477 317 2508 323
rect 2532 317 2572 323
rect 2596 317 2844 323
rect 2868 317 2908 323
rect 3028 317 3228 323
rect 3236 317 3340 323
rect 3540 317 3596 323
rect 4228 317 4476 323
rect 4500 317 5020 323
rect 5092 317 5404 323
rect 5556 317 5596 323
rect 148 297 172 303
rect 196 297 236 303
rect 244 297 284 303
rect 324 297 444 303
rect 500 297 812 303
rect 1012 297 1116 303
rect 1332 297 1356 303
rect 1613 297 1676 303
rect 1613 284 1619 297
rect 1732 297 1836 303
rect 1972 297 1980 303
rect 1988 297 2108 303
rect 2116 297 2188 303
rect 2244 297 2492 303
rect 2500 297 2620 303
rect 2628 297 2732 303
rect 2820 297 2956 303
rect 3124 297 3276 303
rect 3300 297 3356 303
rect 3684 297 3804 303
rect 4132 297 4220 303
rect 4228 297 4252 303
rect 4276 297 4684 303
rect 4708 297 4732 303
rect 4852 297 5116 303
rect 5124 297 5148 303
rect 5156 297 5436 303
rect 5508 297 5628 303
rect 5700 297 5788 303
rect 100 277 252 283
rect 452 277 588 283
rect 900 277 1004 283
rect 1428 277 1612 283
rect 1636 277 1980 283
rect 1988 277 2060 283
rect 2148 277 2204 283
rect 2276 277 2556 283
rect 2564 277 2668 283
rect 2852 277 2860 283
rect 2980 277 3068 283
rect 3076 277 3084 283
rect 3156 277 3196 283
rect 3204 277 3244 283
rect 3444 277 3468 283
rect 3620 277 3740 283
rect 4148 277 4284 283
rect 4292 277 4316 283
rect 4340 277 4380 283
rect 4404 277 4620 283
rect 4644 277 5100 283
rect 5108 277 5500 283
rect 5556 277 5644 283
rect 5796 277 5820 283
rect 20 257 172 263
rect 180 257 284 263
rect 420 257 460 263
rect 580 257 1532 263
rect 1828 257 1964 263
rect 2100 257 2172 263
rect 2196 257 2780 263
rect 3469 263 3475 276
rect 3172 257 3612 263
rect 4084 257 4124 263
rect 4132 257 4508 263
rect 4516 257 4764 263
rect 4772 257 5052 263
rect 5076 257 5084 263
rect 5092 257 5180 263
rect 5620 257 5756 263
rect 660 237 1020 243
rect 1236 237 1292 243
rect 1348 237 2300 243
rect 2308 237 2316 243
rect 2324 237 2652 243
rect 2660 237 2764 243
rect 2877 237 3004 243
rect 1252 217 1420 223
rect 1604 217 1724 223
rect 1796 217 1852 223
rect 1940 217 2172 223
rect 2180 217 2332 223
rect 2340 217 2396 223
rect 2452 217 2540 223
rect 2877 223 2883 237
rect 3060 237 3372 243
rect 3380 237 3420 243
rect 3940 237 4643 243
rect 4637 224 4643 237
rect 4676 237 4780 243
rect 4820 237 4908 243
rect 4980 237 5148 243
rect 5156 237 5260 243
rect 5524 237 5772 243
rect 2660 217 2883 223
rect 3572 217 4108 223
rect 4116 217 4188 223
rect 4196 217 4419 223
rect 2904 214 2952 216
rect 2904 206 2908 214
rect 2918 206 2924 214
rect 2932 206 2938 214
rect 2948 206 2952 214
rect 2904 204 2952 206
rect 4413 204 4419 217
rect 4532 217 4572 223
rect 4644 217 4812 223
rect 4820 217 5011 223
rect 5005 204 5011 217
rect 5060 217 5084 223
rect 5188 217 5196 223
rect 5284 217 5420 223
rect 5428 217 5484 223
rect 5492 217 5660 223
rect 5764 217 5772 223
rect 20 197 44 203
rect 356 197 636 203
rect 772 197 1772 203
rect 1892 197 2028 203
rect 2036 197 2492 203
rect 2500 197 2652 203
rect 3028 197 3100 203
rect 3252 197 3452 203
rect 4100 197 4268 203
rect 4292 197 4332 203
rect 4420 197 4444 203
rect 4564 197 4748 203
rect 4756 197 4828 203
rect 5012 197 5068 203
rect 5140 197 5388 203
rect 5604 197 5692 203
rect 212 177 380 183
rect 964 177 1020 183
rect 1156 177 1404 183
rect 1492 177 1740 183
rect 1748 177 1868 183
rect 1924 177 1980 183
rect 2004 177 2108 183
rect 2164 177 2204 183
rect 2260 177 2444 183
rect 2468 177 2524 183
rect 2548 177 2652 183
rect 2669 177 2876 183
rect 1524 157 1548 163
rect 1604 157 1644 163
rect 1716 157 1948 163
rect 1956 157 2636 163
rect 2669 163 2675 177
rect 2900 177 3100 183
rect 3108 177 3324 183
rect 3332 177 3372 183
rect 4244 177 5228 183
rect 5236 177 5484 183
rect 5652 177 5724 183
rect 5732 177 5820 183
rect 2644 157 2675 163
rect 2692 157 2748 163
rect 2772 157 2972 163
rect 3012 157 3068 163
rect 3092 157 3164 163
rect 3236 157 3276 163
rect 3764 157 4028 163
rect 4036 157 4140 163
rect 4164 157 4332 163
rect 4340 157 4572 163
rect 4596 157 4668 163
rect 4692 157 4924 163
rect 5076 157 5100 163
rect 5124 157 5356 163
rect 5476 157 5708 163
rect 36 137 172 143
rect 1508 137 1612 143
rect 1828 137 2124 143
rect 2324 137 2444 143
rect 2484 137 2492 143
rect 2548 137 2604 143
rect 2612 137 3260 143
rect 3508 137 3692 143
rect 3700 137 3852 143
rect 4020 137 4124 143
rect 4141 143 4147 156
rect 4141 137 4172 143
rect 4228 137 4300 143
rect 4468 137 4524 143
rect 4797 137 4956 143
rect 132 117 268 123
rect 516 117 604 123
rect 708 117 892 123
rect 900 117 988 123
rect 1796 117 1996 123
rect 2004 117 2060 123
rect 2125 123 2131 136
rect 4797 124 4803 137
rect 4964 137 5020 143
rect 5037 137 5155 143
rect 2125 117 2812 123
rect 3060 117 3196 123
rect 3380 117 3820 123
rect 3956 117 4652 123
rect 4660 117 4796 123
rect 4868 117 4940 123
rect 5037 123 5043 137
rect 4996 117 5043 123
rect 5108 117 5116 123
rect 5149 123 5155 137
rect 5172 137 5276 143
rect 5300 137 5340 143
rect 5348 137 5436 143
rect 5460 137 5500 143
rect 5508 137 5548 143
rect 5149 117 5356 123
rect 5364 117 5404 123
rect 5412 117 5468 123
rect 5652 117 5740 123
rect 100 97 156 103
rect 356 97 828 103
rect 1732 97 2780 103
rect 2788 97 3020 103
rect 4132 97 4620 103
rect 4628 97 4684 103
rect 4772 97 5212 103
rect 5220 97 5532 103
rect 5540 97 5564 103
rect 5572 97 5612 103
rect 5780 97 5804 103
rect 5860 97 5891 103
rect 84 77 108 83
rect 244 77 444 83
rect 2020 77 2092 83
rect 2100 77 2252 83
rect 2276 77 2396 83
rect 2436 77 2524 83
rect 2564 77 2652 83
rect 2724 77 3628 83
rect 4260 77 4300 83
rect 2020 57 2332 63
rect 2404 57 3436 63
rect 1352 14 1400 16
rect 1352 6 1356 14
rect 1366 6 1372 14
rect 1380 6 1386 14
rect 1396 6 1400 14
rect 1352 4 1400 6
rect 4440 14 4488 16
rect 4440 6 4444 14
rect 4454 6 4460 14
rect 4468 6 4474 14
rect 4484 6 4488 14
rect 4440 4 4488 6
<< m4contact >>
rect 2908 4206 2910 4214
rect 2910 4206 2916 4214
rect 2924 4206 2932 4214
rect 2940 4206 2946 4214
rect 2946 4206 2948 4214
rect 1948 4196 1956 4204
rect 4764 4196 4772 4204
rect 380 4116 388 4124
rect 2428 4036 2436 4044
rect 4636 4036 4644 4044
rect 2012 4016 2020 4024
rect 1356 4006 1358 4014
rect 1358 4006 1364 4014
rect 1372 4006 1380 4014
rect 1388 4006 1394 4014
rect 1394 4006 1396 4014
rect 4444 4006 4446 4014
rect 4446 4006 4452 4014
rect 4460 4006 4468 4014
rect 4476 4006 4482 4014
rect 4482 4006 4484 4014
rect 4380 3996 4388 4004
rect 4732 3996 4740 4004
rect 2012 3976 2020 3984
rect 1148 3916 1156 3924
rect 2268 3916 2276 3924
rect 2428 3916 2436 3924
rect 4764 3916 4772 3924
rect 1980 3896 1988 3904
rect 1244 3876 1252 3884
rect 1916 3856 1924 3864
rect 2876 3836 2884 3844
rect 5148 3836 5156 3844
rect 636 3796 644 3804
rect 5340 3816 5348 3824
rect 2908 3806 2910 3814
rect 2910 3806 2916 3814
rect 2924 3806 2932 3814
rect 2940 3806 2946 3814
rect 2946 3806 2948 3814
rect 4348 3796 4356 3804
rect 5116 3796 5124 3804
rect 892 3776 900 3784
rect 2428 3776 2436 3784
rect 316 3756 324 3764
rect 2268 3736 2276 3744
rect 636 3716 644 3724
rect 4348 3716 4356 3724
rect 60 3656 68 3664
rect 1916 3656 1924 3664
rect 988 3636 996 3644
rect 4124 3636 4132 3644
rect 5180 3636 5188 3644
rect 1356 3606 1358 3614
rect 1358 3606 1364 3614
rect 1372 3606 1380 3614
rect 1388 3606 1394 3614
rect 1394 3606 1396 3614
rect 4444 3606 4446 3614
rect 4446 3606 4452 3614
rect 4460 3606 4468 3614
rect 4476 3606 4482 3614
rect 4482 3606 4484 3614
rect 2876 3596 2884 3604
rect 4732 3576 4740 3584
rect 2700 3556 2708 3564
rect 4924 3556 4932 3564
rect 1980 3536 1988 3544
rect 2332 3516 2340 3524
rect 2684 3516 2692 3524
rect 60 3496 68 3504
rect 5148 3496 5156 3504
rect 476 3476 484 3484
rect 796 3476 804 3484
rect 380 3456 388 3464
rect 2908 3406 2910 3414
rect 2910 3406 2916 3414
rect 2924 3406 2932 3414
rect 2940 3406 2946 3414
rect 2946 3406 2948 3414
rect 3964 3396 3972 3404
rect 5116 3376 5124 3384
rect 316 3356 324 3364
rect 3868 3356 3876 3364
rect 4380 3336 4388 3344
rect 4604 3336 4612 3344
rect 5372 3336 5380 3344
rect 572 3316 580 3324
rect 1948 3316 1956 3324
rect 5660 3316 5668 3324
rect 604 3296 612 3304
rect 4636 3276 4644 3284
rect 1468 3236 1476 3244
rect 5532 3236 5540 3244
rect 1356 3206 1358 3214
rect 1358 3206 1364 3214
rect 1372 3206 1380 3214
rect 1388 3206 1394 3214
rect 1394 3206 1396 3214
rect 4444 3206 4446 3214
rect 4446 3206 4452 3214
rect 4460 3206 4468 3214
rect 4476 3206 4482 3214
rect 4482 3206 4484 3214
rect 476 3176 484 3184
rect 2332 3176 2340 3184
rect 1276 3156 1284 3164
rect 4124 3156 4132 3164
rect 188 3136 196 3144
rect 4604 3136 4612 3144
rect 924 3116 932 3124
rect 124 3096 132 3104
rect 892 3096 900 3104
rect 604 3076 612 3084
rect 796 3076 804 3084
rect 1532 3076 1540 3084
rect 3868 3076 3876 3084
rect 5340 3056 5348 3064
rect 5820 3036 5828 3044
rect 1564 3016 1572 3024
rect 2908 3006 2910 3014
rect 2910 3006 2916 3014
rect 2924 3006 2932 3014
rect 2940 3006 2946 3014
rect 2946 3006 2948 3014
rect 1084 2996 1092 3004
rect 1180 2996 1188 3004
rect 60 2976 68 2984
rect 476 2976 484 2984
rect 764 2976 772 2984
rect 380 2956 388 2964
rect 540 2956 548 2964
rect 1180 2956 1188 2964
rect 5788 2956 5796 2964
rect 188 2936 196 2944
rect 1084 2936 1092 2944
rect 1212 2936 1220 2944
rect 1244 2936 1252 2944
rect 3868 2936 3876 2944
rect 4924 2936 4932 2944
rect 892 2916 900 2924
rect 1148 2896 1156 2904
rect 1564 2896 1572 2904
rect 3964 2896 3972 2904
rect 1532 2876 1540 2884
rect 1212 2856 1220 2864
rect 924 2836 932 2844
rect 1308 2836 1316 2844
rect 1356 2806 1358 2814
rect 1358 2806 1364 2814
rect 1372 2806 1380 2814
rect 1388 2806 1394 2814
rect 1394 2806 1396 2814
rect 4444 2806 4446 2814
rect 4446 2806 4452 2814
rect 4460 2806 4468 2814
rect 4476 2806 4482 2814
rect 4482 2806 4484 2814
rect 988 2796 996 2804
rect 5628 2776 5636 2784
rect 1308 2736 1316 2744
rect 156 2716 164 2724
rect 1212 2716 1220 2724
rect 1564 2716 1572 2724
rect 4380 2716 4388 2724
rect 4988 2716 4996 2724
rect 604 2696 612 2704
rect 540 2676 548 2684
rect 3036 2656 3044 2664
rect 3068 2656 3076 2664
rect 4380 2616 4388 2624
rect 2908 2606 2910 2614
rect 2910 2606 2916 2614
rect 2924 2606 2932 2614
rect 2940 2606 2946 2614
rect 2946 2606 2948 2614
rect 4636 2596 4644 2604
rect 156 2556 164 2564
rect 892 2556 900 2564
rect 476 2536 484 2544
rect 604 2536 612 2544
rect 3228 2536 3236 2544
rect 5084 2516 5092 2524
rect 3228 2496 3236 2504
rect 1436 2476 1444 2484
rect 1468 2476 1476 2484
rect 4572 2476 4580 2484
rect 1468 2436 1476 2444
rect 1356 2406 1358 2414
rect 1358 2406 1364 2414
rect 1372 2406 1380 2414
rect 1388 2406 1394 2414
rect 1394 2406 1396 2414
rect 4444 2406 4446 2414
rect 4446 2406 4452 2414
rect 4460 2406 4468 2414
rect 4476 2406 4482 2414
rect 4482 2406 4484 2414
rect 1564 2336 1572 2344
rect 764 2276 772 2284
rect 1212 2276 1220 2284
rect 4636 2276 4644 2284
rect 4924 2276 4932 2284
rect 1820 2256 1828 2264
rect 1948 2256 1956 2264
rect 4380 2256 4388 2264
rect 4572 2256 4580 2264
rect 28 2236 36 2244
rect 924 2236 932 2244
rect 2844 2236 2852 2244
rect 892 2216 900 2224
rect 2908 2206 2910 2214
rect 2910 2206 2916 2214
rect 2924 2206 2932 2214
rect 2940 2206 2946 2214
rect 2946 2206 2948 2214
rect 572 2196 580 2204
rect 2844 2176 2852 2184
rect 4572 2136 4580 2144
rect 60 2116 68 2124
rect 1276 2116 1284 2124
rect 4636 2116 4644 2124
rect 5084 2116 5092 2124
rect 1116 2036 1124 2044
rect 1356 2006 1358 2014
rect 1358 2006 1364 2014
rect 1372 2006 1380 2014
rect 1388 2006 1394 2014
rect 1394 2006 1396 2014
rect 4444 2006 4446 2014
rect 4446 2006 4452 2014
rect 4460 2006 4468 2014
rect 4476 2006 4482 2014
rect 4482 2006 4484 2014
rect 348 1936 356 1944
rect 4540 1916 4548 1924
rect 1436 1896 1444 1904
rect 1468 1896 1476 1904
rect 988 1876 996 1884
rect 1500 1836 1508 1844
rect 5660 1836 5668 1844
rect 2908 1806 2910 1814
rect 2910 1806 2916 1814
rect 2924 1806 2932 1814
rect 2940 1806 2946 1814
rect 2946 1806 2948 1814
rect 1820 1796 1828 1804
rect 124 1756 132 1764
rect 3580 1736 3588 1744
rect 4092 1716 4100 1724
rect 1820 1696 1828 1704
rect 3068 1696 3076 1704
rect 4316 1696 4324 1704
rect 5084 1696 5092 1704
rect 5308 1696 5316 1704
rect 5532 1636 5540 1644
rect 2684 1616 2692 1624
rect 1356 1606 1358 1614
rect 1358 1606 1364 1614
rect 1372 1606 1380 1614
rect 1388 1606 1394 1614
rect 1394 1606 1396 1614
rect 4444 1606 4446 1614
rect 4446 1606 4452 1614
rect 4460 1606 4468 1614
rect 4476 1606 4482 1614
rect 4482 1606 4484 1614
rect 124 1536 132 1544
rect 3452 1536 3460 1544
rect 4732 1516 4740 1524
rect 5308 1516 5316 1524
rect 2140 1496 2148 1504
rect 4924 1496 4932 1504
rect 4988 1476 4996 1484
rect 5532 1456 5540 1464
rect 4092 1436 4100 1444
rect 988 1416 996 1424
rect 5500 1416 5508 1424
rect 2908 1406 2910 1414
rect 2910 1406 2916 1414
rect 2924 1406 2932 1414
rect 2940 1406 2946 1414
rect 2946 1406 2948 1414
rect 284 1396 292 1404
rect 2236 1396 2244 1404
rect 3420 1376 3428 1384
rect 700 1356 708 1364
rect 1564 1356 1572 1364
rect 3676 1356 3684 1364
rect 2140 1336 2148 1344
rect 2620 1336 2628 1344
rect 2684 1336 2692 1344
rect 1564 1316 1572 1324
rect 2876 1296 2884 1304
rect 3452 1276 3460 1284
rect 3580 1276 3588 1284
rect 956 1256 964 1264
rect 1116 1256 1124 1264
rect 3068 1256 3076 1264
rect 5404 1236 5412 1244
rect 1020 1216 1028 1224
rect 1356 1206 1358 1214
rect 1358 1206 1364 1214
rect 1372 1206 1380 1214
rect 1388 1206 1394 1214
rect 1394 1206 1396 1214
rect 4444 1206 4446 1214
rect 4446 1206 4452 1214
rect 4460 1206 4468 1214
rect 4476 1206 4482 1214
rect 4482 1206 4484 1214
rect 2748 1196 2756 1204
rect 4316 1196 4324 1204
rect 2236 1176 2244 1184
rect 4540 1176 4548 1184
rect 5084 1176 5092 1184
rect 5788 1176 5796 1184
rect 5276 1156 5284 1164
rect 5372 1156 5380 1164
rect 2620 1136 2628 1144
rect 4764 1136 4772 1144
rect 764 1116 772 1124
rect 892 1116 900 1124
rect 3676 1116 3684 1124
rect 4604 1116 4612 1124
rect 4092 1096 4100 1104
rect 5212 1096 5220 1104
rect 5628 1076 5636 1084
rect 924 1056 932 1064
rect 4092 1056 4100 1064
rect 1020 1036 1028 1044
rect 2876 1016 2884 1024
rect 2908 1006 2910 1014
rect 2910 1006 2916 1014
rect 2924 1006 2932 1014
rect 2940 1006 2946 1014
rect 2946 1006 2948 1014
rect 28 996 36 1004
rect 4796 996 4804 1004
rect 1020 976 1028 984
rect 1052 976 1060 984
rect 2172 976 2180 984
rect 2748 976 2756 984
rect 4636 976 4644 984
rect 4764 976 4772 984
rect 572 956 580 964
rect 2780 956 2788 964
rect 3292 956 3300 964
rect 4732 956 4740 964
rect 636 936 644 944
rect 700 936 708 944
rect 1436 936 1444 944
rect 2972 936 2980 944
rect 124 916 132 924
rect 1052 916 1060 924
rect 3036 916 3044 924
rect 3420 916 3428 924
rect 4604 916 4612 924
rect 508 896 516 904
rect 380 876 388 884
rect 1436 896 1444 904
rect 1468 896 1476 904
rect 1020 816 1028 824
rect 1356 806 1358 814
rect 1358 806 1364 814
rect 1372 806 1380 814
rect 1388 806 1394 814
rect 1394 806 1396 814
rect 4444 806 4446 814
rect 4446 806 4452 814
rect 4460 806 4468 814
rect 4476 806 4482 814
rect 4482 806 4484 814
rect 348 796 356 804
rect 4636 736 4644 744
rect 764 716 772 724
rect 4796 716 4804 724
rect 4956 716 4964 724
rect 3068 696 3076 704
rect 4604 696 4612 704
rect 4988 696 4996 704
rect 956 676 964 684
rect 988 676 996 684
rect 1020 676 1028 684
rect 2812 676 2820 684
rect 5084 676 5092 684
rect 2620 656 2628 664
rect 1500 636 1508 644
rect 1724 636 1732 644
rect 2812 636 2820 644
rect 3004 636 3012 644
rect 4348 656 4356 664
rect 4988 656 4996 664
rect 3292 636 3300 644
rect 5404 636 5412 644
rect 2908 606 2910 614
rect 2910 606 2916 614
rect 2924 606 2932 614
rect 2940 606 2946 614
rect 2946 606 2948 614
rect 1468 596 1476 604
rect 2780 596 2788 604
rect 3004 596 3012 604
rect 2812 576 2820 584
rect 284 556 292 564
rect 2172 556 2180 564
rect 2812 536 2820 544
rect 3004 536 3012 544
rect 3036 536 3044 544
rect 4348 536 4356 544
rect 5084 536 5092 544
rect 4380 516 4388 524
rect 5212 516 5220 524
rect 5756 516 5764 524
rect 508 496 516 504
rect 988 496 996 504
rect 2972 496 2980 504
rect 4956 496 4964 504
rect 5276 496 5284 504
rect 5500 496 5508 504
rect 4508 456 4516 464
rect 5532 436 5540 444
rect 1356 406 1358 414
rect 1358 406 1364 414
rect 1372 406 1380 414
rect 1388 406 1394 414
rect 1394 406 1396 414
rect 4444 406 4446 414
rect 4446 406 4452 414
rect 4460 406 4468 414
rect 4476 406 4482 414
rect 4482 406 4484 414
rect 4252 376 4260 384
rect 4604 376 4612 384
rect 4732 376 4740 384
rect 2268 356 2276 364
rect 4284 356 4292 364
rect 4588 356 4596 364
rect 2460 336 2468 344
rect 380 316 388 324
rect 2396 316 2404 324
rect 2492 336 2500 344
rect 4348 336 4356 344
rect 2524 316 2532 324
rect 2844 316 2852 324
rect 284 296 292 304
rect 1980 296 1988 304
rect 2236 296 2244 304
rect 4732 296 4740 304
rect 5116 296 5124 304
rect 5692 296 5700 304
rect 2268 276 2276 284
rect 2844 276 2852 284
rect 3068 276 3076 284
rect 5820 276 5828 284
rect 4508 256 4516 264
rect 5084 256 5092 264
rect 2652 216 2660 224
rect 2908 206 2910 214
rect 2910 206 2916 214
rect 2924 206 2932 214
rect 2940 206 2946 214
rect 2946 206 2948 214
rect 5084 216 5092 224
rect 5180 216 5188 224
rect 5756 216 5764 224
rect 636 196 644 204
rect 4284 196 4292 204
rect 4348 196 4356 204
rect 4380 196 4388 204
rect 5692 196 5700 204
rect 1020 176 1028 184
rect 1980 176 1988 184
rect 2524 176 2532 184
rect 2652 176 2660 184
rect 2684 156 2692 164
rect 2236 136 2244 144
rect 2460 136 2468 144
rect 2492 136 2500 144
rect 636 116 644 124
rect 5116 116 5124 124
rect 1724 96 1732 104
rect 2396 76 2404 84
rect 2652 76 2660 84
rect 4252 76 4260 84
rect 1356 6 1358 14
rect 1358 6 1364 14
rect 1372 6 1380 14
rect 1388 6 1394 14
rect 1394 6 1396 14
rect 4444 6 4446 14
rect 4446 6 4452 14
rect 4460 6 4468 14
rect 4476 6 4482 14
rect 4482 6 4484 14
<< metal4 >>
rect 378 4124 390 4126
rect 378 4116 380 4124
rect 388 4116 390 4124
rect 314 3764 326 3766
rect 314 3756 316 3764
rect 324 3756 326 3764
rect 58 3664 70 3666
rect 58 3656 60 3664
rect 68 3656 70 3664
rect 58 3504 70 3656
rect 58 3496 60 3504
rect 68 3496 70 3504
rect 58 3494 70 3496
rect 314 3364 326 3756
rect 314 3356 316 3364
rect 324 3356 326 3364
rect 314 3354 326 3356
rect 378 3464 390 4116
rect 1352 4014 1400 4240
rect 2904 4214 2952 4240
rect 2904 4206 2908 4214
rect 2916 4206 2924 4214
rect 2932 4206 2940 4214
rect 2948 4206 2952 4214
rect 1352 4006 1356 4014
rect 1364 4006 1372 4014
rect 1380 4006 1388 4014
rect 1396 4006 1400 4014
rect 1146 3924 1158 3926
rect 1146 3916 1148 3924
rect 1156 3916 1158 3924
rect 634 3804 646 3806
rect 634 3796 636 3804
rect 644 3796 646 3804
rect 634 3724 646 3796
rect 634 3716 636 3724
rect 644 3716 646 3724
rect 634 3714 646 3716
rect 890 3784 902 3786
rect 890 3776 892 3784
rect 900 3776 902 3784
rect 378 3456 380 3464
rect 388 3456 390 3464
rect 186 3144 198 3146
rect 186 3136 188 3144
rect 196 3136 198 3144
rect 122 3104 134 3106
rect 122 3096 124 3104
rect 132 3096 134 3104
rect 58 2984 70 2986
rect 58 2976 60 2984
rect 68 2976 70 2984
rect 26 2244 38 2246
rect 26 2236 28 2244
rect 36 2236 38 2244
rect 26 1004 38 2236
rect 58 2124 70 2976
rect 58 2116 60 2124
rect 68 2116 70 2124
rect 58 2114 70 2116
rect 122 1764 134 3096
rect 186 2944 198 3136
rect 378 2964 390 3456
rect 474 3484 486 3486
rect 474 3476 476 3484
rect 484 3476 486 3484
rect 474 3184 486 3476
rect 794 3484 806 3486
rect 794 3476 796 3484
rect 804 3476 806 3484
rect 474 3176 476 3184
rect 484 3176 486 3184
rect 474 3174 486 3176
rect 570 3324 582 3326
rect 570 3316 572 3324
rect 580 3316 582 3324
rect 378 2956 380 2964
rect 388 2956 390 2964
rect 378 2954 390 2956
rect 474 2984 486 2986
rect 474 2976 476 2984
rect 484 2976 486 2984
rect 186 2936 188 2944
rect 196 2936 198 2944
rect 186 2934 198 2936
rect 154 2724 166 2726
rect 154 2716 156 2724
rect 164 2716 166 2724
rect 154 2564 166 2716
rect 154 2556 156 2564
rect 164 2556 166 2564
rect 154 2554 166 2556
rect 474 2544 486 2976
rect 538 2964 550 2966
rect 538 2956 540 2964
rect 548 2956 550 2964
rect 538 2684 550 2956
rect 538 2676 540 2684
rect 548 2676 550 2684
rect 538 2674 550 2676
rect 474 2536 476 2544
rect 484 2536 486 2544
rect 474 2534 486 2536
rect 570 2204 582 3316
rect 602 3304 614 3306
rect 602 3296 604 3304
rect 612 3296 614 3304
rect 602 3084 614 3296
rect 602 3076 604 3084
rect 612 3076 614 3084
rect 602 3074 614 3076
rect 794 3084 806 3476
rect 890 3104 902 3776
rect 986 3644 998 3646
rect 986 3636 988 3644
rect 996 3636 998 3644
rect 890 3096 892 3104
rect 900 3096 902 3104
rect 890 3094 902 3096
rect 922 3124 934 3126
rect 922 3116 924 3124
rect 932 3116 934 3124
rect 794 3076 796 3084
rect 804 3076 806 3084
rect 794 3074 806 3076
rect 762 2984 774 2986
rect 762 2976 764 2984
rect 772 2976 774 2984
rect 602 2704 614 2706
rect 602 2696 604 2704
rect 612 2696 614 2704
rect 602 2544 614 2696
rect 602 2536 604 2544
rect 612 2536 614 2544
rect 602 2534 614 2536
rect 762 2284 774 2976
rect 890 2924 902 2926
rect 890 2916 892 2924
rect 900 2916 902 2924
rect 890 2564 902 2916
rect 922 2844 934 3116
rect 922 2836 924 2844
rect 932 2836 934 2844
rect 922 2834 934 2836
rect 986 2804 998 3636
rect 1082 3004 1094 3006
rect 1082 2996 1084 3004
rect 1092 2996 1094 3004
rect 1082 2944 1094 2996
rect 1082 2936 1084 2944
rect 1092 2936 1094 2944
rect 1082 2934 1094 2936
rect 1146 2904 1158 3916
rect 1242 3884 1254 3886
rect 1242 3876 1244 3884
rect 1252 3876 1254 3884
rect 1178 3004 1190 3006
rect 1178 2996 1180 3004
rect 1188 2996 1190 3004
rect 1178 2964 1190 2996
rect 1178 2956 1180 2964
rect 1188 2956 1190 2964
rect 1178 2954 1190 2956
rect 1146 2896 1148 2904
rect 1156 2896 1158 2904
rect 1146 2894 1158 2896
rect 1210 2944 1222 2946
rect 1210 2936 1212 2944
rect 1220 2936 1222 2944
rect 1210 2864 1222 2936
rect 1242 2944 1254 3876
rect 1352 3614 1400 4006
rect 1946 4204 1958 4206
rect 1946 4196 1948 4204
rect 1956 4196 1958 4204
rect 1914 3864 1926 3866
rect 1914 3856 1916 3864
rect 1924 3856 1926 3864
rect 1914 3664 1926 3856
rect 1914 3656 1916 3664
rect 1924 3656 1926 3664
rect 1914 3654 1926 3656
rect 1352 3606 1356 3614
rect 1364 3606 1372 3614
rect 1380 3606 1388 3614
rect 1396 3606 1400 3614
rect 1352 3214 1400 3606
rect 1946 3324 1958 4196
rect 2426 4044 2438 4046
rect 2426 4036 2428 4044
rect 2436 4036 2438 4044
rect 2010 4024 2022 4026
rect 2010 4016 2012 4024
rect 2020 4016 2022 4024
rect 2010 3984 2022 4016
rect 2010 3976 2012 3984
rect 2020 3976 2022 3984
rect 2010 3974 2022 3976
rect 2266 3924 2278 3926
rect 2266 3916 2268 3924
rect 2276 3916 2278 3924
rect 1978 3904 1990 3906
rect 1978 3896 1980 3904
rect 1988 3896 1990 3904
rect 1978 3544 1990 3896
rect 2266 3744 2278 3916
rect 2426 3924 2438 4036
rect 2426 3916 2428 3924
rect 2436 3916 2438 3924
rect 2426 3784 2438 3916
rect 2426 3776 2428 3784
rect 2436 3776 2438 3784
rect 2426 3774 2438 3776
rect 2874 3844 2886 3846
rect 2874 3836 2876 3844
rect 2884 3836 2886 3844
rect 2266 3736 2268 3744
rect 2276 3736 2278 3744
rect 2266 3734 2278 3736
rect 2874 3604 2886 3836
rect 2874 3596 2876 3604
rect 2884 3596 2886 3604
rect 2874 3594 2886 3596
rect 2904 3814 2952 4206
rect 4440 4014 4488 4240
rect 4762 4204 4774 4206
rect 4762 4196 4764 4204
rect 4772 4196 4774 4204
rect 4440 4006 4444 4014
rect 4452 4006 4460 4014
rect 4468 4006 4476 4014
rect 4484 4006 4488 4014
rect 2904 3806 2908 3814
rect 2916 3806 2924 3814
rect 2932 3806 2940 3814
rect 2948 3806 2952 3814
rect 4378 4004 4390 4006
rect 4378 3996 4380 4004
rect 4388 3996 4390 4004
rect 1978 3536 1980 3544
rect 1988 3536 1990 3544
rect 1978 3534 1990 3536
rect 2682 3564 2710 3566
rect 2682 3556 2700 3564
rect 2708 3556 2710 3564
rect 2682 3554 2710 3556
rect 1946 3316 1948 3324
rect 1956 3316 1958 3324
rect 1352 3206 1356 3214
rect 1364 3206 1372 3214
rect 1380 3206 1388 3214
rect 1396 3206 1400 3214
rect 1242 2936 1244 2944
rect 1252 2936 1254 2944
rect 1242 2934 1254 2936
rect 1274 3164 1286 3166
rect 1274 3156 1276 3164
rect 1284 3156 1286 3164
rect 1210 2856 1212 2864
rect 1220 2856 1222 2864
rect 1210 2854 1222 2856
rect 986 2796 988 2804
rect 996 2796 998 2804
rect 986 2794 998 2796
rect 890 2556 892 2564
rect 900 2556 902 2564
rect 890 2554 902 2556
rect 1210 2724 1222 2726
rect 1210 2716 1212 2724
rect 1220 2716 1222 2724
rect 762 2276 764 2284
rect 772 2276 774 2284
rect 762 2274 774 2276
rect 1210 2284 1222 2716
rect 1210 2276 1212 2284
rect 1220 2276 1222 2284
rect 1210 2274 1222 2276
rect 922 2244 934 2246
rect 922 2236 924 2244
rect 932 2236 934 2244
rect 570 2196 572 2204
rect 580 2196 582 2204
rect 570 2194 582 2196
rect 890 2224 902 2226
rect 890 2216 892 2224
rect 900 2216 902 2224
rect 122 1756 124 1764
rect 132 1756 134 1764
rect 122 1754 134 1756
rect 346 1944 358 1946
rect 346 1936 348 1944
rect 356 1936 358 1944
rect 26 996 28 1004
rect 36 996 38 1004
rect 26 994 38 996
rect 122 1544 134 1546
rect 122 1536 124 1544
rect 132 1536 134 1544
rect 122 924 134 1536
rect 122 916 124 924
rect 132 916 134 924
rect 122 914 134 916
rect 282 1404 294 1406
rect 282 1396 284 1404
rect 292 1396 294 1404
rect 282 564 294 1396
rect 346 804 358 1936
rect 698 1364 710 1366
rect 698 1356 700 1364
rect 708 1356 710 1364
rect 570 964 646 966
rect 570 956 572 964
rect 580 956 646 964
rect 570 954 646 956
rect 634 944 646 954
rect 634 936 636 944
rect 644 936 646 944
rect 634 934 646 936
rect 698 944 710 1356
rect 698 936 700 944
rect 708 936 710 944
rect 698 934 710 936
rect 762 1124 774 1126
rect 762 1116 764 1124
rect 772 1116 774 1124
rect 506 904 518 906
rect 506 896 508 904
rect 516 896 518 904
rect 346 796 348 804
rect 356 796 358 804
rect 346 794 358 796
rect 378 884 390 886
rect 378 876 380 884
rect 388 876 390 884
rect 282 556 284 564
rect 292 556 294 564
rect 282 304 294 556
rect 378 324 390 876
rect 506 504 518 896
rect 762 724 774 1116
rect 890 1124 902 2216
rect 890 1116 892 1124
rect 900 1116 902 1124
rect 890 1114 902 1116
rect 922 1064 934 2236
rect 1274 2124 1286 3156
rect 1306 2844 1318 2846
rect 1306 2836 1308 2844
rect 1316 2836 1318 2844
rect 1306 2744 1318 2836
rect 1306 2736 1308 2744
rect 1316 2736 1318 2744
rect 1306 2734 1318 2736
rect 1352 2814 1400 3206
rect 1352 2806 1356 2814
rect 1364 2806 1372 2814
rect 1380 2806 1388 2814
rect 1396 2806 1400 2814
rect 1274 2116 1276 2124
rect 1284 2116 1286 2124
rect 1274 2114 1286 2116
rect 1352 2414 1400 2806
rect 1466 3244 1478 3246
rect 1466 3236 1468 3244
rect 1476 3236 1478 3244
rect 1352 2406 1356 2414
rect 1364 2406 1372 2414
rect 1380 2406 1388 2414
rect 1396 2406 1400 2414
rect 1114 2044 1126 2046
rect 1114 2036 1116 2044
rect 1124 2036 1126 2044
rect 986 1884 998 1886
rect 986 1876 988 1884
rect 996 1876 998 1884
rect 986 1424 998 1876
rect 986 1416 988 1424
rect 996 1416 998 1424
rect 986 1414 998 1416
rect 922 1056 924 1064
rect 932 1056 934 1064
rect 922 1054 934 1056
rect 954 1264 966 1266
rect 954 1256 956 1264
rect 964 1256 966 1264
rect 762 716 764 724
rect 772 716 774 724
rect 762 714 774 716
rect 954 684 966 1256
rect 1114 1264 1126 2036
rect 1114 1256 1116 1264
rect 1124 1256 1126 1264
rect 1114 1254 1126 1256
rect 1352 2014 1400 2406
rect 1352 2006 1356 2014
rect 1364 2006 1372 2014
rect 1380 2006 1388 2014
rect 1396 2006 1400 2014
rect 1352 1614 1400 2006
rect 1434 2484 1446 2486
rect 1434 2476 1436 2484
rect 1444 2476 1446 2484
rect 1434 1904 1446 2476
rect 1466 2484 1478 3236
rect 1530 3084 1542 3086
rect 1530 3076 1532 3084
rect 1540 3076 1542 3084
rect 1530 2884 1542 3076
rect 1562 3024 1574 3026
rect 1562 3016 1564 3024
rect 1572 3016 1574 3024
rect 1562 2904 1574 3016
rect 1562 2896 1564 2904
rect 1572 2896 1574 2904
rect 1562 2894 1574 2896
rect 1530 2876 1532 2884
rect 1540 2876 1542 2884
rect 1530 2874 1542 2876
rect 1466 2476 1468 2484
rect 1476 2476 1478 2484
rect 1466 2474 1478 2476
rect 1562 2724 1574 2726
rect 1562 2716 1564 2724
rect 1572 2716 1574 2724
rect 1434 1896 1436 1904
rect 1444 1896 1446 1904
rect 1434 1894 1446 1896
rect 1466 2444 1478 2446
rect 1466 2436 1468 2444
rect 1476 2436 1478 2444
rect 1466 1904 1478 2436
rect 1562 2344 1574 2716
rect 1562 2336 1564 2344
rect 1572 2336 1574 2344
rect 1562 2334 1574 2336
rect 1466 1896 1468 1904
rect 1476 1896 1478 1904
rect 1466 1894 1478 1896
rect 1818 2264 1830 2266
rect 1818 2256 1820 2264
rect 1828 2256 1830 2264
rect 1352 1606 1356 1614
rect 1364 1606 1372 1614
rect 1380 1606 1388 1614
rect 1396 1606 1400 1614
rect 1018 1224 1030 1226
rect 1018 1216 1020 1224
rect 1028 1216 1030 1224
rect 1018 1044 1030 1216
rect 1018 1036 1020 1044
rect 1028 1036 1030 1044
rect 1018 1034 1030 1036
rect 1352 1214 1400 1606
rect 1352 1206 1356 1214
rect 1364 1206 1372 1214
rect 1380 1206 1388 1214
rect 1396 1206 1400 1214
rect 1018 984 1030 986
rect 1018 976 1020 984
rect 1028 976 1030 984
rect 1018 824 1030 976
rect 1050 984 1062 986
rect 1050 976 1052 984
rect 1060 976 1062 984
rect 1050 924 1062 976
rect 1050 916 1052 924
rect 1060 916 1062 924
rect 1050 914 1062 916
rect 1018 816 1020 824
rect 1028 816 1030 824
rect 1018 814 1030 816
rect 1352 814 1400 1206
rect 1498 1844 1510 1846
rect 1498 1836 1500 1844
rect 1508 1836 1510 1844
rect 1434 944 1446 946
rect 1434 936 1436 944
rect 1444 936 1446 944
rect 1434 904 1446 936
rect 1434 896 1436 904
rect 1444 896 1446 904
rect 1434 894 1446 896
rect 1466 904 1478 906
rect 1466 896 1468 904
rect 1476 896 1478 904
rect 1352 806 1356 814
rect 1364 806 1372 814
rect 1380 806 1388 814
rect 1396 806 1400 814
rect 954 676 956 684
rect 964 676 966 684
rect 954 674 966 676
rect 986 684 998 686
rect 986 676 988 684
rect 996 676 998 684
rect 506 496 508 504
rect 516 496 518 504
rect 506 494 518 496
rect 986 504 998 676
rect 986 496 988 504
rect 996 496 998 504
rect 986 494 998 496
rect 1018 684 1030 686
rect 1018 676 1020 684
rect 1028 676 1030 684
rect 378 316 380 324
rect 388 316 390 324
rect 378 314 390 316
rect 282 296 284 304
rect 292 296 294 304
rect 282 294 294 296
rect 634 204 646 206
rect 634 196 636 204
rect 644 196 646 204
rect 634 124 646 196
rect 1018 184 1030 676
rect 1018 176 1020 184
rect 1028 176 1030 184
rect 1018 174 1030 176
rect 1352 414 1400 806
rect 1466 604 1478 896
rect 1498 644 1510 1836
rect 1818 1804 1830 2256
rect 1946 2264 1958 3316
rect 2330 3524 2342 3526
rect 2330 3516 2332 3524
rect 2340 3516 2342 3524
rect 2330 3184 2342 3516
rect 2682 3524 2694 3554
rect 2682 3516 2684 3524
rect 2692 3516 2694 3524
rect 2682 3514 2694 3516
rect 2330 3176 2332 3184
rect 2340 3176 2342 3184
rect 2330 3174 2342 3176
rect 2904 3414 2952 3806
rect 4346 3804 4358 3806
rect 4346 3796 4348 3804
rect 4356 3796 4358 3804
rect 4346 3724 4358 3796
rect 4346 3716 4348 3724
rect 4356 3716 4358 3724
rect 4346 3714 4358 3716
rect 2904 3406 2908 3414
rect 2916 3406 2924 3414
rect 2932 3406 2940 3414
rect 2948 3406 2952 3414
rect 4122 3644 4134 3646
rect 4122 3636 4124 3644
rect 4132 3636 4134 3644
rect 1946 2256 1948 2264
rect 1956 2256 1958 2264
rect 1946 2254 1958 2256
rect 2904 3014 2952 3406
rect 3962 3404 3974 3406
rect 3962 3396 3964 3404
rect 3972 3396 3974 3404
rect 2904 3006 2908 3014
rect 2916 3006 2924 3014
rect 2932 3006 2940 3014
rect 2948 3006 2952 3014
rect 2904 2614 2952 3006
rect 3866 3364 3878 3366
rect 3866 3356 3868 3364
rect 3876 3356 3878 3364
rect 3866 3084 3878 3356
rect 3866 3076 3868 3084
rect 3876 3076 3878 3084
rect 3866 2944 3878 3076
rect 3866 2936 3868 2944
rect 3876 2936 3878 2944
rect 3866 2934 3878 2936
rect 3962 2904 3974 3396
rect 4122 3164 4134 3636
rect 4378 3344 4390 3996
rect 4378 3336 4380 3344
rect 4388 3336 4390 3344
rect 4378 3334 4390 3336
rect 4440 3614 4488 4006
rect 4440 3606 4444 3614
rect 4452 3606 4460 3614
rect 4468 3606 4476 3614
rect 4484 3606 4488 3614
rect 4122 3156 4124 3164
rect 4132 3156 4134 3164
rect 4122 3154 4134 3156
rect 4440 3214 4488 3606
rect 4634 4044 4646 4046
rect 4634 4036 4636 4044
rect 4644 4036 4646 4044
rect 4440 3206 4444 3214
rect 4452 3206 4460 3214
rect 4468 3206 4476 3214
rect 4484 3206 4488 3214
rect 3962 2896 3964 2904
rect 3972 2896 3974 2904
rect 3962 2894 3974 2896
rect 4440 2814 4488 3206
rect 4602 3344 4614 3346
rect 4602 3336 4604 3344
rect 4612 3336 4614 3344
rect 4602 3144 4614 3336
rect 4634 3284 4646 4036
rect 4730 4004 4742 4006
rect 4730 3996 4732 4004
rect 4740 3996 4742 4004
rect 4730 3584 4742 3996
rect 4762 3924 4774 4196
rect 4762 3916 4764 3924
rect 4772 3916 4774 3924
rect 4762 3914 4774 3916
rect 5146 3844 5158 3846
rect 5146 3836 5148 3844
rect 5156 3836 5158 3844
rect 4730 3576 4732 3584
rect 4740 3576 4742 3584
rect 4730 3574 4742 3576
rect 5114 3804 5126 3806
rect 5114 3796 5116 3804
rect 5124 3796 5126 3804
rect 4634 3276 4636 3284
rect 4644 3276 4646 3284
rect 4634 3274 4646 3276
rect 4922 3564 4934 3566
rect 4922 3556 4924 3564
rect 4932 3556 4934 3564
rect 4602 3136 4604 3144
rect 4612 3136 4614 3144
rect 4602 3134 4614 3136
rect 4922 2944 4934 3556
rect 5114 3384 5126 3796
rect 5146 3504 5158 3836
rect 5338 3824 5350 3826
rect 5338 3816 5340 3824
rect 5348 3816 5350 3824
rect 5146 3496 5148 3504
rect 5156 3496 5158 3504
rect 5146 3494 5158 3496
rect 5178 3644 5190 3646
rect 5178 3636 5180 3644
rect 5188 3636 5190 3644
rect 5114 3376 5116 3384
rect 5124 3376 5126 3384
rect 5114 3374 5126 3376
rect 4922 2936 4924 2944
rect 4932 2936 4934 2944
rect 4922 2934 4934 2936
rect 4440 2806 4444 2814
rect 4452 2806 4460 2814
rect 4468 2806 4476 2814
rect 4484 2806 4488 2814
rect 4378 2724 4390 2726
rect 4378 2716 4380 2724
rect 4388 2716 4390 2724
rect 3034 2674 3078 2686
rect 3034 2664 3046 2674
rect 3034 2656 3036 2664
rect 3044 2656 3046 2664
rect 3034 2654 3046 2656
rect 3066 2664 3078 2674
rect 3066 2656 3068 2664
rect 3076 2656 3078 2664
rect 3066 2654 3078 2656
rect 2904 2606 2908 2614
rect 2916 2606 2924 2614
rect 2932 2606 2940 2614
rect 2948 2606 2952 2614
rect 2842 2244 2854 2246
rect 2842 2236 2844 2244
rect 2852 2236 2854 2244
rect 2842 2184 2854 2236
rect 2842 2176 2844 2184
rect 2852 2176 2854 2184
rect 2842 2174 2854 2176
rect 2904 2214 2952 2606
rect 4378 2624 4390 2716
rect 4378 2616 4380 2624
rect 4388 2616 4390 2624
rect 3226 2544 3238 2546
rect 3226 2536 3228 2544
rect 3236 2536 3238 2544
rect 3226 2504 3238 2536
rect 3226 2496 3228 2504
rect 3236 2496 3238 2504
rect 3226 2494 3238 2496
rect 4378 2264 4390 2616
rect 4378 2256 4380 2264
rect 4388 2256 4390 2264
rect 4378 2254 4390 2256
rect 4440 2414 4488 2806
rect 4986 2724 4998 2726
rect 4986 2716 4988 2724
rect 4996 2716 4998 2724
rect 4634 2604 4646 2606
rect 4634 2596 4636 2604
rect 4644 2596 4646 2604
rect 4440 2406 4444 2414
rect 4452 2406 4460 2414
rect 4468 2406 4476 2414
rect 4484 2406 4488 2414
rect 2904 2206 2908 2214
rect 2916 2206 2924 2214
rect 2932 2206 2940 2214
rect 2948 2206 2952 2214
rect 1818 1796 1820 1804
rect 1828 1796 1830 1804
rect 1818 1704 1830 1796
rect 1818 1696 1820 1704
rect 1828 1696 1830 1704
rect 1818 1694 1830 1696
rect 2904 1814 2952 2206
rect 2904 1806 2908 1814
rect 2916 1806 2924 1814
rect 2932 1806 2940 1814
rect 2948 1806 2952 1814
rect 2682 1624 2694 1626
rect 2682 1616 2684 1624
rect 2692 1616 2694 1624
rect 2138 1504 2150 1506
rect 2138 1496 2140 1504
rect 2148 1496 2150 1504
rect 1562 1364 1574 1366
rect 1562 1356 1564 1364
rect 1572 1356 1574 1364
rect 1562 1324 1574 1356
rect 2138 1344 2150 1496
rect 2138 1336 2140 1344
rect 2148 1336 2150 1344
rect 2138 1334 2150 1336
rect 2234 1404 2246 1406
rect 2234 1396 2236 1404
rect 2244 1396 2246 1404
rect 1562 1316 1564 1324
rect 1572 1316 1574 1324
rect 1562 1314 1574 1316
rect 2234 1184 2246 1396
rect 2234 1176 2236 1184
rect 2244 1176 2246 1184
rect 2234 1174 2246 1176
rect 2618 1344 2630 1346
rect 2618 1336 2620 1344
rect 2628 1336 2630 1344
rect 2618 1144 2630 1336
rect 2682 1344 2694 1616
rect 2682 1336 2684 1344
rect 2692 1336 2694 1344
rect 2682 1334 2694 1336
rect 2904 1414 2952 1806
rect 4440 2014 4488 2406
rect 4570 2484 4582 2486
rect 4570 2476 4572 2484
rect 4580 2476 4582 2484
rect 4570 2264 4582 2476
rect 4570 2256 4572 2264
rect 4580 2256 4582 2264
rect 4570 2144 4582 2256
rect 4570 2136 4572 2144
rect 4580 2136 4582 2144
rect 4570 2134 4582 2136
rect 4634 2284 4646 2596
rect 4634 2276 4636 2284
rect 4644 2276 4646 2284
rect 4634 2124 4646 2276
rect 4634 2116 4636 2124
rect 4644 2116 4646 2124
rect 4634 2114 4646 2116
rect 4922 2284 4934 2286
rect 4922 2276 4924 2284
rect 4932 2276 4934 2284
rect 4440 2006 4444 2014
rect 4452 2006 4460 2014
rect 4468 2006 4476 2014
rect 4484 2006 4488 2014
rect 3578 1744 3590 1746
rect 3578 1736 3580 1744
rect 3588 1736 3590 1744
rect 2904 1406 2908 1414
rect 2916 1406 2924 1414
rect 2932 1406 2940 1414
rect 2948 1406 2952 1414
rect 2874 1304 2886 1306
rect 2874 1296 2876 1304
rect 2884 1296 2886 1304
rect 2618 1136 2620 1144
rect 2628 1136 2630 1144
rect 2170 984 2182 986
rect 2170 976 2172 984
rect 2180 976 2182 984
rect 1498 636 1500 644
rect 1508 636 1510 644
rect 1498 634 1510 636
rect 1722 644 1734 646
rect 1722 636 1724 644
rect 1732 636 1734 644
rect 1466 596 1468 604
rect 1476 596 1478 604
rect 1466 594 1478 596
rect 1352 406 1356 414
rect 1364 406 1372 414
rect 1380 406 1388 414
rect 1396 406 1400 414
rect 634 116 636 124
rect 644 116 646 124
rect 634 114 646 116
rect 1352 14 1400 406
rect 1722 104 1734 636
rect 2170 564 2182 976
rect 2618 664 2630 1136
rect 2746 1204 2758 1206
rect 2746 1196 2748 1204
rect 2756 1196 2758 1204
rect 2746 984 2758 1196
rect 2874 1024 2886 1296
rect 2874 1016 2876 1024
rect 2884 1016 2886 1024
rect 2874 1014 2886 1016
rect 2904 1014 2952 1406
rect 3066 1704 3078 1706
rect 3066 1696 3068 1704
rect 3076 1696 3078 1704
rect 3066 1264 3078 1696
rect 3450 1544 3462 1546
rect 3450 1536 3452 1544
rect 3460 1536 3462 1544
rect 3066 1256 3068 1264
rect 3076 1256 3078 1264
rect 3066 1254 3078 1256
rect 3418 1384 3430 1386
rect 3418 1376 3420 1384
rect 3428 1376 3430 1384
rect 2746 976 2748 984
rect 2756 976 2758 984
rect 2746 974 2758 976
rect 2904 1006 2908 1014
rect 2916 1006 2924 1014
rect 2932 1006 2940 1014
rect 2948 1006 2952 1014
rect 2618 656 2620 664
rect 2628 656 2630 664
rect 2618 654 2630 656
rect 2778 964 2790 966
rect 2778 956 2780 964
rect 2788 956 2790 964
rect 2778 604 2790 956
rect 2810 684 2822 686
rect 2810 676 2812 684
rect 2820 676 2822 684
rect 2810 644 2822 676
rect 2810 636 2812 644
rect 2820 636 2822 644
rect 2810 634 2822 636
rect 2778 596 2780 604
rect 2788 596 2790 604
rect 2778 594 2790 596
rect 2904 614 2952 1006
rect 3290 964 3302 966
rect 3290 956 3292 964
rect 3300 956 3302 964
rect 2904 606 2908 614
rect 2916 606 2924 614
rect 2932 606 2940 614
rect 2948 606 2952 614
rect 2170 556 2172 564
rect 2180 556 2182 564
rect 2170 554 2182 556
rect 2810 584 2822 586
rect 2810 576 2812 584
rect 2820 576 2822 584
rect 2810 544 2822 576
rect 2810 536 2812 544
rect 2820 536 2822 544
rect 2810 534 2822 536
rect 2266 364 2278 366
rect 2266 356 2268 364
rect 2276 356 2278 364
rect 1978 304 1990 306
rect 1978 296 1980 304
rect 1988 296 1990 304
rect 1978 184 1990 296
rect 1978 176 1980 184
rect 1988 176 1990 184
rect 1978 174 1990 176
rect 2234 304 2246 306
rect 2234 296 2236 304
rect 2244 296 2246 304
rect 2234 144 2246 296
rect 2266 284 2278 356
rect 2458 344 2470 346
rect 2458 336 2460 344
rect 2468 336 2470 344
rect 2266 276 2268 284
rect 2276 276 2278 284
rect 2266 274 2278 276
rect 2394 324 2406 326
rect 2394 316 2396 324
rect 2404 316 2406 324
rect 2234 136 2236 144
rect 2244 136 2246 144
rect 2234 134 2246 136
rect 1722 96 1724 104
rect 1732 96 1734 104
rect 1722 94 1734 96
rect 2394 84 2406 316
rect 2458 144 2470 336
rect 2458 136 2460 144
rect 2468 136 2470 144
rect 2458 134 2470 136
rect 2490 344 2502 346
rect 2490 336 2492 344
rect 2500 336 2502 344
rect 2490 144 2502 336
rect 2522 324 2534 326
rect 2522 316 2524 324
rect 2532 316 2534 324
rect 2522 184 2534 316
rect 2842 324 2854 326
rect 2842 316 2844 324
rect 2852 316 2854 324
rect 2842 284 2854 316
rect 2842 276 2844 284
rect 2852 276 2854 284
rect 2842 274 2854 276
rect 2522 176 2524 184
rect 2532 176 2534 184
rect 2522 174 2534 176
rect 2650 224 2662 226
rect 2650 216 2652 224
rect 2660 216 2662 224
rect 2650 184 2662 216
rect 2650 176 2652 184
rect 2660 176 2662 184
rect 2650 174 2662 176
rect 2904 214 2952 606
rect 2970 944 2982 946
rect 2970 936 2972 944
rect 2980 936 2982 944
rect 2970 504 2982 936
rect 3034 924 3046 926
rect 3034 916 3036 924
rect 3044 916 3046 924
rect 3002 644 3014 646
rect 3002 636 3004 644
rect 3012 636 3014 644
rect 3002 604 3014 636
rect 3002 596 3004 604
rect 3012 596 3014 604
rect 3002 544 3014 596
rect 3002 536 3004 544
rect 3012 536 3014 544
rect 3002 534 3014 536
rect 3034 544 3046 916
rect 3034 536 3036 544
rect 3044 536 3046 544
rect 3034 534 3046 536
rect 3066 704 3078 706
rect 3066 696 3068 704
rect 3076 696 3078 704
rect 2970 496 2972 504
rect 2980 496 2982 504
rect 2970 494 2982 496
rect 3066 284 3078 696
rect 3290 644 3302 956
rect 3418 924 3430 1376
rect 3450 1284 3462 1536
rect 3450 1276 3452 1284
rect 3460 1276 3462 1284
rect 3450 1274 3462 1276
rect 3578 1284 3590 1736
rect 4090 1724 4102 1726
rect 4090 1716 4092 1724
rect 4100 1716 4102 1724
rect 4090 1444 4102 1716
rect 4090 1436 4092 1444
rect 4100 1436 4102 1444
rect 4090 1434 4102 1436
rect 4314 1704 4326 1706
rect 4314 1696 4316 1704
rect 4324 1696 4326 1704
rect 3578 1276 3580 1284
rect 3588 1276 3590 1284
rect 3578 1274 3590 1276
rect 3674 1364 3686 1366
rect 3674 1356 3676 1364
rect 3684 1356 3686 1364
rect 3674 1124 3686 1356
rect 4314 1204 4326 1696
rect 4314 1196 4316 1204
rect 4324 1196 4326 1204
rect 4314 1194 4326 1196
rect 4440 1614 4488 2006
rect 4440 1606 4444 1614
rect 4452 1606 4460 1614
rect 4468 1606 4476 1614
rect 4484 1606 4488 1614
rect 4440 1214 4488 1606
rect 4440 1206 4444 1214
rect 4452 1206 4460 1214
rect 4468 1206 4476 1214
rect 4484 1206 4488 1214
rect 3674 1116 3676 1124
rect 3684 1116 3686 1124
rect 3674 1114 3686 1116
rect 4090 1104 4102 1106
rect 4090 1096 4092 1104
rect 4100 1096 4102 1104
rect 4090 1064 4102 1096
rect 4090 1056 4092 1064
rect 4100 1056 4102 1064
rect 4090 1054 4102 1056
rect 3418 916 3420 924
rect 3428 916 3430 924
rect 3418 914 3430 916
rect 4440 814 4488 1206
rect 4538 1924 4550 1926
rect 4538 1916 4540 1924
rect 4548 1916 4550 1924
rect 4538 1184 4550 1916
rect 4538 1176 4540 1184
rect 4548 1176 4550 1184
rect 4538 1174 4550 1176
rect 4730 1524 4742 1526
rect 4730 1516 4732 1524
rect 4740 1516 4742 1524
rect 4440 806 4444 814
rect 4452 806 4460 814
rect 4468 806 4476 814
rect 4484 806 4488 814
rect 3290 636 3292 644
rect 3300 636 3302 644
rect 3290 634 3302 636
rect 4346 664 4358 666
rect 4346 656 4348 664
rect 4356 656 4358 664
rect 4346 544 4358 656
rect 4346 536 4348 544
rect 4356 536 4358 544
rect 4346 534 4358 536
rect 4378 524 4390 526
rect 4378 516 4380 524
rect 4388 516 4390 524
rect 3066 276 3068 284
rect 3076 276 3078 284
rect 3066 274 3078 276
rect 4250 384 4262 386
rect 4250 376 4252 384
rect 4260 376 4262 384
rect 2904 206 2908 214
rect 2916 206 2924 214
rect 2932 206 2940 214
rect 2948 206 2952 214
rect 2490 136 2492 144
rect 2500 136 2502 144
rect 2490 134 2502 136
rect 2682 164 2694 166
rect 2682 156 2684 164
rect 2692 156 2694 164
rect 2682 126 2694 156
rect 2394 76 2396 84
rect 2404 76 2406 84
rect 2394 74 2406 76
rect 2650 114 2694 126
rect 2650 84 2662 114
rect 2650 76 2652 84
rect 2660 76 2662 84
rect 2650 74 2662 76
rect 1352 6 1356 14
rect 1364 6 1372 14
rect 1380 6 1388 14
rect 1396 6 1400 14
rect 1352 0 1400 6
rect 2904 0 2952 206
rect 4250 84 4262 376
rect 4282 364 4294 366
rect 4282 356 4284 364
rect 4292 356 4294 364
rect 4282 204 4294 356
rect 4282 196 4284 204
rect 4292 196 4294 204
rect 4282 194 4294 196
rect 4346 344 4358 346
rect 4346 336 4348 344
rect 4356 336 4358 344
rect 4346 204 4358 336
rect 4346 196 4348 204
rect 4356 196 4358 204
rect 4346 194 4358 196
rect 4378 204 4390 516
rect 4378 196 4380 204
rect 4388 196 4390 204
rect 4378 194 4390 196
rect 4440 414 4488 806
rect 4602 1124 4614 1126
rect 4602 1116 4604 1124
rect 4612 1116 4614 1124
rect 4602 924 4614 1116
rect 4602 916 4604 924
rect 4612 916 4614 924
rect 4602 704 4614 916
rect 4634 984 4646 986
rect 4634 976 4636 984
rect 4644 976 4646 984
rect 4634 744 4646 976
rect 4730 964 4742 1516
rect 4922 1504 4934 2276
rect 4922 1496 4924 1504
rect 4932 1496 4934 1504
rect 4922 1494 4934 1496
rect 4986 1484 4998 2716
rect 5082 2524 5094 2526
rect 5082 2516 5084 2524
rect 5092 2516 5094 2524
rect 5082 2124 5094 2516
rect 5082 2116 5084 2124
rect 5092 2116 5094 2124
rect 5082 2114 5094 2116
rect 4986 1476 4988 1484
rect 4996 1476 4998 1484
rect 4986 1474 4998 1476
rect 5082 1704 5094 1706
rect 5082 1696 5084 1704
rect 5092 1696 5094 1704
rect 5082 1184 5094 1696
rect 5082 1176 5084 1184
rect 5092 1176 5094 1184
rect 5082 1174 5094 1176
rect 4762 1144 4774 1146
rect 4762 1136 4764 1144
rect 4772 1136 4774 1144
rect 4762 984 4774 1136
rect 4762 976 4764 984
rect 4772 976 4774 984
rect 4762 974 4774 976
rect 4794 1004 4806 1006
rect 4794 996 4796 1004
rect 4804 996 4806 1004
rect 4730 956 4732 964
rect 4740 956 4742 964
rect 4730 954 4742 956
rect 4634 736 4636 744
rect 4644 736 4646 744
rect 4634 734 4646 736
rect 4794 724 4806 996
rect 4794 716 4796 724
rect 4804 716 4806 724
rect 4794 714 4806 716
rect 4954 724 4966 726
rect 4954 716 4956 724
rect 4964 716 4966 724
rect 4602 696 4604 704
rect 4612 696 4614 704
rect 4602 694 4614 696
rect 4954 504 4966 716
rect 4986 704 4998 706
rect 4986 696 4988 704
rect 4996 696 4998 704
rect 4986 664 4998 696
rect 4986 656 4988 664
rect 4996 656 4998 664
rect 4986 654 4998 656
rect 5082 684 5094 686
rect 5082 676 5084 684
rect 5092 676 5094 684
rect 5082 544 5094 676
rect 5082 536 5084 544
rect 5092 536 5094 544
rect 5082 534 5094 536
rect 4954 496 4956 504
rect 4964 496 4966 504
rect 4954 494 4966 496
rect 4440 406 4444 414
rect 4452 406 4460 414
rect 4468 406 4476 414
rect 4484 406 4488 414
rect 4250 76 4252 84
rect 4260 76 4262 84
rect 4250 74 4262 76
rect 4440 14 4488 406
rect 4506 464 4518 466
rect 4506 456 4508 464
rect 4516 456 4518 464
rect 4506 264 4518 456
rect 4602 384 4614 386
rect 4602 376 4604 384
rect 4612 376 4614 384
rect 4602 366 4614 376
rect 4586 364 4614 366
rect 4586 356 4588 364
rect 4596 356 4614 364
rect 4586 354 4614 356
rect 4730 384 4742 386
rect 4730 376 4732 384
rect 4740 376 4742 384
rect 4730 304 4742 376
rect 4730 296 4732 304
rect 4740 296 4742 304
rect 4730 294 4742 296
rect 5114 304 5126 306
rect 5114 296 5116 304
rect 5124 296 5126 304
rect 4506 256 4508 264
rect 4516 256 4518 264
rect 4506 254 4518 256
rect 5082 264 5094 266
rect 5082 256 5084 264
rect 5092 256 5094 264
rect 5082 224 5094 256
rect 5082 216 5084 224
rect 5092 216 5094 224
rect 5082 214 5094 216
rect 5114 124 5126 296
rect 5178 224 5190 3636
rect 5338 3064 5350 3816
rect 5338 3056 5340 3064
rect 5348 3056 5350 3064
rect 5338 3054 5350 3056
rect 5370 3344 5382 3346
rect 5370 3336 5372 3344
rect 5380 3336 5382 3344
rect 5306 1704 5318 1706
rect 5306 1696 5308 1704
rect 5316 1696 5318 1704
rect 5306 1524 5318 1696
rect 5306 1516 5308 1524
rect 5316 1516 5318 1524
rect 5306 1514 5318 1516
rect 5274 1164 5286 1166
rect 5274 1156 5276 1164
rect 5284 1156 5286 1164
rect 5210 1104 5222 1106
rect 5210 1096 5212 1104
rect 5220 1096 5222 1104
rect 5210 524 5222 1096
rect 5210 516 5212 524
rect 5220 516 5222 524
rect 5210 514 5222 516
rect 5274 504 5286 1156
rect 5370 1164 5382 3336
rect 5658 3324 5670 3326
rect 5658 3316 5660 3324
rect 5668 3316 5670 3324
rect 5530 3244 5542 3246
rect 5530 3236 5532 3244
rect 5540 3236 5542 3244
rect 5530 1644 5542 3236
rect 5530 1636 5532 1644
rect 5540 1636 5542 1644
rect 5530 1634 5542 1636
rect 5626 2784 5638 2786
rect 5626 2776 5628 2784
rect 5636 2776 5638 2784
rect 5530 1464 5542 1466
rect 5530 1456 5532 1464
rect 5540 1456 5542 1464
rect 5498 1424 5510 1426
rect 5498 1416 5500 1424
rect 5508 1416 5510 1424
rect 5370 1156 5372 1164
rect 5380 1156 5382 1164
rect 5370 1154 5382 1156
rect 5402 1244 5414 1246
rect 5402 1236 5404 1244
rect 5412 1236 5414 1244
rect 5402 644 5414 1236
rect 5402 636 5404 644
rect 5412 636 5414 644
rect 5402 634 5414 636
rect 5274 496 5276 504
rect 5284 496 5286 504
rect 5274 494 5286 496
rect 5498 504 5510 1416
rect 5498 496 5500 504
rect 5508 496 5510 504
rect 5498 494 5510 496
rect 5530 444 5542 1456
rect 5626 1084 5638 2776
rect 5658 1844 5670 3316
rect 5818 3044 5830 3046
rect 5818 3036 5820 3044
rect 5828 3036 5830 3044
rect 5658 1836 5660 1844
rect 5668 1836 5670 1844
rect 5658 1834 5670 1836
rect 5786 2964 5798 2966
rect 5786 2956 5788 2964
rect 5796 2956 5798 2964
rect 5786 1184 5798 2956
rect 5786 1176 5788 1184
rect 5796 1176 5798 1184
rect 5786 1174 5798 1176
rect 5626 1076 5628 1084
rect 5636 1076 5638 1084
rect 5626 1074 5638 1076
rect 5530 436 5532 444
rect 5540 436 5542 444
rect 5530 434 5542 436
rect 5754 524 5766 526
rect 5754 516 5756 524
rect 5764 516 5766 524
rect 5178 216 5180 224
rect 5188 216 5190 224
rect 5178 214 5190 216
rect 5690 304 5702 306
rect 5690 296 5692 304
rect 5700 296 5702 304
rect 5690 204 5702 296
rect 5754 224 5766 516
rect 5818 284 5830 3036
rect 5818 276 5820 284
rect 5828 276 5830 284
rect 5818 274 5830 276
rect 5754 216 5756 224
rect 5764 216 5766 224
rect 5754 214 5766 216
rect 5690 196 5692 204
rect 5700 196 5702 204
rect 5690 194 5702 196
rect 5114 116 5116 124
rect 5124 116 5126 124
rect 5114 114 5126 116
rect 4440 6 4444 14
rect 4452 6 4460 14
rect 4468 6 4476 14
rect 4484 6 4488 14
rect 4440 0 4488 6
use NAND2X1  NAND2X1_61
timestamp 1744230924
transform 1 0 88 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_62
timestamp 1744230924
transform 1 0 40 0 1 210
box -4 -6 52 206
use INVX1  INVX1_51
timestamp 1744230924
transform 1 0 8 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_74
timestamp 1744230924
transform -1 0 168 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_4
timestamp 1744230924
transform -1 0 104 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_50
timestamp 1744230924
transform 1 0 8 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_73
timestamp 1744230924
transform -1 0 264 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_11
timestamp 1744230924
transform -1 0 200 0 1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_30
timestamp 1744230924
transform -1 0 280 0 -1 210
box -4 -6 116 206
use OAI21X1  OAI21X1_86
timestamp 1744230924
transform -1 0 424 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_67
timestamp 1744230924
transform 1 0 312 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_1
timestamp 1744230924
transform -1 0 312 0 1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_28
timestamp 1744230924
transform -1 0 392 0 -1 210
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_134
timestamp 1744230924
transform 1 0 392 0 -1 210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_136
timestamp 1744230924
transform 1 0 584 0 -1 210
box -4 -6 196 206
use AOI21X1  AOI21X1_13
timestamp 1744230924
transform 1 0 424 0 1 210
box -4 -6 68 206
use INVX1  INVX1_58
timestamp 1744230924
transform 1 0 488 0 1 210
box -4 -6 36 206
use BUFX4  BUFX4_7
timestamp 1744230924
transform 1 0 520 0 1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_31
timestamp 1744230924
transform -1 0 696 0 1 210
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_75
timestamp 1744230924
transform 1 0 696 0 1 210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_133
timestamp 1744230924
transform 1 0 776 0 -1 210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_135
timestamp 1744230924
transform 1 0 968 0 -1 210
box -4 -6 196 206
use XNOR2X1  XNOR2X1_90
timestamp 1744230924
transform 1 0 888 0 1 210
box -4 -6 116 206
use OAI21X1  OAI21X1_259
timestamp 1744230924
transform -1 0 1064 0 1 210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_76
timestamp 1744230924
transform 1 0 1064 0 1 210
box -4 -6 196 206
use XNOR2X1  XNOR2X1_93
timestamp 1744230924
transform -1 0 1368 0 1 210
box -4 -6 116 206
use XOR2X1  XOR2X1_26
timestamp 1744230924
transform -1 0 1528 0 1 210
box -4 -6 116 206
use FILL  FILL_1_0_2
timestamp 1744230924
transform -1 0 1416 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1744230924
transform -1 0 1400 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_0
timestamp 1744230924
transform -1 0 1384 0 1 210
box -4 -6 20 206
use XNOR2X1  XNOR2X1_87
timestamp 1744230924
transform 1 0 1400 0 -1 210
box -4 -6 116 206
use FILL  FILL_0_0_2
timestamp 1744230924
transform 1 0 1384 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1744230924
transform 1 0 1368 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_0
timestamp 1744230924
transform 1 0 1352 0 -1 210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_78
timestamp 1744230924
transform 1 0 1160 0 -1 210
box -4 -6 196 206
use NAND2X1  NAND2X1_176
timestamp 1744230924
transform 1 0 1528 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_244
timestamp 1744230924
transform 1 0 1512 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_178
timestamp 1744230924
transform 1 0 1608 0 1 210
box -4 -6 52 206
use INVX1  INVX1_152
timestamp 1744230924
transform 1 0 1576 0 1 210
box -4 -6 36 206
use INVX1  INVX1_153
timestamp 1744230924
transform 1 0 1608 0 -1 210
box -4 -6 36 206
use INVX1  INVX1_158
timestamp 1744230924
transform -1 0 1608 0 -1 210
box -4 -6 36 206
use OAI22X1  OAI22X1_11
timestamp 1744230924
transform -1 0 1736 0 1 210
box -4 -6 84 206
use AOI21X1  AOI21X1_52
timestamp 1744230924
transform -1 0 1752 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_129
timestamp 1744230924
transform -1 0 1688 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_234
timestamp 1744230924
transform -1 0 1864 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_233
timestamp 1744230924
transform 1 0 1736 0 1 210
box -4 -6 68 206
use BUFX4  BUFX4_25
timestamp 1744230924
transform 1 0 1752 0 -1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_82
timestamp 1744230924
transform -1 0 1976 0 1 210
box -4 -6 116 206
use OAI21X1  OAI21X1_236
timestamp 1744230924
transform 1 0 1928 0 -1 210
box -4 -6 68 206
use XOR2X1  XOR2X1_27
timestamp 1744230924
transform 1 0 1816 0 -1 210
box -4 -6 116 206
use AND2X2  AND2X2_11
timestamp 1744230924
transform 1 0 2040 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_53
timestamp 1744230924
transform 1 0 1976 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_238
timestamp 1744230924
transform 1 0 1992 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_184
timestamp 1744230924
transform 1 0 2152 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_182
timestamp 1744230924
transform -1 0 2152 0 1 210
box -4 -6 52 206
use INVX1  INVX1_155
timestamp 1744230924
transform -1 0 2200 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_130
timestamp 1744230924
transform 1 0 2120 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_237
timestamp 1744230924
transform -1 0 2120 0 -1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_85
timestamp 1744230924
transform 1 0 2200 0 1 210
box -4 -6 116 206
use NAND2X1  NAND2X1_188
timestamp 1744230924
transform 1 0 2248 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_183
timestamp 1744230924
transform -1 0 2248 0 -1 210
box -4 -6 52 206
use AOI22X1  AOI22X1_27
timestamp 1744230924
transform -1 0 2488 0 1 210
box -4 -6 84 206
use NOR2X1  NOR2X1_134
timestamp 1744230924
transform 1 0 2360 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_186
timestamp 1744230924
transform -1 0 2360 0 1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_84
timestamp 1744230924
transform 1 0 2328 0 -1 210
box -4 -6 116 206
use INVX1  INVX1_154
timestamp 1744230924
transform -1 0 2328 0 -1 210
box -4 -6 36 206
use AOI22X1  AOI22X1_29
timestamp 1744230924
transform 1 0 2488 0 1 210
box -4 -6 84 206
use NAND2X1  NAND2X1_185
timestamp 1744230924
transform 1 0 2488 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_180
timestamp 1744230924
transform -1 0 2488 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_179
timestamp 1744230924
transform -1 0 2664 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_181
timestamp 1744230924
transform -1 0 2616 0 1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_83
timestamp 1744230924
transform -1 0 2760 0 -1 210
box -4 -6 116 206
use NAND2X1  NAND2X1_177
timestamp 1744230924
transform 1 0 2600 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_235
timestamp 1744230924
transform 1 0 2536 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_241
timestamp 1744230924
transform -1 0 2792 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_242
timestamp 1744230924
transform 1 0 2664 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_249
timestamp 1744230924
transform 1 0 2760 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_240
timestamp 1744230924
transform 1 0 2856 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_239
timestamp 1744230924
transform 1 0 2792 0 1 210
box -4 -6 68 206
use XOR2X1  XOR2X1_28
timestamp 1744230924
transform -1 0 2936 0 -1 210
box -4 -6 116 206
use OAI21X1  OAI21X1_251
timestamp 1744230924
transform -1 0 3032 0 1 210
box -4 -6 68 206
use FILL  FILL_1_1_2
timestamp 1744230924
transform -1 0 2968 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_1
timestamp 1744230924
transform -1 0 2952 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_0
timestamp 1744230924
transform -1 0 2936 0 1 210
box -4 -6 20 206
use NAND2X1  NAND2X1_189
timestamp 1744230924
transform 1 0 2984 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_1_2
timestamp 1744230924
transform 1 0 2968 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1744230924
transform 1 0 2952 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_0
timestamp 1744230924
transform 1 0 2936 0 -1 210
box -4 -6 20 206
use OAI21X1  OAI21X1_246
timestamp 1744230924
transform 1 0 3080 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_131
timestamp 1744230924
transform 1 0 3032 0 1 210
box -4 -6 52 206
use INVX1  INVX1_161
timestamp 1744230924
transform 1 0 3096 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_245
timestamp 1744230924
transform -1 0 3096 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_247
timestamp 1744230924
transform -1 0 3208 0 1 210
box -4 -6 68 206
use MUX2X1  MUX2X1_11
timestamp 1744230924
transform -1 0 3272 0 -1 210
box -4 -6 100 206
use NAND2X1  NAND2X1_191
timestamp 1744230924
transform -1 0 3176 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_162
timestamp 1744230924
transform 1 0 3240 0 1 210
box -4 -6 36 206
use INVX1  INVX1_166
timestamp 1744230924
transform -1 0 3240 0 1 210
box -4 -6 36 206
use AOI21X1  AOI21X1_54
timestamp 1744230924
transform -1 0 3496 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_133
timestamp 1744230924
transform -1 0 3432 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_250
timestamp 1744230924
transform -1 0 3384 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_132
timestamp 1744230924
transform 1 0 3272 0 1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_88
timestamp 1744230924
transform 1 0 3272 0 -1 210
box -4 -6 116 206
use INVX1  INVX1_157
timestamp 1744230924
transform 1 0 3608 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_243
timestamp 1744230924
transform 1 0 3544 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_187
timestamp 1744230924
transform -1 0 3544 0 1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_85
timestamp 1744230924
transform 1 0 3576 0 -1 210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_86
timestamp 1744230924
transform 1 0 3384 0 -1 210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_88
timestamp 1744230924
transform 1 0 3768 0 -1 210
box -4 -6 196 206
use BUFX4  BUFX4_18
timestamp 1744230924
transform 1 0 3960 0 -1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_86
timestamp 1744230924
transform -1 0 3752 0 1 210
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_87
timestamp 1744230924
transform 1 0 3752 0 1 210
box -4 -6 196 206
use BUFX4  BUFX4_17
timestamp 1744230924
transform 1 0 3944 0 1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_61
timestamp 1744230924
transform 1 0 4008 0 1 210
box -4 -6 116 206
use XOR2X1  XOR2X1_19
timestamp 1744230924
transform -1 0 4136 0 -1 210
box -4 -6 116 206
use OAI21X1  OAI21X1_180
timestamp 1744230924
transform 1 0 4168 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_141
timestamp 1744230924
transform 1 0 4120 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_182
timestamp 1744230924
transform 1 0 4168 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_125
timestamp 1744230924
transform 1 0 4136 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_110
timestamp 1744230924
transform 1 0 4328 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_143
timestamp 1744230924
transform 1 0 4280 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_145
timestamp 1744230924
transform 1 0 4232 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_142
timestamp 1744230924
transform 1 0 4296 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_183
timestamp 1744230924
transform -1 0 4296 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_177
timestamp 1744230924
transform 1 0 4376 0 1 210
box -4 -6 68 206
use BUFX4  BUFX4_19
timestamp 1744230924
transform 1 0 4344 0 -1 210
box -4 -6 68 206
use FILL  FILL_1_2_2
timestamp 1744230924
transform 1 0 4472 0 1 210
box -4 -6 20 206
use FILL  FILL_1_2_1
timestamp 1744230924
transform 1 0 4456 0 1 210
box -4 -6 20 206
use FILL  FILL_1_2_0
timestamp 1744230924
transform 1 0 4440 0 1 210
box -4 -6 20 206
use FILL  FILL_0_2_2
timestamp 1744230924
transform 1 0 4472 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_2_1
timestamp 1744230924
transform 1 0 4456 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_2_0
timestamp 1744230924
transform 1 0 4440 0 -1 210
box -4 -6 20 206
use INVX1  INVX1_124
timestamp 1744230924
transform 1 0 4408 0 -1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_140
timestamp 1744230924
transform 1 0 4536 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_138
timestamp 1744230924
transform 1 0 4488 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_147
timestamp 1744230924
transform -1 0 4584 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_139
timestamp 1744230924
transform 1 0 4488 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_181
timestamp 1744230924
transform -1 0 4648 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_98
timestamp 1744230924
transform -1 0 4632 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_144
timestamp 1744230924
transform -1 0 4696 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_192
timestamp 1744230924
transform 1 0 4632 0 -1 210
box -4 -6 68 206
use AOI22X1  AOI22X1_19
timestamp 1744230924
transform -1 0 4856 0 1 210
box -4 -6 84 206
use AOI22X1  AOI22X1_20
timestamp 1744230924
transform -1 0 4776 0 1 210
box -4 -6 84 206
use OAI21X1  OAI21X1_187
timestamp 1744230924
transform 1 0 4808 0 -1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_63
timestamp 1744230924
transform 1 0 4696 0 -1 210
box -4 -6 116 206
use OAI21X1  OAI21X1_194
timestamp 1744230924
transform -1 0 4984 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_178
timestamp 1744230924
transform 1 0 4856 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_189
timestamp 1744230924
transform -1 0 4936 0 -1 210
box -4 -6 68 206
use AOI22X1  AOI22X1_21
timestamp 1744230924
transform 1 0 5048 0 1 210
box -4 -6 84 206
use OAI21X1  OAI21X1_179
timestamp 1744230924
transform -1 0 5048 0 1 210
box -4 -6 68 206
use OR2X2  OR2X2_12
timestamp 1744230924
transform 1 0 5000 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_188
timestamp 1744230924
transform 1 0 4936 0 -1 210
box -4 -6 68 206
use AOI22X1  AOI22X1_18
timestamp 1744230924
transform 1 0 5160 0 1 210
box -4 -6 84 206
use INVX1  INVX1_133
timestamp 1744230924
transform -1 0 5160 0 1 210
box -4 -6 36 206
use BUFX4  BUFX4_20
timestamp 1744230924
transform -1 0 5208 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_126
timestamp 1744230924
transform 1 0 5112 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_100
timestamp 1744230924
transform 1 0 5064 0 -1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_60
timestamp 1744230924
transform -1 0 5400 0 1 210
box -4 -6 116 206
use NOR2X1  NOR2X1_107
timestamp 1744230924
transform 1 0 5240 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_193
timestamp 1744230924
transform -1 0 5304 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_128
timestamp 1744230924
transform 1 0 5208 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_103
timestamp 1744230924
transform -1 0 5448 0 1 210
box -4 -6 52 206
use INVX2  INVX2_20
timestamp 1744230924
transform 1 0 5400 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_99
timestamp 1744230924
transform 1 0 5352 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_101
timestamp 1744230924
transform -1 0 5352 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_146
timestamp 1744230924
transform -1 0 5560 0 1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_40
timestamp 1744230924
transform -1 0 5512 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_102
timestamp 1744230924
transform -1 0 5544 0 -1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_39
timestamp 1744230924
transform -1 0 5496 0 -1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_62
timestamp 1744230924
transform -1 0 5768 0 1 210
box -4 -6 116 206
use OAI21X1  OAI21X1_184
timestamp 1744230924
transform -1 0 5656 0 1 210
box -4 -6 68 206
use INVX1  INVX1_137
timestamp 1744230924
transform -1 0 5592 0 1 210
box -4 -6 36 206
use XNOR2X1  XNOR2X1_64
timestamp 1744230924
transform -1 0 5720 0 -1 210
box -4 -6 116 206
use AND2X2  AND2X2_9
timestamp 1744230924
transform 1 0 5544 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_185
timestamp 1744230924
transform 1 0 5768 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_186
timestamp 1744230924
transform 1 0 5720 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_26
timestamp 1744230924
transform 1 0 5784 0 -1 210
box -4 -6 52 206
use FILL  FILL_1_1
timestamp 1744230924
transform -1 0 5848 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_2
timestamp 1744230924
transform -1 0 5864 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_1
timestamp 1744230924
transform 1 0 5832 0 1 210
box -4 -6 20 206
use FILL  FILL_2_2
timestamp 1744230924
transform 1 0 5848 0 1 210
box -4 -6 20 206
use NOR2X1  NOR2X1_40
timestamp 1744230924
transform -1 0 56 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_64
timestamp 1744230924
transform 1 0 56 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_60
timestamp 1744230924
transform 1 0 104 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_36
timestamp 1744230924
transform 1 0 152 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_58
timestamp 1744230924
transform 1 0 200 0 -1 610
box -4 -6 52 206
use AOI22X1  AOI22X1_6
timestamp 1744230924
transform -1 0 328 0 -1 610
box -4 -6 84 206
use INVX1  INVX1_55
timestamp 1744230924
transform 1 0 328 0 -1 610
box -4 -6 36 206
use AOI22X1  AOI22X1_5
timestamp 1744230924
transform -1 0 440 0 -1 610
box -4 -6 84 206
use NAND3X1  NAND3X1_6
timestamp 1744230924
transform -1 0 504 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_79
timestamp 1744230924
transform -1 0 568 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_53
timestamp 1744230924
transform 1 0 568 0 -1 610
box -4 -6 36 206
use INVX1  INVX1_61
timestamp 1744230924
transform 1 0 600 0 -1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_14
timestamp 1744230924
transform -1 0 696 0 -1 610
box -4 -6 68 206
use MUX2X1  MUX2X1_1
timestamp 1744230924
transform -1 0 792 0 -1 610
box -4 -6 100 206
use OAI21X1  OAI21X1_78
timestamp 1744230924
transform 1 0 792 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_63
timestamp 1744230924
transform -1 0 904 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_195
timestamp 1744230924
transform -1 0 952 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_193
timestamp 1744230924
transform -1 0 1000 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_258
timestamp 1744230924
transform 1 0 1000 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_54
timestamp 1744230924
transform 1 0 1064 0 -1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_142
timestamp 1744230924
transform 1 0 1160 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_261
timestamp 1744230924
transform 1 0 1096 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_169
timestamp 1744230924
transform -1 0 1240 0 -1 610
box -4 -6 36 206
use INVX1  INVX1_168
timestamp 1744230924
transform -1 0 1336 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_263
timestamp 1744230924
transform -1 0 1304 0 -1 610
box -4 -6 68 206
use FILL  FILL_2_0_2
timestamp 1744230924
transform 1 0 1368 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1744230924
transform 1 0 1352 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_0
timestamp 1744230924
transform 1 0 1336 0 -1 610
box -4 -6 20 206
use INVX1  INVX1_170
timestamp 1744230924
transform -1 0 1480 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_260
timestamp 1744230924
transform 1 0 1384 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_57
timestamp 1744230924
transform -1 0 1544 0 -1 610
box -4 -6 68 206
use XOR2X1  XOR2X1_29
timestamp 1744230924
transform -1 0 1656 0 -1 610
box -4 -6 116 206
use XNOR2X1  XNOR2X1_92
timestamp 1744230924
transform -1 0 1768 0 -1 610
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_77
timestamp 1744230924
transform 1 0 1768 0 -1 610
box -4 -6 196 206
use INVX2  INVX2_9
timestamp 1744230924
transform -1 0 1992 0 -1 610
box -4 -6 36 206
use XOR2X1  XOR2X1_25
timestamp 1744230924
transform -1 0 2104 0 -1 610
box -4 -6 116 206
use OAI21X1  OAI21X1_130
timestamp 1744230924
transform -1 0 2168 0 -1 610
box -4 -6 68 206
use INVX2  INVX2_10
timestamp 1744230924
transform 1 0 2168 0 -1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_67
timestamp 1744230924
transform -1 0 2248 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_68
timestamp 1744230924
transform -1 0 2296 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_66
timestamp 1744230924
transform 1 0 2296 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_134
timestamp 1744230924
transform 1 0 2344 0 -1 610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_44
timestamp 1744230924
transform 1 0 2408 0 -1 610
box -4 -6 116 206
use BUFX4  BUFX4_24
timestamp 1744230924
transform 1 0 2520 0 -1 610
box -4 -6 68 206
use BUFX2  BUFX2_6
timestamp 1744230924
transform 1 0 2584 0 -1 610
box -4 -6 52 206
use BUFX4  BUFX4_26
timestamp 1744230924
transform 1 0 2632 0 -1 610
box -4 -6 68 206
use BUFX2  BUFX2_7
timestamp 1744230924
transform -1 0 2744 0 -1 610
box -4 -6 52 206
use INVX2  INVX2_26
timestamp 1744230924
transform -1 0 2776 0 -1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_135
timestamp 1744230924
transform -1 0 2824 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_136
timestamp 1744230924
transform -1 0 2872 0 -1 610
box -4 -6 52 206
use FILL  FILL_2_1_0
timestamp 1744230924
transform 1 0 2872 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1744230924
transform 1 0 2888 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1744230924
transform 1 0 2904 0 -1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_255
timestamp 1744230924
transform 1 0 2920 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_56
timestamp 1744230924
transform -1 0 3048 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_190
timestamp 1744230924
transform 1 0 3048 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_156
timestamp 1744230924
transform -1 0 3128 0 -1 610
box -4 -6 36 206
use AOI22X1  AOI22X1_30
timestamp 1744230924
transform 1 0 3128 0 -1 610
box -4 -6 84 206
use AOI22X1  AOI22X1_28
timestamp 1744230924
transform 1 0 3208 0 -1 610
box -4 -6 84 206
use NOR2X1  NOR2X1_139
timestamp 1744230924
transform -1 0 3336 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_8
timestamp 1744230924
transform 1 0 3336 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_248
timestamp 1744230924
transform 1 0 3384 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_252
timestamp 1744230924
transform -1 0 3512 0 -1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_89
timestamp 1744230924
transform 1 0 3512 0 -1 610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_144
timestamp 1744230924
transform 1 0 3704 0 -1 610
box -4 -6 196 206
use INVX1  INVX1_62
timestamp 1744230924
transform 1 0 3896 0 -1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_69
timestamp 1744230924
transform -1 0 3976 0 -1 610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_84
timestamp 1744230924
transform 1 0 3976 0 -1 610
box -4 -6 196 206
use BUFX4  BUFX4_16
timestamp 1744230924
transform 1 0 4168 0 -1 610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_65
timestamp 1744230924
transform 1 0 4232 0 -1 610
box -4 -6 116 206
use OAI21X1  OAI21X1_191
timestamp 1744230924
transform 1 0 4344 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_129
timestamp 1744230924
transform 1 0 4408 0 -1 610
box -4 -6 36 206
use FILL  FILL_2_2_0
timestamp 1744230924
transform 1 0 4440 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_2_1
timestamp 1744230924
transform 1 0 4456 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_2_2
timestamp 1744230924
transform 1 0 4472 0 -1 610
box -4 -6 20 206
use NAND2X1  NAND2X1_136
timestamp 1744230924
transform 1 0 4488 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_176
timestamp 1744230924
transform -1 0 4600 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_137
timestamp 1744230924
transform 1 0 4600 0 -1 610
box -4 -6 52 206
use AND2X2  AND2X2_8
timestamp 1744230924
transform -1 0 4712 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_38
timestamp 1744230924
transform 1 0 4712 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_104
timestamp 1744230924
transform 1 0 4776 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_106
timestamp 1744230924
transform 1 0 4824 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_196
timestamp 1744230924
transform 1 0 4872 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_132
timestamp 1744230924
transform 1 0 4936 0 -1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_42
timestamp 1744230924
transform -1 0 5032 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_41
timestamp 1744230924
transform -1 0 5096 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_127
timestamp 1744230924
transform -1 0 5128 0 -1 610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_66
timestamp 1744230924
transform -1 0 5240 0 -1 610
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_94
timestamp 1744230924
transform 1 0 5240 0 -1 610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_95
timestamp 1744230924
transform -1 0 5624 0 -1 610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_96
timestamp 1744230924
transform -1 0 5816 0 -1 610
box -4 -6 196 206
use FILL  FILL_3_1
timestamp 1744230924
transform -1 0 5832 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_2
timestamp 1744230924
transform -1 0 5848 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_3
timestamp 1744230924
transform -1 0 5864 0 -1 610
box -4 -6 20 206
use XNOR2X1  XNOR2X1_29
timestamp 1744230924
transform 1 0 8 0 1 610
box -4 -6 116 206
use NAND2X1  NAND2X1_59
timestamp 1744230924
transform -1 0 168 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_77
timestamp 1744230924
transform 1 0 168 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_66
timestamp 1744230924
transform 1 0 232 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_83
timestamp 1744230924
transform -1 0 344 0 1 610
box -4 -6 68 206
use INVX2  INVX2_6
timestamp 1744230924
transform -1 0 376 0 1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_38
timestamp 1744230924
transform 1 0 376 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_85
timestamp 1744230924
transform 1 0 424 0 1 610
box -4 -6 68 206
use INVX1  INVX1_59
timestamp 1744230924
transform -1 0 520 0 1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_39
timestamp 1744230924
transform -1 0 568 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_37
timestamp 1744230924
transform -1 0 616 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_84
timestamp 1744230924
transform 1 0 616 0 1 610
box -4 -6 68 206
use INVX8  INVX8_2
timestamp 1744230924
transform -1 0 760 0 1 610
box -4 -6 84 206
use INVX1  INVX1_52
timestamp 1744230924
transform 1 0 760 0 1 610
box -4 -6 36 206
use BUFX4  BUFX4_5
timestamp 1744230924
transform 1 0 792 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_194
timestamp 1744230924
transform 1 0 856 0 1 610
box -4 -6 52 206
use INVX1  INVX1_167
timestamp 1744230924
transform -1 0 936 0 1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_196
timestamp 1744230924
transform 1 0 936 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_197
timestamp 1744230924
transform 1 0 984 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_262
timestamp 1744230924
transform 1 0 1032 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_143
timestamp 1744230924
transform -1 0 1144 0 1 610
box -4 -6 52 206
use AOI21X1  AOI21X1_58
timestamp 1744230924
transform -1 0 1208 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_265
timestamp 1744230924
transform 1 0 1208 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_202
timestamp 1744230924
transform -1 0 1320 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_266
timestamp 1744230924
transform -1 0 1384 0 1 610
box -4 -6 68 206
use FILL  FILL_3_0_0
timestamp 1744230924
transform -1 0 1400 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1744230924
transform -1 0 1416 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1744230924
transform -1 0 1432 0 1 610
box -4 -6 20 206
use XNOR2X1  XNOR2X1_91
timestamp 1744230924
transform -1 0 1544 0 1 610
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_79
timestamp 1744230924
transform 1 0 1544 0 1 610
box -4 -6 196 206
use OAI21X1  OAI21X1_127
timestamp 1744230924
transform 1 0 1736 0 1 610
box -4 -6 68 206
use INVX1  INVX1_83
timestamp 1744230924
transform 1 0 1800 0 1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_63
timestamp 1744230924
transform -1 0 1880 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_100
timestamp 1744230924
transform 1 0 1880 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_60
timestamp 1744230924
transform -1 0 1976 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_132
timestamp 1744230924
transform 1 0 1976 0 1 610
box -4 -6 68 206
use INVX1  INVX1_89
timestamp 1744230924
transform -1 0 2072 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_131
timestamp 1744230924
transform -1 0 2136 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_21
timestamp 1744230924
transform -1 0 2200 0 1 610
box -4 -6 68 206
use INVX1  INVX1_87
timestamp 1744230924
transform 1 0 2200 0 1 610
box -4 -6 36 206
use INVX1  INVX1_93
timestamp 1744230924
transform 1 0 2232 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_135
timestamp 1744230924
transform 1 0 2264 0 1 610
box -4 -6 68 206
use INVX1  INVX1_91
timestamp 1744230924
transform -1 0 2360 0 1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_22
timestamp 1744230924
transform -1 0 2424 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_8
timestamp 1744230924
transform -1 0 2488 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_136
timestamp 1744230924
transform 1 0 2488 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_101
timestamp 1744230924
transform 1 0 2552 0 1 610
box -4 -6 52 206
use INVX1  INVX1_92
timestamp 1744230924
transform -1 0 2632 0 1 610
box -4 -6 36 206
use INVX1  INVX1_159
timestamp 1744230924
transform 1 0 2632 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_253
timestamp 1744230924
transform 1 0 2664 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_257
timestamp 1744230924
transform -1 0 2792 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_137
timestamp 1744230924
transform 1 0 2792 0 1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_18
timestamp 1744230924
transform 1 0 2840 0 1 610
box -4 -6 68 206
use INVX1  INVX1_164
timestamp 1744230924
transform 1 0 2952 0 1 610
box -4 -6 36 206
use FILL  FILL_3_1_2
timestamp 1744230924
transform 1 0 2936 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1744230924
transform 1 0 2920 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_0
timestamp 1744230924
transform 1 0 2904 0 1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_256
timestamp 1744230924
transform -1 0 3048 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_254
timestamp 1744230924
transform 1 0 3080 0 1 610
box -4 -6 68 206
use INVX1  INVX1_165
timestamp 1744230924
transform -1 0 3080 0 1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_55
timestamp 1744230924
transform -1 0 3240 0 1 610
box -4 -6 68 206
use INVX1  INVX1_163
timestamp 1744230924
transform -1 0 3176 0 1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_138
timestamp 1744230924
transform -1 0 3288 0 1 610
box -4 -6 52 206
use INVX1  INVX1_160
timestamp 1744230924
transform -1 0 3320 0 1 610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_89
timestamp 1744230924
transform -1 0 3432 0 1 610
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_83
timestamp 1744230924
transform 1 0 3432 0 1 610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_137
timestamp 1744230924
transform 1 0 3624 0 1 610
box -4 -6 196 206
use NAND2X1  NAND2X1_73
timestamp 1744230924
transform 1 0 3816 0 1 610
box -4 -6 52 206
use INVX1  INVX1_63
timestamp 1744230924
transform 1 0 3864 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_88
timestamp 1744230924
transform 1 0 3896 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_87
timestamp 1744230924
transform -1 0 4024 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_68
timestamp 1744230924
transform 1 0 4024 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_70
timestamp 1744230924
transform 1 0 4072 0 1 610
box -4 -6 52 206
use INVX2  INVX2_7
timestamp 1744230924
transform 1 0 4120 0 1 610
box -4 -6 36 206
use INVX1  INVX1_123
timestamp 1744230924
transform 1 0 4152 0 1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_97
timestamp 1744230924
transform -1 0 4232 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_135
timestamp 1744230924
transform 1 0 4232 0 1 610
box -4 -6 52 206
use INVX1  INVX1_122
timestamp 1744230924
transform -1 0 4312 0 1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_37
timestamp 1744230924
transform 1 0 4312 0 1 610
box -4 -6 68 206
use XOR2X1  XOR2X1_18
timestamp 1744230924
transform -1 0 4488 0 1 610
box -4 -6 116 206
use FILL  FILL_3_2_0
timestamp 1744230924
transform -1 0 4504 0 1 610
box -4 -6 20 206
use FILL  FILL_3_2_1
timestamp 1744230924
transform -1 0 4520 0 1 610
box -4 -6 20 206
use FILL  FILL_3_2_2
timestamp 1744230924
transform -1 0 4536 0 1 610
box -4 -6 20 206
use OAI22X1  OAI22X1_9
timestamp 1744230924
transform -1 0 4616 0 1 610
box -4 -6 84 206
use XNOR2X1  XNOR2X1_59
timestamp 1744230924
transform 1 0 4616 0 1 610
box -4 -6 116 206
use OAI21X1  OAI21X1_198
timestamp 1744230924
transform 1 0 4728 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_105
timestamp 1744230924
transform 1 0 4792 0 1 610
box -4 -6 52 206
use INVX1  INVX1_131
timestamp 1744230924
transform 1 0 4840 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_199
timestamp 1744230924
transform -1 0 4936 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_200
timestamp 1744230924
transform -1 0 5000 0 1 610
box -4 -6 68 206
use INVX1  INVX1_130
timestamp 1744230924
transform 1 0 5000 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_197
timestamp 1744230924
transform -1 0 5096 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_109
timestamp 1744230924
transform -1 0 5144 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_108
timestamp 1744230924
transform 1 0 5144 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_190
timestamp 1744230924
transform 1 0 5192 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_195
timestamp 1744230924
transform -1 0 5320 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_5
timestamp 1744230924
transform -1 0 5368 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_2
timestamp 1744230924
transform 1 0 5368 0 1 610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_104
timestamp 1744230924
transform 1 0 5416 0 1 610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_41
timestamp 1744230924
transform 1 0 5608 0 1 610
box -4 -6 196 206
use BUFX2  BUFX2_24
timestamp 1744230924
transform 1 0 5800 0 1 610
box -4 -6 52 206
use FILL  FILL_4_1
timestamp 1744230924
transform 1 0 5848 0 1 610
box -4 -6 20 206
use INVX2  INVX2_5
timestamp 1744230924
transform 1 0 8 0 -1 1010
box -4 -6 36 206
use INVX1  INVX1_56
timestamp 1744230924
transform 1 0 40 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_5
timestamp 1744230924
transform 1 0 72 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_82
timestamp 1744230924
transform 1 0 136 0 -1 1010
box -4 -6 68 206
use BUFX4  BUFX4_6
timestamp 1744230924
transform -1 0 264 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_147
timestamp 1744230924
transform 1 0 264 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_60
timestamp 1744230924
transform 1 0 312 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_280
timestamp 1744230924
transform 1 0 344 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_181
timestamp 1744230924
transform 1 0 408 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_281
timestamp 1744230924
transform -1 0 504 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_182
timestamp 1744230924
transform 1 0 504 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_19
timestamp 1744230924
transform 1 0 536 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_66
timestamp 1744230924
transform -1 0 664 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_282
timestamp 1744230924
transform 1 0 664 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_209
timestamp 1744230924
transform 1 0 728 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_199
timestamp 1744230924
transform 1 0 776 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_171
timestamp 1744230924
transform -1 0 856 0 -1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_201
timestamp 1744230924
transform -1 0 904 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_200
timestamp 1744230924
transform 1 0 904 0 -1 1010
box -4 -6 52 206
use AOI21X1  AOI21X1_59
timestamp 1744230924
transform 1 0 952 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_60
timestamp 1744230924
transform 1 0 1016 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_64
timestamp 1744230924
transform 1 0 1080 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_174
timestamp 1744230924
transform 1 0 1144 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_268
timestamp 1744230924
transform -1 0 1240 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_61
timestamp 1744230924
transform -1 0 1304 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_145
timestamp 1744230924
transform 1 0 1304 0 -1 1010
box -4 -6 52 206
use FILL  FILL_4_0_0
timestamp 1744230924
transform -1 0 1368 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_1
timestamp 1744230924
transform -1 0 1384 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_2
timestamp 1744230924
transform -1 0 1400 0 -1 1010
box -4 -6 20 206
use OAI21X1  OAI21X1_264
timestamp 1744230924
transform -1 0 1464 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_273
timestamp 1744230924
transform -1 0 1528 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_206
timestamp 1744230924
transform -1 0 1576 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_82
timestamp 1744230924
transform 1 0 1576 0 -1 1010
box -4 -6 196 206
use NOR2X1  NOR2X1_62
timestamp 1744230924
transform -1 0 1816 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_64
timestamp 1744230924
transform 1 0 1816 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_59
timestamp 1744230924
transform -1 0 1912 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_61
timestamp 1744230924
transform 1 0 1912 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_128
timestamp 1744230924
transform 1 0 1960 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_129
timestamp 1744230924
transform -1 0 2088 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_88
timestamp 1744230924
transform 1 0 2088 0 -1 1010
box -4 -6 36 206
use AOI22X1  AOI22X1_14
timestamp 1744230924
transform -1 0 2200 0 -1 1010
box -4 -6 84 206
use NAND2X1  NAND2X1_99
timestamp 1744230924
transform 1 0 2200 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_133
timestamp 1744230924
transform -1 0 2312 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_90
timestamp 1744230924
transform -1 0 2344 0 -1 1010
box -4 -6 36 206
use AOI22X1  AOI22X1_12
timestamp 1744230924
transform 1 0 2344 0 -1 1010
box -4 -6 84 206
use NOR2X1  NOR2X1_69
timestamp 1744230924
transform 1 0 2424 0 -1 1010
box -4 -6 52 206
use MUX2X1  MUX2X1_7
timestamp 1744230924
transform 1 0 2472 0 -1 1010
box -4 -6 100 206
use XNOR2X1  XNOR2X1_43
timestamp 1744230924
transform -1 0 2680 0 -1 1010
box -4 -6 116 206
use NAND2X1  NAND2X1_86
timestamp 1744230924
transform 1 0 2680 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_79
timestamp 1744230924
transform -1 0 2760 0 -1 1010
box -4 -6 36 206
use BUFX4  BUFX4_27
timestamp 1744230924
transform -1 0 2824 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_192
timestamp 1744230924
transform -1 0 2872 0 -1 1010
box -4 -6 52 206
use FILL  FILL_4_1_0
timestamp 1744230924
transform -1 0 2888 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_1
timestamp 1744230924
transform -1 0 2904 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_2
timestamp 1744230924
transform -1 0 2920 0 -1 1010
box -4 -6 20 206
use OAI21X1  OAI21X1_112
timestamp 1744230924
transform -1 0 2984 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_85
timestamp 1744230924
transform 1 0 2984 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_78
timestamp 1744230924
transform 1 0 3032 0 -1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_87
timestamp 1744230924
transform 1 0 3064 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_143
timestamp 1744230924
transform 1 0 3112 0 -1 1010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_90
timestamp 1744230924
transform 1 0 3304 0 -1 1010
box -4 -6 196 206
use BUFX4  BUFX4_12
timestamp 1744230924
transform 1 0 3496 0 -1 1010
box -4 -6 68 206
use OR2X2  OR2X2_7
timestamp 1744230924
transform 1 0 3560 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_72
timestamp 1744230924
transform -1 0 3672 0 -1 1010
box -4 -6 52 206
use XOR2X1  XOR2X1_6
timestamp 1744230924
transform -1 0 3784 0 -1 1010
box -4 -6 116 206
use NOR2X1  NOR2X1_43
timestamp 1744230924
transform 1 0 3784 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_91
timestamp 1744230924
transform 1 0 3832 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_15
timestamp 1744230924
transform 1 0 3896 0 -1 1010
box -4 -6 68 206
use AND2X2  AND2X2_4
timestamp 1744230924
transform 1 0 3960 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_89
timestamp 1744230924
transform 1 0 4024 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_74
timestamp 1744230924
transform -1 0 4136 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_4
timestamp 1744230924
transform -1 0 4184 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_174
timestamp 1744230924
transform -1 0 4248 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_175
timestamp 1744230924
transform -1 0 4312 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_145
timestamp 1744230924
transform 1 0 4312 0 -1 1010
box -4 -6 196 206
use FILL  FILL_4_2_0
timestamp 1744230924
transform -1 0 4520 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_2_1
timestamp 1744230924
transform -1 0 4536 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_2_2
timestamp 1744230924
transform -1 0 4552 0 -1 1010
box -4 -6 20 206
use XNOR2X1  XNOR2X1_58
timestamp 1744230924
transform -1 0 4664 0 -1 1010
box -4 -6 116 206
use XNOR2X1  XNOR2X1_38
timestamp 1744230924
transform 1 0 4664 0 -1 1010
box -4 -6 116 206
use INVX1  INVX1_76
timestamp 1744230924
transform 1 0 4776 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_13
timestamp 1744230924
transform 1 0 4808 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_148
timestamp 1744230924
transform 1 0 4872 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_93
timestamp 1744230924
transform 1 0 4920 0 -1 1010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_97
timestamp 1744230924
transform -1 0 5304 0 -1 1010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_102
timestamp 1744230924
transform 1 0 5304 0 -1 1010
box -4 -6 196 206
use INVX2  INVX2_23
timestamp 1744230924
transform -1 0 5528 0 -1 1010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_39
timestamp 1744230924
transform 1 0 5528 0 -1 1010
box -4 -6 196 206
use BUFX2  BUFX2_22
timestamp 1744230924
transform 1 0 5720 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_25
timestamp 1744230924
transform 1 0 5768 0 -1 1010
box -4 -6 52 206
use FILL  FILL_5_1
timestamp 1744230924
transform -1 0 5832 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_2
timestamp 1744230924
transform -1 0 5848 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_3
timestamp 1744230924
transform -1 0 5864 0 -1 1010
box -4 -6 20 206
use OAI21X1  OAI21X1_81
timestamp 1744230924
transform 1 0 8 0 1 1010
box -4 -6 68 206
use AOI22X1  AOI22X1_4
timestamp 1744230924
transform 1 0 72 0 1 1010
box -4 -6 84 206
use AOI21X1  AOI21X1_12
timestamp 1744230924
transform -1 0 216 0 1 1010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_32
timestamp 1744230924
transform 1 0 216 0 1 1010
box -4 -6 116 206
use NOR2X1  NOR2X1_149
timestamp 1744230924
transform 1 0 328 0 1 1010
box -4 -6 52 206
use INVX2  INVX2_4
timestamp 1744230924
transform 1 0 376 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_276
timestamp 1744230924
transform 1 0 408 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_148
timestamp 1744230924
transform 1 0 472 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_179
timestamp 1744230924
transform -1 0 552 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_277
timestamp 1744230924
transform -1 0 616 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_176
timestamp 1744230924
transform 1 0 616 0 1 1010
box -4 -6 36 206
use AOI21X1  AOI21X1_65
timestamp 1744230924
transform -1 0 712 0 1 1010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_98
timestamp 1744230924
transform -1 0 824 0 1 1010
box -4 -6 116 206
use AND2X2  AND2X2_12
timestamp 1744230924
transform 1 0 824 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_198
timestamp 1744230924
transform 1 0 888 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_140
timestamp 1744230924
transform 1 0 936 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_141
timestamp 1744230924
transform -1 0 1032 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_267
timestamp 1744230924
transform 1 0 1032 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_271
timestamp 1744230924
transform 1 0 1160 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_270
timestamp 1744230924
transform 1 0 1096 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_146
timestamp 1744230924
transform 1 0 1224 0 1 1010
box -4 -6 52 206
use AOI21X1  AOI21X1_62
timestamp 1744230924
transform 1 0 1304 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_175
timestamp 1744230924
transform 1 0 1272 0 1 1010
box -4 -6 36 206
use FILL  FILL_5_0_0
timestamp 1744230924
transform -1 0 1384 0 1 1010
box -4 -6 20 206
use NOR2X1  NOR2X1_144
timestamp 1744230924
transform 1 0 1448 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_173
timestamp 1744230924
transform -1 0 1448 0 1 1010
box -4 -6 36 206
use FILL  FILL_5_0_2
timestamp 1744230924
transform -1 0 1416 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_1
timestamp 1744230924
transform -1 0 1400 0 1 1010
box -4 -6 20 206
use XOR2X1  XOR2X1_30
timestamp 1744230924
transform 1 0 1496 0 1 1010
box -4 -6 116 206
use INVX1  INVX1_172
timestamp 1744230924
transform -1 0 1640 0 1 1010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_81
timestamp 1744230924
transform 1 0 1640 0 1 1010
box -4 -6 196 206
use INVX4  INVX4_6
timestamp 1744230924
transform 1 0 1832 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_93
timestamp 1744230924
transform 1 0 1880 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_86
timestamp 1744230924
transform 1 0 1928 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_124
timestamp 1744230924
transform -1 0 2024 0 1 1010
box -4 -6 68 206
use AOI22X1  AOI22X1_13
timestamp 1744230924
transform 1 0 2024 0 1 1010
box -4 -6 84 206
use NAND2X1  NAND2X1_98
timestamp 1744230924
transform -1 0 2152 0 1 1010
box -4 -6 52 206
use AOI21X1  AOI21X1_20
timestamp 1744230924
transform -1 0 2216 0 1 1010
box -4 -6 68 206
use AOI22X1  AOI22X1_11
timestamp 1744230924
transform 1 0 2216 0 1 1010
box -4 -6 84 206
use OAI21X1  OAI21X1_126
timestamp 1744230924
transform -1 0 2360 0 1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_6
timestamp 1744230924
transform -1 0 2456 0 1 1010
box -4 -6 100 206
use XOR2X1  XOR2X1_13
timestamp 1744230924
transform -1 0 2568 0 1 1010
box -4 -6 116 206
use INVX1  INVX1_84
timestamp 1744230924
transform 1 0 2568 0 1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_97
timestamp 1744230924
transform -1 0 2648 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_125
timestamp 1744230924
transform -1 0 2712 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_91
timestamp 1744230924
transform 1 0 2712 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_117
timestamp 1744230924
transform 1 0 2760 0 1 1010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_42
timestamp 1744230924
transform -1 0 2936 0 1 1010
box -4 -6 116 206
use FILL  FILL_5_1_0
timestamp 1744230924
transform 1 0 2936 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_1
timestamp 1744230924
transform 1 0 2952 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_2
timestamp 1744230924
transform 1 0 2968 0 1 1010
box -4 -6 20 206
use INVX4  INVX4_3
timestamp 1744230924
transform 1 0 2984 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_9
timestamp 1744230924
transform 1 0 3032 0 1 1010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_138
timestamp 1744230924
transform 1 0 3080 0 1 1010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_141
timestamp 1744230924
transform 1 0 3272 0 1 1010
box -4 -6 196 206
use BUFX4  BUFX4_14
timestamp 1744230924
transform -1 0 3528 0 1 1010
box -4 -6 68 206
use BUFX4  BUFX4_15
timestamp 1744230924
transform 1 0 3528 0 1 1010
box -4 -6 68 206
use BUFX4  BUFX4_13
timestamp 1744230924
transform 1 0 3592 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_94
timestamp 1744230924
transform 1 0 3656 0 1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_2
timestamp 1744230924
transform -1 0 3816 0 1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_95
timestamp 1744230924
transform -1 0 3880 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_93
timestamp 1744230924
transform 1 0 3880 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_71
timestamp 1744230924
transform -1 0 3992 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_44
timestamp 1744230924
transform 1 0 3992 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_64
timestamp 1744230924
transform -1 0 4072 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_90
timestamp 1744230924
transform 1 0 4072 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_92
timestamp 1744230924
transform -1 0 4200 0 1 1010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_35
timestamp 1744230924
transform -1 0 4312 0 1 1010
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_148
timestamp 1744230924
transform 1 0 4312 0 1 1010
box -4 -6 196 206
use FILL  FILL_5_2_0
timestamp 1744230924
transform -1 0 4520 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_2_1
timestamp 1744230924
transform -1 0 4536 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_2_2
timestamp 1744230924
transform -1 0 4552 0 1 1010
box -4 -6 20 206
use INVX4  INVX4_5
timestamp 1744230924
transform -1 0 4600 0 1 1010
box -4 -6 52 206
use INVX2  INVX2_8
timestamp 1744230924
transform -1 0 4632 0 1 1010
box -4 -6 36 206
use BUFX2  BUFX2_3
timestamp 1744230924
transform -1 0 4680 0 1 1010
box -4 -6 52 206
use XOR2X1  XOR2X1_17
timestamp 1744230924
transform -1 0 4792 0 1 1010
box -4 -6 116 206
use INVX4  INVX4_2
timestamp 1744230924
transform 1 0 4792 0 1 1010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_92
timestamp 1744230924
transform 1 0 4840 0 1 1010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_91
timestamp 1744230924
transform 1 0 5032 0 1 1010
box -4 -6 196 206
use XNOR2X1  XNOR2X1_68
timestamp 1744230924
transform 1 0 5224 0 1 1010
box -4 -6 116 206
use XNOR2X1  XNOR2X1_70
timestamp 1744230924
transform 1 0 5336 0 1 1010
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_101
timestamp 1744230924
transform 1 0 5448 0 1 1010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_38
timestamp 1744230924
transform 1 0 5640 0 1 1010
box -4 -6 196 206
use FILL  FILL_6_1
timestamp 1744230924
transform 1 0 5832 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_2
timestamp 1744230924
transform 1 0 5848 0 1 1010
box -4 -6 20 206
use INVX1  INVX1_49
timestamp 1744230924
transform 1 0 8 0 -1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_32
timestamp 1744230924
transform -1 0 88 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_80
timestamp 1744230924
transform 1 0 88 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_41
timestamp 1744230924
transform 1 0 152 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_42
timestamp 1744230924
transform 1 0 200 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_35
timestamp 1744230924
transform -1 0 296 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_34
timestamp 1744230924
transform -1 0 344 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_48
timestamp 1744230924
transform 1 0 344 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_54
timestamp 1744230924
transform 1 0 376 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_55
timestamp 1744230924
transform -1 0 472 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_53
timestamp 1744230924
transform 1 0 472 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_69
timestamp 1744230924
transform 1 0 520 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_57
timestamp 1744230924
transform 1 0 584 0 -1 1410
box -4 -6 52 206
use INVX2  INVX2_27
timestamp 1744230924
transform -1 0 664 0 -1 1410
box -4 -6 36 206
use MUX2X1  MUX2X1_12
timestamp 1744230924
transform -1 0 760 0 -1 1410
box -4 -6 100 206
use OAI21X1  OAI21X1_278
timestamp 1744230924
transform 1 0 760 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_279
timestamp 1744230924
transform -1 0 888 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_180
timestamp 1744230924
transform -1 0 920 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_274
timestamp 1744230924
transform 1 0 920 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_275
timestamp 1744230924
transform -1 0 1048 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_203
timestamp 1744230924
transform -1 0 1096 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_269
timestamp 1744230924
transform -1 0 1160 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_205
timestamp 1744230924
transform 1 0 1160 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_272
timestamp 1744230924
transform -1 0 1272 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_204
timestamp 1744230924
transform -1 0 1320 0 -1 1410
box -4 -6 52 206
use FILL  FILL_6_0_0
timestamp 1744230924
transform -1 0 1336 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_1
timestamp 1744230924
transform -1 0 1352 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_2
timestamp 1744230924
transform -1 0 1368 0 -1 1410
box -4 -6 20 206
use XNOR2X1  XNOR2X1_96
timestamp 1744230924
transform -1 0 1480 0 -1 1410
box -4 -6 116 206
use XNOR2X1  XNOR2X1_95
timestamp 1744230924
transform 1 0 1480 0 -1 1410
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_80
timestamp 1744230924
transform 1 0 1592 0 -1 1410
box -4 -6 196 206
use NAND2X1  NAND2X1_94
timestamp 1744230924
transform 1 0 1784 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_95
timestamp 1744230924
transform 1 0 1832 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_85
timestamp 1744230924
transform 1 0 1880 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_123
timestamp 1744230924
transform 1 0 1912 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_96
timestamp 1744230924
transform 1 0 1976 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_70
timestamp 1744230924
transform -1 0 2072 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_120
timestamp 1744230924
transform -1 0 2136 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_121
timestamp 1744230924
transform 1 0 2136 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_122
timestamp 1744230924
transform -1 0 2264 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_118
timestamp 1744230924
transform 1 0 2264 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_119
timestamp 1744230924
transform 1 0 2328 0 -1 1410
box -4 -6 68 206
use MUX2X1  MUX2X1_5
timestamp 1744230924
transform -1 0 2488 0 -1 1410
box -4 -6 100 206
use AOI21X1  AOI21X1_19
timestamp 1744230924
transform 1 0 2488 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_58
timestamp 1744230924
transform 1 0 2552 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_81
timestamp 1744230924
transform 1 0 2600 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_115
timestamp 1744230924
transform 1 0 2632 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_114
timestamp 1744230924
transform 1 0 2696 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_90
timestamp 1744230924
transform -1 0 2808 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_80
timestamp 1744230924
transform 1 0 2808 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_113
timestamp 1744230924
transform 1 0 2840 0 -1 1410
box -4 -6 68 206
use FILL  FILL_6_1_0
timestamp 1744230924
transform -1 0 2920 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_1
timestamp 1744230924
transform -1 0 2936 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_2
timestamp 1744230924
transform -1 0 2952 0 -1 1410
box -4 -6 20 206
use XOR2X1  XOR2X1_10
timestamp 1744230924
transform -1 0 3064 0 -1 1410
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_142
timestamp 1744230924
transform 1 0 3064 0 -1 1410
box -4 -6 196 206
use XOR2X1  XOR2X1_7
timestamp 1744230924
transform -1 0 3368 0 -1 1410
box -4 -6 116 206
use XOR2X1  XOR2X1_8
timestamp 1744230924
transform -1 0 3480 0 -1 1410
box -4 -6 116 206
use XNOR2X1  XNOR2X1_33
timestamp 1744230924
transform 1 0 3480 0 -1 1410
box -4 -6 116 206
use NAND2X1  NAND2X1_77
timestamp 1744230924
transform 1 0 3592 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_78
timestamp 1744230924
transform 1 0 3640 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_68
timestamp 1744230924
transform 1 0 3688 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_76
timestamp 1744230924
transform -1 0 3768 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_65
timestamp 1744230924
transform 1 0 3768 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_75
timestamp 1744230924
transform -1 0 3848 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_81
timestamp 1744230924
transform -1 0 3896 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_79
timestamp 1744230924
transform 1 0 3896 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_56
timestamp 1744230924
transform -1 0 3992 0 -1 1410
box -4 -6 52 206
use AOI22X1  AOI22X1_9
timestamp 1744230924
transform -1 0 4072 0 -1 1410
box -4 -6 84 206
use AOI22X1  AOI22X1_7
timestamp 1744230924
transform 1 0 4072 0 -1 1410
box -4 -6 84 206
use NOR2X1  NOR2X1_51
timestamp 1744230924
transform -1 0 4200 0 -1 1410
box -4 -6 52 206
use XNOR2X1  XNOR2X1_34
timestamp 1744230924
transform -1 0 4312 0 -1 1410
box -4 -6 116 206
use OAI21X1  OAI21X1_109
timestamp 1744230924
transform -1 0 4376 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_52
timestamp 1744230924
transform 1 0 4376 0 -1 1410
box -4 -6 52 206
use FILL  FILL_6_2_0
timestamp 1744230924
transform 1 0 4424 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_2_1
timestamp 1744230924
transform 1 0 4440 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_2_2
timestamp 1744230924
transform 1 0 4456 0 -1 1410
box -4 -6 20 206
use NOR2X1  NOR2X1_54
timestamp 1744230924
transform 1 0 4472 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_53
timestamp 1744230924
transform 1 0 4520 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_105
timestamp 1744230924
transform 1 0 4568 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_73
timestamp 1744230924
transform 1 0 4632 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_106
timestamp 1744230924
transform 1 0 4664 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_7
timestamp 1744230924
transform 1 0 4728 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_98
timestamp 1744230924
transform -1 0 4984 0 -1 1410
box -4 -6 196 206
use CLKBUF1  CLKBUF1_7
timestamp 1744230924
transform 1 0 4984 0 -1 1410
box -4 -6 148 206
use NAND2X1  NAND2X1_154
timestamp 1744230924
transform 1 0 5128 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_155
timestamp 1744230924
transform 1 0 5176 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_153
timestamp 1744230924
transform 1 0 5224 0 -1 1410
box -4 -6 52 206
use INVX4  INVX4_8
timestamp 1744230924
transform 1 0 5272 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_158
timestamp 1744230924
transform 1 0 5320 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_136
timestamp 1744230924
transform -1 0 5400 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_160
timestamp 1744230924
transform -1 0 5448 0 -1 1410
box -4 -6 52 206
use OR2X2  OR2X2_13
timestamp 1744230924
transform -1 0 5512 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_38
timestamp 1744230924
transform -1 0 5560 0 -1 1410
box -4 -6 52 206
use XOR2X1  XOR2X1_20
timestamp 1744230924
transform -1 0 5672 0 -1 1410
box -4 -6 116 206
use XOR2X1  XOR2X1_21
timestamp 1744230924
transform -1 0 5784 0 -1 1410
box -4 -6 116 206
use BUFX2  BUFX2_48
timestamp 1744230924
transform 1 0 5784 0 -1 1410
box -4 -6 52 206
use FILL  FILL_7_1
timestamp 1744230924
transform -1 0 5848 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_2
timestamp 1744230924
transform -1 0 5864 0 -1 1410
box -4 -6 20 206
use AND2X2  AND2X2_3
timestamp 1744230924
transform 1 0 8 0 1 1410
box -4 -6 68 206
use OR2X2  OR2X2_6
timestamp 1744230924
transform 1 0 72 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_71
timestamp 1744230924
transform 1 0 136 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_10
timestamp 1744230924
transform -1 0 264 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_9
timestamp 1744230924
transform -1 0 328 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_72
timestamp 1744230924
transform -1 0 392 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_67
timestamp 1744230924
transform 1 0 392 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_52
timestamp 1744230924
transform 1 0 456 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_56
timestamp 1744230924
transform 1 0 504 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_68
timestamp 1744230924
transform 1 0 552 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_70
timestamp 1744230924
transform 1 0 616 0 1 1410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_27
timestamp 1744230924
transform -1 0 792 0 1 1410
box -4 -6 116 206
use AOI22X1  AOI22X1_32
timestamp 1744230924
transform 1 0 792 0 1 1410
box -4 -6 84 206
use AOI22X1  AOI22X1_33
timestamp 1744230924
transform 1 0 872 0 1 1410
box -4 -6 84 206
use INVX1  INVX1_178
timestamp 1744230924
transform -1 0 984 0 1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_150
timestamp 1744230924
transform 1 0 984 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_208
timestamp 1744230924
transform -1 0 1080 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_177
timestamp 1744230924
transform -1 0 1112 0 1 1410
box -4 -6 36 206
use XNOR2X1  XNOR2X1_94
timestamp 1744230924
transform -1 0 1224 0 1 1410
box -4 -6 116 206
use AOI21X1  AOI21X1_63
timestamp 1744230924
transform 1 0 1224 0 1 1410
box -4 -6 68 206
use AOI22X1  AOI22X1_31
timestamp 1744230924
transform 1 0 1288 0 1 1410
box -4 -6 84 206
use FILL  FILL_7_0_0
timestamp 1744230924
transform -1 0 1384 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_1
timestamp 1744230924
transform -1 0 1400 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_2
timestamp 1744230924
transform -1 0 1416 0 1 1410
box -4 -6 20 206
use XNOR2X1  XNOR2X1_97
timestamp 1744230924
transform -1 0 1528 0 1 1410
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_132
timestamp 1744230924
transform 1 0 1528 0 1 1410
box -4 -6 196 206
use CLKBUF1  CLKBUF1_1
timestamp 1744230924
transform -1 0 1864 0 1 1410
box -4 -6 148 206
use XNOR2X1  XNOR2X1_39
timestamp 1744230924
transform 1 0 1864 0 1 1410
box -4 -6 116 206
use XOR2X1  XOR2X1_12
timestamp 1744230924
transform 1 0 1976 0 1 1410
box -4 -6 116 206
use NAND2X1  NAND2X1_92
timestamp 1744230924
transform -1 0 2136 0 1 1410
box -4 -6 52 206
use XOR2X1  XOR2X1_11
timestamp 1744230924
transform -1 0 2248 0 1 1410
box -4 -6 116 206
use NOR2X1  NOR2X1_65
timestamp 1744230924
transform -1 0 2296 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_82
timestamp 1744230924
transform -1 0 2328 0 1 1410
box -4 -6 36 206
use XNOR2X1  XNOR2X1_41
timestamp 1744230924
transform -1 0 2440 0 1 1410
box -4 -6 116 206
use OR2X2  OR2X2_8
timestamp 1744230924
transform 1 0 2440 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_89
timestamp 1744230924
transform -1 0 2552 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_88
timestamp 1744230924
transform -1 0 2600 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_57
timestamp 1744230924
transform 1 0 2600 0 1 1410
box -4 -6 52 206
use AND2X2  AND2X2_5
timestamp 1744230924
transform 1 0 2648 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_116
timestamp 1744230924
transform -1 0 2776 0 1 1410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_40
timestamp 1744230924
transform -1 0 2888 0 1 1410
box -4 -6 116 206
use FILL  FILL_7_1_0
timestamp 1744230924
transform 1 0 2888 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_1
timestamp 1744230924
transform 1 0 2904 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_2
timestamp 1744230924
transform 1 0 2920 0 1 1410
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_140
timestamp 1744230924
transform 1 0 2936 0 1 1410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_139
timestamp 1744230924
transform 1 0 3128 0 1 1410
box -4 -6 196 206
use CLKBUF1  CLKBUF1_5
timestamp 1744230924
transform 1 0 3320 0 1 1410
box -4 -6 148 206
use OAI21X1  OAI21X1_98
timestamp 1744230924
transform 1 0 3464 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_99
timestamp 1744230924
transform -1 0 3592 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_69
timestamp 1744230924
transform -1 0 3624 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_96
timestamp 1744230924
transform 1 0 3624 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_102
timestamp 1744230924
transform 1 0 3688 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_103
timestamp 1744230924
transform 1 0 3752 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_104
timestamp 1744230924
transform -1 0 3880 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_97
timestamp 1744230924
transform -1 0 3944 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_72
timestamp 1744230924
transform 1 0 3944 0 1 1410
box -4 -6 36 206
use AOI22X1  AOI22X1_10
timestamp 1744230924
transform -1 0 4056 0 1 1410
box -4 -6 84 206
use AOI22X1  AOI22X1_8
timestamp 1744230924
transform 1 0 4056 0 1 1410
box -4 -6 84 206
use MUX2X1  MUX2X1_4
timestamp 1744230924
transform 1 0 4136 0 1 1410
box -4 -6 100 206
use AOI21X1  AOI21X1_18
timestamp 1744230924
transform 1 0 4232 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_77
timestamp 1744230924
transform -1 0 4328 0 1 1410
box -4 -6 36 206
use INVX1  INVX1_75
timestamp 1744230924
transform 1 0 4328 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_110
timestamp 1744230924
transform -1 0 4424 0 1 1410
box -4 -6 68 206
use FILL  FILL_7_2_0
timestamp 1744230924
transform -1 0 4440 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_2_1
timestamp 1744230924
transform -1 0 4456 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_2_2
timestamp 1744230924
transform -1 0 4472 0 1 1410
box -4 -6 20 206
use INVX1  INVX1_71
timestamp 1744230924
transform -1 0 4504 0 1 1410
box -4 -6 36 206
use AOI21X1  AOI21X1_17
timestamp 1744230924
transform 1 0 4504 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_111
timestamp 1744230924
transform 1 0 4568 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_84
timestamp 1744230924
transform -1 0 4680 0 1 1410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_152
timestamp 1744230924
transform 1 0 4680 0 1 1410
box -4 -6 196 206
use CLKBUF1  CLKBUF1_10
timestamp 1744230924
transform -1 0 5016 0 1 1410
box -4 -6 148 206
use NAND2X1  NAND2X1_156
timestamp 1744230924
transform -1 0 5064 0 1 1410
box -4 -6 52 206
use AOI22X1  AOI22X1_23
timestamp 1744230924
transform -1 0 5144 0 1 1410
box -4 -6 84 206
use OAI21X1  OAI21X1_201
timestamp 1744230924
transform 1 0 5144 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_159
timestamp 1744230924
transform 1 0 5208 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_202
timestamp 1744230924
transform 1 0 5256 0 1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_115
timestamp 1744230924
transform 1 0 5320 0 1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_15
timestamp 1744230924
transform -1 0 5432 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_161
timestamp 1744230924
transform 1 0 5432 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_113
timestamp 1744230924
transform -1 0 5528 0 1 1410
box -4 -6 52 206
use XNOR2X1  XNOR2X1_71
timestamp 1744230924
transform 1 0 5528 0 1 1410
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_42
timestamp 1744230924
transform 1 0 5640 0 1 1410
box -4 -6 196 206
use FILL  FILL_8_1
timestamp 1744230924
transform 1 0 5832 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_2
timestamp 1744230924
transform 1 0 5848 0 1 1410
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_124
timestamp 1744230924
transform -1 0 200 0 -1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_76
timestamp 1744230924
transform -1 0 264 0 -1 1810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_25
timestamp 1744230924
transform -1 0 376 0 -1 1810
box -4 -6 116 206
use XNOR2X1  XNOR2X1_26
timestamp 1744230924
transform -1 0 488 0 -1 1810
box -4 -6 116 206
use OAI21X1  OAI21X1_65
timestamp 1744230924
transform -1 0 552 0 -1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_8
timestamp 1744230924
transform -1 0 616 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_66
timestamp 1744230924
transform -1 0 680 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_47
timestamp 1744230924
transform -1 0 712 0 -1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_31
timestamp 1744230924
transform 1 0 712 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_64
timestamp 1744230924
transform 1 0 760 0 -1 1810
box -4 -6 68 206
use XOR2X1  XOR2X1_5
timestamp 1744230924
transform -1 0 936 0 -1 1810
box -4 -6 116 206
use XOR2X1  XOR2X1_31
timestamp 1744230924
transform 1 0 936 0 -1 1810
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_130
timestamp 1744230924
transform 1 0 1048 0 -1 1810
box -4 -6 196 206
use NAND2X1  NAND2X1_48
timestamp 1744230924
transform 1 0 1240 0 -1 1810
box -4 -6 52 206
use FILL  FILL_8_0_0
timestamp 1744230924
transform 1 0 1288 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_1
timestamp 1744230924
transform 1 0 1304 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_2
timestamp 1744230924
transform 1 0 1320 0 -1 1810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_131
timestamp 1744230924
transform 1 0 1336 0 -1 1810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_129
timestamp 1744230924
transform 1 0 1528 0 -1 1810
box -4 -6 196 206
use XNOR2X1  XNOR2X1_10
timestamp 1744230924
transform -1 0 1832 0 -1 1810
box -4 -6 116 206
use OAI21X1  OAI21X1_25
timestamp 1744230924
transform 1 0 1832 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_20
timestamp 1744230924
transform 1 0 1896 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_26
timestamp 1744230924
transform 1 0 1944 0 -1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_2
timestamp 1744230924
transform -1 0 2072 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_20
timestamp 1744230924
transform -1 0 2104 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_27
timestamp 1744230924
transform 1 0 2104 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_28
timestamp 1744230924
transform -1 0 2232 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_21
timestamp 1744230924
transform 1 0 2232 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_22
timestamp 1744230924
transform 1 0 2280 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_26
timestamp 1744230924
transform 1 0 2328 0 -1 1810
box -4 -6 196 206
use CLKBUF1  CLKBUF1_3
timestamp 1744230924
transform 1 0 2520 0 -1 1810
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_25
timestamp 1744230924
transform 1 0 2664 0 -1 1810
box -4 -6 196 206
use FILL  FILL_8_1_0
timestamp 1744230924
transform 1 0 2856 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_1
timestamp 1744230924
transform 1 0 2872 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_2
timestamp 1744230924
transform 1 0 2888 0 -1 1810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_24
timestamp 1744230924
transform 1 0 2904 0 -1 1810
box -4 -6 196 206
use NAND2X1  NAND2X1_10
timestamp 1744230924
transform -1 0 3144 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_11
timestamp 1744230924
transform 1 0 3144 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_11
timestamp 1744230924
transform 1 0 3208 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_12
timestamp 1744230924
transform -1 0 3320 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_10
timestamp 1744230924
transform -1 0 3384 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_11
timestamp 1744230924
transform -1 0 3416 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_13
timestamp 1744230924
transform 1 0 3416 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_12
timestamp 1744230924
transform 1 0 3480 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_45
timestamp 1744230924
transform -1 0 3576 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_47
timestamp 1744230924
transform 1 0 3576 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_66
timestamp 1744230924
transform -1 0 3656 0 -1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_46
timestamp 1744230924
transform -1 0 3704 0 -1 1810
box -4 -6 52 206
use AOI21X1  AOI21X1_16
timestamp 1744230924
transform -1 0 3768 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_48
timestamp 1744230924
transform 1 0 3768 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_82
timestamp 1744230924
transform 1 0 3816 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_107
timestamp 1744230924
transform 1 0 3864 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_70
timestamp 1744230924
transform 1 0 3928 0 -1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_83
timestamp 1744230924
transform 1 0 3960 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_108
timestamp 1744230924
transform -1 0 4072 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_74
timestamp 1744230924
transform -1 0 4104 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_100
timestamp 1744230924
transform 1 0 4104 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_80
timestamp 1744230924
transform -1 0 4216 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_146
timestamp 1744230924
transform 1 0 4216 0 -1 1810
box -4 -6 196 206
use FILL  FILL_8_2_0
timestamp 1744230924
transform 1 0 4408 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_2_1
timestamp 1744230924
transform 1 0 4424 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_2_2
timestamp 1744230924
transform 1 0 4440 0 -1 1810
box -4 -6 20 206
use XNOR2X1  XNOR2X1_37
timestamp 1744230924
transform 1 0 4456 0 -1 1810
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_151
timestamp 1744230924
transform 1 0 4568 0 -1 1810
box -4 -6 196 206
use INVX2  INVX2_2
timestamp 1744230924
transform -1 0 4792 0 -1 1810
box -4 -6 36 206
use XNOR2X1  XNOR2X1_15
timestamp 1744230924
transform 1 0 4792 0 -1 1810
box -4 -6 116 206
use INVX2  INVX2_21
timestamp 1744230924
transform 1 0 4904 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_205
timestamp 1744230924
transform 1 0 4936 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_206
timestamp 1744230924
transform -1 0 5064 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_163
timestamp 1744230924
transform 1 0 5064 0 -1 1810
box -4 -6 52 206
use AOI22X1  AOI22X1_24
timestamp 1744230924
transform -1 0 5192 0 -1 1810
box -4 -6 84 206
use OAI21X1  OAI21X1_203
timestamp 1744230924
transform -1 0 5256 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_116
timestamp 1744230924
transform -1 0 5304 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_162
timestamp 1744230924
transform -1 0 5352 0 -1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_16
timestamp 1744230924
transform -1 0 5416 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_117
timestamp 1744230924
transform 1 0 5416 0 -1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_14
timestamp 1744230924
transform 1 0 5464 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_112
timestamp 1744230924
transform -1 0 5576 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_40
timestamp 1744230924
transform 1 0 5576 0 -1 1810
box -4 -6 196 206
use BUFX2  BUFX2_23
timestamp 1744230924
transform 1 0 5768 0 -1 1810
box -4 -6 52 206
use FILL  FILL_9_1
timestamp 1744230924
transform -1 0 5832 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_2
timestamp 1744230924
transform -1 0 5848 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_3
timestamp 1744230924
transform -1 0 5864 0 -1 1810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_74
timestamp 1744230924
transform 1 0 8 0 1 1810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_73
timestamp 1744230924
transform 1 0 200 0 1 1810
box -4 -6 196 206
use NAND2X1  NAND2X1_65
timestamp 1744230924
transform -1 0 440 0 1 1810
box -4 -6 52 206
use OR2X2  OR2X2_5
timestamp 1744230924
transform 1 0 440 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_33
timestamp 1744230924
transform 1 0 504 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_50
timestamp 1744230924
transform -1 0 600 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_49
timestamp 1744230924
transform -1 0 648 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_75
timestamp 1744230924
transform -1 0 712 0 1 1810
box -4 -6 68 206
use AND2X2  AND2X2_2
timestamp 1744230924
transform 1 0 712 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_57
timestamp 1744230924
transform 1 0 776 0 1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_207
timestamp 1744230924
transform -1 0 856 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_44
timestamp 1744230924
transform -1 0 888 0 1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_51
timestamp 1744230924
transform -1 0 936 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_46
timestamp 1744230924
transform 1 0 936 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_63
timestamp 1744230924
transform 1 0 968 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_62
timestamp 1744230924
transform -1 0 1096 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_46
timestamp 1744230924
transform -1 0 1144 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_45
timestamp 1744230924
transform 1 0 1144 0 1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_47
timestamp 1744230924
transform -1 0 1224 0 1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_68
timestamp 1744230924
transform 1 0 1224 0 1 1810
box -4 -6 196 206
use FILL  FILL_9_0_0
timestamp 1744230924
transform 1 0 1416 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_1
timestamp 1744230924
transform 1 0 1432 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_2
timestamp 1744230924
transform 1 0 1448 0 1 1810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_70
timestamp 1744230924
transform 1 0 1464 0 1 1810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_17
timestamp 1744230924
transform 1 0 1656 0 1 1810
box -4 -6 196 206
use INVX1  INVX1_21
timestamp 1744230924
transform 1 0 1848 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_21
timestamp 1744230924
transform -1 0 1944 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_19
timestamp 1744230924
transform -1 0 1992 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_23
timestamp 1744230924
transform -1 0 2056 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_18
timestamp 1744230924
transform -1 0 2104 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_19
timestamp 1744230924
transform -1 0 2136 0 1 1810
box -4 -6 36 206
use XNOR2X1  XNOR2X1_9
timestamp 1744230924
transform -1 0 2248 0 1 1810
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_22
timestamp 1744230924
transform 1 0 2248 0 1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_7
timestamp 1744230924
transform -1 0 2504 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_10
timestamp 1744230924
transform 1 0 2504 0 1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_7
timestamp 1744230924
transform -1 0 2584 0 1 1810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_1
timestamp 1744230924
transform 1 0 2584 0 1 1810
box -4 -6 116 206
use NAND2X1  NAND2X1_5
timestamp 1744230924
transform 1 0 2696 0 1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_23
timestamp 1744230924
transform 1 0 2744 0 1 1810
box -4 -6 196 206
use FILL  FILL_9_1_0
timestamp 1744230924
transform 1 0 2936 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_1
timestamp 1744230924
transform 1 0 2952 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_2
timestamp 1744230924
transform 1 0 2968 0 1 1810
box -4 -6 20 206
use NAND2X1  NAND2X1_6
timestamp 1744230924
transform 1 0 2984 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_7
timestamp 1744230924
transform -1 0 3080 0 1 1810
box -4 -6 52 206
use INVX2  INVX2_1
timestamp 1744230924
transform -1 0 3112 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_8
timestamp 1744230924
transform -1 0 3176 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_8
timestamp 1744230924
transform 1 0 3176 0 1 1810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_2
timestamp 1744230924
transform 1 0 3224 0 1 1810
box -4 -6 116 206
use OAI21X1  OAI21X1_9
timestamp 1744230924
transform 1 0 3336 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_9
timestamp 1744230924
transform 1 0 3400 0 1 1810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_3
timestamp 1744230924
transform -1 0 3560 0 1 1810
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_34
timestamp 1744230924
transform 1 0 3560 0 1 1810
box -4 -6 196 206
use MUX2X1  MUX2X1_3
timestamp 1744230924
transform 1 0 3752 0 1 1810
box -4 -6 100 206
use OAI21X1  OAI21X1_101
timestamp 1744230924
transform -1 0 3912 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_50
timestamp 1744230924
transform 1 0 3912 0 1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_49
timestamp 1744230924
transform -1 0 4008 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_67
timestamp 1744230924
transform 1 0 4008 0 1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_55
timestamp 1744230924
transform 1 0 4040 0 1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_33
timestamp 1744230924
transform -1 0 4280 0 1 1810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_147
timestamp 1744230924
transform 1 0 4280 0 1 1810
box -4 -6 196 206
use FILL  FILL_9_2_0
timestamp 1744230924
transform 1 0 4472 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_2_1
timestamp 1744230924
transform 1 0 4488 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_2_2
timestamp 1744230924
transform 1 0 4504 0 1 1810
box -4 -6 20 206
use AOI21X1  AOI21X1_3
timestamp 1744230924
transform 1 0 4520 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_36
timestamp 1744230924
transform -1 0 4648 0 1 1810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_12
timestamp 1744230924
transform 1 0 4648 0 1 1810
box -4 -6 116 206
use OAI21X1  OAI21X1_43
timestamp 1744230924
transform 1 0 4760 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_30
timestamp 1744230924
transform -1 0 4856 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_44
timestamp 1744230924
transform 1 0 4856 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_5
timestamp 1744230924
transform 1 0 4920 0 1 1810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_16
timestamp 1744230924
transform -1 0 5096 0 1 1810
box -4 -6 116 206
use INVX1  INVX1_135
timestamp 1744230924
transform 1 0 5096 0 1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_111
timestamp 1744230924
transform 1 0 5128 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_157
timestamp 1744230924
transform -1 0 5224 0 1 1810
box -4 -6 52 206
use INVX4  INVX4_4
timestamp 1744230924
transform -1 0 5272 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_152
timestamp 1744230924
transform -1 0 5320 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_134
timestamp 1744230924
transform 1 0 5320 0 1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_149
timestamp 1744230924
transform 1 0 5352 0 1 1810
box -4 -6 52 206
use INVX2  INVX2_22
timestamp 1744230924
transform -1 0 5432 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_204
timestamp 1744230924
transform 1 0 5432 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_114
timestamp 1744230924
transform -1 0 5544 0 1 1810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_69
timestamp 1744230924
transform -1 0 5656 0 1 1810
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_103
timestamp 1744230924
transform 1 0 5656 0 1 1810
box -4 -6 196 206
use FILL  FILL_10_1
timestamp 1744230924
transform 1 0 5848 0 1 1810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_123
timestamp 1744230924
transform 1 0 8 0 -1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_72
timestamp 1744230924
transform 1 0 200 0 -1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_122
timestamp 1744230924
transform -1 0 584 0 -1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_71
timestamp 1744230924
transform 1 0 584 0 -1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_128
timestamp 1744230924
transform -1 0 968 0 -1 2210
box -4 -6 196 206
use CLKBUF1  CLKBUF1_6
timestamp 1744230924
transform -1 0 1112 0 -1 2210
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_67
timestamp 1744230924
transform -1 0 1304 0 -1 2210
box -4 -6 196 206
use FILL  FILL_10_0_0
timestamp 1744230924
transform 1 0 1304 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_0_1
timestamp 1744230924
transform 1 0 1320 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_0_2
timestamp 1744230924
transform 1 0 1336 0 -1 2210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_16
timestamp 1744230924
transform 1 0 1352 0 -1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_15
timestamp 1744230924
transform 1 0 1544 0 -1 2210
box -4 -6 196 206
use INVX1  INVX1_18
timestamp 1744230924
transform 1 0 1736 0 -1 2210
box -4 -6 36 206
use NOR2X1  NOR2X1_14
timestamp 1744230924
transform 1 0 1768 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_22
timestamp 1744230924
transform 1 0 1816 0 -1 2210
box -4 -6 68 206
use NOR2X1  NOR2X1_13
timestamp 1744230924
transform 1 0 1880 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_17
timestamp 1744230924
transform 1 0 1928 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_24
timestamp 1744230924
transform 1 0 1960 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_21
timestamp 1744230924
transform 1 0 2024 0 -1 2210
box -4 -6 196 206
use NOR2X1  NOR2X1_5
timestamp 1744230924
transform -1 0 2264 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_9
timestamp 1744230924
transform 1 0 2264 0 -1 2210
box -4 -6 36 206
use NOR2X1  NOR2X1_6
timestamp 1744230924
transform 1 0 2296 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_5
timestamp 1744230924
transform 1 0 2344 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_6
timestamp 1744230924
transform 1 0 2408 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_4
timestamp 1744230924
transform 1 0 2472 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_29
timestamp 1744230924
transform 1 0 2536 0 -1 2210
box -4 -6 196 206
use INVX1  INVX1_1
timestamp 1744230924
transform 1 0 2728 0 -1 2210
box -4 -6 36 206
use NOR2X1  NOR2X1_1
timestamp 1744230924
transform 1 0 2760 0 -1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_1
timestamp 1744230924
transform 1 0 2808 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_2
timestamp 1744230924
transform -1 0 2888 0 -1 2210
box -4 -6 36 206
use FILL  FILL_10_1_0
timestamp 1744230924
transform 1 0 2888 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_1_1
timestamp 1744230924
transform 1 0 2904 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_1_2
timestamp 1744230924
transform 1 0 2920 0 -1 2210
box -4 -6 20 206
use NOR2X1  NOR2X1_2
timestamp 1744230924
transform 1 0 2936 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_27
timestamp 1744230924
transform -1 0 3176 0 -1 2210
box -4 -6 196 206
use BUFX2  BUFX2_10
timestamp 1744230924
transform -1 0 3224 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_19
timestamp 1744230924
transform -1 0 3416 0 -1 2210
box -4 -6 196 206
use BUFX2  BUFX2_11
timestamp 1744230924
transform -1 0 3464 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_32
timestamp 1744230924
transform 1 0 3464 0 -1 2210
box -4 -6 196 206
use INVX1  INVX1_5
timestamp 1744230924
transform 1 0 3656 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_1
timestamp 1744230924
transform 1 0 3688 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_2
timestamp 1744230924
transform 1 0 3752 0 -1 2210
box -4 -6 68 206
use XOR2X1  XOR2X1_9
timestamp 1744230924
transform 1 0 3816 0 -1 2210
box -4 -6 116 206
use INVX1  INVX1_7
timestamp 1744230924
transform 1 0 3928 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_3
timestamp 1744230924
transform -1 0 4024 0 -1 2210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_36
timestamp 1744230924
transform -1 0 4136 0 -1 2210
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_35
timestamp 1744230924
transform 1 0 4136 0 -1 2210
box -4 -6 196 206
use OR2X2  OR2X2_3
timestamp 1744230924
transform -1 0 4392 0 -1 2210
box -4 -6 68 206
use NOR2X1  NOR2X1_21
timestamp 1744230924
transform -1 0 4440 0 -1 2210
box -4 -6 52 206
use FILL  FILL_10_2_0
timestamp 1744230924
transform 1 0 4440 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_2_1
timestamp 1744230924
transform 1 0 4456 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_2_2
timestamp 1744230924
transform 1 0 4472 0 -1 2210
box -4 -6 20 206
use NAND2X1  NAND2X1_30
timestamp 1744230924
transform 1 0 4488 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_20
timestamp 1744230924
transform -1 0 4584 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_38
timestamp 1744230924
transform 1 0 4584 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_26
timestamp 1744230924
transform -1 0 4696 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_37
timestamp 1744230924
transform 1 0 4696 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_39
timestamp 1744230924
transform 1 0 4760 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_29
timestamp 1744230924
transform 1 0 4824 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_26
timestamp 1744230924
transform 1 0 4872 0 -1 2210
box -4 -6 36 206
use OAI22X1  OAI22X1_4
timestamp 1744230924
transform 1 0 4904 0 -1 2210
box -4 -6 84 206
use NAND2X1  NAND2X1_27
timestamp 1744230924
transform 1 0 4984 0 -1 2210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_17
timestamp 1744230924
transform 1 0 5032 0 -1 2210
box -4 -6 116 206
use XNOR2X1  XNOR2X1_67
timestamp 1744230924
transform -1 0 5256 0 -1 2210
box -4 -6 116 206
use AOI22X1  AOI22X1_22
timestamp 1744230924
transform 1 0 5256 0 -1 2210
box -4 -6 84 206
use NAND2X1  NAND2X1_150
timestamp 1744230924
transform -1 0 5384 0 -1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_151
timestamp 1744230924
transform 1 0 5384 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_159
timestamp 1744230924
transform 1 0 5432 0 -1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_50
timestamp 1744230924
transform 1 0 5624 0 -1 2210
box -4 -6 196 206
use BUFX2  BUFX2_34
timestamp 1744230924
transform 1 0 5816 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_125
timestamp 1744230924
transform -1 0 200 0 1 2210
box -4 -6 196 206
use XNOR2X1  XNOR2X1_81
timestamp 1744230924
transform -1 0 312 0 1 2210
box -4 -6 116 206
use XNOR2X1  XNOR2X1_80
timestamp 1744230924
transform -1 0 424 0 1 2210
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_126
timestamp 1744230924
transform -1 0 616 0 1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_127
timestamp 1744230924
transform 1 0 616 0 1 2210
box -4 -6 196 206
use XNOR2X1  XNOR2X1_51
timestamp 1744230924
transform 1 0 808 0 1 2210
box -4 -6 116 206
use NAND2X1  NAND2X1_123
timestamp 1744230924
transform -1 0 968 0 1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_69
timestamp 1744230924
transform -1 0 1160 0 1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_18
timestamp 1744230924
transform -1 0 1352 0 1 2210
box -4 -6 196 206
use FILL  FILL_11_0_0
timestamp 1744230924
transform 1 0 1352 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_0_1
timestamp 1744230924
transform 1 0 1368 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_0_2
timestamp 1744230924
transform 1 0 1384 0 1 2210
box -4 -6 20 206
use XNOR2X1  XNOR2X1_11
timestamp 1744230924
transform 1 0 1400 0 1 2210
box -4 -6 116 206
use OAI21X1  OAI21X1_32
timestamp 1744230924
transform 1 0 1512 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_31
timestamp 1744230924
transform 1 0 1576 0 1 2210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_14
timestamp 1744230924
transform -1 0 1832 0 1 2210
box -4 -6 196 206
use CLKBUF1  CLKBUF1_11
timestamp 1744230924
transform 1 0 1832 0 1 2210
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_13
timestamp 1744230924
transform -1 0 2168 0 1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_20
timestamp 1744230924
transform -1 0 2360 0 1 2210
box -4 -6 196 206
use INVX1  INVX1_8
timestamp 1744230924
transform 1 0 2360 0 1 2210
box -4 -6 36 206
use BUFX2  BUFX2_12
timestamp 1744230924
transform -1 0 2440 0 1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_28
timestamp 1744230924
transform 1 0 2440 0 1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_30
timestamp 1744230924
transform 1 0 2632 0 1 2210
box -4 -6 196 206
use INVX1  INVX1_3
timestamp 1744230924
transform 1 0 2824 0 1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_2
timestamp 1744230924
transform 1 0 2856 0 1 2210
box -4 -6 52 206
use FILL  FILL_11_1_0
timestamp 1744230924
transform -1 0 2920 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_1_1
timestamp 1744230924
transform -1 0 2936 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_1_2
timestamp 1744230924
transform -1 0 2952 0 1 2210
box -4 -6 20 206
use NOR2X1  NOR2X1_4
timestamp 1744230924
transform -1 0 3000 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_4
timestamp 1744230924
transform -1 0 3032 0 1 2210
box -4 -6 36 206
use NOR2X1  NOR2X1_3
timestamp 1744230924
transform 1 0 3032 0 1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_31
timestamp 1744230924
transform 1 0 3080 0 1 2210
box -4 -6 196 206
use NAND2X1  NAND2X1_4
timestamp 1744230924
transform -1 0 3320 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_6
timestamp 1744230924
transform 1 0 3320 0 1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_3
timestamp 1744230924
transform 1 0 3352 0 1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_3
timestamp 1744230924
transform 1 0 3400 0 1 2210
box -4 -6 196 206
use BUFX2  BUFX2_13
timestamp 1744230924
transform 1 0 3592 0 1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_11
timestamp 1744230924
transform -1 0 3832 0 1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_150
timestamp 1744230924
transform 1 0 3832 0 1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_149
timestamp 1744230924
transform 1 0 4024 0 1 2210
box -4 -6 196 206
use NAND2X1  NAND2X1_33
timestamp 1744230924
transform 1 0 4216 0 1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_24
timestamp 1744230924
transform 1 0 4264 0 1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_25
timestamp 1744230924
transform -1 0 4360 0 1 2210
box -4 -6 52 206
use NAND3X1  NAND3X1_1
timestamp 1744230924
transform -1 0 4456 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_25
timestamp 1744230924
transform 1 0 4360 0 1 2210
box -4 -6 36 206
use INVX1  INVX1_28
timestamp 1744230924
transform -1 0 4536 0 1 2210
box -4 -6 36 206
use FILL  FILL_11_2_2
timestamp 1744230924
transform -1 0 4504 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_2_1
timestamp 1744230924
transform -1 0 4488 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_2_0
timestamp 1744230924
transform -1 0 4472 0 1 2210
box -4 -6 20 206
use NAND2X1  NAND2X1_28
timestamp 1744230924
transform -1 0 4632 0 1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_18
timestamp 1744230924
transform -1 0 4584 0 1 2210
box -4 -6 52 206
use OAI22X1  OAI22X1_5
timestamp 1744230924
transform -1 0 4760 0 1 2210
box -4 -6 84 206
use NAND2X1  NAND2X1_35
timestamp 1744230924
transform 1 0 4632 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_27
timestamp 1744230924
transform 1 0 4760 0 1 2210
box -4 -6 36 206
use XNOR2X1  XNOR2X1_13
timestamp 1744230924
transform -1 0 4904 0 1 2210
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_156
timestamp 1744230924
transform 1 0 4904 0 1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_47
timestamp 1744230924
transform 1 0 5096 0 1 2210
box -4 -6 196 206
use BUFX2  BUFX2_31
timestamp 1744230924
transform 1 0 5288 0 1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_100
timestamp 1744230924
transform 1 0 5336 0 1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_37
timestamp 1744230924
transform 1 0 5528 0 1 2210
box -4 -6 196 206
use BUFX2  BUFX2_20
timestamp 1744230924
transform 1 0 5720 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_30
timestamp 1744230924
transform 1 0 5768 0 1 2210
box -4 -6 52 206
use FILL  FILL_12_1
timestamp 1744230924
transform 1 0 5816 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_2
timestamp 1744230924
transform 1 0 5832 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_3
timestamp 1744230924
transform 1 0 5848 0 1 2210
box -4 -6 20 206
use OAI21X1  OAI21X1_232
timestamp 1744230924
transform 1 0 8 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_175
timestamp 1744230924
transform -1 0 120 0 -1 2610
box -4 -6 52 206
use INVX2  INVX2_24
timestamp 1744230924
transform 1 0 120 0 -1 2610
box -4 -6 36 206
use INVX1  INVX1_144
timestamp 1744230924
transform 1 0 152 0 -1 2610
box -4 -6 36 206
use AOI21X1  AOI21X1_50
timestamp 1744230924
transform 1 0 184 0 -1 2610
box -4 -6 68 206
use MUX2X1  MUX2X1_10
timestamp 1744230924
transform 1 0 248 0 -1 2610
box -4 -6 100 206
use OAI21X1  OAI21X1_221
timestamp 1744230924
transform -1 0 408 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_174
timestamp 1744230924
transform -1 0 456 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_128
timestamp 1744230924
transform -1 0 504 0 -1 2610
box -4 -6 52 206
use XNOR2X1  XNOR2X1_79
timestamp 1744230924
transform -1 0 616 0 -1 2610
box -4 -6 116 206
use XNOR2X1  XNOR2X1_52
timestamp 1744230924
transform 1 0 616 0 -1 2610
box -4 -6 116 206
use AOI21X1  AOI21X1_28
timestamp 1744230924
transform 1 0 728 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_106
timestamp 1744230924
transform -1 0 824 0 -1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_156
timestamp 1744230924
transform 1 0 824 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_111
timestamp 1744230924
transform -1 0 920 0 -1 2610
box -4 -6 36 206
use INVX1  INVX1_104
timestamp 1744230924
transform -1 0 952 0 -1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_11
timestamp 1744230924
transform 1 0 952 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_162
timestamp 1744230924
transform 1 0 1016 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_112
timestamp 1744230924
transform -1 0 1112 0 -1 2610
box -4 -6 36 206
use NOR2X1  NOR2X1_83
timestamp 1744230924
transform -1 0 1160 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_155
timestamp 1744230924
transform -1 0 1224 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_81
timestamp 1744230924
transform -1 0 1272 0 -1 2610
box -4 -6 52 206
use XNOR2X1  XNOR2X1_75
timestamp 1744230924
transform 1 0 1272 0 -1 2610
box -4 -6 116 206
use FILL  FILL_12_0_0
timestamp 1744230924
transform 1 0 1384 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_0_1
timestamp 1744230924
transform 1 0 1400 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_0_2
timestamp 1744230924
transform 1 0 1416 0 -1 2610
box -4 -6 20 206
use XNOR2X1  XNOR2X1_76
timestamp 1744230924
transform 1 0 1432 0 -1 2610
box -4 -6 116 206
use NAND2X1  NAND2X1_24
timestamp 1744230924
transform 1 0 1544 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_29
timestamp 1744230924
transform 1 0 1592 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_23
timestamp 1744230924
transform -1 0 1704 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_33
timestamp 1744230924
transform -1 0 1768 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_16
timestamp 1744230924
transform -1 0 1816 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_30
timestamp 1744230924
transform -1 0 1880 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_23
timestamp 1744230924
transform -1 0 1912 0 -1 2610
box -4 -6 36 206
use INVX1  INVX1_22
timestamp 1744230924
transform -1 0 1944 0 -1 2610
box -4 -6 36 206
use NOR2X1  NOR2X1_15
timestamp 1744230924
transform -1 0 1992 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_6
timestamp 1744230924
transform -1 0 2184 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_8
timestamp 1744230924
transform -1 0 2376 0 -1 2610
box -4 -6 196 206
use BUFX2  BUFX2_15
timestamp 1744230924
transform -1 0 2424 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_12
timestamp 1744230924
transform -1 0 2616 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_5
timestamp 1744230924
transform -1 0 2808 0 -1 2610
box -4 -6 196 206
use BUFX2  BUFX2_14
timestamp 1744230924
transform -1 0 2856 0 -1 2610
box -4 -6 52 206
use FILL  FILL_12_1_0
timestamp 1744230924
transform -1 0 2872 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_1_1
timestamp 1744230924
transform -1 0 2888 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_1_2
timestamp 1744230924
transform -1 0 2904 0 -1 2610
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_4
timestamp 1744230924
transform -1 0 3096 0 -1 2610
box -4 -6 196 206
use XNOR2X1  XNOR2X1_4
timestamp 1744230924
transform 1 0 3096 0 -1 2610
box -4 -6 116 206
use OAI21X1  OAI21X1_15
timestamp 1744230924
transform -1 0 3272 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_14
timestamp 1744230924
transform 1 0 3272 0 -1 2610
box -4 -6 52 206
use OAI22X1  OAI22X1_1
timestamp 1744230924
transform 1 0 3320 0 -1 2610
box -4 -6 84 206
use NOR2X1  NOR2X1_9
timestamp 1744230924
transform 1 0 3400 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_13
timestamp 1744230924
transform -1 0 3496 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_8
timestamp 1744230924
transform 1 0 3496 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_12
timestamp 1744230924
transform -1 0 3576 0 -1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_14
timestamp 1744230924
transform -1 0 3640 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_13
timestamp 1744230924
transform -1 0 3672 0 -1 2610
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_170
timestamp 1744230924
transform -1 0 3864 0 -1 2610
box -4 -6 196 206
use AOI22X1  AOI22X1_2
timestamp 1744230924
transform 1 0 3864 0 -1 2610
box -4 -6 84 206
use NOR2X1  NOR2X1_26
timestamp 1744230924
transform 1 0 3944 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_169
timestamp 1744230924
transform -1 0 4184 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_161
timestamp 1744230924
transform -1 0 4376 0 -1 2610
box -4 -6 196 206
use AOI21X1  AOI21X1_4
timestamp 1744230924
transform 1 0 4376 0 -1 2610
box -4 -6 68 206
use FILL  FILL_12_2_0
timestamp 1744230924
transform -1 0 4456 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_2_1
timestamp 1744230924
transform -1 0 4472 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_2_2
timestamp 1744230924
transform -1 0 4488 0 -1 2610
box -4 -6 20 206
use NAND3X1  NAND3X1_2
timestamp 1744230924
transform -1 0 4552 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_23
timestamp 1744230924
transform -1 0 4600 0 -1 2610
box -4 -6 52 206
use AOI22X1  AOI22X1_1
timestamp 1744230924
transform 1 0 4600 0 -1 2610
box -4 -6 84 206
use INVX1  INVX1_29
timestamp 1744230924
transform 1 0 4680 0 -1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_42
timestamp 1744230924
transform -1 0 4776 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_32
timestamp 1744230924
transform -1 0 4824 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_40
timestamp 1744230924
transform -1 0 4888 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_31
timestamp 1744230924
transform -1 0 4936 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_17
timestamp 1744230924
transform 1 0 4936 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_19
timestamp 1744230924
transform -1 0 5032 0 -1 2610
box -4 -6 52 206
use XOR2X1  XOR2X1_2
timestamp 1744230924
transform -1 0 5144 0 -1 2610
box -4 -6 116 206
use XOR2X1  XOR2X1_3
timestamp 1744230924
transform 1 0 5144 0 -1 2610
box -4 -6 116 206
use XNOR2X1  XNOR2X1_72
timestamp 1744230924
transform -1 0 5368 0 -1 2610
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_99
timestamp 1744230924
transform 1 0 5368 0 -1 2610
box -4 -6 196 206
use BUFX2  BUFX2_29
timestamp 1744230924
transform 1 0 5560 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_36
timestamp 1744230924
transform 1 0 5608 0 -1 2610
box -4 -6 196 206
use BUFX2  BUFX2_19
timestamp 1744230924
transform 1 0 5800 0 -1 2610
box -4 -6 52 206
use FILL  FILL_13_1
timestamp 1744230924
transform -1 0 5864 0 -1 2610
box -4 -6 20 206
use AOI21X1  AOI21X1_51
timestamp 1744230924
transform -1 0 72 0 1 2610
box -4 -6 68 206
use XOR2X1  XOR2X1_24
timestamp 1744230924
transform -1 0 184 0 1 2610
box -4 -6 116 206
use INVX1  INVX1_113
timestamp 1744230924
transform 1 0 184 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_223
timestamp 1744230924
transform -1 0 280 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_147
timestamp 1744230924
transform 1 0 280 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_219
timestamp 1744230924
transform -1 0 376 0 1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_48
timestamp 1744230924
transform -1 0 440 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_143
timestamp 1744230924
transform -1 0 472 0 1 2610
box -4 -6 36 206
use AOI22X1  AOI22X1_25
timestamp 1744230924
transform 1 0 472 0 1 2610
box -4 -6 84 206
use INVX1  INVX1_149
timestamp 1744230924
transform 1 0 552 0 1 2610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_77
timestamp 1744230924
transform -1 0 696 0 1 2610
box -4 -6 116 206
use MUX2X1  MUX2X1_8
timestamp 1744230924
transform 1 0 696 0 1 2610
box -4 -6 100 206
use OAI21X1  OAI21X1_163
timestamp 1744230924
transform -1 0 856 0 1 2610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_53
timestamp 1744230924
transform 1 0 856 0 1 2610
box -4 -6 116 206
use AOI21X1  AOI21X1_29
timestamp 1744230924
transform 1 0 968 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_114
timestamp 1744230924
transform -1 0 1064 0 1 2610
box -4 -6 36 206
use NOR2X1  NOR2X1_82
timestamp 1744230924
transform 1 0 1064 0 1 2610
box -4 -6 52 206
use BUFX4  BUFX4_1
timestamp 1744230924
transform 1 0 1112 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_161
timestamp 1744230924
transform -1 0 1240 0 1 2610
box -4 -6 68 206
use INVX2  INVX2_15
timestamp 1744230924
transform 1 0 1240 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_211
timestamp 1744230924
transform -1 0 1336 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_172
timestamp 1744230924
transform 1 0 1336 0 1 2610
box -4 -6 52 206
use FILL  FILL_13_0_0
timestamp 1744230924
transform 1 0 1384 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_0_1
timestamp 1744230924
transform 1 0 1400 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_0_2
timestamp 1744230924
transform 1 0 1416 0 1 2610
box -4 -6 20 206
use OAI21X1  OAI21X1_220
timestamp 1744230924
transform 1 0 1432 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_35
timestamp 1744230924
transform -1 0 1560 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_24
timestamp 1744230924
transform -1 0 1592 0 1 2610
box -4 -6 36 206
use OAI22X1  OAI22X1_3
timestamp 1744230924
transform -1 0 1672 0 1 2610
box -4 -6 84 206
use OAI21X1  OAI21X1_34
timestamp 1744230924
transform 1 0 1672 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_25
timestamp 1744230924
transform -1 0 1784 0 1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_9
timestamp 1744230924
transform -1 0 1976 0 1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_10
timestamp 1744230924
transform -1 0 2168 0 1 2610
box -4 -6 196 206
use XNOR2X1  XNOR2X1_8
timestamp 1744230924
transform 1 0 2168 0 1 2610
box -4 -6 116 206
use AOI21X1  AOI21X1_1
timestamp 1744230924
transform 1 0 2280 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_12
timestamp 1744230924
transform 1 0 2344 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_20
timestamp 1744230924
transform -1 0 2456 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_19
timestamp 1744230924
transform -1 0 2520 0 1 2610
box -4 -6 68 206
use AND2X2  AND2X2_1
timestamp 1744230924
transform -1 0 2584 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_17
timestamp 1744230924
transform -1 0 2632 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_18
timestamp 1744230924
transform 1 0 2632 0 1 2610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_7
timestamp 1744230924
transform 1 0 2696 0 1 2610
box -4 -6 116 206
use INVX1  INVX1_16
timestamp 1744230924
transform -1 0 2840 0 1 2610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_5
timestamp 1744230924
transform 1 0 2840 0 1 2610
box -4 -6 116 206
use FILL  FILL_13_1_0
timestamp 1744230924
transform -1 0 2968 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_1_1
timestamp 1744230924
transform -1 0 2984 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_1_2
timestamp 1744230924
transform -1 0 3000 0 1 2610
box -4 -6 20 206
use NOR2X1  NOR2X1_11
timestamp 1744230924
transform -1 0 3048 0 1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_10
timestamp 1744230924
transform 1 0 3048 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_15
timestamp 1744230924
transform -1 0 3128 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_17
timestamp 1744230924
transform -1 0 3192 0 1 2610
box -4 -6 68 206
use OAI22X1  OAI22X1_2
timestamp 1744230924
transform -1 0 3272 0 1 2610
box -4 -6 84 206
use INVX1  INVX1_14
timestamp 1744230924
transform -1 0 3304 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_15
timestamp 1744230924
transform -1 0 3352 0 1 2610
box -4 -6 52 206
use OR2X2  OR2X2_1
timestamp 1744230924
transform -1 0 3416 0 1 2610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_171
timestamp 1744230924
transform -1 0 3608 0 1 2610
box -4 -6 196 206
use XNOR2X1  XNOR2X1_18
timestamp 1744230924
transform 1 0 3608 0 1 2610
box -4 -6 116 206
use OAI21X1  OAI21X1_45
timestamp 1744230924
transform -1 0 3784 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_34
timestamp 1744230924
transform -1 0 3816 0 1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_3
timestamp 1744230924
transform 1 0 3816 0 1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_6
timestamp 1744230924
transform 1 0 3880 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_33
timestamp 1744230924
transform -1 0 3976 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_36
timestamp 1744230924
transform -1 0 4024 0 1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_27
timestamp 1744230924
transform 1 0 4024 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_32
timestamp 1744230924
transform 1 0 4072 0 1 2610
box -4 -6 36 206
use INVX1  INVX1_31
timestamp 1744230924
transform -1 0 4136 0 1 2610
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_162
timestamp 1744230924
transform -1 0 4328 0 1 2610
box -4 -6 196 206
use NOR2X1  NOR2X1_22
timestamp 1744230924
transform -1 0 4376 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_41
timestamp 1744230924
transform -1 0 4440 0 1 2610
box -4 -6 68 206
use FILL  FILL_13_2_0
timestamp 1744230924
transform 1 0 4440 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_2_1
timestamp 1744230924
transform 1 0 4456 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_2_2
timestamp 1744230924
transform 1 0 4472 0 1 2610
box -4 -6 20 206
use XOR2X1  XOR2X1_1
timestamp 1744230924
transform 1 0 4488 0 1 2610
box -4 -6 116 206
use NAND2X1  NAND2X1_34
timestamp 1744230924
transform 1 0 4600 0 1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_154
timestamp 1744230924
transform 1 0 4648 0 1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_45
timestamp 1744230924
transform 1 0 4840 0 1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_155
timestamp 1744230924
transform 1 0 5032 0 1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_46
timestamp 1744230924
transform 1 0 5224 0 1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_160
timestamp 1744230924
transform 1 0 5416 0 1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_51
timestamp 1744230924
transform 1 0 5608 0 1 2610
box -4 -6 196 206
use BUFX2  BUFX2_35
timestamp 1744230924
transform 1 0 5800 0 1 2610
box -4 -6 52 206
use FILL  FILL_14_1
timestamp 1744230924
transform 1 0 5848 0 1 2610
box -4 -6 20 206
use INVX1  INVX1_150
timestamp 1744230924
transform 1 0 8 0 -1 3010
box -4 -6 36 206
use INVX1  INVX1_151
timestamp 1744230924
transform -1 0 72 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_231
timestamp 1744230924
transform -1 0 136 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_17
timestamp 1744230924
transform -1 0 200 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_227
timestamp 1744230924
transform 1 0 200 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_148
timestamp 1744230924
transform -1 0 296 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_222
timestamp 1744230924
transform -1 0 360 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_46
timestamp 1744230924
transform -1 0 424 0 -1 3010
box -4 -6 68 206
use AOI22X1  AOI22X1_26
timestamp 1744230924
transform 1 0 424 0 -1 3010
box -4 -6 84 206
use OAI21X1  OAI21X1_228
timestamp 1744230924
transform 1 0 504 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_229
timestamp 1744230924
transform -1 0 632 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_218
timestamp 1744230924
transform 1 0 632 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_171
timestamp 1744230924
transform -1 0 744 0 -1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_84
timestamp 1744230924
transform -1 0 792 0 -1 3010
box -4 -6 52 206
use AOI22X1  AOI22X1_17
timestamp 1744230924
transform -1 0 872 0 -1 3010
box -4 -6 84 206
use NAND2X1  NAND2X1_120
timestamp 1744230924
transform 1 0 872 0 -1 3010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_50
timestamp 1744230924
transform -1 0 1032 0 -1 3010
box -4 -6 116 206
use INVX2  INVX2_12
timestamp 1744230924
transform -1 0 1064 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_216
timestamp 1744230924
transform 1 0 1064 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_146
timestamp 1744230924
transform 1 0 1128 0 -1 3010
box -4 -6 36 206
use AOI21X1  AOI21X1_49
timestamp 1744230924
transform -1 0 1224 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_225
timestamp 1744230924
transform -1 0 1288 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_166
timestamp 1744230924
transform 1 0 1288 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_168
timestamp 1744230924
transform 1 0 1336 0 -1 3010
box -4 -6 52 206
use FILL  FILL_14_0_0
timestamp 1744230924
transform -1 0 1400 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_0_1
timestamp 1744230924
transform -1 0 1416 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_0_2
timestamp 1744230924
transform -1 0 1432 0 -1 3010
box -4 -6 20 206
use NAND2X1  NAND2X1_167
timestamp 1744230924
transform -1 0 1480 0 -1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_123
timestamp 1744230924
transform -1 0 1528 0 -1 3010
box -4 -6 52 206
use AOI21X1  AOI21X1_45
timestamp 1744230924
transform 1 0 1528 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_217
timestamp 1744230924
transform 1 0 1592 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_142
timestamp 1744230924
transform -1 0 1688 0 -1 3010
box -4 -6 36 206
use AOI21X1  AOI21X1_47
timestamp 1744230924
transform -1 0 1752 0 -1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_119
timestamp 1744230924
transform -1 0 1800 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_224
timestamp 1744230924
transform 1 0 1800 0 -1 3010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_78
timestamp 1744230924
transform 1 0 1864 0 -1 3010
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_119
timestamp 1744230924
transform -1 0 2168 0 -1 3010
box -4 -6 196 206
use BUFX2  BUFX2_49
timestamp 1744230924
transform -1 0 2216 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_36
timestamp 1744230924
transform 1 0 2216 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_58
timestamp 1744230924
transform 1 0 2264 0 -1 3010
box -4 -6 196 206
use XOR2X1  XOR2X1_16
timestamp 1744230924
transform -1 0 2568 0 -1 3010
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_1
timestamp 1744230924
transform -1 0 2760 0 -1 3010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_7
timestamp 1744230924
transform -1 0 2952 0 -1 3010
box -4 -6 196 206
use FILL  FILL_14_1_0
timestamp 1744230924
transform 1 0 2952 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_1_1
timestamp 1744230924
transform 1 0 2968 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_1_2
timestamp 1744230924
transform 1 0 2984 0 -1 3010
box -4 -6 20 206
use NAND2X1  NAND2X1_16
timestamp 1744230924
transform 1 0 3000 0 -1 3010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_6
timestamp 1744230924
transform -1 0 3160 0 -1 3010
box -4 -6 116 206
use OAI21X1  OAI21X1_16
timestamp 1744230924
transform -1 0 3224 0 -1 3010
box -4 -6 68 206
use OR2X2  OR2X2_2
timestamp 1744230924
transform -1 0 3288 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_172
timestamp 1744230924
transform -1 0 3480 0 -1 3010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_173
timestamp 1744230924
transform -1 0 3672 0 -1 3010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_167
timestamp 1744230924
transform -1 0 3864 0 -1 3010
box -4 -6 196 206
use XNOR2X1  XNOR2X1_19
timestamp 1744230924
transform -1 0 3976 0 -1 3010
box -4 -6 116 206
use OAI21X1  OAI21X1_47
timestamp 1744230924
transform -1 0 4040 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_36
timestamp 1744230924
transform 1 0 4040 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_46
timestamp 1744230924
transform -1 0 4136 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_168
timestamp 1744230924
transform -1 0 4328 0 -1 3010
box -4 -6 196 206
use XNOR2X1  XNOR2X1_24
timestamp 1744230924
transform -1 0 4440 0 -1 3010
box -4 -6 116 206
use FILL  FILL_14_2_0
timestamp 1744230924
transform 1 0 4440 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_2_1
timestamp 1744230924
transform 1 0 4456 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_2_2
timestamp 1744230924
transform 1 0 4472 0 -1 3010
box -4 -6 20 206
use INVX1  INVX1_43
timestamp 1744230924
transform 1 0 4488 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_60
timestamp 1744230924
transform 1 0 4520 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_59
timestamp 1744230924
transform 1 0 4584 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_158
timestamp 1744230924
transform 1 0 4648 0 -1 3010
box -4 -6 196 206
use XNOR2X1  XNOR2X1_14
timestamp 1744230924
transform -1 0 4952 0 -1 3010
box -4 -6 116 206
use CLKBUF1  CLKBUF1_4
timestamp 1744230924
transform 1 0 4952 0 -1 3010
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_49
timestamp 1744230924
transform 1 0 5096 0 -1 3010
box -4 -6 196 206
use BUFX2  BUFX2_17
timestamp 1744230924
transform -1 0 5336 0 -1 3010
box -4 -6 52 206
use DFFSR  DFFSR_1
timestamp 1744230924
transform -1 0 5688 0 -1 3010
box -4 -6 356 206
use NAND2X1  NAND2X1_226
timestamp 1744230924
transform 1 0 5688 0 -1 3010
box -4 -6 52 206
use OR2X2  OR2X2_15
timestamp 1744230924
transform -1 0 5800 0 -1 3010
box -4 -6 68 206
use BUFX2  BUFX2_33
timestamp 1744230924
transform 1 0 5800 0 -1 3010
box -4 -6 52 206
use FILL  FILL_15_1
timestamp 1744230924
transform -1 0 5864 0 -1 3010
box -4 -6 20 206
use OAI21X1  OAI21X1_230
timestamp 1744230924
transform -1 0 72 0 1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_125
timestamp 1744230924
transform 1 0 72 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_127
timestamp 1744230924
transform 1 0 120 0 1 3010
box -4 -6 52 206
use INVX2  INVX2_25
timestamp 1744230924
transform 1 0 168 0 1 3010
box -4 -6 36 206
use NOR2X1  NOR2X1_126
timestamp 1744230924
transform -1 0 248 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_226
timestamp 1744230924
transform -1 0 312 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_173
timestamp 1744230924
transform -1 0 360 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_124
timestamp 1744230924
transform -1 0 408 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_117
timestamp 1744230924
transform 1 0 408 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_150
timestamp 1744230924
transform -1 0 520 0 1 3010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_49
timestamp 1744230924
transform 1 0 520 0 1 3010
box -4 -6 116 206
use NAND2X1  NAND2X1_122
timestamp 1744230924
transform -1 0 680 0 1 3010
box -4 -6 52 206
use INVX1  INVX1_108
timestamp 1744230924
transform 1 0 680 0 1 3010
box -4 -6 36 206
use BUFX4  BUFX4_2
timestamp 1744230924
transform 1 0 712 0 1 3010
box -4 -6 68 206
use AOI22X1  AOI22X1_16
timestamp 1744230924
transform -1 0 856 0 1 3010
box -4 -6 84 206
use NAND2X1  NAND2X1_119
timestamp 1744230924
transform 1 0 856 0 1 3010
box -4 -6 52 206
use INVX1  INVX1_107
timestamp 1744230924
transform -1 0 936 0 1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_160
timestamp 1744230924
transform 1 0 936 0 1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_121
timestamp 1744230924
transform 1 0 1000 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_215
timestamp 1744230924
transform 1 0 1048 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_44
timestamp 1744230924
transform 1 0 1112 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_213
timestamp 1744230924
transform 1 0 1176 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_145
timestamp 1744230924
transform 1 0 1240 0 1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_165
timestamp 1744230924
transform -1 0 1320 0 1 3010
box -4 -6 52 206
use INVX1  INVX1_141
timestamp 1744230924
transform -1 0 1352 0 1 3010
box -4 -6 36 206
use FILL  FILL_15_0_0
timestamp 1744230924
transform -1 0 1368 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_0_1
timestamp 1744230924
transform -1 0 1384 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_0_2
timestamp 1744230924
transform -1 0 1400 0 1 3010
box -4 -6 20 206
use OAI21X1  OAI21X1_214
timestamp 1744230924
transform -1 0 1464 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_169
timestamp 1744230924
transform 1 0 1464 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_212
timestamp 1744230924
transform -1 0 1576 0 1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_122
timestamp 1744230924
transform -1 0 1624 0 1 3010
box -4 -6 52 206
use OR2X2  OR2X2_14
timestamp 1744230924
transform -1 0 1688 0 1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_118
timestamp 1744230924
transform -1 0 1736 0 1 3010
box -4 -6 52 206
use AND2X2  AND2X2_10
timestamp 1744230924
transform 1 0 1736 0 1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_120
timestamp 1744230924
transform -1 0 1992 0 1 3010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_61
timestamp 1744230924
transform -1 0 2184 0 1 3010
box -4 -6 196 206
use BUFX2  BUFX2_37
timestamp 1744230924
transform -1 0 2232 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_59
timestamp 1744230924
transform -1 0 2280 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_173
timestamp 1744230924
transform -1 0 2344 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_172
timestamp 1744230924
transform -1 0 2408 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_35
timestamp 1744230924
transform -1 0 2472 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_121
timestamp 1744230924
transform -1 0 2504 0 1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_170
timestamp 1744230924
transform 1 0 2504 0 1 3010
box -4 -6 68 206
use MUX2X1  MUX2X1_9
timestamp 1744230924
transform -1 0 2664 0 1 3010
box -4 -6 100 206
use BUFX4  BUFX4_11
timestamp 1744230924
transform -1 0 2728 0 1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_2
timestamp 1744230924
transform -1 0 2920 0 1 3010
box -4 -6 196 206
use FILL  FILL_15_1_0
timestamp 1744230924
transform -1 0 2936 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_1_1
timestamp 1744230924
transform -1 0 2952 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_1_2
timestamp 1744230924
transform -1 0 2968 0 1 3010
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_174
timestamp 1744230924
transform -1 0 3160 0 1 3010
box -4 -6 196 206
use BUFX4  BUFX4_10
timestamp 1744230924
transform 1 0 3160 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_40
timestamp 1744230924
transform -1 0 3272 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_39
timestamp 1744230924
transform -1 0 3320 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_51
timestamp 1744230924
transform -1 0 3384 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_50
timestamp 1744230924
transform -1 0 3448 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_49
timestamp 1744230924
transform -1 0 3512 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_37
timestamp 1744230924
transform -1 0 3544 0 1 3010
box -4 -6 36 206
use XNOR2X1  XNOR2X1_20
timestamp 1744230924
transform -1 0 3656 0 1 3010
box -4 -6 116 206
use XOR2X1  XOR2X1_4
timestamp 1744230924
transform 1 0 3656 0 1 3010
box -4 -6 116 206
use NAND2X1  NAND2X1_38
timestamp 1744230924
transform 1 0 3768 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_28
timestamp 1744230924
transform 1 0 3816 0 1 3010
box -4 -6 52 206
use OAI22X1  OAI22X1_6
timestamp 1744230924
transform -1 0 3944 0 1 3010
box -4 -6 84 206
use INVX1  INVX1_35
timestamp 1744230924
transform -1 0 3976 0 1 3010
box -4 -6 36 206
use OR2X2  OR2X2_4
timestamp 1744230924
transform -1 0 4040 0 1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_166
timestamp 1744230924
transform -1 0 4232 0 1 3010
box -4 -6 196 206
use AOI22X1  AOI22X1_3
timestamp 1744230924
transform -1 0 4312 0 1 3010
box -4 -6 84 206
use INVX1  INVX1_41
timestamp 1744230924
transform 1 0 4312 0 1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_61
timestamp 1744230924
transform -1 0 4408 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_45
timestamp 1744230924
transform 1 0 4408 0 1 3010
box -4 -6 52 206
use FILL  FILL_15_2_0
timestamp 1744230924
transform 1 0 4456 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_2_1
timestamp 1744230924
transform 1 0 4472 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_2_2
timestamp 1744230924
transform 1 0 4488 0 1 3010
box -4 -6 20 206
use NAND2X1  NAND2X1_44
timestamp 1744230924
transform 1 0 4504 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_58
timestamp 1744230924
transform -1 0 4616 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_42
timestamp 1744230924
transform -1 0 4648 0 1 3010
box -4 -6 36 206
use XNOR2X1  XNOR2X1_23
timestamp 1744230924
transform -1 0 4760 0 1 3010
box -4 -6 116 206
use INVX1  INVX1_38
timestamp 1744230924
transform -1 0 4792 0 1 3010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_153
timestamp 1744230924
transform 1 0 4792 0 1 3010
box -4 -6 196 206
use DFFSR  DFFSR_2
timestamp 1744230924
transform -1 0 5336 0 1 3010
box -4 -6 356 206
use NAND2X1  NAND2X1_227
timestamp 1744230924
transform -1 0 5384 0 1 3010
box -4 -6 52 206
use OR2X2  OR2X2_16
timestamp 1744230924
transform -1 0 5448 0 1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_106
timestamp 1744230924
transform 1 0 5448 0 1 3010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_43
timestamp 1744230924
transform 1 0 5640 0 1 3010
box -4 -6 196 206
use FILL  FILL_16_1
timestamp 1744230924
transform 1 0 5832 0 1 3010
box -4 -6 20 206
use FILL  FILL_16_2
timestamp 1744230924
transform 1 0 5848 0 1 3010
box -4 -6 20 206
use XNOR2X1  XNOR2X1_47
timestamp 1744230924
transform 1 0 8 0 -1 3410
box -4 -6 116 206
use INVX8  INVX8_3
timestamp 1744230924
transform -1 0 200 0 -1 3410
box -4 -6 84 206
use BUFX4  BUFX4_4
timestamp 1744230924
transform -1 0 264 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_103
timestamp 1744230924
transform 1 0 264 0 -1 3410
box -4 -6 36 206
use BUFX4  BUFX4_3
timestamp 1744230924
transform 1 0 296 0 -1 3410
box -4 -6 68 206
use AOI22X1  AOI22X1_15
timestamp 1744230924
transform 1 0 360 0 -1 3410
box -4 -6 84 206
use OAI21X1  OAI21X1_153
timestamp 1744230924
transform -1 0 504 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_10
timestamp 1744230924
transform -1 0 568 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_109
timestamp 1744230924
transform -1 0 600 0 -1 3410
box -4 -6 36 206
use INVX1  INVX1_105
timestamp 1744230924
transform 1 0 600 0 -1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_118
timestamp 1744230924
transform 1 0 632 0 -1 3410
box -4 -6 52 206
use NAND3X1  NAND3X1_9
timestamp 1744230924
transform -1 0 744 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_151
timestamp 1744230924
transform -1 0 808 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_116
timestamp 1744230924
transform 1 0 808 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_114
timestamp 1744230924
transform -1 0 904 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_154
timestamp 1744230924
transform -1 0 968 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_159
timestamp 1744230924
transform -1 0 1032 0 -1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_120
timestamp 1744230924
transform 1 0 1032 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_210
timestamp 1744230924
transform 1 0 1080 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_139
timestamp 1744230924
transform -1 0 1176 0 -1 3410
box -4 -6 36 206
use OAI22X1  OAI22X1_10
timestamp 1744230924
transform -1 0 1256 0 -1 3410
box -4 -6 84 206
use OAI21X1  OAI21X1_207
timestamp 1744230924
transform 1 0 1256 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_208
timestamp 1744230924
transform -1 0 1384 0 -1 3410
box -4 -6 68 206
use FILL  FILL_16_0_0
timestamp 1744230924
transform 1 0 1384 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_0_1
timestamp 1744230924
transform 1 0 1400 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_0_2
timestamp 1744230924
transform 1 0 1416 0 -1 3410
box -4 -6 20 206
use XNOR2X1  XNOR2X1_73
timestamp 1744230924
transform 1 0 1432 0 -1 3410
box -4 -6 116 206
use AOI21X1  AOI21X1_43
timestamp 1744230924
transform 1 0 1544 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_138
timestamp 1744230924
transform -1 0 1640 0 -1 3410
box -4 -6 36 206
use INVX1  INVX1_140
timestamp 1744230924
transform 1 0 1640 0 -1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_209
timestamp 1744230924
transform -1 0 1736 0 -1 3410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_74
timestamp 1744230924
transform -1 0 1848 0 -1 3410
box -4 -6 116 206
use CLKBUF1  CLKBUF1_13
timestamp 1744230924
transform -1 0 1992 0 -1 3410
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_118
timestamp 1744230924
transform -1 0 2184 0 -1 3410
box -4 -6 196 206
use XNOR2X1  XNOR2X1_57
timestamp 1744230924
transform -1 0 2296 0 -1 3410
box -4 -6 116 206
use XOR2X1  XOR2X1_15
timestamp 1744230924
transform -1 0 2408 0 -1 3410
box -4 -6 116 206
use OAI21X1  OAI21X1_171
timestamp 1744230924
transform -1 0 2472 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_133
timestamp 1744230924
transform -1 0 2520 0 -1 3410
box -4 -6 52 206
use NAND3X1  NAND3X1_12
timestamp 1744230924
transform 1 0 2520 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_134
timestamp 1744230924
transform -1 0 2632 0 -1 3410
box -4 -6 52 206
use AOI21X1  AOI21X1_36
timestamp 1744230924
transform 1 0 2632 0 -1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_96
timestamp 1744230924
transform 1 0 2696 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_169
timestamp 1744230924
transform 1 0 2744 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_120
timestamp 1744230924
transform 1 0 2808 0 -1 3410
box -4 -6 36 206
use AOI21X1  AOI21X1_34
timestamp 1744230924
transform 1 0 2840 0 -1 3410
box -4 -6 68 206
use FILL  FILL_16_1_0
timestamp 1744230924
transform -1 0 2920 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_1_1
timestamp 1744230924
transform -1 0 2936 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_1_2
timestamp 1744230924
transform -1 0 2952 0 -1 3410
box -4 -6 20 206
use NOR2X1  NOR2X1_95
timestamp 1744230924
transform -1 0 3000 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_168
timestamp 1744230924
transform 1 0 3000 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_130
timestamp 1744230924
transform 1 0 3064 0 -1 3410
box -4 -6 52 206
use AOI21X1  AOI21X1_33
timestamp 1744230924
transform -1 0 3176 0 -1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_94
timestamp 1744230924
transform 1 0 3176 0 -1 3410
box -4 -6 52 206
use XNOR2X1  XNOR2X1_100
timestamp 1744230924
transform 1 0 3224 0 -1 3410
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_112
timestamp 1744230924
transform -1 0 3528 0 -1 3410
box -4 -6 196 206
use INVX1  INVX1_96
timestamp 1744230924
transform -1 0 3560 0 -1 3410
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_110
timestamp 1744230924
transform -1 0 3752 0 -1 3410
box -4 -6 196 206
use OAI22X1  OAI22X1_7
timestamp 1744230924
transform 1 0 3752 0 -1 3410
box -4 -6 84 206
use OAI21X1  OAI21X1_48
timestamp 1744230924
transform -1 0 3896 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_37
timestamp 1744230924
transform 1 0 3896 0 -1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_165
timestamp 1744230924
transform -1 0 4136 0 -1 3410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_164
timestamp 1744230924
transform -1 0 4328 0 -1 3410
box -4 -6 196 206
use XNOR2X1  XNOR2X1_21
timestamp 1744230924
transform 1 0 4328 0 -1 3410
box -4 -6 116 206
use FILL  FILL_16_2_0
timestamp 1744230924
transform 1 0 4440 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_2_1
timestamp 1744230924
transform 1 0 4456 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_2_2
timestamp 1744230924
transform 1 0 4472 0 -1 3410
box -4 -6 20 206
use BUFX2  BUFX2_42
timestamp 1744230924
transform 1 0 4488 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_57
timestamp 1744230924
transform 1 0 4536 0 -1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_30
timestamp 1744230924
transform -1 0 4648 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_43
timestamp 1744230924
transform -1 0 4696 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_56
timestamp 1744230924
transform 1 0 4696 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_157
timestamp 1744230924
transform 1 0 4760 0 -1 3410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_44
timestamp 1744230924
transform 1 0 4952 0 -1 3410
box -4 -6 196 206
use BUFX2  BUFX2_50
timestamp 1744230924
transform 1 0 5144 0 -1 3410
box -4 -6 52 206
use DFFSR  DFFSR_16
timestamp 1744230924
transform -1 0 5544 0 -1 3410
box -4 -6 356 206
use DFFPOSX1  DFFPOSX1_105
timestamp 1744230924
transform -1 0 5736 0 -1 3410
box -4 -6 196 206
use BUFX2  BUFX2_21
timestamp 1744230924
transform 1 0 5736 0 -1 3410
box -4 -6 52 206
use BUFX2  BUFX2_27
timestamp 1744230924
transform 1 0 5784 0 -1 3410
box -4 -6 52 206
use FILL  FILL_17_1
timestamp 1744230924
transform -1 0 5848 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_2
timestamp 1744230924
transform -1 0 5864 0 -1 3410
box -4 -6 20 206
use NOR2X1  NOR2X1_78
timestamp 1744230924
transform -1 0 168 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_146
timestamp 1744230924
transform -1 0 120 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_113
timestamp 1744230924
transform 1 0 8 0 -1 3810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_48
timestamp 1744230924
transform 1 0 72 0 1 3410
box -4 -6 116 206
use OAI21X1  OAI21X1_147
timestamp 1744230924
transform -1 0 72 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_145
timestamp 1744230924
transform -1 0 264 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_102
timestamp 1744230924
transform -1 0 200 0 -1 3810
box -4 -6 36 206
use XNOR2X1  XNOR2X1_46
timestamp 1744230924
transform 1 0 216 0 1 3410
box -4 -6 116 206
use INVX1  INVX1_101
timestamp 1744230924
transform 1 0 184 0 1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_158
timestamp 1744230924
transform 1 0 360 0 -1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_85
timestamp 1744230924
transform 1 0 312 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_109
timestamp 1744230924
transform -1 0 312 0 -1 3810
box -4 -6 52 206
use OR2X2  OR2X2_10
timestamp 1744230924
transform 1 0 360 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_110
timestamp 1744230924
transform 1 0 328 0 1 3410
box -4 -6 36 206
use AOI21X1  AOI21X1_25
timestamp 1744230924
transform -1 0 488 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_148
timestamp 1744230924
transform -1 0 552 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_149
timestamp 1744230924
transform 1 0 552 0 1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_24
timestamp 1744230924
transform 1 0 616 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_79
timestamp 1744230924
transform -1 0 728 0 1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_76
timestamp 1744230924
transform 1 0 728 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_157
timestamp 1744230924
transform -1 0 488 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_115
timestamp 1744230924
transform -1 0 680 0 -1 3810
box -4 -6 196 206
use AND2X2  AND2X2_7
timestamp 1744230924
transform -1 0 744 0 -1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_26
timestamp 1744230924
transform 1 0 776 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_80
timestamp 1744230924
transform 1 0 840 0 1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_115
timestamp 1744230924
transform -1 0 936 0 1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_66
timestamp 1744230924
transform -1 0 1128 0 1 3410
box -4 -6 196 206
use INVX2  INVX2_14
timestamp 1744230924
transform -1 0 776 0 -1 3810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_121
timestamp 1744230924
transform -1 0 968 0 -1 3810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_65
timestamp 1744230924
transform -1 0 1160 0 -1 3810
box -4 -6 196 206
use XOR2X1  XOR2X1_22
timestamp 1744230924
transform 1 0 1208 0 1 3410
box -4 -6 116 206
use INVX2  INVX2_13
timestamp 1744230924
transform -1 0 1208 0 1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_170
timestamp 1744230924
transform -1 0 1176 0 1 3410
box -4 -6 52 206
use FILL  FILL_18_0_2
timestamp 1744230924
transform -1 0 1400 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_0_1
timestamp 1744230924
transform -1 0 1384 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_0_0
timestamp 1744230924
transform -1 0 1368 0 -1 3810
box -4 -6 20 206
use XOR2X1  XOR2X1_23
timestamp 1744230924
transform 1 0 1416 0 1 3410
box -4 -6 116 206
use FILL  FILL_17_0_2
timestamp 1744230924
transform 1 0 1400 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_0_1
timestamp 1744230924
transform 1 0 1384 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_0_0
timestamp 1744230924
transform 1 0 1368 0 1 3410
box -4 -6 20 206
use NAND2X1  NAND2X1_164
timestamp 1744230924
transform 1 0 1320 0 1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_59
timestamp 1744230924
transform -1 0 1592 0 -1 3810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_116
timestamp 1744230924
transform -1 0 1352 0 -1 3810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_60
timestamp 1744230924
transform -1 0 1720 0 1 3410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_117
timestamp 1744230924
transform -1 0 1912 0 1 3410
box -4 -6 196 206
use XNOR2X1  XNOR2X1_104
timestamp 1744230924
transform -1 0 1704 0 -1 3810
box -4 -6 116 206
use MUX2X1  MUX2X1_13
timestamp 1744230924
transform -1 0 1800 0 -1 3810
box -4 -6 100 206
use NOR2X1  NOR2X1_155
timestamp 1744230924
transform 1 0 1800 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_217
timestamp 1744230924
transform -1 0 1960 0 -1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_69
timestamp 1744230924
transform 1 0 1848 0 -1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_156
timestamp 1744230924
transform -1 0 1960 0 1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_215
timestamp 1744230924
transform 1 0 2008 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_225
timestamp 1744230924
transform 1 0 1960 0 -1 3810
box -4 -6 52 206
use XOR2X1  XOR2X1_34
timestamp 1744230924
transform 1 0 1960 0 1 3410
box -4 -6 116 206
use NAND2X1  NAND2X1_221
timestamp 1744230924
transform -1 0 2216 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_222
timestamp 1744230924
transform 1 0 2120 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_296
timestamp 1744230924
transform 1 0 2056 0 -1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_70
timestamp 1744230924
transform -1 0 2216 0 1 3410
box -4 -6 68 206
use OAI22X1  OAI22X1_12
timestamp 1744230924
transform -1 0 2152 0 1 3410
box -4 -6 84 206
use NAND2X1  NAND2X1_220
timestamp 1744230924
transform -1 0 2296 0 -1 3810
box -4 -6 52 206
use INVX2  INVX2_18
timestamp 1744230924
transform -1 0 2248 0 -1 3810
box -4 -6 36 206
use XOR2X1  XOR2X1_33
timestamp 1744230924
transform 1 0 2216 0 1 3410
box -4 -6 116 206
use INVX1  INVX1_116
timestamp 1744230924
transform -1 0 2440 0 -1 3810
box -4 -6 36 206
use XOR2X1  XOR2X1_32
timestamp 1744230924
transform 1 0 2296 0 -1 3810
box -4 -6 116 206
use NAND2X1  NAND2X1_131
timestamp 1744230924
transform -1 0 2440 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_298
timestamp 1744230924
transform -1 0 2392 0 1 3410
box -4 -6 68 206
use OAI22X1  OAI22X1_8
timestamp 1744230924
transform -1 0 2584 0 -1 3810
box -4 -6 84 206
use BUFX4  BUFX4_9
timestamp 1744230924
transform -1 0 2504 0 -1 3810
box -4 -6 68 206
use INVX4  INVX4_7
timestamp 1744230924
transform 1 0 2488 0 1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_132
timestamp 1744230924
transform 1 0 2440 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_164
timestamp 1744230924
transform -1 0 2696 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_124
timestamp 1744230924
transform 1 0 2584 0 -1 3810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_56
timestamp 1744230924
transform 1 0 2648 0 1 3410
box -4 -6 116 206
use INVX8  INVX8_1
timestamp 1744230924
transform -1 0 2648 0 1 3410
box -4 -6 84 206
use INVX2  INVX2_19
timestamp 1744230924
transform 1 0 2536 0 1 3410
box -4 -6 36 206
use INVX1  INVX1_117
timestamp 1744230924
transform -1 0 2792 0 -1 3810
box -4 -6 36 206
use AOI21X1  AOI21X1_31
timestamp 1744230924
transform -1 0 2760 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_167
timestamp 1744230924
transform 1 0 2760 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_127
timestamp 1744230924
transform -1 0 2904 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_283
timestamp 1744230924
transform 1 0 2792 0 -1 3810
box -4 -6 68 206
use FILL  FILL_17_1_1
timestamp 1744230924
transform 1 0 2888 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_1_0
timestamp 1744230924
transform 1 0 2872 0 1 3410
box -4 -6 20 206
use NAND2X1  NAND2X1_129
timestamp 1744230924
transform -1 0 2872 0 1 3410
box -4 -6 52 206
use FILL  FILL_17_1_2
timestamp 1744230924
transform 1 0 2904 0 1 3410
box -4 -6 20 206
use AOI21X1  AOI21X1_32
timestamp 1744230924
transform 1 0 2920 0 1 3410
box -4 -6 68 206
use FILL  FILL_18_1_0
timestamp 1744230924
transform 1 0 2904 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_1_1
timestamp 1744230924
transform 1 0 2920 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_1_2
timestamp 1744230924
transform 1 0 2936 0 -1 3810
box -4 -6 20 206
use BUFX4  BUFX4_8
timestamp 1744230924
transform 1 0 2952 0 -1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_93
timestamp 1744230924
transform -1 0 3032 0 1 3410
box -4 -6 52 206
use OR2X2  OR2X2_11
timestamp 1744230924
transform -1 0 3096 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_184
timestamp 1744230924
transform 1 0 3016 0 -1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_286
timestamp 1744230924
transform 1 0 3048 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_297
timestamp 1744230924
transform -1 0 3288 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_92
timestamp 1744230924
transform -1 0 3224 0 1 3410
box -4 -6 52 206
use INVX1  INVX1_119
timestamp 1744230924
transform 1 0 3144 0 1 3410
box -4 -6 36 206
use NOR2X1  NOR2X1_91
timestamp 1744230924
transform 1 0 3096 0 1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_55
timestamp 1744230924
transform -1 0 3304 0 -1 3810
box -4 -6 196 206
use INVX1  INVX1_118
timestamp 1744230924
transform -1 0 3320 0 1 3410
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_57
timestamp 1744230924
transform -1 0 3512 0 1 3410
box -4 -6 196 206
use INVX1  INVX1_186
timestamp 1744230924
transform -1 0 3544 0 1 3410
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_111
timestamp 1744230924
transform -1 0 3736 0 1 3410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_52
timestamp 1744230924
transform -1 0 3496 0 -1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_299
timestamp 1744230924
transform 1 0 3496 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_54
timestamp 1744230924
transform -1 0 3608 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_138
timestamp 1744230924
transform 1 0 3608 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_47
timestamp 1744230924
transform 1 0 3736 0 1 3410
box -4 -6 52 206
use XNOR2X1  XNOR2X1_45
timestamp 1744230924
transform 1 0 3784 0 1 3410
box -4 -6 116 206
use INVX2  INVX2_3
timestamp 1744230924
transform -1 0 3928 0 1 3410
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_163
timestamp 1744230924
transform -1 0 4120 0 1 3410
box -4 -6 196 206
use NOR2X1  NOR2X1_74
timestamp 1744230924
transform -1 0 3720 0 -1 3810
box -4 -6 52 206
use NOR2X1  NOR2X1_72
timestamp 1744230924
transform 1 0 3720 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_137
timestamp 1744230924
transform -1 0 3832 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_94
timestamp 1744230924
transform -1 0 3864 0 -1 3810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_107
timestamp 1744230924
transform -1 0 4056 0 -1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_54
timestamp 1744230924
transform -1 0 4184 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_52
timestamp 1744230924
transform -1 0 4248 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_55
timestamp 1744230924
transform 1 0 4248 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_53
timestamp 1744230924
transform -1 0 4376 0 1 3410
box -4 -6 68 206
use INVX4  INVX4_1
timestamp 1744230924
transform -1 0 4104 0 -1 3810
box -4 -6 52 206
use DFFSR  DFFSR_7
timestamp 1744230924
transform -1 0 4456 0 -1 3810
box -4 -6 356 206
use INVX1  INVX1_39
timestamp 1744230924
transform -1 0 4408 0 1 3410
box -4 -6 36 206
use INVX1  INVX1_40
timestamp 1744230924
transform -1 0 4440 0 1 3410
box -4 -6 36 206
use FILL  FILL_17_2_0
timestamp 1744230924
transform 1 0 4440 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_2_1
timestamp 1744230924
transform 1 0 4456 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_2_2
timestamp 1744230924
transform 1 0 4472 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_2_0
timestamp 1744230924
transform -1 0 4472 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_2_1
timestamp 1744230924
transform -1 0 4488 0 -1 3810
box -4 -6 20 206
use NOR2X1  NOR2X1_29
timestamp 1744230924
transform 1 0 4488 0 1 3410
box -4 -6 52 206
use FILL  FILL_18_2_2
timestamp 1744230924
transform -1 0 4504 0 -1 3810
box -4 -6 20 206
use OR2X2  OR2X2_21
timestamp 1744230924
transform -1 0 4568 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_42
timestamp 1744230924
transform 1 0 4648 0 1 3410
box -4 -6 52 206
use AOI21X1  AOI21X1_7
timestamp 1744230924
transform -1 0 4648 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_41
timestamp 1744230924
transform 1 0 4536 0 1 3410
box -4 -6 52 206
use DFFSR  DFFSR_5
timestamp 1744230924
transform -1 0 4920 0 -1 3810
box -4 -6 356 206
use XNOR2X1  XNOR2X1_22
timestamp 1744230924
transform -1 0 4808 0 1 3410
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_48
timestamp 1744230924
transform -1 0 5000 0 1 3410
box -4 -6 196 206
use CLKBUF1  CLKBUF1_2
timestamp 1744230924
transform 1 0 5000 0 1 3410
box -4 -6 148 206
use OR2X2  OR2X2_19
timestamp 1744230924
transform -1 0 4984 0 -1 3810
box -4 -6 68 206
use DFFSR  DFFSR_10
timestamp 1744230924
transform 1 0 4984 0 -1 3810
box -4 -6 356 206
use DFFSR  DFFSR_17
timestamp 1744230924
transform 1 0 5144 0 1 3410
box -4 -6 356 206
use INVX8  INVX8_4
timestamp 1744230924
transform 1 0 5336 0 -1 3810
box -4 -6 84 206
use DFFSR  DFFSR_9
timestamp 1744230924
transform 1 0 5496 0 1 3410
box -4 -6 356 206
use BUFX4  BUFX4_22
timestamp 1744230924
transform 1 0 5416 0 -1 3810
box -4 -6 68 206
use DFFSR  DFFSR_14
timestamp 1744230924
transform 1 0 5480 0 -1 3810
box -4 -6 356 206
use FILL  FILL_18_1
timestamp 1744230924
transform 1 0 5848 0 1 3410
box -4 -6 20 206
use FILL  FILL_19_1
timestamp 1744230924
transform -1 0 5848 0 -1 3810
box -4 -6 20 206
use FILL  FILL_19_2
timestamp 1744230924
transform -1 0 5864 0 -1 3810
box -4 -6 20 206
use OAI21X1  OAI21X1_144
timestamp 1744230924
transform 1 0 8 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_108
timestamp 1744230924
transform 1 0 72 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_110
timestamp 1744230924
transform -1 0 168 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_111
timestamp 1744230924
transform -1 0 216 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_112
timestamp 1744230924
transform 1 0 216 0 1 3810
box -4 -6 52 206
use NOR2X1  NOR2X1_86
timestamp 1744230924
transform -1 0 312 0 1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_27
timestamp 1744230924
transform 1 0 312 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_152
timestamp 1744230924
transform -1 0 440 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_121
timestamp 1744230924
transform -1 0 488 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_106
timestamp 1744230924
transform 1 0 488 0 1 3810
box -4 -6 52 206
use NOR2X1  NOR2X1_77
timestamp 1744230924
transform -1 0 584 0 1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_23
timestamp 1744230924
transform -1 0 648 0 1 3810
box -4 -6 68 206
use XOR2X1  XOR2X1_14
timestamp 1744230924
transform -1 0 760 0 1 3810
box -4 -6 116 206
use INVX1  INVX1_99
timestamp 1744230924
transform 1 0 760 0 1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_140
timestamp 1744230924
transform 1 0 792 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_139
timestamp 1744230924
transform -1 0 920 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_104
timestamp 1744230924
transform -1 0 968 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_102
timestamp 1744230924
transform -1 0 1016 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_98
timestamp 1744230924
transform 1 0 1016 0 1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_103
timestamp 1744230924
transform -1 0 1096 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_97
timestamp 1744230924
transform -1 0 1128 0 1 3810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_64
timestamp 1744230924
transform -1 0 1320 0 1 3810
box -4 -6 196 206
use FILL  FILL_19_0_0
timestamp 1744230924
transform 1 0 1320 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_0_1
timestamp 1744230924
transform 1 0 1336 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_0_2
timestamp 1744230924
transform 1 0 1352 0 1 3810
box -4 -6 20 206
use XNOR2X1  XNOR2X1_103
timestamp 1744230924
transform 1 0 1368 0 1 3810
box -4 -6 116 206
use XNOR2X1  XNOR2X1_54
timestamp 1744230924
transform 1 0 1480 0 1 3810
box -4 -6 116 206
use OAI21X1  OAI21X1_294
timestamp 1744230924
transform 1 0 1592 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_291
timestamp 1744230924
transform -1 0 1720 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_224
timestamp 1744230924
transform -1 0 1768 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_293
timestamp 1744230924
transform 1 0 1768 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_292
timestamp 1744230924
transform -1 0 1896 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_216
timestamp 1744230924
transform 1 0 1896 0 1 3810
box -4 -6 52 206
use INVX2  INVX2_17
timestamp 1744230924
transform -1 0 1976 0 1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_295
timestamp 1744230924
transform 1 0 1976 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_153
timestamp 1744230924
transform 1 0 2040 0 1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_68
timestamp 1744230924
transform 1 0 2088 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_154
timestamp 1744230924
transform -1 0 2200 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_212
timestamp 1744230924
transform -1 0 2248 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_213
timestamp 1744230924
transform -1 0 2296 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_185
timestamp 1744230924
transform 1 0 2296 0 1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_289
timestamp 1744230924
transform 1 0 2328 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_211
timestamp 1744230924
transform -1 0 2440 0 1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_30
timestamp 1744230924
transform -1 0 2504 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_90
timestamp 1744230924
transform 1 0 2504 0 1 3810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_55
timestamp 1744230924
transform 1 0 2552 0 1 3810
box -4 -6 116 206
use NAND2X1  NAND2X1_126
timestamp 1744230924
transform -1 0 2712 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_128
timestamp 1744230924
transform -1 0 2760 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_166
timestamp 1744230924
transform 1 0 2760 0 1 3810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_99
timestamp 1744230924
transform 1 0 2824 0 1 3810
box -4 -6 116 206
use FILL  FILL_19_1_0
timestamp 1744230924
transform 1 0 2936 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_1_1
timestamp 1744230924
transform 1 0 2952 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_1_2
timestamp 1744230924
transform 1 0 2968 0 1 3810
box -4 -6 20 206
use NOR2X1  NOR2X1_151
timestamp 1744230924
transform 1 0 2984 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_214
timestamp 1744230924
transform 1 0 3032 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_210
timestamp 1744230924
transform -1 0 3128 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_285
timestamp 1744230924
transform -1 0 3192 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_284
timestamp 1744230924
transform 1 0 3192 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_183
timestamp 1744230924
transform -1 0 3288 0 1 3810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_53
timestamp 1744230924
transform -1 0 3480 0 1 3810
box -4 -6 196 206
use NOR2X1  NOR2X1_71
timestamp 1744230924
transform -1 0 3528 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_46
timestamp 1744230924
transform 1 0 3528 0 1 3810
box -4 -6 52 206
use INVX2  INVX2_11
timestamp 1744230924
transform 1 0 3576 0 1 3810
box -4 -6 36 206
use NOR2X1  NOR2X1_73
timestamp 1744230924
transform -1 0 3656 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_51
timestamp 1744230924
transform -1 0 3704 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_53
timestamp 1744230924
transform -1 0 3752 0 1 3810
box -4 -6 52 206
use CLKBUF1  CLKBUF1_12
timestamp 1744230924
transform -1 0 3896 0 1 3810
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_108
timestamp 1744230924
transform -1 0 4088 0 1 3810
box -4 -6 196 206
use BUFX2  BUFX2_39
timestamp 1744230924
transform -1 0 4136 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_41
timestamp 1744230924
transform 1 0 4136 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_16
timestamp 1744230924
transform 1 0 4184 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_43
timestamp 1744230924
transform 1 0 4232 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_40
timestamp 1744230924
transform 1 0 4280 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_232
timestamp 1744230924
transform 1 0 4328 0 1 3810
box -4 -6 52 206
use FILL  FILL_19_2_0
timestamp 1744230924
transform -1 0 4392 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_2_1
timestamp 1744230924
transform -1 0 4408 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_2_2
timestamp 1744230924
transform -1 0 4424 0 1 3810
box -4 -6 20 206
use DFFSR  DFFSR_3
timestamp 1744230924
transform -1 0 4776 0 1 3810
box -4 -6 356 206
use NAND2X1  NAND2X1_228
timestamp 1744230924
transform -1 0 4824 0 1 3810
box -4 -6 52 206
use OR2X2  OR2X2_17
timestamp 1744230924
transform -1 0 4888 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_230
timestamp 1744230924
transform -1 0 4936 0 1 3810
box -4 -6 52 206
use BUFX4  BUFX4_21
timestamp 1744230924
transform -1 0 5000 0 1 3810
box -4 -6 68 206
use BUFX4  BUFX4_23
timestamp 1744230924
transform -1 0 5064 0 1 3810
box -4 -6 68 206
use BUFX2  BUFX2_28
timestamp 1744230924
transform -1 0 5112 0 1 3810
box -4 -6 52 206
use DFFSR  DFFSR_11
timestamp 1744230924
transform 1 0 5112 0 1 3810
box -4 -6 356 206
use DFFSR  DFFSR_13
timestamp 1744230924
transform 1 0 5464 0 1 3810
box -4 -6 356 206
use FILL  FILL_20_1
timestamp 1744230924
transform 1 0 5816 0 1 3810
box -4 -6 20 206
use FILL  FILL_20_2
timestamp 1744230924
transform 1 0 5832 0 1 3810
box -4 -6 20 206
use FILL  FILL_20_3
timestamp 1744230924
transform 1 0 5848 0 1 3810
box -4 -6 20 206
use OAI21X1  OAI21X1_142
timestamp 1744230924
transform -1 0 72 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_100
timestamp 1744230924
transform -1 0 104 0 -1 4210
box -4 -6 36 206
use OR2X2  OR2X2_9
timestamp 1744230924
transform 1 0 104 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_105
timestamp 1744230924
transform 1 0 168 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_143
timestamp 1744230924
transform -1 0 280 0 -1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_75
timestamp 1744230924
transform 1 0 280 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_141
timestamp 1744230924
transform 1 0 328 0 -1 4210
box -4 -6 68 206
use AND2X2  AND2X2_6
timestamp 1744230924
transform -1 0 456 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_114
timestamp 1744230924
transform -1 0 648 0 -1 4210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_63
timestamp 1744230924
transform -1 0 840 0 -1 4210
box -4 -6 196 206
use CLKBUF1  CLKBUF1_9
timestamp 1744230924
transform -1 0 984 0 -1 4210
box -4 -6 148 206
use NAND2X1  NAND2X1_107
timestamp 1744230924
transform 1 0 984 0 -1 4210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_62
timestamp 1744230924
transform -1 0 1224 0 -1 4210
box -4 -6 196 206
use XNOR2X1  XNOR2X1_102
timestamp 1744230924
transform 1 0 1224 0 -1 4210
box -4 -6 116 206
use FILL  FILL_20_0_0
timestamp 1744230924
transform -1 0 1352 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_0_1
timestamp 1744230924
transform -1 0 1368 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_0_2
timestamp 1744230924
transform -1 0 1384 0 -1 4210
box -4 -6 20 206
use OAI21X1  OAI21X1_290
timestamp 1744230924
transform -1 0 1448 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_219
timestamp 1744230924
transform -1 0 1496 0 -1 4210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_101
timestamp 1744230924
transform 1 0 1496 0 -1 4210
box -4 -6 116 206
use NAND2X1  NAND2X1_223
timestamp 1744230924
transform 1 0 1608 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_218
timestamp 1744230924
transform -1 0 1704 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_287
timestamp 1744230924
transform 1 0 1704 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_288
timestamp 1744230924
transform -1 0 1832 0 -1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_152
timestamp 1744230924
transform 1 0 1832 0 -1 4210
box -4 -6 52 206
use AOI21X1  AOI21X1_67
timestamp 1744230924
transform -1 0 1944 0 -1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_89
timestamp 1744230924
transform -1 0 1992 0 -1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_88
timestamp 1744230924
transform -1 0 2040 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_57
timestamp 1744230924
transform -1 0 2088 0 -1 4210
box -4 -6 52 206
use INVX1  INVX1_115
timestamp 1744230924
transform -1 0 2120 0 -1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_87
timestamp 1744230924
transform 1 0 2120 0 -1 4210
box -4 -6 52 206
use INVX2  INVX2_16
timestamp 1744230924
transform 1 0 2168 0 -1 4210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_54
timestamp 1744230924
transform -1 0 2392 0 -1 4210
box -4 -6 196 206
use INVX1  INVX1_95
timestamp 1744230924
transform -1 0 2424 0 -1 4210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_56
timestamp 1744230924
transform -1 0 2616 0 -1 4210
box -4 -6 196 206
use BUFX2  BUFX2_58
timestamp 1744230924
transform -1 0 2664 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_125
timestamp 1744230924
transform 1 0 2664 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_165
timestamp 1744230924
transform 1 0 2712 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_113
timestamp 1744230924
transform -1 0 2968 0 -1 4210
box -4 -6 196 206
use FILL  FILL_20_1_0
timestamp 1744230924
transform -1 0 2984 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_1_1
timestamp 1744230924
transform -1 0 3000 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_1_2
timestamp 1744230924
transform -1 0 3016 0 -1 4210
box -4 -6 20 206
use CLKBUF1  CLKBUF1_8
timestamp 1744230924
transform -1 0 3160 0 -1 4210
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_109
timestamp 1744230924
transform -1 0 3352 0 -1 4210
box -4 -6 196 206
use BUFX2  BUFX2_45
timestamp 1744230924
transform -1 0 3400 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_18
timestamp 1744230924
transform -1 0 3448 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_52
timestamp 1744230924
transform 1 0 3448 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_55
timestamp 1744230924
transform -1 0 3544 0 -1 4210
box -4 -6 52 206
use DFFSR  DFFSR_8
timestamp 1744230924
transform -1 0 3896 0 -1 4210
box -4 -6 356 206
use NAND2X1  NAND2X1_233
timestamp 1744230924
transform -1 0 3944 0 -1 4210
box -4 -6 52 206
use OR2X2  OR2X2_22
timestamp 1744230924
transform -1 0 4008 0 -1 4210
box -4 -6 68 206
use DFFSR  DFFSR_4
timestamp 1744230924
transform -1 0 4360 0 -1 4210
box -4 -6 356 206
use NAND2X1  NAND2X1_229
timestamp 1744230924
transform -1 0 4408 0 -1 4210
box -4 -6 52 206
use FILL  FILL_20_2_0
timestamp 1744230924
transform -1 0 4424 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_2_1
timestamp 1744230924
transform -1 0 4440 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_2_2
timestamp 1744230924
transform -1 0 4456 0 -1 4210
box -4 -6 20 206
use OR2X2  OR2X2_18
timestamp 1744230924
transform -1 0 4520 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_44
timestamp 1744230924
transform -1 0 4568 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_32
timestamp 1744230924
transform 1 0 4568 0 -1 4210
box -4 -6 52 206
use DFFSR  DFFSR_6
timestamp 1744230924
transform -1 0 4968 0 -1 4210
box -4 -6 356 206
use NAND2X1  NAND2X1_231
timestamp 1744230924
transform -1 0 5016 0 -1 4210
box -4 -6 52 206
use OR2X2  OR2X2_20
timestamp 1744230924
transform -1 0 5080 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_56
timestamp 1744230924
transform 1 0 5080 0 -1 4210
box -4 -6 52 206
use DFFSR  DFFSR_12
timestamp 1744230924
transform 1 0 5128 0 -1 4210
box -4 -6 356 206
use DFFSR  DFFSR_15
timestamp 1744230924
transform -1 0 5832 0 -1 4210
box -4 -6 356 206
use FILL  FILL_21_1
timestamp 1744230924
transform -1 0 5848 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_2
timestamp 1744230924
transform -1 0 5864 0 -1 4210
box -4 -6 20 206
<< labels >>
flabel metal4 s 1352 0 1400 24 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 2904 0 2952 24 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 973 4237 979 4243 3 FreeSans 24 90 0 0 clk
port 2 nsew
flabel metal2 s 3933 4237 3939 4243 3 FreeSans 24 90 0 0 rst
port 3 nsew
flabel metal3 s 5885 2937 5891 2943 3 FreeSans 24 0 0 0 theta[0]
port 4 nsew
flabel metal3 s 5885 3097 5891 3103 3 FreeSans 24 0 0 0 theta[1]
port 5 nsew
flabel metal2 s 4781 4237 4787 4243 3 FreeSans 24 90 0 0 theta[2]
port 6 nsew
flabel metal2 s 4221 4237 4227 4243 3 FreeSans 24 90 0 0 theta[3]
port 7 nsew
flabel metal2 s 4893 4237 4899 4243 3 FreeSans 24 90 0 0 theta[4]
port 8 nsew
flabel metal2 s 4829 4237 4835 4243 3 FreeSans 24 90 0 0 theta[5]
port 9 nsew
flabel metal2 s 4381 4237 4387 4243 3 FreeSans 24 90 0 0 theta[6]
port 10 nsew
flabel metal2 s 3757 4237 3763 4243 3 FreeSans 24 90 0 0 theta[7]
port 11 nsew
flabel metal2 s 5085 4237 5091 4243 3 FreeSans 24 90 0 0 sine[0]
port 12 nsew
flabel metal3 s 5885 2497 5891 2503 3 FreeSans 24 0 0 0 sine[1]
port 13 nsew
flabel metal3 s 5885 2377 5891 2383 3 FreeSans 24 0 0 0 sine[2]
port 14 nsew
flabel metal3 s 5885 2337 5891 2343 3 FreeSans 24 0 0 0 sine[3]
port 15 nsew
flabel metal2 s 4589 4237 4595 4243 3 FreeSans 24 90 0 0 sine[4]
port 16 nsew
flabel metal3 s 5885 2897 5891 2903 3 FreeSans 24 0 0 0 sine[5]
port 17 nsew
flabel metal3 s 5885 2097 5891 2103 3 FreeSans 24 0 0 0 sine[6]
port 18 nsew
flabel metal3 s 5885 2697 5891 2703 3 FreeSans 24 0 0 0 sine[7]
port 19 nsew
flabel metal3 s 5885 2537 5891 2543 3 FreeSans 24 0 0 0 cosine[0]
port 20 nsew
flabel metal3 s 5885 2297 5891 2303 3 FreeSans 24 0 0 0 cosine[1]
port 21 nsew
flabel metal3 s 5885 3297 5891 3303 3 FreeSans 24 0 0 0 cosine[2]
port 22 nsew
flabel metal3 s 5885 897 5891 903 3 FreeSans 24 0 0 0 cosine[3]
port 23 nsew
flabel metal3 s 5885 1697 5891 1703 3 FreeSans 24 0 0 0 cosine[4]
port 24 nsew
flabel metal3 s 5885 697 5891 703 3 FreeSans 24 0 0 0 cosine[5]
port 25 nsew
flabel metal3 s 5885 937 5891 943 3 FreeSans 24 0 0 0 cosine[6]
port 26 nsew
flabel metal3 s 5885 97 5891 103 3 FreeSans 24 0 0 0 cosine[7]
port 27 nsew
flabel metal3 s 5885 3337 5891 3343 3 FreeSans 24 0 0 0 done
port 28 nsew
<< end >>

magic
tech scmos
timestamp 0
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 450 1500
string LEFsymmetry Y
string LEFview TRUE
<< end >>

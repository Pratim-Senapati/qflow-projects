VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sincos
  CLASS BLOCK ;
  FOREIGN sincos ;
  ORIGIN -0.400 0.000 ;
  SIZE 588.700 BY 424.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 290.800 412.400 291.600 412.600 ;
        RECT 293.400 412.400 294.200 412.600 ;
        RECT 289.200 411.800 294.200 412.400 ;
        RECT 289.200 411.600 290.000 411.800 ;
        RECT 455.600 411.600 456.400 413.200 ;
        RECT 508.400 411.600 509.200 413.200 ;
        RECT 542.600 410.800 543.400 411.000 ;
        RECT 516.400 410.200 543.400 410.800 ;
        RECT 552.600 410.800 553.400 411.000 ;
        RECT 552.600 410.200 579.600 410.800 ;
        RECT 1.800 401.600 2.600 406.200 ;
        RECT 6.000 401.600 6.800 410.200 ;
        RECT 9.200 401.600 10.000 406.200 ;
        RECT 13.400 401.600 14.200 410.200 ;
        RECT 17.200 401.600 18.000 406.200 ;
        RECT 20.400 401.600 21.200 406.200 ;
        RECT 22.600 401.600 23.400 406.200 ;
        RECT 26.800 401.600 27.600 410.200 ;
        RECT 28.400 401.600 29.200 410.200 ;
        RECT 33.200 401.600 34.000 410.200 ;
        RECT 37.400 401.600 38.200 406.200 ;
        RECT 41.200 401.600 42.000 409.800 ;
        RECT 44.400 401.600 45.200 406.200 ;
        RECT 47.600 401.600 48.400 410.200 ;
        RECT 53.200 401.600 54.000 406.200 ;
        RECT 56.400 401.600 57.200 406.200 ;
        RECT 62.000 401.600 62.800 410.000 ;
        RECT 66.800 401.600 67.600 410.200 ;
        RECT 72.400 401.600 73.200 406.200 ;
        RECT 75.600 401.600 76.400 406.200 ;
        RECT 81.200 401.600 82.000 410.000 ;
        RECT 84.400 401.600 85.200 410.200 ;
        RECT 87.600 401.600 88.400 410.200 ;
        RECT 90.800 401.600 91.600 410.200 ;
        RECT 94.000 401.600 94.800 410.200 ;
        RECT 97.200 401.600 98.000 410.200 ;
        RECT 98.800 401.600 99.600 406.200 ;
        RECT 102.000 401.600 102.800 406.200 ;
        RECT 105.200 401.600 106.000 410.200 ;
        RECT 110.800 401.600 111.600 406.200 ;
        RECT 114.000 401.600 114.800 406.200 ;
        RECT 119.600 401.600 120.400 410.000 ;
        RECT 124.400 402.200 125.400 408.800 ;
        RECT 124.600 401.600 125.400 402.200 ;
        RECT 130.600 401.600 131.600 408.800 ;
        RECT 139.400 401.600 140.200 406.200 ;
        RECT 143.600 401.600 144.400 410.200 ;
        RECT 145.200 401.600 146.000 406.200 ;
        RECT 148.400 401.600 149.200 406.200 ;
        RECT 151.600 402.200 152.600 408.800 ;
        RECT 151.800 401.600 152.600 402.200 ;
        RECT 157.800 401.600 158.800 408.800 ;
        RECT 161.200 401.600 162.000 406.200 ;
        RECT 164.400 401.600 165.200 406.200 ;
        RECT 166.000 401.600 166.800 406.200 ;
        RECT 169.200 401.600 170.000 406.200 ;
        RECT 170.800 401.600 171.600 410.200 ;
        RECT 175.000 401.600 175.800 406.200 ;
        RECT 177.800 401.600 178.600 406.200 ;
        RECT 182.000 401.600 182.800 410.200 ;
        RECT 183.600 401.600 184.400 410.200 ;
        RECT 191.600 401.600 192.400 409.000 ;
        RECT 198.000 401.600 198.800 410.200 ;
        RECT 202.800 401.600 203.600 410.200 ;
        RECT 206.000 401.600 206.800 409.000 ;
        RECT 210.800 401.600 211.600 406.200 ;
        RECT 212.400 401.600 213.200 410.200 ;
        RECT 217.200 401.600 218.000 410.200 ;
        RECT 222.000 401.600 222.800 410.200 ;
        RECT 227.600 401.600 228.400 406.200 ;
        RECT 230.800 401.600 231.600 406.200 ;
        RECT 236.400 401.600 237.200 410.000 ;
        RECT 241.200 401.600 242.000 406.200 ;
        RECT 244.400 401.600 245.200 410.200 ;
        RECT 250.000 401.600 250.800 406.200 ;
        RECT 253.200 401.600 254.000 406.200 ;
        RECT 258.800 401.600 259.600 410.000 ;
        RECT 263.600 401.600 264.400 409.000 ;
        RECT 266.800 401.600 267.600 406.200 ;
        RECT 270.000 401.600 270.800 406.200 ;
        RECT 271.600 401.600 272.400 410.200 ;
        RECT 275.800 401.600 276.600 406.200 ;
        RECT 279.600 401.600 280.400 410.200 ;
        RECT 285.200 401.600 286.000 406.200 ;
        RECT 288.400 401.600 289.200 406.200 ;
        RECT 294.000 401.600 294.800 410.000 ;
        RECT 302.000 401.600 302.800 410.200 ;
        RECT 305.200 401.600 306.000 410.200 ;
        RECT 308.400 401.600 309.200 410.200 ;
        RECT 311.600 401.600 312.400 410.200 ;
        RECT 314.800 401.600 315.600 410.200 ;
        RECT 318.000 401.600 318.800 410.200 ;
        RECT 323.600 401.600 324.400 406.200 ;
        RECT 326.800 401.600 327.600 406.200 ;
        RECT 332.400 401.600 333.200 410.000 ;
        RECT 337.200 401.600 338.000 409.000 ;
        RECT 342.000 401.600 342.800 409.000 ;
        RECT 346.800 401.600 347.600 409.000 ;
        RECT 351.600 401.600 352.400 409.000 ;
        RECT 354.800 401.600 355.600 406.200 ;
        RECT 358.000 401.600 358.800 406.200 ;
        RECT 361.200 401.600 362.000 406.200 ;
        RECT 364.400 401.600 365.200 406.200 ;
        RECT 372.400 401.600 373.200 406.200 ;
        RECT 375.600 401.600 376.400 406.200 ;
        RECT 382.000 401.600 382.800 406.200 ;
        RECT 385.200 401.600 386.000 406.200 ;
        RECT 388.400 401.600 389.200 406.200 ;
        RECT 390.000 401.600 390.800 406.200 ;
        RECT 393.200 401.600 394.000 406.200 ;
        RECT 397.000 401.600 397.800 410.200 ;
        RECT 401.200 401.600 402.000 406.200 ;
        RECT 404.400 401.600 405.200 406.200 ;
        RECT 407.600 401.600 408.400 406.200 ;
        RECT 410.800 401.600 411.600 406.200 ;
        RECT 418.800 401.600 419.600 406.200 ;
        RECT 422.000 401.600 422.800 406.200 ;
        RECT 428.400 401.600 429.200 406.200 ;
        RECT 431.600 401.600 432.400 406.200 ;
        RECT 434.800 401.600 435.600 406.200 ;
        RECT 436.400 401.600 437.200 406.200 ;
        RECT 439.600 401.600 440.400 406.200 ;
        RECT 448.200 401.600 449.000 410.200 ;
        RECT 454.000 401.600 454.800 409.000 ;
        RECT 458.800 401.600 459.600 409.000 ;
        RECT 462.000 401.600 462.800 406.200 ;
        RECT 465.200 401.600 466.000 406.200 ;
        RECT 468.400 401.600 469.200 406.200 ;
        RECT 471.600 401.600 472.400 406.200 ;
        RECT 479.600 401.600 480.400 406.200 ;
        RECT 482.800 401.600 483.600 406.200 ;
        RECT 489.200 401.600 490.000 406.200 ;
        RECT 492.400 401.600 493.200 406.200 ;
        RECT 495.600 401.600 496.400 406.200 ;
        RECT 497.200 401.600 498.000 406.200 ;
        RECT 500.400 401.600 501.200 406.200 ;
        RECT 504.200 401.600 505.000 410.200 ;
        RECT 516.400 409.600 517.200 410.200 ;
        RECT 519.600 410.000 520.600 410.200 ;
        RECT 575.400 410.000 576.200 410.200 ;
        RECT 578.800 409.600 579.600 410.200 ;
        RECT 510.000 401.600 510.800 409.000 ;
        RECT 513.200 401.600 514.000 406.200 ;
        RECT 516.400 401.600 517.200 406.200 ;
        RECT 519.600 401.600 520.400 406.200 ;
        RECT 526.000 401.600 526.800 406.200 ;
        RECT 529.200 401.600 530.000 406.200 ;
        RECT 537.200 401.600 538.000 406.200 ;
        RECT 540.400 401.600 541.200 406.200 ;
        RECT 543.600 401.600 544.400 406.200 ;
        RECT 546.800 401.600 547.600 406.200 ;
        RECT 548.400 401.600 549.200 406.200 ;
        RECT 551.600 401.600 552.400 406.200 ;
        RECT 554.800 401.600 555.600 406.200 ;
        RECT 558.000 401.600 558.800 406.200 ;
        RECT 566.000 401.600 566.800 406.200 ;
        RECT 569.200 401.600 570.000 406.200 ;
        RECT 575.600 401.600 576.400 406.200 ;
        RECT 578.800 401.600 579.600 406.200 ;
        RECT 582.000 401.600 582.800 406.200 ;
        RECT 0.400 400.400 586.800 401.600 ;
        RECT 1.200 391.800 2.000 400.400 ;
        RECT 5.400 395.800 6.200 400.400 ;
        RECT 7.600 395.800 8.400 400.400 ;
        RECT 10.800 395.800 11.600 400.400 ;
        RECT 12.400 395.800 13.200 400.400 ;
        RECT 15.600 395.800 16.400 400.400 ;
        RECT 17.200 395.800 18.000 400.400 ;
        RECT 20.400 395.800 21.200 400.400 ;
        RECT 22.000 395.800 22.800 400.400 ;
        RECT 25.200 395.800 26.000 400.400 ;
        RECT 30.000 391.800 30.800 400.400 ;
        RECT 33.200 393.000 34.000 400.400 ;
        RECT 38.600 395.800 39.400 400.400 ;
        RECT 42.800 391.800 43.600 400.400 ;
        RECT 44.400 395.800 45.200 400.400 ;
        RECT 47.600 395.800 48.400 400.400 ;
        RECT 49.200 395.800 50.000 400.400 ;
        RECT 52.400 395.800 53.200 400.400 ;
        RECT 57.200 391.800 58.000 400.400 ;
        RECT 62.000 393.000 62.800 400.400 ;
        RECT 66.800 393.200 67.800 400.400 ;
        RECT 73.000 399.800 73.800 400.400 ;
        RECT 73.000 393.200 74.000 399.800 ;
        RECT 76.400 395.800 77.200 400.400 ;
        RECT 79.600 391.800 80.400 400.400 ;
        RECT 83.800 395.800 84.600 400.400 ;
        RECT 86.600 395.800 87.400 400.400 ;
        RECT 90.800 391.800 91.600 400.400 ;
        RECT 92.400 395.800 93.200 400.400 ;
        RECT 95.600 395.800 96.400 400.400 ;
        RECT 97.200 395.800 98.000 400.400 ;
        RECT 100.400 395.800 101.200 400.400 ;
        RECT 102.000 395.800 102.800 400.400 ;
        RECT 105.200 395.800 106.000 400.400 ;
        RECT 108.400 395.800 109.200 400.400 ;
        RECT 111.600 395.800 112.400 400.400 ;
        RECT 114.800 391.800 115.600 400.400 ;
        RECT 120.400 395.800 121.200 400.400 ;
        RECT 123.600 395.800 124.400 400.400 ;
        RECT 129.200 392.000 130.000 400.400 ;
        RECT 139.000 399.800 139.800 400.400 ;
        RECT 138.800 393.200 139.800 399.800 ;
        RECT 145.000 393.200 146.000 400.400 ;
        RECT 150.200 399.800 151.000 400.400 ;
        RECT 150.000 393.200 151.000 399.800 ;
        RECT 156.200 393.200 157.200 400.400 ;
        RECT 159.600 391.800 160.400 400.400 ;
        RECT 163.800 395.800 164.600 400.400 ;
        RECT 166.600 395.800 167.400 400.400 ;
        RECT 170.800 391.800 171.600 400.400 ;
        RECT 172.400 395.800 173.200 400.400 ;
        RECT 175.600 395.800 176.400 400.400 ;
        RECT 177.200 391.800 178.000 400.400 ;
        RECT 181.400 395.800 182.200 400.400 ;
        RECT 184.200 395.800 185.000 400.400 ;
        RECT 188.400 391.800 189.200 400.400 ;
        RECT 190.000 395.800 190.800 400.400 ;
        RECT 193.200 395.800 194.000 400.400 ;
        RECT 196.400 391.800 197.200 400.400 ;
        RECT 198.000 391.800 198.800 400.400 ;
        RECT 202.200 395.800 203.000 400.400 ;
        RECT 204.400 391.800 205.200 400.400 ;
        RECT 210.800 393.000 211.600 400.400 ;
        RECT 218.800 391.800 219.600 400.400 ;
        RECT 220.400 395.800 221.200 400.400 ;
        RECT 223.600 395.800 224.400 400.400 ;
        RECT 225.200 395.800 226.000 400.400 ;
        RECT 228.400 395.800 229.200 400.400 ;
        RECT 230.000 395.800 230.800 400.400 ;
        RECT 233.200 391.800 234.000 400.400 ;
        RECT 237.400 395.800 238.200 400.400 ;
        RECT 239.600 395.800 240.400 400.400 ;
        RECT 242.800 395.800 243.600 400.400 ;
        RECT 247.600 393.000 248.400 400.400 ;
        RECT 250.800 391.800 251.600 400.400 ;
        RECT 257.400 399.800 258.200 400.400 ;
        RECT 257.200 393.200 258.200 399.800 ;
        RECT 263.400 393.200 264.400 400.400 ;
        RECT 266.800 395.800 267.600 400.400 ;
        RECT 270.000 395.800 270.800 400.400 ;
        RECT 271.600 395.800 272.400 400.400 ;
        RECT 274.800 395.800 275.600 400.400 ;
        RECT 276.400 391.800 277.200 400.400 ;
        RECT 280.600 395.800 281.400 400.400 ;
        RECT 284.600 399.800 285.400 400.400 ;
        RECT 284.400 393.200 285.400 399.800 ;
        RECT 290.600 393.200 291.600 400.400 ;
        RECT 298.800 391.800 299.600 400.400 ;
        RECT 303.600 395.800 304.400 400.400 ;
        RECT 306.800 395.800 307.600 400.400 ;
        RECT 308.400 395.800 309.200 400.400 ;
        RECT 311.600 395.800 312.400 400.400 ;
        RECT 313.800 395.800 314.600 400.400 ;
        RECT 318.000 391.800 318.800 400.400 ;
        RECT 319.600 391.800 320.400 400.400 ;
        RECT 323.800 395.800 324.600 400.400 ;
        RECT 327.600 395.800 328.400 400.400 ;
        RECT 330.800 391.800 331.600 400.400 ;
        RECT 336.400 395.800 337.200 400.400 ;
        RECT 339.600 395.800 340.400 400.400 ;
        RECT 345.200 392.000 346.000 400.400 ;
        RECT 351.600 391.800 352.400 400.400 ;
        RECT 354.800 393.000 355.600 400.400 ;
        RECT 358.000 391.800 358.800 400.400 ;
        RECT 364.400 391.800 365.200 400.400 ;
        RECT 367.600 393.000 368.400 400.400 ;
        RECT 372.400 393.000 373.200 400.400 ;
        RECT 375.600 391.800 376.400 400.400 ;
        RECT 378.800 391.800 379.600 400.400 ;
        RECT 382.000 391.800 382.800 400.400 ;
        RECT 385.200 391.800 386.000 400.400 ;
        RECT 388.400 391.800 389.200 400.400 ;
        RECT 391.600 391.800 392.400 400.400 ;
        RECT 397.200 395.800 398.000 400.400 ;
        RECT 400.400 395.800 401.200 400.400 ;
        RECT 406.000 392.000 406.800 400.400 ;
        RECT 410.800 393.000 411.600 400.400 ;
        RECT 415.600 393.000 416.400 400.400 ;
        RECT 420.400 393.000 421.200 400.400 ;
        RECT 425.200 393.000 426.000 400.400 ;
        RECT 430.000 393.000 430.800 400.400 ;
        RECT 433.200 395.800 434.000 400.400 ;
        RECT 436.400 395.800 437.200 400.400 ;
        RECT 442.800 395.800 443.600 400.400 ;
        RECT 446.000 395.800 446.800 400.400 ;
        RECT 449.200 395.800 450.000 400.400 ;
        RECT 452.400 395.800 453.200 400.400 ;
        RECT 460.400 395.800 461.200 400.400 ;
        RECT 463.600 395.800 464.400 400.400 ;
        RECT 470.000 395.800 470.800 400.400 ;
        RECT 473.200 395.800 474.000 400.400 ;
        RECT 476.400 395.800 477.200 400.400 ;
        RECT 478.000 395.800 478.800 400.400 ;
        RECT 481.200 395.800 482.000 400.400 ;
        RECT 485.000 391.800 485.800 400.400 ;
        RECT 489.200 395.800 490.000 400.400 ;
        RECT 492.400 395.800 493.200 400.400 ;
        RECT 494.000 391.800 494.800 400.400 ;
        RECT 497.200 393.000 498.000 400.400 ;
        RECT 500.400 391.800 501.200 400.400 ;
        RECT 503.600 393.000 504.400 400.400 ;
        RECT 508.400 393.000 509.200 400.400 ;
        RECT 511.600 395.800 512.400 400.400 ;
        RECT 514.800 395.800 515.600 400.400 ;
        RECT 518.000 395.800 518.800 400.400 ;
        RECT 524.400 395.800 525.200 400.400 ;
        RECT 527.600 395.800 528.400 400.400 ;
        RECT 535.600 395.800 536.400 400.400 ;
        RECT 538.800 395.800 539.600 400.400 ;
        RECT 542.000 395.800 542.800 400.400 ;
        RECT 545.200 395.800 546.000 400.400 ;
        RECT 546.800 395.800 547.600 400.400 ;
        RECT 550.000 395.800 550.800 400.400 ;
        RECT 553.200 395.800 554.000 400.400 ;
        RECT 559.600 395.800 560.400 400.400 ;
        RECT 562.800 395.800 563.600 400.400 ;
        RECT 570.800 395.800 571.600 400.400 ;
        RECT 574.000 395.800 574.800 400.400 ;
        RECT 577.200 395.800 578.000 400.400 ;
        RECT 580.400 395.800 581.200 400.400 ;
        RECT 514.800 391.800 515.600 392.400 ;
        RECT 518.000 391.800 519.000 392.000 ;
        RECT 550.000 391.800 550.800 392.400 ;
        RECT 553.200 391.800 554.200 392.000 ;
        RECT 514.800 391.200 541.800 391.800 ;
        RECT 550.000 391.200 577.000 391.800 ;
        RECT 541.000 391.000 541.800 391.200 ;
        RECT 576.200 391.000 577.000 391.200 ;
        RECT 511.600 373.600 512.400 375.200 ;
        RECT 528.200 370.800 529.000 371.000 ;
        RECT 577.800 370.800 578.600 371.000 ;
        RECT 502.000 370.200 529.000 370.800 ;
        RECT 551.600 370.200 578.600 370.800 ;
        RECT 1.200 361.600 2.000 366.200 ;
        RECT 4.400 361.600 5.200 366.200 ;
        RECT 6.600 361.600 7.400 366.200 ;
        RECT 10.800 361.600 11.600 370.200 ;
        RECT 15.600 361.600 16.400 370.200 ;
        RECT 18.800 361.600 19.600 366.200 ;
        RECT 21.000 361.600 21.800 366.200 ;
        RECT 25.200 361.600 26.000 370.200 ;
        RECT 26.800 361.600 27.600 366.200 ;
        RECT 30.000 361.600 30.800 366.200 ;
        RECT 31.600 361.600 32.400 370.200 ;
        RECT 36.400 361.600 37.200 370.200 ;
        RECT 40.600 361.600 41.400 366.200 ;
        RECT 43.400 361.600 44.200 366.200 ;
        RECT 47.600 361.600 48.400 370.200 ;
        RECT 50.800 361.600 51.600 370.200 ;
        RECT 56.400 361.600 57.200 366.200 ;
        RECT 59.600 361.600 60.400 366.200 ;
        RECT 65.200 361.600 66.000 370.000 ;
        RECT 70.000 361.600 70.800 369.800 ;
        RECT 73.200 361.600 74.000 366.200 ;
        RECT 76.400 361.600 77.200 370.200 ;
        RECT 79.600 361.600 80.400 370.200 ;
        RECT 85.200 361.600 86.000 366.200 ;
        RECT 88.400 361.600 89.200 366.200 ;
        RECT 94.000 361.600 94.800 370.000 ;
        RECT 98.800 361.600 99.600 370.200 ;
        RECT 104.400 361.600 105.200 366.200 ;
        RECT 107.600 361.600 108.400 366.200 ;
        RECT 113.200 361.600 114.000 370.000 ;
        RECT 118.000 361.600 118.800 370.200 ;
        RECT 123.600 361.600 124.400 366.200 ;
        RECT 126.800 361.600 127.600 366.200 ;
        RECT 132.400 361.600 133.200 370.000 ;
        RECT 142.000 361.600 142.800 370.200 ;
        RECT 147.600 361.600 148.400 366.200 ;
        RECT 150.800 361.600 151.600 366.200 ;
        RECT 156.400 361.600 157.200 370.000 ;
        RECT 161.200 361.600 162.200 368.800 ;
        RECT 167.400 362.200 168.400 368.800 ;
        RECT 167.400 361.600 168.200 362.200 ;
        RECT 172.000 361.600 172.800 370.200 ;
        RECT 177.200 361.600 178.000 369.800 ;
        RECT 180.400 361.600 181.200 370.200 ;
        RECT 186.800 361.600 187.600 369.000 ;
        RECT 191.600 361.600 192.400 366.200 ;
        RECT 194.800 361.600 195.600 366.200 ;
        RECT 196.400 361.600 197.200 366.200 ;
        RECT 199.600 361.600 200.400 366.200 ;
        RECT 201.200 361.600 202.000 366.200 ;
        RECT 204.400 361.600 205.200 366.200 ;
        RECT 206.000 361.600 206.800 370.200 ;
        RECT 210.200 361.600 211.000 366.200 ;
        RECT 212.400 361.600 213.200 366.200 ;
        RECT 215.600 361.600 216.400 366.200 ;
        RECT 217.200 361.600 218.000 366.200 ;
        RECT 220.400 361.600 221.200 366.200 ;
        RECT 223.600 361.600 224.400 370.200 ;
        RECT 225.200 361.600 226.000 366.200 ;
        RECT 228.400 361.600 229.200 366.200 ;
        RECT 231.600 362.200 232.600 368.800 ;
        RECT 231.800 361.600 232.600 362.200 ;
        RECT 237.800 361.600 238.800 368.800 ;
        RECT 242.800 361.600 243.600 366.200 ;
        RECT 244.400 361.600 245.200 370.200 ;
        RECT 247.600 361.600 248.400 369.000 ;
        RECT 250.800 361.600 251.600 370.200 ;
        RECT 257.200 361.600 258.000 370.200 ;
        RECT 258.800 361.600 259.600 366.200 ;
        RECT 262.000 361.600 262.800 366.200 ;
        RECT 264.200 361.600 265.000 366.200 ;
        RECT 268.400 361.600 269.200 370.200 ;
        RECT 273.200 361.600 274.000 369.000 ;
        RECT 278.000 361.600 278.800 366.200 ;
        RECT 279.600 361.600 280.400 370.200 ;
        RECT 283.800 361.600 284.600 366.200 ;
        RECT 286.000 361.600 286.800 366.200 ;
        RECT 289.200 361.600 290.000 366.200 ;
        RECT 297.200 361.600 298.000 369.000 ;
        RECT 300.400 361.600 301.200 370.200 ;
        RECT 302.000 361.600 302.800 366.200 ;
        RECT 305.200 361.600 306.000 370.200 ;
        RECT 309.400 361.600 310.200 366.200 ;
        RECT 313.200 361.600 314.000 370.200 ;
        RECT 318.800 361.600 319.600 366.200 ;
        RECT 322.000 361.600 322.800 366.200 ;
        RECT 327.600 361.600 328.400 370.000 ;
        RECT 332.400 361.600 333.200 370.200 ;
        RECT 338.000 361.600 338.800 366.200 ;
        RECT 341.200 361.600 342.000 366.200 ;
        RECT 346.800 361.600 347.600 370.000 ;
        RECT 350.000 361.600 350.800 370.200 ;
        RECT 354.200 361.600 355.000 366.200 ;
        RECT 358.000 361.600 358.800 369.000 ;
        RECT 361.200 361.600 362.000 370.200 ;
        RECT 365.400 361.600 366.200 366.200 ;
        RECT 370.800 361.600 371.600 370.200 ;
        RECT 372.400 361.600 373.200 370.200 ;
        RECT 377.800 361.600 378.600 366.200 ;
        RECT 382.000 361.600 382.800 370.200 ;
        RECT 385.200 361.600 386.000 366.200 ;
        RECT 388.400 361.600 389.200 370.200 ;
        RECT 394.000 361.600 394.800 366.200 ;
        RECT 397.200 361.600 398.000 366.200 ;
        RECT 402.800 361.600 403.600 370.000 ;
        RECT 406.000 361.600 406.800 370.200 ;
        RECT 409.200 361.600 410.000 370.200 ;
        RECT 410.800 361.600 411.600 366.200 ;
        RECT 414.000 361.600 414.800 366.200 ;
        RECT 417.200 361.600 418.000 366.200 ;
        RECT 420.400 361.600 421.200 366.200 ;
        RECT 428.400 361.600 429.200 366.200 ;
        RECT 431.600 361.600 432.400 366.200 ;
        RECT 438.000 361.600 438.800 366.200 ;
        RECT 441.200 361.600 442.000 366.200 ;
        RECT 444.400 361.600 445.200 366.200 ;
        RECT 453.000 361.600 453.800 370.200 ;
        RECT 457.200 361.600 458.000 366.200 ;
        RECT 460.400 361.600 461.200 366.200 ;
        RECT 463.600 361.600 464.400 366.200 ;
        RECT 466.800 361.600 467.600 366.200 ;
        RECT 474.800 361.600 475.600 366.200 ;
        RECT 478.000 361.600 478.800 366.200 ;
        RECT 484.400 361.600 485.200 366.200 ;
        RECT 487.600 361.600 488.400 366.200 ;
        RECT 490.800 361.600 491.600 366.200 ;
        RECT 494.600 361.600 495.400 370.200 ;
        RECT 502.000 369.600 502.800 370.200 ;
        RECT 505.400 370.000 506.200 370.200 ;
        RECT 498.800 361.600 499.600 366.200 ;
        RECT 502.000 361.600 502.800 366.200 ;
        RECT 505.200 361.600 506.000 366.200 ;
        RECT 511.600 361.600 512.400 366.200 ;
        RECT 514.800 361.600 515.600 366.200 ;
        RECT 522.800 361.600 523.600 366.200 ;
        RECT 526.000 361.600 526.800 366.200 ;
        RECT 529.200 361.600 530.000 366.200 ;
        RECT 532.400 361.600 533.200 366.200 ;
        RECT 534.000 361.600 534.800 370.200 ;
        RECT 537.200 361.600 538.000 370.200 ;
        RECT 540.400 361.600 541.200 370.200 ;
        RECT 543.600 361.600 544.400 369.000 ;
        RECT 546.800 361.600 547.600 370.200 ;
        RECT 551.600 369.600 552.400 370.200 ;
        RECT 554.800 370.000 555.800 370.200 ;
        RECT 548.400 361.600 549.200 366.200 ;
        RECT 551.600 361.600 552.400 366.200 ;
        RECT 554.800 361.600 555.600 366.200 ;
        RECT 561.200 361.600 562.000 366.200 ;
        RECT 564.400 361.600 565.200 366.200 ;
        RECT 572.400 361.600 573.200 366.200 ;
        RECT 575.600 361.600 576.400 366.200 ;
        RECT 578.800 361.600 579.600 366.200 ;
        RECT 582.000 361.600 582.800 366.200 ;
        RECT 0.400 360.400 586.800 361.600 ;
        RECT 1.800 355.800 2.600 360.400 ;
        RECT 6.000 351.800 6.800 360.400 ;
        RECT 9.400 359.800 10.200 360.400 ;
        RECT 9.200 353.200 10.200 359.800 ;
        RECT 15.400 353.200 16.400 360.400 ;
        RECT 18.800 355.800 19.600 360.400 ;
        RECT 23.800 359.800 24.600 360.400 ;
        RECT 23.600 353.200 24.600 359.800 ;
        RECT 29.800 353.200 30.800 360.400 ;
        RECT 33.200 355.800 34.000 360.400 ;
        RECT 39.000 351.800 39.800 360.400 ;
        RECT 46.000 353.000 46.800 360.400 ;
        RECT 49.800 355.800 50.600 360.400 ;
        RECT 54.000 351.800 54.800 360.400 ;
        RECT 55.600 351.800 56.400 360.400 ;
        RECT 59.800 355.800 60.600 360.400 ;
        RECT 63.600 353.000 64.400 360.400 ;
        RECT 71.600 351.800 72.400 360.400 ;
        RECT 73.200 351.800 74.000 360.400 ;
        RECT 79.600 353.000 80.400 360.400 ;
        RECT 84.400 351.800 85.200 360.400 ;
        RECT 89.200 355.800 90.000 360.400 ;
        RECT 92.400 355.800 93.200 360.400 ;
        RECT 95.600 351.800 96.400 360.400 ;
        RECT 101.200 355.800 102.000 360.400 ;
        RECT 104.400 355.800 105.200 360.400 ;
        RECT 110.000 352.000 110.800 360.400 ;
        RECT 113.200 355.800 114.000 360.400 ;
        RECT 116.400 355.800 117.200 360.400 ;
        RECT 119.600 351.800 120.400 360.400 ;
        RECT 123.000 359.800 123.800 360.400 ;
        RECT 122.800 353.200 123.800 359.800 ;
        RECT 129.000 353.200 130.000 360.400 ;
        RECT 132.400 355.800 133.200 360.400 ;
        RECT 135.600 355.800 136.400 360.400 ;
        RECT 143.800 359.800 144.600 360.400 ;
        RECT 143.600 353.200 144.600 359.800 ;
        RECT 149.800 353.200 150.800 360.400 ;
        RECT 154.800 351.800 155.600 360.400 ;
        RECT 160.400 355.800 161.200 360.400 ;
        RECT 163.600 355.800 164.400 360.400 ;
        RECT 169.200 352.000 170.000 360.400 ;
        RECT 174.000 351.800 174.800 360.400 ;
        RECT 179.600 355.800 180.400 360.400 ;
        RECT 182.800 355.800 183.600 360.400 ;
        RECT 188.400 352.000 189.200 360.400 ;
        RECT 194.800 351.800 195.600 360.400 ;
        RECT 198.200 359.800 199.000 360.400 ;
        RECT 198.000 353.200 199.000 359.800 ;
        RECT 204.200 353.200 205.200 360.400 ;
        RECT 207.600 351.800 208.400 360.400 ;
        RECT 214.000 351.800 214.800 360.400 ;
        RECT 218.800 353.000 219.600 360.400 ;
        RECT 223.800 359.800 224.600 360.400 ;
        RECT 223.600 353.200 224.600 359.800 ;
        RECT 229.800 353.200 230.800 360.400 ;
        RECT 233.800 355.800 234.600 360.400 ;
        RECT 238.000 351.800 238.800 360.400 ;
        RECT 239.600 355.800 240.400 360.400 ;
        RECT 242.800 355.800 243.600 360.400 ;
        RECT 244.400 355.800 245.200 360.400 ;
        RECT 247.600 355.800 248.400 360.400 ;
        RECT 249.200 351.800 250.000 360.400 ;
        RECT 252.400 351.800 253.200 360.400 ;
        RECT 254.000 351.800 254.800 360.400 ;
        RECT 257.200 351.800 258.000 360.400 ;
        RECT 260.400 351.800 261.200 360.400 ;
        RECT 263.600 351.800 264.400 360.400 ;
        RECT 267.000 359.800 267.800 360.400 ;
        RECT 266.800 353.200 267.800 359.800 ;
        RECT 273.000 353.200 274.000 360.400 ;
        RECT 276.400 351.800 277.200 360.400 ;
        RECT 280.600 355.800 281.400 360.400 ;
        RECT 282.800 355.800 283.600 360.400 ;
        RECT 286.000 355.800 286.800 360.400 ;
        RECT 294.000 353.000 294.800 360.400 ;
        RECT 302.000 351.800 302.800 360.400 ;
        RECT 305.800 351.800 306.600 360.400 ;
        RECT 310.000 351.800 310.800 360.400 ;
        RECT 314.800 355.800 315.600 360.400 ;
        RECT 321.200 351.800 322.000 360.400 ;
        RECT 323.400 355.800 324.200 360.400 ;
        RECT 327.600 351.800 328.400 360.400 ;
        RECT 330.800 355.800 331.600 360.400 ;
        RECT 334.000 351.800 334.800 360.400 ;
        RECT 339.600 355.800 340.400 360.400 ;
        RECT 342.800 355.800 343.600 360.400 ;
        RECT 348.400 352.000 349.200 360.400 ;
        RECT 353.200 355.800 354.000 360.400 ;
        RECT 356.400 351.800 357.200 360.400 ;
        RECT 362.000 355.800 362.800 360.400 ;
        RECT 365.200 355.800 366.000 360.400 ;
        RECT 370.800 352.000 371.600 360.400 ;
        RECT 375.600 353.000 376.400 360.400 ;
        RECT 380.600 359.800 381.400 360.400 ;
        RECT 380.400 353.200 381.400 359.800 ;
        RECT 386.600 353.200 387.600 360.400 ;
        RECT 391.600 351.800 392.400 360.400 ;
        RECT 394.800 351.800 395.600 360.400 ;
        RECT 400.400 355.800 401.200 360.400 ;
        RECT 403.600 355.800 404.400 360.400 ;
        RECT 409.200 352.000 410.000 360.400 ;
        RECT 413.000 355.800 413.800 360.400 ;
        RECT 417.200 351.800 418.000 360.400 ;
        RECT 419.400 355.800 420.200 360.400 ;
        RECT 423.600 351.800 424.400 360.400 ;
        RECT 425.200 351.800 426.000 360.400 ;
        RECT 429.400 355.800 430.200 360.400 ;
        RECT 432.200 355.800 433.000 360.400 ;
        RECT 436.400 351.800 437.200 360.400 ;
        RECT 439.600 355.800 440.400 360.400 ;
        RECT 442.800 355.800 443.600 360.400 ;
        RECT 449.200 351.800 450.000 360.400 ;
        RECT 454.000 355.800 454.800 360.400 ;
        RECT 457.200 355.800 458.000 360.400 ;
        RECT 462.000 353.000 462.800 360.400 ;
        RECT 465.200 355.800 466.000 360.400 ;
        RECT 468.400 355.800 469.200 360.400 ;
        RECT 471.600 353.200 472.600 360.400 ;
        RECT 477.800 359.800 478.600 360.400 ;
        RECT 477.800 353.200 478.800 359.800 ;
        RECT 482.800 351.800 483.600 360.400 ;
        RECT 488.400 355.800 489.200 360.400 ;
        RECT 491.600 355.800 492.400 360.400 ;
        RECT 497.200 352.000 498.000 360.400 ;
        RECT 500.400 351.800 501.200 360.400 ;
        RECT 503.600 351.800 504.400 360.400 ;
        RECT 506.800 351.800 507.600 360.400 ;
        RECT 510.000 351.800 510.800 360.400 ;
        RECT 513.200 351.800 514.000 360.400 ;
        RECT 514.800 355.800 515.600 360.400 ;
        RECT 518.000 355.800 518.800 360.400 ;
        RECT 521.200 355.800 522.000 360.400 ;
        RECT 527.600 355.800 528.400 360.400 ;
        RECT 530.800 355.800 531.600 360.400 ;
        RECT 538.800 355.800 539.600 360.400 ;
        RECT 542.000 355.800 542.800 360.400 ;
        RECT 545.200 355.800 546.000 360.400 ;
        RECT 548.400 355.800 549.200 360.400 ;
        RECT 550.000 355.800 550.800 360.400 ;
        RECT 553.200 355.800 554.000 360.400 ;
        RECT 556.400 355.800 557.200 360.400 ;
        RECT 562.800 355.800 563.600 360.400 ;
        RECT 566.000 355.800 566.800 360.400 ;
        RECT 574.000 355.800 574.800 360.400 ;
        RECT 577.200 355.800 578.000 360.400 ;
        RECT 580.400 355.800 581.200 360.400 ;
        RECT 583.600 355.800 584.400 360.400 ;
        RECT 518.000 351.800 518.800 352.400 ;
        RECT 521.200 351.800 522.200 352.000 ;
        RECT 553.200 351.800 554.000 352.400 ;
        RECT 556.600 351.800 557.400 352.000 ;
        RECT 518.000 351.200 545.000 351.800 ;
        RECT 553.200 351.200 580.200 351.800 ;
        RECT 544.200 351.000 545.000 351.200 ;
        RECT 579.400 351.000 580.200 351.200 ;
        RECT 514.800 331.600 515.600 333.200 ;
        RECT 523.800 330.800 524.600 331.000 ;
        RECT 523.800 330.200 550.800 330.800 ;
        RECT 2.800 322.200 3.800 328.800 ;
        RECT 3.000 321.600 3.800 322.200 ;
        RECT 9.000 321.600 10.000 328.800 ;
        RECT 12.400 321.600 13.200 330.200 ;
        RECT 15.600 321.600 16.400 330.200 ;
        RECT 18.800 321.600 19.600 330.200 ;
        RECT 20.400 321.600 21.200 330.200 ;
        RECT 23.600 321.600 24.400 329.000 ;
        RECT 26.800 321.600 27.600 326.200 ;
        RECT 31.600 321.600 32.400 329.000 ;
        RECT 34.800 321.600 35.600 330.200 ;
        RECT 38.000 321.600 38.800 329.000 ;
        RECT 45.000 321.600 45.800 326.200 ;
        RECT 49.200 321.600 50.000 330.200 ;
        RECT 52.400 321.600 53.200 325.800 ;
        RECT 55.600 321.600 56.400 326.200 ;
        RECT 58.800 321.600 59.600 326.200 ;
        RECT 60.400 321.600 61.200 326.200 ;
        RECT 63.600 321.600 64.400 326.200 ;
        RECT 66.800 321.600 67.600 326.200 ;
        RECT 70.000 321.600 70.800 325.800 ;
        RECT 73.200 321.600 74.000 326.200 ;
        RECT 75.400 321.600 76.200 326.200 ;
        RECT 79.600 321.600 80.400 330.200 ;
        RECT 81.200 321.600 82.000 326.200 ;
        RECT 84.400 321.600 85.200 326.200 ;
        RECT 86.000 321.600 86.800 326.200 ;
        RECT 89.200 321.600 90.000 326.200 ;
        RECT 91.400 321.600 92.200 326.200 ;
        RECT 95.600 321.600 96.400 330.200 ;
        RECT 97.800 321.600 98.600 326.200 ;
        RECT 102.000 321.600 102.800 330.200 ;
        RECT 103.600 321.600 104.400 330.200 ;
        RECT 108.400 321.600 109.200 330.200 ;
        RECT 112.600 321.600 113.400 326.200 ;
        RECT 116.400 321.600 117.200 326.200 ;
        RECT 118.000 321.600 118.800 330.200 ;
        RECT 124.400 321.600 125.200 330.200 ;
        RECT 126.000 321.600 126.800 330.200 ;
        RECT 130.200 321.600 131.000 326.200 ;
        RECT 133.000 321.600 133.800 326.200 ;
        RECT 137.200 321.600 138.000 330.200 ;
        RECT 145.200 322.200 146.200 328.800 ;
        RECT 145.400 321.600 146.200 322.200 ;
        RECT 151.400 321.600 152.400 328.800 ;
        RECT 156.400 321.600 157.200 329.000 ;
        RECT 162.800 321.600 163.600 326.200 ;
        RECT 164.400 321.600 165.200 326.200 ;
        RECT 168.200 321.600 169.000 326.200 ;
        RECT 172.400 321.600 173.200 330.200 ;
        RECT 175.600 321.600 176.600 328.800 ;
        RECT 181.800 322.200 182.800 328.800 ;
        RECT 181.800 321.600 182.600 322.200 ;
        RECT 185.200 321.600 186.000 330.200 ;
        RECT 188.400 321.600 189.200 330.200 ;
        RECT 191.600 321.600 192.400 330.200 ;
        RECT 194.800 321.600 195.600 330.200 ;
        RECT 198.000 321.600 198.800 330.200 ;
        RECT 201.200 321.600 202.000 330.200 ;
        RECT 206.800 321.600 207.600 326.200 ;
        RECT 210.000 321.600 210.800 326.200 ;
        RECT 215.600 321.600 216.400 330.000 ;
        RECT 220.400 321.600 221.400 328.800 ;
        RECT 226.600 322.200 227.600 328.800 ;
        RECT 226.600 321.600 227.400 322.200 ;
        RECT 231.600 321.600 232.600 328.800 ;
        RECT 237.800 322.200 238.800 328.800 ;
        RECT 237.800 321.600 238.600 322.200 ;
        RECT 241.800 321.600 242.600 326.200 ;
        RECT 246.000 321.600 246.800 330.200 ;
        RECT 247.600 321.600 248.400 326.200 ;
        RECT 250.800 321.600 251.600 326.200 ;
        RECT 252.400 321.600 253.200 326.200 ;
        RECT 255.600 321.600 256.400 325.800 ;
        RECT 258.800 321.600 259.600 326.200 ;
        RECT 262.000 321.600 262.800 326.200 ;
        RECT 265.200 321.600 266.000 329.000 ;
        RECT 270.000 321.600 270.800 330.200 ;
        RECT 274.800 321.600 275.600 330.200 ;
        RECT 279.000 321.600 279.800 326.200 ;
        RECT 281.200 321.600 282.000 326.200 ;
        RECT 286.000 321.600 286.800 329.000 ;
        RECT 298.800 321.600 299.600 330.200 ;
        RECT 300.400 321.600 301.200 330.200 ;
        RECT 304.600 321.600 305.400 326.200 ;
        RECT 306.800 321.600 307.600 326.200 ;
        RECT 310.000 321.600 310.800 326.200 ;
        RECT 314.800 321.600 315.600 329.000 ;
        RECT 318.000 321.600 318.800 330.200 ;
        RECT 324.400 322.200 325.400 328.800 ;
        RECT 324.600 321.600 325.400 322.200 ;
        RECT 330.600 321.600 331.600 328.800 ;
        RECT 335.600 321.600 336.400 330.200 ;
        RECT 341.200 321.600 342.000 326.200 ;
        RECT 344.400 321.600 345.200 326.200 ;
        RECT 350.000 321.600 350.800 330.000 ;
        RECT 354.800 321.600 355.600 326.200 ;
        RECT 358.000 321.600 358.800 330.200 ;
        RECT 363.600 321.600 364.400 326.200 ;
        RECT 366.800 321.600 367.600 326.200 ;
        RECT 372.400 321.600 373.200 330.000 ;
        RECT 375.600 321.600 376.400 330.200 ;
        RECT 382.000 321.600 382.800 330.200 ;
        RECT 384.200 321.600 385.000 326.200 ;
        RECT 388.400 321.600 389.200 330.200 ;
        RECT 390.000 321.600 390.800 326.200 ;
        RECT 393.200 321.600 394.000 326.200 ;
        RECT 396.400 321.600 397.200 330.200 ;
        RECT 402.000 321.600 402.800 326.200 ;
        RECT 405.200 321.600 406.000 326.200 ;
        RECT 410.800 321.600 411.600 330.000 ;
        RECT 415.600 321.600 416.400 330.200 ;
        RECT 421.200 321.600 422.000 326.200 ;
        RECT 424.400 321.600 425.200 326.200 ;
        RECT 430.000 321.600 430.800 330.000 ;
        RECT 434.800 322.200 435.800 328.800 ;
        RECT 435.000 321.600 435.800 322.200 ;
        RECT 441.000 321.600 442.000 328.800 ;
        RECT 450.800 321.600 451.600 329.000 ;
        RECT 454.000 321.600 454.800 330.200 ;
        RECT 458.200 321.600 459.000 326.200 ;
        RECT 463.600 321.600 464.400 330.200 ;
        RECT 465.200 321.600 466.000 326.200 ;
        RECT 468.400 321.600 469.200 326.200 ;
        RECT 470.000 321.600 470.800 330.200 ;
        RECT 474.200 321.600 475.000 326.200 ;
        RECT 478.000 321.600 478.800 330.000 ;
        RECT 483.600 321.600 484.400 326.200 ;
        RECT 486.800 321.600 487.600 326.200 ;
        RECT 492.400 321.600 493.200 330.200 ;
        RECT 497.200 321.600 498.000 330.000 ;
        RECT 502.800 321.600 503.600 326.200 ;
        RECT 506.000 321.600 506.800 326.200 ;
        RECT 511.600 321.600 512.400 330.200 ;
        RECT 546.600 330.000 547.400 330.200 ;
        RECT 550.000 329.600 550.800 330.200 ;
        RECT 516.400 321.600 517.200 329.000 ;
        RECT 519.600 321.600 520.400 326.200 ;
        RECT 522.800 321.600 523.600 326.200 ;
        RECT 526.000 321.600 526.800 326.200 ;
        RECT 529.200 321.600 530.000 326.200 ;
        RECT 537.200 321.600 538.000 326.200 ;
        RECT 540.400 321.600 541.200 326.200 ;
        RECT 546.800 321.600 547.600 326.200 ;
        RECT 550.000 321.600 550.800 326.200 ;
        RECT 553.200 321.600 554.000 326.200 ;
        RECT 556.400 321.600 557.200 330.200 ;
        RECT 562.000 321.600 562.800 326.200 ;
        RECT 565.200 321.600 566.000 326.200 ;
        RECT 570.800 321.600 571.600 330.000 ;
        RECT 575.600 321.600 576.400 329.000 ;
        RECT 580.400 321.600 581.200 329.000 ;
        RECT 0.400 320.400 586.800 321.600 ;
        RECT 1.800 315.800 2.600 320.400 ;
        RECT 6.000 311.800 6.800 320.400 ;
        RECT 7.600 311.800 8.400 320.400 ;
        RECT 12.400 311.800 13.200 320.400 ;
        RECT 17.200 311.800 18.000 320.400 ;
        RECT 23.600 311.800 24.400 320.400 ;
        RECT 25.800 315.800 26.600 320.400 ;
        RECT 30.000 311.800 30.800 320.400 ;
        RECT 31.600 315.800 32.400 320.400 ;
        RECT 34.800 315.800 35.600 320.400 ;
        RECT 39.600 311.800 40.400 320.400 ;
        RECT 41.200 315.800 42.000 320.400 ;
        RECT 44.400 315.800 45.200 320.400 ;
        RECT 46.600 315.800 47.400 320.400 ;
        RECT 50.800 311.800 51.600 320.400 ;
        RECT 54.200 319.800 55.000 320.400 ;
        RECT 54.000 313.200 55.000 319.800 ;
        RECT 60.200 313.200 61.200 320.400 ;
        RECT 63.600 315.800 64.400 320.400 ;
        RECT 66.800 315.800 67.600 320.400 ;
        RECT 68.400 315.800 69.200 320.400 ;
        RECT 73.200 313.000 74.000 320.400 ;
        RECT 76.400 311.800 77.200 320.400 ;
        RECT 82.800 313.000 83.600 320.400 ;
        RECT 86.000 315.800 86.800 320.400 ;
        RECT 89.200 315.800 90.000 320.400 ;
        RECT 92.400 315.800 93.200 320.400 ;
        RECT 94.000 311.800 94.800 320.400 ;
        RECT 98.200 315.800 99.000 320.400 ;
        RECT 100.400 311.800 101.200 320.400 ;
        RECT 105.200 311.800 106.000 320.400 ;
        RECT 109.400 315.800 110.200 320.400 ;
        RECT 113.200 313.000 114.000 320.400 ;
        RECT 118.000 311.800 118.800 320.400 ;
        RECT 122.200 315.800 123.000 320.400 ;
        RECT 124.400 315.800 125.200 320.400 ;
        RECT 127.600 315.800 128.400 320.400 ;
        RECT 130.800 315.800 131.600 320.400 ;
        RECT 134.000 315.800 134.800 320.400 ;
        RECT 141.000 315.800 141.800 320.400 ;
        RECT 145.200 311.800 146.000 320.400 ;
        RECT 146.800 315.800 147.600 320.400 ;
        RECT 150.000 315.800 150.800 320.400 ;
        RECT 152.200 315.800 153.000 320.400 ;
        RECT 156.400 311.800 157.200 320.400 ;
        RECT 161.200 311.800 162.000 320.400 ;
        RECT 165.000 311.800 165.800 320.400 ;
        RECT 172.400 311.800 173.200 320.400 ;
        RECT 174.000 315.800 174.800 320.400 ;
        RECT 177.200 312.200 178.000 320.400 ;
        RECT 182.000 311.800 182.800 320.400 ;
        RECT 187.600 315.800 188.400 320.400 ;
        RECT 190.800 315.800 191.600 320.400 ;
        RECT 196.400 312.000 197.200 320.400 ;
        RECT 201.200 311.800 202.000 320.400 ;
        RECT 206.800 315.800 207.600 320.400 ;
        RECT 210.000 315.800 210.800 320.400 ;
        RECT 215.600 312.000 216.400 320.400 ;
        RECT 220.400 313.000 221.200 320.400 ;
        RECT 225.200 313.000 226.000 320.400 ;
        RECT 229.000 315.800 229.800 320.400 ;
        RECT 233.200 311.800 234.000 320.400 ;
        RECT 235.400 315.800 236.200 320.400 ;
        RECT 239.600 311.800 240.400 320.400 ;
        RECT 244.400 313.000 245.200 320.400 ;
        RECT 249.200 315.800 250.000 320.400 ;
        RECT 250.800 311.800 251.600 320.400 ;
        RECT 255.000 315.800 255.800 320.400 ;
        RECT 258.400 311.800 259.200 320.400 ;
        RECT 263.600 312.200 264.400 320.400 ;
        RECT 266.800 311.800 267.600 320.400 ;
        RECT 270.000 313.000 270.800 320.400 ;
        RECT 274.800 311.800 275.600 320.400 ;
        RECT 280.400 315.800 281.200 320.400 ;
        RECT 283.600 315.800 284.400 320.400 ;
        RECT 289.200 312.000 290.000 320.400 ;
        RECT 298.800 311.800 299.600 320.400 ;
        RECT 304.400 315.800 305.200 320.400 ;
        RECT 307.600 315.800 308.400 320.400 ;
        RECT 313.200 312.000 314.000 320.400 ;
        RECT 318.000 313.000 318.800 320.400 ;
        RECT 321.200 311.800 322.000 320.400 ;
        RECT 322.800 315.800 323.600 320.400 ;
        RECT 326.000 315.800 326.800 320.400 ;
        RECT 327.600 315.800 328.400 320.400 ;
        RECT 330.800 315.800 331.600 320.400 ;
        RECT 333.000 315.800 333.800 320.400 ;
        RECT 337.200 311.800 338.000 320.400 ;
        RECT 339.400 315.800 340.200 320.400 ;
        RECT 343.600 311.800 344.400 320.400 ;
        RECT 345.800 315.800 346.600 320.400 ;
        RECT 350.000 311.800 350.800 320.400 ;
        RECT 353.200 315.800 354.000 320.400 ;
        RECT 356.400 313.200 357.400 320.400 ;
        RECT 362.600 319.800 363.400 320.400 ;
        RECT 367.800 319.800 368.600 320.400 ;
        RECT 362.600 313.200 363.600 319.800 ;
        RECT 367.600 313.200 368.600 319.800 ;
        RECT 373.800 313.200 374.800 320.400 ;
        RECT 377.200 315.800 378.000 320.400 ;
        RECT 380.400 315.800 381.200 320.400 ;
        RECT 382.000 311.800 382.800 320.400 ;
        RECT 386.800 311.800 387.600 320.400 ;
        RECT 393.200 311.800 394.000 320.400 ;
        RECT 396.400 315.800 397.200 320.400 ;
        RECT 400.200 311.800 401.000 320.400 ;
        RECT 406.000 311.800 406.800 320.400 ;
        RECT 411.600 315.800 412.400 320.400 ;
        RECT 414.800 315.800 415.600 320.400 ;
        RECT 420.400 312.000 421.200 320.400 ;
        RECT 428.400 313.000 429.200 320.400 ;
        RECT 431.600 315.800 432.400 320.400 ;
        RECT 435.400 315.800 436.200 320.400 ;
        RECT 439.600 311.800 440.400 320.400 ;
        RECT 441.200 315.800 442.000 320.400 ;
        RECT 444.400 315.800 445.200 320.400 ;
        RECT 450.800 315.800 451.600 320.400 ;
        RECT 454.000 315.800 454.800 320.400 ;
        RECT 456.200 315.800 457.000 320.400 ;
        RECT 460.400 311.800 461.200 320.400 ;
        RECT 463.600 315.800 464.400 320.400 ;
        RECT 466.800 313.200 467.800 320.400 ;
        RECT 473.000 319.800 473.800 320.400 ;
        RECT 473.000 313.200 474.000 319.800 ;
        RECT 478.000 315.800 478.800 320.400 ;
        RECT 481.200 312.000 482.000 320.400 ;
        RECT 486.800 315.800 487.600 320.400 ;
        RECT 490.000 315.800 490.800 320.400 ;
        RECT 495.600 311.800 496.400 320.400 ;
        RECT 498.800 315.800 499.600 320.400 ;
        RECT 502.000 315.800 502.800 320.400 ;
        RECT 505.200 315.800 506.000 320.400 ;
        RECT 508.400 315.800 509.200 320.400 ;
        RECT 516.400 315.800 517.200 320.400 ;
        RECT 519.600 315.800 520.400 320.400 ;
        RECT 526.000 315.800 526.800 320.400 ;
        RECT 529.200 315.800 530.000 320.400 ;
        RECT 532.400 315.800 533.200 320.400 ;
        RECT 534.000 315.800 534.800 320.400 ;
        RECT 537.200 315.800 538.000 320.400 ;
        RECT 541.000 311.800 541.800 320.400 ;
        RECT 546.800 312.000 547.600 320.400 ;
        RECT 552.400 315.800 553.200 320.400 ;
        RECT 555.600 315.800 556.400 320.400 ;
        RECT 561.200 311.800 562.000 320.400 ;
        RECT 566.000 312.000 566.800 320.400 ;
        RECT 571.600 315.800 572.400 320.400 ;
        RECT 574.800 315.800 575.600 320.400 ;
        RECT 580.400 311.800 581.200 320.400 ;
        RECT 1.200 281.600 2.000 286.200 ;
        RECT 6.000 281.600 6.800 286.200 ;
        RECT 8.200 281.600 9.000 286.200 ;
        RECT 12.400 281.600 13.200 290.200 ;
        RECT 15.600 281.600 16.400 285.800 ;
        RECT 18.800 281.600 19.600 286.200 ;
        RECT 20.400 281.600 21.200 290.200 ;
        RECT 24.600 281.600 25.400 286.200 ;
        RECT 28.400 281.600 29.200 286.200 ;
        RECT 30.600 281.600 31.400 286.200 ;
        RECT 34.800 281.600 35.600 290.200 ;
        RECT 39.600 281.600 40.400 289.000 ;
        RECT 44.400 281.600 45.200 289.000 ;
        RECT 50.800 281.600 51.600 290.200 ;
        RECT 55.000 281.600 55.800 286.200 ;
        RECT 57.800 281.600 58.600 286.200 ;
        RECT 62.000 281.600 62.800 290.200 ;
        RECT 63.600 281.600 64.400 290.200 ;
        RECT 67.800 281.600 68.600 286.200 ;
        RECT 70.000 281.600 70.800 286.200 ;
        RECT 73.200 281.600 74.000 286.200 ;
        RECT 78.000 281.600 78.800 290.200 ;
        RECT 84.400 281.600 85.200 289.000 ;
        RECT 87.600 281.600 88.400 286.200 ;
        RECT 90.800 281.600 91.600 286.200 ;
        RECT 94.000 281.600 95.000 288.800 ;
        RECT 100.200 282.200 101.200 288.800 ;
        RECT 100.200 281.600 101.000 282.200 ;
        RECT 105.200 281.600 106.000 290.200 ;
        RECT 106.800 281.600 107.600 290.200 ;
        RECT 111.000 281.600 111.800 286.200 ;
        RECT 113.200 281.600 114.000 286.200 ;
        RECT 119.600 281.600 120.400 289.000 ;
        RECT 123.400 281.600 124.200 286.200 ;
        RECT 127.600 281.600 128.400 290.200 ;
        RECT 129.200 281.600 130.000 286.200 ;
        RECT 132.400 281.600 133.200 286.200 ;
        RECT 134.000 281.600 134.800 286.200 ;
        RECT 137.200 281.600 138.000 286.200 ;
        RECT 143.600 281.600 144.400 286.200 ;
        RECT 146.800 281.600 147.600 286.200 ;
        RECT 151.600 281.600 152.400 290.200 ;
        RECT 154.800 281.600 155.600 289.000 ;
        RECT 159.600 281.600 160.400 290.200 ;
        RECT 163.800 281.600 164.600 286.200 ;
        RECT 167.600 281.600 168.400 286.200 ;
        RECT 172.400 281.600 173.200 289.000 ;
        RECT 178.800 281.600 179.600 290.200 ;
        RECT 180.400 281.600 181.200 290.200 ;
        RECT 184.600 281.600 185.400 286.200 ;
        RECT 188.400 282.200 189.400 288.800 ;
        RECT 188.600 281.600 189.400 282.200 ;
        RECT 194.600 281.600 195.600 288.800 ;
        RECT 199.600 281.600 200.400 290.200 ;
        RECT 205.200 281.600 206.000 286.200 ;
        RECT 208.400 281.600 209.200 286.200 ;
        RECT 214.000 281.600 214.800 290.000 ;
        RECT 218.800 281.600 219.600 289.000 ;
        RECT 223.600 281.600 224.400 289.000 ;
        RECT 228.400 281.600 229.200 290.000 ;
        RECT 234.000 281.600 234.800 286.200 ;
        RECT 237.200 281.600 238.000 286.200 ;
        RECT 242.800 281.600 243.600 290.200 ;
        RECT 247.600 281.600 248.600 288.800 ;
        RECT 253.800 282.200 254.800 288.800 ;
        RECT 253.800 281.600 254.600 282.200 ;
        RECT 258.800 281.600 259.600 290.200 ;
        RECT 264.400 281.600 265.200 286.200 ;
        RECT 267.600 281.600 268.400 286.200 ;
        RECT 273.200 281.600 274.000 290.000 ;
        RECT 278.000 281.600 278.800 290.200 ;
        RECT 283.600 281.600 284.400 286.200 ;
        RECT 286.800 281.600 287.600 286.200 ;
        RECT 292.400 281.600 293.200 290.000 ;
        RECT 300.400 281.600 301.200 286.200 ;
        RECT 303.600 281.600 304.400 286.200 ;
        RECT 306.800 281.600 307.800 288.800 ;
        RECT 313.000 282.200 314.000 288.800 ;
        RECT 313.000 281.600 313.800 282.200 ;
        RECT 317.000 281.600 317.800 286.200 ;
        RECT 321.200 281.600 322.000 290.200 ;
        RECT 325.000 281.600 325.800 290.200 ;
        RECT 330.800 281.600 331.600 290.200 ;
        RECT 336.400 281.600 337.200 286.200 ;
        RECT 339.600 281.600 340.400 286.200 ;
        RECT 345.200 281.600 346.000 290.000 ;
        RECT 350.000 281.600 350.800 290.200 ;
        RECT 355.600 281.600 356.400 286.200 ;
        RECT 358.800 281.600 359.600 286.200 ;
        RECT 364.400 281.600 365.200 290.000 ;
        RECT 369.200 281.600 370.000 290.200 ;
        RECT 374.800 281.600 375.600 286.200 ;
        RECT 378.000 281.600 378.800 286.200 ;
        RECT 383.600 281.600 384.400 290.000 ;
        RECT 388.400 281.600 389.400 288.800 ;
        RECT 394.600 282.200 395.600 288.800 ;
        RECT 394.600 281.600 395.400 282.200 ;
        RECT 398.600 281.600 399.400 286.200 ;
        RECT 402.800 281.600 403.600 290.200 ;
        RECT 404.400 281.600 405.200 286.200 ;
        RECT 408.200 281.600 409.000 286.200 ;
        RECT 412.400 281.600 413.200 290.200 ;
        RECT 415.600 281.600 416.400 290.200 ;
        RECT 421.200 281.600 422.000 286.200 ;
        RECT 424.400 281.600 425.200 286.200 ;
        RECT 430.000 281.600 430.800 290.000 ;
        RECT 434.800 281.600 435.800 288.800 ;
        RECT 441.000 282.200 442.000 288.800 ;
        RECT 441.000 281.600 441.800 282.200 ;
        RECT 449.200 281.600 450.000 286.200 ;
        RECT 452.400 281.600 453.200 290.200 ;
        RECT 456.600 281.600 457.400 286.200 ;
        RECT 458.800 281.600 459.600 290.200 ;
        RECT 463.000 281.600 463.800 286.200 ;
        RECT 466.800 281.600 467.600 290.000 ;
        RECT 472.400 281.600 473.200 286.200 ;
        RECT 475.600 281.600 476.400 286.200 ;
        RECT 481.200 281.600 482.000 290.200 ;
        RECT 486.000 281.600 487.000 288.800 ;
        RECT 492.200 282.200 493.200 288.800 ;
        RECT 492.200 281.600 493.000 282.200 ;
        RECT 495.600 281.600 496.400 290.200 ;
        RECT 498.800 281.600 499.600 290.200 ;
        RECT 502.000 281.600 502.800 290.200 ;
        RECT 505.200 281.600 506.000 290.200 ;
        RECT 508.400 281.600 509.200 290.200 ;
        RECT 511.600 281.600 512.400 290.000 ;
        RECT 517.200 281.600 518.000 286.200 ;
        RECT 520.400 281.600 521.200 286.200 ;
        RECT 526.000 281.600 526.800 290.200 ;
        RECT 530.800 281.600 531.600 289.000 ;
        RECT 534.000 281.600 534.800 286.200 ;
        RECT 537.200 281.600 538.000 286.200 ;
        RECT 540.400 281.600 541.200 286.200 ;
        RECT 543.600 281.600 544.400 286.200 ;
        RECT 551.600 281.600 552.400 286.200 ;
        RECT 554.800 281.600 555.600 286.200 ;
        RECT 561.200 281.600 562.000 286.200 ;
        RECT 564.400 281.600 565.200 286.200 ;
        RECT 567.600 281.600 568.400 286.200 ;
        RECT 569.200 281.600 570.000 286.200 ;
        RECT 572.400 281.600 573.200 286.200 ;
        RECT 576.200 281.600 577.000 290.200 ;
        RECT 582.000 281.600 582.800 289.000 ;
        RECT 0.400 280.400 586.800 281.600 ;
        RECT 4.400 273.000 5.200 280.400 ;
        RECT 9.200 273.200 10.200 280.400 ;
        RECT 15.400 279.800 16.200 280.400 ;
        RECT 15.400 273.200 16.400 279.800 ;
        RECT 18.800 275.800 19.600 280.400 ;
        RECT 22.600 275.800 23.400 280.400 ;
        RECT 26.800 271.800 27.600 280.400 ;
        RECT 28.400 275.800 29.200 280.400 ;
        RECT 32.200 275.800 33.000 280.400 ;
        RECT 36.400 271.800 37.200 280.400 ;
        RECT 41.200 273.000 42.000 280.400 ;
        RECT 46.000 275.800 46.800 280.400 ;
        RECT 49.200 273.000 50.000 280.400 ;
        RECT 55.600 275.800 56.400 280.400 ;
        RECT 60.400 273.200 61.400 280.400 ;
        RECT 66.600 279.800 67.400 280.400 ;
        RECT 66.600 273.200 67.600 279.800 ;
        RECT 71.600 272.200 72.400 280.400 ;
        RECT 76.800 271.800 77.600 280.400 ;
        RECT 80.200 275.800 81.000 280.400 ;
        RECT 84.400 271.800 85.200 280.400 ;
        RECT 87.800 279.800 88.600 280.400 ;
        RECT 87.600 273.200 88.600 279.800 ;
        RECT 93.800 273.200 94.800 280.400 ;
        RECT 98.800 273.000 99.600 280.400 ;
        RECT 105.200 275.800 106.000 280.400 ;
        RECT 106.800 271.800 107.600 280.400 ;
        RECT 113.200 273.000 114.000 280.400 ;
        RECT 116.400 271.800 117.200 280.400 ;
        RECT 118.600 275.800 119.400 280.400 ;
        RECT 122.800 271.800 123.600 280.400 ;
        RECT 124.400 271.800 125.200 280.400 ;
        RECT 128.200 275.800 129.000 280.400 ;
        RECT 132.400 271.800 133.200 280.400 ;
        RECT 134.000 275.800 134.800 280.400 ;
        RECT 137.200 275.800 138.000 280.400 ;
        RECT 143.600 271.800 144.400 280.400 ;
        RECT 147.800 275.800 148.600 280.400 ;
        RECT 150.600 275.800 151.400 280.400 ;
        RECT 154.800 271.800 155.600 280.400 ;
        RECT 158.000 275.800 158.800 280.400 ;
        RECT 159.600 271.800 160.400 280.400 ;
        RECT 166.000 271.800 166.800 280.400 ;
        RECT 167.600 271.800 168.400 280.400 ;
        RECT 171.800 275.800 172.600 280.400 ;
        RECT 174.000 275.800 174.800 280.400 ;
        RECT 177.200 275.800 178.000 280.400 ;
        RECT 180.400 271.800 181.200 280.400 ;
        RECT 186.000 275.800 186.800 280.400 ;
        RECT 189.200 275.800 190.000 280.400 ;
        RECT 194.800 272.000 195.600 280.400 ;
        RECT 199.600 271.800 200.400 280.400 ;
        RECT 205.200 275.800 206.000 280.400 ;
        RECT 208.400 275.800 209.200 280.400 ;
        RECT 214.000 272.000 214.800 280.400 ;
        RECT 219.000 279.800 219.800 280.400 ;
        RECT 218.800 273.200 219.800 279.800 ;
        RECT 225.000 273.200 226.000 280.400 ;
        RECT 230.000 273.000 230.800 280.400 ;
        RECT 234.800 271.800 235.600 280.400 ;
        RECT 240.200 275.800 241.000 280.400 ;
        RECT 244.400 271.800 245.200 280.400 ;
        RECT 246.600 275.800 247.400 280.400 ;
        RECT 250.800 271.800 251.600 280.400 ;
        RECT 254.000 272.200 254.800 280.400 ;
        RECT 257.200 275.800 258.000 280.400 ;
        RECT 258.800 275.800 259.600 280.400 ;
        RECT 262.000 275.800 262.800 280.400 ;
        RECT 263.600 271.800 264.400 280.400 ;
        RECT 267.800 275.800 268.600 280.400 ;
        RECT 271.800 279.800 272.600 280.400 ;
        RECT 271.600 273.200 272.600 279.800 ;
        RECT 277.800 273.200 278.800 280.400 ;
        RECT 282.800 275.800 283.600 280.400 ;
        RECT 286.200 279.800 287.000 280.400 ;
        RECT 286.000 273.200 287.000 279.800 ;
        RECT 292.200 273.200 293.200 280.400 ;
        RECT 303.600 271.800 304.400 280.400 ;
        RECT 305.200 271.800 306.000 280.400 ;
        RECT 311.600 275.800 312.400 280.400 ;
        RECT 313.800 275.800 314.600 280.400 ;
        RECT 318.000 271.800 318.800 280.400 ;
        RECT 319.600 271.800 320.400 280.400 ;
        RECT 326.000 271.800 326.800 280.400 ;
        RECT 329.200 275.800 330.000 280.400 ;
        RECT 330.800 275.800 331.600 280.400 ;
        RECT 334.000 275.800 334.800 280.400 ;
        RECT 337.800 271.800 338.600 280.400 ;
        RECT 343.600 271.800 344.400 280.400 ;
        RECT 349.200 275.800 350.000 280.400 ;
        RECT 352.400 275.800 353.200 280.400 ;
        RECT 358.000 272.000 358.800 280.400 ;
        RECT 363.000 279.800 363.800 280.400 ;
        RECT 362.800 273.200 363.800 279.800 ;
        RECT 369.000 273.200 370.000 280.400 ;
        RECT 373.000 275.800 373.800 280.400 ;
        RECT 377.200 271.800 378.000 280.400 ;
        RECT 380.400 275.800 381.200 280.400 ;
        RECT 382.000 275.800 382.800 280.400 ;
        RECT 385.200 276.200 386.000 280.400 ;
        RECT 390.000 273.000 390.800 280.400 ;
        RECT 396.400 275.800 397.200 280.400 ;
        RECT 398.000 275.800 398.800 280.400 ;
        RECT 401.200 275.800 402.000 280.400 ;
        RECT 402.800 271.800 403.600 280.400 ;
        RECT 407.600 275.800 408.400 280.400 ;
        RECT 412.400 275.800 413.200 280.400 ;
        RECT 415.600 271.800 416.400 280.400 ;
        RECT 421.200 275.800 422.000 280.400 ;
        RECT 424.400 275.800 425.200 280.400 ;
        RECT 430.000 272.000 430.800 280.400 ;
        RECT 436.400 271.800 437.200 280.400 ;
        RECT 438.600 275.800 439.400 280.400 ;
        RECT 442.800 271.800 443.600 280.400 ;
        RECT 451.000 279.800 451.800 280.400 ;
        RECT 450.800 273.200 451.800 279.800 ;
        RECT 457.000 273.200 458.000 280.400 ;
        RECT 460.400 275.800 461.200 280.400 ;
        RECT 463.600 275.800 464.400 280.400 ;
        RECT 466.800 272.000 467.600 280.400 ;
        RECT 472.400 275.800 473.200 280.400 ;
        RECT 475.600 275.800 476.400 280.400 ;
        RECT 481.200 271.800 482.000 280.400 ;
        RECT 486.000 272.000 486.800 280.400 ;
        RECT 491.600 275.800 492.400 280.400 ;
        RECT 494.800 275.800 495.600 280.400 ;
        RECT 500.400 271.800 501.200 280.400 ;
        RECT 505.200 272.000 506.000 280.400 ;
        RECT 510.800 275.800 511.600 280.400 ;
        RECT 514.000 275.800 514.800 280.400 ;
        RECT 519.600 271.800 520.400 280.400 ;
        RECT 524.400 272.000 525.200 280.400 ;
        RECT 530.000 275.800 530.800 280.400 ;
        RECT 533.200 275.800 534.000 280.400 ;
        RECT 538.800 271.800 539.600 280.400 ;
        RECT 543.600 272.000 544.400 280.400 ;
        RECT 549.200 275.800 550.000 280.400 ;
        RECT 552.400 275.800 553.200 280.400 ;
        RECT 558.000 271.800 558.800 280.400 ;
        RECT 562.800 272.000 563.600 280.400 ;
        RECT 568.400 275.800 569.200 280.400 ;
        RECT 571.600 275.800 572.400 280.400 ;
        RECT 577.200 271.800 578.000 280.400 ;
        RECT 582.000 273.000 582.800 280.400 ;
        RECT 1.200 241.600 2.000 250.200 ;
        RECT 5.400 241.600 6.200 246.200 ;
        RECT 7.600 241.600 8.400 246.200 ;
        RECT 10.800 241.600 11.600 246.200 ;
        RECT 12.400 241.600 13.200 250.200 ;
        RECT 15.600 241.600 16.400 246.200 ;
        RECT 20.400 241.600 21.200 249.000 ;
        RECT 26.800 241.600 27.600 249.800 ;
        RECT 32.000 241.600 32.800 250.200 ;
        RECT 35.400 241.600 36.200 246.200 ;
        RECT 39.600 241.600 40.400 250.200 ;
        RECT 41.200 241.600 42.000 246.200 ;
        RECT 44.400 241.600 45.200 246.200 ;
        RECT 49.200 241.600 50.000 250.200 ;
        RECT 52.400 241.600 53.400 248.800 ;
        RECT 58.600 242.200 59.600 248.800 ;
        RECT 63.600 242.200 64.600 248.800 ;
        RECT 58.600 241.600 59.400 242.200 ;
        RECT 63.800 241.600 64.600 242.200 ;
        RECT 69.800 241.600 70.800 248.800 ;
        RECT 74.800 241.600 75.600 249.000 ;
        RECT 81.200 241.600 82.000 246.200 ;
        RECT 82.800 241.600 83.600 250.200 ;
        RECT 87.000 241.600 87.800 246.200 ;
        RECT 90.800 241.600 91.600 246.200 ;
        RECT 94.000 241.600 94.800 246.200 ;
        RECT 95.600 241.600 96.400 246.200 ;
        RECT 98.800 241.600 99.600 245.800 ;
        RECT 102.000 241.600 102.800 250.200 ;
        RECT 106.200 241.600 107.000 246.200 ;
        RECT 110.000 241.600 110.800 246.200 ;
        RECT 114.800 241.600 115.600 250.200 ;
        RECT 117.000 241.600 117.800 246.200 ;
        RECT 121.200 241.600 122.000 250.200 ;
        RECT 126.000 241.600 126.800 250.200 ;
        RECT 129.200 242.200 130.200 248.800 ;
        RECT 129.400 241.600 130.200 242.200 ;
        RECT 135.400 241.600 136.400 248.800 ;
        RECT 145.200 242.200 146.200 248.800 ;
        RECT 145.400 241.600 146.200 242.200 ;
        RECT 151.400 241.600 152.400 248.800 ;
        RECT 154.800 241.600 155.600 246.200 ;
        RECT 158.000 241.600 158.800 246.200 ;
        RECT 159.600 241.600 160.400 250.200 ;
        RECT 163.800 241.600 164.600 246.200 ;
        RECT 166.000 241.600 166.800 246.200 ;
        RECT 169.200 241.600 170.000 246.200 ;
        RECT 171.400 241.600 172.200 246.200 ;
        RECT 175.600 241.600 176.400 250.200 ;
        RECT 180.400 241.600 181.200 250.200 ;
        RECT 182.600 241.600 183.400 246.200 ;
        RECT 186.800 241.600 187.600 250.200 ;
        RECT 190.000 241.600 190.800 246.200 ;
        RECT 193.200 241.600 194.000 246.200 ;
        RECT 198.000 241.600 198.800 250.200 ;
        RECT 201.200 241.600 202.000 250.200 ;
        RECT 206.800 241.600 207.600 246.200 ;
        RECT 210.000 241.600 210.800 246.200 ;
        RECT 215.600 241.600 216.400 250.000 ;
        RECT 220.400 241.600 221.200 250.200 ;
        RECT 226.000 241.600 226.800 246.200 ;
        RECT 229.200 241.600 230.000 246.200 ;
        RECT 234.800 241.600 235.600 250.000 ;
        RECT 239.600 241.600 240.400 249.000 ;
        RECT 244.400 241.600 245.200 250.200 ;
        RECT 250.000 241.600 250.800 246.200 ;
        RECT 253.200 241.600 254.000 246.200 ;
        RECT 258.800 241.600 259.600 250.000 ;
        RECT 263.600 241.600 264.400 250.200 ;
        RECT 269.200 241.600 270.000 246.200 ;
        RECT 272.400 241.600 273.200 246.200 ;
        RECT 278.000 241.600 278.800 250.000 ;
        RECT 282.800 241.600 283.600 249.000 ;
        RECT 292.400 241.600 293.200 250.200 ;
        RECT 298.000 241.600 298.800 246.200 ;
        RECT 301.200 241.600 302.000 246.200 ;
        RECT 306.800 241.600 307.600 250.000 ;
        RECT 311.600 242.200 312.600 248.800 ;
        RECT 311.800 241.600 312.600 242.200 ;
        RECT 317.800 241.600 318.800 248.800 ;
        RECT 321.800 241.600 322.600 246.200 ;
        RECT 326.000 241.600 326.800 250.200 ;
        RECT 327.600 241.600 328.400 246.200 ;
        RECT 330.800 241.600 331.600 246.200 ;
        RECT 332.400 241.600 333.200 250.200 ;
        RECT 338.800 241.600 339.600 250.200 ;
        RECT 340.400 241.600 341.200 250.200 ;
        RECT 345.200 241.600 346.000 246.200 ;
        RECT 348.400 241.600 349.200 246.200 ;
        RECT 350.000 241.600 350.800 250.200 ;
        RECT 356.400 241.600 357.200 246.200 ;
        RECT 358.600 241.600 359.400 246.200 ;
        RECT 362.800 241.600 363.600 250.200 ;
        RECT 366.000 241.600 366.800 246.200 ;
        RECT 369.200 241.600 370.000 250.200 ;
        RECT 374.800 241.600 375.600 246.200 ;
        RECT 378.000 241.600 378.800 246.200 ;
        RECT 383.600 241.600 384.400 250.000 ;
        RECT 388.400 241.600 389.200 249.000 ;
        RECT 394.800 241.600 395.600 250.200 ;
        RECT 401.200 241.600 402.000 250.200 ;
        RECT 406.800 241.600 407.600 246.200 ;
        RECT 410.000 241.600 410.800 246.200 ;
        RECT 415.600 241.600 416.400 250.000 ;
        RECT 420.400 241.600 421.200 250.200 ;
        RECT 426.000 241.600 426.800 246.200 ;
        RECT 429.200 241.600 430.000 246.200 ;
        RECT 434.800 241.600 435.600 250.000 ;
        RECT 439.600 241.600 440.400 249.000 ;
        RECT 450.800 241.600 451.600 245.800 ;
        RECT 454.000 241.600 454.800 246.200 ;
        RECT 458.800 241.600 459.600 250.200 ;
        RECT 462.000 241.600 462.800 249.000 ;
        RECT 468.400 241.600 469.200 246.200 ;
        RECT 472.200 241.600 473.000 246.200 ;
        RECT 476.400 241.600 477.200 250.200 ;
        RECT 478.000 241.600 478.800 246.200 ;
        RECT 481.200 241.600 482.000 246.200 ;
        RECT 483.400 241.600 484.200 246.200 ;
        RECT 487.600 241.600 488.400 250.200 ;
        RECT 489.200 241.600 490.000 246.200 ;
        RECT 492.400 241.600 493.200 246.200 ;
        RECT 494.000 241.600 494.800 250.200 ;
        RECT 502.000 241.600 502.800 250.200 ;
        RECT 505.200 241.600 506.200 248.800 ;
        RECT 511.400 242.200 512.400 248.800 ;
        RECT 516.400 242.200 517.400 248.800 ;
        RECT 511.400 241.600 512.200 242.200 ;
        RECT 516.600 241.600 517.400 242.200 ;
        RECT 522.600 241.600 523.600 248.800 ;
        RECT 527.600 241.600 528.600 248.800 ;
        RECT 533.800 242.200 534.800 248.800 ;
        RECT 533.800 241.600 534.600 242.200 ;
        RECT 538.800 241.600 539.600 250.000 ;
        RECT 544.400 241.600 545.200 246.200 ;
        RECT 547.600 241.600 548.400 246.200 ;
        RECT 553.200 241.600 554.000 250.200 ;
        RECT 558.000 241.600 558.800 249.000 ;
        RECT 562.800 241.600 563.600 250.000 ;
        RECT 568.400 241.600 569.200 246.200 ;
        RECT 571.600 241.600 572.400 246.200 ;
        RECT 577.200 241.600 578.000 250.200 ;
        RECT 582.000 241.600 582.800 249.000 ;
        RECT 0.400 240.400 586.800 241.600 ;
        RECT 2.800 231.800 3.600 240.400 ;
        RECT 8.400 235.800 9.200 240.400 ;
        RECT 11.600 235.800 12.400 240.400 ;
        RECT 17.200 232.000 18.000 240.400 ;
        RECT 22.000 233.200 23.000 240.400 ;
        RECT 28.200 239.800 29.000 240.400 ;
        RECT 28.200 233.200 29.200 239.800 ;
        RECT 33.200 233.200 34.200 240.400 ;
        RECT 39.400 239.800 40.200 240.400 ;
        RECT 39.400 233.200 40.400 239.800 ;
        RECT 44.400 231.800 45.200 240.400 ;
        RECT 50.000 235.800 50.800 240.400 ;
        RECT 53.200 235.800 54.000 240.400 ;
        RECT 58.800 232.000 59.600 240.400 ;
        RECT 63.600 232.000 64.400 240.400 ;
        RECT 69.200 235.800 70.000 240.400 ;
        RECT 72.400 235.800 73.200 240.400 ;
        RECT 78.000 231.800 78.800 240.400 ;
        RECT 83.000 239.800 83.800 240.400 ;
        RECT 82.800 233.200 83.800 239.800 ;
        RECT 89.000 233.200 90.000 240.400 ;
        RECT 92.400 235.800 93.200 240.400 ;
        RECT 95.600 235.800 96.400 240.400 ;
        RECT 98.800 231.800 99.600 240.400 ;
        RECT 104.400 235.800 105.200 240.400 ;
        RECT 107.600 235.800 108.400 240.400 ;
        RECT 113.200 232.000 114.000 240.400 ;
        RECT 118.000 231.800 118.800 240.400 ;
        RECT 123.600 235.800 124.400 240.400 ;
        RECT 126.800 235.800 127.600 240.400 ;
        RECT 132.400 232.000 133.200 240.400 ;
        RECT 142.200 239.800 143.000 240.400 ;
        RECT 142.000 233.200 143.000 239.800 ;
        RECT 148.200 233.200 149.200 240.400 ;
        RECT 151.600 231.800 152.400 240.400 ;
        RECT 155.800 235.800 156.600 240.400 ;
        RECT 158.000 231.800 158.800 240.400 ;
        RECT 162.200 235.800 163.000 240.400 ;
        RECT 166.000 231.800 166.800 240.400 ;
        RECT 171.600 235.800 172.400 240.400 ;
        RECT 174.800 235.800 175.600 240.400 ;
        RECT 180.400 232.000 181.200 240.400 ;
        RECT 183.600 231.800 184.400 240.400 ;
        RECT 186.800 231.800 187.600 240.400 ;
        RECT 190.000 231.800 190.800 240.400 ;
        RECT 193.200 231.800 194.000 240.400 ;
        RECT 196.400 231.800 197.200 240.400 ;
        RECT 199.600 231.800 200.400 240.400 ;
        RECT 205.200 235.800 206.000 240.400 ;
        RECT 208.400 235.800 209.200 240.400 ;
        RECT 214.000 232.000 214.800 240.400 ;
        RECT 218.800 231.800 219.600 240.400 ;
        RECT 224.400 235.800 225.200 240.400 ;
        RECT 227.600 235.800 228.400 240.400 ;
        RECT 233.200 232.000 234.000 240.400 ;
        RECT 236.400 235.800 237.200 240.400 ;
        RECT 241.200 233.000 242.000 240.400 ;
        RECT 246.000 232.000 246.800 240.400 ;
        RECT 251.600 235.800 252.400 240.400 ;
        RECT 254.800 235.800 255.600 240.400 ;
        RECT 260.400 231.800 261.200 240.400 ;
        RECT 265.200 232.000 266.000 240.400 ;
        RECT 270.800 235.800 271.600 240.400 ;
        RECT 274.000 235.800 274.800 240.400 ;
        RECT 279.600 231.800 280.400 240.400 ;
        RECT 282.800 235.800 283.600 240.400 ;
        RECT 286.000 235.800 286.800 240.400 ;
        RECT 289.200 235.800 290.000 240.400 ;
        RECT 298.800 231.800 299.600 240.400 ;
        RECT 302.000 235.800 302.800 240.400 ;
        RECT 303.600 231.800 304.400 240.400 ;
        RECT 310.000 232.000 310.800 240.400 ;
        RECT 315.600 235.800 316.400 240.400 ;
        RECT 318.800 235.800 319.600 240.400 ;
        RECT 324.400 231.800 325.200 240.400 ;
        RECT 327.600 235.800 328.400 240.400 ;
        RECT 330.800 235.800 331.600 240.400 ;
        RECT 332.400 235.800 333.200 240.400 ;
        RECT 335.600 235.800 336.400 240.400 ;
        RECT 338.800 235.800 339.600 240.400 ;
        RECT 342.000 232.000 342.800 240.400 ;
        RECT 347.600 235.800 348.400 240.400 ;
        RECT 350.800 235.800 351.600 240.400 ;
        RECT 356.400 231.800 357.200 240.400 ;
        RECT 361.200 233.000 362.000 240.400 ;
        RECT 366.000 231.800 366.800 240.400 ;
        RECT 371.600 235.800 372.400 240.400 ;
        RECT 374.800 235.800 375.600 240.400 ;
        RECT 380.400 232.000 381.200 240.400 ;
        RECT 385.200 232.000 386.000 240.400 ;
        RECT 390.800 235.800 391.600 240.400 ;
        RECT 394.000 235.800 394.800 240.400 ;
        RECT 399.600 231.800 400.400 240.400 ;
        RECT 404.400 232.000 405.200 240.400 ;
        RECT 410.000 235.800 410.800 240.400 ;
        RECT 413.200 235.800 414.000 240.400 ;
        RECT 418.800 231.800 419.600 240.400 ;
        RECT 422.000 235.800 422.800 240.400 ;
        RECT 425.200 235.800 426.000 240.400 ;
        RECT 426.800 231.800 427.600 240.400 ;
        RECT 434.800 231.800 435.600 240.400 ;
        RECT 436.400 235.800 437.200 240.400 ;
        RECT 441.200 236.200 442.000 240.400 ;
        RECT 444.400 235.800 445.200 240.400 ;
        RECT 452.400 235.800 453.200 240.400 ;
        RECT 457.200 231.800 458.000 240.400 ;
        RECT 458.800 235.800 459.600 240.400 ;
        RECT 462.000 235.800 462.800 240.400 ;
        RECT 463.600 235.800 464.400 240.400 ;
        RECT 466.800 235.800 467.600 240.400 ;
        RECT 468.400 231.800 469.200 240.400 ;
        RECT 474.800 231.800 475.600 240.400 ;
        RECT 476.400 235.800 477.200 240.400 ;
        RECT 481.200 233.200 482.200 240.400 ;
        RECT 487.400 239.800 488.200 240.400 ;
        RECT 487.400 233.200 488.400 239.800 ;
        RECT 492.400 232.000 493.200 240.400 ;
        RECT 498.000 235.800 498.800 240.400 ;
        RECT 501.200 235.800 502.000 240.400 ;
        RECT 506.800 231.800 507.600 240.400 ;
        RECT 511.600 232.000 512.400 240.400 ;
        RECT 517.200 235.800 518.000 240.400 ;
        RECT 520.400 235.800 521.200 240.400 ;
        RECT 526.000 231.800 526.800 240.400 ;
        RECT 530.800 233.000 531.600 240.400 ;
        RECT 535.600 232.000 536.400 240.400 ;
        RECT 541.200 235.800 542.000 240.400 ;
        RECT 544.400 235.800 545.200 240.400 ;
        RECT 550.000 231.800 550.800 240.400 ;
        RECT 554.800 232.000 555.600 240.400 ;
        RECT 560.400 235.800 561.200 240.400 ;
        RECT 563.600 235.800 564.400 240.400 ;
        RECT 569.200 231.800 570.000 240.400 ;
        RECT 574.000 233.000 574.800 240.400 ;
        RECT 578.800 233.000 579.600 240.400 ;
        RECT 2.800 201.600 3.600 210.000 ;
        RECT 8.400 201.600 9.200 206.200 ;
        RECT 11.600 201.600 12.400 206.200 ;
        RECT 17.200 201.600 18.000 210.200 ;
        RECT 22.000 201.600 22.800 210.000 ;
        RECT 27.600 201.600 28.400 206.200 ;
        RECT 30.800 201.600 31.600 206.200 ;
        RECT 36.400 201.600 37.200 210.200 ;
        RECT 41.200 201.600 42.000 210.200 ;
        RECT 46.800 201.600 47.600 206.200 ;
        RECT 50.000 201.600 50.800 206.200 ;
        RECT 55.600 201.600 56.400 210.000 ;
        RECT 60.400 201.600 61.200 210.000 ;
        RECT 66.000 201.600 66.800 206.200 ;
        RECT 69.200 201.600 70.000 206.200 ;
        RECT 74.800 201.600 75.600 210.200 ;
        RECT 79.600 201.600 80.400 210.200 ;
        RECT 85.200 201.600 86.000 206.200 ;
        RECT 88.400 201.600 89.200 206.200 ;
        RECT 94.000 201.600 94.800 210.000 ;
        RECT 97.200 201.600 98.000 210.200 ;
        RECT 100.400 201.600 101.200 210.200 ;
        RECT 103.600 201.600 104.400 210.200 ;
        RECT 106.800 201.600 107.600 210.200 ;
        RECT 110.000 201.600 110.800 210.200 ;
        RECT 113.200 201.600 114.000 210.200 ;
        RECT 118.800 201.600 119.600 206.200 ;
        RECT 122.000 201.600 122.800 206.200 ;
        RECT 127.600 201.600 128.400 210.000 ;
        RECT 137.200 201.600 138.000 210.000 ;
        RECT 142.800 201.600 143.600 206.200 ;
        RECT 146.000 201.600 146.800 206.200 ;
        RECT 151.600 201.600 152.400 210.200 ;
        RECT 156.400 201.600 157.200 210.000 ;
        RECT 162.000 201.600 162.800 206.200 ;
        RECT 165.200 201.600 166.000 206.200 ;
        RECT 170.800 201.600 171.600 210.200 ;
        RECT 174.000 201.600 174.800 206.200 ;
        RECT 177.200 201.600 178.000 210.200 ;
        RECT 182.000 201.600 182.800 210.200 ;
        RECT 186.200 201.600 187.000 206.200 ;
        RECT 188.400 201.600 189.200 210.200 ;
        RECT 193.200 201.600 194.000 206.200 ;
        RECT 196.400 201.600 197.200 210.200 ;
        RECT 200.600 201.600 201.400 206.200 ;
        RECT 204.400 201.600 205.200 210.000 ;
        RECT 210.000 201.600 210.800 206.200 ;
        RECT 213.200 201.600 214.000 206.200 ;
        RECT 218.800 201.600 219.600 210.200 ;
        RECT 225.200 201.600 226.000 210.200 ;
        RECT 226.800 201.600 227.600 206.200 ;
        RECT 230.000 201.600 230.800 210.200 ;
        RECT 234.800 201.600 235.600 210.200 ;
        RECT 239.000 201.600 239.800 206.200 ;
        RECT 241.200 201.600 242.000 210.200 ;
        RECT 245.400 201.600 246.200 206.200 ;
        RECT 247.600 201.600 248.400 210.200 ;
        RECT 251.800 201.600 252.600 206.200 ;
        RECT 255.600 201.600 256.400 210.000 ;
        RECT 261.200 201.600 262.000 206.200 ;
        RECT 264.400 201.600 265.200 206.200 ;
        RECT 270.000 201.600 270.800 210.200 ;
        RECT 273.200 201.600 274.000 206.200 ;
        RECT 276.400 201.600 277.200 210.200 ;
        RECT 281.200 201.600 282.000 206.200 ;
        RECT 284.400 201.600 285.200 206.200 ;
        RECT 287.600 201.600 288.400 206.200 ;
        RECT 294.000 201.600 294.800 210.200 ;
        RECT 300.400 201.600 301.200 210.200 ;
        RECT 306.000 201.600 306.800 206.200 ;
        RECT 309.200 201.600 310.000 206.200 ;
        RECT 314.800 201.600 315.600 210.000 ;
        RECT 319.600 201.600 320.400 209.000 ;
        RECT 324.400 201.600 325.200 210.200 ;
        RECT 330.000 201.600 330.800 206.200 ;
        RECT 333.200 201.600 334.000 206.200 ;
        RECT 338.800 201.600 339.600 210.000 ;
        RECT 343.600 201.600 344.400 209.000 ;
        RECT 348.400 201.600 349.200 210.000 ;
        RECT 354.000 201.600 354.800 206.200 ;
        RECT 357.200 201.600 358.000 206.200 ;
        RECT 362.800 201.600 363.600 210.200 ;
        RECT 366.000 201.600 366.800 206.200 ;
        RECT 369.200 201.600 370.000 210.200 ;
        RECT 373.400 201.600 374.200 206.200 ;
        RECT 375.600 201.600 376.400 210.200 ;
        RECT 379.800 201.600 380.600 206.200 ;
        RECT 383.600 202.200 384.600 208.800 ;
        RECT 383.800 201.600 384.600 202.200 ;
        RECT 389.800 201.600 390.800 208.800 ;
        RECT 393.200 201.600 394.000 206.200 ;
        RECT 397.000 201.600 397.800 206.200 ;
        RECT 401.200 201.600 402.000 210.200 ;
        RECT 404.400 201.600 405.400 208.800 ;
        RECT 410.600 202.200 411.600 208.800 ;
        RECT 410.600 201.600 411.400 202.200 ;
        RECT 415.600 201.600 416.400 210.000 ;
        RECT 421.200 201.600 422.000 206.200 ;
        RECT 424.400 201.600 425.200 206.200 ;
        RECT 430.000 201.600 430.800 210.200 ;
        RECT 435.400 201.600 436.200 210.200 ;
        RECT 442.800 201.600 443.600 210.200 ;
        RECT 449.200 201.600 450.000 206.200 ;
        RECT 452.400 201.600 453.200 206.200 ;
        RECT 457.200 201.600 458.000 210.200 ;
        RECT 458.800 201.600 459.600 210.200 ;
        RECT 463.000 201.600 463.800 206.200 ;
        RECT 465.200 201.600 466.000 206.200 ;
        RECT 468.400 201.600 469.200 206.200 ;
        RECT 470.000 201.600 470.800 210.200 ;
        RECT 474.200 201.600 475.000 206.200 ;
        RECT 476.400 201.600 477.200 210.200 ;
        RECT 480.600 201.600 481.400 206.200 ;
        RECT 482.800 201.600 483.600 206.200 ;
        RECT 486.000 201.600 486.800 206.200 ;
        RECT 487.600 201.600 488.400 206.200 ;
        RECT 490.800 201.600 491.600 210.200 ;
        RECT 497.200 201.600 498.000 210.200 ;
        RECT 498.800 201.600 499.600 206.200 ;
        RECT 502.000 201.600 502.800 206.200 ;
        RECT 505.200 202.200 506.200 208.800 ;
        RECT 505.400 201.600 506.200 202.200 ;
        RECT 511.400 201.600 512.400 208.800 ;
        RECT 516.400 201.600 517.400 208.800 ;
        RECT 522.600 202.200 523.600 208.800 ;
        RECT 522.600 201.600 523.400 202.200 ;
        RECT 527.600 201.600 528.400 209.000 ;
        RECT 534.000 201.600 534.800 206.200 ;
        RECT 537.200 201.600 538.000 206.200 ;
        RECT 538.800 201.600 539.600 206.200 ;
        RECT 542.000 201.600 542.800 206.200 ;
        RECT 545.200 201.600 546.000 210.000 ;
        RECT 550.800 201.600 551.600 206.200 ;
        RECT 554.000 201.600 554.800 206.200 ;
        RECT 559.600 201.600 560.400 210.200 ;
        RECT 564.400 201.600 565.200 210.000 ;
        RECT 570.000 201.600 570.800 206.200 ;
        RECT 573.200 201.600 574.000 206.200 ;
        RECT 578.800 201.600 579.600 210.200 ;
        RECT 583.600 201.600 584.400 209.000 ;
        RECT 0.400 200.400 586.800 201.600 ;
        RECT 2.800 192.000 3.600 200.400 ;
        RECT 8.400 195.800 9.200 200.400 ;
        RECT 11.600 195.800 12.400 200.400 ;
        RECT 17.200 191.800 18.000 200.400 ;
        RECT 22.000 192.000 22.800 200.400 ;
        RECT 27.600 195.800 28.400 200.400 ;
        RECT 30.800 195.800 31.600 200.400 ;
        RECT 36.400 191.800 37.200 200.400 ;
        RECT 39.600 195.800 40.400 200.400 ;
        RECT 42.800 195.800 43.600 200.400 ;
        RECT 47.000 191.800 47.800 200.400 ;
        RECT 50.800 191.800 51.600 200.400 ;
        RECT 55.600 195.800 56.400 200.400 ;
        RECT 58.800 195.800 59.600 200.400 ;
        RECT 60.400 195.800 61.200 200.400 ;
        RECT 63.600 195.800 64.400 200.400 ;
        RECT 65.800 195.800 66.600 200.400 ;
        RECT 70.000 191.800 70.800 200.400 ;
        RECT 71.600 195.800 72.400 200.400 ;
        RECT 74.800 192.200 75.600 200.400 ;
        RECT 78.000 195.800 78.800 200.400 ;
        RECT 81.200 195.800 82.000 200.400 ;
        RECT 84.400 195.800 85.200 200.400 ;
        RECT 87.600 195.800 88.400 200.400 ;
        RECT 89.200 195.800 90.000 200.400 ;
        RECT 92.400 195.800 93.200 200.400 ;
        RECT 94.000 195.800 94.800 200.400 ;
        RECT 97.200 191.800 98.000 200.400 ;
        RECT 101.400 195.800 102.200 200.400 ;
        RECT 104.200 195.800 105.000 200.400 ;
        RECT 108.400 191.800 109.200 200.400 ;
        RECT 110.000 195.800 110.800 200.400 ;
        RECT 113.200 195.800 114.000 200.400 ;
        RECT 114.800 195.800 115.600 200.400 ;
        RECT 118.000 195.800 118.800 200.400 ;
        RECT 121.200 195.800 122.000 200.400 ;
        RECT 124.400 192.000 125.200 200.400 ;
        RECT 130.000 195.800 130.800 200.400 ;
        RECT 133.200 195.800 134.000 200.400 ;
        RECT 138.800 191.800 139.600 200.400 ;
        RECT 148.400 192.000 149.200 200.400 ;
        RECT 154.000 195.800 154.800 200.400 ;
        RECT 157.200 195.800 158.000 200.400 ;
        RECT 162.800 191.800 163.600 200.400 ;
        RECT 167.600 192.000 168.400 200.400 ;
        RECT 173.200 195.800 174.000 200.400 ;
        RECT 176.400 195.800 177.200 200.400 ;
        RECT 182.000 191.800 182.800 200.400 ;
        RECT 185.200 195.800 186.000 200.400 ;
        RECT 189.000 195.800 189.800 200.400 ;
        RECT 193.200 191.800 194.000 200.400 ;
        RECT 194.800 195.800 195.600 200.400 ;
        RECT 198.000 195.800 198.800 200.400 ;
        RECT 200.200 195.800 201.000 200.400 ;
        RECT 204.400 191.800 205.200 200.400 ;
        RECT 206.000 195.800 206.800 200.400 ;
        RECT 209.200 195.800 210.000 200.400 ;
        RECT 212.400 195.800 213.200 200.400 ;
        RECT 215.600 193.200 216.600 200.400 ;
        RECT 221.800 199.800 222.600 200.400 ;
        RECT 221.800 193.200 222.800 199.800 ;
        RECT 226.800 192.000 227.600 200.400 ;
        RECT 232.400 195.800 233.200 200.400 ;
        RECT 235.600 195.800 236.400 200.400 ;
        RECT 241.200 191.800 242.000 200.400 ;
        RECT 245.000 195.800 245.800 200.400 ;
        RECT 249.200 191.800 250.000 200.400 ;
        RECT 250.800 195.800 251.600 200.400 ;
        RECT 257.200 191.800 258.000 200.400 ;
        RECT 260.600 199.800 261.400 200.400 ;
        RECT 260.400 193.200 261.400 199.800 ;
        RECT 266.600 193.200 267.600 200.400 ;
        RECT 270.000 195.800 270.800 200.400 ;
        RECT 273.200 195.800 274.000 200.400 ;
        RECT 276.400 192.000 277.200 200.400 ;
        RECT 282.000 195.800 282.800 200.400 ;
        RECT 285.200 195.800 286.000 200.400 ;
        RECT 290.800 191.800 291.600 200.400 ;
        RECT 298.800 195.800 299.600 200.400 ;
        RECT 302.000 195.800 302.800 200.400 ;
        RECT 303.600 195.800 304.400 200.400 ;
        RECT 306.800 195.800 307.600 200.400 ;
        RECT 310.000 191.800 310.800 200.400 ;
        RECT 312.200 195.800 313.000 200.400 ;
        RECT 316.400 191.800 317.200 200.400 ;
        RECT 318.000 195.800 318.800 200.400 ;
        RECT 321.200 195.800 322.000 200.400 ;
        RECT 324.600 199.800 325.400 200.400 ;
        RECT 324.400 193.200 325.400 199.800 ;
        RECT 330.600 193.200 331.600 200.400 ;
        RECT 334.000 191.800 334.800 200.400 ;
        RECT 338.200 195.800 339.000 200.400 ;
        RECT 340.400 195.800 341.200 200.400 ;
        RECT 343.600 195.800 344.400 200.400 ;
        RECT 346.800 193.200 347.800 200.400 ;
        RECT 353.000 199.800 353.800 200.400 ;
        RECT 353.000 193.200 354.000 199.800 ;
        RECT 358.000 192.000 358.800 200.400 ;
        RECT 363.600 195.800 364.400 200.400 ;
        RECT 366.800 195.800 367.600 200.400 ;
        RECT 372.400 191.800 373.200 200.400 ;
        RECT 377.200 192.200 378.000 200.400 ;
        RECT 382.400 191.800 383.200 200.400 ;
        RECT 385.800 195.800 386.600 200.400 ;
        RECT 390.000 191.800 390.800 200.400 ;
        RECT 391.600 191.800 392.400 200.400 ;
        RECT 399.600 191.800 400.400 200.400 ;
        RECT 401.200 195.800 402.000 200.400 ;
        RECT 404.400 191.800 405.200 200.400 ;
        RECT 410.800 191.800 411.600 200.400 ;
        RECT 416.400 195.800 417.200 200.400 ;
        RECT 419.600 195.800 420.400 200.400 ;
        RECT 425.200 192.000 426.000 200.400 ;
        RECT 430.000 192.000 430.800 200.400 ;
        RECT 435.600 195.800 436.400 200.400 ;
        RECT 438.800 195.800 439.600 200.400 ;
        RECT 444.400 191.800 445.200 200.400 ;
        RECT 454.000 193.000 454.800 200.400 ;
        RECT 459.400 195.800 460.200 200.400 ;
        RECT 463.600 191.800 464.400 200.400 ;
        RECT 467.000 199.800 467.800 200.400 ;
        RECT 466.800 193.200 467.800 199.800 ;
        RECT 473.000 193.200 474.000 200.400 ;
        RECT 476.400 191.800 477.200 200.400 ;
        RECT 480.600 195.800 481.400 200.400 ;
        RECT 484.400 195.800 485.200 200.400 ;
        RECT 486.000 191.800 486.800 200.400 ;
        RECT 490.200 195.800 491.000 200.400 ;
        RECT 494.000 193.000 494.800 200.400 ;
        RECT 500.400 193.200 501.400 200.400 ;
        RECT 506.600 199.800 507.400 200.400 ;
        RECT 506.600 193.200 507.600 199.800 ;
        RECT 510.000 195.800 510.800 200.400 ;
        RECT 513.200 191.800 514.000 200.400 ;
        RECT 518.000 195.800 518.800 200.400 ;
        RECT 521.200 195.800 522.000 200.400 ;
        RECT 522.800 191.800 523.600 200.400 ;
        RECT 526.000 191.800 526.800 200.400 ;
        RECT 527.600 195.800 528.400 200.400 ;
        RECT 530.800 195.800 531.600 200.400 ;
        RECT 532.400 195.800 533.200 200.400 ;
        RECT 535.600 195.800 536.400 200.400 ;
        RECT 538.800 195.800 539.600 200.400 ;
        RECT 542.000 191.800 542.800 200.400 ;
        RECT 543.600 191.800 544.400 200.400 ;
        RECT 547.800 195.800 548.600 200.400 ;
        RECT 553.200 191.800 554.000 200.400 ;
        RECT 556.400 193.200 557.400 200.400 ;
        RECT 562.600 199.800 563.400 200.400 ;
        RECT 562.600 193.200 563.600 199.800 ;
        RECT 567.600 192.000 568.400 200.400 ;
        RECT 573.200 195.800 574.000 200.400 ;
        RECT 576.400 195.800 577.200 200.400 ;
        RECT 582.000 191.800 582.800 200.400 ;
        RECT 2.800 161.600 3.600 170.200 ;
        RECT 8.400 161.600 9.200 166.200 ;
        RECT 11.600 161.600 12.400 166.200 ;
        RECT 17.200 161.600 18.000 170.000 ;
        RECT 21.000 161.600 21.800 166.200 ;
        RECT 25.200 161.600 26.000 170.200 ;
        RECT 28.400 161.600 29.400 168.800 ;
        RECT 34.600 162.200 35.600 168.800 ;
        RECT 34.600 161.600 35.400 162.200 ;
        RECT 39.600 161.600 40.600 168.800 ;
        RECT 45.800 162.200 46.800 168.800 ;
        RECT 45.800 161.600 46.600 162.200 ;
        RECT 49.800 161.600 50.600 166.200 ;
        RECT 54.000 161.600 54.800 170.200 ;
        RECT 58.800 161.600 59.600 169.000 ;
        RECT 62.600 161.600 63.400 166.200 ;
        RECT 66.800 161.600 67.600 170.200 ;
        RECT 70.000 161.600 70.800 166.200 ;
        RECT 71.600 161.600 72.400 170.200 ;
        RECT 76.400 161.600 77.200 170.200 ;
        RECT 80.600 161.600 81.400 166.200 ;
        RECT 84.400 161.600 85.400 168.800 ;
        RECT 90.600 162.200 91.600 168.800 ;
        RECT 95.600 162.200 96.600 168.800 ;
        RECT 90.600 161.600 91.400 162.200 ;
        RECT 95.800 161.600 96.600 162.200 ;
        RECT 101.800 161.600 102.800 168.800 ;
        RECT 106.800 161.600 107.600 170.000 ;
        RECT 112.400 161.600 113.200 166.200 ;
        RECT 115.600 161.600 116.400 166.200 ;
        RECT 121.200 161.600 122.000 170.200 ;
        RECT 124.400 161.600 125.200 166.200 ;
        RECT 127.600 161.600 128.400 166.200 ;
        RECT 135.600 161.600 136.400 170.000 ;
        RECT 141.200 161.600 142.000 166.200 ;
        RECT 144.400 161.600 145.200 166.200 ;
        RECT 150.000 161.600 150.800 170.200 ;
        RECT 154.800 161.600 155.600 170.000 ;
        RECT 160.400 161.600 161.200 166.200 ;
        RECT 163.600 161.600 164.400 166.200 ;
        RECT 169.200 161.600 170.000 170.200 ;
        RECT 174.000 161.600 175.000 168.800 ;
        RECT 180.200 162.200 181.200 168.800 ;
        RECT 180.200 161.600 181.000 162.200 ;
        RECT 183.600 161.600 184.400 170.200 ;
        RECT 187.800 161.600 188.600 166.200 ;
        RECT 190.000 161.600 190.800 166.200 ;
        RECT 193.200 161.600 194.000 166.200 ;
        RECT 194.800 161.600 195.600 170.200 ;
        RECT 199.000 161.600 199.800 166.200 ;
        RECT 204.400 161.600 205.200 169.000 ;
        RECT 209.200 161.600 210.000 166.200 ;
        RECT 210.800 161.600 211.600 170.200 ;
        RECT 215.000 161.600 215.800 166.200 ;
        RECT 217.800 161.600 218.600 166.200 ;
        RECT 222.000 161.600 222.800 170.200 ;
        RECT 223.600 161.600 224.400 166.200 ;
        RECT 226.800 161.600 227.600 166.200 ;
        RECT 228.400 161.600 229.200 166.200 ;
        RECT 231.600 161.600 232.400 166.200 ;
        RECT 234.800 161.600 235.600 170.000 ;
        RECT 240.400 161.600 241.200 166.200 ;
        RECT 243.600 161.600 244.400 166.200 ;
        RECT 249.200 161.600 250.000 170.200 ;
        RECT 252.400 161.600 253.200 170.200 ;
        RECT 255.600 161.600 256.400 170.200 ;
        RECT 258.800 161.600 259.600 170.200 ;
        RECT 262.000 161.600 262.800 170.200 ;
        RECT 265.200 161.600 266.000 170.200 ;
        RECT 268.400 161.600 269.200 170.000 ;
        RECT 274.000 161.600 274.800 166.200 ;
        RECT 277.200 161.600 278.000 166.200 ;
        RECT 282.800 161.600 283.600 170.200 ;
        RECT 292.400 161.600 293.200 170.000 ;
        RECT 298.000 161.600 298.800 166.200 ;
        RECT 301.200 161.600 302.000 166.200 ;
        RECT 306.800 161.600 307.600 170.200 ;
        RECT 310.000 161.600 310.800 166.200 ;
        RECT 313.200 161.600 314.000 166.200 ;
        RECT 314.800 161.600 315.600 170.200 ;
        RECT 319.000 161.600 319.800 166.200 ;
        RECT 321.200 161.600 322.000 166.200 ;
        RECT 324.400 161.600 325.200 166.200 ;
        RECT 326.600 161.600 327.400 166.200 ;
        RECT 330.800 161.600 331.600 170.200 ;
        RECT 333.000 161.600 333.800 166.200 ;
        RECT 337.200 161.600 338.000 170.200 ;
        RECT 340.400 161.600 341.200 166.200 ;
        RECT 342.000 161.600 342.800 170.200 ;
        RECT 346.200 161.600 347.000 166.200 ;
        RECT 348.400 161.600 349.200 166.200 ;
        RECT 351.600 161.600 352.400 166.200 ;
        RECT 356.400 161.600 357.200 170.200 ;
        RECT 358.000 161.600 358.800 170.200 ;
        RECT 364.400 161.600 365.200 166.200 ;
        RECT 369.200 161.600 370.000 170.200 ;
        RECT 374.000 161.600 374.800 169.000 ;
        RECT 377.200 161.600 378.000 170.200 ;
        RECT 382.000 161.600 382.800 166.200 ;
        RECT 385.200 161.600 386.000 166.200 ;
        RECT 386.800 161.600 387.600 170.200 ;
        RECT 391.000 161.600 391.800 166.200 ;
        RECT 393.200 161.600 394.000 166.200 ;
        RECT 396.400 161.600 397.200 166.200 ;
        RECT 399.600 161.600 400.400 166.200 ;
        RECT 401.800 161.600 402.600 166.200 ;
        RECT 406.000 161.600 406.800 170.200 ;
        RECT 409.200 161.600 410.000 166.200 ;
        RECT 410.800 161.600 411.600 170.200 ;
        RECT 415.000 161.600 415.800 166.200 ;
        RECT 417.200 161.600 418.000 166.200 ;
        RECT 420.400 161.600 421.200 166.200 ;
        RECT 423.600 161.600 424.400 170.000 ;
        RECT 429.200 161.600 430.000 166.200 ;
        RECT 432.400 161.600 433.200 166.200 ;
        RECT 438.000 161.600 438.800 170.200 ;
        RECT 447.600 162.200 448.600 168.800 ;
        RECT 447.800 161.600 448.600 162.200 ;
        RECT 453.800 161.600 454.800 168.800 ;
        RECT 458.800 161.600 459.600 170.000 ;
        RECT 464.400 161.600 465.200 166.200 ;
        RECT 467.600 161.600 468.400 166.200 ;
        RECT 473.200 161.600 474.000 170.200 ;
        RECT 478.000 161.600 478.800 170.200 ;
        RECT 481.200 162.200 482.200 168.800 ;
        RECT 481.400 161.600 482.200 162.200 ;
        RECT 487.400 161.600 488.400 168.800 ;
        RECT 490.800 161.600 491.600 170.200 ;
        RECT 494.000 161.600 494.800 170.200 ;
        RECT 498.200 161.600 499.000 166.200 ;
        RECT 501.000 161.600 501.800 166.200 ;
        RECT 505.200 161.600 506.000 170.200 ;
        RECT 506.800 161.600 507.600 166.200 ;
        RECT 510.000 161.600 510.800 166.200 ;
        RECT 516.400 161.600 517.200 169.000 ;
        RECT 520.200 161.600 521.000 166.200 ;
        RECT 524.400 161.600 525.200 170.200 ;
        RECT 529.200 161.600 530.000 170.200 ;
        RECT 530.800 161.600 531.600 166.200 ;
        RECT 534.000 161.600 534.800 166.200 ;
        RECT 537.200 161.600 538.000 165.800 ;
        RECT 540.400 161.600 541.200 166.200 ;
        RECT 542.000 161.600 542.800 170.200 ;
        RECT 546.800 161.600 547.600 166.200 ;
        RECT 550.000 161.600 550.800 165.800 ;
        RECT 556.400 161.600 557.200 170.200 ;
        RECT 559.600 161.600 560.400 170.000 ;
        RECT 565.200 161.600 566.000 166.200 ;
        RECT 568.400 161.600 569.200 166.200 ;
        RECT 574.000 161.600 574.800 170.200 ;
        RECT 578.800 161.600 579.600 169.000 ;
        RECT 0.400 160.400 586.800 161.600 ;
        RECT 1.200 155.800 2.000 160.400 ;
        RECT 4.400 152.200 5.200 160.400 ;
        RECT 10.200 151.800 11.000 160.400 ;
        RECT 14.000 151.800 14.800 160.400 ;
        RECT 18.200 155.800 19.000 160.400 ;
        RECT 23.600 153.000 24.400 160.400 ;
        RECT 30.000 153.000 30.800 160.400 ;
        RECT 33.800 155.800 34.600 160.400 ;
        RECT 38.000 151.800 38.800 160.400 ;
        RECT 39.600 151.800 40.400 160.400 ;
        RECT 43.800 155.800 44.600 160.400 ;
        RECT 46.000 155.800 46.800 160.400 ;
        RECT 49.200 155.800 50.000 160.400 ;
        RECT 50.800 155.800 51.600 160.400 ;
        RECT 54.000 155.800 54.800 160.400 ;
        RECT 55.600 151.800 56.400 160.400 ;
        RECT 59.800 155.800 60.600 160.400 ;
        RECT 62.000 151.800 62.800 160.400 ;
        RECT 66.200 155.800 67.000 160.400 ;
        RECT 70.000 153.200 71.000 160.400 ;
        RECT 76.200 159.800 77.000 160.400 ;
        RECT 76.200 153.200 77.200 159.800 ;
        RECT 81.200 153.000 82.000 160.400 ;
        RECT 89.200 153.000 90.000 160.400 ;
        RECT 97.200 155.800 98.000 160.400 ;
        RECT 98.800 151.800 99.600 160.400 ;
        RECT 103.600 155.800 104.400 160.400 ;
        RECT 106.800 155.800 107.600 160.400 ;
        RECT 110.000 155.800 110.800 160.400 ;
        RECT 113.200 153.200 114.200 160.400 ;
        RECT 119.400 159.800 120.200 160.400 ;
        RECT 119.400 153.200 120.400 159.800 ;
        RECT 124.400 153.000 125.200 160.400 ;
        RECT 130.800 153.000 131.600 160.400 ;
        RECT 143.600 153.200 144.600 160.400 ;
        RECT 149.800 159.800 150.600 160.400 ;
        RECT 149.800 153.200 150.800 159.800 ;
        RECT 154.800 152.000 155.600 160.400 ;
        RECT 160.400 155.800 161.200 160.400 ;
        RECT 163.600 155.800 164.400 160.400 ;
        RECT 169.200 151.800 170.000 160.400 ;
        RECT 172.400 151.800 173.200 160.400 ;
        RECT 175.600 151.800 176.400 160.400 ;
        RECT 178.800 151.800 179.600 160.400 ;
        RECT 182.000 151.800 182.800 160.400 ;
        RECT 185.200 151.800 186.000 160.400 ;
        RECT 188.600 159.800 189.400 160.400 ;
        RECT 188.400 153.200 189.400 159.800 ;
        RECT 194.600 153.200 195.600 160.400 ;
        RECT 199.800 159.800 200.600 160.400 ;
        RECT 199.600 153.200 200.600 159.800 ;
        RECT 205.800 153.200 206.800 160.400 ;
        RECT 209.200 155.800 210.000 160.400 ;
        RECT 212.400 155.800 213.200 160.400 ;
        RECT 215.600 153.200 216.600 160.400 ;
        RECT 221.800 159.800 222.600 160.400 ;
        RECT 221.800 153.200 222.800 159.800 ;
        RECT 228.400 151.800 229.200 160.400 ;
        RECT 231.600 155.800 232.400 160.400 ;
        RECT 234.800 153.200 235.800 160.400 ;
        RECT 241.000 159.800 241.800 160.400 ;
        RECT 241.000 153.200 242.000 159.800 ;
        RECT 247.000 151.800 247.800 160.400 ;
        RECT 250.800 155.800 251.600 160.400 ;
        RECT 254.000 155.800 254.800 160.400 ;
        RECT 255.600 155.800 256.400 160.400 ;
        RECT 258.800 155.800 259.600 160.400 ;
        RECT 260.400 151.800 261.200 160.400 ;
        RECT 265.200 155.800 266.000 160.400 ;
        RECT 268.400 152.200 269.200 160.400 ;
        RECT 272.200 155.800 273.000 160.400 ;
        RECT 276.400 151.800 277.200 160.400 ;
        RECT 279.600 153.200 280.600 160.400 ;
        RECT 285.800 159.800 286.600 160.400 ;
        RECT 285.800 153.200 286.800 159.800 ;
        RECT 295.600 152.000 296.400 160.400 ;
        RECT 301.200 155.800 302.000 160.400 ;
        RECT 304.400 155.800 305.200 160.400 ;
        RECT 310.000 151.800 310.800 160.400 ;
        RECT 314.800 152.000 315.600 160.400 ;
        RECT 320.400 155.800 321.200 160.400 ;
        RECT 323.600 155.800 324.400 160.400 ;
        RECT 329.200 151.800 330.000 160.400 ;
        RECT 332.400 151.800 333.200 160.400 ;
        RECT 335.600 151.800 336.400 160.400 ;
        RECT 338.800 151.800 339.600 160.400 ;
        RECT 342.000 151.800 342.800 160.400 ;
        RECT 345.200 151.800 346.000 160.400 ;
        RECT 346.800 151.800 347.600 160.400 ;
        RECT 351.000 155.800 351.800 160.400 ;
        RECT 353.800 155.800 354.600 160.400 ;
        RECT 358.000 151.800 358.800 160.400 ;
        RECT 361.200 155.800 362.000 160.400 ;
        RECT 362.800 151.800 363.600 160.400 ;
        RECT 367.000 155.800 367.800 160.400 ;
        RECT 369.200 151.800 370.000 160.400 ;
        RECT 373.400 155.800 374.200 160.400 ;
        RECT 375.600 151.800 376.400 160.400 ;
        RECT 379.800 155.800 380.600 160.400 ;
        RECT 382.600 155.800 383.400 160.400 ;
        RECT 386.800 151.800 387.600 160.400 ;
        RECT 389.000 155.800 389.800 160.400 ;
        RECT 393.200 151.800 394.000 160.400 ;
        RECT 394.800 155.800 395.600 160.400 ;
        RECT 402.800 153.000 403.600 160.400 ;
        RECT 407.600 153.000 408.400 160.400 ;
        RECT 415.600 152.200 416.400 160.400 ;
        RECT 420.800 151.800 421.600 160.400 ;
        RECT 425.200 153.000 426.000 160.400 ;
        RECT 431.600 155.800 432.400 160.400 ;
        RECT 433.200 155.800 434.000 160.400 ;
        RECT 437.000 155.800 437.800 160.400 ;
        RECT 441.200 151.800 442.000 160.400 ;
        RECT 449.200 155.800 450.000 160.400 ;
        RECT 452.400 153.000 453.200 160.400 ;
        RECT 457.200 151.800 458.000 160.400 ;
        RECT 461.400 155.800 462.200 160.400 ;
        RECT 463.600 155.800 464.400 160.400 ;
        RECT 466.800 155.800 467.600 160.400 ;
        RECT 470.000 152.000 470.800 160.400 ;
        RECT 475.600 155.800 476.400 160.400 ;
        RECT 478.800 155.800 479.600 160.400 ;
        RECT 484.400 151.800 485.200 160.400 ;
        RECT 487.600 151.800 488.400 160.400 ;
        RECT 490.800 151.800 491.600 160.400 ;
        RECT 494.000 151.800 494.800 160.400 ;
        RECT 497.200 151.800 498.000 160.400 ;
        RECT 500.400 151.800 501.200 160.400 ;
        RECT 502.000 155.800 502.800 160.400 ;
        RECT 505.200 155.800 506.000 160.400 ;
        RECT 511.600 153.000 512.400 160.400 ;
        RECT 514.800 151.800 515.600 160.400 ;
        RECT 519.000 155.800 519.800 160.400 ;
        RECT 521.200 155.800 522.000 160.400 ;
        RECT 524.400 155.800 525.200 160.400 ;
        RECT 526.000 151.800 526.800 160.400 ;
        RECT 530.200 155.800 531.000 160.400 ;
        RECT 532.400 151.800 533.200 160.400 ;
        RECT 538.800 156.200 539.600 160.400 ;
        RECT 542.000 155.800 542.800 160.400 ;
        RECT 543.600 155.800 544.400 160.400 ;
        RECT 546.800 155.800 547.600 160.400 ;
        RECT 551.600 151.800 552.400 160.400 ;
        RECT 555.000 159.800 555.800 160.400 ;
        RECT 554.800 153.200 555.800 159.800 ;
        RECT 561.000 153.200 562.000 160.400 ;
        RECT 566.000 152.000 566.800 160.400 ;
        RECT 571.600 155.800 572.400 160.400 ;
        RECT 574.800 155.800 575.600 160.400 ;
        RECT 580.400 151.800 581.200 160.400 ;
        RECT 554.800 131.600 555.600 133.200 ;
        RECT 578.800 131.600 579.600 133.200 ;
        RECT 1.200 121.600 2.000 126.200 ;
        RECT 7.600 121.600 8.400 130.200 ;
        RECT 9.200 121.600 10.000 130.200 ;
        RECT 13.400 121.600 14.200 126.200 ;
        RECT 15.600 121.600 16.400 130.200 ;
        RECT 20.400 121.600 21.200 130.200 ;
        RECT 28.400 121.600 29.200 130.200 ;
        RECT 33.200 121.600 34.000 130.200 ;
        RECT 34.800 121.600 35.600 126.200 ;
        RECT 38.000 121.600 38.800 126.200 ;
        RECT 41.200 121.600 42.000 126.200 ;
        RECT 42.800 121.600 43.600 126.200 ;
        RECT 46.000 121.600 46.800 126.200 ;
        RECT 47.600 121.600 48.400 126.200 ;
        RECT 50.800 121.600 51.600 126.200 ;
        RECT 52.400 121.600 53.200 130.200 ;
        RECT 56.600 121.600 57.400 126.200 ;
        RECT 58.800 121.600 59.600 126.200 ;
        RECT 62.000 121.600 62.800 126.200 ;
        RECT 65.200 121.600 66.000 130.200 ;
        RECT 68.000 121.600 68.800 130.200 ;
        RECT 73.200 121.600 74.000 129.800 ;
        RECT 76.400 121.600 77.200 130.200 ;
        RECT 80.600 121.600 81.400 126.200 ;
        RECT 83.400 121.600 84.200 126.200 ;
        RECT 87.600 121.600 88.400 130.200 ;
        RECT 90.800 121.600 91.600 126.200 ;
        RECT 92.400 121.600 93.200 130.200 ;
        RECT 96.600 121.600 97.400 126.200 ;
        RECT 99.400 121.600 100.200 126.200 ;
        RECT 103.600 121.600 104.400 130.200 ;
        RECT 105.200 121.600 106.000 126.200 ;
        RECT 108.400 121.600 109.200 126.200 ;
        RECT 110.600 121.600 111.400 126.200 ;
        RECT 114.800 121.600 115.600 130.200 ;
        RECT 116.400 121.600 117.200 126.200 ;
        RECT 119.600 121.600 120.400 126.200 ;
        RECT 121.800 121.600 122.600 126.200 ;
        RECT 126.000 121.600 126.800 130.200 ;
        RECT 127.600 121.600 128.400 126.200 ;
        RECT 130.800 121.600 131.600 126.200 ;
        RECT 138.800 121.600 139.800 128.800 ;
        RECT 145.000 122.200 146.000 128.800 ;
        RECT 150.000 122.200 151.000 128.800 ;
        RECT 145.000 121.600 145.800 122.200 ;
        RECT 150.200 121.600 151.000 122.200 ;
        RECT 156.200 121.600 157.200 128.800 ;
        RECT 161.200 121.600 162.000 130.000 ;
        RECT 166.800 121.600 167.600 126.200 ;
        RECT 170.000 121.600 170.800 126.200 ;
        RECT 175.600 121.600 176.400 130.200 ;
        RECT 178.800 121.600 179.600 126.200 ;
        RECT 182.000 121.600 182.800 126.200 ;
        RECT 183.600 121.600 184.400 126.200 ;
        RECT 186.800 121.600 187.600 126.200 ;
        RECT 188.400 121.600 189.200 126.200 ;
        RECT 191.600 121.600 192.400 130.200 ;
        RECT 195.800 121.600 196.600 126.200 ;
        RECT 198.000 121.600 198.800 126.200 ;
        RECT 201.200 121.600 202.000 126.200 ;
        RECT 206.000 121.600 206.800 130.200 ;
        RECT 208.200 121.600 209.000 126.200 ;
        RECT 212.400 121.600 213.200 130.200 ;
        RECT 214.000 121.600 214.800 130.200 ;
        RECT 218.200 121.600 219.000 126.200 ;
        RECT 221.000 121.600 221.800 126.200 ;
        RECT 225.200 121.600 226.000 130.200 ;
        RECT 226.800 121.600 227.600 130.200 ;
        RECT 231.000 121.600 231.800 126.200 ;
        RECT 233.200 121.600 234.000 130.200 ;
        RECT 237.400 121.600 238.200 126.200 ;
        RECT 240.800 121.600 241.600 130.200 ;
        RECT 246.000 121.600 246.800 129.800 ;
        RECT 250.800 121.600 251.600 129.000 ;
        RECT 255.600 121.600 256.400 130.200 ;
        RECT 260.400 121.600 261.200 126.200 ;
        RECT 263.600 121.600 264.400 130.200 ;
        RECT 267.800 121.600 268.600 126.200 ;
        RECT 270.000 121.600 270.800 130.200 ;
        RECT 274.200 121.600 275.000 126.200 ;
        RECT 276.400 121.600 277.200 126.200 ;
        RECT 279.600 121.600 280.400 126.200 ;
        RECT 281.200 121.600 282.000 126.200 ;
        RECT 284.400 121.600 285.200 130.200 ;
        RECT 288.600 121.600 289.400 126.200 ;
        RECT 297.200 121.600 298.200 128.800 ;
        RECT 303.400 122.200 304.400 128.800 ;
        RECT 303.400 121.600 304.200 122.200 ;
        RECT 308.400 121.600 309.200 130.000 ;
        RECT 314.000 121.600 314.800 126.200 ;
        RECT 317.200 121.600 318.000 126.200 ;
        RECT 322.800 121.600 323.600 130.200 ;
        RECT 327.600 121.600 328.600 128.800 ;
        RECT 333.800 122.200 334.800 128.800 ;
        RECT 333.800 121.600 334.600 122.200 ;
        RECT 338.800 121.600 339.800 128.800 ;
        RECT 345.000 122.200 346.000 128.800 ;
        RECT 350.000 122.200 351.000 128.800 ;
        RECT 345.000 121.600 345.800 122.200 ;
        RECT 350.200 121.600 351.000 122.200 ;
        RECT 356.200 121.600 357.200 128.800 ;
        RECT 359.600 121.600 360.400 126.200 ;
        RECT 362.800 121.600 363.600 126.200 ;
        RECT 364.400 121.600 365.200 126.200 ;
        RECT 367.600 121.600 368.400 126.200 ;
        RECT 369.200 121.600 370.000 126.200 ;
        RECT 372.400 121.600 373.200 126.200 ;
        RECT 375.600 121.600 376.400 126.200 ;
        RECT 377.200 121.600 378.000 126.200 ;
        RECT 380.400 121.600 381.200 126.200 ;
        RECT 383.600 121.600 384.400 126.200 ;
        RECT 385.200 121.600 386.000 126.200 ;
        RECT 388.400 121.600 389.200 126.200 ;
        RECT 390.000 121.600 390.800 126.200 ;
        RECT 393.200 121.600 394.000 126.200 ;
        RECT 398.000 121.600 398.800 130.200 ;
        RECT 404.400 121.600 405.200 129.000 ;
        RECT 409.200 121.600 410.000 129.000 ;
        RECT 418.800 121.600 419.600 130.200 ;
        RECT 422.000 121.600 423.000 128.800 ;
        RECT 428.200 122.200 429.200 128.800 ;
        RECT 428.200 121.600 429.000 122.200 ;
        RECT 432.200 121.600 433.000 126.200 ;
        RECT 436.400 121.600 437.200 130.200 ;
        RECT 438.000 121.600 438.800 130.200 ;
        RECT 447.600 121.600 448.400 130.200 ;
        RECT 452.400 121.600 453.200 130.200 ;
        RECT 457.200 121.600 458.000 130.200 ;
        RECT 461.400 121.600 462.200 126.200 ;
        RECT 463.600 121.600 464.400 126.200 ;
        RECT 466.800 121.600 467.600 130.200 ;
        RECT 471.000 121.600 471.800 126.200 ;
        RECT 473.200 121.600 474.000 126.200 ;
        RECT 476.400 121.600 477.200 125.800 ;
        RECT 481.200 121.600 482.000 130.200 ;
        RECT 486.800 121.600 487.600 126.200 ;
        RECT 490.000 121.600 490.800 126.200 ;
        RECT 495.600 121.600 496.400 130.000 ;
        RECT 498.800 121.600 499.600 130.200 ;
        RECT 502.000 121.600 502.800 130.200 ;
        RECT 505.200 121.600 506.000 130.200 ;
        RECT 508.400 121.600 509.200 130.200 ;
        RECT 511.600 121.600 512.400 130.200 ;
        RECT 513.200 121.600 514.000 126.200 ;
        RECT 516.400 121.600 517.200 126.200 ;
        RECT 518.000 121.600 518.800 126.200 ;
        RECT 521.200 121.600 522.000 126.200 ;
        RECT 522.800 121.600 523.600 126.200 ;
        RECT 526.000 121.600 526.800 126.200 ;
        RECT 527.600 121.600 528.400 130.200 ;
        RECT 530.800 121.600 531.600 130.200 ;
        RECT 532.400 121.600 533.200 126.200 ;
        RECT 535.600 121.600 536.400 126.200 ;
        RECT 538.800 121.600 539.600 126.200 ;
        RECT 540.400 121.600 541.200 126.200 ;
        RECT 543.600 121.600 544.400 126.200 ;
        RECT 547.400 121.600 548.200 130.200 ;
        RECT 553.200 121.600 554.000 129.000 ;
        RECT 558.000 121.600 559.000 128.800 ;
        RECT 564.200 122.200 565.200 128.800 ;
        RECT 564.200 121.600 565.000 122.200 ;
        RECT 569.200 121.600 570.200 128.800 ;
        RECT 575.400 122.200 576.400 128.800 ;
        RECT 575.400 121.600 576.200 122.200 ;
        RECT 580.400 121.600 581.200 129.000 ;
        RECT 0.400 120.400 586.800 121.600 ;
        RECT 1.200 111.800 2.000 120.400 ;
        RECT 5.400 115.800 6.200 120.400 ;
        RECT 9.200 113.000 10.000 120.400 ;
        RECT 18.800 113.000 19.600 120.400 ;
        RECT 23.800 119.800 24.600 120.400 ;
        RECT 23.600 113.200 24.600 119.800 ;
        RECT 29.800 113.200 30.800 120.400 ;
        RECT 33.200 111.800 34.000 120.400 ;
        RECT 38.000 111.800 38.800 120.400 ;
        RECT 41.200 111.800 42.000 120.400 ;
        RECT 45.400 115.800 46.200 120.400 ;
        RECT 47.600 111.800 48.400 120.400 ;
        RECT 54.000 115.800 54.800 120.400 ;
        RECT 56.200 115.800 57.000 120.400 ;
        RECT 60.400 111.800 61.200 120.400 ;
        RECT 62.000 115.800 62.800 120.400 ;
        RECT 68.400 113.000 69.200 120.400 ;
        RECT 73.200 113.200 74.200 120.400 ;
        RECT 79.400 119.800 80.200 120.400 ;
        RECT 79.400 113.200 80.400 119.800 ;
        RECT 82.800 115.800 83.600 120.400 ;
        RECT 86.000 112.200 86.800 120.400 ;
        RECT 89.200 115.800 90.000 120.400 ;
        RECT 92.400 115.800 93.200 120.400 ;
        RECT 94.000 111.800 94.800 120.400 ;
        RECT 102.000 111.800 102.800 120.400 ;
        RECT 103.600 111.800 104.400 120.400 ;
        RECT 107.800 115.800 108.600 120.400 ;
        RECT 110.000 111.800 110.800 120.400 ;
        RECT 114.200 115.800 115.000 120.400 ;
        RECT 116.400 111.800 117.200 120.400 ;
        RECT 120.600 115.800 121.400 120.400 ;
        RECT 122.800 111.800 123.600 120.400 ;
        RECT 127.600 115.800 128.400 120.400 ;
        RECT 132.400 113.000 133.200 120.400 ;
        RECT 143.600 115.800 144.400 120.400 ;
        RECT 145.200 111.800 146.000 120.400 ;
        RECT 151.800 119.800 152.600 120.400 ;
        RECT 151.600 113.200 152.600 119.800 ;
        RECT 157.800 113.200 158.800 120.400 ;
        RECT 162.800 115.800 163.600 120.400 ;
        RECT 166.000 112.000 166.800 120.400 ;
        RECT 171.600 115.800 172.400 120.400 ;
        RECT 174.800 115.800 175.600 120.400 ;
        RECT 180.400 111.800 181.200 120.400 ;
        RECT 183.600 111.800 184.400 120.400 ;
        RECT 186.800 111.800 187.600 120.400 ;
        RECT 188.400 115.800 189.200 120.400 ;
        RECT 191.600 115.800 192.400 120.400 ;
        RECT 193.200 115.800 194.000 120.400 ;
        RECT 197.000 115.800 197.800 120.400 ;
        RECT 201.200 111.800 202.000 120.400 ;
        RECT 204.400 113.000 205.200 120.400 ;
        RECT 210.800 115.800 211.600 120.400 ;
        RECT 214.000 115.800 214.800 120.400 ;
        RECT 218.800 113.000 219.600 120.400 ;
        RECT 223.600 113.000 224.400 120.400 ;
        RECT 230.600 115.800 231.400 120.400 ;
        RECT 234.800 111.800 235.600 120.400 ;
        RECT 237.600 111.800 238.400 120.400 ;
        RECT 242.800 112.200 243.600 120.400 ;
        RECT 247.600 113.200 248.600 120.400 ;
        RECT 253.800 119.800 254.600 120.400 ;
        RECT 253.800 113.200 254.800 119.800 ;
        RECT 257.200 115.800 258.000 120.400 ;
        RECT 260.400 115.800 261.200 120.400 ;
        RECT 263.600 115.800 264.400 120.400 ;
        RECT 265.800 115.800 266.600 120.400 ;
        RECT 270.000 111.800 270.800 120.400 ;
        RECT 271.600 115.800 272.400 120.400 ;
        RECT 274.800 115.800 275.600 120.400 ;
        RECT 276.400 111.800 277.200 120.400 ;
        RECT 280.600 115.800 281.400 120.400 ;
        RECT 284.400 113.200 285.400 120.400 ;
        RECT 290.600 119.800 291.400 120.400 ;
        RECT 290.600 113.200 291.600 119.800 ;
        RECT 298.800 111.800 299.600 120.400 ;
        RECT 302.000 111.800 302.800 120.400 ;
        RECT 305.200 113.000 306.000 120.400 ;
        RECT 310.000 112.000 310.800 120.400 ;
        RECT 315.600 115.800 316.400 120.400 ;
        RECT 318.800 115.800 319.600 120.400 ;
        RECT 324.400 111.800 325.200 120.400 ;
        RECT 329.200 112.000 330.000 120.400 ;
        RECT 334.800 115.800 335.600 120.400 ;
        RECT 338.000 115.800 338.800 120.400 ;
        RECT 343.600 111.800 344.400 120.400 ;
        RECT 346.800 111.800 347.600 120.400 ;
        RECT 350.000 113.000 350.800 120.400 ;
        RECT 354.800 113.000 355.600 120.400 ;
        RECT 358.000 111.800 358.800 120.400 ;
        RECT 361.200 113.000 362.000 120.400 ;
        RECT 364.400 111.800 365.200 120.400 ;
        RECT 366.000 111.800 366.800 120.400 ;
        RECT 370.200 115.800 371.000 120.400 ;
        RECT 373.600 111.800 374.400 120.400 ;
        RECT 378.800 112.200 379.600 120.400 ;
        RECT 382.600 115.800 383.400 120.400 ;
        RECT 386.800 111.800 387.600 120.400 ;
        RECT 388.400 111.800 389.200 120.400 ;
        RECT 392.600 115.800 393.400 120.400 ;
        RECT 394.800 115.800 395.600 120.400 ;
        RECT 398.000 115.800 398.800 120.400 ;
        RECT 399.600 111.800 400.400 120.400 ;
        RECT 406.000 115.800 406.800 120.400 ;
        RECT 407.600 111.800 408.400 120.400 ;
        RECT 411.800 115.800 412.600 120.400 ;
        RECT 414.600 115.800 415.400 120.400 ;
        RECT 418.800 111.800 419.600 120.400 ;
        RECT 422.000 113.200 423.000 120.400 ;
        RECT 428.200 119.800 429.000 120.400 ;
        RECT 428.200 113.200 429.200 119.800 ;
        RECT 433.200 112.000 434.000 120.400 ;
        RECT 438.800 115.800 439.600 120.400 ;
        RECT 442.000 115.800 442.800 120.400 ;
        RECT 447.600 111.800 448.400 120.400 ;
        RECT 455.600 111.800 456.400 120.400 ;
        RECT 458.800 111.800 459.600 120.400 ;
        RECT 462.000 111.800 462.800 120.400 ;
        RECT 465.200 113.000 466.000 120.400 ;
        RECT 470.000 113.200 471.000 120.400 ;
        RECT 476.200 119.800 477.000 120.400 ;
        RECT 476.200 113.200 477.200 119.800 ;
        RECT 479.600 111.800 480.400 120.400 ;
        RECT 482.800 111.800 483.600 120.400 ;
        RECT 486.000 112.000 486.800 120.400 ;
        RECT 491.600 115.800 492.400 120.400 ;
        RECT 494.800 115.800 495.600 120.400 ;
        RECT 500.400 111.800 501.200 120.400 ;
        RECT 505.200 112.000 506.000 120.400 ;
        RECT 510.800 115.800 511.600 120.400 ;
        RECT 514.000 115.800 514.800 120.400 ;
        RECT 519.600 111.800 520.400 120.400 ;
        RECT 524.600 119.800 525.400 120.400 ;
        RECT 524.400 113.200 525.400 119.800 ;
        RECT 530.600 113.200 531.600 120.400 ;
        RECT 535.800 119.800 536.600 120.400 ;
        RECT 535.600 113.200 536.600 119.800 ;
        RECT 541.800 113.200 542.800 120.400 ;
        RECT 546.800 112.000 547.600 120.400 ;
        RECT 552.400 115.800 553.200 120.400 ;
        RECT 555.600 115.800 556.400 120.400 ;
        RECT 561.200 111.800 562.000 120.400 ;
        RECT 566.000 112.000 566.800 120.400 ;
        RECT 571.600 115.800 572.400 120.400 ;
        RECT 574.800 115.800 575.600 120.400 ;
        RECT 580.400 111.800 581.200 120.400 ;
        RECT 1.200 81.600 2.000 90.200 ;
        RECT 4.400 81.600 5.200 86.200 ;
        RECT 7.600 81.600 8.400 86.200 ;
        RECT 10.800 81.600 11.600 85.800 ;
        RECT 14.000 81.600 14.800 90.200 ;
        RECT 18.200 81.600 19.000 86.200 ;
        RECT 20.400 81.600 21.200 90.200 ;
        RECT 23.600 81.600 24.400 89.000 ;
        RECT 26.800 81.600 27.600 90.200 ;
        RECT 31.600 81.600 32.400 86.200 ;
        RECT 34.800 81.600 35.600 90.200 ;
        RECT 39.000 81.600 39.800 86.200 ;
        RECT 41.200 81.600 42.000 86.200 ;
        RECT 45.000 81.600 45.800 86.200 ;
        RECT 49.200 81.600 50.000 90.200 ;
        RECT 50.800 81.600 51.600 86.200 ;
        RECT 54.000 81.600 54.800 86.200 ;
        RECT 57.200 81.600 58.000 85.800 ;
        RECT 63.600 81.600 64.400 89.000 ;
        RECT 66.800 81.600 67.600 90.200 ;
        RECT 71.000 81.600 71.800 86.200 ;
        RECT 73.200 81.600 74.000 86.200 ;
        RECT 76.400 81.600 77.200 86.200 ;
        RECT 78.000 81.600 78.800 86.200 ;
        RECT 81.200 81.600 82.000 86.200 ;
        RECT 84.400 81.600 85.200 86.200 ;
        RECT 86.000 81.600 86.800 86.200 ;
        RECT 89.200 81.600 90.000 86.200 ;
        RECT 90.800 81.600 91.600 86.200 ;
        RECT 94.000 81.600 94.800 86.200 ;
        RECT 97.200 81.600 98.000 89.000 ;
        RECT 103.600 81.600 104.400 89.000 ;
        RECT 110.000 81.600 110.800 89.000 ;
        RECT 114.800 81.600 115.600 86.200 ;
        RECT 118.600 81.600 119.400 86.200 ;
        RECT 122.800 81.600 123.600 90.200 ;
        RECT 127.600 81.600 128.400 89.000 ;
        RECT 130.800 81.600 131.600 90.200 ;
        RECT 141.000 81.600 141.800 86.200 ;
        RECT 145.200 81.600 146.000 90.200 ;
        RECT 147.400 81.600 148.200 86.200 ;
        RECT 151.600 81.600 152.400 90.200 ;
        RECT 153.200 81.600 154.000 86.200 ;
        RECT 156.400 81.600 157.200 86.200 ;
        RECT 159.600 81.600 160.400 90.000 ;
        RECT 165.200 81.600 166.000 86.200 ;
        RECT 168.400 81.600 169.200 86.200 ;
        RECT 174.000 81.600 174.800 90.200 ;
        RECT 180.400 81.600 181.200 90.200 ;
        RECT 182.000 81.600 182.800 90.200 ;
        RECT 190.000 81.600 190.800 90.200 ;
        RECT 191.600 81.600 192.400 90.200 ;
        RECT 196.400 81.600 197.200 90.200 ;
        RECT 200.600 81.600 201.400 86.200 ;
        RECT 203.400 81.600 204.200 86.200 ;
        RECT 207.600 81.600 208.400 90.200 ;
        RECT 209.200 81.600 210.000 86.200 ;
        RECT 217.200 81.600 218.000 89.000 ;
        RECT 220.400 81.600 221.200 86.200 ;
        RECT 223.600 81.600 224.400 86.200 ;
        RECT 225.800 81.600 226.600 86.200 ;
        RECT 230.000 81.600 230.800 90.200 ;
        RECT 233.200 81.600 234.000 86.200 ;
        RECT 236.400 81.600 237.200 89.000 ;
        RECT 242.800 81.600 243.600 90.200 ;
        RECT 249.200 81.600 250.000 89.800 ;
        RECT 254.400 81.600 255.200 90.200 ;
        RECT 258.800 81.600 259.800 88.800 ;
        RECT 265.000 82.200 266.000 88.800 ;
        RECT 265.000 81.600 265.800 82.200 ;
        RECT 268.400 81.600 269.200 86.200 ;
        RECT 271.600 81.600 272.400 86.200 ;
        RECT 274.800 81.600 275.600 86.200 ;
        RECT 276.400 81.600 277.200 90.200 ;
        RECT 279.600 81.600 280.400 89.000 ;
        RECT 282.800 81.600 283.600 86.200 ;
        RECT 286.000 81.600 286.800 86.200 ;
        RECT 293.000 81.600 293.800 86.200 ;
        RECT 297.200 81.600 298.000 90.200 ;
        RECT 298.800 81.600 299.600 86.200 ;
        RECT 302.000 81.600 302.800 86.200 ;
        RECT 303.600 81.600 304.400 86.200 ;
        RECT 306.800 81.600 307.600 86.200 ;
        RECT 310.000 81.600 310.800 86.200 ;
        RECT 313.200 81.600 314.000 90.000 ;
        RECT 318.800 81.600 319.600 86.200 ;
        RECT 322.000 81.600 322.800 86.200 ;
        RECT 327.600 81.600 328.400 90.200 ;
        RECT 332.400 81.600 333.200 90.000 ;
        RECT 338.000 81.600 338.800 86.200 ;
        RECT 341.200 81.600 342.000 86.200 ;
        RECT 346.800 81.600 347.600 90.200 ;
        RECT 351.600 81.600 352.400 89.000 ;
        RECT 354.800 81.600 355.600 90.200 ;
        RECT 359.000 81.600 359.800 90.200 ;
        RECT 362.800 81.600 363.600 86.200 ;
        RECT 366.000 81.600 366.800 86.200 ;
        RECT 369.200 81.600 370.200 88.800 ;
        RECT 375.400 82.200 376.400 88.800 ;
        RECT 375.400 81.600 376.200 82.200 ;
        RECT 378.800 81.600 379.600 90.200 ;
        RECT 383.600 81.600 384.400 90.200 ;
        RECT 387.800 81.600 388.600 86.200 ;
        RECT 391.600 81.600 392.400 89.000 ;
        RECT 396.400 81.600 397.200 86.200 ;
        RECT 399.600 81.600 400.400 89.800 ;
        RECT 402.800 81.600 403.600 90.200 ;
        RECT 407.000 81.600 407.800 86.200 ;
        RECT 409.200 81.600 410.000 86.200 ;
        RECT 412.400 81.600 413.200 86.200 ;
        RECT 415.600 81.600 416.400 89.000 ;
        RECT 419.400 81.600 420.200 86.200 ;
        RECT 423.600 81.600 424.400 90.200 ;
        RECT 425.800 81.600 426.600 86.200 ;
        RECT 430.000 81.600 430.800 90.200 ;
        RECT 433.200 81.600 434.000 90.000 ;
        RECT 438.800 81.600 439.600 86.200 ;
        RECT 442.000 81.600 442.800 86.200 ;
        RECT 447.600 81.600 448.400 90.200 ;
        RECT 457.200 81.600 458.200 88.800 ;
        RECT 463.400 82.200 464.400 88.800 ;
        RECT 468.400 82.200 469.400 88.800 ;
        RECT 463.400 81.600 464.200 82.200 ;
        RECT 468.600 81.600 469.400 82.200 ;
        RECT 474.600 81.600 475.600 88.800 ;
        RECT 478.000 81.600 478.800 86.200 ;
        RECT 481.200 81.600 482.000 86.200 ;
        RECT 484.400 81.600 485.200 85.800 ;
        RECT 487.600 81.600 488.400 86.200 ;
        RECT 490.800 81.600 491.600 86.200 ;
        RECT 494.000 81.600 494.800 90.000 ;
        RECT 499.600 81.600 500.400 86.200 ;
        RECT 502.800 81.600 503.600 86.200 ;
        RECT 508.400 81.600 509.200 90.200 ;
        RECT 513.200 81.600 514.000 90.200 ;
        RECT 518.800 81.600 519.600 86.200 ;
        RECT 522.000 81.600 522.800 86.200 ;
        RECT 527.600 81.600 528.400 90.000 ;
        RECT 532.400 81.600 533.200 90.000 ;
        RECT 538.000 81.600 538.800 86.200 ;
        RECT 541.200 81.600 542.000 86.200 ;
        RECT 546.800 81.600 547.600 90.200 ;
        RECT 551.600 81.600 552.400 90.200 ;
        RECT 554.800 81.600 555.600 90.000 ;
        RECT 560.400 81.600 561.200 86.200 ;
        RECT 563.600 81.600 564.400 86.200 ;
        RECT 569.200 81.600 570.000 90.200 ;
        RECT 574.000 81.600 574.800 89.000 ;
        RECT 578.800 81.600 579.600 89.000 ;
        RECT 0.400 80.400 586.800 81.600 ;
        RECT 3.000 79.800 3.800 80.400 ;
        RECT 2.800 73.200 3.800 79.800 ;
        RECT 9.000 73.200 10.000 80.400 ;
        RECT 12.400 75.800 13.200 80.400 ;
        RECT 15.600 75.800 16.400 80.400 ;
        RECT 17.200 71.800 18.000 80.400 ;
        RECT 21.400 75.800 22.200 80.400 ;
        RECT 23.600 75.800 24.400 80.400 ;
        RECT 26.800 75.800 27.600 80.400 ;
        RECT 29.000 75.800 29.800 80.400 ;
        RECT 33.200 71.800 34.000 80.400 ;
        RECT 36.400 71.800 37.200 80.400 ;
        RECT 38.000 71.800 38.800 80.400 ;
        RECT 42.800 71.800 43.600 80.400 ;
        RECT 47.000 75.800 47.800 80.400 ;
        RECT 50.800 75.800 51.600 80.400 ;
        RECT 55.600 71.800 56.400 80.400 ;
        RECT 60.400 71.800 61.200 80.400 ;
        RECT 62.000 71.800 62.800 80.400 ;
        RECT 66.200 75.800 67.000 80.400 ;
        RECT 68.400 71.800 69.200 80.400 ;
        RECT 71.600 71.800 72.400 80.400 ;
        RECT 74.800 71.800 75.600 80.400 ;
        RECT 76.400 75.800 77.200 80.400 ;
        RECT 81.200 73.000 82.000 80.400 ;
        RECT 84.400 71.800 85.200 80.400 ;
        RECT 86.000 75.800 86.800 80.400 ;
        RECT 89.200 75.800 90.000 80.400 ;
        RECT 92.400 75.800 93.200 80.400 ;
        RECT 94.000 75.800 94.800 80.400 ;
        RECT 97.200 75.800 98.000 80.400 ;
        RECT 98.800 75.800 99.600 80.400 ;
        RECT 102.000 75.800 102.800 80.400 ;
        RECT 103.600 71.800 104.400 80.400 ;
        RECT 107.800 75.800 108.600 80.400 ;
        RECT 113.200 71.800 114.000 80.400 ;
        RECT 118.000 73.000 118.800 80.400 ;
        RECT 121.200 71.800 122.000 80.400 ;
        RECT 125.400 75.800 126.200 80.400 ;
        RECT 127.600 75.800 128.400 80.400 ;
        RECT 130.800 75.800 131.600 80.400 ;
        RECT 133.000 75.800 133.800 80.400 ;
        RECT 137.200 71.800 138.000 80.400 ;
        RECT 145.200 73.200 146.200 80.400 ;
        RECT 151.400 79.800 152.200 80.400 ;
        RECT 151.400 73.200 152.400 79.800 ;
        RECT 156.400 72.000 157.200 80.400 ;
        RECT 162.000 75.800 162.800 80.400 ;
        RECT 165.200 75.800 166.000 80.400 ;
        RECT 170.800 71.800 171.600 80.400 ;
        RECT 174.000 71.800 174.800 80.400 ;
        RECT 178.200 75.800 179.000 80.400 ;
        RECT 180.400 75.800 181.200 80.400 ;
        RECT 186.800 71.800 187.600 80.400 ;
        RECT 188.400 75.800 189.200 80.400 ;
        RECT 191.600 75.800 192.400 80.400 ;
        RECT 196.400 71.800 197.200 80.400 ;
        RECT 198.000 71.800 198.800 80.400 ;
        RECT 202.200 75.800 203.000 80.400 ;
        RECT 206.000 75.800 206.800 80.400 ;
        RECT 208.200 75.800 209.000 80.400 ;
        RECT 212.400 71.800 213.200 80.400 ;
        RECT 217.200 73.000 218.000 80.400 ;
        RECT 220.400 75.800 221.200 80.400 ;
        RECT 223.600 75.800 224.400 80.400 ;
        RECT 226.800 71.800 227.600 80.400 ;
        RECT 231.000 75.800 231.800 80.400 ;
        RECT 234.800 75.800 235.600 80.400 ;
        RECT 239.600 73.000 240.400 80.400 ;
        RECT 244.400 76.200 245.200 80.400 ;
        RECT 247.600 75.800 248.400 80.400 ;
        RECT 249.200 71.800 250.000 80.400 ;
        RECT 253.400 75.800 254.200 80.400 ;
        RECT 255.600 75.800 256.400 80.400 ;
        RECT 258.800 75.800 259.600 80.400 ;
        RECT 262.000 75.800 262.800 80.400 ;
        RECT 263.600 75.800 264.400 80.400 ;
        RECT 266.800 71.800 267.600 80.400 ;
        RECT 271.000 75.800 271.800 80.400 ;
        RECT 273.800 75.800 274.600 80.400 ;
        RECT 278.000 71.800 278.800 80.400 ;
        RECT 279.600 71.800 280.400 80.400 ;
        RECT 284.400 75.800 285.200 80.400 ;
        RECT 287.600 76.200 288.400 80.400 ;
        RECT 295.600 75.800 296.400 80.400 ;
        RECT 299.400 75.800 300.200 80.400 ;
        RECT 303.600 71.800 304.400 80.400 ;
        RECT 306.800 75.800 307.600 80.400 ;
        RECT 308.400 71.800 309.200 80.400 ;
        RECT 312.600 75.800 313.400 80.400 ;
        RECT 316.400 75.800 317.200 80.400 ;
        RECT 321.200 73.000 322.000 80.400 ;
        RECT 327.600 71.800 328.400 80.400 ;
        RECT 330.800 75.800 331.600 80.400 ;
        RECT 334.000 73.200 335.000 80.400 ;
        RECT 340.200 79.800 341.000 80.400 ;
        RECT 340.200 73.200 341.200 79.800 ;
        RECT 345.200 72.000 346.000 80.400 ;
        RECT 350.800 75.800 351.600 80.400 ;
        RECT 354.000 75.800 354.800 80.400 ;
        RECT 359.600 71.800 360.400 80.400 ;
        RECT 364.400 72.000 365.200 80.400 ;
        RECT 370.000 75.800 370.800 80.400 ;
        RECT 373.200 75.800 374.000 80.400 ;
        RECT 378.800 71.800 379.600 80.400 ;
        RECT 382.000 75.800 382.800 80.400 ;
        RECT 385.200 75.800 386.000 80.400 ;
        RECT 386.800 75.800 387.600 80.400 ;
        RECT 390.000 71.800 390.800 80.400 ;
        RECT 394.200 75.800 395.000 80.400 ;
        RECT 397.000 75.800 397.800 80.400 ;
        RECT 401.200 71.800 402.000 80.400 ;
        RECT 402.800 75.800 403.600 80.400 ;
        RECT 406.000 75.800 406.800 80.400 ;
        RECT 407.600 75.800 408.400 80.400 ;
        RECT 410.800 75.800 411.600 80.400 ;
        RECT 412.400 71.800 413.200 80.400 ;
        RECT 415.600 75.800 416.400 80.400 ;
        RECT 422.000 71.800 422.800 80.400 ;
        RECT 423.600 75.800 424.400 80.400 ;
        RECT 426.800 75.800 427.600 80.400 ;
        RECT 430.000 75.800 430.800 80.400 ;
        RECT 433.200 73.000 434.000 80.400 ;
        RECT 439.600 73.200 440.600 80.400 ;
        RECT 445.800 79.800 446.600 80.400 ;
        RECT 445.800 73.200 446.800 79.800 ;
        RECT 454.000 71.800 454.800 80.400 ;
        RECT 460.400 71.800 461.200 80.400 ;
        RECT 463.800 79.800 464.600 80.400 ;
        RECT 463.600 73.200 464.600 79.800 ;
        RECT 469.800 73.200 470.800 80.400 ;
        RECT 473.200 71.800 474.000 80.400 ;
        RECT 477.400 75.800 478.200 80.400 ;
        RECT 479.600 71.800 480.400 80.400 ;
        RECT 484.400 75.800 485.200 80.400 ;
        RECT 488.200 75.800 489.000 80.400 ;
        RECT 492.400 71.800 493.200 80.400 ;
        RECT 494.600 75.800 495.400 80.400 ;
        RECT 498.800 71.800 499.600 80.400 ;
        RECT 500.400 75.800 501.200 80.400 ;
        RECT 504.200 75.800 505.000 80.400 ;
        RECT 508.400 71.800 509.200 80.400 ;
        RECT 513.200 71.800 514.000 80.400 ;
        RECT 514.800 71.800 515.600 80.400 ;
        RECT 519.600 71.800 520.400 80.400 ;
        RECT 523.800 75.800 524.600 80.400 ;
        RECT 526.600 75.800 527.400 80.400 ;
        RECT 530.800 71.800 531.600 80.400 ;
        RECT 534.000 73.000 534.800 80.400 ;
        RECT 538.800 73.000 539.600 80.400 ;
        RECT 543.600 72.000 544.400 80.400 ;
        RECT 549.200 75.800 550.000 80.400 ;
        RECT 552.400 75.800 553.200 80.400 ;
        RECT 558.000 71.800 558.800 80.400 ;
        RECT 562.800 72.000 563.600 80.400 ;
        RECT 568.400 75.800 569.200 80.400 ;
        RECT 571.600 75.800 572.400 80.400 ;
        RECT 577.200 71.800 578.000 80.400 ;
        RECT 582.000 73.000 582.800 80.400 ;
        RECT 4.400 41.600 5.200 50.200 ;
        RECT 6.000 41.600 6.800 46.200 ;
        RECT 9.200 41.600 10.000 46.200 ;
        RECT 10.800 41.600 11.600 46.200 ;
        RECT 14.000 41.600 14.800 46.200 ;
        RECT 15.600 41.600 16.400 50.200 ;
        RECT 20.400 41.600 21.200 46.200 ;
        RECT 23.600 41.600 24.400 46.200 ;
        RECT 30.000 41.600 30.800 49.000 ;
        RECT 33.200 41.600 34.000 46.200 ;
        RECT 41.200 41.600 42.000 49.000 ;
        RECT 46.000 41.600 46.800 45.800 ;
        RECT 49.200 41.600 50.000 46.200 ;
        RECT 51.400 41.600 52.200 46.200 ;
        RECT 55.600 41.600 56.400 50.200 ;
        RECT 57.200 41.600 58.000 46.200 ;
        RECT 60.400 41.600 61.200 46.200 ;
        RECT 66.800 41.600 67.600 49.000 ;
        RECT 71.200 41.600 72.000 50.200 ;
        RECT 76.400 41.600 77.200 49.800 ;
        RECT 79.600 41.600 80.400 50.200 ;
        RECT 83.800 41.600 84.600 46.200 ;
        RECT 86.000 41.600 86.800 46.200 ;
        RECT 89.200 41.600 90.000 46.200 ;
        RECT 90.800 41.600 91.600 46.200 ;
        RECT 94.000 41.600 94.800 46.200 ;
        RECT 95.600 41.600 96.400 46.200 ;
        RECT 98.800 41.600 99.600 46.200 ;
        RECT 100.400 41.600 101.200 50.200 ;
        RECT 104.600 41.600 105.400 46.200 ;
        RECT 106.800 41.600 107.600 46.200 ;
        RECT 110.000 41.600 110.800 50.200 ;
        RECT 114.200 41.600 115.000 46.200 ;
        RECT 116.400 41.600 117.200 50.200 ;
        RECT 122.800 41.600 123.600 46.200 ;
        RECT 125.000 41.600 125.800 46.200 ;
        RECT 129.200 41.600 130.000 50.200 ;
        RECT 132.400 41.600 133.200 46.200 ;
        RECT 138.800 41.600 139.600 50.200 ;
        RECT 143.000 41.600 143.800 46.200 ;
        RECT 146.800 41.600 147.600 46.200 ;
        RECT 151.600 41.600 152.400 49.000 ;
        RECT 156.400 41.600 157.400 48.800 ;
        RECT 162.600 42.200 163.600 48.800 ;
        RECT 162.600 41.600 163.400 42.200 ;
        RECT 167.600 41.600 168.600 48.800 ;
        RECT 173.800 42.200 174.800 48.800 ;
        RECT 173.800 41.600 174.600 42.200 ;
        RECT 178.800 41.600 179.600 50.000 ;
        RECT 184.400 41.600 185.200 46.200 ;
        RECT 187.600 41.600 188.400 46.200 ;
        RECT 193.200 41.600 194.000 50.200 ;
        RECT 198.000 41.600 198.800 50.200 ;
        RECT 201.200 41.600 202.200 48.800 ;
        RECT 207.400 42.200 208.400 48.800 ;
        RECT 207.400 41.600 208.200 42.200 ;
        RECT 211.400 41.600 212.200 46.200 ;
        RECT 215.600 41.600 216.400 50.200 ;
        RECT 217.200 41.600 218.000 50.200 ;
        RECT 223.600 41.600 224.400 50.200 ;
        RECT 228.400 41.600 229.200 50.200 ;
        RECT 230.000 41.600 230.800 50.200 ;
        RECT 234.800 41.600 235.600 50.200 ;
        RECT 239.000 41.600 239.800 46.200 ;
        RECT 242.800 42.200 243.800 48.800 ;
        RECT 243.000 41.600 243.800 42.200 ;
        RECT 249.000 41.600 250.000 48.800 ;
        RECT 254.000 41.600 254.800 49.000 ;
        RECT 257.200 41.600 258.000 50.200 ;
        RECT 260.400 41.600 261.200 49.000 ;
        RECT 265.200 41.600 266.000 49.000 ;
        RECT 268.400 41.600 269.200 50.200 ;
        RECT 271.600 41.600 272.400 49.000 ;
        RECT 276.400 41.600 277.200 50.200 ;
        RECT 281.200 41.600 282.000 50.200 ;
        RECT 286.000 41.600 286.800 50.200 ;
        RECT 292.400 41.600 293.200 50.200 ;
        RECT 296.600 41.600 297.400 46.200 ;
        RECT 302.000 41.600 302.800 49.000 ;
        RECT 305.200 41.600 306.000 46.200 ;
        RECT 308.400 41.600 309.200 46.200 ;
        RECT 311.600 41.600 312.400 46.200 ;
        RECT 314.800 41.600 315.600 49.000 ;
        RECT 322.800 41.600 323.600 49.000 ;
        RECT 332.400 41.600 333.200 50.200 ;
        RECT 335.600 41.600 336.400 49.000 ;
        RECT 338.800 41.600 339.600 50.200 ;
        RECT 343.000 41.600 343.800 46.200 ;
        RECT 345.800 41.600 346.600 46.200 ;
        RECT 350.000 41.600 350.800 50.200 ;
        RECT 353.200 41.600 354.000 50.000 ;
        RECT 358.800 41.600 359.600 46.200 ;
        RECT 362.000 41.600 362.800 46.200 ;
        RECT 367.600 41.600 368.400 50.200 ;
        RECT 372.400 41.600 373.200 50.000 ;
        RECT 378.000 41.600 378.800 46.200 ;
        RECT 381.200 41.600 382.000 46.200 ;
        RECT 386.800 41.600 387.600 50.200 ;
        RECT 390.000 41.600 390.800 46.200 ;
        RECT 393.200 41.600 394.000 46.200 ;
        RECT 396.400 41.600 397.200 46.200 ;
        RECT 399.600 41.600 400.400 50.000 ;
        RECT 405.200 41.600 406.000 46.200 ;
        RECT 408.400 41.600 409.200 46.200 ;
        RECT 414.000 41.600 414.800 50.200 ;
        RECT 418.800 41.600 419.600 49.000 ;
        RECT 422.000 41.600 422.800 50.200 ;
        RECT 425.200 42.200 426.200 48.800 ;
        RECT 425.400 41.600 426.200 42.200 ;
        RECT 431.400 41.600 432.400 48.800 ;
        RECT 434.800 41.600 435.600 50.200 ;
        RECT 439.000 41.600 439.800 46.200 ;
        RECT 441.200 41.600 442.000 46.200 ;
        RECT 449.200 41.600 450.000 46.200 ;
        RECT 452.400 41.600 453.200 46.200 ;
        RECT 454.600 41.600 455.400 46.200 ;
        RECT 458.800 41.600 459.600 50.200 ;
        RECT 460.400 41.600 461.200 46.200 ;
        RECT 463.600 41.600 464.400 46.200 ;
        RECT 466.800 41.600 467.600 49.800 ;
        RECT 470.000 41.600 470.800 46.200 ;
        RECT 473.200 41.600 474.000 49.000 ;
        RECT 478.000 41.600 478.800 50.200 ;
        RECT 482.800 41.600 483.600 50.200 ;
        RECT 487.600 41.600 488.400 50.200 ;
        RECT 491.800 41.600 492.600 46.200 ;
        RECT 494.000 41.600 494.800 46.200 ;
        RECT 500.400 41.600 501.200 49.000 ;
        RECT 506.800 41.600 507.600 49.000 ;
        RECT 511.600 41.600 512.400 46.200 ;
        RECT 514.800 41.600 515.800 48.800 ;
        RECT 521.000 42.200 522.000 48.800 ;
        RECT 521.000 41.600 521.800 42.200 ;
        RECT 526.000 41.600 526.800 50.000 ;
        RECT 531.600 41.600 532.400 46.200 ;
        RECT 534.800 41.600 535.600 46.200 ;
        RECT 540.400 41.600 541.200 50.200 ;
        RECT 545.200 41.600 546.000 50.200 ;
        RECT 550.800 41.600 551.600 46.200 ;
        RECT 554.000 41.600 554.800 46.200 ;
        RECT 559.600 41.600 560.400 50.000 ;
        RECT 564.400 41.600 565.200 50.200 ;
        RECT 570.000 41.600 570.800 46.200 ;
        RECT 573.200 41.600 574.000 46.200 ;
        RECT 578.800 41.600 579.600 50.000 ;
        RECT 0.400 40.400 586.800 41.600 ;
        RECT 1.200 35.800 2.000 40.400 ;
        RECT 4.400 35.800 5.200 40.400 ;
        RECT 7.600 35.800 8.400 40.400 ;
        RECT 9.200 35.800 10.000 40.400 ;
        RECT 12.400 35.800 13.200 40.400 ;
        RECT 17.200 33.000 18.000 40.400 ;
        RECT 21.000 35.800 21.800 40.400 ;
        RECT 25.200 31.800 26.000 40.400 ;
        RECT 28.400 33.000 29.200 40.400 ;
        RECT 31.600 35.800 32.400 40.400 ;
        RECT 34.800 35.800 35.600 40.400 ;
        RECT 37.000 35.800 37.800 40.400 ;
        RECT 41.200 31.800 42.000 40.400 ;
        RECT 44.400 33.000 45.200 40.400 ;
        RECT 49.200 35.800 50.000 40.400 ;
        RECT 54.000 33.000 54.800 40.400 ;
        RECT 57.200 31.800 58.000 40.400 ;
        RECT 60.400 33.200 61.400 40.400 ;
        RECT 66.600 39.800 67.400 40.400 ;
        RECT 66.600 33.200 67.600 39.800 ;
        RECT 71.600 32.000 72.400 40.400 ;
        RECT 77.200 35.800 78.000 40.400 ;
        RECT 80.400 35.800 81.200 40.400 ;
        RECT 86.000 31.800 86.800 40.400 ;
        RECT 91.000 39.800 91.800 40.400 ;
        RECT 90.800 33.200 91.800 39.800 ;
        RECT 97.000 33.200 98.000 40.400 ;
        RECT 101.000 35.800 101.800 40.400 ;
        RECT 105.200 31.800 106.000 40.400 ;
        RECT 108.400 32.000 109.200 40.400 ;
        RECT 114.000 35.800 114.800 40.400 ;
        RECT 117.200 35.800 118.000 40.400 ;
        RECT 122.800 31.800 123.600 40.400 ;
        RECT 127.600 33.200 128.600 40.400 ;
        RECT 133.800 39.800 134.600 40.400 ;
        RECT 133.800 33.200 134.800 39.800 ;
        RECT 143.600 33.200 144.600 40.400 ;
        RECT 149.800 39.800 150.600 40.400 ;
        RECT 149.800 33.200 150.800 39.800 ;
        RECT 153.200 35.800 154.000 40.400 ;
        RECT 156.400 35.800 157.200 40.400 ;
        RECT 158.000 35.800 158.800 40.400 ;
        RECT 161.200 35.800 162.000 40.400 ;
        RECT 164.400 35.800 165.200 40.400 ;
        RECT 166.000 31.800 166.800 40.400 ;
        RECT 172.400 31.800 173.200 40.400 ;
        RECT 174.000 31.800 174.800 40.400 ;
        RECT 178.200 35.800 179.000 40.400 ;
        RECT 181.000 35.800 181.800 40.400 ;
        RECT 185.200 31.800 186.000 40.400 ;
        RECT 188.400 33.200 189.400 40.400 ;
        RECT 194.600 39.800 195.400 40.400 ;
        RECT 194.600 33.200 195.600 39.800 ;
        RECT 199.600 33.000 200.400 40.400 ;
        RECT 204.400 35.800 205.200 40.400 ;
        RECT 207.600 32.200 208.400 40.400 ;
        RECT 210.800 35.800 211.600 40.400 ;
        RECT 214.000 35.800 214.800 40.400 ;
        RECT 215.600 35.800 216.400 40.400 ;
        RECT 218.800 35.800 219.600 40.400 ;
        RECT 222.200 39.800 223.000 40.400 ;
        RECT 222.000 33.200 223.000 39.800 ;
        RECT 228.200 33.200 229.200 40.400 ;
        RECT 231.600 35.800 232.400 40.400 ;
        RECT 234.800 35.800 235.600 40.400 ;
        RECT 236.400 31.800 237.200 40.400 ;
        RECT 246.000 33.000 246.800 40.400 ;
        RECT 250.800 33.000 251.600 40.400 ;
        RECT 257.200 35.800 258.000 40.400 ;
        RECT 260.400 35.800 261.200 40.400 ;
        RECT 262.000 35.800 262.800 40.400 ;
        RECT 265.200 35.800 266.000 40.400 ;
        RECT 266.800 31.800 267.600 40.400 ;
        RECT 271.000 35.800 271.800 40.400 ;
        RECT 273.800 35.800 274.600 40.400 ;
        RECT 278.000 31.800 278.800 40.400 ;
        RECT 279.600 31.800 280.400 40.400 ;
        RECT 283.800 35.800 284.600 40.400 ;
        RECT 286.000 31.800 286.800 40.400 ;
        RECT 290.200 35.800 291.000 40.400 ;
        RECT 297.800 35.800 298.600 40.400 ;
        RECT 302.000 31.800 302.800 40.400 ;
        RECT 303.600 31.800 304.400 40.400 ;
        RECT 308.400 31.800 309.200 40.400 ;
        RECT 312.600 35.800 313.400 40.400 ;
        RECT 315.400 35.800 316.200 40.400 ;
        RECT 319.600 31.800 320.400 40.400 ;
        RECT 322.800 35.800 323.600 40.400 ;
        RECT 324.400 35.800 325.200 40.400 ;
        RECT 327.600 31.800 328.400 40.400 ;
        RECT 333.000 35.800 333.800 40.400 ;
        RECT 337.200 31.800 338.000 40.400 ;
        RECT 342.000 31.800 342.800 40.400 ;
        RECT 346.800 33.000 347.600 40.400 ;
        RECT 350.000 35.800 350.800 40.400 ;
        RECT 353.200 35.800 354.000 40.400 ;
        RECT 354.800 31.800 355.600 40.400 ;
        RECT 359.000 35.800 359.800 40.400 ;
        RECT 361.200 35.800 362.000 40.400 ;
        RECT 366.000 33.200 367.000 40.400 ;
        RECT 372.200 39.800 373.000 40.400 ;
        RECT 372.200 33.200 373.200 39.800 ;
        RECT 377.200 32.000 378.000 40.400 ;
        RECT 382.800 35.800 383.600 40.400 ;
        RECT 386.000 35.800 386.800 40.400 ;
        RECT 391.600 31.800 392.400 40.400 ;
        RECT 396.400 33.000 397.200 40.400 ;
        RECT 399.600 31.800 400.400 40.400 ;
        RECT 403.000 39.800 403.800 40.400 ;
        RECT 402.800 33.200 403.800 39.800 ;
        RECT 409.000 33.200 410.000 40.400 ;
        RECT 412.400 35.800 413.200 40.400 ;
        RECT 415.600 35.800 416.400 40.400 ;
        RECT 417.200 31.800 418.000 40.400 ;
        RECT 421.400 35.800 422.200 40.400 ;
        RECT 423.600 35.800 424.400 40.400 ;
        RECT 426.800 35.800 427.600 40.400 ;
        RECT 428.400 35.800 429.200 40.400 ;
        RECT 431.600 35.800 432.400 40.400 ;
        RECT 433.200 31.800 434.000 40.400 ;
        RECT 438.000 31.800 438.800 40.400 ;
        RECT 442.200 35.800 443.000 40.400 ;
        RECT 449.200 35.800 450.000 40.400 ;
        RECT 452.400 35.800 453.200 40.400 ;
        RECT 454.000 35.800 454.800 40.400 ;
        RECT 457.200 35.800 458.000 40.400 ;
        RECT 459.400 35.800 460.200 40.400 ;
        RECT 463.600 31.800 464.400 40.400 ;
        RECT 465.200 35.800 466.000 40.400 ;
        RECT 468.400 35.800 469.200 40.400 ;
        RECT 474.800 33.000 475.600 40.400 ;
        RECT 482.800 33.000 483.600 40.400 ;
        RECT 486.000 31.800 486.800 40.400 ;
        RECT 490.200 35.800 491.000 40.400 ;
        RECT 493.000 35.800 493.800 40.400 ;
        RECT 497.200 31.800 498.000 40.400 ;
        RECT 499.400 35.800 500.200 40.400 ;
        RECT 503.600 31.800 504.400 40.400 ;
        RECT 506.800 33.000 507.600 40.400 ;
        RECT 514.800 35.800 515.600 40.400 ;
        RECT 518.000 33.000 518.800 40.400 ;
        RECT 524.400 31.800 525.200 40.400 ;
        RECT 530.800 33.200 531.800 40.400 ;
        RECT 537.000 39.800 537.800 40.400 ;
        RECT 537.000 33.200 538.000 39.800 ;
        RECT 543.600 31.800 544.400 40.400 ;
        RECT 548.400 33.000 549.200 40.400 ;
        RECT 551.600 35.800 552.400 40.400 ;
        RECT 554.800 35.800 555.600 40.400 ;
        RECT 558.000 35.800 558.800 40.400 ;
        RECT 560.200 35.800 561.000 40.400 ;
        RECT 564.400 31.800 565.200 40.400 ;
        RECT 567.600 33.200 568.600 40.400 ;
        RECT 573.800 39.800 574.600 40.400 ;
        RECT 573.800 33.200 574.800 39.800 ;
        RECT 577.200 31.800 578.000 40.400 ;
        RECT 581.400 35.800 582.200 40.400 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 6.000 1.600 6.800 5.800 ;
        RECT 9.200 1.600 10.000 6.200 ;
        RECT 11.400 1.600 12.200 6.200 ;
        RECT 15.600 1.600 16.400 10.200 ;
        RECT 18.800 1.600 19.800 8.800 ;
        RECT 25.000 2.200 26.000 8.800 ;
        RECT 25.000 1.600 25.800 2.200 ;
        RECT 30.000 1.600 31.000 8.800 ;
        RECT 36.200 2.200 37.200 8.800 ;
        RECT 36.200 1.600 37.000 2.200 ;
        RECT 41.200 1.600 42.000 10.000 ;
        RECT 46.800 1.600 47.600 6.200 ;
        RECT 50.000 1.600 50.800 6.200 ;
        RECT 55.600 1.600 56.400 10.200 ;
        RECT 60.400 1.600 61.200 10.000 ;
        RECT 66.000 1.600 66.800 6.200 ;
        RECT 69.200 1.600 70.000 6.200 ;
        RECT 74.800 1.600 75.600 10.200 ;
        RECT 79.600 1.600 80.400 10.000 ;
        RECT 85.200 1.600 86.000 6.200 ;
        RECT 88.400 1.600 89.200 6.200 ;
        RECT 94.000 1.600 94.800 10.200 ;
        RECT 98.800 1.600 99.600 10.000 ;
        RECT 104.400 1.600 105.200 6.200 ;
        RECT 107.600 1.600 108.400 6.200 ;
        RECT 113.200 1.600 114.000 10.200 ;
        RECT 118.000 1.600 118.800 10.000 ;
        RECT 123.600 1.600 124.400 6.200 ;
        RECT 126.800 1.600 127.600 6.200 ;
        RECT 132.400 1.600 133.200 10.200 ;
        RECT 142.000 2.200 143.000 8.800 ;
        RECT 142.200 1.600 143.000 2.200 ;
        RECT 148.200 1.600 149.200 8.800 ;
        RECT 151.600 1.600 152.400 10.200 ;
        RECT 155.800 1.600 156.600 6.200 ;
        RECT 159.600 1.600 160.400 6.200 ;
        RECT 161.200 1.600 162.000 6.200 ;
        RECT 167.600 1.600 168.400 10.200 ;
        RECT 172.400 1.600 173.200 9.000 ;
        RECT 177.200 1.600 178.000 9.000 ;
        RECT 180.400 1.600 181.200 10.200 ;
        RECT 183.600 2.200 184.600 8.800 ;
        RECT 183.800 1.600 184.600 2.200 ;
        RECT 189.800 1.600 190.800 8.800 ;
        RECT 193.200 1.600 194.000 10.200 ;
        RECT 197.400 1.600 198.200 6.200 ;
        RECT 199.600 1.600 200.400 10.200 ;
        RECT 203.800 1.600 204.600 6.200 ;
        RECT 206.600 1.600 207.400 6.200 ;
        RECT 210.800 1.600 211.600 10.200 ;
        RECT 212.400 1.600 213.200 10.200 ;
        RECT 218.800 1.600 219.600 6.200 ;
        RECT 220.400 1.600 221.200 6.200 ;
        RECT 223.600 1.600 224.400 6.200 ;
        RECT 225.200 1.600 226.000 6.200 ;
        RECT 228.400 1.600 229.200 6.200 ;
        RECT 231.600 1.600 232.400 6.200 ;
        RECT 234.800 2.200 235.800 8.800 ;
        RECT 235.000 1.600 235.800 2.200 ;
        RECT 241.000 1.600 242.000 8.800 ;
        RECT 244.400 1.600 245.200 6.200 ;
        RECT 247.600 1.600 248.400 6.200 ;
        RECT 249.200 1.600 250.000 6.200 ;
        RECT 252.400 1.600 253.200 6.200 ;
        RECT 254.000 1.600 254.800 10.200 ;
        RECT 258.200 1.600 259.000 6.200 ;
        RECT 260.400 1.600 261.200 6.200 ;
        RECT 263.600 1.600 264.400 6.200 ;
        RECT 266.800 1.600 267.800 8.800 ;
        RECT 273.000 2.200 274.000 8.800 ;
        RECT 273.000 1.600 273.800 2.200 ;
        RECT 276.400 1.600 277.200 10.200 ;
        RECT 280.600 1.600 281.400 6.200 ;
        RECT 284.400 1.600 285.400 8.800 ;
        RECT 290.600 2.200 291.600 8.800 ;
        RECT 290.600 1.600 291.400 2.200 ;
        RECT 298.800 1.600 299.600 6.200 ;
        RECT 302.000 1.600 302.800 6.200 ;
        RECT 304.200 1.600 305.000 6.200 ;
        RECT 308.400 1.600 309.200 10.200 ;
        RECT 310.000 1.600 310.800 6.200 ;
        RECT 313.200 1.600 314.000 6.200 ;
        RECT 316.400 1.600 317.200 6.200 ;
        RECT 319.200 1.600 320.000 10.200 ;
        RECT 324.400 1.600 325.200 9.800 ;
        RECT 329.200 2.200 330.200 8.800 ;
        RECT 329.400 1.600 330.200 2.200 ;
        RECT 335.400 1.600 336.400 8.800 ;
        RECT 340.400 1.600 341.200 10.000 ;
        RECT 346.000 1.600 346.800 6.200 ;
        RECT 349.200 1.600 350.000 6.200 ;
        RECT 354.800 1.600 355.600 10.200 ;
        RECT 359.600 1.600 360.400 10.000 ;
        RECT 365.200 1.600 366.000 6.200 ;
        RECT 368.400 1.600 369.200 6.200 ;
        RECT 374.000 1.600 374.800 10.200 ;
        RECT 378.800 1.600 379.600 10.000 ;
        RECT 384.400 1.600 385.200 6.200 ;
        RECT 387.600 1.600 388.400 6.200 ;
        RECT 393.200 1.600 394.000 10.200 ;
        RECT 398.000 1.600 398.800 9.000 ;
        RECT 401.200 1.600 402.000 10.200 ;
        RECT 404.400 1.600 405.400 8.800 ;
        RECT 410.600 2.200 411.600 8.800 ;
        RECT 410.600 1.600 411.400 2.200 ;
        RECT 414.000 1.600 414.800 6.200 ;
        RECT 417.200 1.600 418.000 10.200 ;
        RECT 421.400 1.600 422.200 6.200 ;
        RECT 424.200 1.600 425.000 6.200 ;
        RECT 428.400 1.600 429.200 10.200 ;
        RECT 430.000 1.600 430.800 6.200 ;
        RECT 433.200 1.600 434.000 6.200 ;
        RECT 436.400 1.600 437.200 9.000 ;
        RECT 439.600 1.600 440.400 10.200 ;
        RECT 441.200 1.600 442.000 6.200 ;
        RECT 449.200 1.600 450.000 6.200 ;
        RECT 452.400 1.600 453.200 6.200 ;
        RECT 454.000 1.600 454.800 6.200 ;
        RECT 457.200 1.600 458.000 6.200 ;
        RECT 462.000 1.600 462.800 10.200 ;
        RECT 463.600 1.600 464.400 10.200 ;
        RECT 467.800 1.600 468.600 6.200 ;
        RECT 471.600 2.200 472.600 8.800 ;
        RECT 471.800 1.600 472.600 2.200 ;
        RECT 477.800 1.600 478.800 8.800 ;
        RECT 481.200 1.600 482.000 10.200 ;
        RECT 485.400 1.600 486.200 6.200 ;
        RECT 488.200 1.600 489.000 6.200 ;
        RECT 492.400 1.600 493.200 10.200 ;
        RECT 494.000 1.600 494.800 10.200 ;
        RECT 498.200 1.600 499.000 6.200 ;
        RECT 503.000 1.600 503.800 10.200 ;
        RECT 506.800 1.600 507.600 10.200 ;
        RECT 511.600 1.600 512.400 6.200 ;
        RECT 514.800 1.600 515.600 10.200 ;
        RECT 518.000 1.600 518.800 9.000 ;
        RECT 521.200 1.600 522.000 6.200 ;
        RECT 525.000 1.600 525.800 6.200 ;
        RECT 529.200 1.600 530.000 10.200 ;
        RECT 534.000 1.600 534.800 10.200 ;
        RECT 535.600 1.600 536.400 10.200 ;
        RECT 540.400 1.600 541.200 10.200 ;
        RECT 546.800 1.600 547.600 9.000 ;
        RECT 553.200 1.600 554.000 10.200 ;
        RECT 554.800 1.600 555.600 6.200 ;
        RECT 558.000 1.600 558.800 9.800 ;
        RECT 562.800 1.600 563.800 8.800 ;
        RECT 569.000 2.200 570.000 8.800 ;
        RECT 569.000 1.600 569.800 2.200 ;
        RECT 572.400 1.600 573.200 10.200 ;
        RECT 576.600 1.600 577.400 6.200 ;
        RECT 580.400 1.600 581.200 9.000 ;
        RECT 0.400 0.400 586.800 1.600 ;
      LAYER via1 ;
        RECT 290.800 411.800 291.600 412.600 ;
        RECT 454.000 407.600 454.800 408.400 ;
        RECT 519.600 403.600 520.400 404.400 ;
        RECT 578.800 403.600 579.600 404.400 ;
        RECT 135.800 400.600 136.600 401.400 ;
        RECT 137.200 400.600 138.000 401.400 ;
        RECT 138.600 400.600 139.400 401.400 ;
        RECT 444.600 400.600 445.400 401.400 ;
        RECT 446.000 400.600 446.800 401.400 ;
        RECT 447.400 400.600 448.200 401.400 ;
        RECT 290.800 399.600 291.600 400.400 ;
        RECT 508.400 399.600 509.200 400.400 ;
        RECT 518.000 391.200 518.800 392.000 ;
        RECT 553.200 391.200 554.000 392.000 ;
        RECT 502.000 363.600 502.800 364.400 ;
        RECT 554.800 363.600 555.600 364.400 ;
        RECT 135.800 360.600 136.600 361.400 ;
        RECT 137.200 360.600 138.000 361.400 ;
        RECT 138.600 360.600 139.400 361.400 ;
        RECT 444.600 360.600 445.400 361.400 ;
        RECT 446.000 360.600 446.800 361.400 ;
        RECT 447.400 360.600 448.200 361.400 ;
        RECT 553.200 357.600 554.000 358.400 ;
        RECT 521.200 351.200 522.000 352.000 ;
        RECT 553.200 351.600 554.000 352.400 ;
        RECT 550.000 323.600 550.800 324.400 ;
        RECT 135.800 320.600 136.600 321.400 ;
        RECT 137.200 320.600 138.000 321.400 ;
        RECT 138.600 320.600 139.400 321.400 ;
        RECT 444.600 320.600 445.400 321.400 ;
        RECT 446.000 320.600 446.800 321.400 ;
        RECT 447.400 320.600 448.200 321.400 ;
        RECT 135.800 280.600 136.600 281.400 ;
        RECT 137.200 280.600 138.000 281.400 ;
        RECT 138.600 280.600 139.400 281.400 ;
        RECT 444.600 280.600 445.400 281.400 ;
        RECT 446.000 280.600 446.800 281.400 ;
        RECT 447.400 280.600 448.200 281.400 ;
        RECT 135.800 240.600 136.600 241.400 ;
        RECT 137.200 240.600 138.000 241.400 ;
        RECT 138.600 240.600 139.400 241.400 ;
        RECT 444.600 240.600 445.400 241.400 ;
        RECT 446.000 240.600 446.800 241.400 ;
        RECT 447.400 240.600 448.200 241.400 ;
        RECT 135.800 200.600 136.600 201.400 ;
        RECT 137.200 200.600 138.000 201.400 ;
        RECT 138.600 200.600 139.400 201.400 ;
        RECT 444.600 200.600 445.400 201.400 ;
        RECT 446.000 200.600 446.800 201.400 ;
        RECT 447.400 200.600 448.200 201.400 ;
        RECT 135.800 160.600 136.600 161.400 ;
        RECT 137.200 160.600 138.000 161.400 ;
        RECT 138.600 160.600 139.400 161.400 ;
        RECT 444.600 160.600 445.400 161.400 ;
        RECT 446.000 160.600 446.800 161.400 ;
        RECT 447.400 160.600 448.200 161.400 ;
        RECT 553.200 127.600 554.000 128.400 ;
        RECT 580.400 127.600 581.200 128.400 ;
        RECT 135.800 120.600 136.600 121.400 ;
        RECT 137.200 120.600 138.000 121.400 ;
        RECT 138.600 120.600 139.400 121.400 ;
        RECT 444.600 120.600 445.400 121.400 ;
        RECT 446.000 120.600 446.800 121.400 ;
        RECT 447.400 120.600 448.200 121.400 ;
        RECT 135.800 80.600 136.600 81.400 ;
        RECT 137.200 80.600 138.000 81.400 ;
        RECT 138.600 80.600 139.400 81.400 ;
        RECT 444.600 80.600 445.400 81.400 ;
        RECT 446.000 80.600 446.800 81.400 ;
        RECT 447.400 80.600 448.200 81.400 ;
        RECT 135.800 40.600 136.600 41.400 ;
        RECT 137.200 40.600 138.000 41.400 ;
        RECT 138.600 40.600 139.400 41.400 ;
        RECT 444.600 40.600 445.400 41.400 ;
        RECT 446.000 40.600 446.800 41.400 ;
        RECT 447.400 40.600 448.200 41.400 ;
        RECT 135.800 0.600 136.600 1.400 ;
        RECT 137.200 0.600 138.000 1.400 ;
        RECT 138.600 0.600 139.400 1.400 ;
        RECT 444.600 0.600 445.400 1.400 ;
        RECT 446.000 0.600 446.800 1.400 ;
        RECT 447.400 0.600 448.200 1.400 ;
      LAYER metal2 ;
        RECT 290.800 411.800 291.600 412.600 ;
        RECT 135.200 400.600 140.000 401.400 ;
        RECT 290.900 400.400 291.500 411.800 ;
        RECT 455.600 411.600 456.400 412.400 ;
        RECT 508.400 411.600 509.200 412.400 ;
        RECT 454.000 408.300 454.800 408.400 ;
        RECT 455.700 408.300 456.300 411.600 ;
        RECT 454.000 407.700 456.300 408.300 ;
        RECT 454.000 407.600 454.800 407.700 ;
        RECT 444.000 400.600 448.800 401.400 ;
        RECT 508.500 400.400 509.100 411.600 ;
        RECT 519.600 410.000 520.400 410.800 ;
        RECT 519.700 404.400 520.300 410.000 ;
        RECT 578.800 409.600 579.600 410.400 ;
        RECT 578.900 404.400 579.500 409.600 ;
        RECT 519.600 403.600 520.400 404.400 ;
        RECT 578.800 403.600 579.600 404.400 ;
        RECT 290.800 399.600 291.600 400.400 ;
        RECT 508.400 399.600 509.200 400.400 ;
        RECT 511.600 395.800 512.400 396.600 ;
        RECT 518.000 395.800 518.800 396.600 ;
        RECT 553.200 395.800 554.000 396.600 ;
        RECT 511.700 374.400 512.300 395.800 ;
        RECT 518.100 392.000 518.700 395.800 ;
        RECT 553.300 392.000 553.900 395.800 ;
        RECT 518.000 391.200 518.800 392.000 ;
        RECT 553.200 391.200 554.000 392.000 ;
        RECT 511.600 373.600 512.400 374.400 ;
        RECT 502.000 369.600 502.800 370.400 ;
        RECT 554.800 370.000 555.600 370.800 ;
        RECT 502.100 364.400 502.700 369.600 ;
        RECT 554.900 364.400 555.500 370.000 ;
        RECT 502.000 363.600 502.800 364.400 ;
        RECT 554.800 363.600 555.600 364.400 ;
        RECT 135.200 360.600 140.000 361.400 ;
        RECT 444.000 360.600 448.800 361.400 ;
        RECT 553.200 357.600 554.000 358.400 ;
        RECT 514.800 355.800 515.600 356.600 ;
        RECT 521.200 355.800 522.000 356.600 ;
        RECT 514.900 332.400 515.500 355.800 ;
        RECT 521.300 352.000 521.900 355.800 ;
        RECT 553.300 352.400 553.900 357.600 ;
        RECT 521.200 351.200 522.000 352.000 ;
        RECT 553.200 351.600 554.000 352.400 ;
        RECT 514.800 331.600 515.600 332.400 ;
        RECT 550.000 329.600 550.800 330.400 ;
        RECT 550.100 324.400 550.700 329.600 ;
        RECT 550.000 323.600 550.800 324.400 ;
        RECT 135.200 320.600 140.000 321.400 ;
        RECT 444.000 320.600 448.800 321.400 ;
        RECT 135.200 280.600 140.000 281.400 ;
        RECT 444.000 280.600 448.800 281.400 ;
        RECT 135.200 240.600 140.000 241.400 ;
        RECT 444.000 240.600 448.800 241.400 ;
        RECT 135.200 200.600 140.000 201.400 ;
        RECT 444.000 200.600 448.800 201.400 ;
        RECT 135.200 160.600 140.000 161.400 ;
        RECT 444.000 160.600 448.800 161.400 ;
        RECT 554.800 131.600 555.600 132.400 ;
        RECT 578.800 131.600 579.600 132.400 ;
        RECT 553.200 128.300 554.000 128.400 ;
        RECT 554.900 128.300 555.500 131.600 ;
        RECT 553.200 127.700 555.500 128.300 ;
        RECT 578.900 128.300 579.500 131.600 ;
        RECT 580.400 128.300 581.200 128.400 ;
        RECT 578.900 127.700 581.200 128.300 ;
        RECT 553.200 127.600 554.000 127.700 ;
        RECT 580.400 127.600 581.200 127.700 ;
        RECT 135.200 120.600 140.000 121.400 ;
        RECT 444.000 120.600 448.800 121.400 ;
        RECT 135.200 80.600 140.000 81.400 ;
        RECT 444.000 80.600 448.800 81.400 ;
        RECT 135.200 40.600 140.000 41.400 ;
        RECT 444.000 40.600 448.800 41.400 ;
        RECT 135.200 0.600 140.000 1.400 ;
        RECT 444.000 0.600 448.800 1.400 ;
      LAYER via2 ;
        RECT 135.800 400.600 136.600 401.400 ;
        RECT 137.200 400.600 138.000 401.400 ;
        RECT 138.600 400.600 139.400 401.400 ;
        RECT 444.600 400.600 445.400 401.400 ;
        RECT 446.000 400.600 446.800 401.400 ;
        RECT 447.400 400.600 448.200 401.400 ;
        RECT 135.800 360.600 136.600 361.400 ;
        RECT 137.200 360.600 138.000 361.400 ;
        RECT 138.600 360.600 139.400 361.400 ;
        RECT 444.600 360.600 445.400 361.400 ;
        RECT 446.000 360.600 446.800 361.400 ;
        RECT 447.400 360.600 448.200 361.400 ;
        RECT 135.800 320.600 136.600 321.400 ;
        RECT 137.200 320.600 138.000 321.400 ;
        RECT 138.600 320.600 139.400 321.400 ;
        RECT 444.600 320.600 445.400 321.400 ;
        RECT 446.000 320.600 446.800 321.400 ;
        RECT 447.400 320.600 448.200 321.400 ;
        RECT 135.800 280.600 136.600 281.400 ;
        RECT 137.200 280.600 138.000 281.400 ;
        RECT 138.600 280.600 139.400 281.400 ;
        RECT 444.600 280.600 445.400 281.400 ;
        RECT 446.000 280.600 446.800 281.400 ;
        RECT 447.400 280.600 448.200 281.400 ;
        RECT 135.800 240.600 136.600 241.400 ;
        RECT 137.200 240.600 138.000 241.400 ;
        RECT 138.600 240.600 139.400 241.400 ;
        RECT 444.600 240.600 445.400 241.400 ;
        RECT 446.000 240.600 446.800 241.400 ;
        RECT 447.400 240.600 448.200 241.400 ;
        RECT 135.800 200.600 136.600 201.400 ;
        RECT 137.200 200.600 138.000 201.400 ;
        RECT 138.600 200.600 139.400 201.400 ;
        RECT 444.600 200.600 445.400 201.400 ;
        RECT 446.000 200.600 446.800 201.400 ;
        RECT 447.400 200.600 448.200 201.400 ;
        RECT 135.800 160.600 136.600 161.400 ;
        RECT 137.200 160.600 138.000 161.400 ;
        RECT 138.600 160.600 139.400 161.400 ;
        RECT 444.600 160.600 445.400 161.400 ;
        RECT 446.000 160.600 446.800 161.400 ;
        RECT 447.400 160.600 448.200 161.400 ;
        RECT 135.800 120.600 136.600 121.400 ;
        RECT 137.200 120.600 138.000 121.400 ;
        RECT 138.600 120.600 139.400 121.400 ;
        RECT 444.600 120.600 445.400 121.400 ;
        RECT 446.000 120.600 446.800 121.400 ;
        RECT 447.400 120.600 448.200 121.400 ;
        RECT 135.800 80.600 136.600 81.400 ;
        RECT 137.200 80.600 138.000 81.400 ;
        RECT 138.600 80.600 139.400 81.400 ;
        RECT 444.600 80.600 445.400 81.400 ;
        RECT 446.000 80.600 446.800 81.400 ;
        RECT 447.400 80.600 448.200 81.400 ;
        RECT 135.800 40.600 136.600 41.400 ;
        RECT 137.200 40.600 138.000 41.400 ;
        RECT 138.600 40.600 139.400 41.400 ;
        RECT 444.600 40.600 445.400 41.400 ;
        RECT 446.000 40.600 446.800 41.400 ;
        RECT 447.400 40.600 448.200 41.400 ;
        RECT 135.800 0.600 136.600 1.400 ;
        RECT 137.200 0.600 138.000 1.400 ;
        RECT 138.600 0.600 139.400 1.400 ;
        RECT 444.600 0.600 445.400 1.400 ;
        RECT 446.000 0.600 446.800 1.400 ;
        RECT 447.400 0.600 448.200 1.400 ;
      LAYER metal3 ;
        RECT 135.200 400.400 140.000 401.600 ;
        RECT 444.000 400.400 448.800 401.600 ;
        RECT 135.200 360.400 140.000 361.600 ;
        RECT 444.000 360.400 448.800 361.600 ;
        RECT 135.200 320.400 140.000 321.600 ;
        RECT 444.000 320.400 448.800 321.600 ;
        RECT 135.200 280.400 140.000 281.600 ;
        RECT 444.000 280.400 448.800 281.600 ;
        RECT 135.200 240.400 140.000 241.600 ;
        RECT 444.000 240.400 448.800 241.600 ;
        RECT 135.200 200.400 140.000 201.600 ;
        RECT 444.000 200.400 448.800 201.600 ;
        RECT 135.200 160.400 140.000 161.600 ;
        RECT 444.000 160.400 448.800 161.600 ;
        RECT 135.200 120.400 140.000 121.600 ;
        RECT 444.000 120.400 448.800 121.600 ;
        RECT 135.200 80.400 140.000 81.600 ;
        RECT 444.000 80.400 448.800 81.600 ;
        RECT 135.200 40.400 140.000 41.600 ;
        RECT 444.000 40.400 448.800 41.600 ;
        RECT 135.200 0.400 140.000 1.600 ;
        RECT 444.000 0.400 448.800 1.600 ;
      LAYER via3 ;
        RECT 135.600 400.600 136.400 401.400 ;
        RECT 137.200 400.600 138.000 401.400 ;
        RECT 138.800 400.600 139.600 401.400 ;
        RECT 444.400 400.600 445.200 401.400 ;
        RECT 446.000 400.600 446.800 401.400 ;
        RECT 447.600 400.600 448.400 401.400 ;
        RECT 135.600 360.600 136.400 361.400 ;
        RECT 137.200 360.600 138.000 361.400 ;
        RECT 138.800 360.600 139.600 361.400 ;
        RECT 444.400 360.600 445.200 361.400 ;
        RECT 446.000 360.600 446.800 361.400 ;
        RECT 447.600 360.600 448.400 361.400 ;
        RECT 135.600 320.600 136.400 321.400 ;
        RECT 137.200 320.600 138.000 321.400 ;
        RECT 138.800 320.600 139.600 321.400 ;
        RECT 444.400 320.600 445.200 321.400 ;
        RECT 446.000 320.600 446.800 321.400 ;
        RECT 447.600 320.600 448.400 321.400 ;
        RECT 135.600 280.600 136.400 281.400 ;
        RECT 137.200 280.600 138.000 281.400 ;
        RECT 138.800 280.600 139.600 281.400 ;
        RECT 444.400 280.600 445.200 281.400 ;
        RECT 446.000 280.600 446.800 281.400 ;
        RECT 447.600 280.600 448.400 281.400 ;
        RECT 135.600 240.600 136.400 241.400 ;
        RECT 137.200 240.600 138.000 241.400 ;
        RECT 138.800 240.600 139.600 241.400 ;
        RECT 444.400 240.600 445.200 241.400 ;
        RECT 446.000 240.600 446.800 241.400 ;
        RECT 447.600 240.600 448.400 241.400 ;
        RECT 135.600 200.600 136.400 201.400 ;
        RECT 137.200 200.600 138.000 201.400 ;
        RECT 138.800 200.600 139.600 201.400 ;
        RECT 444.400 200.600 445.200 201.400 ;
        RECT 446.000 200.600 446.800 201.400 ;
        RECT 447.600 200.600 448.400 201.400 ;
        RECT 135.600 160.600 136.400 161.400 ;
        RECT 137.200 160.600 138.000 161.400 ;
        RECT 138.800 160.600 139.600 161.400 ;
        RECT 444.400 160.600 445.200 161.400 ;
        RECT 446.000 160.600 446.800 161.400 ;
        RECT 447.600 160.600 448.400 161.400 ;
        RECT 135.600 120.600 136.400 121.400 ;
        RECT 137.200 120.600 138.000 121.400 ;
        RECT 138.800 120.600 139.600 121.400 ;
        RECT 444.400 120.600 445.200 121.400 ;
        RECT 446.000 120.600 446.800 121.400 ;
        RECT 447.600 120.600 448.400 121.400 ;
        RECT 135.600 80.600 136.400 81.400 ;
        RECT 137.200 80.600 138.000 81.400 ;
        RECT 138.800 80.600 139.600 81.400 ;
        RECT 444.400 80.600 445.200 81.400 ;
        RECT 446.000 80.600 446.800 81.400 ;
        RECT 447.600 80.600 448.400 81.400 ;
        RECT 135.600 40.600 136.400 41.400 ;
        RECT 137.200 40.600 138.000 41.400 ;
        RECT 138.800 40.600 139.600 41.400 ;
        RECT 444.400 40.600 445.200 41.400 ;
        RECT 446.000 40.600 446.800 41.400 ;
        RECT 447.600 40.600 448.400 41.400 ;
        RECT 135.600 0.600 136.400 1.400 ;
        RECT 137.200 0.600 138.000 1.400 ;
        RECT 138.800 0.600 139.600 1.400 ;
        RECT 444.400 0.600 445.200 1.400 ;
        RECT 446.000 0.600 446.800 1.400 ;
        RECT 447.600 0.600 448.400 1.400 ;
      LAYER metal4 ;
        RECT 135.200 0.000 140.000 424.000 ;
        RECT 444.000 0.000 448.800 424.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.400 420.400 586.800 421.600 ;
        RECT 4.400 416.600 5.200 420.400 ;
        RECT 9.200 417.800 10.000 420.400 ;
        RECT 10.800 417.800 11.600 420.400 ;
        RECT 14.000 416.200 14.800 420.400 ;
        RECT 17.200 415.800 18.000 420.400 ;
        RECT 25.200 416.600 26.000 420.400 ;
        RECT 28.400 417.800 29.200 420.400 ;
        RECT 31.600 417.800 32.400 420.400 ;
        RECT 34.800 416.600 35.600 420.400 ;
        RECT 41.800 416.000 42.600 420.400 ;
        RECT 47.600 416.000 48.400 420.400 ;
        RECT 53.200 417.800 54.000 420.400 ;
        RECT 56.400 417.800 57.400 420.400 ;
        RECT 62.000 415.800 62.800 420.400 ;
        RECT 66.800 416.000 67.600 420.400 ;
        RECT 72.400 417.800 73.200 420.400 ;
        RECT 75.600 417.800 76.600 420.400 ;
        RECT 81.200 415.800 82.000 420.400 ;
        RECT 84.400 415.800 85.200 420.400 ;
        RECT 87.600 415.800 88.400 420.400 ;
        RECT 90.800 415.800 91.600 420.400 ;
        RECT 94.000 415.800 94.800 420.400 ;
        RECT 97.200 415.800 98.000 420.400 ;
        RECT 98.800 415.800 99.600 420.400 ;
        RECT 105.200 416.000 106.000 420.400 ;
        RECT 110.800 417.800 111.600 420.400 ;
        RECT 114.000 417.800 115.000 420.400 ;
        RECT 119.600 415.800 120.400 420.400 ;
        RECT 124.600 419.800 125.400 420.400 ;
        RECT 124.400 416.400 125.400 419.800 ;
        RECT 130.600 416.400 131.600 420.400 ;
        RECT 142.000 416.600 142.800 420.400 ;
        RECT 148.400 415.800 149.200 420.400 ;
        RECT 151.800 419.800 152.600 420.400 ;
        RECT 151.600 416.400 152.600 419.800 ;
        RECT 157.800 416.400 158.800 420.400 ;
        RECT 161.200 415.800 162.000 420.400 ;
        RECT 169.200 415.800 170.000 420.400 ;
        RECT 172.400 416.600 173.200 420.400 ;
        RECT 180.400 416.600 181.200 420.400 ;
        RECT 183.600 417.800 184.400 420.400 ;
        RECT 186.800 417.800 187.600 420.400 ;
        RECT 188.400 417.800 189.200 420.400 ;
        RECT 192.600 415.800 193.400 420.400 ;
        RECT 194.800 417.800 195.600 420.400 ;
        RECT 198.000 417.800 198.800 420.400 ;
        RECT 199.600 417.800 200.400 420.400 ;
        RECT 202.800 417.800 203.600 420.400 ;
        RECT 206.000 415.800 206.800 420.400 ;
        RECT 210.800 417.800 211.600 420.400 ;
        RECT 212.400 417.800 213.200 420.400 ;
        RECT 215.600 417.800 216.400 420.400 ;
        RECT 217.200 415.800 218.000 420.400 ;
        RECT 222.000 416.000 222.800 420.400 ;
        RECT 227.600 417.800 228.400 420.400 ;
        RECT 230.800 417.800 231.800 420.400 ;
        RECT 236.400 415.800 237.200 420.400 ;
        RECT 241.200 417.800 242.000 420.400 ;
        RECT 244.400 416.000 245.200 420.400 ;
        RECT 250.000 417.800 250.800 420.400 ;
        RECT 253.200 417.800 254.200 420.400 ;
        RECT 258.800 415.800 259.600 420.400 ;
        RECT 263.600 415.800 264.400 420.400 ;
        RECT 266.800 415.800 267.600 420.400 ;
        RECT 273.200 416.600 274.000 420.400 ;
        RECT 279.600 416.000 280.400 420.400 ;
        RECT 285.200 417.800 286.000 420.400 ;
        RECT 288.400 417.800 289.400 420.400 ;
        RECT 294.000 415.800 294.800 420.400 ;
        RECT 302.000 415.800 302.800 420.400 ;
        RECT 305.200 415.800 306.000 420.400 ;
        RECT 308.400 415.800 309.200 420.400 ;
        RECT 311.600 415.800 312.400 420.400 ;
        RECT 314.800 415.800 315.600 420.400 ;
        RECT 318.000 416.000 318.800 420.400 ;
        RECT 323.600 417.800 324.400 420.400 ;
        RECT 326.800 417.800 327.800 420.400 ;
        RECT 332.400 415.800 333.200 420.400 ;
        RECT 337.200 415.800 338.000 420.400 ;
        RECT 342.000 415.800 342.800 420.400 ;
        RECT 346.800 415.800 347.600 420.400 ;
        RECT 351.600 415.800 352.400 420.400 ;
        RECT 354.800 417.800 355.600 420.400 ;
        RECT 361.200 415.800 362.000 420.400 ;
        RECT 372.400 417.800 373.200 420.400 ;
        RECT 375.600 417.800 376.400 420.400 ;
        RECT 385.200 415.800 386.000 420.400 ;
        RECT 393.200 415.800 394.000 420.400 ;
        RECT 396.400 416.200 397.200 420.400 ;
        RECT 399.600 417.800 400.400 420.400 ;
        RECT 401.200 417.800 402.000 420.400 ;
        RECT 407.600 415.800 408.400 420.400 ;
        RECT 418.800 417.800 419.600 420.400 ;
        RECT 422.000 417.800 422.800 420.400 ;
        RECT 431.600 415.800 432.400 420.400 ;
        RECT 439.600 415.800 440.400 420.400 ;
        RECT 447.600 416.200 448.400 420.400 ;
        RECT 450.800 417.800 451.600 420.400 ;
        RECT 454.000 415.800 454.800 420.400 ;
        RECT 458.800 415.800 459.600 420.400 ;
        RECT 462.000 417.800 462.800 420.400 ;
        RECT 468.400 415.800 469.200 420.400 ;
        RECT 479.600 417.800 480.400 420.400 ;
        RECT 482.800 417.800 483.600 420.400 ;
        RECT 492.400 415.800 493.200 420.400 ;
        RECT 500.400 415.800 501.200 420.400 ;
        RECT 503.600 416.200 504.400 420.400 ;
        RECT 506.800 417.800 507.600 420.400 ;
        RECT 510.000 415.800 510.800 420.400 ;
        RECT 516.400 415.800 517.200 420.400 ;
        RECT 526.000 417.800 526.800 420.400 ;
        RECT 529.200 417.800 530.000 420.400 ;
        RECT 540.400 415.800 541.200 420.400 ;
        RECT 546.800 417.800 547.600 420.400 ;
        RECT 548.400 417.800 549.200 420.400 ;
        RECT 554.800 415.800 555.600 420.400 ;
        RECT 566.000 417.800 566.800 420.400 ;
        RECT 569.200 417.800 570.000 420.400 ;
        RECT 578.800 415.800 579.600 420.400 ;
        RECT 2.800 381.600 3.600 385.400 ;
        RECT 7.600 381.600 8.400 386.200 ;
        RECT 15.600 381.600 16.400 386.200 ;
        RECT 20.400 381.600 21.200 386.200 ;
        RECT 22.000 381.600 22.800 386.200 ;
        RECT 26.800 381.600 27.600 384.200 ;
        RECT 30.000 381.600 30.800 384.200 ;
        RECT 32.200 381.600 33.000 386.200 ;
        RECT 36.400 381.600 37.200 384.200 ;
        RECT 41.200 381.600 42.000 385.400 ;
        RECT 47.600 381.600 48.400 386.200 ;
        RECT 49.200 381.600 50.000 386.200 ;
        RECT 54.000 381.600 54.800 384.200 ;
        RECT 57.200 381.600 58.000 384.200 ;
        RECT 58.800 381.600 59.600 384.200 ;
        RECT 63.000 381.600 63.800 386.200 ;
        RECT 66.800 381.600 67.800 385.600 ;
        RECT 73.000 382.200 74.000 385.600 ;
        RECT 73.000 381.600 73.800 382.200 ;
        RECT 76.400 381.600 77.200 384.200 ;
        RECT 81.200 381.600 82.000 385.400 ;
        RECT 89.200 381.600 90.000 385.400 ;
        RECT 95.600 381.600 96.400 386.200 ;
        RECT 100.400 381.600 101.200 386.200 ;
        RECT 102.000 381.600 102.800 384.200 ;
        RECT 108.400 381.600 109.200 386.200 ;
        RECT 111.600 381.600 112.400 384.200 ;
        RECT 114.800 381.600 115.600 386.000 ;
        RECT 120.400 381.600 121.200 384.200 ;
        RECT 123.600 381.600 124.600 384.200 ;
        RECT 129.200 381.600 130.000 386.200 ;
        RECT 138.800 382.200 139.800 385.600 ;
        RECT 139.000 381.600 139.800 382.200 ;
        RECT 145.000 381.600 146.000 385.600 ;
        RECT 150.000 382.200 151.000 385.600 ;
        RECT 150.200 381.600 151.000 382.200 ;
        RECT 156.200 381.600 157.200 385.600 ;
        RECT 161.200 381.600 162.000 385.400 ;
        RECT 169.200 381.600 170.000 385.400 ;
        RECT 175.600 381.600 176.400 386.200 ;
        RECT 178.800 381.600 179.600 385.400 ;
        RECT 186.800 381.600 187.600 385.400 ;
        RECT 190.000 381.600 190.800 386.200 ;
        RECT 196.400 381.600 197.200 386.200 ;
        RECT 199.600 381.600 200.400 385.400 ;
        RECT 204.400 381.600 205.200 384.200 ;
        RECT 207.600 381.600 208.400 384.200 ;
        RECT 209.800 381.600 210.600 386.200 ;
        RECT 214.000 381.600 214.800 384.200 ;
        RECT 215.600 381.600 216.400 384.200 ;
        RECT 218.800 381.600 219.600 384.200 ;
        RECT 223.600 381.600 224.400 386.200 ;
        RECT 228.400 381.600 229.200 386.200 ;
        RECT 230.000 381.600 230.800 384.200 ;
        RECT 234.800 381.600 235.600 385.400 ;
        RECT 242.800 381.600 243.600 386.200 ;
        RECT 244.400 381.600 245.200 384.200 ;
        RECT 248.600 381.600 249.400 386.200 ;
        RECT 250.800 381.600 251.600 384.200 ;
        RECT 254.000 381.600 254.800 384.200 ;
        RECT 257.200 382.200 258.200 385.600 ;
        RECT 257.400 381.600 258.200 382.200 ;
        RECT 263.400 381.600 264.400 385.600 ;
        RECT 270.000 381.600 270.800 386.200 ;
        RECT 274.800 381.600 275.600 386.200 ;
        RECT 278.000 381.600 278.800 385.400 ;
        RECT 284.400 382.200 285.400 385.600 ;
        RECT 284.600 381.600 285.400 382.200 ;
        RECT 290.600 381.600 291.600 385.600 ;
        RECT 298.800 381.600 299.600 384.200 ;
        RECT 302.000 381.600 302.800 384.200 ;
        RECT 303.600 381.600 304.400 386.200 ;
        RECT 311.600 381.600 312.400 386.200 ;
        RECT 316.400 381.600 317.200 385.400 ;
        RECT 321.200 381.600 322.000 385.400 ;
        RECT 327.600 381.600 328.400 384.200 ;
        RECT 330.800 381.600 331.600 386.000 ;
        RECT 336.400 381.600 337.200 384.200 ;
        RECT 339.600 381.600 340.600 384.200 ;
        RECT 345.200 381.600 346.000 386.200 ;
        RECT 348.400 381.600 349.200 384.200 ;
        RECT 351.600 381.600 352.400 384.200 ;
        RECT 354.800 381.600 355.600 386.200 ;
        RECT 358.000 381.600 358.800 386.200 ;
        RECT 361.200 381.600 362.000 384.200 ;
        RECT 364.400 381.600 365.200 384.200 ;
        RECT 367.600 381.600 368.400 386.200 ;
        RECT 372.400 381.600 373.200 386.200 ;
        RECT 375.600 381.600 376.400 386.200 ;
        RECT 378.800 381.600 379.600 386.200 ;
        RECT 382.000 381.600 382.800 386.200 ;
        RECT 385.200 381.600 386.000 386.200 ;
        RECT 388.400 381.600 389.200 386.200 ;
        RECT 391.600 381.600 392.400 386.000 ;
        RECT 397.200 381.600 398.000 384.200 ;
        RECT 400.400 381.600 401.400 384.200 ;
        RECT 406.000 381.600 406.800 386.200 ;
        RECT 410.800 381.600 411.600 386.200 ;
        RECT 415.600 381.600 416.400 386.200 ;
        RECT 420.400 381.600 421.200 386.200 ;
        RECT 425.200 381.600 426.000 386.200 ;
        RECT 430.000 381.600 430.800 386.200 ;
        RECT 433.200 381.600 434.000 386.200 ;
        RECT 442.800 381.600 443.600 384.200 ;
        RECT 449.200 381.600 450.000 386.200 ;
        RECT 460.400 381.600 461.200 384.200 ;
        RECT 463.600 381.600 464.400 384.200 ;
        RECT 473.200 381.600 474.000 386.200 ;
        RECT 481.200 381.600 482.000 386.200 ;
        RECT 484.400 381.600 485.200 385.800 ;
        RECT 487.600 381.600 488.400 384.200 ;
        RECT 492.400 381.600 493.200 386.200 ;
        RECT 494.000 381.600 494.800 386.200 ;
        RECT 497.200 381.600 498.000 386.200 ;
        RECT 500.400 381.600 501.200 386.200 ;
        RECT 503.600 381.600 504.400 386.200 ;
        RECT 508.400 381.600 509.200 386.200 ;
        RECT 514.800 381.600 515.600 386.200 ;
        RECT 524.400 381.600 525.200 384.200 ;
        RECT 527.600 381.600 528.400 384.200 ;
        RECT 538.800 381.600 539.600 386.200 ;
        RECT 545.200 381.600 546.000 384.200 ;
        RECT 550.000 381.600 550.800 386.200 ;
        RECT 559.600 381.600 560.400 384.200 ;
        RECT 562.800 381.600 563.600 384.200 ;
        RECT 574.000 381.600 574.800 386.200 ;
        RECT 580.400 381.600 581.200 384.200 ;
        RECT 0.400 380.400 586.800 381.600 ;
        RECT 1.200 375.800 2.000 380.400 ;
        RECT 9.200 376.600 10.000 380.400 ;
        RECT 12.400 377.800 13.200 380.400 ;
        RECT 15.600 377.800 16.400 380.400 ;
        RECT 18.800 377.800 19.600 380.400 ;
        RECT 23.600 376.600 24.400 380.400 ;
        RECT 30.000 375.800 30.800 380.400 ;
        RECT 31.600 377.800 32.400 380.400 ;
        RECT 34.800 377.800 35.600 380.400 ;
        RECT 38.000 376.600 38.800 380.400 ;
        RECT 46.000 376.600 46.800 380.400 ;
        RECT 50.800 376.000 51.600 380.400 ;
        RECT 56.400 377.800 57.200 380.400 ;
        RECT 59.600 377.800 60.600 380.400 ;
        RECT 65.200 375.800 66.000 380.400 ;
        RECT 70.600 376.000 71.400 380.400 ;
        RECT 76.400 375.800 77.200 380.400 ;
        RECT 79.600 376.000 80.400 380.400 ;
        RECT 85.200 377.800 86.000 380.400 ;
        RECT 88.400 377.800 89.400 380.400 ;
        RECT 94.000 375.800 94.800 380.400 ;
        RECT 98.800 376.000 99.600 380.400 ;
        RECT 104.400 377.800 105.200 380.400 ;
        RECT 107.600 377.800 108.600 380.400 ;
        RECT 113.200 375.800 114.000 380.400 ;
        RECT 118.000 376.000 118.800 380.400 ;
        RECT 123.600 377.800 124.400 380.400 ;
        RECT 126.800 377.800 127.800 380.400 ;
        RECT 132.400 375.800 133.200 380.400 ;
        RECT 142.000 376.000 142.800 380.400 ;
        RECT 147.600 377.800 148.400 380.400 ;
        RECT 150.800 377.800 151.800 380.400 ;
        RECT 156.400 375.800 157.200 380.400 ;
        RECT 161.200 376.400 162.200 380.400 ;
        RECT 167.400 379.800 168.200 380.400 ;
        RECT 167.400 376.400 168.400 379.800 ;
        RECT 172.000 375.000 172.800 380.400 ;
        RECT 177.200 375.400 178.000 380.400 ;
        RECT 180.400 377.800 181.200 380.400 ;
        RECT 183.600 377.800 184.400 380.400 ;
        RECT 185.800 375.800 186.600 380.400 ;
        RECT 190.000 377.800 190.800 380.400 ;
        RECT 194.800 375.800 195.600 380.400 ;
        RECT 196.400 375.800 197.200 380.400 ;
        RECT 201.200 375.800 202.000 380.400 ;
        RECT 207.600 376.600 208.400 380.400 ;
        RECT 212.400 375.800 213.200 380.400 ;
        RECT 220.400 375.800 221.200 380.400 ;
        RECT 223.600 375.800 224.400 380.400 ;
        RECT 228.400 375.800 229.200 380.400 ;
        RECT 231.800 379.800 232.600 380.400 ;
        RECT 231.600 376.400 232.600 379.800 ;
        RECT 237.800 376.400 238.800 380.400 ;
        RECT 242.800 377.800 243.600 380.400 ;
        RECT 244.400 375.800 245.200 380.400 ;
        RECT 247.600 375.800 248.400 380.400 ;
        RECT 255.600 376.600 256.400 380.400 ;
        RECT 258.800 375.800 259.600 380.400 ;
        RECT 266.800 376.600 267.600 380.400 ;
        RECT 270.000 377.800 270.800 380.400 ;
        RECT 274.200 375.800 275.000 380.400 ;
        RECT 278.000 377.800 278.800 380.400 ;
        RECT 281.200 376.600 282.000 380.400 ;
        RECT 289.200 375.800 290.000 380.400 ;
        RECT 297.200 375.800 298.000 380.400 ;
        RECT 300.400 375.800 301.200 380.400 ;
        RECT 302.000 377.800 302.800 380.400 ;
        RECT 306.800 376.600 307.600 380.400 ;
        RECT 313.200 376.000 314.000 380.400 ;
        RECT 318.800 377.800 319.600 380.400 ;
        RECT 322.000 377.800 323.000 380.400 ;
        RECT 327.600 375.800 328.400 380.400 ;
        RECT 332.400 376.000 333.200 380.400 ;
        RECT 338.000 377.800 338.800 380.400 ;
        RECT 341.200 377.800 342.200 380.400 ;
        RECT 346.800 375.800 347.600 380.400 ;
        RECT 351.600 376.600 352.400 380.400 ;
        RECT 358.000 375.800 358.800 380.400 ;
        RECT 362.800 376.600 363.600 380.400 ;
        RECT 367.600 377.800 368.400 380.400 ;
        RECT 370.800 377.800 371.600 380.400 ;
        RECT 372.400 377.800 373.200 380.400 ;
        RECT 375.600 377.800 376.400 380.400 ;
        RECT 380.400 376.600 381.200 380.400 ;
        RECT 385.200 377.800 386.000 380.400 ;
        RECT 388.400 376.000 389.200 380.400 ;
        RECT 394.000 377.800 394.800 380.400 ;
        RECT 397.200 377.800 398.200 380.400 ;
        RECT 402.800 375.800 403.600 380.400 ;
        RECT 406.000 375.800 406.800 380.400 ;
        RECT 409.200 375.800 410.000 380.400 ;
        RECT 410.800 377.800 411.600 380.400 ;
        RECT 417.200 375.800 418.000 380.400 ;
        RECT 428.400 377.800 429.200 380.400 ;
        RECT 431.600 377.800 432.400 380.400 ;
        RECT 441.200 375.800 442.000 380.400 ;
        RECT 452.400 376.200 453.200 380.400 ;
        RECT 455.600 377.800 456.400 380.400 ;
        RECT 457.200 377.800 458.000 380.400 ;
        RECT 463.600 375.800 464.400 380.400 ;
        RECT 474.800 377.800 475.600 380.400 ;
        RECT 478.000 377.800 478.800 380.400 ;
        RECT 487.600 375.800 488.400 380.400 ;
        RECT 494.000 376.200 494.800 380.400 ;
        RECT 497.200 377.800 498.000 380.400 ;
        RECT 502.000 375.800 502.800 380.400 ;
        RECT 511.600 377.800 512.400 380.400 ;
        RECT 514.800 377.800 515.600 380.400 ;
        RECT 526.000 375.800 526.800 380.400 ;
        RECT 532.400 377.800 533.200 380.400 ;
        RECT 534.000 375.800 534.800 380.400 ;
        RECT 537.200 375.800 538.000 380.400 ;
        RECT 540.400 375.800 541.200 380.400 ;
        RECT 543.600 375.800 544.400 380.400 ;
        RECT 546.800 375.800 547.600 380.400 ;
        RECT 551.600 375.800 552.400 380.400 ;
        RECT 561.200 377.800 562.000 380.400 ;
        RECT 564.400 377.800 565.200 380.400 ;
        RECT 575.600 375.800 576.400 380.400 ;
        RECT 582.000 377.800 582.800 380.400 ;
        RECT 4.400 341.600 5.200 345.400 ;
        RECT 9.200 342.200 10.200 345.600 ;
        RECT 9.400 341.600 10.200 342.200 ;
        RECT 15.400 341.600 16.400 345.600 ;
        RECT 18.800 341.600 19.600 344.200 ;
        RECT 23.600 342.200 24.600 345.600 ;
        RECT 23.800 341.600 24.600 342.200 ;
        RECT 29.800 341.600 30.800 345.600 ;
        RECT 33.200 341.600 34.000 344.200 ;
        RECT 36.400 341.600 37.200 344.200 ;
        RECT 39.600 341.600 40.400 345.800 ;
        RECT 42.800 341.600 43.600 344.200 ;
        RECT 47.000 341.600 47.800 346.200 ;
        RECT 52.400 341.600 53.200 345.400 ;
        RECT 57.200 341.600 58.000 345.400 ;
        RECT 62.600 341.600 63.400 346.200 ;
        RECT 66.800 341.600 67.600 344.200 ;
        RECT 68.400 341.600 69.200 344.200 ;
        RECT 71.600 341.600 72.400 344.200 ;
        RECT 73.200 341.600 74.000 344.200 ;
        RECT 76.400 341.600 77.200 344.200 ;
        RECT 78.600 341.600 79.400 346.200 ;
        RECT 82.800 341.600 83.600 344.200 ;
        RECT 84.400 341.600 85.200 344.200 ;
        RECT 87.600 341.600 88.400 344.200 ;
        RECT 92.400 341.600 93.200 346.200 ;
        RECT 95.600 341.600 96.400 346.000 ;
        RECT 101.200 341.600 102.000 344.200 ;
        RECT 104.400 341.600 105.400 344.200 ;
        RECT 110.000 341.600 110.800 346.200 ;
        RECT 116.400 341.600 117.200 346.200 ;
        RECT 119.600 341.600 120.400 346.200 ;
        RECT 122.800 342.200 123.800 345.600 ;
        RECT 123.000 341.600 123.800 342.200 ;
        RECT 129.000 341.600 130.000 345.600 ;
        RECT 132.400 341.600 133.200 346.200 ;
        RECT 143.600 342.200 144.600 345.600 ;
        RECT 143.800 341.600 144.600 342.200 ;
        RECT 149.800 341.600 150.800 345.600 ;
        RECT 154.800 341.600 155.600 346.000 ;
        RECT 160.400 341.600 161.200 344.200 ;
        RECT 163.600 341.600 164.600 344.200 ;
        RECT 169.200 341.600 170.000 346.200 ;
        RECT 174.000 341.600 174.800 346.000 ;
        RECT 179.600 341.600 180.400 344.200 ;
        RECT 182.800 341.600 183.800 344.200 ;
        RECT 188.400 341.600 189.200 346.200 ;
        RECT 191.600 341.600 192.400 344.200 ;
        RECT 194.800 341.600 195.600 344.200 ;
        RECT 198.000 342.200 199.000 345.600 ;
        RECT 198.200 341.600 199.000 342.200 ;
        RECT 204.200 341.600 205.200 345.600 ;
        RECT 212.400 341.600 213.200 345.400 ;
        RECT 215.600 341.600 216.400 344.200 ;
        RECT 219.800 341.600 220.600 346.200 ;
        RECT 223.600 342.200 224.600 345.600 ;
        RECT 223.800 341.600 224.600 342.200 ;
        RECT 229.800 341.600 230.800 345.600 ;
        RECT 236.400 341.600 237.200 345.400 ;
        RECT 242.800 341.600 243.600 346.200 ;
        RECT 244.400 341.600 245.200 346.200 ;
        RECT 249.200 341.600 250.000 346.200 ;
        RECT 252.400 341.600 253.200 346.200 ;
        RECT 254.000 341.600 254.800 346.200 ;
        RECT 257.200 341.600 258.000 346.200 ;
        RECT 260.400 341.600 261.200 346.200 ;
        RECT 263.600 341.600 264.400 346.200 ;
        RECT 266.800 342.200 267.800 345.600 ;
        RECT 267.000 341.600 267.800 342.200 ;
        RECT 273.000 341.600 274.000 345.600 ;
        RECT 278.000 341.600 278.800 345.400 ;
        RECT 286.000 341.600 286.800 346.200 ;
        RECT 293.000 341.600 293.800 346.200 ;
        RECT 297.200 341.600 298.000 344.200 ;
        RECT 298.800 341.600 299.600 344.200 ;
        RECT 302.000 341.600 302.800 344.200 ;
        RECT 305.200 341.600 306.000 345.800 ;
        RECT 308.400 341.600 309.200 344.200 ;
        RECT 310.000 341.600 310.800 344.200 ;
        RECT 313.200 341.600 314.000 344.200 ;
        RECT 314.800 341.600 315.600 344.200 ;
        RECT 318.000 341.600 318.800 344.200 ;
        RECT 321.200 341.600 322.000 344.200 ;
        RECT 326.000 341.600 326.800 345.400 ;
        RECT 330.800 341.600 331.600 344.200 ;
        RECT 334.000 341.600 334.800 346.000 ;
        RECT 339.600 341.600 340.400 344.200 ;
        RECT 342.800 341.600 343.800 344.200 ;
        RECT 348.400 341.600 349.200 346.200 ;
        RECT 353.200 341.600 354.000 344.200 ;
        RECT 356.400 341.600 357.200 346.000 ;
        RECT 362.000 341.600 362.800 344.200 ;
        RECT 365.200 341.600 366.200 344.200 ;
        RECT 370.800 341.600 371.600 346.200 ;
        RECT 375.600 341.600 376.400 346.200 ;
        RECT 380.400 342.200 381.400 345.600 ;
        RECT 380.600 341.600 381.400 342.200 ;
        RECT 386.600 341.600 387.600 345.600 ;
        RECT 391.600 341.600 392.400 346.200 ;
        RECT 394.800 341.600 395.600 346.000 ;
        RECT 400.400 341.600 401.200 344.200 ;
        RECT 403.600 341.600 404.600 344.200 ;
        RECT 409.200 341.600 410.000 346.200 ;
        RECT 415.600 341.600 416.400 345.400 ;
        RECT 422.000 341.600 422.800 345.400 ;
        RECT 426.800 341.600 427.600 345.400 ;
        RECT 434.800 341.600 435.600 345.400 ;
        RECT 439.600 341.600 440.400 344.200 ;
        RECT 442.800 341.600 443.600 344.200 ;
        RECT 449.200 341.600 450.000 344.200 ;
        RECT 452.400 341.600 453.200 344.200 ;
        RECT 454.000 341.600 454.800 346.200 ;
        RECT 458.800 341.600 459.600 344.200 ;
        RECT 463.000 341.600 463.800 346.200 ;
        RECT 465.200 341.600 466.000 346.200 ;
        RECT 471.600 341.600 472.600 345.600 ;
        RECT 477.800 342.200 478.800 345.600 ;
        RECT 477.800 341.600 478.600 342.200 ;
        RECT 482.800 341.600 483.600 346.000 ;
        RECT 488.400 341.600 489.200 344.200 ;
        RECT 491.600 341.600 492.600 344.200 ;
        RECT 497.200 341.600 498.000 346.200 ;
        RECT 500.400 341.600 501.200 346.200 ;
        RECT 503.600 341.600 504.400 346.200 ;
        RECT 506.800 341.600 507.600 346.200 ;
        RECT 510.000 341.600 510.800 346.200 ;
        RECT 513.200 341.600 514.000 346.200 ;
        RECT 518.000 341.600 518.800 346.200 ;
        RECT 527.600 341.600 528.400 344.200 ;
        RECT 530.800 341.600 531.600 344.200 ;
        RECT 542.000 341.600 542.800 346.200 ;
        RECT 548.400 341.600 549.200 344.200 ;
        RECT 553.200 341.600 554.000 346.200 ;
        RECT 562.800 341.600 563.600 344.200 ;
        RECT 566.000 341.600 566.800 344.200 ;
        RECT 577.200 341.600 578.000 346.200 ;
        RECT 583.600 341.600 584.400 344.200 ;
        RECT 0.400 340.400 586.800 341.600 ;
        RECT 3.000 339.800 3.800 340.400 ;
        RECT 2.800 336.400 3.800 339.800 ;
        RECT 9.000 336.400 10.000 340.400 ;
        RECT 12.400 335.800 13.200 340.400 ;
        RECT 15.600 335.800 16.400 340.400 ;
        RECT 18.800 335.800 19.600 340.400 ;
        RECT 20.400 335.800 21.200 340.400 ;
        RECT 23.600 335.800 24.400 340.400 ;
        RECT 26.800 337.800 27.600 340.400 ;
        RECT 31.600 335.800 32.400 340.400 ;
        RECT 34.800 335.800 35.600 340.400 ;
        RECT 36.800 335.800 37.600 340.400 ;
        RECT 42.800 335.800 43.600 340.400 ;
        RECT 47.600 336.600 48.400 340.400 ;
        RECT 55.600 333.800 56.400 340.400 ;
        RECT 58.800 337.800 59.600 340.400 ;
        RECT 60.400 337.800 61.200 340.400 ;
        RECT 63.600 335.800 64.400 340.400 ;
        RECT 73.200 333.800 74.000 340.400 ;
        RECT 78.000 336.600 78.800 340.400 ;
        RECT 81.200 335.800 82.000 340.400 ;
        RECT 89.200 335.800 90.000 340.400 ;
        RECT 94.000 336.600 94.800 340.400 ;
        RECT 100.400 336.600 101.200 340.400 ;
        RECT 103.600 337.800 104.400 340.400 ;
        RECT 106.800 337.800 107.600 340.400 ;
        RECT 110.000 336.600 110.800 340.400 ;
        RECT 116.400 337.800 117.200 340.400 ;
        RECT 122.800 336.600 123.600 340.400 ;
        RECT 127.600 336.600 128.400 340.400 ;
        RECT 135.600 336.600 136.400 340.400 ;
        RECT 145.400 339.800 146.200 340.400 ;
        RECT 145.200 336.400 146.200 339.800 ;
        RECT 151.400 336.400 152.400 340.400 ;
        RECT 155.400 335.800 156.200 340.400 ;
        RECT 159.600 337.800 160.400 340.400 ;
        RECT 162.800 337.800 163.600 340.400 ;
        RECT 164.400 337.800 165.200 340.400 ;
        RECT 170.800 336.600 171.600 340.400 ;
        RECT 175.600 336.400 176.600 340.400 ;
        RECT 181.800 339.800 182.600 340.400 ;
        RECT 181.800 336.400 182.800 339.800 ;
        RECT 185.200 335.800 186.000 340.400 ;
        RECT 188.400 335.800 189.200 340.400 ;
        RECT 191.600 335.800 192.400 340.400 ;
        RECT 194.800 335.800 195.600 340.400 ;
        RECT 198.000 335.800 198.800 340.400 ;
        RECT 201.200 336.000 202.000 340.400 ;
        RECT 206.800 337.800 207.600 340.400 ;
        RECT 210.000 337.800 211.000 340.400 ;
        RECT 215.600 335.800 216.400 340.400 ;
        RECT 220.400 336.400 221.400 340.400 ;
        RECT 226.600 339.800 227.400 340.400 ;
        RECT 226.600 336.400 227.600 339.800 ;
        RECT 231.600 336.400 232.600 340.400 ;
        RECT 237.800 339.800 238.600 340.400 ;
        RECT 237.800 336.400 238.800 339.800 ;
        RECT 244.400 336.600 245.200 340.400 ;
        RECT 250.800 335.800 251.600 340.400 ;
        RECT 252.400 333.800 253.200 340.400 ;
        RECT 262.000 335.800 262.800 340.400 ;
        RECT 264.200 335.800 265.000 340.400 ;
        RECT 268.400 337.800 269.200 340.400 ;
        RECT 270.000 337.800 270.800 340.400 ;
        RECT 273.200 337.800 274.000 340.400 ;
        RECT 276.400 336.600 277.200 340.400 ;
        RECT 281.200 337.800 282.000 340.400 ;
        RECT 285.000 335.800 285.800 340.400 ;
        RECT 289.200 337.800 290.000 340.400 ;
        RECT 295.600 337.800 296.400 340.400 ;
        RECT 298.800 337.800 299.600 340.400 ;
        RECT 302.000 336.600 302.800 340.400 ;
        RECT 306.800 335.800 307.600 340.400 ;
        RECT 311.600 337.800 312.400 340.400 ;
        RECT 315.800 335.800 316.600 340.400 ;
        RECT 318.000 337.800 318.800 340.400 ;
        RECT 321.200 337.800 322.000 340.400 ;
        RECT 324.600 339.800 325.400 340.400 ;
        RECT 324.400 336.400 325.400 339.800 ;
        RECT 330.600 336.400 331.600 340.400 ;
        RECT 335.600 336.000 336.400 340.400 ;
        RECT 341.200 337.800 342.000 340.400 ;
        RECT 344.400 337.800 345.400 340.400 ;
        RECT 350.000 335.800 350.800 340.400 ;
        RECT 354.800 337.800 355.600 340.400 ;
        RECT 358.000 336.000 358.800 340.400 ;
        RECT 363.600 337.800 364.400 340.400 ;
        RECT 366.800 337.800 367.800 340.400 ;
        RECT 372.400 335.800 373.200 340.400 ;
        RECT 377.200 336.600 378.000 340.400 ;
        RECT 386.800 336.600 387.600 340.400 ;
        RECT 390.000 335.800 390.800 340.400 ;
        RECT 396.400 336.000 397.200 340.400 ;
        RECT 402.000 337.800 402.800 340.400 ;
        RECT 405.200 337.800 406.200 340.400 ;
        RECT 410.800 335.800 411.600 340.400 ;
        RECT 415.600 336.000 416.400 340.400 ;
        RECT 421.200 337.800 422.000 340.400 ;
        RECT 424.400 337.800 425.400 340.400 ;
        RECT 430.000 335.800 430.800 340.400 ;
        RECT 435.000 339.800 435.800 340.400 ;
        RECT 434.800 336.400 435.800 339.800 ;
        RECT 441.000 336.400 442.000 340.400 ;
        RECT 450.800 335.800 451.600 340.400 ;
        RECT 455.600 336.600 456.400 340.400 ;
        RECT 460.400 337.800 461.200 340.400 ;
        RECT 463.600 337.800 464.400 340.400 ;
        RECT 468.400 335.800 469.200 340.400 ;
        RECT 471.600 336.600 472.400 340.400 ;
        RECT 478.000 335.800 478.800 340.400 ;
        RECT 483.400 337.800 484.400 340.400 ;
        RECT 486.800 337.800 487.600 340.400 ;
        RECT 492.400 336.000 493.200 340.400 ;
        RECT 497.200 335.800 498.000 340.400 ;
        RECT 502.600 337.800 503.600 340.400 ;
        RECT 506.000 337.800 506.800 340.400 ;
        RECT 511.600 336.000 512.400 340.400 ;
        RECT 516.400 335.800 517.200 340.400 ;
        RECT 519.600 337.800 520.400 340.400 ;
        RECT 526.000 335.800 526.800 340.400 ;
        RECT 537.200 337.800 538.000 340.400 ;
        RECT 540.400 337.800 541.200 340.400 ;
        RECT 550.000 335.800 550.800 340.400 ;
        RECT 556.400 336.000 557.200 340.400 ;
        RECT 562.000 337.800 562.800 340.400 ;
        RECT 565.200 337.800 566.200 340.400 ;
        RECT 570.800 335.800 571.600 340.400 ;
        RECT 575.600 335.800 576.400 340.400 ;
        RECT 580.400 335.800 581.200 340.400 ;
        RECT 222.000 308.800 222.800 310.400 ;
        RECT 4.400 301.600 5.200 305.400 ;
        RECT 7.600 301.600 8.400 304.200 ;
        RECT 10.800 301.600 11.600 304.200 ;
        RECT 12.400 301.600 13.200 304.200 ;
        RECT 15.600 301.600 16.400 304.200 ;
        RECT 17.200 301.600 18.000 306.200 ;
        RECT 20.400 301.600 21.200 304.200 ;
        RECT 23.600 301.600 24.400 304.200 ;
        RECT 28.400 301.600 29.200 305.400 ;
        RECT 34.800 301.600 35.600 306.200 ;
        RECT 36.400 301.600 37.200 304.200 ;
        RECT 39.600 301.600 40.400 304.200 ;
        RECT 41.200 301.600 42.000 306.200 ;
        RECT 49.200 301.600 50.000 305.400 ;
        RECT 54.000 302.200 55.000 305.600 ;
        RECT 54.200 301.600 55.000 302.200 ;
        RECT 60.200 301.600 61.200 305.600 ;
        RECT 66.800 301.600 67.600 306.200 ;
        RECT 68.400 301.600 69.200 304.200 ;
        RECT 73.200 301.600 74.000 306.200 ;
        RECT 76.400 301.600 77.200 306.200 ;
        RECT 78.000 301.600 78.800 306.200 ;
        RECT 84.000 301.600 84.800 306.200 ;
        RECT 86.000 301.600 86.800 306.200 ;
        RECT 92.400 301.600 93.200 304.200 ;
        RECT 95.600 301.600 96.400 305.400 ;
        RECT 100.400 301.600 101.200 304.200 ;
        RECT 103.600 301.600 104.400 304.200 ;
        RECT 106.800 301.600 107.600 305.400 ;
        RECT 112.200 301.600 113.000 306.200 ;
        RECT 116.400 301.600 117.200 304.200 ;
        RECT 119.600 301.600 120.400 305.400 ;
        RECT 124.400 301.600 125.200 304.200 ;
        RECT 130.800 301.600 131.600 306.200 ;
        RECT 134.000 301.600 134.800 304.200 ;
        RECT 143.600 301.600 144.400 305.400 ;
        RECT 146.800 301.600 147.600 306.200 ;
        RECT 154.800 301.600 155.600 305.400 ;
        RECT 158.000 301.600 158.800 304.200 ;
        RECT 161.200 301.600 162.000 304.200 ;
        RECT 164.400 301.600 165.200 305.800 ;
        RECT 167.600 301.600 168.400 304.200 ;
        RECT 169.200 301.600 170.000 304.200 ;
        RECT 172.400 301.600 173.200 304.200 ;
        RECT 176.600 301.600 177.400 306.000 ;
        RECT 182.000 301.600 182.800 306.000 ;
        RECT 187.600 301.600 188.400 304.200 ;
        RECT 190.800 301.600 191.800 304.200 ;
        RECT 196.400 301.600 197.200 306.200 ;
        RECT 201.200 301.600 202.000 306.000 ;
        RECT 206.800 301.600 207.600 304.200 ;
        RECT 210.000 301.600 211.000 304.200 ;
        RECT 215.600 301.600 216.400 306.200 ;
        RECT 220.400 301.600 221.200 306.200 ;
        RECT 225.200 301.600 226.000 306.200 ;
        RECT 231.600 301.600 232.400 305.400 ;
        RECT 238.000 301.600 238.800 305.400 ;
        RECT 241.200 301.600 242.000 304.200 ;
        RECT 245.400 301.600 246.200 306.200 ;
        RECT 249.200 301.600 250.000 304.200 ;
        RECT 252.400 301.600 253.200 305.400 ;
        RECT 258.400 301.600 259.200 307.000 ;
        RECT 263.600 301.600 264.400 306.600 ;
        RECT 266.800 301.600 267.600 306.200 ;
        RECT 270.000 301.600 270.800 306.200 ;
        RECT 274.800 301.600 275.600 306.000 ;
        RECT 280.400 301.600 281.200 304.200 ;
        RECT 283.600 301.600 284.600 304.200 ;
        RECT 289.200 301.600 290.000 306.200 ;
        RECT 298.800 301.600 299.600 306.000 ;
        RECT 304.400 301.600 305.200 304.200 ;
        RECT 307.600 301.600 308.600 304.200 ;
        RECT 313.200 301.600 314.000 306.200 ;
        RECT 318.000 301.600 318.800 306.200 ;
        RECT 321.200 301.600 322.000 306.200 ;
        RECT 326.000 301.600 326.800 306.200 ;
        RECT 330.800 301.600 331.600 306.200 ;
        RECT 335.600 301.600 336.400 305.400 ;
        RECT 342.000 301.600 342.800 305.400 ;
        RECT 348.400 301.600 349.200 305.400 ;
        RECT 353.200 301.600 354.000 304.200 ;
        RECT 356.400 301.600 357.400 305.600 ;
        RECT 362.600 302.200 363.600 305.600 ;
        RECT 367.600 302.200 368.600 305.600 ;
        RECT 362.600 301.600 363.400 302.200 ;
        RECT 367.800 301.600 368.600 302.200 ;
        RECT 373.800 301.600 374.800 305.600 ;
        RECT 377.200 301.600 378.000 306.200 ;
        RECT 382.000 301.600 382.800 304.200 ;
        RECT 385.200 301.600 386.000 304.200 ;
        RECT 391.600 301.600 392.400 305.400 ;
        RECT 396.400 301.600 397.200 304.200 ;
        RECT 399.600 301.600 400.400 305.800 ;
        RECT 402.800 301.600 403.600 304.200 ;
        RECT 406.000 301.600 406.800 306.000 ;
        RECT 411.600 301.600 412.400 304.200 ;
        RECT 414.800 301.600 415.800 304.200 ;
        RECT 420.400 301.600 421.200 306.200 ;
        RECT 423.600 301.600 424.400 306.200 ;
        RECT 429.600 301.600 430.400 306.200 ;
        RECT 431.600 301.600 432.400 304.200 ;
        RECT 438.000 301.600 438.800 305.400 ;
        RECT 441.200 301.600 442.000 306.200 ;
        RECT 450.800 301.600 451.600 306.200 ;
        RECT 458.800 301.600 459.600 305.400 ;
        RECT 463.600 301.600 464.400 304.200 ;
        RECT 466.800 301.600 467.800 305.600 ;
        RECT 473.000 302.200 474.000 305.600 ;
        RECT 473.000 301.600 473.800 302.200 ;
        RECT 478.000 301.600 478.800 304.200 ;
        RECT 481.200 301.600 482.000 306.200 ;
        RECT 486.600 301.600 487.600 304.200 ;
        RECT 490.000 301.600 490.800 304.200 ;
        RECT 495.600 301.600 496.400 306.000 ;
        RECT 498.800 301.600 499.600 304.200 ;
        RECT 505.200 301.600 506.000 306.200 ;
        RECT 516.400 301.600 517.200 304.200 ;
        RECT 519.600 301.600 520.400 304.200 ;
        RECT 529.200 301.600 530.000 306.200 ;
        RECT 537.200 301.600 538.000 306.200 ;
        RECT 540.400 301.600 541.200 305.800 ;
        RECT 543.600 301.600 544.400 304.200 ;
        RECT 546.800 301.600 547.600 306.200 ;
        RECT 552.200 301.600 553.200 304.200 ;
        RECT 555.600 301.600 556.400 304.200 ;
        RECT 561.200 301.600 562.000 306.000 ;
        RECT 566.000 301.600 566.800 306.200 ;
        RECT 571.400 301.600 572.400 304.200 ;
        RECT 574.800 301.600 575.600 304.200 ;
        RECT 580.400 301.600 581.200 306.000 ;
        RECT 0.400 300.400 586.800 301.600 ;
        RECT 1.200 297.800 2.000 300.400 ;
        RECT 6.000 297.800 6.800 300.400 ;
        RECT 10.800 296.600 11.600 300.400 ;
        RECT 18.800 293.800 19.600 300.400 ;
        RECT 22.000 296.600 22.800 300.400 ;
        RECT 28.400 297.800 29.200 300.400 ;
        RECT 33.200 296.600 34.000 300.400 ;
        RECT 36.400 297.800 37.200 300.400 ;
        RECT 40.600 295.800 41.400 300.400 ;
        RECT 43.200 295.800 44.000 300.400 ;
        RECT 49.200 295.800 50.000 300.400 ;
        RECT 52.400 296.600 53.200 300.400 ;
        RECT 60.400 296.600 61.200 300.400 ;
        RECT 65.200 296.600 66.000 300.400 ;
        RECT 73.200 295.800 74.000 300.400 ;
        RECT 74.800 297.800 75.600 300.400 ;
        RECT 78.000 297.800 78.800 300.400 ;
        RECT 79.600 295.800 80.400 300.400 ;
        RECT 85.600 295.800 86.400 300.400 ;
        RECT 87.600 295.800 88.400 300.400 ;
        RECT 94.000 296.400 95.000 300.400 ;
        RECT 100.200 299.800 101.000 300.400 ;
        RECT 100.200 296.400 101.200 299.800 ;
        RECT 105.200 295.800 106.000 300.400 ;
        RECT 108.400 296.600 109.200 300.400 ;
        RECT 113.200 297.800 114.000 300.400 ;
        RECT 116.400 297.800 117.200 300.400 ;
        RECT 120.600 295.800 121.400 300.400 ;
        RECT 126.000 296.600 126.800 300.400 ;
        RECT 129.200 295.800 130.000 300.400 ;
        RECT 134.000 295.800 134.800 300.400 ;
        RECT 146.800 295.800 147.600 300.400 ;
        RECT 148.400 297.800 149.200 300.400 ;
        RECT 151.600 297.800 152.400 300.400 ;
        RECT 153.800 295.800 154.600 300.400 ;
        RECT 158.000 297.800 158.800 300.400 ;
        RECT 161.200 296.600 162.000 300.400 ;
        RECT 167.600 297.800 168.400 300.400 ;
        RECT 169.200 297.800 170.000 300.400 ;
        RECT 173.400 295.800 174.200 300.400 ;
        RECT 175.600 297.800 176.400 300.400 ;
        RECT 178.800 297.800 179.600 300.400 ;
        RECT 182.000 296.600 182.800 300.400 ;
        RECT 188.600 299.800 189.400 300.400 ;
        RECT 188.400 296.400 189.400 299.800 ;
        RECT 194.600 296.400 195.600 300.400 ;
        RECT 199.600 296.000 200.400 300.400 ;
        RECT 205.200 297.800 206.000 300.400 ;
        RECT 208.400 297.800 209.400 300.400 ;
        RECT 214.000 295.800 214.800 300.400 ;
        RECT 218.800 295.800 219.600 300.400 ;
        RECT 223.600 295.800 224.400 300.400 ;
        RECT 228.400 295.800 229.200 300.400 ;
        RECT 233.800 297.800 234.800 300.400 ;
        RECT 237.200 297.800 238.000 300.400 ;
        RECT 242.800 296.000 243.600 300.400 ;
        RECT 247.600 296.400 248.600 300.400 ;
        RECT 253.800 299.800 254.600 300.400 ;
        RECT 253.800 296.400 254.800 299.800 ;
        RECT 258.800 296.000 259.600 300.400 ;
        RECT 264.400 297.800 265.200 300.400 ;
        RECT 267.600 297.800 268.600 300.400 ;
        RECT 273.200 295.800 274.000 300.400 ;
        RECT 278.000 296.000 278.800 300.400 ;
        RECT 283.600 297.800 284.400 300.400 ;
        RECT 286.800 297.800 287.800 300.400 ;
        RECT 292.400 295.800 293.200 300.400 ;
        RECT 300.400 295.800 301.200 300.400 ;
        RECT 306.800 296.400 307.800 300.400 ;
        RECT 313.000 299.800 313.800 300.400 ;
        RECT 313.000 296.400 314.000 299.800 ;
        RECT 319.600 296.600 320.400 300.400 ;
        RECT 324.400 296.200 325.200 300.400 ;
        RECT 327.600 297.800 328.400 300.400 ;
        RECT 330.800 296.000 331.600 300.400 ;
        RECT 336.400 297.800 337.200 300.400 ;
        RECT 339.600 297.800 340.600 300.400 ;
        RECT 345.200 295.800 346.000 300.400 ;
        RECT 350.000 296.000 350.800 300.400 ;
        RECT 355.600 297.800 356.400 300.400 ;
        RECT 358.800 297.800 359.800 300.400 ;
        RECT 364.400 295.800 365.200 300.400 ;
        RECT 369.200 296.000 370.000 300.400 ;
        RECT 374.800 297.800 375.600 300.400 ;
        RECT 378.000 297.800 379.000 300.400 ;
        RECT 383.600 295.800 384.400 300.400 ;
        RECT 388.400 296.400 389.400 300.400 ;
        RECT 394.600 299.800 395.400 300.400 ;
        RECT 394.600 296.400 395.600 299.800 ;
        RECT 401.200 296.600 402.000 300.400 ;
        RECT 404.400 297.800 405.200 300.400 ;
        RECT 410.800 296.600 411.600 300.400 ;
        RECT 415.600 296.000 416.400 300.400 ;
        RECT 421.200 297.800 422.000 300.400 ;
        RECT 424.400 297.800 425.400 300.400 ;
        RECT 430.000 295.800 430.800 300.400 ;
        RECT 434.800 296.400 435.800 300.400 ;
        RECT 441.000 299.800 441.800 300.400 ;
        RECT 441.000 296.400 442.000 299.800 ;
        RECT 449.200 297.800 450.000 300.400 ;
        RECT 454.000 296.600 454.800 300.400 ;
        RECT 460.400 296.600 461.200 300.400 ;
        RECT 466.800 295.800 467.600 300.400 ;
        RECT 472.200 297.800 473.200 300.400 ;
        RECT 475.600 297.800 476.400 300.400 ;
        RECT 481.200 296.000 482.000 300.400 ;
        RECT 486.000 296.400 487.000 300.400 ;
        RECT 492.200 299.800 493.000 300.400 ;
        RECT 492.200 296.400 493.200 299.800 ;
        RECT 495.600 295.800 496.400 300.400 ;
        RECT 498.800 295.800 499.600 300.400 ;
        RECT 502.000 295.800 502.800 300.400 ;
        RECT 505.200 295.800 506.000 300.400 ;
        RECT 508.400 295.800 509.200 300.400 ;
        RECT 511.600 295.800 512.400 300.400 ;
        RECT 517.000 297.800 518.000 300.400 ;
        RECT 520.400 297.800 521.200 300.400 ;
        RECT 526.000 296.000 526.800 300.400 ;
        RECT 530.800 295.800 531.600 300.400 ;
        RECT 534.000 297.800 534.800 300.400 ;
        RECT 540.400 295.800 541.200 300.400 ;
        RECT 551.600 297.800 552.400 300.400 ;
        RECT 554.800 297.800 555.600 300.400 ;
        RECT 564.400 295.800 565.200 300.400 ;
        RECT 569.200 295.800 570.000 300.400 ;
        RECT 575.600 296.200 576.400 300.400 ;
        RECT 578.800 297.800 579.600 300.400 ;
        RECT 582.000 295.800 582.800 300.400 ;
        RECT 220.400 291.600 221.200 293.200 ;
        RECT 222.000 291.600 222.800 293.200 ;
        RECT 229.000 292.400 229.800 292.600 ;
        RECT 229.000 291.800 234.000 292.400 ;
        RECT 233.200 291.600 234.000 291.800 ;
        RECT 1.200 261.600 2.000 264.200 ;
        RECT 5.400 261.600 6.200 266.200 ;
        RECT 9.200 261.600 10.200 265.600 ;
        RECT 15.400 262.200 16.400 265.600 ;
        RECT 15.400 261.600 16.200 262.200 ;
        RECT 18.800 261.600 19.600 264.200 ;
        RECT 25.200 261.600 26.000 265.400 ;
        RECT 28.400 261.600 29.200 264.200 ;
        RECT 34.800 261.600 35.600 265.400 ;
        RECT 38.000 261.600 38.800 264.200 ;
        RECT 42.200 261.600 43.000 266.200 ;
        RECT 46.000 261.600 46.800 264.200 ;
        RECT 48.000 261.600 48.800 266.200 ;
        RECT 54.000 261.600 54.800 266.200 ;
        RECT 55.600 261.600 56.400 264.200 ;
        RECT 60.400 261.600 61.400 265.600 ;
        RECT 66.600 262.200 67.600 265.600 ;
        RECT 66.600 261.600 67.400 262.200 ;
        RECT 71.600 261.600 72.400 266.600 ;
        RECT 76.800 261.600 77.600 267.000 ;
        RECT 82.800 261.600 83.600 265.400 ;
        RECT 87.600 262.200 88.600 265.600 ;
        RECT 87.800 261.600 88.600 262.200 ;
        RECT 93.800 261.600 94.800 265.600 ;
        RECT 97.800 261.600 98.600 266.200 ;
        RECT 102.000 261.600 102.800 264.200 ;
        RECT 105.200 261.600 106.000 264.200 ;
        RECT 106.800 261.600 107.600 264.200 ;
        RECT 110.000 261.600 110.800 264.200 ;
        RECT 113.200 261.600 114.000 266.200 ;
        RECT 116.400 261.600 117.200 266.200 ;
        RECT 121.200 261.600 122.000 265.400 ;
        RECT 124.400 261.600 125.200 266.200 ;
        RECT 130.800 261.600 131.600 265.400 ;
        RECT 134.000 261.600 134.800 266.200 ;
        RECT 145.200 261.600 146.000 265.400 ;
        RECT 153.200 261.600 154.000 265.400 ;
        RECT 158.000 261.600 158.800 264.200 ;
        RECT 164.400 261.600 165.200 265.400 ;
        RECT 169.200 261.600 170.000 265.400 ;
        RECT 177.200 261.600 178.000 266.200 ;
        RECT 180.400 261.600 181.200 266.000 ;
        RECT 186.000 261.600 186.800 264.200 ;
        RECT 189.200 261.600 190.200 264.200 ;
        RECT 194.800 261.600 195.600 266.200 ;
        RECT 199.600 261.600 200.400 266.000 ;
        RECT 205.200 261.600 206.000 264.200 ;
        RECT 208.400 261.600 209.400 264.200 ;
        RECT 214.000 261.600 214.800 266.200 ;
        RECT 218.800 262.200 219.800 265.600 ;
        RECT 219.000 261.600 219.800 262.200 ;
        RECT 225.000 261.600 226.000 265.600 ;
        RECT 229.000 261.600 229.800 266.200 ;
        RECT 233.200 261.600 234.000 264.200 ;
        RECT 234.800 261.600 235.600 264.200 ;
        RECT 238.000 261.600 238.800 264.200 ;
        RECT 242.800 261.600 243.600 265.400 ;
        RECT 249.200 261.600 250.000 265.400 ;
        RECT 254.600 261.600 255.400 266.000 ;
        RECT 262.000 261.600 262.800 266.200 ;
        RECT 265.200 261.600 266.000 265.400 ;
        RECT 271.600 262.200 272.600 265.600 ;
        RECT 271.800 261.600 272.600 262.200 ;
        RECT 277.800 261.600 278.800 265.600 ;
        RECT 282.800 261.600 283.600 264.200 ;
        RECT 286.000 262.200 287.000 265.600 ;
        RECT 286.200 261.600 287.000 262.200 ;
        RECT 292.200 261.600 293.200 265.600 ;
        RECT 300.400 261.600 301.200 264.200 ;
        RECT 303.600 261.600 304.400 264.200 ;
        RECT 305.200 261.600 306.000 264.200 ;
        RECT 308.400 261.600 309.200 264.200 ;
        RECT 311.600 261.600 312.400 264.200 ;
        RECT 316.400 261.600 317.200 265.400 ;
        RECT 324.400 261.600 325.200 265.400 ;
        RECT 329.200 261.600 330.000 264.200 ;
        RECT 334.000 261.600 334.800 266.200 ;
        RECT 337.200 261.600 338.000 265.800 ;
        RECT 340.400 261.600 341.200 264.200 ;
        RECT 343.600 261.600 344.400 266.000 ;
        RECT 349.200 261.600 350.000 264.200 ;
        RECT 352.400 261.600 353.400 264.200 ;
        RECT 358.000 261.600 358.800 266.200 ;
        RECT 362.800 262.200 363.800 265.600 ;
        RECT 363.000 261.600 363.800 262.200 ;
        RECT 369.000 261.600 370.000 265.600 ;
        RECT 375.600 261.600 376.400 265.400 ;
        RECT 380.400 261.600 381.200 264.200 ;
        RECT 382.000 261.600 382.800 268.200 ;
        RECT 389.000 261.600 389.800 266.200 ;
        RECT 393.200 261.600 394.000 264.200 ;
        RECT 396.400 261.600 397.200 264.200 ;
        RECT 401.200 261.600 402.000 266.200 ;
        RECT 402.800 261.600 403.600 264.200 ;
        RECT 406.000 261.600 406.800 264.200 ;
        RECT 407.600 261.600 408.400 264.200 ;
        RECT 412.400 261.600 413.200 264.200 ;
        RECT 415.600 261.600 416.400 266.000 ;
        RECT 421.200 261.600 422.000 264.200 ;
        RECT 424.400 261.600 425.400 264.200 ;
        RECT 430.000 261.600 430.800 266.200 ;
        RECT 433.200 261.600 434.000 264.200 ;
        RECT 436.400 261.600 437.200 264.200 ;
        RECT 441.200 261.600 442.000 265.400 ;
        RECT 450.800 262.200 451.800 265.600 ;
        RECT 451.000 261.600 451.800 262.200 ;
        RECT 457.000 261.600 458.000 265.600 ;
        RECT 460.400 261.600 461.200 266.200 ;
        RECT 466.800 261.600 467.600 266.200 ;
        RECT 472.200 261.600 473.200 264.200 ;
        RECT 475.600 261.600 476.400 264.200 ;
        RECT 481.200 261.600 482.000 266.000 ;
        RECT 486.000 261.600 486.800 266.200 ;
        RECT 491.400 261.600 492.400 264.200 ;
        RECT 494.800 261.600 495.600 264.200 ;
        RECT 500.400 261.600 501.200 266.000 ;
        RECT 505.200 261.600 506.000 266.200 ;
        RECT 510.600 261.600 511.600 264.200 ;
        RECT 514.000 261.600 514.800 264.200 ;
        RECT 519.600 261.600 520.400 266.000 ;
        RECT 524.400 261.600 525.200 266.200 ;
        RECT 529.800 261.600 530.800 264.200 ;
        RECT 533.200 261.600 534.000 264.200 ;
        RECT 538.800 261.600 539.600 266.000 ;
        RECT 543.600 261.600 544.400 266.200 ;
        RECT 549.000 261.600 550.000 264.200 ;
        RECT 552.400 261.600 553.200 264.200 ;
        RECT 558.000 261.600 558.800 266.000 ;
        RECT 562.800 261.600 563.600 266.200 ;
        RECT 568.200 261.600 569.200 264.200 ;
        RECT 571.600 261.600 572.400 264.200 ;
        RECT 577.200 261.600 578.000 266.000 ;
        RECT 582.000 261.600 582.800 266.200 ;
        RECT 0.400 260.400 586.800 261.600 ;
        RECT 2.800 256.600 3.600 260.400 ;
        RECT 10.800 255.800 11.600 260.400 ;
        RECT 12.400 255.800 13.200 260.400 ;
        RECT 15.600 257.800 16.400 260.400 ;
        RECT 19.400 255.800 20.200 260.400 ;
        RECT 23.600 257.800 24.400 260.400 ;
        RECT 26.800 255.400 27.600 260.400 ;
        RECT 32.000 255.000 32.800 260.400 ;
        RECT 38.000 256.600 38.800 260.400 ;
        RECT 44.400 255.800 45.200 260.400 ;
        RECT 46.000 257.800 46.800 260.400 ;
        RECT 49.200 257.800 50.000 260.400 ;
        RECT 52.400 256.400 53.400 260.400 ;
        RECT 58.600 259.800 59.400 260.400 ;
        RECT 63.800 259.800 64.600 260.400 ;
        RECT 58.600 256.400 59.600 259.800 ;
        RECT 63.600 256.400 64.600 259.800 ;
        RECT 69.800 256.400 70.800 260.400 ;
        RECT 73.800 255.800 74.600 260.400 ;
        RECT 78.000 257.800 78.800 260.400 ;
        RECT 81.200 257.800 82.000 260.400 ;
        RECT 84.400 256.600 85.200 260.400 ;
        RECT 90.800 257.800 91.600 260.400 ;
        RECT 94.000 257.800 94.800 260.400 ;
        RECT 95.600 253.800 96.400 260.400 ;
        RECT 103.600 256.600 104.400 260.400 ;
        RECT 110.000 257.800 110.800 260.400 ;
        RECT 111.600 257.800 112.400 260.400 ;
        RECT 114.800 257.800 115.600 260.400 ;
        RECT 119.600 256.600 120.400 260.400 ;
        RECT 122.800 257.800 123.600 260.400 ;
        RECT 126.000 257.800 126.800 260.400 ;
        RECT 129.400 259.800 130.200 260.400 ;
        RECT 129.200 256.400 130.200 259.800 ;
        RECT 135.400 256.400 136.400 260.400 ;
        RECT 145.400 259.800 146.200 260.400 ;
        RECT 145.200 256.400 146.200 259.800 ;
        RECT 151.400 256.400 152.400 260.400 ;
        RECT 154.800 255.800 155.600 260.400 ;
        RECT 161.200 256.600 162.000 260.400 ;
        RECT 169.200 255.800 170.000 260.400 ;
        RECT 174.000 256.600 174.800 260.400 ;
        RECT 177.200 257.800 178.000 260.400 ;
        RECT 180.400 257.800 181.200 260.400 ;
        RECT 185.200 256.600 186.000 260.400 ;
        RECT 190.000 257.800 190.800 260.400 ;
        RECT 193.200 257.800 194.000 260.400 ;
        RECT 194.800 257.800 195.600 260.400 ;
        RECT 198.000 257.800 198.800 260.400 ;
        RECT 201.200 256.000 202.000 260.400 ;
        RECT 206.800 257.800 207.600 260.400 ;
        RECT 210.000 257.800 211.000 260.400 ;
        RECT 215.600 255.800 216.400 260.400 ;
        RECT 220.400 256.000 221.200 260.400 ;
        RECT 226.000 257.800 226.800 260.400 ;
        RECT 229.200 257.800 230.200 260.400 ;
        RECT 234.800 255.800 235.600 260.400 ;
        RECT 239.600 255.800 240.400 260.400 ;
        RECT 244.400 256.000 245.200 260.400 ;
        RECT 250.000 257.800 250.800 260.400 ;
        RECT 253.200 257.800 254.200 260.400 ;
        RECT 258.800 255.800 259.600 260.400 ;
        RECT 263.600 256.000 264.400 260.400 ;
        RECT 269.200 257.800 270.000 260.400 ;
        RECT 272.400 257.800 273.400 260.400 ;
        RECT 278.000 255.800 278.800 260.400 ;
        RECT 282.800 255.800 283.600 260.400 ;
        RECT 292.400 256.000 293.200 260.400 ;
        RECT 298.000 257.800 298.800 260.400 ;
        RECT 301.200 257.800 302.200 260.400 ;
        RECT 306.800 255.800 307.600 260.400 ;
        RECT 311.800 259.800 312.600 260.400 ;
        RECT 311.600 256.400 312.600 259.800 ;
        RECT 317.800 256.400 318.800 260.400 ;
        RECT 324.400 256.600 325.200 260.400 ;
        RECT 327.600 255.800 328.400 260.400 ;
        RECT 334.000 256.600 334.800 260.400 ;
        RECT 340.400 257.800 341.200 260.400 ;
        RECT 343.600 257.800 344.400 260.400 ;
        RECT 348.400 255.800 349.200 260.400 ;
        RECT 350.000 257.800 350.800 260.400 ;
        RECT 353.200 257.800 354.000 260.400 ;
        RECT 356.400 257.800 357.200 260.400 ;
        RECT 361.200 256.600 362.000 260.400 ;
        RECT 366.000 257.800 366.800 260.400 ;
        RECT 369.200 256.000 370.000 260.400 ;
        RECT 374.800 257.800 375.600 260.400 ;
        RECT 378.000 257.800 379.000 260.400 ;
        RECT 383.600 255.800 384.400 260.400 ;
        RECT 387.200 255.800 388.000 260.400 ;
        RECT 393.200 255.800 394.000 260.400 ;
        RECT 394.800 257.800 395.600 260.400 ;
        RECT 398.000 257.800 398.800 260.400 ;
        RECT 401.200 256.000 402.000 260.400 ;
        RECT 406.800 257.800 407.600 260.400 ;
        RECT 410.000 257.800 411.000 260.400 ;
        RECT 415.600 255.800 416.400 260.400 ;
        RECT 420.400 256.000 421.200 260.400 ;
        RECT 426.000 257.800 426.800 260.400 ;
        RECT 429.200 257.800 430.200 260.400 ;
        RECT 434.800 255.800 435.600 260.400 ;
        RECT 438.600 255.800 439.400 260.400 ;
        RECT 442.800 257.800 443.600 260.400 ;
        RECT 454.000 253.800 454.800 260.400 ;
        RECT 455.600 257.800 456.400 260.400 ;
        RECT 458.800 257.800 459.600 260.400 ;
        RECT 460.800 255.800 461.600 260.400 ;
        RECT 466.800 255.800 467.600 260.400 ;
        RECT 468.400 257.800 469.200 260.400 ;
        RECT 474.800 256.600 475.600 260.400 ;
        RECT 481.200 255.800 482.000 260.400 ;
        RECT 486.000 256.600 486.800 260.400 ;
        RECT 492.400 255.800 493.200 260.400 ;
        RECT 494.000 257.800 494.800 260.400 ;
        RECT 497.200 257.800 498.000 260.400 ;
        RECT 498.800 257.800 499.600 260.400 ;
        RECT 502.000 257.800 502.800 260.400 ;
        RECT 505.200 256.400 506.200 260.400 ;
        RECT 511.400 259.800 512.200 260.400 ;
        RECT 516.600 259.800 517.400 260.400 ;
        RECT 511.400 256.400 512.400 259.800 ;
        RECT 516.400 256.400 517.400 259.800 ;
        RECT 522.600 256.400 523.600 260.400 ;
        RECT 527.600 256.400 528.600 260.400 ;
        RECT 533.800 259.800 534.600 260.400 ;
        RECT 533.800 256.400 534.800 259.800 ;
        RECT 538.800 255.800 539.600 260.400 ;
        RECT 544.200 257.800 545.200 260.400 ;
        RECT 547.600 257.800 548.400 260.400 ;
        RECT 553.200 256.000 554.000 260.400 ;
        RECT 558.000 255.800 558.800 260.400 ;
        RECT 562.800 255.800 563.600 260.400 ;
        RECT 568.200 257.800 569.200 260.400 ;
        RECT 571.600 257.800 572.400 260.400 ;
        RECT 577.200 256.000 578.000 260.400 ;
        RECT 582.000 255.800 582.800 260.400 ;
        RECT 2.800 221.600 3.600 226.000 ;
        RECT 8.400 221.600 9.200 224.200 ;
        RECT 11.600 221.600 12.600 224.200 ;
        RECT 17.200 221.600 18.000 226.200 ;
        RECT 22.000 221.600 23.000 225.600 ;
        RECT 28.200 222.200 29.200 225.600 ;
        RECT 28.200 221.600 29.000 222.200 ;
        RECT 33.200 221.600 34.200 225.600 ;
        RECT 39.400 222.200 40.400 225.600 ;
        RECT 39.400 221.600 40.200 222.200 ;
        RECT 44.400 221.600 45.200 226.000 ;
        RECT 50.000 221.600 50.800 224.200 ;
        RECT 53.200 221.600 54.200 224.200 ;
        RECT 58.800 221.600 59.600 226.200 ;
        RECT 63.600 221.600 64.400 226.200 ;
        RECT 69.000 221.600 70.000 224.200 ;
        RECT 72.400 221.600 73.200 224.200 ;
        RECT 78.000 221.600 78.800 226.000 ;
        RECT 82.800 222.200 83.800 225.600 ;
        RECT 83.000 221.600 83.800 222.200 ;
        RECT 89.000 221.600 90.000 225.600 ;
        RECT 95.600 221.600 96.400 226.200 ;
        RECT 98.800 221.600 99.600 226.000 ;
        RECT 104.400 221.600 105.200 224.200 ;
        RECT 107.600 221.600 108.600 224.200 ;
        RECT 113.200 221.600 114.000 226.200 ;
        RECT 118.000 221.600 118.800 226.000 ;
        RECT 123.600 221.600 124.400 224.200 ;
        RECT 126.800 221.600 127.800 224.200 ;
        RECT 132.400 221.600 133.200 226.200 ;
        RECT 142.000 222.200 143.000 225.600 ;
        RECT 142.200 221.600 143.000 222.200 ;
        RECT 148.200 221.600 149.200 225.600 ;
        RECT 153.200 221.600 154.000 225.400 ;
        RECT 159.600 221.600 160.400 225.400 ;
        RECT 166.000 221.600 166.800 226.000 ;
        RECT 171.600 221.600 172.400 224.200 ;
        RECT 174.800 221.600 175.800 224.200 ;
        RECT 180.400 221.600 181.200 226.200 ;
        RECT 183.600 221.600 184.400 226.200 ;
        RECT 186.800 221.600 187.600 226.200 ;
        RECT 190.000 221.600 190.800 226.200 ;
        RECT 193.200 221.600 194.000 226.200 ;
        RECT 196.400 221.600 197.200 226.200 ;
        RECT 199.600 221.600 200.400 226.000 ;
        RECT 205.200 221.600 206.000 224.200 ;
        RECT 208.400 221.600 209.400 224.200 ;
        RECT 214.000 221.600 214.800 226.200 ;
        RECT 218.800 221.600 219.600 226.000 ;
        RECT 224.400 221.600 225.200 224.200 ;
        RECT 227.600 221.600 228.600 224.200 ;
        RECT 233.200 221.600 234.000 226.200 ;
        RECT 236.400 221.600 237.200 224.200 ;
        RECT 241.200 221.600 242.000 226.200 ;
        RECT 246.000 221.600 246.800 226.200 ;
        RECT 251.400 221.600 252.400 224.200 ;
        RECT 254.800 221.600 255.600 224.200 ;
        RECT 260.400 221.600 261.200 226.000 ;
        RECT 265.200 221.600 266.000 226.200 ;
        RECT 270.600 221.600 271.600 224.200 ;
        RECT 274.000 221.600 274.800 224.200 ;
        RECT 279.600 221.600 280.400 226.000 ;
        RECT 282.800 221.600 283.600 224.200 ;
        RECT 286.000 221.600 286.800 226.200 ;
        RECT 295.600 221.600 296.400 224.200 ;
        RECT 298.800 221.600 299.600 224.200 ;
        RECT 302.000 221.600 302.800 224.200 ;
        RECT 303.600 221.600 304.400 224.200 ;
        RECT 306.800 221.600 307.600 224.200 ;
        RECT 310.000 221.600 310.800 226.200 ;
        RECT 315.400 221.600 316.400 224.200 ;
        RECT 318.800 221.600 319.600 224.200 ;
        RECT 324.400 221.600 325.200 226.000 ;
        RECT 330.800 221.600 331.600 226.200 ;
        RECT 332.400 221.600 333.200 224.200 ;
        RECT 335.600 221.600 336.400 226.200 ;
        RECT 342.000 221.600 342.800 226.200 ;
        RECT 347.400 221.600 348.400 224.200 ;
        RECT 350.800 221.600 351.600 224.200 ;
        RECT 356.400 221.600 357.200 226.000 ;
        RECT 361.200 221.600 362.000 226.200 ;
        RECT 366.000 221.600 366.800 226.000 ;
        RECT 371.600 221.600 372.400 224.200 ;
        RECT 374.800 221.600 375.800 224.200 ;
        RECT 380.400 221.600 381.200 226.200 ;
        RECT 385.200 221.600 386.000 226.200 ;
        RECT 390.600 221.600 391.600 224.200 ;
        RECT 394.000 221.600 394.800 224.200 ;
        RECT 399.600 221.600 400.400 226.000 ;
        RECT 404.400 221.600 405.200 226.200 ;
        RECT 409.800 221.600 410.800 224.200 ;
        RECT 413.200 221.600 414.000 224.200 ;
        RECT 418.800 221.600 419.600 226.000 ;
        RECT 422.000 221.600 422.800 226.200 ;
        RECT 426.800 221.600 427.600 224.200 ;
        RECT 430.000 221.600 430.800 224.200 ;
        RECT 431.600 221.600 432.400 224.200 ;
        RECT 434.800 221.600 435.600 224.200 ;
        RECT 436.400 221.600 437.200 224.200 ;
        RECT 444.400 221.600 445.200 228.200 ;
        RECT 452.400 221.600 453.200 224.200 ;
        RECT 454.000 221.600 454.800 224.200 ;
        RECT 457.200 221.600 458.000 224.200 ;
        RECT 462.000 221.600 462.800 226.200 ;
        RECT 463.600 221.600 464.400 226.200 ;
        RECT 473.200 221.600 474.000 225.400 ;
        RECT 476.400 221.600 477.200 224.200 ;
        RECT 481.200 221.600 482.200 225.600 ;
        RECT 487.400 222.200 488.400 225.600 ;
        RECT 487.400 221.600 488.200 222.200 ;
        RECT 492.400 221.600 493.200 226.200 ;
        RECT 497.800 221.600 498.800 224.200 ;
        RECT 501.200 221.600 502.000 224.200 ;
        RECT 506.800 221.600 507.600 226.000 ;
        RECT 511.600 221.600 512.400 226.200 ;
        RECT 517.000 221.600 518.000 224.200 ;
        RECT 520.400 221.600 521.200 224.200 ;
        RECT 526.000 221.600 526.800 226.000 ;
        RECT 530.800 221.600 531.600 226.200 ;
        RECT 535.600 221.600 536.400 226.200 ;
        RECT 541.000 221.600 542.000 224.200 ;
        RECT 544.400 221.600 545.200 224.200 ;
        RECT 550.000 221.600 550.800 226.000 ;
        RECT 554.800 221.600 555.600 226.200 ;
        RECT 560.200 221.600 561.200 224.200 ;
        RECT 563.600 221.600 564.400 224.200 ;
        RECT 569.200 221.600 570.000 226.000 ;
        RECT 574.000 221.600 574.800 226.200 ;
        RECT 578.800 221.600 579.600 226.200 ;
        RECT 0.400 220.400 586.800 221.600 ;
        RECT 2.800 215.800 3.600 220.400 ;
        RECT 8.200 217.800 9.200 220.400 ;
        RECT 11.600 217.800 12.400 220.400 ;
        RECT 17.200 216.000 18.000 220.400 ;
        RECT 22.000 215.800 22.800 220.400 ;
        RECT 27.400 217.800 28.400 220.400 ;
        RECT 30.800 217.800 31.600 220.400 ;
        RECT 36.400 216.000 37.200 220.400 ;
        RECT 41.200 216.000 42.000 220.400 ;
        RECT 46.800 217.800 47.600 220.400 ;
        RECT 50.000 217.800 51.000 220.400 ;
        RECT 55.600 215.800 56.400 220.400 ;
        RECT 60.400 215.800 61.200 220.400 ;
        RECT 65.800 217.800 66.800 220.400 ;
        RECT 69.200 217.800 70.000 220.400 ;
        RECT 74.800 216.000 75.600 220.400 ;
        RECT 79.600 216.000 80.400 220.400 ;
        RECT 85.200 217.800 86.000 220.400 ;
        RECT 88.400 217.800 89.400 220.400 ;
        RECT 94.000 215.800 94.800 220.400 ;
        RECT 97.200 215.800 98.000 220.400 ;
        RECT 100.400 215.800 101.200 220.400 ;
        RECT 103.600 215.800 104.400 220.400 ;
        RECT 106.800 215.800 107.600 220.400 ;
        RECT 110.000 215.800 110.800 220.400 ;
        RECT 113.200 216.000 114.000 220.400 ;
        RECT 118.800 217.800 119.600 220.400 ;
        RECT 122.000 217.800 123.000 220.400 ;
        RECT 127.600 215.800 128.400 220.400 ;
        RECT 137.200 215.800 138.000 220.400 ;
        RECT 142.600 217.800 143.600 220.400 ;
        RECT 146.000 217.800 146.800 220.400 ;
        RECT 151.600 216.000 152.400 220.400 ;
        RECT 156.400 215.800 157.200 220.400 ;
        RECT 161.800 217.800 162.800 220.400 ;
        RECT 165.200 217.800 166.000 220.400 ;
        RECT 170.800 216.000 171.600 220.400 ;
        RECT 174.000 217.800 174.800 220.400 ;
        RECT 177.200 217.800 178.000 220.400 ;
        RECT 180.400 217.800 181.200 220.400 ;
        RECT 183.600 216.600 184.400 220.400 ;
        RECT 188.400 217.800 189.200 220.400 ;
        RECT 191.600 217.800 192.400 220.400 ;
        RECT 193.200 217.800 194.000 220.400 ;
        RECT 198.000 216.600 198.800 220.400 ;
        RECT 204.400 215.800 205.200 220.400 ;
        RECT 209.800 217.800 210.800 220.400 ;
        RECT 213.200 217.800 214.000 220.400 ;
        RECT 218.800 216.000 219.600 220.400 ;
        RECT 222.000 217.800 222.800 220.400 ;
        RECT 225.200 217.800 226.000 220.400 ;
        RECT 226.800 217.800 227.600 220.400 ;
        RECT 230.000 217.800 230.800 220.400 ;
        RECT 233.200 217.800 234.000 220.400 ;
        RECT 236.400 216.600 237.200 220.400 ;
        RECT 242.800 216.600 243.600 220.400 ;
        RECT 249.200 216.600 250.000 220.400 ;
        RECT 255.600 215.800 256.400 220.400 ;
        RECT 261.000 217.800 262.000 220.400 ;
        RECT 264.400 217.800 265.200 220.400 ;
        RECT 270.000 216.000 270.800 220.400 ;
        RECT 273.200 217.800 274.000 220.400 ;
        RECT 276.400 217.800 277.200 220.400 ;
        RECT 279.600 217.800 280.400 220.400 ;
        RECT 281.200 215.800 282.000 220.400 ;
        RECT 287.600 217.800 288.400 220.400 ;
        RECT 294.000 217.800 294.800 220.400 ;
        RECT 297.200 217.800 298.000 220.400 ;
        RECT 300.400 216.000 301.200 220.400 ;
        RECT 306.000 217.800 306.800 220.400 ;
        RECT 309.200 217.800 310.200 220.400 ;
        RECT 314.800 215.800 315.600 220.400 ;
        RECT 319.600 215.800 320.400 220.400 ;
        RECT 324.400 216.000 325.200 220.400 ;
        RECT 330.000 217.800 330.800 220.400 ;
        RECT 333.200 217.800 334.200 220.400 ;
        RECT 338.800 215.800 339.600 220.400 ;
        RECT 343.600 215.800 344.400 220.400 ;
        RECT 348.400 215.800 349.200 220.400 ;
        RECT 353.800 217.800 354.800 220.400 ;
        RECT 357.200 217.800 358.000 220.400 ;
        RECT 362.800 216.000 363.600 220.400 ;
        RECT 366.000 217.800 366.800 220.400 ;
        RECT 370.800 216.600 371.600 220.400 ;
        RECT 377.200 216.600 378.000 220.400 ;
        RECT 383.800 219.800 384.600 220.400 ;
        RECT 383.600 216.400 384.600 219.800 ;
        RECT 389.800 216.400 390.800 220.400 ;
        RECT 393.200 217.800 394.000 220.400 ;
        RECT 399.600 216.600 400.400 220.400 ;
        RECT 404.400 216.400 405.400 220.400 ;
        RECT 410.600 219.800 411.400 220.400 ;
        RECT 410.600 216.400 411.600 219.800 ;
        RECT 415.600 215.800 416.400 220.400 ;
        RECT 421.000 217.800 422.000 220.400 ;
        RECT 424.400 217.800 425.200 220.400 ;
        RECT 430.000 216.000 430.800 220.400 ;
        RECT 434.800 216.200 435.600 220.400 ;
        RECT 438.000 217.800 438.800 220.400 ;
        RECT 439.600 217.800 440.400 220.400 ;
        RECT 442.800 217.800 443.600 220.400 ;
        RECT 449.200 215.800 450.000 220.400 ;
        RECT 454.000 217.800 454.800 220.400 ;
        RECT 457.200 217.800 458.000 220.400 ;
        RECT 460.400 216.600 461.200 220.400 ;
        RECT 468.400 215.800 469.200 220.400 ;
        RECT 471.600 216.600 472.400 220.400 ;
        RECT 478.000 216.600 478.800 220.400 ;
        RECT 482.800 215.800 483.600 220.400 ;
        RECT 487.600 217.800 488.400 220.400 ;
        RECT 492.400 216.600 493.200 220.400 ;
        RECT 498.800 215.800 499.600 220.400 ;
        RECT 505.400 219.800 506.200 220.400 ;
        RECT 505.200 216.400 506.200 219.800 ;
        RECT 511.400 216.400 512.400 220.400 ;
        RECT 516.400 216.400 517.400 220.400 ;
        RECT 522.600 219.800 523.400 220.400 ;
        RECT 522.600 216.400 523.600 219.800 ;
        RECT 526.400 215.800 527.200 220.400 ;
        RECT 532.400 215.800 533.200 220.400 ;
        RECT 537.200 215.800 538.000 220.400 ;
        RECT 538.800 215.800 539.600 220.400 ;
        RECT 545.200 215.800 546.000 220.400 ;
        RECT 550.600 217.800 551.600 220.400 ;
        RECT 554.000 217.800 554.800 220.400 ;
        RECT 559.600 216.000 560.400 220.400 ;
        RECT 564.400 215.800 565.200 220.400 ;
        RECT 569.800 217.800 570.800 220.400 ;
        RECT 573.200 217.800 574.000 220.400 ;
        RECT 578.800 216.000 579.600 220.400 ;
        RECT 583.600 215.800 584.400 220.400 ;
        RECT 2.800 181.600 3.600 186.200 ;
        RECT 8.200 181.600 9.200 184.200 ;
        RECT 11.600 181.600 12.400 184.200 ;
        RECT 17.200 181.600 18.000 186.000 ;
        RECT 22.000 181.600 22.800 186.200 ;
        RECT 27.400 181.600 28.400 184.200 ;
        RECT 30.800 181.600 31.600 184.200 ;
        RECT 36.400 181.600 37.200 186.000 ;
        RECT 42.800 181.600 43.600 186.200 ;
        RECT 44.400 181.600 45.200 184.200 ;
        RECT 47.600 181.600 48.400 185.800 ;
        RECT 50.800 181.600 51.600 184.200 ;
        RECT 54.000 181.600 54.800 184.200 ;
        RECT 58.800 181.600 59.600 186.200 ;
        RECT 63.600 181.600 64.400 186.200 ;
        RECT 68.400 181.600 69.200 185.400 ;
        RECT 74.200 181.600 75.000 186.000 ;
        RECT 78.000 181.600 78.800 184.200 ;
        RECT 84.400 181.600 85.200 186.200 ;
        RECT 87.600 181.600 88.400 184.200 ;
        RECT 92.400 181.600 93.200 186.200 ;
        RECT 94.000 181.600 94.800 184.200 ;
        RECT 98.800 181.600 99.600 185.400 ;
        RECT 106.800 181.600 107.600 185.400 ;
        RECT 113.200 181.600 114.000 186.200 ;
        RECT 114.800 181.600 115.600 184.200 ;
        RECT 121.200 181.600 122.000 186.200 ;
        RECT 124.400 181.600 125.200 186.200 ;
        RECT 129.800 181.600 130.800 184.200 ;
        RECT 133.200 181.600 134.000 184.200 ;
        RECT 138.800 181.600 139.600 186.000 ;
        RECT 148.400 181.600 149.200 186.200 ;
        RECT 153.800 181.600 154.800 184.200 ;
        RECT 157.200 181.600 158.000 184.200 ;
        RECT 162.800 181.600 163.600 186.000 ;
        RECT 167.600 181.600 168.400 186.200 ;
        RECT 173.000 181.600 174.000 184.200 ;
        RECT 176.400 181.600 177.200 184.200 ;
        RECT 182.000 181.600 182.800 186.000 ;
        RECT 185.200 181.600 186.000 184.200 ;
        RECT 191.600 181.600 192.400 185.400 ;
        RECT 198.000 181.600 198.800 186.200 ;
        RECT 202.800 181.600 203.600 185.400 ;
        RECT 209.200 181.600 210.000 186.200 ;
        RECT 212.400 181.600 213.200 184.200 ;
        RECT 215.600 181.600 216.600 185.600 ;
        RECT 221.800 182.200 222.800 185.600 ;
        RECT 221.800 181.600 222.600 182.200 ;
        RECT 226.800 181.600 227.600 186.200 ;
        RECT 232.200 181.600 233.200 184.200 ;
        RECT 235.600 181.600 236.400 184.200 ;
        RECT 241.200 181.600 242.000 186.000 ;
        RECT 247.600 181.600 248.400 185.400 ;
        RECT 250.800 181.600 251.600 184.200 ;
        RECT 254.000 181.600 254.800 184.200 ;
        RECT 257.200 181.600 258.000 184.200 ;
        RECT 260.400 182.200 261.400 185.600 ;
        RECT 260.600 181.600 261.400 182.200 ;
        RECT 266.600 181.600 267.600 185.600 ;
        RECT 270.000 181.600 270.800 186.200 ;
        RECT 276.400 181.600 277.200 186.200 ;
        RECT 281.800 181.600 282.800 184.200 ;
        RECT 285.200 181.600 286.000 184.200 ;
        RECT 290.800 181.600 291.600 186.000 ;
        RECT 298.800 181.600 299.600 186.200 ;
        RECT 306.800 181.600 307.600 186.200 ;
        RECT 310.000 181.600 310.800 186.200 ;
        RECT 314.800 181.600 315.600 185.400 ;
        RECT 318.000 181.600 318.800 186.200 ;
        RECT 324.400 182.200 325.400 185.600 ;
        RECT 324.600 181.600 325.400 182.200 ;
        RECT 330.600 181.600 331.600 185.600 ;
        RECT 335.600 181.600 336.400 185.400 ;
        RECT 340.400 181.600 341.200 186.200 ;
        RECT 346.800 181.600 347.800 185.600 ;
        RECT 353.000 182.200 354.000 185.600 ;
        RECT 353.000 181.600 353.800 182.200 ;
        RECT 358.000 181.600 358.800 186.200 ;
        RECT 363.400 181.600 364.400 184.200 ;
        RECT 366.800 181.600 367.600 184.200 ;
        RECT 372.400 181.600 373.200 186.000 ;
        RECT 377.200 181.600 378.000 186.600 ;
        RECT 382.400 181.600 383.200 187.000 ;
        RECT 388.400 181.600 389.200 185.400 ;
        RECT 391.600 181.600 392.400 184.200 ;
        RECT 394.800 181.600 395.600 184.200 ;
        RECT 396.400 181.600 397.200 184.200 ;
        RECT 399.600 181.600 400.400 184.200 ;
        RECT 401.200 181.600 402.000 184.200 ;
        RECT 404.400 181.600 405.200 184.200 ;
        RECT 407.600 181.600 408.400 184.200 ;
        RECT 410.800 181.600 411.600 186.000 ;
        RECT 416.400 181.600 417.200 184.200 ;
        RECT 419.600 181.600 420.600 184.200 ;
        RECT 425.200 181.600 426.000 186.200 ;
        RECT 430.000 181.600 430.800 186.200 ;
        RECT 435.400 181.600 436.400 184.200 ;
        RECT 438.800 181.600 439.600 184.200 ;
        RECT 444.400 181.600 445.200 186.000 ;
        RECT 453.000 181.600 453.800 186.200 ;
        RECT 457.200 181.600 458.000 184.200 ;
        RECT 462.000 181.600 462.800 185.400 ;
        RECT 466.800 182.200 467.800 185.600 ;
        RECT 467.000 181.600 467.800 182.200 ;
        RECT 473.000 181.600 474.000 185.600 ;
        RECT 478.000 181.600 478.800 185.400 ;
        RECT 484.400 181.600 485.200 184.200 ;
        RECT 487.600 181.600 488.400 185.400 ;
        RECT 493.000 181.600 493.800 186.200 ;
        RECT 497.200 181.600 498.000 184.200 ;
        RECT 500.400 181.600 501.400 185.600 ;
        RECT 506.600 182.200 507.600 185.600 ;
        RECT 506.600 181.600 507.400 182.200 ;
        RECT 510.000 181.600 510.800 184.200 ;
        RECT 513.200 181.600 514.000 184.200 ;
        RECT 516.400 181.600 517.200 184.200 ;
        RECT 521.200 181.600 522.000 186.200 ;
        RECT 522.800 181.600 523.600 186.200 ;
        RECT 526.000 181.600 526.800 186.200 ;
        RECT 530.800 181.600 531.600 186.200 ;
        RECT 532.400 181.600 533.200 184.200 ;
        RECT 535.600 181.600 536.400 186.200 ;
        RECT 542.000 181.600 542.800 186.200 ;
        RECT 545.200 181.600 546.000 185.400 ;
        RECT 550.000 181.600 550.800 184.200 ;
        RECT 553.200 181.600 554.000 184.200 ;
        RECT 556.400 181.600 557.400 185.600 ;
        RECT 562.600 182.200 563.600 185.600 ;
        RECT 562.600 181.600 563.400 182.200 ;
        RECT 567.600 181.600 568.400 186.200 ;
        RECT 573.000 181.600 574.000 184.200 ;
        RECT 576.400 181.600 577.200 184.200 ;
        RECT 582.000 181.600 582.800 186.000 ;
        RECT 0.400 180.400 586.800 181.600 ;
        RECT 2.800 176.000 3.600 180.400 ;
        RECT 8.400 177.800 9.200 180.400 ;
        RECT 11.600 177.800 12.600 180.400 ;
        RECT 17.200 175.800 18.000 180.400 ;
        RECT 23.600 176.600 24.400 180.400 ;
        RECT 28.400 176.400 29.400 180.400 ;
        RECT 34.600 179.800 35.400 180.400 ;
        RECT 34.600 176.400 35.600 179.800 ;
        RECT 39.600 176.400 40.600 180.400 ;
        RECT 45.800 179.800 46.600 180.400 ;
        RECT 45.800 176.400 46.800 179.800 ;
        RECT 52.400 176.600 53.200 180.400 ;
        RECT 55.600 177.800 56.400 180.400 ;
        RECT 59.800 175.800 60.600 180.400 ;
        RECT 65.200 176.600 66.000 180.400 ;
        RECT 70.000 177.800 70.800 180.400 ;
        RECT 71.600 177.800 72.400 180.400 ;
        RECT 74.800 177.800 75.600 180.400 ;
        RECT 78.000 176.600 78.800 180.400 ;
        RECT 84.400 176.400 85.400 180.400 ;
        RECT 90.600 179.800 91.400 180.400 ;
        RECT 95.800 179.800 96.600 180.400 ;
        RECT 90.600 176.400 91.600 179.800 ;
        RECT 95.600 176.400 96.600 179.800 ;
        RECT 101.800 176.400 102.800 180.400 ;
        RECT 106.800 175.800 107.600 180.400 ;
        RECT 112.200 177.800 113.200 180.400 ;
        RECT 115.600 177.800 116.400 180.400 ;
        RECT 121.200 176.000 122.000 180.400 ;
        RECT 124.400 175.800 125.200 180.400 ;
        RECT 135.600 175.800 136.400 180.400 ;
        RECT 141.000 177.800 142.000 180.400 ;
        RECT 144.400 177.800 145.200 180.400 ;
        RECT 150.000 176.000 150.800 180.400 ;
        RECT 154.800 175.800 155.600 180.400 ;
        RECT 160.200 177.800 161.200 180.400 ;
        RECT 163.600 177.800 164.400 180.400 ;
        RECT 169.200 176.000 170.000 180.400 ;
        RECT 174.000 176.400 175.000 180.400 ;
        RECT 180.200 179.800 181.000 180.400 ;
        RECT 180.200 176.400 181.200 179.800 ;
        RECT 185.200 176.600 186.000 180.400 ;
        RECT 190.000 175.800 190.800 180.400 ;
        RECT 196.400 176.600 197.200 180.400 ;
        RECT 201.200 177.800 202.000 180.400 ;
        RECT 205.400 175.800 206.200 180.400 ;
        RECT 209.200 177.800 210.000 180.400 ;
        RECT 212.400 176.600 213.200 180.400 ;
        RECT 220.400 176.600 221.200 180.400 ;
        RECT 223.600 175.800 224.400 180.400 ;
        RECT 228.400 175.800 229.200 180.400 ;
        RECT 234.800 175.800 235.600 180.400 ;
        RECT 240.200 177.800 241.200 180.400 ;
        RECT 243.600 177.800 244.400 180.400 ;
        RECT 249.200 176.000 250.000 180.400 ;
        RECT 252.400 175.800 253.200 180.400 ;
        RECT 255.600 175.800 256.400 180.400 ;
        RECT 258.800 175.800 259.600 180.400 ;
        RECT 262.000 175.800 262.800 180.400 ;
        RECT 265.200 175.800 266.000 180.400 ;
        RECT 268.400 175.800 269.200 180.400 ;
        RECT 273.800 177.800 274.800 180.400 ;
        RECT 277.200 177.800 278.000 180.400 ;
        RECT 282.800 176.000 283.600 180.400 ;
        RECT 292.400 175.800 293.200 180.400 ;
        RECT 297.800 177.800 298.800 180.400 ;
        RECT 301.200 177.800 302.000 180.400 ;
        RECT 306.800 176.000 307.600 180.400 ;
        RECT 313.200 175.800 314.000 180.400 ;
        RECT 316.400 176.600 317.200 180.400 ;
        RECT 321.200 175.800 322.000 180.400 ;
        RECT 329.200 176.600 330.000 180.400 ;
        RECT 335.600 176.600 336.400 180.400 ;
        RECT 340.400 177.800 341.200 180.400 ;
        RECT 343.600 176.600 344.400 180.400 ;
        RECT 348.400 175.800 349.200 180.400 ;
        RECT 353.200 177.800 354.000 180.400 ;
        RECT 356.400 177.800 357.200 180.400 ;
        RECT 358.000 177.800 358.800 180.400 ;
        RECT 361.200 177.800 362.000 180.400 ;
        RECT 364.400 177.800 365.200 180.400 ;
        RECT 366.000 177.800 366.800 180.400 ;
        RECT 369.200 177.800 370.000 180.400 ;
        RECT 370.800 177.800 371.600 180.400 ;
        RECT 375.000 175.800 375.800 180.400 ;
        RECT 377.200 177.800 378.000 180.400 ;
        RECT 380.400 177.800 381.200 180.400 ;
        RECT 382.000 175.800 382.800 180.400 ;
        RECT 388.400 176.600 389.200 180.400 ;
        RECT 393.200 177.800 394.000 180.400 ;
        RECT 396.400 175.800 397.200 180.400 ;
        RECT 404.400 176.600 405.200 180.400 ;
        RECT 409.200 177.800 410.000 180.400 ;
        RECT 412.400 176.600 413.200 180.400 ;
        RECT 420.400 175.800 421.200 180.400 ;
        RECT 423.600 175.800 424.400 180.400 ;
        RECT 429.000 177.800 430.000 180.400 ;
        RECT 432.400 177.800 433.200 180.400 ;
        RECT 438.000 176.000 438.800 180.400 ;
        RECT 447.800 179.800 448.600 180.400 ;
        RECT 447.600 176.400 448.600 179.800 ;
        RECT 453.800 176.400 454.800 180.400 ;
        RECT 458.800 175.800 459.600 180.400 ;
        RECT 464.200 177.800 465.200 180.400 ;
        RECT 467.600 177.800 468.400 180.400 ;
        RECT 473.200 176.000 474.000 180.400 ;
        RECT 478.000 175.800 478.800 180.400 ;
        RECT 481.400 179.800 482.200 180.400 ;
        RECT 481.200 176.400 482.200 179.800 ;
        RECT 487.400 176.400 488.400 180.400 ;
        RECT 490.800 175.800 491.600 180.400 ;
        RECT 495.600 176.600 496.400 180.400 ;
        RECT 503.600 176.600 504.400 180.400 ;
        RECT 506.800 175.800 507.600 180.400 ;
        RECT 511.600 175.800 512.400 180.400 ;
        RECT 517.600 175.800 518.400 180.400 ;
        RECT 522.800 176.600 523.600 180.400 ;
        RECT 526.000 177.800 526.800 180.400 ;
        RECT 529.200 177.800 530.000 180.400 ;
        RECT 534.000 175.800 534.800 180.400 ;
        RECT 540.400 173.800 541.200 180.400 ;
        RECT 542.000 177.800 542.800 180.400 ;
        RECT 545.200 177.800 546.000 180.400 ;
        RECT 546.800 173.800 547.600 180.400 ;
        RECT 553.200 177.800 554.000 180.400 ;
        RECT 556.400 177.800 557.200 180.400 ;
        RECT 559.600 175.800 560.400 180.400 ;
        RECT 565.000 177.800 566.000 180.400 ;
        RECT 568.400 177.800 569.200 180.400 ;
        RECT 574.000 176.000 574.800 180.400 ;
        RECT 578.800 175.800 579.600 180.400 ;
        RECT 3.800 141.600 4.600 146.000 ;
        RECT 7.600 141.600 8.400 144.200 ;
        RECT 10.800 141.600 11.600 145.800 ;
        RECT 15.600 141.600 16.400 145.400 ;
        RECT 20.400 141.600 21.200 144.200 ;
        RECT 24.600 141.600 25.400 146.200 ;
        RECT 26.800 141.600 27.600 144.200 ;
        RECT 31.000 141.600 31.800 146.200 ;
        RECT 36.400 141.600 37.200 145.400 ;
        RECT 41.200 141.600 42.000 145.400 ;
        RECT 46.000 141.600 46.800 146.200 ;
        RECT 50.800 141.600 51.600 146.200 ;
        RECT 57.200 141.600 58.000 145.400 ;
        RECT 63.600 141.600 64.400 145.400 ;
        RECT 70.000 141.600 71.000 145.600 ;
        RECT 76.200 142.200 77.200 145.600 ;
        RECT 76.200 141.600 77.000 142.200 ;
        RECT 80.000 141.600 80.800 146.200 ;
        RECT 86.000 141.600 86.800 146.200 ;
        RECT 88.000 141.600 88.800 146.200 ;
        RECT 94.000 141.600 94.800 146.200 ;
        RECT 97.200 141.600 98.000 144.200 ;
        RECT 98.800 141.600 99.600 144.200 ;
        RECT 102.000 141.600 102.800 144.200 ;
        RECT 106.800 141.600 107.600 146.200 ;
        RECT 110.000 141.600 110.800 144.200 ;
        RECT 113.200 141.600 114.200 145.600 ;
        RECT 119.400 142.200 120.400 145.600 ;
        RECT 119.400 141.600 120.200 142.200 ;
        RECT 123.400 141.600 124.200 146.200 ;
        RECT 127.600 141.600 128.400 144.200 ;
        RECT 129.600 141.600 130.400 146.200 ;
        RECT 135.600 141.600 136.400 146.200 ;
        RECT 143.600 141.600 144.600 145.600 ;
        RECT 149.800 142.200 150.800 145.600 ;
        RECT 149.800 141.600 150.600 142.200 ;
        RECT 154.800 141.600 155.600 146.200 ;
        RECT 160.200 141.600 161.200 144.200 ;
        RECT 163.600 141.600 164.400 144.200 ;
        RECT 169.200 141.600 170.000 146.000 ;
        RECT 172.400 141.600 173.200 146.200 ;
        RECT 175.600 141.600 176.400 146.200 ;
        RECT 178.800 141.600 179.600 146.200 ;
        RECT 182.000 141.600 182.800 146.200 ;
        RECT 185.200 141.600 186.000 146.200 ;
        RECT 188.400 142.200 189.400 145.600 ;
        RECT 188.600 141.600 189.400 142.200 ;
        RECT 194.600 141.600 195.600 145.600 ;
        RECT 199.600 142.200 200.600 145.600 ;
        RECT 199.800 141.600 200.600 142.200 ;
        RECT 205.800 141.600 206.800 145.600 ;
        RECT 212.400 141.600 213.200 146.200 ;
        RECT 215.600 141.600 216.600 145.600 ;
        RECT 221.800 142.200 222.800 145.600 ;
        RECT 221.800 141.600 222.600 142.200 ;
        RECT 225.200 141.600 226.000 144.200 ;
        RECT 228.400 141.600 229.200 144.200 ;
        RECT 231.600 141.600 232.400 144.200 ;
        RECT 234.800 141.600 235.800 145.600 ;
        RECT 241.000 142.200 242.000 145.600 ;
        RECT 241.000 141.600 241.800 142.200 ;
        RECT 244.400 141.600 245.200 144.200 ;
        RECT 247.600 141.600 248.400 145.800 ;
        RECT 254.000 141.600 254.800 146.200 ;
        RECT 258.800 141.600 259.600 146.200 ;
        RECT 260.400 141.600 261.200 144.200 ;
        RECT 263.600 141.600 264.400 144.200 ;
        RECT 267.800 141.600 268.600 146.000 ;
        RECT 274.800 141.600 275.600 145.400 ;
        RECT 279.600 141.600 280.600 145.600 ;
        RECT 285.800 142.200 286.800 145.600 ;
        RECT 285.800 141.600 286.600 142.200 ;
        RECT 295.600 141.600 296.400 146.200 ;
        RECT 301.000 141.600 302.000 144.200 ;
        RECT 304.400 141.600 305.200 144.200 ;
        RECT 310.000 141.600 310.800 146.000 ;
        RECT 314.800 141.600 315.600 146.200 ;
        RECT 320.200 141.600 321.200 144.200 ;
        RECT 323.600 141.600 324.400 144.200 ;
        RECT 329.200 141.600 330.000 146.000 ;
        RECT 332.400 141.600 333.200 146.200 ;
        RECT 335.600 141.600 336.400 146.200 ;
        RECT 338.800 141.600 339.600 146.200 ;
        RECT 342.000 141.600 342.800 146.200 ;
        RECT 345.200 141.600 346.000 146.200 ;
        RECT 348.400 141.600 349.200 145.400 ;
        RECT 356.400 141.600 357.200 145.400 ;
        RECT 361.200 141.600 362.000 144.200 ;
        RECT 364.400 141.600 365.200 145.400 ;
        RECT 370.800 141.600 371.600 145.400 ;
        RECT 377.200 141.600 378.000 145.400 ;
        RECT 385.200 141.600 386.000 145.400 ;
        RECT 391.600 141.600 392.400 145.400 ;
        RECT 394.800 141.600 395.600 144.200 ;
        RECT 398.000 141.600 398.800 146.200 ;
        RECT 404.000 141.600 404.800 146.200 ;
        RECT 406.400 141.600 407.200 146.200 ;
        RECT 412.400 141.600 413.200 146.200 ;
        RECT 415.600 141.600 416.400 146.600 ;
        RECT 420.800 141.600 421.600 147.000 ;
        RECT 424.200 141.600 425.000 146.200 ;
        RECT 428.400 141.600 429.200 144.200 ;
        RECT 431.600 141.600 432.400 144.200 ;
        RECT 433.200 141.600 434.000 144.200 ;
        RECT 439.600 141.600 440.400 145.400 ;
        RECT 449.200 141.600 450.000 144.200 ;
        RECT 451.400 141.600 452.200 146.200 ;
        RECT 455.600 141.600 456.400 144.200 ;
        RECT 458.800 141.600 459.600 145.400 ;
        RECT 466.800 141.600 467.600 146.200 ;
        RECT 470.000 141.600 470.800 146.200 ;
        RECT 475.400 141.600 476.400 144.200 ;
        RECT 478.800 141.600 479.600 144.200 ;
        RECT 484.400 141.600 485.200 146.000 ;
        RECT 487.600 141.600 488.400 146.200 ;
        RECT 490.800 141.600 491.600 146.200 ;
        RECT 494.000 141.600 494.800 146.200 ;
        RECT 497.200 141.600 498.000 146.200 ;
        RECT 500.400 141.600 501.200 146.200 ;
        RECT 505.200 141.600 506.000 146.200 ;
        RECT 506.800 141.600 507.600 146.200 ;
        RECT 512.800 141.600 513.600 146.200 ;
        RECT 516.400 141.600 517.200 145.400 ;
        RECT 521.200 141.600 522.000 146.200 ;
        RECT 527.600 141.600 528.400 145.400 ;
        RECT 532.400 141.600 533.200 144.200 ;
        RECT 535.600 141.600 536.400 144.200 ;
        RECT 542.000 141.600 542.800 148.200 ;
        RECT 543.600 141.600 544.400 146.200 ;
        RECT 548.400 141.600 549.200 144.200 ;
        RECT 551.600 141.600 552.400 144.200 ;
        RECT 554.800 142.200 555.800 145.600 ;
        RECT 555.000 141.600 555.800 142.200 ;
        RECT 561.000 141.600 562.000 145.600 ;
        RECT 566.000 141.600 566.800 146.200 ;
        RECT 571.400 141.600 572.400 144.200 ;
        RECT 574.800 141.600 575.600 144.200 ;
        RECT 580.400 141.600 581.200 146.000 ;
        RECT 0.400 140.400 586.800 141.600 ;
        RECT 1.200 137.800 2.000 140.400 ;
        RECT 4.400 137.800 5.200 140.400 ;
        RECT 7.600 137.800 8.400 140.400 ;
        RECT 10.800 136.600 11.600 140.400 ;
        RECT 15.600 137.800 16.400 140.400 ;
        RECT 18.800 137.800 19.600 140.400 ;
        RECT 20.400 137.800 21.200 140.400 ;
        RECT 23.600 137.800 24.400 140.400 ;
        RECT 25.200 137.800 26.000 140.400 ;
        RECT 28.400 137.800 29.200 140.400 ;
        RECT 30.000 137.800 30.800 140.400 ;
        RECT 33.200 137.800 34.000 140.400 ;
        RECT 34.800 137.800 35.600 140.400 ;
        RECT 38.000 135.800 38.800 140.400 ;
        RECT 46.000 135.800 46.800 140.400 ;
        RECT 47.600 135.800 48.400 140.400 ;
        RECT 54.000 136.600 54.800 140.400 ;
        RECT 58.800 135.800 59.600 140.400 ;
        RECT 65.200 135.800 66.000 140.400 ;
        RECT 68.000 135.000 68.800 140.400 ;
        RECT 73.200 135.400 74.000 140.400 ;
        RECT 78.000 136.600 78.800 140.400 ;
        RECT 86.000 136.600 86.800 140.400 ;
        RECT 90.800 137.800 91.600 140.400 ;
        RECT 94.000 136.600 94.800 140.400 ;
        RECT 102.000 136.600 102.800 140.400 ;
        RECT 108.400 135.800 109.200 140.400 ;
        RECT 113.200 136.600 114.000 140.400 ;
        RECT 116.400 135.800 117.200 140.400 ;
        RECT 124.400 136.600 125.200 140.400 ;
        RECT 130.800 135.800 131.600 140.400 ;
        RECT 138.800 136.400 139.800 140.400 ;
        RECT 145.000 139.800 145.800 140.400 ;
        RECT 150.200 139.800 151.000 140.400 ;
        RECT 145.000 136.400 146.000 139.800 ;
        RECT 150.000 136.400 151.000 139.800 ;
        RECT 156.200 136.400 157.200 140.400 ;
        RECT 161.200 135.800 162.000 140.400 ;
        RECT 166.600 137.800 167.600 140.400 ;
        RECT 170.000 137.800 170.800 140.400 ;
        RECT 175.600 136.000 176.400 140.400 ;
        RECT 178.800 135.800 179.600 140.400 ;
        RECT 183.600 135.800 184.400 140.400 ;
        RECT 188.400 137.800 189.200 140.400 ;
        RECT 193.200 136.600 194.000 140.400 ;
        RECT 198.000 135.800 198.800 140.400 ;
        RECT 202.800 137.800 203.600 140.400 ;
        RECT 206.000 137.800 206.800 140.400 ;
        RECT 210.800 136.600 211.600 140.400 ;
        RECT 215.600 136.600 216.400 140.400 ;
        RECT 223.600 136.600 224.400 140.400 ;
        RECT 228.400 136.600 229.200 140.400 ;
        RECT 234.800 136.600 235.600 140.400 ;
        RECT 240.800 135.000 241.600 140.400 ;
        RECT 246.000 135.400 246.800 140.400 ;
        RECT 249.800 135.800 250.600 140.400 ;
        RECT 254.000 137.800 254.800 140.400 ;
        RECT 255.600 137.800 256.400 140.400 ;
        RECT 258.800 137.800 259.600 140.400 ;
        RECT 260.400 137.800 261.200 140.400 ;
        RECT 265.200 136.600 266.000 140.400 ;
        RECT 271.600 136.600 272.400 140.400 ;
        RECT 279.600 135.800 280.400 140.400 ;
        RECT 281.200 137.800 282.000 140.400 ;
        RECT 286.000 136.600 286.800 140.400 ;
        RECT 297.200 136.400 298.200 140.400 ;
        RECT 303.400 139.800 304.200 140.400 ;
        RECT 303.400 136.400 304.400 139.800 ;
        RECT 308.400 135.800 309.200 140.400 ;
        RECT 313.800 137.800 314.800 140.400 ;
        RECT 317.200 137.800 318.000 140.400 ;
        RECT 322.800 136.000 323.600 140.400 ;
        RECT 327.600 136.400 328.600 140.400 ;
        RECT 333.800 139.800 334.600 140.400 ;
        RECT 333.800 136.400 334.800 139.800 ;
        RECT 338.800 136.400 339.800 140.400 ;
        RECT 345.000 139.800 345.800 140.400 ;
        RECT 350.200 139.800 351.000 140.400 ;
        RECT 345.000 136.400 346.000 139.800 ;
        RECT 350.000 136.400 351.000 139.800 ;
        RECT 356.200 136.400 357.200 140.400 ;
        RECT 359.600 135.800 360.400 140.400 ;
        RECT 364.400 135.800 365.200 140.400 ;
        RECT 369.200 137.800 370.000 140.400 ;
        RECT 375.600 135.800 376.400 140.400 ;
        RECT 377.200 137.800 378.000 140.400 ;
        RECT 383.600 135.800 384.400 140.400 ;
        RECT 388.400 135.800 389.200 140.400 ;
        RECT 390.000 135.800 390.800 140.400 ;
        RECT 394.800 137.800 395.600 140.400 ;
        RECT 398.000 137.800 398.800 140.400 ;
        RECT 399.600 135.800 400.400 140.400 ;
        RECT 405.600 135.800 406.400 140.400 ;
        RECT 408.000 135.800 408.800 140.400 ;
        RECT 414.000 135.800 414.800 140.400 ;
        RECT 415.600 137.800 416.400 140.400 ;
        RECT 418.800 137.800 419.600 140.400 ;
        RECT 422.000 136.400 423.000 140.400 ;
        RECT 428.200 139.800 429.000 140.400 ;
        RECT 428.200 136.400 429.200 139.800 ;
        RECT 434.800 136.600 435.600 140.400 ;
        RECT 438.000 137.800 438.800 140.400 ;
        RECT 441.200 137.800 442.000 140.400 ;
        RECT 447.600 137.800 448.400 140.400 ;
        RECT 450.800 137.800 451.600 140.400 ;
        RECT 452.400 137.800 453.200 140.400 ;
        RECT 455.600 137.800 456.400 140.400 ;
        RECT 458.800 136.600 459.600 140.400 ;
        RECT 463.600 137.800 464.400 140.400 ;
        RECT 468.400 136.600 469.200 140.400 ;
        RECT 473.200 133.800 474.000 140.400 ;
        RECT 481.200 136.000 482.000 140.400 ;
        RECT 486.800 137.800 487.600 140.400 ;
        RECT 490.000 137.800 491.000 140.400 ;
        RECT 495.600 135.800 496.400 140.400 ;
        RECT 498.800 135.800 499.600 140.400 ;
        RECT 502.000 135.800 502.800 140.400 ;
        RECT 505.200 135.800 506.000 140.400 ;
        RECT 508.400 135.800 509.200 140.400 ;
        RECT 511.600 135.800 512.400 140.400 ;
        RECT 513.200 135.800 514.000 140.400 ;
        RECT 518.000 135.800 518.800 140.400 ;
        RECT 522.800 135.800 523.600 140.400 ;
        RECT 527.600 135.800 528.400 140.400 ;
        RECT 530.800 135.800 531.600 140.400 ;
        RECT 532.400 135.800 533.200 140.400 ;
        RECT 538.800 137.800 539.600 140.400 ;
        RECT 543.600 135.800 544.400 140.400 ;
        RECT 546.800 136.200 547.600 140.400 ;
        RECT 550.000 137.800 550.800 140.400 ;
        RECT 553.200 135.800 554.000 140.400 ;
        RECT 558.000 136.400 559.000 140.400 ;
        RECT 564.200 139.800 565.000 140.400 ;
        RECT 564.200 136.400 565.200 139.800 ;
        RECT 569.200 136.400 570.200 140.400 ;
        RECT 575.400 139.800 576.200 140.400 ;
        RECT 575.400 136.400 576.400 139.800 ;
        RECT 580.400 135.800 581.200 140.400 ;
        RECT 2.800 101.600 3.600 105.400 ;
        RECT 8.000 101.600 8.800 106.200 ;
        RECT 14.000 101.600 14.800 106.200 ;
        RECT 15.600 101.600 16.400 104.200 ;
        RECT 19.800 101.600 20.600 106.200 ;
        RECT 23.600 102.200 24.600 105.600 ;
        RECT 23.800 101.600 24.600 102.200 ;
        RECT 29.800 101.600 30.800 105.600 ;
        RECT 33.200 101.600 34.000 104.200 ;
        RECT 36.400 101.600 37.200 104.200 ;
        RECT 38.000 101.600 38.800 106.200 ;
        RECT 42.800 101.600 43.600 105.400 ;
        RECT 47.600 101.600 48.400 104.200 ;
        RECT 50.800 101.600 51.600 104.200 ;
        RECT 54.000 101.600 54.800 104.200 ;
        RECT 58.800 101.600 59.600 105.400 ;
        RECT 62.000 101.600 62.800 104.200 ;
        RECT 65.200 101.600 66.000 104.200 ;
        RECT 69.400 101.600 70.200 106.200 ;
        RECT 73.200 101.600 74.200 105.600 ;
        RECT 79.400 102.200 80.400 105.600 ;
        RECT 79.400 101.600 80.200 102.200 ;
        RECT 85.400 101.600 86.200 106.000 ;
        RECT 89.200 101.600 90.000 106.200 ;
        RECT 94.000 101.600 94.800 104.200 ;
        RECT 97.200 101.600 98.000 104.200 ;
        RECT 98.800 101.600 99.600 104.200 ;
        RECT 102.000 101.600 102.800 104.200 ;
        RECT 105.200 101.600 106.000 105.400 ;
        RECT 111.600 101.600 112.400 105.400 ;
        RECT 118.000 101.600 118.800 105.400 ;
        RECT 122.800 101.600 123.600 104.200 ;
        RECT 126.000 101.600 126.800 104.200 ;
        RECT 127.600 101.600 128.400 104.200 ;
        RECT 131.400 101.600 132.200 106.200 ;
        RECT 135.600 101.600 136.400 104.200 ;
        RECT 143.600 101.600 144.400 104.200 ;
        RECT 145.200 101.600 146.000 104.200 ;
        RECT 148.400 101.600 149.200 104.200 ;
        RECT 151.600 102.200 152.600 105.600 ;
        RECT 151.800 101.600 152.600 102.200 ;
        RECT 157.800 101.600 158.800 105.600 ;
        RECT 162.800 101.600 163.600 104.200 ;
        RECT 166.000 101.600 166.800 106.200 ;
        RECT 171.400 101.600 172.400 104.200 ;
        RECT 174.800 101.600 175.600 104.200 ;
        RECT 180.400 101.600 181.200 106.000 ;
        RECT 183.600 101.600 184.400 106.200 ;
        RECT 186.800 101.600 187.600 106.200 ;
        RECT 188.400 101.600 189.200 106.200 ;
        RECT 193.200 101.600 194.000 104.200 ;
        RECT 199.600 101.600 200.400 105.400 ;
        RECT 203.200 101.600 204.000 106.200 ;
        RECT 209.200 101.600 210.000 106.200 ;
        RECT 214.000 101.600 214.800 106.200 ;
        RECT 215.600 101.600 216.400 104.200 ;
        RECT 219.800 101.600 220.600 106.200 ;
        RECT 222.400 101.600 223.200 106.200 ;
        RECT 228.400 101.600 229.200 106.200 ;
        RECT 233.200 101.600 234.000 105.400 ;
        RECT 237.600 101.600 238.400 107.000 ;
        RECT 242.800 101.600 243.600 106.600 ;
        RECT 247.600 101.600 248.600 105.600 ;
        RECT 253.800 102.200 254.800 105.600 ;
        RECT 253.800 101.600 254.600 102.200 ;
        RECT 257.200 101.600 258.000 104.200 ;
        RECT 263.600 101.600 264.400 106.200 ;
        RECT 268.400 101.600 269.200 105.400 ;
        RECT 271.600 101.600 272.400 106.200 ;
        RECT 278.000 101.600 278.800 105.400 ;
        RECT 284.400 101.600 285.400 105.600 ;
        RECT 290.600 102.200 291.600 105.600 ;
        RECT 290.600 101.600 291.400 102.200 ;
        RECT 298.800 101.600 299.600 106.200 ;
        RECT 302.000 101.600 302.800 106.200 ;
        RECT 305.200 101.600 306.000 106.200 ;
        RECT 310.000 101.600 310.800 106.200 ;
        RECT 315.400 101.600 316.400 104.200 ;
        RECT 318.800 101.600 319.600 104.200 ;
        RECT 324.400 101.600 325.200 106.000 ;
        RECT 329.200 101.600 330.000 106.200 ;
        RECT 334.600 101.600 335.600 104.200 ;
        RECT 338.000 101.600 338.800 104.200 ;
        RECT 343.600 101.600 344.400 106.000 ;
        RECT 346.800 101.600 347.600 106.200 ;
        RECT 350.000 101.600 350.800 106.200 ;
        RECT 354.800 101.600 355.600 106.200 ;
        RECT 358.000 101.600 358.800 106.200 ;
        RECT 361.200 101.600 362.000 106.200 ;
        RECT 364.400 101.600 365.200 106.200 ;
        RECT 367.600 101.600 368.400 105.400 ;
        RECT 373.600 101.600 374.400 107.000 ;
        RECT 378.800 101.600 379.600 106.600 ;
        RECT 385.200 101.600 386.000 105.400 ;
        RECT 390.000 101.600 390.800 105.400 ;
        RECT 398.000 101.600 398.800 106.200 ;
        RECT 399.600 101.600 400.400 104.200 ;
        RECT 402.800 101.600 403.600 104.200 ;
        RECT 406.000 101.600 406.800 104.200 ;
        RECT 409.200 101.600 410.000 105.400 ;
        RECT 417.200 101.600 418.000 105.400 ;
        RECT 422.000 101.600 423.000 105.600 ;
        RECT 428.200 102.200 429.200 105.600 ;
        RECT 428.200 101.600 429.000 102.200 ;
        RECT 433.200 101.600 434.000 106.200 ;
        RECT 438.600 101.600 439.600 104.200 ;
        RECT 442.000 101.600 442.800 104.200 ;
        RECT 447.600 101.600 448.400 106.000 ;
        RECT 455.600 101.600 456.400 106.200 ;
        RECT 458.800 101.600 459.600 106.200 ;
        RECT 462.000 101.600 462.800 106.200 ;
        RECT 465.200 101.600 466.000 106.200 ;
        RECT 470.000 101.600 471.000 105.600 ;
        RECT 476.200 102.200 477.200 105.600 ;
        RECT 476.200 101.600 477.000 102.200 ;
        RECT 479.600 101.600 480.400 106.200 ;
        RECT 482.800 101.600 483.600 106.200 ;
        RECT 486.000 101.600 486.800 106.200 ;
        RECT 491.400 101.600 492.400 104.200 ;
        RECT 494.800 101.600 495.600 104.200 ;
        RECT 500.400 101.600 501.200 106.000 ;
        RECT 505.200 101.600 506.000 106.200 ;
        RECT 510.600 101.600 511.600 104.200 ;
        RECT 514.000 101.600 514.800 104.200 ;
        RECT 519.600 101.600 520.400 106.000 ;
        RECT 524.400 102.200 525.400 105.600 ;
        RECT 524.600 101.600 525.400 102.200 ;
        RECT 530.600 101.600 531.600 105.600 ;
        RECT 535.600 102.200 536.600 105.600 ;
        RECT 535.800 101.600 536.600 102.200 ;
        RECT 541.800 101.600 542.800 105.600 ;
        RECT 546.800 101.600 547.600 106.200 ;
        RECT 552.200 101.600 553.200 104.200 ;
        RECT 555.600 101.600 556.400 104.200 ;
        RECT 561.200 101.600 562.000 106.000 ;
        RECT 566.000 101.600 566.800 106.200 ;
        RECT 571.400 101.600 572.400 104.200 ;
        RECT 574.800 101.600 575.600 104.200 ;
        RECT 580.400 101.600 581.200 106.000 ;
        RECT 0.400 100.400 586.800 101.600 ;
        RECT 1.200 95.800 2.000 100.400 ;
        RECT 4.400 97.800 5.200 100.400 ;
        RECT 7.600 93.800 8.400 100.400 ;
        RECT 15.600 96.600 16.400 100.400 ;
        RECT 20.400 95.800 21.200 100.400 ;
        RECT 23.600 95.800 24.400 100.400 ;
        RECT 26.800 97.800 27.600 100.400 ;
        RECT 30.000 97.800 30.800 100.400 ;
        RECT 31.600 97.800 32.400 100.400 ;
        RECT 36.400 96.600 37.200 100.400 ;
        RECT 41.200 97.800 42.000 100.400 ;
        RECT 47.600 96.600 48.400 100.400 ;
        RECT 50.800 97.800 51.600 100.400 ;
        RECT 54.000 93.800 54.800 100.400 ;
        RECT 60.400 97.800 61.200 100.400 ;
        RECT 64.600 95.800 65.400 100.400 ;
        RECT 68.400 96.600 69.200 100.400 ;
        RECT 73.200 95.800 74.000 100.400 ;
        RECT 78.000 95.800 78.800 100.400 ;
        RECT 84.400 97.800 85.200 100.400 ;
        RECT 89.200 95.800 90.000 100.400 ;
        RECT 90.800 95.800 91.600 100.400 ;
        RECT 96.200 95.800 97.000 100.400 ;
        RECT 100.400 97.800 101.200 100.400 ;
        RECT 102.600 95.800 103.400 100.400 ;
        RECT 106.800 97.800 107.600 100.400 ;
        RECT 109.000 95.800 109.800 100.400 ;
        RECT 113.200 97.800 114.000 100.400 ;
        RECT 114.800 97.800 115.600 100.400 ;
        RECT 121.200 96.600 122.000 100.400 ;
        RECT 124.400 97.800 125.200 100.400 ;
        RECT 128.600 95.800 129.400 100.400 ;
        RECT 130.800 97.800 131.600 100.400 ;
        RECT 134.000 97.800 134.800 100.400 ;
        RECT 143.600 96.600 144.400 100.400 ;
        RECT 150.000 96.600 150.800 100.400 ;
        RECT 156.400 95.800 157.200 100.400 ;
        RECT 159.600 95.800 160.400 100.400 ;
        RECT 165.000 97.800 166.000 100.400 ;
        RECT 168.400 97.800 169.200 100.400 ;
        RECT 174.000 96.000 174.800 100.400 ;
        RECT 177.200 97.800 178.000 100.400 ;
        RECT 180.400 97.800 181.200 100.400 ;
        RECT 182.000 97.800 182.800 100.400 ;
        RECT 185.200 97.800 186.000 100.400 ;
        RECT 186.800 97.800 187.600 100.400 ;
        RECT 190.000 97.800 190.800 100.400 ;
        RECT 191.600 97.800 192.400 100.400 ;
        RECT 194.800 97.800 195.600 100.400 ;
        RECT 198.000 96.600 198.800 100.400 ;
        RECT 206.000 96.600 206.800 100.400 ;
        RECT 209.200 97.800 210.000 100.400 ;
        RECT 212.400 95.800 213.200 100.400 ;
        RECT 218.400 95.800 219.200 100.400 ;
        RECT 220.400 95.800 221.200 100.400 ;
        RECT 228.400 96.600 229.200 100.400 ;
        RECT 233.200 97.800 234.000 100.400 ;
        RECT 235.200 95.800 236.000 100.400 ;
        RECT 241.200 95.800 242.000 100.400 ;
        RECT 242.800 97.800 243.600 100.400 ;
        RECT 246.000 97.800 246.800 100.400 ;
        RECT 249.200 95.400 250.000 100.400 ;
        RECT 254.400 95.000 255.200 100.400 ;
        RECT 258.800 96.400 259.800 100.400 ;
        RECT 265.000 99.800 265.800 100.400 ;
        RECT 265.000 96.400 266.000 99.800 ;
        RECT 268.400 95.800 269.200 100.400 ;
        RECT 274.800 97.800 275.600 100.400 ;
        RECT 276.400 95.800 277.200 100.400 ;
        RECT 279.600 95.800 280.400 100.400 ;
        RECT 286.000 95.800 286.800 100.400 ;
        RECT 295.600 96.600 296.400 100.400 ;
        RECT 298.800 95.800 299.600 100.400 ;
        RECT 303.600 97.800 304.400 100.400 ;
        RECT 306.800 95.800 307.600 100.400 ;
        RECT 313.200 95.800 314.000 100.400 ;
        RECT 318.600 97.800 319.600 100.400 ;
        RECT 322.000 97.800 322.800 100.400 ;
        RECT 327.600 96.000 328.400 100.400 ;
        RECT 332.400 95.800 333.200 100.400 ;
        RECT 337.800 97.800 338.800 100.400 ;
        RECT 341.200 97.800 342.000 100.400 ;
        RECT 346.800 96.000 347.600 100.400 ;
        RECT 351.600 95.800 352.400 100.400 ;
        RECT 354.800 95.800 355.600 100.400 ;
        RECT 356.400 97.800 357.200 100.400 ;
        RECT 359.600 96.200 360.400 100.400 ;
        RECT 366.000 95.800 366.800 100.400 ;
        RECT 369.200 96.400 370.200 100.400 ;
        RECT 375.400 99.800 376.200 100.400 ;
        RECT 375.400 96.400 376.400 99.800 ;
        RECT 378.800 97.800 379.600 100.400 ;
        RECT 382.000 97.800 382.800 100.400 ;
        RECT 385.200 96.600 386.000 100.400 ;
        RECT 390.600 95.800 391.400 100.400 ;
        RECT 394.800 97.800 395.600 100.400 ;
        RECT 399.000 96.000 399.800 100.400 ;
        RECT 404.400 96.600 405.200 100.400 ;
        RECT 412.400 95.800 413.200 100.400 ;
        RECT 415.600 95.800 416.400 100.400 ;
        RECT 422.000 96.600 422.800 100.400 ;
        RECT 428.400 96.600 429.200 100.400 ;
        RECT 433.200 95.800 434.000 100.400 ;
        RECT 438.600 97.800 439.600 100.400 ;
        RECT 442.000 97.800 442.800 100.400 ;
        RECT 447.600 96.000 448.400 100.400 ;
        RECT 457.200 96.400 458.200 100.400 ;
        RECT 463.400 99.800 464.200 100.400 ;
        RECT 468.600 99.800 469.400 100.400 ;
        RECT 463.400 96.400 464.400 99.800 ;
        RECT 468.400 96.400 469.400 99.800 ;
        RECT 474.600 96.400 475.600 100.400 ;
        RECT 478.000 97.800 478.800 100.400 ;
        RECT 481.200 93.800 482.000 100.400 ;
        RECT 487.600 95.800 488.400 100.400 ;
        RECT 494.000 95.800 494.800 100.400 ;
        RECT 499.400 97.800 500.400 100.400 ;
        RECT 502.800 97.800 503.600 100.400 ;
        RECT 508.400 96.000 509.200 100.400 ;
        RECT 513.200 96.000 514.000 100.400 ;
        RECT 518.800 97.800 519.600 100.400 ;
        RECT 522.000 97.800 523.000 100.400 ;
        RECT 527.600 95.800 528.400 100.400 ;
        RECT 532.400 95.800 533.200 100.400 ;
        RECT 537.800 97.800 538.800 100.400 ;
        RECT 541.200 97.800 542.000 100.400 ;
        RECT 546.800 96.000 547.600 100.400 ;
        RECT 551.600 95.800 552.400 100.400 ;
        RECT 554.800 95.800 555.600 100.400 ;
        RECT 560.200 97.800 561.200 100.400 ;
        RECT 563.600 97.800 564.400 100.400 ;
        RECT 569.200 96.000 570.000 100.400 ;
        RECT 574.000 95.800 574.800 100.400 ;
        RECT 578.800 95.800 579.600 100.400 ;
        RECT 2.800 62.200 3.800 65.600 ;
        RECT 3.000 61.600 3.800 62.200 ;
        RECT 9.000 61.600 10.000 65.600 ;
        RECT 15.600 61.600 16.400 66.200 ;
        RECT 18.800 61.600 19.600 65.400 ;
        RECT 23.600 61.600 24.400 66.200 ;
        RECT 31.600 61.600 32.400 65.400 ;
        RECT 36.400 61.600 37.200 66.200 ;
        RECT 38.000 61.600 38.800 64.200 ;
        RECT 41.200 61.600 42.000 64.200 ;
        RECT 44.400 61.600 45.200 65.400 ;
        RECT 50.800 61.600 51.600 64.200 ;
        RECT 52.400 61.600 53.200 64.200 ;
        RECT 55.600 61.600 56.400 64.200 ;
        RECT 57.200 61.600 58.000 64.200 ;
        RECT 60.400 61.600 61.200 64.200 ;
        RECT 63.600 61.600 64.400 65.400 ;
        RECT 68.400 61.600 69.200 66.200 ;
        RECT 71.600 61.600 72.400 66.200 ;
        RECT 74.800 61.600 75.600 66.200 ;
        RECT 76.400 61.600 77.200 64.200 ;
        RECT 81.200 61.600 82.000 66.200 ;
        RECT 84.400 61.600 85.200 66.200 ;
        RECT 86.000 61.600 86.800 66.200 ;
        RECT 92.400 61.600 93.200 64.200 ;
        RECT 94.000 61.600 94.800 66.200 ;
        RECT 98.800 61.600 99.600 66.200 ;
        RECT 105.200 61.600 106.000 65.400 ;
        RECT 110.000 61.600 110.800 64.200 ;
        RECT 113.200 61.600 114.000 64.200 ;
        RECT 114.800 61.600 115.600 64.200 ;
        RECT 119.000 61.600 119.800 66.200 ;
        RECT 122.800 61.600 123.600 65.400 ;
        RECT 130.800 61.600 131.600 66.200 ;
        RECT 135.600 61.600 136.400 65.400 ;
        RECT 145.200 61.600 146.200 65.600 ;
        RECT 151.400 62.200 152.400 65.600 ;
        RECT 151.400 61.600 152.200 62.200 ;
        RECT 156.400 61.600 157.200 66.200 ;
        RECT 161.800 61.600 162.800 64.200 ;
        RECT 165.200 61.600 166.000 64.200 ;
        RECT 170.800 61.600 171.600 66.000 ;
        RECT 175.600 61.600 176.400 65.400 ;
        RECT 180.400 61.600 181.200 64.200 ;
        RECT 183.600 61.600 184.400 64.200 ;
        RECT 186.800 61.600 187.600 64.200 ;
        RECT 188.400 61.600 189.200 66.200 ;
        RECT 193.200 61.600 194.000 64.200 ;
        RECT 196.400 61.600 197.200 64.200 ;
        RECT 199.600 61.600 200.400 65.400 ;
        RECT 206.000 61.600 206.800 64.200 ;
        RECT 210.800 61.600 211.600 65.400 ;
        RECT 214.000 61.600 214.800 64.200 ;
        RECT 218.200 61.600 219.000 66.200 ;
        RECT 220.400 61.600 221.200 64.200 ;
        RECT 223.600 61.600 224.400 64.200 ;
        RECT 228.400 61.600 229.200 65.400 ;
        RECT 234.800 61.600 235.600 64.200 ;
        RECT 236.400 61.600 237.200 64.200 ;
        RECT 240.600 61.600 241.400 66.200 ;
        RECT 247.600 61.600 248.400 68.200 ;
        RECT 250.800 61.600 251.600 65.400 ;
        RECT 255.600 61.600 256.400 66.200 ;
        RECT 262.000 61.600 262.800 64.200 ;
        RECT 263.600 61.600 264.400 64.200 ;
        RECT 268.400 61.600 269.200 65.400 ;
        RECT 276.400 61.600 277.200 65.400 ;
        RECT 279.600 61.600 280.400 64.200 ;
        RECT 282.800 61.600 283.600 64.200 ;
        RECT 284.400 61.600 285.200 68.200 ;
        RECT 295.600 61.600 296.400 64.200 ;
        RECT 302.000 61.600 302.800 65.400 ;
        RECT 306.800 61.600 307.600 64.200 ;
        RECT 310.000 61.600 310.800 65.400 ;
        RECT 316.400 61.600 317.200 64.200 ;
        RECT 318.000 61.600 318.800 64.200 ;
        RECT 322.200 61.600 323.000 66.200 ;
        RECT 324.400 61.600 325.200 64.200 ;
        RECT 327.600 61.600 328.400 64.200 ;
        RECT 330.800 61.600 331.600 64.200 ;
        RECT 334.000 61.600 335.000 65.600 ;
        RECT 340.200 62.200 341.200 65.600 ;
        RECT 340.200 61.600 341.000 62.200 ;
        RECT 345.200 61.600 346.000 66.200 ;
        RECT 350.600 61.600 351.600 64.200 ;
        RECT 354.000 61.600 354.800 64.200 ;
        RECT 359.600 61.600 360.400 66.000 ;
        RECT 364.400 61.600 365.200 66.200 ;
        RECT 369.800 61.600 370.800 64.200 ;
        RECT 373.200 61.600 374.000 64.200 ;
        RECT 378.800 61.600 379.600 66.000 ;
        RECT 382.000 61.600 382.800 66.200 ;
        RECT 386.800 61.600 387.600 64.200 ;
        RECT 391.600 61.600 392.400 65.400 ;
        RECT 399.600 61.600 400.400 65.400 ;
        RECT 402.800 61.600 403.600 66.200 ;
        RECT 407.600 61.600 408.400 66.200 ;
        RECT 412.400 61.600 413.200 66.200 ;
        RECT 415.600 61.600 416.400 64.200 ;
        RECT 418.800 61.600 419.600 64.200 ;
        RECT 422.000 61.600 422.800 64.200 ;
        RECT 423.600 61.600 424.400 66.200 ;
        RECT 430.000 61.600 430.800 64.200 ;
        RECT 432.200 61.600 433.000 66.200 ;
        RECT 436.400 61.600 437.200 64.200 ;
        RECT 439.600 61.600 440.600 65.600 ;
        RECT 445.800 62.200 446.800 65.600 ;
        RECT 445.800 61.600 446.600 62.200 ;
        RECT 458.800 61.600 459.600 65.400 ;
        RECT 463.600 62.200 464.600 65.600 ;
        RECT 463.800 61.600 464.600 62.200 ;
        RECT 469.800 61.600 470.800 65.600 ;
        RECT 474.800 61.600 475.600 65.400 ;
        RECT 479.600 61.600 480.400 64.200 ;
        RECT 482.800 61.600 483.600 64.200 ;
        RECT 484.400 61.600 485.200 64.200 ;
        RECT 490.800 61.600 491.600 65.400 ;
        RECT 497.200 61.600 498.000 65.400 ;
        RECT 500.400 61.600 501.200 64.200 ;
        RECT 506.800 61.600 507.600 65.400 ;
        RECT 510.000 61.600 510.800 64.200 ;
        RECT 513.200 61.600 514.000 64.200 ;
        RECT 514.800 61.600 515.600 64.200 ;
        RECT 518.000 61.600 518.800 64.200 ;
        RECT 521.200 61.600 522.000 65.400 ;
        RECT 529.200 61.600 530.000 65.400 ;
        RECT 534.000 61.600 534.800 66.200 ;
        RECT 538.800 61.600 539.600 66.200 ;
        RECT 543.600 61.600 544.400 66.200 ;
        RECT 549.000 61.600 550.000 64.200 ;
        RECT 552.400 61.600 553.200 64.200 ;
        RECT 558.000 61.600 558.800 66.000 ;
        RECT 562.800 61.600 563.600 66.200 ;
        RECT 568.200 61.600 569.200 64.200 ;
        RECT 571.600 61.600 572.400 64.200 ;
        RECT 577.200 61.600 578.000 66.000 ;
        RECT 582.000 61.600 582.800 66.200 ;
        RECT 0.400 60.400 586.800 61.600 ;
        RECT 1.200 57.800 2.000 60.400 ;
        RECT 4.400 57.800 5.200 60.400 ;
        RECT 6.000 55.800 6.800 60.400 ;
        RECT 10.800 55.800 11.600 60.400 ;
        RECT 15.600 57.800 16.400 60.400 ;
        RECT 18.800 57.800 19.600 60.400 ;
        RECT 20.400 55.800 21.200 60.400 ;
        RECT 25.200 55.800 26.000 60.400 ;
        RECT 31.200 55.800 32.000 60.400 ;
        RECT 33.200 57.800 34.000 60.400 ;
        RECT 36.400 55.800 37.200 60.400 ;
        RECT 42.400 55.800 43.200 60.400 ;
        RECT 49.200 53.800 50.000 60.400 ;
        RECT 54.000 56.600 54.800 60.400 ;
        RECT 57.200 57.800 58.000 60.400 ;
        RECT 60.400 57.800 61.200 60.400 ;
        RECT 63.600 57.800 64.400 60.400 ;
        RECT 67.800 55.800 68.600 60.400 ;
        RECT 71.200 55.000 72.000 60.400 ;
        RECT 76.400 55.400 77.200 60.400 ;
        RECT 81.200 56.600 82.000 60.400 ;
        RECT 89.200 55.800 90.000 60.400 ;
        RECT 94.000 55.800 94.800 60.400 ;
        RECT 98.800 55.800 99.600 60.400 ;
        RECT 102.000 56.600 102.800 60.400 ;
        RECT 106.800 57.800 107.600 60.400 ;
        RECT 111.600 56.600 112.400 60.400 ;
        RECT 116.400 57.800 117.200 60.400 ;
        RECT 119.600 57.800 120.400 60.400 ;
        RECT 122.800 57.800 123.600 60.400 ;
        RECT 127.600 56.600 128.400 60.400 ;
        RECT 132.400 57.800 133.200 60.400 ;
        RECT 140.400 56.600 141.200 60.400 ;
        RECT 146.800 57.800 147.600 60.400 ;
        RECT 148.400 57.800 149.200 60.400 ;
        RECT 152.600 55.800 153.400 60.400 ;
        RECT 156.400 56.400 157.400 60.400 ;
        RECT 162.600 59.800 163.400 60.400 ;
        RECT 162.600 56.400 163.600 59.800 ;
        RECT 167.600 56.400 168.600 60.400 ;
        RECT 173.800 59.800 174.600 60.400 ;
        RECT 173.800 56.400 174.800 59.800 ;
        RECT 178.800 55.800 179.600 60.400 ;
        RECT 184.200 57.800 185.200 60.400 ;
        RECT 187.600 57.800 188.400 60.400 ;
        RECT 193.200 56.000 194.000 60.400 ;
        RECT 198.000 55.800 198.800 60.400 ;
        RECT 201.200 56.400 202.200 60.400 ;
        RECT 207.400 59.800 208.200 60.400 ;
        RECT 207.400 56.400 208.400 59.800 ;
        RECT 214.000 56.600 214.800 60.400 ;
        RECT 217.200 55.800 218.000 60.400 ;
        RECT 220.400 57.800 221.200 60.400 ;
        RECT 223.600 57.800 224.400 60.400 ;
        RECT 225.200 57.800 226.000 60.400 ;
        RECT 228.400 57.800 229.200 60.400 ;
        RECT 230.000 57.800 230.800 60.400 ;
        RECT 233.200 57.800 234.000 60.400 ;
        RECT 236.400 56.600 237.200 60.400 ;
        RECT 243.000 59.800 243.800 60.400 ;
        RECT 242.800 56.400 243.800 59.800 ;
        RECT 249.000 56.400 250.000 60.400 ;
        RECT 254.000 55.800 254.800 60.400 ;
        RECT 257.200 55.800 258.000 60.400 ;
        RECT 260.400 55.800 261.200 60.400 ;
        RECT 265.200 55.800 266.000 60.400 ;
        RECT 268.400 55.800 269.200 60.400 ;
        RECT 271.600 55.800 272.400 60.400 ;
        RECT 276.400 55.800 277.200 60.400 ;
        RECT 278.000 57.800 278.800 60.400 ;
        RECT 281.200 57.800 282.000 60.400 ;
        RECT 282.800 57.800 283.600 60.400 ;
        RECT 286.000 57.800 286.800 60.400 ;
        RECT 294.000 56.600 294.800 60.400 ;
        RECT 298.800 57.800 299.600 60.400 ;
        RECT 303.000 55.800 303.800 60.400 ;
        RECT 305.200 55.800 306.000 60.400 ;
        RECT 311.600 57.800 312.400 60.400 ;
        RECT 313.600 55.800 314.400 60.400 ;
        RECT 319.600 55.800 320.400 60.400 ;
        RECT 321.600 55.800 322.400 60.400 ;
        RECT 327.600 55.800 328.400 60.400 ;
        RECT 329.200 57.800 330.000 60.400 ;
        RECT 332.400 57.800 333.200 60.400 ;
        RECT 335.600 55.800 336.400 60.400 ;
        RECT 340.400 56.600 341.200 60.400 ;
        RECT 348.400 56.600 349.200 60.400 ;
        RECT 353.200 55.800 354.000 60.400 ;
        RECT 358.600 57.800 359.600 60.400 ;
        RECT 362.000 57.800 362.800 60.400 ;
        RECT 367.600 56.000 368.400 60.400 ;
        RECT 372.400 55.800 373.200 60.400 ;
        RECT 377.800 57.800 378.800 60.400 ;
        RECT 381.200 57.800 382.000 60.400 ;
        RECT 386.800 56.000 387.600 60.400 ;
        RECT 390.000 57.800 390.800 60.400 ;
        RECT 396.400 55.800 397.200 60.400 ;
        RECT 399.600 55.800 400.400 60.400 ;
        RECT 405.000 57.800 406.000 60.400 ;
        RECT 408.400 57.800 409.200 60.400 ;
        RECT 414.000 56.000 414.800 60.400 ;
        RECT 418.800 55.800 419.600 60.400 ;
        RECT 422.000 55.800 422.800 60.400 ;
        RECT 425.400 59.800 426.200 60.400 ;
        RECT 425.200 56.400 426.200 59.800 ;
        RECT 431.400 56.400 432.400 60.400 ;
        RECT 436.400 56.600 437.200 60.400 ;
        RECT 441.200 57.800 442.000 60.400 ;
        RECT 449.200 55.800 450.000 60.400 ;
        RECT 457.200 56.600 458.000 60.400 ;
        RECT 460.400 55.800 461.200 60.400 ;
        RECT 467.400 56.000 468.200 60.400 ;
        RECT 472.200 55.800 473.000 60.400 ;
        RECT 476.400 57.800 477.200 60.400 ;
        RECT 478.000 57.800 478.800 60.400 ;
        RECT 481.200 57.800 482.000 60.400 ;
        RECT 482.800 57.800 483.600 60.400 ;
        RECT 486.000 57.800 486.800 60.400 ;
        RECT 489.200 56.600 490.000 60.400 ;
        RECT 494.000 57.800 494.800 60.400 ;
        RECT 497.200 57.800 498.000 60.400 ;
        RECT 501.400 55.800 502.200 60.400 ;
        RECT 503.600 57.800 504.400 60.400 ;
        RECT 507.800 55.800 508.600 60.400 ;
        RECT 511.600 57.800 512.400 60.400 ;
        RECT 514.800 56.400 515.800 60.400 ;
        RECT 521.000 59.800 521.800 60.400 ;
        RECT 521.000 56.400 522.000 59.800 ;
        RECT 526.000 55.800 526.800 60.400 ;
        RECT 531.400 57.800 532.400 60.400 ;
        RECT 534.800 57.800 535.600 60.400 ;
        RECT 540.400 56.000 541.200 60.400 ;
        RECT 545.200 56.000 546.000 60.400 ;
        RECT 550.800 57.800 551.600 60.400 ;
        RECT 554.000 57.800 555.000 60.400 ;
        RECT 559.600 55.800 560.400 60.400 ;
        RECT 564.400 56.000 565.200 60.400 ;
        RECT 570.000 57.800 570.800 60.400 ;
        RECT 573.200 57.800 574.200 60.400 ;
        RECT 578.800 55.800 579.600 60.400 ;
        RECT 1.200 21.600 2.000 24.200 ;
        RECT 4.400 21.600 5.200 26.200 ;
        RECT 9.200 21.600 10.000 26.200 ;
        RECT 14.000 21.600 14.800 24.200 ;
        RECT 18.200 21.600 19.000 26.200 ;
        RECT 23.600 21.600 24.400 25.400 ;
        RECT 28.400 21.600 29.200 26.200 ;
        RECT 31.600 21.600 32.400 26.200 ;
        RECT 39.600 21.600 40.400 25.400 ;
        RECT 43.400 21.600 44.200 26.200 ;
        RECT 47.600 21.600 48.400 24.200 ;
        RECT 49.200 21.600 50.000 24.200 ;
        RECT 54.000 21.600 54.800 26.200 ;
        RECT 57.200 21.600 58.000 26.200 ;
        RECT 60.400 21.600 61.400 25.600 ;
        RECT 66.600 22.200 67.600 25.600 ;
        RECT 66.600 21.600 67.400 22.200 ;
        RECT 71.600 21.600 72.400 26.200 ;
        RECT 77.000 21.600 78.000 24.200 ;
        RECT 80.400 21.600 81.200 24.200 ;
        RECT 86.000 21.600 86.800 26.000 ;
        RECT 90.800 22.200 91.800 25.600 ;
        RECT 91.000 21.600 91.800 22.200 ;
        RECT 97.000 21.600 98.000 25.600 ;
        RECT 103.600 21.600 104.400 25.400 ;
        RECT 108.400 21.600 109.200 26.200 ;
        RECT 113.800 21.600 114.800 24.200 ;
        RECT 117.200 21.600 118.000 24.200 ;
        RECT 122.800 21.600 123.600 26.000 ;
        RECT 127.600 21.600 128.600 25.600 ;
        RECT 133.800 22.200 134.800 25.600 ;
        RECT 133.800 21.600 134.600 22.200 ;
        RECT 143.600 21.600 144.600 25.600 ;
        RECT 149.800 22.200 150.800 25.600 ;
        RECT 149.800 21.600 150.600 22.200 ;
        RECT 153.200 21.600 154.000 26.200 ;
        RECT 158.000 21.600 158.800 24.200 ;
        RECT 161.200 21.600 162.000 26.200 ;
        RECT 170.800 21.600 171.600 25.400 ;
        RECT 175.600 21.600 176.400 25.400 ;
        RECT 183.600 21.600 184.400 25.400 ;
        RECT 188.400 21.600 189.400 25.600 ;
        RECT 194.600 22.200 195.600 25.600 ;
        RECT 194.600 21.600 195.400 22.200 ;
        RECT 198.600 21.600 199.400 26.200 ;
        RECT 202.800 21.600 203.600 24.200 ;
        RECT 207.000 21.600 207.800 26.000 ;
        RECT 214.000 21.600 214.800 26.200 ;
        RECT 215.600 21.600 216.400 26.200 ;
        RECT 222.000 22.200 223.000 25.600 ;
        RECT 222.200 21.600 223.000 22.200 ;
        RECT 228.200 21.600 229.200 25.600 ;
        RECT 234.800 21.600 235.600 26.200 ;
        RECT 236.400 21.600 237.200 24.200 ;
        RECT 239.600 21.600 240.400 24.200 ;
        RECT 241.200 21.600 242.000 26.200 ;
        RECT 247.200 21.600 248.000 26.200 ;
        RECT 249.600 21.600 250.400 26.200 ;
        RECT 255.600 21.600 256.400 26.200 ;
        RECT 260.400 21.600 261.200 26.200 ;
        RECT 265.200 21.600 266.000 26.200 ;
        RECT 268.400 21.600 269.200 25.400 ;
        RECT 276.400 21.600 277.200 25.400 ;
        RECT 281.200 21.600 282.000 25.400 ;
        RECT 287.600 21.600 288.400 25.400 ;
        RECT 300.400 21.600 301.200 25.400 ;
        RECT 303.600 21.600 304.400 24.200 ;
        RECT 306.800 21.600 307.600 24.200 ;
        RECT 310.000 21.600 310.800 25.400 ;
        RECT 318.000 21.600 318.800 25.400 ;
        RECT 322.800 21.600 323.600 24.200 ;
        RECT 324.400 21.600 325.200 24.200 ;
        RECT 327.600 21.600 328.400 24.200 ;
        RECT 330.800 21.600 331.600 24.200 ;
        RECT 335.600 21.600 336.400 25.400 ;
        RECT 338.800 21.600 339.600 24.200 ;
        RECT 342.000 21.600 342.800 24.200 ;
        RECT 343.600 21.600 344.400 24.200 ;
        RECT 347.800 21.600 348.600 26.200 ;
        RECT 353.200 21.600 354.000 26.200 ;
        RECT 356.400 21.600 357.200 25.400 ;
        RECT 361.200 21.600 362.000 24.200 ;
        RECT 366.000 21.600 367.000 25.600 ;
        RECT 372.200 22.200 373.200 25.600 ;
        RECT 372.200 21.600 373.000 22.200 ;
        RECT 377.200 21.600 378.000 26.200 ;
        RECT 382.600 21.600 383.600 24.200 ;
        RECT 386.000 21.600 386.800 24.200 ;
        RECT 391.600 21.600 392.400 26.000 ;
        RECT 396.400 21.600 397.200 26.200 ;
        RECT 399.600 21.600 400.400 26.200 ;
        RECT 402.800 22.200 403.800 25.600 ;
        RECT 403.000 21.600 403.800 22.200 ;
        RECT 409.000 21.600 410.000 25.600 ;
        RECT 412.400 21.600 413.200 26.200 ;
        RECT 418.800 21.600 419.600 25.400 ;
        RECT 423.600 21.600 424.400 26.200 ;
        RECT 428.400 21.600 429.200 26.200 ;
        RECT 433.200 21.600 434.000 24.200 ;
        RECT 436.400 21.600 437.200 24.200 ;
        RECT 439.600 21.600 440.400 25.400 ;
        RECT 449.200 21.600 450.000 26.200 ;
        RECT 454.000 21.600 454.800 26.200 ;
        RECT 462.000 21.600 462.800 25.400 ;
        RECT 468.400 21.600 469.200 26.200 ;
        RECT 470.000 21.600 470.800 26.200 ;
        RECT 476.000 21.600 476.800 26.200 ;
        RECT 478.000 21.600 478.800 26.200 ;
        RECT 484.000 21.600 484.800 26.200 ;
        RECT 487.600 21.600 488.400 25.400 ;
        RECT 495.600 21.600 496.400 25.400 ;
        RECT 502.000 21.600 502.800 25.400 ;
        RECT 505.600 21.600 506.400 26.200 ;
        RECT 511.600 21.600 512.400 26.200 ;
        RECT 514.800 21.600 515.600 24.200 ;
        RECT 516.800 21.600 517.600 26.200 ;
        RECT 522.800 21.600 523.600 26.200 ;
        RECT 524.400 21.600 525.200 24.200 ;
        RECT 527.600 21.600 528.400 24.200 ;
        RECT 530.800 21.600 531.800 25.600 ;
        RECT 537.000 22.200 538.000 25.600 ;
        RECT 537.000 21.600 537.800 22.200 ;
        RECT 540.400 21.600 541.200 24.200 ;
        RECT 543.600 21.600 544.400 24.200 ;
        RECT 545.200 21.600 546.000 24.200 ;
        RECT 549.400 21.600 550.200 26.200 ;
        RECT 554.800 21.600 555.600 26.200 ;
        RECT 558.000 21.600 558.800 24.200 ;
        RECT 562.800 21.600 563.600 25.400 ;
        RECT 567.600 21.600 568.600 25.600 ;
        RECT 573.800 22.200 574.800 25.600 ;
        RECT 573.800 21.600 574.600 22.200 ;
        RECT 578.800 21.600 579.600 25.400 ;
        RECT 0.400 20.400 586.800 21.600 ;
        RECT 1.200 17.800 2.000 20.400 ;
        RECT 9.200 13.800 10.000 20.400 ;
        RECT 14.000 16.600 14.800 20.400 ;
        RECT 18.800 16.400 19.800 20.400 ;
        RECT 25.000 19.800 25.800 20.400 ;
        RECT 25.000 16.400 26.000 19.800 ;
        RECT 30.000 16.400 31.000 20.400 ;
        RECT 36.200 19.800 37.000 20.400 ;
        RECT 36.200 16.400 37.200 19.800 ;
        RECT 41.200 15.800 42.000 20.400 ;
        RECT 46.600 17.800 47.600 20.400 ;
        RECT 50.000 17.800 50.800 20.400 ;
        RECT 55.600 16.000 56.400 20.400 ;
        RECT 60.400 15.800 61.200 20.400 ;
        RECT 65.800 17.800 66.800 20.400 ;
        RECT 69.200 17.800 70.000 20.400 ;
        RECT 74.800 16.000 75.600 20.400 ;
        RECT 79.600 15.800 80.400 20.400 ;
        RECT 85.000 17.800 86.000 20.400 ;
        RECT 88.400 17.800 89.200 20.400 ;
        RECT 94.000 16.000 94.800 20.400 ;
        RECT 98.800 15.800 99.600 20.400 ;
        RECT 104.200 17.800 105.200 20.400 ;
        RECT 107.600 17.800 108.400 20.400 ;
        RECT 113.200 16.000 114.000 20.400 ;
        RECT 118.000 15.800 118.800 20.400 ;
        RECT 123.400 17.800 124.400 20.400 ;
        RECT 126.800 17.800 127.600 20.400 ;
        RECT 132.400 16.000 133.200 20.400 ;
        RECT 142.200 19.800 143.000 20.400 ;
        RECT 142.000 16.400 143.000 19.800 ;
        RECT 148.200 16.400 149.200 20.400 ;
        RECT 153.200 16.600 154.000 20.400 ;
        RECT 159.600 17.800 160.400 20.400 ;
        RECT 161.200 17.800 162.000 20.400 ;
        RECT 164.400 17.800 165.200 20.400 ;
        RECT 167.600 17.800 168.400 20.400 ;
        RECT 169.200 17.800 170.000 20.400 ;
        RECT 173.400 15.800 174.200 20.400 ;
        RECT 177.200 15.800 178.000 20.400 ;
        RECT 180.400 15.800 181.200 20.400 ;
        RECT 183.800 19.800 184.600 20.400 ;
        RECT 183.600 16.400 184.600 19.800 ;
        RECT 189.800 16.400 190.800 20.400 ;
        RECT 194.800 16.600 195.600 20.400 ;
        RECT 201.200 16.600 202.000 20.400 ;
        RECT 209.200 16.600 210.000 20.400 ;
        RECT 212.400 17.800 213.200 20.400 ;
        RECT 215.600 17.800 216.400 20.400 ;
        RECT 218.800 17.800 219.600 20.400 ;
        RECT 223.600 15.800 224.400 20.400 ;
        RECT 225.200 15.800 226.000 20.400 ;
        RECT 231.600 17.800 232.400 20.400 ;
        RECT 235.000 19.800 235.800 20.400 ;
        RECT 234.800 16.400 235.800 19.800 ;
        RECT 241.000 16.400 242.000 20.400 ;
        RECT 247.600 15.800 248.400 20.400 ;
        RECT 249.200 15.800 250.000 20.400 ;
        RECT 255.600 16.600 256.400 20.400 ;
        RECT 260.400 15.800 261.200 20.400 ;
        RECT 266.800 16.400 267.800 20.400 ;
        RECT 273.000 19.800 273.800 20.400 ;
        RECT 273.000 16.400 274.000 19.800 ;
        RECT 278.000 16.600 278.800 20.400 ;
        RECT 284.400 16.400 285.400 20.400 ;
        RECT 290.600 19.800 291.400 20.400 ;
        RECT 290.600 16.400 291.600 19.800 ;
        RECT 298.800 15.800 299.600 20.400 ;
        RECT 306.800 16.600 307.600 20.400 ;
        RECT 310.000 17.800 310.800 20.400 ;
        RECT 316.400 15.800 317.200 20.400 ;
        RECT 319.200 15.000 320.000 20.400 ;
        RECT 324.400 15.400 325.200 20.400 ;
        RECT 329.400 19.800 330.200 20.400 ;
        RECT 329.200 16.400 330.200 19.800 ;
        RECT 335.400 16.400 336.400 20.400 ;
        RECT 340.400 15.800 341.200 20.400 ;
        RECT 345.800 17.800 346.800 20.400 ;
        RECT 349.200 17.800 350.000 20.400 ;
        RECT 354.800 16.000 355.600 20.400 ;
        RECT 359.600 15.800 360.400 20.400 ;
        RECT 365.000 17.800 366.000 20.400 ;
        RECT 368.400 17.800 369.200 20.400 ;
        RECT 374.000 16.000 374.800 20.400 ;
        RECT 378.800 15.800 379.600 20.400 ;
        RECT 384.200 17.800 385.200 20.400 ;
        RECT 387.600 17.800 388.400 20.400 ;
        RECT 393.200 16.000 394.000 20.400 ;
        RECT 398.000 15.800 398.800 20.400 ;
        RECT 401.200 15.800 402.000 20.400 ;
        RECT 404.400 16.400 405.400 20.400 ;
        RECT 410.600 19.800 411.400 20.400 ;
        RECT 410.600 16.400 411.600 19.800 ;
        RECT 414.000 17.800 414.800 20.400 ;
        RECT 418.800 16.600 419.600 20.400 ;
        RECT 426.800 16.600 427.600 20.400 ;
        RECT 430.000 15.800 430.800 20.400 ;
        RECT 436.400 15.800 437.200 20.400 ;
        RECT 439.600 15.800 440.400 20.400 ;
        RECT 441.200 17.800 442.000 20.400 ;
        RECT 449.200 15.800 450.000 20.400 ;
        RECT 457.200 15.800 458.000 20.400 ;
        RECT 458.800 17.800 459.600 20.400 ;
        RECT 462.000 17.800 462.800 20.400 ;
        RECT 465.200 16.600 466.000 20.400 ;
        RECT 471.800 19.800 472.600 20.400 ;
        RECT 471.600 16.400 472.600 19.800 ;
        RECT 477.800 16.400 478.800 20.400 ;
        RECT 482.800 16.600 483.600 20.400 ;
        RECT 490.800 16.600 491.600 20.400 ;
        RECT 495.600 16.600 496.400 20.400 ;
        RECT 500.400 17.800 501.200 20.400 ;
        RECT 503.600 16.200 504.400 20.400 ;
        RECT 506.800 17.800 507.600 20.400 ;
        RECT 510.000 17.800 510.800 20.400 ;
        RECT 511.600 17.800 512.400 20.400 ;
        RECT 514.800 15.800 515.600 20.400 ;
        RECT 518.000 15.800 518.800 20.400 ;
        RECT 521.200 17.800 522.000 20.400 ;
        RECT 527.600 16.600 528.400 20.400 ;
        RECT 530.800 17.800 531.600 20.400 ;
        RECT 534.000 17.800 534.800 20.400 ;
        RECT 535.600 17.800 536.400 20.400 ;
        RECT 538.800 17.800 539.600 20.400 ;
        RECT 540.400 15.800 541.200 20.400 ;
        RECT 543.600 17.800 544.400 20.400 ;
        RECT 547.800 15.800 548.600 20.400 ;
        RECT 550.000 17.800 550.800 20.400 ;
        RECT 553.200 17.800 554.000 20.400 ;
        RECT 557.400 16.000 558.200 20.400 ;
        RECT 562.800 16.400 563.800 20.400 ;
        RECT 569.000 19.800 569.800 20.400 ;
        RECT 569.000 16.400 570.000 19.800 ;
        RECT 574.000 16.600 574.800 20.400 ;
        RECT 580.400 15.800 581.200 20.400 ;
      LAYER via1 ;
        RECT 291.000 420.600 291.800 421.400 ;
        RECT 292.400 420.600 293.200 421.400 ;
        RECT 293.800 420.600 294.600 421.400 ;
        RECT 291.000 380.600 291.800 381.400 ;
        RECT 292.400 380.600 293.200 381.400 ;
        RECT 293.800 380.600 294.600 381.400 ;
        RECT 291.000 340.600 291.800 341.400 ;
        RECT 292.400 340.600 293.200 341.400 ;
        RECT 293.800 340.600 294.600 341.400 ;
        RECT 222.000 309.600 222.800 310.400 ;
        RECT 220.400 305.400 221.200 306.200 ;
        RECT 291.000 300.600 291.800 301.400 ;
        RECT 292.400 300.600 293.200 301.400 ;
        RECT 293.800 300.600 294.600 301.400 ;
        RECT 291.000 260.600 291.800 261.400 ;
        RECT 292.400 260.600 293.200 261.400 ;
        RECT 293.800 260.600 294.600 261.400 ;
        RECT 291.000 220.600 291.800 221.400 ;
        RECT 292.400 220.600 293.200 221.400 ;
        RECT 293.800 220.600 294.600 221.400 ;
        RECT 291.000 180.600 291.800 181.400 ;
        RECT 292.400 180.600 293.200 181.400 ;
        RECT 293.800 180.600 294.600 181.400 ;
        RECT 291.000 140.600 291.800 141.400 ;
        RECT 292.400 140.600 293.200 141.400 ;
        RECT 293.800 140.600 294.600 141.400 ;
        RECT 291.000 100.600 291.800 101.400 ;
        RECT 292.400 100.600 293.200 101.400 ;
        RECT 293.800 100.600 294.600 101.400 ;
        RECT 291.000 60.600 291.800 61.400 ;
        RECT 292.400 60.600 293.200 61.400 ;
        RECT 293.800 60.600 294.600 61.400 ;
        RECT 291.000 20.600 291.800 21.400 ;
        RECT 292.400 20.600 293.200 21.400 ;
        RECT 293.800 20.600 294.600 21.400 ;
      LAYER metal2 ;
        RECT 290.400 420.600 295.200 421.400 ;
        RECT 290.400 380.600 295.200 381.400 ;
        RECT 290.400 340.600 295.200 341.400 ;
        RECT 222.000 309.600 222.800 310.400 ;
        RECT 222.100 306.300 222.700 309.600 ;
        RECT 220.500 306.200 222.700 306.300 ;
        RECT 220.400 305.700 222.700 306.200 ;
        RECT 220.400 305.400 221.200 305.700 ;
        RECT 220.500 292.400 221.100 305.400 ;
        RECT 231.600 302.300 232.400 302.400 ;
        RECT 231.600 301.700 233.900 302.300 ;
        RECT 231.600 301.600 232.400 301.700 ;
        RECT 223.600 296.300 224.400 296.600 ;
        RECT 222.100 295.800 224.400 296.300 ;
        RECT 222.100 295.700 224.300 295.800 ;
        RECT 222.100 292.400 222.700 295.700 ;
        RECT 233.300 292.400 233.900 301.700 ;
        RECT 290.400 300.600 295.200 301.400 ;
        RECT 220.400 291.600 221.200 292.400 ;
        RECT 222.000 291.600 222.800 292.400 ;
        RECT 233.200 291.600 234.000 292.400 ;
        RECT 290.400 260.600 295.200 261.400 ;
        RECT 290.400 220.600 295.200 221.400 ;
        RECT 290.400 180.600 295.200 181.400 ;
        RECT 290.400 140.600 295.200 141.400 ;
        RECT 290.400 100.600 295.200 101.400 ;
        RECT 290.400 60.600 295.200 61.400 ;
        RECT 290.400 20.600 295.200 21.400 ;
      LAYER via2 ;
        RECT 291.000 420.600 291.800 421.400 ;
        RECT 292.400 420.600 293.200 421.400 ;
        RECT 293.800 420.600 294.600 421.400 ;
        RECT 291.000 380.600 291.800 381.400 ;
        RECT 292.400 380.600 293.200 381.400 ;
        RECT 293.800 380.600 294.600 381.400 ;
        RECT 291.000 340.600 291.800 341.400 ;
        RECT 292.400 340.600 293.200 341.400 ;
        RECT 293.800 340.600 294.600 341.400 ;
        RECT 291.000 300.600 291.800 301.400 ;
        RECT 292.400 300.600 293.200 301.400 ;
        RECT 293.800 300.600 294.600 301.400 ;
        RECT 291.000 260.600 291.800 261.400 ;
        RECT 292.400 260.600 293.200 261.400 ;
        RECT 293.800 260.600 294.600 261.400 ;
        RECT 291.000 220.600 291.800 221.400 ;
        RECT 292.400 220.600 293.200 221.400 ;
        RECT 293.800 220.600 294.600 221.400 ;
        RECT 291.000 180.600 291.800 181.400 ;
        RECT 292.400 180.600 293.200 181.400 ;
        RECT 293.800 180.600 294.600 181.400 ;
        RECT 291.000 140.600 291.800 141.400 ;
        RECT 292.400 140.600 293.200 141.400 ;
        RECT 293.800 140.600 294.600 141.400 ;
        RECT 291.000 100.600 291.800 101.400 ;
        RECT 292.400 100.600 293.200 101.400 ;
        RECT 293.800 100.600 294.600 101.400 ;
        RECT 291.000 60.600 291.800 61.400 ;
        RECT 292.400 60.600 293.200 61.400 ;
        RECT 293.800 60.600 294.600 61.400 ;
        RECT 291.000 20.600 291.800 21.400 ;
        RECT 292.400 20.600 293.200 21.400 ;
        RECT 293.800 20.600 294.600 21.400 ;
      LAYER metal3 ;
        RECT 290.400 420.400 295.200 421.600 ;
        RECT 290.400 380.400 295.200 381.600 ;
        RECT 290.400 340.400 295.200 341.600 ;
        RECT 290.400 300.400 295.200 301.600 ;
        RECT 290.400 260.400 295.200 261.600 ;
        RECT 290.400 220.400 295.200 221.600 ;
        RECT 290.400 180.400 295.200 181.600 ;
        RECT 290.400 140.400 295.200 141.600 ;
        RECT 290.400 100.400 295.200 101.600 ;
        RECT 290.400 60.400 295.200 61.600 ;
        RECT 290.400 20.400 295.200 21.600 ;
      LAYER via3 ;
        RECT 290.800 420.600 291.600 421.400 ;
        RECT 292.400 420.600 293.200 421.400 ;
        RECT 294.000 420.600 294.800 421.400 ;
        RECT 290.800 380.600 291.600 381.400 ;
        RECT 292.400 380.600 293.200 381.400 ;
        RECT 294.000 380.600 294.800 381.400 ;
        RECT 290.800 340.600 291.600 341.400 ;
        RECT 292.400 340.600 293.200 341.400 ;
        RECT 294.000 340.600 294.800 341.400 ;
        RECT 290.800 300.600 291.600 301.400 ;
        RECT 292.400 300.600 293.200 301.400 ;
        RECT 294.000 300.600 294.800 301.400 ;
        RECT 290.800 260.600 291.600 261.400 ;
        RECT 292.400 260.600 293.200 261.400 ;
        RECT 294.000 260.600 294.800 261.400 ;
        RECT 290.800 220.600 291.600 221.400 ;
        RECT 292.400 220.600 293.200 221.400 ;
        RECT 294.000 220.600 294.800 221.400 ;
        RECT 290.800 180.600 291.600 181.400 ;
        RECT 292.400 180.600 293.200 181.400 ;
        RECT 294.000 180.600 294.800 181.400 ;
        RECT 290.800 140.600 291.600 141.400 ;
        RECT 292.400 140.600 293.200 141.400 ;
        RECT 294.000 140.600 294.800 141.400 ;
        RECT 290.800 100.600 291.600 101.400 ;
        RECT 292.400 100.600 293.200 101.400 ;
        RECT 294.000 100.600 294.800 101.400 ;
        RECT 290.800 60.600 291.600 61.400 ;
        RECT 292.400 60.600 293.200 61.400 ;
        RECT 294.000 60.600 294.800 61.400 ;
        RECT 290.800 20.600 291.600 21.400 ;
        RECT 292.400 20.600 293.200 21.400 ;
        RECT 294.000 20.600 294.800 21.400 ;
      LAYER metal4 ;
        RECT 290.400 0.000 295.200 424.000 ;
    END
  END gnd
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 97.200 413.800 98.000 414.400 ;
        RECT 314.800 413.800 315.600 414.400 ;
        RECT 96.200 413.000 98.000 413.800 ;
        RECT 313.800 413.000 315.600 413.800 ;
        RECT 387.400 388.200 389.200 389.000 ;
        RECT 388.400 387.600 389.200 388.200 ;
        RECT 500.400 348.200 502.200 349.000 ;
        RECT 500.400 347.600 501.200 348.200 ;
        RECT 198.000 333.800 198.800 334.400 ;
        RECT 197.000 333.000 198.800 333.800 ;
        RECT 495.600 293.800 496.400 294.400 ;
        RECT 495.600 293.000 497.400 293.800 ;
        RECT 183.600 228.200 185.400 229.000 ;
        RECT 183.600 227.600 184.400 228.200 ;
        RECT 110.000 213.800 110.800 214.400 ;
        RECT 109.000 213.000 110.800 213.800 ;
        RECT 252.400 173.800 253.200 174.400 ;
        RECT 252.400 173.000 254.200 173.800 ;
        RECT 184.200 148.200 186.000 149.000 ;
        RECT 185.200 147.600 186.000 148.200 ;
        RECT 332.400 148.200 334.200 149.000 ;
        RECT 499.400 148.200 501.200 149.000 ;
        RECT 332.400 147.600 333.200 148.200 ;
        RECT 500.400 147.600 501.200 148.200 ;
        RECT 498.800 133.800 499.600 134.400 ;
        RECT 498.800 133.000 500.600 133.800 ;
      LAYER via1 ;
        RECT 97.200 413.600 98.000 414.400 ;
        RECT 314.800 413.600 315.600 414.400 ;
        RECT 198.000 333.600 198.800 334.400 ;
        RECT 495.600 293.600 496.400 294.400 ;
        RECT 110.000 213.600 110.800 214.400 ;
        RECT 252.400 173.600 253.200 174.400 ;
        RECT 498.800 133.600 499.600 134.400 ;
      LAYER metal2 ;
        RECT 97.300 420.400 97.900 424.300 ;
        RECT 97.200 419.600 98.000 420.400 ;
        RECT 97.300 414.400 97.900 419.600 ;
        RECT 314.800 417.600 315.600 418.400 ;
        RECT 388.400 417.600 389.200 418.400 ;
        RECT 314.900 414.400 315.500 417.600 ;
        RECT 97.200 413.600 98.000 414.400 ;
        RECT 314.800 413.600 315.600 414.400 ;
        RECT 388.500 388.400 389.100 417.600 ;
        RECT 388.400 387.600 389.200 388.400 ;
        RECT 388.500 356.400 389.100 387.600 ;
        RECT 388.400 355.600 389.200 356.400 ;
        RECT 500.400 355.600 501.200 356.400 ;
        RECT 500.500 348.400 501.100 355.600 ;
        RECT 500.400 347.600 501.200 348.400 ;
        RECT 198.000 333.600 198.800 334.400 ;
        RECT 198.100 332.400 198.700 333.600 ;
        RECT 198.000 331.600 198.800 332.400 ;
        RECT 495.600 293.600 496.400 294.400 ;
        RECT 495.700 272.400 496.300 293.600 ;
        RECT 495.600 271.600 496.400 272.400 ;
        RECT 183.600 227.600 184.400 228.400 ;
        RECT 183.700 226.400 184.300 227.600 ;
        RECT 110.000 225.600 110.800 226.400 ;
        RECT 183.600 225.600 184.400 226.400 ;
        RECT 110.100 214.400 110.700 225.600 ;
        RECT 110.000 213.600 110.800 214.400 ;
        RECT 252.400 179.600 253.200 180.400 ;
        RECT 252.500 174.400 253.100 179.600 ;
        RECT 252.400 173.600 253.200 174.400 ;
        RECT 185.200 169.600 186.000 170.400 ;
        RECT 185.300 148.400 185.900 169.600 ;
        RECT 252.500 152.400 253.100 173.600 ;
        RECT 252.400 151.600 253.200 152.400 ;
        RECT 332.400 151.600 333.200 152.400 ;
        RECT 332.500 148.400 333.100 151.600 ;
        RECT 185.200 147.600 186.000 148.400 ;
        RECT 332.400 147.600 333.200 148.400 ;
        RECT 498.800 147.600 499.600 148.400 ;
        RECT 500.400 147.600 501.200 148.400 ;
        RECT 498.900 134.400 499.500 147.600 ;
        RECT 498.800 133.600 499.600 134.400 ;
      LAYER metal3 ;
        RECT 97.200 420.300 98.000 420.400 ;
        RECT 194.800 420.300 195.600 420.400 ;
        RECT 97.200 419.700 195.600 420.300 ;
        RECT 97.200 419.600 98.000 419.700 ;
        RECT 194.800 419.600 195.600 419.700 ;
        RECT 194.900 418.300 195.500 419.600 ;
        RECT 314.800 418.300 315.600 418.400 ;
        RECT 388.400 418.300 389.200 418.400 ;
        RECT 194.900 417.700 389.200 418.300 ;
        RECT 314.800 417.600 315.600 417.700 ;
        RECT 388.400 417.600 389.200 417.700 ;
        RECT 388.400 356.300 389.200 356.400 ;
        RECT 492.400 356.300 493.200 356.400 ;
        RECT 500.400 356.300 501.200 356.400 ;
        RECT 388.400 355.700 501.200 356.300 ;
        RECT 388.400 355.600 389.200 355.700 ;
        RECT 492.400 355.600 493.200 355.700 ;
        RECT 500.400 355.600 501.200 355.700 ;
        RECT 194.800 332.300 195.600 332.400 ;
        RECT 198.000 332.300 198.800 332.400 ;
        RECT 194.800 331.700 198.800 332.300 ;
        RECT 194.800 331.600 195.600 331.700 ;
        RECT 198.000 331.600 198.800 331.700 ;
        RECT 492.400 294.300 493.200 294.400 ;
        RECT 495.600 294.300 496.400 294.400 ;
        RECT 492.400 293.700 496.400 294.300 ;
        RECT 492.400 293.600 493.200 293.700 ;
        RECT 495.600 293.600 496.400 293.700 ;
        RECT 495.600 272.300 496.400 272.400 ;
        RECT 498.800 272.300 499.600 272.400 ;
        RECT 495.600 271.700 499.600 272.300 ;
        RECT 495.600 271.600 496.400 271.700 ;
        RECT 498.800 271.600 499.600 271.700 ;
        RECT 110.000 226.300 110.800 226.400 ;
        RECT 182.000 226.300 182.800 226.400 ;
        RECT 183.600 226.300 184.400 226.400 ;
        RECT 194.800 226.300 195.600 226.400 ;
        RECT 110.000 225.700 195.600 226.300 ;
        RECT 110.000 225.600 110.800 225.700 ;
        RECT 182.000 225.600 182.800 225.700 ;
        RECT 183.600 225.600 184.400 225.700 ;
        RECT 194.800 225.600 195.600 225.700 ;
        RECT 182.000 180.300 182.800 180.400 ;
        RECT 252.400 180.300 253.200 180.400 ;
        RECT 182.000 179.700 253.200 180.300 ;
        RECT 182.000 179.600 182.800 179.700 ;
        RECT 252.400 179.600 253.200 179.700 ;
        RECT 182.000 170.300 182.800 170.400 ;
        RECT 185.200 170.300 186.000 170.400 ;
        RECT 182.000 169.700 186.000 170.300 ;
        RECT 182.000 169.600 182.800 169.700 ;
        RECT 185.200 169.600 186.000 169.700 ;
        RECT 252.400 152.300 253.200 152.400 ;
        RECT 332.400 152.300 333.200 152.400 ;
        RECT 252.400 151.700 333.200 152.300 ;
        RECT 252.400 151.600 253.200 151.700 ;
        RECT 332.400 151.600 333.200 151.700 ;
        RECT 498.800 148.300 499.600 148.400 ;
        RECT 500.400 148.300 501.200 148.400 ;
        RECT 498.800 147.700 501.200 148.300 ;
        RECT 498.800 147.600 499.600 147.700 ;
        RECT 500.400 147.600 501.200 147.700 ;
      LAYER metal4 ;
        RECT 181.800 169.400 183.000 226.600 ;
        RECT 194.600 225.400 195.800 420.600 ;
        RECT 492.200 293.400 493.400 356.600 ;
        RECT 498.600 147.400 499.800 272.600 ;
    END
  END clk
  PIN rst
    PORT
      LAYER metal1 ;
        RECT 393.200 413.600 394.000 415.200 ;
        RECT 439.600 413.600 440.400 415.200 ;
        RECT 500.400 413.600 501.200 415.200 ;
        RECT 433.200 386.800 434.000 388.400 ;
        RECT 481.200 386.800 482.000 388.400 ;
        RECT 492.400 386.800 493.200 388.400 ;
        RECT 532.400 374.300 533.200 374.400 ;
        RECT 534.000 374.300 534.800 375.200 ;
        RECT 532.400 373.700 534.800 374.300 ;
        RECT 532.400 373.600 533.200 373.700 ;
        RECT 534.000 373.600 534.800 373.700 ;
        RECT 537.200 306.800 538.000 308.400 ;
        RECT 569.200 293.600 570.000 295.200 ;
      LAYER via1 ;
        RECT 433.200 387.600 434.000 388.400 ;
        RECT 481.200 387.600 482.000 388.400 ;
        RECT 492.400 387.600 493.200 388.400 ;
        RECT 537.200 307.600 538.000 308.400 ;
      LAYER metal2 ;
        RECT 393.300 418.400 393.900 424.300 ;
        RECT 393.200 417.600 394.000 418.400 ;
        RECT 439.600 417.600 440.400 418.400 ;
        RECT 393.300 414.400 393.900 417.600 ;
        RECT 439.700 414.400 440.300 417.600 ;
        RECT 393.200 413.600 394.000 414.400 ;
        RECT 439.600 413.600 440.400 414.400 ;
        RECT 500.400 413.600 501.200 414.400 ;
        RECT 433.200 387.600 434.000 388.400 ;
        RECT 433.300 382.400 433.900 387.600 ;
        RECT 439.700 382.400 440.300 413.600 ;
        RECT 481.200 387.600 482.000 388.400 ;
        RECT 492.400 387.600 493.200 388.400 ;
        RECT 481.300 382.400 481.900 387.600 ;
        RECT 492.500 382.400 493.100 387.600 ;
        RECT 500.500 382.400 501.100 413.600 ;
        RECT 433.200 381.600 434.000 382.400 ;
        RECT 439.600 381.600 440.400 382.400 ;
        RECT 481.200 381.600 482.000 382.400 ;
        RECT 492.400 381.600 493.200 382.400 ;
        RECT 500.400 381.600 501.200 382.400 ;
        RECT 532.400 381.600 533.200 382.400 ;
        RECT 532.500 374.400 533.100 381.600 ;
        RECT 532.400 373.600 533.200 374.400 ;
        RECT 537.200 307.600 538.000 308.400 ;
        RECT 537.300 306.400 537.900 307.600 ;
        RECT 537.200 305.600 538.000 306.400 ;
        RECT 537.300 296.400 537.900 305.600 ;
        RECT 537.200 295.600 538.000 296.400 ;
        RECT 569.200 295.600 570.000 296.400 ;
        RECT 569.300 294.400 569.900 295.600 ;
        RECT 569.200 293.600 570.000 294.400 ;
      LAYER metal3 ;
        RECT 393.200 418.300 394.000 418.400 ;
        RECT 439.600 418.300 440.400 418.400 ;
        RECT 393.200 417.700 440.400 418.300 ;
        RECT 393.200 417.600 394.000 417.700 ;
        RECT 439.600 417.600 440.400 417.700 ;
        RECT 433.200 382.300 434.000 382.400 ;
        RECT 439.600 382.300 440.400 382.400 ;
        RECT 481.200 382.300 482.000 382.400 ;
        RECT 492.400 382.300 493.200 382.400 ;
        RECT 500.400 382.300 501.200 382.400 ;
        RECT 532.400 382.300 533.200 382.400 ;
        RECT 534.000 382.300 534.800 382.400 ;
        RECT 433.200 381.700 534.800 382.300 ;
        RECT 433.200 381.600 434.000 381.700 ;
        RECT 439.600 381.600 440.400 381.700 ;
        RECT 481.200 381.600 482.000 381.700 ;
        RECT 492.400 381.600 493.200 381.700 ;
        RECT 500.400 381.600 501.200 381.700 ;
        RECT 532.400 381.600 533.200 381.700 ;
        RECT 534.000 381.600 534.800 381.700 ;
        RECT 534.000 306.300 534.800 306.400 ;
        RECT 537.200 306.300 538.000 306.400 ;
        RECT 534.000 305.700 538.000 306.300 ;
        RECT 534.000 305.600 534.800 305.700 ;
        RECT 537.200 305.600 538.000 305.700 ;
        RECT 537.200 296.300 538.000 296.400 ;
        RECT 569.200 296.300 570.000 296.400 ;
        RECT 537.200 295.700 570.000 296.300 ;
        RECT 537.200 295.600 538.000 295.700 ;
        RECT 569.200 295.600 570.000 295.700 ;
      LAYER metal4 ;
        RECT 533.800 305.400 535.000 382.600 ;
    END
  END rst
  PIN theta[0]
    PORT
      LAYER metal1 ;
        RECT 554.800 293.600 555.600 295.200 ;
        RECT 577.000 294.300 578.000 294.400 ;
        RECT 578.800 294.300 579.600 294.400 ;
        RECT 577.000 293.700 579.600 294.300 ;
        RECT 577.000 293.600 578.000 293.700 ;
        RECT 578.800 293.600 579.600 293.700 ;
        RECT 576.800 292.800 577.600 293.600 ;
        RECT 572.400 288.800 573.200 290.400 ;
      LAYER via1 ;
        RECT 572.400 289.600 573.200 290.400 ;
      LAYER metal2 ;
        RECT 554.800 293.600 555.600 294.400 ;
        RECT 572.400 293.600 573.200 294.400 ;
        RECT 578.800 293.600 579.600 294.400 ;
        RECT 572.500 290.400 573.100 293.600 ;
        RECT 572.400 289.600 573.200 290.400 ;
      LAYER metal3 ;
        RECT 554.800 294.300 555.600 294.400 ;
        RECT 572.400 294.300 573.200 294.400 ;
        RECT 578.800 294.300 579.600 294.400 ;
        RECT 554.800 293.700 589.100 294.300 ;
        RECT 554.800 293.600 555.600 293.700 ;
        RECT 572.400 293.600 573.200 293.700 ;
        RECT 578.800 293.600 579.600 293.700 ;
    END
  END theta[0]
  PIN theta[1]
    PORT
      LAYER metal1 ;
        RECT 534.000 311.600 534.800 313.200 ;
        RECT 541.600 308.400 542.400 309.200 ;
        RECT 519.600 306.800 520.400 308.400 ;
        RECT 541.800 307.600 542.800 308.400 ;
      LAYER via1 ;
        RECT 519.600 307.600 520.400 308.400 ;
        RECT 542.000 307.600 542.800 308.400 ;
      LAYER metal2 ;
        RECT 534.000 311.600 534.800 312.400 ;
        RECT 534.100 308.400 534.700 311.600 ;
        RECT 519.600 307.600 520.400 308.400 ;
        RECT 534.000 307.600 534.800 308.400 ;
        RECT 542.000 307.600 542.800 308.400 ;
      LAYER metal3 ;
        RECT 542.100 309.700 589.100 310.300 ;
        RECT 542.100 308.400 542.700 309.700 ;
        RECT 519.600 308.300 520.400 308.400 ;
        RECT 534.000 308.300 534.800 308.400 ;
        RECT 542.000 308.300 542.800 308.400 ;
        RECT 519.600 307.700 542.800 308.300 ;
        RECT 519.600 307.600 520.400 307.700 ;
        RECT 534.000 307.600 534.800 307.700 ;
        RECT 542.000 307.600 542.800 307.700 ;
    END
  END theta[1]
  PIN theta[2]
    PORT
      LAYER metal1 ;
        RECT 478.000 391.600 478.800 393.200 ;
        RECT 485.600 388.400 486.400 389.200 ;
        RECT 463.600 386.800 464.400 388.400 ;
        RECT 485.800 387.600 486.800 388.400 ;
      LAYER via1 ;
        RECT 463.600 387.600 464.400 388.400 ;
        RECT 486.000 387.600 486.800 388.400 ;
      LAYER metal2 ;
        RECT 478.100 420.400 478.700 424.300 ;
        RECT 478.000 419.600 478.800 420.400 ;
        RECT 463.600 391.600 464.400 392.400 ;
        RECT 478.000 391.600 478.800 392.400 ;
        RECT 486.000 391.600 486.800 392.400 ;
        RECT 463.700 388.400 464.300 391.600 ;
        RECT 486.100 388.400 486.700 391.600 ;
        RECT 463.600 387.600 464.400 388.400 ;
        RECT 486.000 387.600 486.800 388.400 ;
      LAYER metal3 ;
        RECT 476.400 420.300 477.200 420.400 ;
        RECT 478.000 420.300 478.800 420.400 ;
        RECT 476.400 419.700 478.800 420.300 ;
        RECT 476.400 419.600 477.200 419.700 ;
        RECT 478.000 419.600 478.800 419.700 ;
        RECT 463.600 392.300 464.400 392.400 ;
        RECT 476.400 392.300 477.200 392.400 ;
        RECT 478.000 392.300 478.800 392.400 ;
        RECT 486.000 392.300 486.800 392.400 ;
        RECT 463.600 391.700 486.800 392.300 ;
        RECT 463.600 391.600 464.400 391.700 ;
        RECT 476.400 391.600 477.200 391.700 ;
        RECT 478.000 391.600 478.800 391.700 ;
        RECT 486.000 391.600 486.800 391.700 ;
      LAYER metal4 ;
        RECT 476.200 391.400 477.400 420.600 ;
    END
  END theta[2]
  PIN theta[3]
    PORT
      LAYER metal1 ;
        RECT 422.000 413.600 422.800 415.200 ;
        RECT 449.000 413.600 450.000 414.400 ;
        RECT 448.800 412.800 449.600 413.600 ;
        RECT 436.400 408.800 437.200 410.400 ;
      LAYER via1 ;
        RECT 449.200 413.600 450.000 414.400 ;
        RECT 436.400 409.600 437.200 410.400 ;
      LAYER metal2 ;
        RECT 422.100 414.400 422.700 424.300 ;
        RECT 422.000 413.600 422.800 414.400 ;
        RECT 449.200 413.600 450.000 414.400 ;
        RECT 422.100 410.400 422.700 413.600 ;
        RECT 449.300 410.400 449.900 413.600 ;
        RECT 422.000 409.600 422.800 410.400 ;
        RECT 436.400 409.600 437.200 410.400 ;
        RECT 449.200 409.600 450.000 410.400 ;
      LAYER metal3 ;
        RECT 422.000 410.300 422.800 410.400 ;
        RECT 436.400 410.300 437.200 410.400 ;
        RECT 449.200 410.300 450.000 410.400 ;
        RECT 422.000 409.700 450.000 410.300 ;
        RECT 422.000 409.600 422.800 409.700 ;
        RECT 436.400 409.600 437.200 409.700 ;
        RECT 449.200 409.600 450.000 409.700 ;
    END
  END theta[3]
  PIN theta[4]
    PORT
      LAYER metal1 ;
        RECT 489.200 391.600 490.000 393.200 ;
        RECT 478.000 373.600 478.800 375.200 ;
        RECT 495.400 373.600 496.400 374.400 ;
        RECT 495.200 372.800 496.000 373.600 ;
      LAYER via1 ;
        RECT 495.600 373.600 496.400 374.400 ;
      LAYER metal2 ;
        RECT 489.300 392.400 489.900 424.300 ;
        RECT 489.200 391.600 490.000 392.400 ;
        RECT 489.300 374.400 489.900 391.600 ;
        RECT 478.000 373.600 478.800 374.400 ;
        RECT 489.200 373.600 490.000 374.400 ;
        RECT 495.600 373.600 496.400 374.400 ;
      LAYER metal3 ;
        RECT 478.000 374.300 478.800 374.400 ;
        RECT 489.200 374.300 490.000 374.400 ;
        RECT 495.600 374.300 496.400 374.400 ;
        RECT 478.000 373.700 496.400 374.300 ;
        RECT 478.000 373.600 478.800 373.700 ;
        RECT 489.200 373.600 490.000 373.700 ;
        RECT 495.600 373.600 496.400 373.700 ;
    END
  END theta[4]
  PIN theta[5]
    PORT
      LAYER metal1 ;
        RECT 482.800 413.600 483.600 415.200 ;
        RECT 505.000 413.600 506.000 414.400 ;
        RECT 504.800 412.800 505.600 413.600 ;
        RECT 497.200 408.800 498.000 410.400 ;
      LAYER via1 ;
        RECT 505.200 413.600 506.000 414.400 ;
        RECT 497.200 409.600 498.000 410.400 ;
      LAYER metal2 ;
        RECT 482.900 414.400 483.500 424.300 ;
        RECT 482.800 413.600 483.600 414.400 ;
        RECT 505.200 413.600 506.000 414.400 ;
        RECT 482.900 410.400 483.500 413.600 ;
        RECT 505.300 410.400 505.900 413.600 ;
        RECT 482.800 409.600 483.600 410.400 ;
        RECT 497.200 409.600 498.000 410.400 ;
        RECT 505.200 409.600 506.000 410.400 ;
      LAYER metal3 ;
        RECT 482.800 410.300 483.600 410.400 ;
        RECT 497.200 410.300 498.000 410.400 ;
        RECT 505.200 410.300 506.000 410.400 ;
        RECT 482.800 409.700 506.000 410.300 ;
        RECT 482.800 409.600 483.600 409.700 ;
        RECT 497.200 409.600 498.000 409.700 ;
        RECT 505.200 409.600 506.000 409.700 ;
    END
  END theta[5]
  PIN theta[6]
    PORT
      LAYER metal1 ;
        RECT 436.400 392.300 437.200 393.200 ;
        RECT 438.000 392.300 438.800 392.400 ;
        RECT 436.400 391.700 438.800 392.300 ;
        RECT 436.400 391.600 437.200 391.700 ;
        RECT 438.000 391.600 438.800 391.700 ;
        RECT 431.600 373.600 432.400 375.200 ;
        RECT 453.800 373.600 454.800 374.400 ;
        RECT 453.600 372.800 454.400 373.600 ;
      LAYER via1 ;
        RECT 454.000 373.600 454.800 374.400 ;
      LAYER metal2 ;
        RECT 438.100 392.400 438.700 424.300 ;
        RECT 438.000 391.600 438.800 392.400 ;
        RECT 438.100 374.400 438.700 391.600 ;
        RECT 431.600 373.600 432.400 374.400 ;
        RECT 438.000 373.600 438.800 374.400 ;
        RECT 454.000 373.600 454.800 374.400 ;
      LAYER metal3 ;
        RECT 431.600 374.300 432.400 374.400 ;
        RECT 438.000 374.300 438.800 374.400 ;
        RECT 454.000 374.300 454.800 374.400 ;
        RECT 431.600 373.700 454.800 374.300 ;
        RECT 431.600 373.600 432.400 373.700 ;
        RECT 438.000 373.600 438.800 373.700 ;
        RECT 454.000 373.600 454.800 373.700 ;
    END
  END theta[6]
  PIN theta[7]
    PORT
      LAYER metal1 ;
        RECT 375.600 413.600 376.400 415.200 ;
        RECT 397.800 413.600 398.800 414.400 ;
        RECT 397.600 412.800 398.400 413.600 ;
        RECT 390.000 408.800 390.800 410.400 ;
      LAYER via1 ;
        RECT 398.000 413.600 398.800 414.400 ;
        RECT 390.000 409.600 390.800 410.400 ;
      LAYER metal2 ;
        RECT 375.700 414.400 376.300 424.300 ;
        RECT 375.600 413.600 376.400 414.400 ;
        RECT 398.000 413.600 398.800 414.400 ;
        RECT 375.700 410.400 376.300 413.600 ;
        RECT 398.100 410.400 398.700 413.600 ;
        RECT 375.600 409.600 376.400 410.400 ;
        RECT 390.000 409.600 390.800 410.400 ;
        RECT 398.000 409.600 398.800 410.400 ;
      LAYER metal3 ;
        RECT 375.600 410.300 376.400 410.400 ;
        RECT 390.000 410.300 390.800 410.400 ;
        RECT 398.000 410.300 398.800 410.400 ;
        RECT 375.600 409.700 398.800 410.300 ;
        RECT 375.600 409.600 376.400 409.700 ;
        RECT 390.000 409.600 390.800 409.700 ;
        RECT 398.000 409.600 398.800 409.700 ;
    END
  END theta[7]
  PIN sine[0]
    PORT
      LAYER metal1 ;
        RECT 506.800 391.800 507.600 399.800 ;
        RECT 506.800 389.600 507.400 391.800 ;
        RECT 506.800 382.200 507.600 389.600 ;
      LAYER via1 ;
        RECT 506.800 397.600 507.600 398.400 ;
      LAYER metal2 ;
        RECT 508.500 414.300 509.100 424.300 ;
        RECT 506.900 413.700 509.100 414.300 ;
        RECT 506.900 398.400 507.500 413.700 ;
        RECT 506.800 397.600 507.600 398.400 ;
    END
  END sine[0]
  PIN sine[1]
    PORT
      LAYER metal1 ;
        RECT 559.600 252.400 560.400 259.800 ;
        RECT 559.800 250.200 560.400 252.400 ;
        RECT 559.600 242.200 560.400 250.200 ;
      LAYER via1 ;
        RECT 559.600 247.600 560.400 248.400 ;
      LAYER metal2 ;
        RECT 559.600 249.600 560.400 250.400 ;
        RECT 559.700 248.400 560.300 249.600 ;
        RECT 559.600 247.600 560.400 248.400 ;
      LAYER metal3 ;
        RECT 559.600 250.300 560.400 250.400 ;
        RECT 559.600 249.700 589.100 250.300 ;
        RECT 559.600 249.600 560.400 249.700 ;
    END
  END sine[1]
  PIN sine[2]
    PORT
      LAYER metal1 ;
        RECT 580.400 238.300 581.200 239.800 ;
        RECT 585.200 238.300 586.000 238.400 ;
        RECT 580.400 237.700 586.000 238.300 ;
        RECT 580.400 231.800 581.200 237.700 ;
        RECT 585.200 237.600 586.000 237.700 ;
        RECT 580.600 229.600 581.200 231.800 ;
        RECT 580.400 222.200 581.200 229.600 ;
      LAYER metal2 ;
        RECT 585.200 237.600 586.000 238.400 ;
      LAYER metal3 ;
        RECT 585.200 238.300 586.000 238.400 ;
        RECT 585.200 237.700 589.100 238.300 ;
        RECT 585.200 237.600 586.000 237.700 ;
    END
  END sine[2]
  PIN sine[3]
    PORT
      LAYER metal1 ;
        RECT 532.400 231.800 533.200 239.800 ;
        RECT 532.600 229.600 533.200 231.800 ;
        RECT 532.400 222.200 533.200 229.600 ;
      LAYER via1 ;
        RECT 532.400 233.600 533.200 234.400 ;
      LAYER metal2 ;
        RECT 532.400 233.600 533.200 234.400 ;
      LAYER metal3 ;
        RECT 532.400 234.300 533.200 234.400 ;
        RECT 532.400 233.700 589.100 234.300 ;
        RECT 532.400 233.600 533.200 233.700 ;
    END
  END sine[3]
  PIN sine[4]
    PORT
      LAYER metal1 ;
        RECT 460.400 412.400 461.200 419.800 ;
        RECT 460.600 410.200 461.200 412.400 ;
        RECT 460.400 402.200 461.200 410.200 ;
      LAYER via1 ;
        RECT 460.400 417.600 461.200 418.400 ;
      LAYER metal2 ;
        RECT 458.900 423.700 461.100 424.300 ;
        RECT 460.500 418.400 461.100 423.700 ;
        RECT 460.400 417.600 461.200 418.400 ;
    END
  END sine[4]
  PIN sine[5]
    PORT
      LAYER metal1 ;
        RECT 583.600 292.400 584.400 299.800 ;
        RECT 583.800 290.200 584.400 292.400 ;
        RECT 583.600 288.300 584.400 290.200 ;
        RECT 585.200 288.300 586.000 288.400 ;
        RECT 583.600 287.700 586.000 288.300 ;
        RECT 583.600 282.200 584.400 287.700 ;
        RECT 585.200 287.600 586.000 287.700 ;
      LAYER metal2 ;
        RECT 585.200 289.600 586.000 290.400 ;
        RECT 585.300 288.400 585.900 289.600 ;
        RECT 585.200 287.600 586.000 288.400 ;
      LAYER metal3 ;
        RECT 585.200 290.300 586.000 290.400 ;
        RECT 585.200 289.700 589.100 290.300 ;
        RECT 585.200 289.600 586.000 289.700 ;
    END
  END sine[5]
  PIN sine[6]
    PORT
      LAYER metal1 ;
        RECT 585.200 212.400 586.000 219.800 ;
        RECT 585.400 210.200 586.000 212.400 ;
        RECT 585.200 202.200 586.000 210.200 ;
      LAYER via1 ;
        RECT 585.200 207.600 586.000 208.400 ;
      LAYER metal2 ;
        RECT 585.200 209.600 586.000 210.400 ;
        RECT 585.300 208.400 585.900 209.600 ;
        RECT 585.200 207.600 586.000 208.400 ;
      LAYER metal3 ;
        RECT 585.200 210.300 586.000 210.400 ;
        RECT 585.200 209.700 589.100 210.300 ;
        RECT 585.200 209.600 586.000 209.700 ;
    END
  END sine[6]
  PIN sine[7]
    PORT
      LAYER metal1 ;
        RECT 583.600 271.800 584.400 279.800 ;
        RECT 583.800 269.600 584.400 271.800 ;
        RECT 583.600 268.300 584.400 269.600 ;
        RECT 585.200 268.300 586.000 268.400 ;
        RECT 583.600 267.700 586.000 268.300 ;
        RECT 583.600 262.200 584.400 267.700 ;
        RECT 585.200 267.600 586.000 267.700 ;
      LAYER metal2 ;
        RECT 585.200 269.600 586.000 270.400 ;
        RECT 585.300 268.400 585.900 269.600 ;
        RECT 585.200 267.600 586.000 268.400 ;
      LAYER metal3 ;
        RECT 585.200 270.300 586.000 270.400 ;
        RECT 585.200 269.700 589.100 270.300 ;
        RECT 585.200 269.600 586.000 269.700 ;
    END
  END sine[7]
  PIN cosine[0]
    PORT
      LAYER metal1 ;
        RECT 583.600 254.300 584.400 259.800 ;
        RECT 585.200 254.300 586.000 254.400 ;
        RECT 583.600 253.700 586.000 254.300 ;
        RECT 583.600 252.400 584.400 253.700 ;
        RECT 585.200 253.600 586.000 253.700 ;
        RECT 583.800 250.200 584.400 252.400 ;
        RECT 583.600 242.200 584.400 250.200 ;
      LAYER metal2 ;
        RECT 585.200 253.600 586.000 254.400 ;
      LAYER metal3 ;
        RECT 585.200 254.300 586.000 254.400 ;
        RECT 585.200 253.700 589.100 254.300 ;
        RECT 585.200 253.600 586.000 253.700 ;
    END
  END cosine[0]
  PIN cosine[1]
    PORT
      LAYER metal1 ;
        RECT 575.600 231.800 576.400 239.800 ;
        RECT 575.800 229.600 576.400 231.800 ;
        RECT 575.600 222.200 576.400 229.600 ;
      LAYER via1 ;
        RECT 575.600 227.600 576.400 228.400 ;
      LAYER metal2 ;
        RECT 575.600 229.600 576.400 230.400 ;
        RECT 575.700 228.400 576.300 229.600 ;
        RECT 575.600 227.600 576.400 228.400 ;
      LAYER metal3 ;
        RECT 575.600 230.300 576.400 230.400 ;
        RECT 575.600 229.700 589.100 230.300 ;
        RECT 575.600 229.600 576.400 229.700 ;
    END
  END cosine[1]
  PIN cosine[2]
    PORT
      LAYER metal1 ;
        RECT 577.200 332.400 578.000 339.800 ;
        RECT 577.400 330.200 578.000 332.400 ;
        RECT 577.200 322.200 578.000 330.200 ;
      LAYER via1 ;
        RECT 577.200 327.600 578.000 328.400 ;
      LAYER metal2 ;
        RECT 577.200 329.600 578.000 330.400 ;
        RECT 577.300 328.400 577.900 329.600 ;
        RECT 577.200 327.600 578.000 328.400 ;
      LAYER metal3 ;
        RECT 577.200 330.300 578.000 330.400 ;
        RECT 577.200 329.700 589.100 330.300 ;
        RECT 577.200 329.600 578.000 329.700 ;
    END
  END cosine[2]
  PIN cosine[3]
    PORT
      LAYER metal1 ;
        RECT 575.600 92.400 576.400 99.800 ;
        RECT 575.800 90.200 576.400 92.400 ;
        RECT 575.600 82.200 576.400 90.200 ;
      LAYER via1 ;
        RECT 575.600 87.600 576.400 88.400 ;
      LAYER metal2 ;
        RECT 575.600 89.600 576.400 90.400 ;
        RECT 575.700 88.400 576.300 89.600 ;
        RECT 575.600 87.600 576.400 88.400 ;
      LAYER metal3 ;
        RECT 575.600 90.300 576.400 90.400 ;
        RECT 575.600 89.700 589.100 90.300 ;
        RECT 575.600 89.600 576.400 89.700 ;
    END
  END cosine[3]
  PIN cosine[4]
    PORT
      LAYER metal1 ;
        RECT 580.400 172.400 581.200 179.800 ;
        RECT 580.600 170.200 581.200 172.400 ;
        RECT 580.400 168.300 581.200 170.200 ;
        RECT 585.200 168.300 586.000 168.400 ;
        RECT 580.400 167.700 586.000 168.300 ;
        RECT 580.400 162.200 581.200 167.700 ;
        RECT 585.200 167.600 586.000 167.700 ;
      LAYER metal2 ;
        RECT 585.200 169.600 586.000 170.400 ;
        RECT 585.300 168.400 585.900 169.600 ;
        RECT 585.200 167.600 586.000 168.400 ;
      LAYER metal3 ;
        RECT 585.200 170.300 586.000 170.400 ;
        RECT 585.200 169.700 589.100 170.300 ;
        RECT 585.200 169.600 586.000 169.700 ;
    END
  END cosine[4]
  PIN cosine[5]
    PORT
      LAYER metal1 ;
        RECT 583.600 71.800 584.400 79.800 ;
        RECT 583.800 69.600 584.400 71.800 ;
        RECT 583.600 68.300 584.400 69.600 ;
        RECT 585.200 68.300 586.000 68.400 ;
        RECT 583.600 67.700 586.000 68.300 ;
        RECT 583.600 62.200 584.400 67.700 ;
        RECT 585.200 67.600 586.000 67.700 ;
      LAYER metal2 ;
        RECT 585.200 69.600 586.000 70.400 ;
        RECT 585.300 68.400 585.900 69.600 ;
        RECT 585.200 67.600 586.000 68.400 ;
      LAYER metal3 ;
        RECT 585.200 70.300 586.000 70.400 ;
        RECT 585.200 69.700 589.100 70.300 ;
        RECT 585.200 69.600 586.000 69.700 ;
    END
  END cosine[5]
  PIN cosine[6]
    PORT
      LAYER metal1 ;
        RECT 580.400 94.300 581.200 99.800 ;
        RECT 585.200 94.300 586.000 94.400 ;
        RECT 580.400 93.700 586.000 94.300 ;
        RECT 580.400 92.400 581.200 93.700 ;
        RECT 585.200 93.600 586.000 93.700 ;
        RECT 580.600 90.200 581.200 92.400 ;
        RECT 580.400 82.200 581.200 90.200 ;
      LAYER metal2 ;
        RECT 585.200 93.600 586.000 94.400 ;
      LAYER metal3 ;
        RECT 585.200 94.300 586.000 94.400 ;
        RECT 585.200 93.700 589.100 94.300 ;
        RECT 585.200 93.600 586.000 93.700 ;
    END
  END cosine[6]
  PIN cosine[7]
    PORT
      LAYER metal1 ;
        RECT 582.000 12.400 582.800 19.800 ;
        RECT 582.200 10.200 582.800 12.400 ;
        RECT 582.000 8.300 582.800 10.200 ;
        RECT 585.200 8.300 586.000 8.400 ;
        RECT 582.000 7.700 586.000 8.300 ;
        RECT 582.000 2.200 582.800 7.700 ;
        RECT 585.200 7.600 586.000 7.700 ;
      LAYER metal2 ;
        RECT 585.200 9.600 586.000 10.400 ;
        RECT 585.300 8.400 585.900 9.600 ;
        RECT 585.200 7.600 586.000 8.400 ;
      LAYER metal3 ;
        RECT 585.200 10.300 586.000 10.400 ;
        RECT 585.200 9.700 589.100 10.300 ;
        RECT 585.200 9.600 586.000 9.700 ;
    END
  END cosine[7]
  PIN done
    PORT
      LAYER metal1 ;
        RECT 582.000 334.300 582.800 339.800 ;
        RECT 585.200 334.300 586.000 334.400 ;
        RECT 582.000 333.700 586.000 334.300 ;
        RECT 582.000 332.400 582.800 333.700 ;
        RECT 585.200 333.600 586.000 333.700 ;
        RECT 582.200 330.200 582.800 332.400 ;
        RECT 582.000 322.200 582.800 330.200 ;
      LAYER metal2 ;
        RECT 585.200 333.600 586.000 334.400 ;
      LAYER metal3 ;
        RECT 585.200 334.300 586.000 334.400 ;
        RECT 585.200 333.700 589.100 334.300 ;
        RECT 585.200 333.600 586.000 333.700 ;
    END
  END done
  OBS
      LAYER metal1 ;
        RECT 1.200 415.800 2.000 419.800 ;
        RECT 2.800 416.000 3.600 419.800 ;
        RECT 6.000 416.000 6.800 419.800 ;
        RECT 2.800 415.800 6.800 416.000 ;
        RECT 1.400 414.400 2.000 415.800 ;
        RECT 3.000 415.400 6.600 415.800 ;
        RECT 5.200 414.400 6.000 414.800 ;
        RECT 1.200 413.600 3.800 414.400 ;
        RECT 5.200 414.300 6.800 414.400 ;
        RECT 7.600 414.300 8.400 419.800 ;
        RECT 12.400 417.800 13.200 419.800 ;
        RECT 9.200 416.300 10.000 417.200 ;
        RECT 10.800 416.300 11.600 417.200 ;
        RECT 9.200 415.700 11.600 416.300 ;
        RECT 9.200 415.600 10.000 415.700 ;
        RECT 10.800 415.600 11.600 415.700 ;
        RECT 12.600 415.600 13.200 417.800 ;
        RECT 15.600 415.800 16.400 419.800 ;
        RECT 19.800 416.400 20.600 419.800 ;
        RECT 12.600 415.000 15.000 415.600 ;
        RECT 5.200 413.800 8.400 414.300 ;
        RECT 6.000 413.700 8.400 413.800 ;
        RECT 6.000 413.600 6.800 413.700 ;
        RECT 3.200 412.400 3.800 413.600 ;
        RECT 2.800 411.600 3.800 412.400 ;
        RECT 4.400 411.600 5.200 413.200 ;
        RECT 1.200 410.200 2.000 410.400 ;
        RECT 3.200 410.200 3.800 411.600 ;
        RECT 1.200 409.600 2.600 410.200 ;
        RECT 3.200 409.600 4.200 410.200 ;
        RECT 2.000 408.400 2.600 409.600 ;
        RECT 2.000 407.600 2.800 408.400 ;
        RECT 3.400 402.200 4.200 409.600 ;
        RECT 7.600 402.200 8.400 413.700 ;
        RECT 9.200 414.300 10.000 414.400 ;
        RECT 12.400 414.300 13.400 414.400 ;
        RECT 9.200 413.700 13.400 414.300 ;
        RECT 9.200 413.600 10.000 413.700 ;
        RECT 12.400 413.600 13.400 413.700 ;
        RECT 12.800 412.800 13.600 413.600 ;
        RECT 14.400 412.000 15.000 415.000 ;
        RECT 15.800 412.400 16.400 415.800 ;
        RECT 18.800 415.800 20.600 416.400 ;
        RECT 22.000 415.800 22.800 419.800 ;
        RECT 23.600 416.000 24.400 419.800 ;
        RECT 26.800 416.000 27.600 419.800 ;
        RECT 30.000 417.800 30.800 419.800 ;
        RECT 23.600 415.800 27.600 416.000 ;
        RECT 17.200 413.600 18.000 415.200 ;
        RECT 14.200 411.400 15.000 412.000 ;
        RECT 15.600 411.600 16.400 412.400 ;
        RECT 10.800 411.200 15.000 411.400 ;
        RECT 10.800 410.800 14.800 411.200 ;
        RECT 10.800 402.200 11.600 410.800 ;
        RECT 15.800 410.200 16.400 411.600 ;
        RECT 15.000 409.600 16.400 410.200 ;
        RECT 18.800 412.300 19.600 415.800 ;
        RECT 22.200 414.400 22.800 415.800 ;
        RECT 23.800 415.400 27.400 415.800 ;
        RECT 28.400 415.600 29.200 417.200 ;
        RECT 26.000 414.400 26.800 414.800 ;
        RECT 30.200 414.400 30.800 417.800 ;
        RECT 33.200 416.000 34.000 419.800 ;
        RECT 36.400 416.000 37.200 419.800 ;
        RECT 33.200 415.800 37.200 416.000 ;
        RECT 38.000 415.800 38.800 419.800 ;
        RECT 40.200 418.400 41.000 419.800 ;
        RECT 39.600 417.600 41.000 418.400 ;
        RECT 40.200 416.800 41.000 417.600 ;
        RECT 39.600 415.800 41.000 416.800 ;
        RECT 44.400 415.800 45.200 419.800 ;
        RECT 33.400 415.400 37.000 415.800 ;
        RECT 34.000 414.400 34.800 414.800 ;
        RECT 38.000 414.400 38.600 415.800 ;
        RECT 22.000 413.600 24.600 414.400 ;
        RECT 26.000 413.800 27.600 414.400 ;
        RECT 26.800 413.600 27.600 413.800 ;
        RECT 30.000 414.300 30.800 414.400 ;
        RECT 33.200 414.300 34.800 414.400 ;
        RECT 30.000 413.800 34.800 414.300 ;
        RECT 30.000 413.700 34.000 413.800 ;
        RECT 30.000 413.600 30.800 413.700 ;
        RECT 33.200 413.600 34.000 413.700 ;
        RECT 36.200 413.600 38.800 414.400 ;
        RECT 24.000 412.400 24.600 413.600 ;
        RECT 18.800 411.700 22.700 412.300 ;
        RECT 15.000 404.400 15.800 409.600 ;
        RECT 15.000 403.600 16.400 404.400 ;
        RECT 15.000 402.200 15.800 403.600 ;
        RECT 18.800 402.200 19.600 411.700 ;
        RECT 22.100 410.400 22.700 411.700 ;
        RECT 23.600 411.600 24.600 412.400 ;
        RECT 25.200 412.300 26.000 413.200 ;
        RECT 30.200 412.300 30.800 413.600 ;
        RECT 25.200 411.700 30.800 412.300 ;
        RECT 25.200 411.600 26.000 411.700 ;
        RECT 20.400 408.800 21.200 410.400 ;
        RECT 22.000 410.200 22.800 410.400 ;
        RECT 24.000 410.200 24.600 411.600 ;
        RECT 30.200 410.200 30.800 411.700 ;
        RECT 31.600 410.800 32.400 412.400 ;
        RECT 34.800 411.600 35.600 413.200 ;
        RECT 36.200 410.400 36.800 413.600 ;
        RECT 39.600 412.400 40.200 415.800 ;
        RECT 44.400 415.600 45.000 415.800 ;
        RECT 43.200 415.200 45.000 415.600 ;
        RECT 40.800 415.000 45.000 415.200 ;
        RECT 46.000 415.400 46.800 419.800 ;
        RECT 50.200 418.400 51.400 419.800 ;
        RECT 50.200 417.800 51.600 418.400 ;
        RECT 54.800 417.800 55.600 419.800 ;
        RECT 59.200 418.400 60.000 419.800 ;
        RECT 59.200 417.800 61.200 418.400 ;
        RECT 50.800 417.000 51.600 417.800 ;
        RECT 55.000 417.200 55.600 417.800 ;
        RECT 55.000 416.600 57.800 417.200 ;
        RECT 57.000 416.400 57.800 416.600 ;
        RECT 58.800 416.400 59.600 417.200 ;
        RECT 60.400 417.000 61.200 417.800 ;
        RECT 49.000 415.400 49.800 415.600 ;
        RECT 40.800 414.600 43.800 415.000 ;
        RECT 46.000 414.800 49.800 415.400 ;
        RECT 40.800 414.400 41.600 414.600 ;
        RECT 39.600 411.600 40.400 412.400 ;
        RECT 22.000 409.600 23.400 410.200 ;
        RECT 24.000 409.600 25.000 410.200 ;
        RECT 22.800 408.400 23.400 409.600 ;
        RECT 22.000 407.600 23.600 408.400 ;
        RECT 24.200 402.200 25.000 409.600 ;
        RECT 30.000 409.400 31.800 410.200 ;
        RECT 34.800 409.600 36.800 410.400 ;
        RECT 38.000 410.200 38.800 410.400 ;
        RECT 37.400 409.600 38.800 410.200 ;
        RECT 39.600 410.200 40.200 411.600 ;
        RECT 41.000 411.000 41.600 414.400 ;
        RECT 42.400 413.800 43.200 414.000 ;
        RECT 42.400 413.200 43.400 413.800 ;
        RECT 42.800 412.400 43.400 413.200 ;
        RECT 44.400 412.800 45.200 414.400 ;
        RECT 42.800 411.600 43.600 412.400 ;
        RECT 46.000 411.400 46.800 414.800 ;
        RECT 53.000 414.200 53.800 414.400 ;
        RECT 58.800 414.200 59.400 416.400 ;
        RECT 63.600 415.000 64.400 419.800 ;
        RECT 65.200 415.400 66.000 419.800 ;
        RECT 69.400 418.400 70.600 419.800 ;
        RECT 69.400 417.800 70.800 418.400 ;
        RECT 74.000 417.800 74.800 419.800 ;
        RECT 78.400 418.400 79.200 419.800 ;
        RECT 78.400 417.800 80.400 418.400 ;
        RECT 70.000 417.000 70.800 417.800 ;
        RECT 74.200 417.200 74.800 417.800 ;
        RECT 74.200 416.600 77.000 417.200 ;
        RECT 76.200 416.400 77.000 416.600 ;
        RECT 78.000 416.400 78.800 417.200 ;
        RECT 79.600 417.000 80.400 417.800 ;
        RECT 68.200 415.400 69.000 415.600 ;
        RECT 65.200 414.800 69.000 415.400 ;
        RECT 62.000 414.200 63.600 414.400 ;
        RECT 52.600 413.600 63.600 414.200 ;
        RECT 50.800 412.800 51.600 413.000 ;
        RECT 47.800 412.200 51.600 412.800 ;
        RECT 47.800 412.000 48.600 412.200 ;
        RECT 49.400 411.400 50.200 411.600 ;
        RECT 41.000 410.400 43.400 411.000 ;
        RECT 31.000 402.200 31.800 409.400 ;
        RECT 35.800 402.200 36.600 409.600 ;
        RECT 37.400 408.400 38.000 409.600 ;
        RECT 37.200 407.600 38.000 408.400 ;
        RECT 39.600 402.200 40.400 410.200 ;
        RECT 42.800 406.200 43.400 410.400 ;
        RECT 46.000 410.800 50.200 411.400 ;
        RECT 42.800 402.200 43.600 406.200 ;
        RECT 46.000 402.200 46.800 410.800 ;
        RECT 52.600 410.400 53.200 413.600 ;
        RECT 59.800 413.400 60.600 413.600 ;
        RECT 58.800 412.400 59.600 412.600 ;
        RECT 61.400 412.400 62.200 412.600 ;
        RECT 57.200 411.800 62.200 412.400 ;
        RECT 57.200 411.600 58.000 411.800 ;
        RECT 65.200 411.400 66.000 414.800 ;
        RECT 72.200 414.200 73.000 414.400 ;
        RECT 78.000 414.200 78.600 416.400 ;
        RECT 82.800 415.000 83.600 419.800 ;
        RECT 86.000 415.200 86.800 419.800 ;
        RECT 89.200 415.200 90.000 419.800 ;
        RECT 92.400 415.200 93.200 419.800 ;
        RECT 95.600 415.200 96.400 419.800 ;
        RECT 101.400 416.400 102.200 419.800 ;
        RECT 100.400 415.800 102.200 416.400 ;
        RECT 84.400 414.400 86.800 415.200 ;
        RECT 87.800 414.400 90.000 415.200 ;
        RECT 91.000 414.400 93.200 415.200 ;
        RECT 94.600 414.400 96.400 415.200 ;
        RECT 81.200 414.200 82.800 414.400 ;
        RECT 71.800 413.600 82.800 414.200 ;
        RECT 70.000 412.800 70.800 413.000 ;
        RECT 67.000 412.200 70.800 412.800 ;
        RECT 67.000 412.000 67.800 412.200 ;
        RECT 68.600 411.400 69.400 411.600 ;
        RECT 58.800 411.000 64.400 411.200 ;
        RECT 58.600 410.800 64.400 411.000 ;
        RECT 50.800 409.800 53.200 410.400 ;
        RECT 54.600 410.600 64.400 410.800 ;
        RECT 54.600 410.200 59.400 410.600 ;
        RECT 50.800 408.800 51.400 409.800 ;
        RECT 50.000 408.000 51.400 408.800 ;
        RECT 53.000 409.000 53.800 409.200 ;
        RECT 54.600 409.000 55.200 410.200 ;
        RECT 53.000 408.400 55.200 409.000 ;
        RECT 55.800 409.000 61.200 409.600 ;
        RECT 55.800 408.800 56.600 409.000 ;
        RECT 60.400 408.800 61.200 409.000 ;
        RECT 54.200 407.400 55.000 407.600 ;
        RECT 57.000 407.400 57.800 407.600 ;
        RECT 50.800 406.200 51.600 407.000 ;
        RECT 54.200 406.800 57.800 407.400 ;
        RECT 55.000 406.200 55.600 406.800 ;
        RECT 60.400 406.200 61.200 407.000 ;
        RECT 50.200 402.200 51.400 406.200 ;
        RECT 54.800 402.200 55.600 406.200 ;
        RECT 59.200 405.600 61.200 406.200 ;
        RECT 59.200 402.200 60.000 405.600 ;
        RECT 63.600 402.200 64.400 410.600 ;
        RECT 65.200 410.800 69.400 411.400 ;
        RECT 65.200 402.200 66.000 410.800 ;
        RECT 71.800 410.400 72.400 413.600 ;
        RECT 79.000 413.400 79.800 413.600 ;
        RECT 78.000 412.400 78.800 412.600 ;
        RECT 80.600 412.400 81.400 412.600 ;
        RECT 76.400 411.800 81.400 412.400 ;
        RECT 76.400 411.600 77.200 411.800 ;
        RECT 84.400 411.600 85.200 414.400 ;
        RECT 87.800 413.800 88.600 414.400 ;
        RECT 91.000 413.800 91.800 414.400 ;
        RECT 94.600 413.800 95.400 414.400 ;
        RECT 86.000 413.000 88.600 413.800 ;
        RECT 89.400 413.000 91.800 413.800 ;
        RECT 92.800 413.000 95.400 413.800 ;
        RECT 98.800 413.600 99.600 415.200 ;
        RECT 87.800 411.600 88.600 413.000 ;
        RECT 91.000 411.600 91.800 413.000 ;
        RECT 94.600 411.600 95.400 413.000 ;
        RECT 78.000 411.000 83.600 411.200 ;
        RECT 77.800 410.800 83.600 411.000 ;
        RECT 84.400 410.800 86.800 411.600 ;
        RECT 87.800 410.800 90.000 411.600 ;
        RECT 91.000 410.800 93.200 411.600 ;
        RECT 94.600 410.800 96.400 411.600 ;
        RECT 70.000 409.800 72.400 410.400 ;
        RECT 73.800 410.600 83.600 410.800 ;
        RECT 73.800 410.200 78.600 410.600 ;
        RECT 70.000 408.800 70.600 409.800 ;
        RECT 69.200 408.000 70.600 408.800 ;
        RECT 72.200 409.000 73.000 409.200 ;
        RECT 73.800 409.000 74.400 410.200 ;
        RECT 72.200 408.400 74.400 409.000 ;
        RECT 75.000 409.000 80.400 409.600 ;
        RECT 75.000 408.800 75.800 409.000 ;
        RECT 79.600 408.800 80.400 409.000 ;
        RECT 73.400 407.400 74.200 407.600 ;
        RECT 76.200 407.400 77.000 407.600 ;
        RECT 70.000 406.200 70.800 407.000 ;
        RECT 73.400 406.800 77.000 407.400 ;
        RECT 74.200 406.200 74.800 406.800 ;
        RECT 79.600 406.200 80.400 407.000 ;
        RECT 69.400 402.200 70.600 406.200 ;
        RECT 74.000 402.200 74.800 406.200 ;
        RECT 78.400 405.600 80.400 406.200 ;
        RECT 78.400 402.200 79.200 405.600 ;
        RECT 82.800 402.200 83.600 410.600 ;
        RECT 86.000 402.200 86.800 410.800 ;
        RECT 89.200 402.200 90.000 410.800 ;
        RECT 92.400 402.200 93.200 410.800 ;
        RECT 95.600 402.200 96.400 410.800 ;
        RECT 100.400 402.200 101.200 415.800 ;
        RECT 103.600 415.400 104.400 419.800 ;
        RECT 107.800 418.400 109.000 419.800 ;
        RECT 107.800 417.800 109.200 418.400 ;
        RECT 112.400 417.800 113.200 419.800 ;
        RECT 116.800 418.400 117.600 419.800 ;
        RECT 116.800 417.800 118.800 418.400 ;
        RECT 108.400 417.000 109.200 417.800 ;
        RECT 112.600 417.200 113.200 417.800 ;
        RECT 112.600 416.600 115.400 417.200 ;
        RECT 114.600 416.400 115.400 416.600 ;
        RECT 116.400 416.400 117.200 417.200 ;
        RECT 118.000 417.000 118.800 417.800 ;
        RECT 106.600 415.400 107.400 415.600 ;
        RECT 103.600 414.800 107.400 415.400 ;
        RECT 103.600 411.400 104.400 414.800 ;
        RECT 110.600 414.200 111.400 414.400 ;
        RECT 116.400 414.200 117.000 416.400 ;
        RECT 121.200 415.000 122.000 419.800 ;
        RECT 122.800 415.800 123.600 419.800 ;
        RECT 127.200 416.200 128.800 419.800 ;
        RECT 122.800 415.200 125.000 415.800 ;
        RECT 126.000 415.400 127.600 415.600 ;
        RECT 124.200 415.000 125.000 415.200 ;
        RECT 125.600 414.800 127.600 415.400 ;
        RECT 125.600 414.400 126.200 414.800 ;
        RECT 119.600 414.200 121.200 414.400 ;
        RECT 110.200 413.600 121.200 414.200 ;
        RECT 122.800 413.800 126.200 414.400 ;
        RECT 122.800 413.600 124.400 413.800 ;
        RECT 108.400 412.800 109.200 413.000 ;
        RECT 105.400 412.200 109.200 412.800 ;
        RECT 110.200 412.400 110.800 413.600 ;
        RECT 117.400 413.400 118.200 413.600 ;
        RECT 126.800 413.400 127.600 414.200 ;
        RECT 126.800 412.800 127.400 413.400 ;
        RECT 116.400 412.400 117.200 412.600 ;
        RECT 119.000 412.400 119.800 412.600 ;
        RECT 105.400 412.000 106.200 412.200 ;
        RECT 110.000 411.600 110.800 412.400 ;
        RECT 114.800 411.800 119.800 412.400 ;
        RECT 124.800 412.200 127.400 412.800 ;
        RECT 128.200 412.800 128.800 416.200 ;
        RECT 132.400 415.800 133.200 419.800 ;
        RECT 138.800 415.800 139.600 419.800 ;
        RECT 140.400 416.000 141.200 419.800 ;
        RECT 143.600 416.000 144.400 419.800 ;
        RECT 145.800 416.400 146.600 419.800 ;
        RECT 140.400 415.800 144.400 416.000 ;
        RECT 129.400 414.800 130.200 415.600 ;
        RECT 130.800 415.200 133.200 415.800 ;
        RECT 130.800 415.000 131.600 415.200 ;
        RECT 129.600 414.400 130.200 414.800 ;
        RECT 139.000 414.400 139.600 415.800 ;
        RECT 140.600 415.400 144.200 415.800 ;
        RECT 145.200 415.600 147.600 416.400 ;
        RECT 142.800 414.400 143.600 414.800 ;
        RECT 129.600 413.600 130.400 414.400 ;
        RECT 131.600 413.600 133.200 414.400 ;
        RECT 134.000 414.300 134.800 414.400 ;
        RECT 138.800 414.300 141.400 414.400 ;
        RECT 134.000 413.700 141.400 414.300 ;
        RECT 142.800 413.800 144.400 414.400 ;
        RECT 134.000 413.600 134.800 413.700 ;
        RECT 138.800 413.600 141.400 413.700 ;
        RECT 143.600 413.600 144.400 413.800 ;
        RECT 128.200 412.400 129.200 412.800 ;
        RECT 128.200 412.200 130.000 412.400 ;
        RECT 124.800 412.000 125.600 412.200 ;
        RECT 114.800 411.600 115.600 411.800 ;
        RECT 128.600 411.600 130.000 412.200 ;
        RECT 107.000 411.400 107.800 411.600 ;
        RECT 103.600 410.800 107.800 411.400 ;
        RECT 102.000 410.300 102.800 410.400 ;
        RECT 103.600 410.300 104.400 410.800 ;
        RECT 110.200 410.400 110.800 411.600 ;
        RECT 127.000 411.400 127.800 411.600 ;
        RECT 116.400 411.000 122.000 411.200 ;
        RECT 116.200 410.800 122.000 411.000 ;
        RECT 102.000 409.700 104.400 410.300 ;
        RECT 102.000 408.800 102.800 409.700 ;
        RECT 103.600 402.200 104.400 409.700 ;
        RECT 108.400 409.800 110.800 410.400 ;
        RECT 112.200 410.600 122.000 410.800 ;
        RECT 112.200 410.200 117.000 410.600 ;
        RECT 108.400 408.800 109.000 409.800 ;
        RECT 107.600 408.000 109.000 408.800 ;
        RECT 110.600 409.000 111.400 409.200 ;
        RECT 112.200 409.000 112.800 410.200 ;
        RECT 110.600 408.400 112.800 409.000 ;
        RECT 113.400 409.000 118.800 409.600 ;
        RECT 113.400 408.800 114.200 409.000 ;
        RECT 118.000 408.800 118.800 409.000 ;
        RECT 111.800 407.400 112.600 407.600 ;
        RECT 114.600 407.400 115.400 407.600 ;
        RECT 108.400 406.200 109.200 407.000 ;
        RECT 111.800 406.800 115.400 407.400 ;
        RECT 112.600 406.200 113.200 406.800 ;
        RECT 118.000 406.200 118.800 407.000 ;
        RECT 107.800 402.200 109.000 406.200 ;
        RECT 112.400 402.200 113.200 406.200 ;
        RECT 116.800 405.600 118.800 406.200 ;
        RECT 116.800 402.200 117.600 405.600 ;
        RECT 121.200 402.200 122.000 410.600 ;
        RECT 124.400 410.800 127.800 411.400 ;
        RECT 124.400 410.200 125.000 410.800 ;
        RECT 128.600 410.200 129.200 411.600 ;
        RECT 138.800 410.200 139.600 410.400 ;
        RECT 140.800 410.200 141.400 413.600 ;
        RECT 142.000 411.600 142.800 413.200 ;
        RECT 122.800 409.600 125.000 410.200 ;
        RECT 122.800 402.200 123.600 409.600 ;
        RECT 124.200 409.400 125.000 409.600 ;
        RECT 127.200 409.600 129.200 410.200 ;
        RECT 130.800 409.600 133.200 410.200 ;
        RECT 138.800 409.600 140.200 410.200 ;
        RECT 140.800 409.600 141.800 410.200 ;
        RECT 127.200 408.400 128.800 409.600 ;
        RECT 130.800 409.400 131.600 409.600 ;
        RECT 126.000 407.600 128.800 408.400 ;
        RECT 127.200 402.200 128.800 407.600 ;
        RECT 132.400 402.200 133.200 409.600 ;
        RECT 139.600 408.400 140.200 409.600 ;
        RECT 139.600 407.600 140.400 408.400 ;
        RECT 141.000 402.200 141.800 409.600 ;
        RECT 145.200 408.800 146.000 410.400 ;
        RECT 146.800 402.200 147.600 415.600 ;
        RECT 150.000 415.800 150.800 419.800 ;
        RECT 154.400 416.200 156.000 419.800 ;
        RECT 150.000 415.200 152.200 415.800 ;
        RECT 153.200 415.400 154.800 415.600 ;
        RECT 148.400 413.600 149.200 415.200 ;
        RECT 151.400 415.000 152.200 415.200 ;
        RECT 152.800 414.800 154.800 415.400 ;
        RECT 152.800 414.400 153.400 414.800 ;
        RECT 150.000 413.800 153.400 414.400 ;
        RECT 150.000 413.600 151.600 413.800 ;
        RECT 154.000 413.400 154.800 414.200 ;
        RECT 154.000 412.800 154.600 413.400 ;
        RECT 152.000 412.200 154.600 412.800 ;
        RECT 155.400 412.800 156.000 416.200 ;
        RECT 159.600 415.800 160.400 419.800 ;
        RECT 163.800 416.400 164.600 419.800 ;
        RECT 156.600 414.800 157.400 415.600 ;
        RECT 158.000 415.200 160.400 415.800 ;
        RECT 162.800 415.800 164.600 416.400 ;
        RECT 166.600 416.400 167.400 419.800 ;
        RECT 166.600 415.800 168.400 416.400 ;
        RECT 170.800 416.000 171.600 419.800 ;
        RECT 174.000 416.000 174.800 419.800 ;
        RECT 170.800 415.800 174.800 416.000 ;
        RECT 175.600 415.800 176.400 419.800 ;
        RECT 177.200 415.800 178.000 419.800 ;
        RECT 178.800 416.000 179.600 419.800 ;
        RECT 182.000 416.000 182.800 419.800 ;
        RECT 185.200 417.800 186.000 419.800 ;
        RECT 178.800 415.800 182.800 416.000 ;
        RECT 158.000 415.000 158.800 415.200 ;
        RECT 156.800 414.400 157.400 414.800 ;
        RECT 156.800 413.600 157.600 414.400 ;
        RECT 158.800 413.600 160.400 414.400 ;
        RECT 161.200 413.600 162.000 415.200 ;
        RECT 155.400 412.400 156.400 412.800 ;
        RECT 155.400 412.200 157.200 412.400 ;
        RECT 152.000 412.000 152.800 412.200 ;
        RECT 155.800 411.600 157.200 412.200 ;
        RECT 154.200 411.400 155.000 411.600 ;
        RECT 151.600 410.800 155.000 411.400 ;
        RECT 151.600 410.200 152.200 410.800 ;
        RECT 155.800 410.200 156.400 411.600 ;
        RECT 150.000 409.600 152.200 410.200 ;
        RECT 150.000 402.200 150.800 409.600 ;
        RECT 151.400 409.400 152.200 409.600 ;
        RECT 154.400 409.600 156.400 410.200 ;
        RECT 158.000 409.600 160.400 410.200 ;
        RECT 154.400 408.400 156.000 409.600 ;
        RECT 158.000 409.400 158.800 409.600 ;
        RECT 153.200 407.600 156.000 408.400 ;
        RECT 154.400 402.200 156.000 407.600 ;
        RECT 159.600 402.200 160.400 409.600 ;
        RECT 162.800 402.200 163.600 415.800 ;
        RECT 164.400 408.800 165.200 410.400 ;
        RECT 166.000 408.800 166.800 410.400 ;
        RECT 167.600 402.200 168.400 415.800 ;
        RECT 171.000 415.400 174.600 415.800 ;
        RECT 169.200 413.600 170.000 415.200 ;
        RECT 171.600 414.400 172.400 414.800 ;
        RECT 175.600 414.400 176.200 415.800 ;
        RECT 177.400 414.400 178.000 415.800 ;
        RECT 179.000 415.400 182.600 415.800 ;
        RECT 183.600 415.600 184.400 417.200 ;
        RECT 185.400 416.300 186.000 417.800 ;
        RECT 188.600 416.400 189.400 417.200 ;
        RECT 188.400 416.300 189.200 416.400 ;
        RECT 185.300 415.700 189.200 416.300 ;
        RECT 190.000 415.800 190.800 419.800 ;
        RECT 181.200 414.400 182.000 414.800 ;
        RECT 170.800 413.800 172.400 414.400 ;
        RECT 170.800 413.600 171.600 413.800 ;
        RECT 173.800 413.600 176.400 414.400 ;
        RECT 177.200 413.600 179.800 414.400 ;
        RECT 181.200 414.300 182.800 414.400 ;
        RECT 183.700 414.300 184.300 415.600 ;
        RECT 185.400 414.400 186.000 415.700 ;
        RECT 188.400 415.600 189.200 415.700 ;
        RECT 181.200 413.800 184.300 414.300 ;
        RECT 182.000 413.700 184.300 413.800 ;
        RECT 182.000 413.600 182.800 413.700 ;
        RECT 185.200 413.600 186.000 414.400 ;
        RECT 169.300 412.300 169.900 413.600 ;
        RECT 172.400 412.300 173.200 413.200 ;
        RECT 169.300 411.700 173.200 412.300 ;
        RECT 172.400 411.600 173.200 411.700 ;
        RECT 173.800 410.200 174.400 413.600 ;
        RECT 179.200 412.400 179.800 413.600 ;
        RECT 178.800 411.600 179.800 412.400 ;
        RECT 180.400 411.600 181.200 413.200 ;
        RECT 175.600 410.200 176.400 410.400 ;
        RECT 173.400 409.600 174.400 410.200 ;
        RECT 175.000 409.600 176.400 410.200 ;
        RECT 177.200 410.200 178.000 410.400 ;
        RECT 179.200 410.200 179.800 411.600 ;
        RECT 185.400 410.200 186.000 413.600 ;
        RECT 186.800 410.800 187.600 412.400 ;
        RECT 188.400 412.200 189.200 412.400 ;
        RECT 190.200 412.200 190.800 415.800 ;
        RECT 196.400 417.800 197.200 419.800 ;
        RECT 201.200 417.800 202.000 419.800 ;
        RECT 196.400 414.400 197.000 417.800 ;
        RECT 198.000 415.600 198.800 417.200 ;
        RECT 201.200 414.400 201.800 417.800 ;
        RECT 202.800 415.600 203.600 417.200 ;
        RECT 191.600 412.800 192.400 414.400 ;
        RECT 193.200 414.300 194.000 414.400 ;
        RECT 196.400 414.300 197.200 414.400 ;
        RECT 193.200 413.700 197.200 414.300 ;
        RECT 193.200 413.600 194.000 413.700 ;
        RECT 196.400 413.600 197.200 413.700 ;
        RECT 201.200 413.600 202.000 414.400 ;
        RECT 193.200 412.200 194.000 412.400 ;
        RECT 188.400 411.600 190.800 412.200 ;
        RECT 192.400 411.600 194.000 412.200 ;
        RECT 188.600 410.200 189.200 411.600 ;
        RECT 192.400 411.200 193.200 411.600 ;
        RECT 194.800 410.800 195.600 412.400 ;
        RECT 196.400 410.200 197.000 413.600 ;
        RECT 201.200 412.400 201.800 413.600 ;
        RECT 204.400 412.400 205.200 419.800 ;
        RECT 207.600 415.200 208.400 419.800 ;
        RECT 206.200 414.600 208.400 415.200 ;
        RECT 199.600 410.800 200.400 412.400 ;
        RECT 201.200 411.600 202.000 412.400 ;
        RECT 201.200 410.200 201.800 411.600 ;
        RECT 204.400 410.200 205.000 412.400 ;
        RECT 206.200 411.600 206.800 414.600 ;
        RECT 207.600 411.600 208.400 413.200 ;
        RECT 205.600 410.800 206.800 411.600 ;
        RECT 206.200 410.200 206.800 410.800 ;
        RECT 177.200 409.600 178.600 410.200 ;
        RECT 179.200 409.600 180.200 410.200 ;
        RECT 173.400 402.200 174.200 409.600 ;
        RECT 175.000 408.400 175.600 409.600 ;
        RECT 174.800 407.600 175.600 408.400 ;
        RECT 178.000 408.400 178.600 409.600 ;
        RECT 178.000 407.600 178.800 408.400 ;
        RECT 179.400 402.200 180.200 409.600 ;
        RECT 185.200 409.400 187.000 410.200 ;
        RECT 186.200 402.200 187.000 409.400 ;
        RECT 188.400 402.200 189.200 410.200 ;
        RECT 190.000 409.600 194.000 410.200 ;
        RECT 190.000 402.200 190.800 409.600 ;
        RECT 193.200 402.200 194.000 409.600 ;
        RECT 195.400 409.400 197.200 410.200 ;
        RECT 200.200 409.400 202.000 410.200 ;
        RECT 195.400 402.200 196.200 409.400 ;
        RECT 200.200 402.200 201.000 409.400 ;
        RECT 204.400 402.200 205.200 410.200 ;
        RECT 206.200 409.600 208.400 410.200 ;
        RECT 207.600 402.200 208.400 409.600 ;
        RECT 209.200 402.200 210.000 419.800 ;
        RECT 214.000 417.800 214.800 419.800 ;
        RECT 210.800 416.300 211.600 417.200 ;
        RECT 212.400 416.300 213.200 417.200 ;
        RECT 210.800 415.700 213.200 416.300 ;
        RECT 210.800 415.600 211.600 415.700 ;
        RECT 212.400 415.600 213.200 415.700 ;
        RECT 214.200 414.400 214.800 417.800 ;
        RECT 212.400 414.300 213.200 414.400 ;
        RECT 214.000 414.300 214.800 414.400 ;
        RECT 212.400 413.700 214.800 414.300 ;
        RECT 212.400 413.600 213.200 413.700 ;
        RECT 214.000 413.600 214.800 413.700 ;
        RECT 217.200 413.600 218.000 415.200 ;
        RECT 214.200 410.200 214.800 413.600 ;
        RECT 215.600 412.300 216.400 412.400 ;
        RECT 217.300 412.300 217.900 413.600 ;
        RECT 215.600 411.700 217.900 412.300 ;
        RECT 215.600 410.800 216.400 411.700 ;
        RECT 214.000 409.400 215.800 410.200 ;
        RECT 215.000 402.200 215.800 409.400 ;
        RECT 218.800 402.200 219.600 419.800 ;
        RECT 220.400 415.400 221.200 419.800 ;
        RECT 224.600 418.400 225.800 419.800 ;
        RECT 224.600 417.800 226.000 418.400 ;
        RECT 229.200 417.800 230.000 419.800 ;
        RECT 233.600 418.400 234.400 419.800 ;
        RECT 233.600 417.800 235.600 418.400 ;
        RECT 225.200 417.000 226.000 417.800 ;
        RECT 229.400 417.200 230.000 417.800 ;
        RECT 229.400 416.600 232.200 417.200 ;
        RECT 231.400 416.400 232.200 416.600 ;
        RECT 233.200 416.400 234.000 417.200 ;
        RECT 234.800 417.000 235.600 417.800 ;
        RECT 223.400 415.400 224.200 415.600 ;
        RECT 220.400 414.800 224.200 415.400 ;
        RECT 220.400 411.400 221.200 414.800 ;
        RECT 227.400 414.200 228.200 414.400 ;
        RECT 233.200 414.200 233.800 416.400 ;
        RECT 238.000 415.000 238.800 419.800 ;
        RECT 236.400 414.200 238.000 414.400 ;
        RECT 227.000 413.600 238.000 414.200 ;
        RECT 225.200 412.800 226.000 413.000 ;
        RECT 222.200 412.200 226.000 412.800 ;
        RECT 227.000 412.300 227.600 413.600 ;
        RECT 234.200 413.400 235.000 413.600 ;
        RECT 233.200 412.400 234.000 412.600 ;
        RECT 235.800 412.400 236.600 412.600 ;
        RECT 228.400 412.300 229.200 412.400 ;
        RECT 222.200 412.000 223.000 412.200 ;
        RECT 226.900 411.700 229.200 412.300 ;
        RECT 223.800 411.400 224.600 411.600 ;
        RECT 220.400 410.800 224.600 411.400 ;
        RECT 220.400 402.200 221.200 410.800 ;
        RECT 227.000 410.400 227.600 411.700 ;
        RECT 228.400 411.600 229.200 411.700 ;
        RECT 231.600 411.800 236.600 412.400 ;
        RECT 231.600 411.600 232.400 411.800 ;
        RECT 233.200 411.000 238.800 411.200 ;
        RECT 233.000 410.800 238.800 411.000 ;
        RECT 225.200 409.800 227.600 410.400 ;
        RECT 229.000 410.600 238.800 410.800 ;
        RECT 229.000 410.200 233.800 410.600 ;
        RECT 225.200 408.800 225.800 409.800 ;
        RECT 224.400 408.000 225.800 408.800 ;
        RECT 227.400 409.000 228.200 409.200 ;
        RECT 229.000 409.000 229.600 410.200 ;
        RECT 227.400 408.400 229.600 409.000 ;
        RECT 230.200 409.000 235.600 409.600 ;
        RECT 230.200 408.800 231.000 409.000 ;
        RECT 234.800 408.800 235.600 409.000 ;
        RECT 228.600 407.400 229.400 407.600 ;
        RECT 231.400 407.400 232.200 407.600 ;
        RECT 225.200 406.200 226.000 407.000 ;
        RECT 228.600 406.800 232.200 407.400 ;
        RECT 229.400 406.200 230.000 406.800 ;
        RECT 234.800 406.200 235.600 407.000 ;
        RECT 224.600 402.200 225.800 406.200 ;
        RECT 229.200 402.200 230.000 406.200 ;
        RECT 233.600 405.600 235.600 406.200 ;
        RECT 233.600 402.200 234.400 405.600 ;
        RECT 238.000 402.200 238.800 410.600 ;
        RECT 239.600 402.200 240.400 419.800 ;
        RECT 241.200 415.600 242.000 417.200 ;
        RECT 242.800 415.400 243.600 419.800 ;
        RECT 247.000 418.400 248.200 419.800 ;
        RECT 247.000 417.800 248.400 418.400 ;
        RECT 251.600 417.800 252.400 419.800 ;
        RECT 256.000 418.400 256.800 419.800 ;
        RECT 256.000 417.800 258.000 418.400 ;
        RECT 247.600 417.000 248.400 417.800 ;
        RECT 251.800 417.200 252.400 417.800 ;
        RECT 251.800 416.600 254.600 417.200 ;
        RECT 253.800 416.400 254.600 416.600 ;
        RECT 255.600 416.400 256.400 417.200 ;
        RECT 257.200 417.000 258.000 417.800 ;
        RECT 245.800 415.400 246.600 415.600 ;
        RECT 242.800 414.800 246.600 415.400 ;
        RECT 242.800 411.400 243.600 414.800 ;
        RECT 249.800 414.200 250.600 414.400 ;
        RECT 255.600 414.200 256.200 416.400 ;
        RECT 260.400 415.000 261.200 419.800 ;
        RECT 258.800 414.200 260.400 414.400 ;
        RECT 249.400 413.600 260.400 414.200 ;
        RECT 247.600 412.800 248.400 413.000 ;
        RECT 244.600 412.200 248.400 412.800 ;
        RECT 249.400 412.400 250.000 413.600 ;
        RECT 256.600 413.400 257.400 413.600 ;
        RECT 255.600 412.400 256.400 412.600 ;
        RECT 258.200 412.400 259.000 412.600 ;
        RECT 244.600 412.000 245.400 412.200 ;
        RECT 249.200 411.600 250.000 412.400 ;
        RECT 254.000 411.800 259.000 412.400 ;
        RECT 262.000 412.400 262.800 419.800 ;
        RECT 265.200 415.200 266.000 419.800 ;
        RECT 269.400 416.400 270.200 419.800 ;
        RECT 268.400 415.800 270.200 416.400 ;
        RECT 271.600 416.000 272.400 419.800 ;
        RECT 274.800 416.000 275.600 419.800 ;
        RECT 271.600 415.800 275.600 416.000 ;
        RECT 276.400 415.800 277.200 419.800 ;
        RECT 263.800 414.600 266.000 415.200 ;
        RECT 254.000 411.600 254.800 411.800 ;
        RECT 246.200 411.400 247.000 411.600 ;
        RECT 242.800 410.800 247.000 411.400 ;
        RECT 242.800 402.200 243.600 410.800 ;
        RECT 249.400 410.400 250.000 411.600 ;
        RECT 255.600 411.000 261.200 411.200 ;
        RECT 255.400 410.800 261.200 411.000 ;
        RECT 247.600 409.800 250.000 410.400 ;
        RECT 251.400 410.600 261.200 410.800 ;
        RECT 251.400 410.200 256.200 410.600 ;
        RECT 247.600 408.800 248.200 409.800 ;
        RECT 246.800 408.000 248.200 408.800 ;
        RECT 249.800 409.000 250.600 409.200 ;
        RECT 251.400 409.000 252.000 410.200 ;
        RECT 249.800 408.400 252.000 409.000 ;
        RECT 252.600 409.000 258.000 409.600 ;
        RECT 252.600 408.800 253.400 409.000 ;
        RECT 257.200 408.800 258.000 409.000 ;
        RECT 251.000 407.400 251.800 407.600 ;
        RECT 253.800 407.400 254.600 407.600 ;
        RECT 247.600 406.200 248.400 407.000 ;
        RECT 251.000 406.800 254.600 407.400 ;
        RECT 251.800 406.200 252.400 406.800 ;
        RECT 257.200 406.200 258.000 407.000 ;
        RECT 247.000 402.200 248.200 406.200 ;
        RECT 251.600 402.200 252.400 406.200 ;
        RECT 256.000 405.600 258.000 406.200 ;
        RECT 256.000 402.200 256.800 405.600 ;
        RECT 260.400 402.200 261.200 410.600 ;
        RECT 262.000 410.200 262.600 412.400 ;
        RECT 263.800 411.600 264.400 414.600 ;
        RECT 266.800 413.600 267.600 415.200 ;
        RECT 268.400 414.300 269.200 415.800 ;
        RECT 271.800 415.400 275.400 415.800 ;
        RECT 272.400 414.400 273.200 414.800 ;
        RECT 276.400 414.400 277.000 415.800 ;
        RECT 278.000 415.400 278.800 419.800 ;
        RECT 282.200 418.400 283.400 419.800 ;
        RECT 282.200 417.800 283.600 418.400 ;
        RECT 286.800 417.800 287.600 419.800 ;
        RECT 291.200 418.400 292.000 419.800 ;
        RECT 291.200 417.800 293.200 418.400 ;
        RECT 282.800 417.000 283.600 417.800 ;
        RECT 287.000 417.200 287.600 417.800 ;
        RECT 287.000 416.600 289.800 417.200 ;
        RECT 289.000 416.400 289.800 416.600 ;
        RECT 290.800 416.400 291.600 417.200 ;
        RECT 292.400 417.000 293.200 417.800 ;
        RECT 281.000 415.400 281.800 415.600 ;
        RECT 278.000 414.800 281.800 415.400 ;
        RECT 270.000 414.300 270.800 414.400 ;
        RECT 268.400 413.700 270.800 414.300 ;
        RECT 265.200 411.600 266.000 413.200 ;
        RECT 263.200 410.800 264.400 411.600 ;
        RECT 263.800 410.200 264.400 410.800 ;
        RECT 262.000 402.200 262.800 410.200 ;
        RECT 263.800 409.600 266.000 410.200 ;
        RECT 265.200 402.200 266.000 409.600 ;
        RECT 268.400 402.200 269.200 413.700 ;
        RECT 270.000 413.600 270.800 413.700 ;
        RECT 271.600 413.800 273.200 414.400 ;
        RECT 271.600 413.600 272.400 413.800 ;
        RECT 274.600 413.600 277.200 414.400 ;
        RECT 273.200 412.300 274.000 413.200 ;
        RECT 270.100 411.700 274.000 412.300 ;
        RECT 270.100 410.400 270.700 411.700 ;
        RECT 273.200 411.600 274.000 411.700 ;
        RECT 274.600 412.400 275.200 413.600 ;
        RECT 274.600 411.600 275.600 412.400 ;
        RECT 270.000 408.800 270.800 410.400 ;
        RECT 274.600 410.200 275.200 411.600 ;
        RECT 278.000 411.400 278.800 414.800 ;
        RECT 285.000 414.200 285.800 414.400 ;
        RECT 290.800 414.200 291.400 416.400 ;
        RECT 295.600 415.000 296.400 419.800 ;
        RECT 303.600 415.200 304.400 419.800 ;
        RECT 306.800 415.200 307.600 419.800 ;
        RECT 310.000 415.200 310.800 419.800 ;
        RECT 313.200 415.200 314.000 419.800 ;
        RECT 302.000 414.400 304.400 415.200 ;
        RECT 305.400 414.400 307.600 415.200 ;
        RECT 308.600 414.400 310.800 415.200 ;
        RECT 312.200 414.400 314.000 415.200 ;
        RECT 316.400 415.400 317.200 419.800 ;
        RECT 320.600 418.400 321.800 419.800 ;
        RECT 320.600 417.800 322.000 418.400 ;
        RECT 325.200 417.800 326.000 419.800 ;
        RECT 329.600 418.400 330.400 419.800 ;
        RECT 329.600 417.800 331.600 418.400 ;
        RECT 321.200 417.000 322.000 417.800 ;
        RECT 325.400 417.200 326.000 417.800 ;
        RECT 325.400 416.600 328.200 417.200 ;
        RECT 327.400 416.400 328.200 416.600 ;
        RECT 329.200 416.400 330.000 417.200 ;
        RECT 330.800 417.000 331.600 417.800 ;
        RECT 319.400 415.400 320.200 415.600 ;
        RECT 316.400 414.800 320.200 415.400 ;
        RECT 294.000 414.200 295.600 414.400 ;
        RECT 284.600 413.600 295.600 414.200 ;
        RECT 282.800 412.800 283.600 413.000 ;
        RECT 279.800 412.200 283.600 412.800 ;
        RECT 279.800 412.000 280.600 412.200 ;
        RECT 281.400 411.400 282.200 411.600 ;
        RECT 278.000 410.800 282.200 411.400 ;
        RECT 276.400 410.200 277.200 410.400 ;
        RECT 274.200 409.600 275.200 410.200 ;
        RECT 275.800 409.600 277.200 410.200 ;
        RECT 274.200 402.200 275.000 409.600 ;
        RECT 275.800 408.400 276.400 409.600 ;
        RECT 275.600 407.600 276.400 408.400 ;
        RECT 278.000 402.200 278.800 410.800 ;
        RECT 284.600 410.400 285.200 413.600 ;
        RECT 291.800 413.400 292.600 413.600 ;
        RECT 302.000 411.600 302.800 414.400 ;
        RECT 305.400 413.800 306.200 414.400 ;
        RECT 308.600 413.800 309.400 414.400 ;
        RECT 312.200 413.800 313.000 414.400 ;
        RECT 303.600 413.000 306.200 413.800 ;
        RECT 307.000 413.000 309.400 413.800 ;
        RECT 310.400 413.000 313.000 413.800 ;
        RECT 305.400 411.600 306.200 413.000 ;
        RECT 308.600 411.600 309.400 413.000 ;
        RECT 312.200 411.600 313.000 413.000 ;
        RECT 290.800 411.000 296.400 411.200 ;
        RECT 290.600 410.800 296.400 411.000 ;
        RECT 302.000 410.800 304.400 411.600 ;
        RECT 305.400 410.800 307.600 411.600 ;
        RECT 308.600 410.800 310.800 411.600 ;
        RECT 312.200 410.800 314.000 411.600 ;
        RECT 282.800 409.800 285.200 410.400 ;
        RECT 286.600 410.600 296.400 410.800 ;
        RECT 286.600 410.200 291.400 410.600 ;
        RECT 282.800 408.800 283.400 409.800 ;
        RECT 282.000 408.000 283.400 408.800 ;
        RECT 285.000 409.000 285.800 409.200 ;
        RECT 286.600 409.000 287.200 410.200 ;
        RECT 285.000 408.400 287.200 409.000 ;
        RECT 287.800 409.000 293.200 409.600 ;
        RECT 287.800 408.800 288.600 409.000 ;
        RECT 292.400 408.800 293.200 409.000 ;
        RECT 286.200 407.400 287.000 407.600 ;
        RECT 289.000 407.400 289.800 407.600 ;
        RECT 282.800 406.200 283.600 407.000 ;
        RECT 286.200 406.800 289.800 407.400 ;
        RECT 287.000 406.200 287.600 406.800 ;
        RECT 292.400 406.200 293.200 407.000 ;
        RECT 282.200 402.200 283.400 406.200 ;
        RECT 286.800 402.200 287.600 406.200 ;
        RECT 291.200 405.600 293.200 406.200 ;
        RECT 291.200 402.200 292.000 405.600 ;
        RECT 295.600 402.200 296.400 410.600 ;
        RECT 303.600 402.200 304.400 410.800 ;
        RECT 306.800 402.200 307.600 410.800 ;
        RECT 310.000 402.200 310.800 410.800 ;
        RECT 313.200 402.200 314.000 410.800 ;
        RECT 316.400 411.400 317.200 414.800 ;
        RECT 323.400 414.200 324.200 414.400 ;
        RECT 329.200 414.200 329.800 416.400 ;
        RECT 334.000 415.000 334.800 419.800 ;
        RECT 332.400 414.200 334.000 414.400 ;
        RECT 323.000 413.600 334.000 414.200 ;
        RECT 321.200 412.800 322.000 413.000 ;
        RECT 318.200 412.200 322.000 412.800 ;
        RECT 323.000 412.400 323.600 413.600 ;
        RECT 330.200 413.400 331.000 413.600 ;
        RECT 329.200 412.400 330.000 412.600 ;
        RECT 331.800 412.400 332.600 412.600 ;
        RECT 318.200 412.000 319.000 412.200 ;
        RECT 322.800 411.600 323.600 412.400 ;
        RECT 327.600 411.800 332.600 412.400 ;
        RECT 335.600 412.400 336.400 419.800 ;
        RECT 338.800 415.200 339.600 419.800 ;
        RECT 337.400 414.600 339.600 415.200 ;
        RECT 327.600 411.600 328.400 411.800 ;
        RECT 319.800 411.400 320.600 411.600 ;
        RECT 316.400 410.800 320.600 411.400 ;
        RECT 316.400 402.200 317.200 410.800 ;
        RECT 323.000 410.400 323.600 411.600 ;
        RECT 329.200 411.000 334.800 411.200 ;
        RECT 329.000 410.800 334.800 411.000 ;
        RECT 321.200 409.800 323.600 410.400 ;
        RECT 325.000 410.600 334.800 410.800 ;
        RECT 325.000 410.200 329.800 410.600 ;
        RECT 321.200 408.800 321.800 409.800 ;
        RECT 320.400 408.000 321.800 408.800 ;
        RECT 323.400 409.000 324.200 409.200 ;
        RECT 325.000 409.000 325.600 410.200 ;
        RECT 323.400 408.400 325.600 409.000 ;
        RECT 326.200 409.000 331.600 409.600 ;
        RECT 326.200 408.800 327.000 409.000 ;
        RECT 330.800 408.800 331.600 409.000 ;
        RECT 324.600 407.400 325.400 407.600 ;
        RECT 327.400 407.400 328.200 407.600 ;
        RECT 321.200 406.200 322.000 407.000 ;
        RECT 324.600 406.800 328.200 407.400 ;
        RECT 325.400 406.200 326.000 406.800 ;
        RECT 330.800 406.200 331.600 407.000 ;
        RECT 320.600 402.200 321.800 406.200 ;
        RECT 325.200 402.200 326.000 406.200 ;
        RECT 329.600 405.600 331.600 406.200 ;
        RECT 329.600 402.200 330.400 405.600 ;
        RECT 334.000 402.200 334.800 410.600 ;
        RECT 335.600 410.200 336.200 412.400 ;
        RECT 337.400 411.600 338.000 414.600 ;
        RECT 338.800 411.600 339.600 413.200 ;
        RECT 340.400 412.400 341.200 419.800 ;
        RECT 343.600 415.200 344.400 419.800 ;
        RECT 342.200 414.600 344.400 415.200 ;
        RECT 345.200 415.200 346.000 419.800 ;
        RECT 345.200 414.600 347.400 415.200 ;
        RECT 336.800 410.800 338.000 411.600 ;
        RECT 337.400 410.200 338.000 410.800 ;
        RECT 340.400 410.200 341.000 412.400 ;
        RECT 342.200 411.600 342.800 414.600 ;
        RECT 343.600 412.300 344.400 413.200 ;
        RECT 345.200 412.300 346.000 413.200 ;
        RECT 343.600 411.700 346.000 412.300 ;
        RECT 343.600 411.600 344.400 411.700 ;
        RECT 345.200 411.600 346.000 411.700 ;
        RECT 346.800 411.600 347.400 414.600 ;
        RECT 348.400 412.400 349.200 419.800 ;
        RECT 341.600 410.800 342.800 411.600 ;
        RECT 342.200 410.200 342.800 410.800 ;
        RECT 346.800 410.800 348.000 411.600 ;
        RECT 346.800 410.200 347.400 410.800 ;
        RECT 348.600 410.200 349.200 412.400 ;
        RECT 335.600 402.200 336.400 410.200 ;
        RECT 337.400 409.600 339.600 410.200 ;
        RECT 338.800 402.200 339.600 409.600 ;
        RECT 340.400 402.200 341.200 410.200 ;
        RECT 342.200 409.600 344.400 410.200 ;
        RECT 343.600 402.200 344.400 409.600 ;
        RECT 345.200 409.600 347.400 410.200 ;
        RECT 345.200 402.200 346.000 409.600 ;
        RECT 348.400 402.200 349.200 410.200 ;
        RECT 350.000 412.400 350.800 419.800 ;
        RECT 353.200 415.200 354.000 419.800 ;
        RECT 356.400 416.000 357.200 419.800 ;
        RECT 351.800 414.600 354.000 415.200 ;
        RECT 356.200 415.200 357.200 416.000 ;
        RECT 350.000 410.200 350.600 412.400 ;
        RECT 351.800 411.600 352.400 414.600 ;
        RECT 353.200 412.300 354.000 413.200 ;
        RECT 354.800 412.300 355.600 412.400 ;
        RECT 353.200 411.700 355.600 412.300 ;
        RECT 353.200 411.600 354.000 411.700 ;
        RECT 354.800 411.600 355.600 411.700 ;
        RECT 351.200 410.800 352.400 411.600 ;
        RECT 351.800 410.200 352.400 410.800 ;
        RECT 356.200 410.800 357.000 415.200 ;
        RECT 358.000 414.600 358.800 419.800 ;
        RECT 364.400 416.600 365.200 419.800 ;
        RECT 366.000 417.000 366.800 419.800 ;
        RECT 367.600 417.000 368.400 419.800 ;
        RECT 369.200 417.000 370.000 419.800 ;
        RECT 370.800 417.000 371.600 419.800 ;
        RECT 374.000 417.000 374.800 419.800 ;
        RECT 377.200 417.000 378.000 419.800 ;
        RECT 378.800 417.000 379.600 419.800 ;
        RECT 380.400 417.000 381.200 419.800 ;
        RECT 362.800 415.800 365.200 416.600 ;
        RECT 382.000 416.600 382.800 419.800 ;
        RECT 362.800 415.200 363.600 415.800 ;
        RECT 357.600 414.000 358.800 414.600 ;
        RECT 361.800 414.600 363.600 415.200 ;
        RECT 367.600 415.600 368.600 416.400 ;
        RECT 371.600 415.600 373.200 416.400 ;
        RECT 374.000 415.800 378.600 416.400 ;
        RECT 382.000 415.800 384.600 416.600 ;
        RECT 374.000 415.600 374.800 415.800 ;
        RECT 357.600 412.000 358.200 414.000 ;
        RECT 361.800 413.400 362.600 414.600 ;
        RECT 358.800 412.600 362.600 413.400 ;
        RECT 367.600 412.800 368.400 415.600 ;
        RECT 374.000 414.800 374.800 415.000 ;
        RECT 370.400 414.200 374.800 414.800 ;
        RECT 370.400 414.000 371.200 414.200 ;
        RECT 377.800 413.400 378.600 415.800 ;
        RECT 383.800 415.200 384.600 415.800 ;
        RECT 383.800 414.400 386.800 415.200 ;
        RECT 388.400 413.800 389.200 419.800 ;
        RECT 390.600 416.400 391.400 419.800 ;
        RECT 390.600 415.800 392.400 416.400 ;
        RECT 370.800 412.600 374.000 413.400 ;
        RECT 377.800 412.600 379.800 413.400 ;
        RECT 380.400 413.000 389.200 413.800 ;
        RECT 390.000 414.300 390.800 414.400 ;
        RECT 391.600 414.300 392.400 415.800 ;
        RECT 390.000 413.700 392.400 414.300 ;
        RECT 390.000 413.600 390.800 413.700 ;
        RECT 364.400 412.000 365.200 412.600 ;
        RECT 382.000 412.000 382.800 412.400 ;
        RECT 385.200 412.000 386.000 412.400 ;
        RECT 387.000 412.000 387.800 412.200 ;
        RECT 357.600 411.400 358.400 412.000 ;
        RECT 364.400 411.400 387.800 412.000 ;
        RECT 350.000 402.200 350.800 410.200 ;
        RECT 351.800 409.600 354.000 410.200 ;
        RECT 356.200 410.000 357.200 410.800 ;
        RECT 353.200 402.200 354.000 409.600 ;
        RECT 356.400 402.200 357.200 410.000 ;
        RECT 357.800 409.600 358.400 411.400 ;
        RECT 359.000 410.800 359.800 411.000 ;
        RECT 359.000 410.300 386.000 410.800 ;
        RECT 386.800 410.300 387.600 410.400 ;
        RECT 359.000 410.200 387.600 410.300 ;
        RECT 381.800 410.000 382.600 410.200 ;
        RECT 385.200 409.700 387.600 410.200 ;
        RECT 385.200 409.600 386.000 409.700 ;
        RECT 386.800 409.600 387.600 409.700 ;
        RECT 357.800 409.000 366.800 409.600 ;
        RECT 357.800 407.400 358.400 409.000 ;
        RECT 366.000 408.800 366.800 409.000 ;
        RECT 369.200 409.000 377.800 409.600 ;
        RECT 369.200 408.800 370.000 409.000 ;
        RECT 361.000 407.600 363.600 408.400 ;
        RECT 357.800 406.800 360.400 407.400 ;
        RECT 359.600 402.200 360.400 406.800 ;
        RECT 362.800 402.200 363.600 407.600 ;
        RECT 364.200 406.800 368.400 407.600 ;
        RECT 366.000 402.200 366.800 405.000 ;
        RECT 367.600 402.200 368.400 405.000 ;
        RECT 369.200 402.200 370.000 405.000 ;
        RECT 370.800 402.200 371.600 408.400 ;
        RECT 374.000 407.600 376.600 408.400 ;
        RECT 377.200 408.200 377.800 409.000 ;
        RECT 378.800 409.400 379.600 409.600 ;
        RECT 378.800 409.000 384.200 409.400 ;
        RECT 378.800 408.800 385.000 409.000 ;
        RECT 383.600 408.200 385.000 408.800 ;
        RECT 377.200 407.600 383.000 408.200 ;
        RECT 386.000 408.000 387.600 408.800 ;
        RECT 386.000 407.600 386.600 408.000 ;
        RECT 374.000 402.200 374.800 407.000 ;
        RECT 377.200 402.200 378.000 407.000 ;
        RECT 382.400 406.800 386.600 407.600 ;
        RECT 388.400 407.400 389.200 413.000 ;
        RECT 387.200 406.800 389.200 407.400 ;
        RECT 378.800 402.200 379.600 405.000 ;
        RECT 380.400 402.200 381.200 405.000 ;
        RECT 383.600 402.200 384.400 406.800 ;
        RECT 387.200 406.200 387.800 406.800 ;
        RECT 386.800 405.600 387.800 406.200 ;
        RECT 386.800 402.200 387.600 405.600 ;
        RECT 391.600 402.200 392.400 413.700 ;
        RECT 394.800 415.800 395.600 419.800 ;
        RECT 398.000 417.800 398.800 419.800 ;
        RECT 394.800 412.400 395.400 415.800 ;
        RECT 398.000 415.600 398.600 417.800 ;
        RECT 399.600 416.300 400.400 417.200 ;
        RECT 401.200 416.300 402.000 416.400 ;
        RECT 399.600 415.700 402.000 416.300 ;
        RECT 402.800 416.000 403.600 419.800 ;
        RECT 399.600 415.600 400.400 415.700 ;
        RECT 401.200 415.600 402.000 415.700 ;
        RECT 396.200 415.000 398.600 415.600 ;
        RECT 402.600 415.200 403.600 416.000 ;
        RECT 393.200 412.300 394.000 412.400 ;
        RECT 394.800 412.300 395.600 412.400 ;
        RECT 393.200 411.700 395.600 412.300 ;
        RECT 393.200 411.600 394.000 411.700 ;
        RECT 394.800 411.600 395.600 411.700 ;
        RECT 396.200 412.000 396.800 415.000 ;
        RECT 394.800 410.200 395.400 411.600 ;
        RECT 396.200 411.400 397.000 412.000 ;
        RECT 396.200 411.200 400.400 411.400 ;
        RECT 396.400 410.800 400.400 411.200 ;
        RECT 394.800 409.600 396.200 410.200 ;
        RECT 395.400 402.200 396.200 409.600 ;
        RECT 399.600 402.200 400.400 410.800 ;
        RECT 402.600 410.800 403.400 415.200 ;
        RECT 404.400 414.600 405.200 419.800 ;
        RECT 410.800 416.600 411.600 419.800 ;
        RECT 412.400 417.000 413.200 419.800 ;
        RECT 414.000 417.000 414.800 419.800 ;
        RECT 415.600 417.000 416.400 419.800 ;
        RECT 417.200 417.000 418.000 419.800 ;
        RECT 420.400 417.000 421.200 419.800 ;
        RECT 423.600 417.000 424.400 419.800 ;
        RECT 425.200 417.000 426.000 419.800 ;
        RECT 426.800 417.000 427.600 419.800 ;
        RECT 409.200 415.800 411.600 416.600 ;
        RECT 428.400 416.600 429.200 419.800 ;
        RECT 409.200 415.200 410.000 415.800 ;
        RECT 404.000 414.000 405.200 414.600 ;
        RECT 408.200 414.600 410.000 415.200 ;
        RECT 414.000 415.600 415.000 416.400 ;
        RECT 418.000 415.600 419.600 416.400 ;
        RECT 420.400 415.800 425.000 416.400 ;
        RECT 428.400 415.800 431.000 416.600 ;
        RECT 420.400 415.600 421.200 415.800 ;
        RECT 404.000 412.000 404.600 414.000 ;
        RECT 408.200 413.400 409.000 414.600 ;
        RECT 405.200 412.600 409.000 413.400 ;
        RECT 414.000 412.800 414.800 415.600 ;
        RECT 420.400 414.800 421.200 415.000 ;
        RECT 416.800 414.200 421.200 414.800 ;
        RECT 416.800 414.000 417.600 414.200 ;
        RECT 424.200 413.400 425.000 415.800 ;
        RECT 430.200 415.200 431.000 415.800 ;
        RECT 430.200 414.400 433.200 415.200 ;
        RECT 434.800 413.800 435.600 419.800 ;
        RECT 437.000 416.400 437.800 419.800 ;
        RECT 437.000 415.800 438.800 416.400 ;
        RECT 417.200 412.600 420.400 413.400 ;
        RECT 424.200 412.600 426.200 413.400 ;
        RECT 426.800 413.000 435.600 413.800 ;
        RECT 436.400 414.300 437.200 414.400 ;
        RECT 438.000 414.300 438.800 415.800 ;
        RECT 436.400 413.700 438.800 414.300 ;
        RECT 436.400 413.600 437.200 413.700 ;
        RECT 410.800 412.000 411.600 412.600 ;
        RECT 428.400 412.000 429.200 412.400 ;
        RECT 431.600 412.000 432.400 412.400 ;
        RECT 433.400 412.000 434.200 412.200 ;
        RECT 404.000 411.400 404.800 412.000 ;
        RECT 410.800 411.400 434.200 412.000 ;
        RECT 402.600 410.000 403.600 410.800 ;
        RECT 402.800 402.200 403.600 410.000 ;
        RECT 404.200 409.600 404.800 411.400 ;
        RECT 405.400 410.800 406.200 411.000 ;
        RECT 405.400 410.300 432.400 410.800 ;
        RECT 433.200 410.300 434.000 410.400 ;
        RECT 405.400 410.200 434.000 410.300 ;
        RECT 428.200 410.000 429.000 410.200 ;
        RECT 431.600 409.700 434.000 410.200 ;
        RECT 431.600 409.600 432.400 409.700 ;
        RECT 433.200 409.600 434.000 409.700 ;
        RECT 404.200 409.000 413.200 409.600 ;
        RECT 404.200 407.400 404.800 409.000 ;
        RECT 412.400 408.800 413.200 409.000 ;
        RECT 415.600 409.000 424.200 409.600 ;
        RECT 415.600 408.800 416.400 409.000 ;
        RECT 407.400 407.600 410.000 408.400 ;
        RECT 404.200 406.800 406.800 407.400 ;
        RECT 406.000 402.200 406.800 406.800 ;
        RECT 409.200 402.200 410.000 407.600 ;
        RECT 410.600 406.800 414.800 407.600 ;
        RECT 412.400 402.200 413.200 405.000 ;
        RECT 414.000 402.200 414.800 405.000 ;
        RECT 415.600 402.200 416.400 405.000 ;
        RECT 417.200 402.200 418.000 408.400 ;
        RECT 420.400 407.600 423.000 408.400 ;
        RECT 423.600 408.200 424.200 409.000 ;
        RECT 425.200 409.400 426.000 409.600 ;
        RECT 425.200 409.000 430.600 409.400 ;
        RECT 425.200 408.800 431.400 409.000 ;
        RECT 430.000 408.200 431.400 408.800 ;
        RECT 423.600 407.600 429.400 408.200 ;
        RECT 432.400 408.000 434.000 408.800 ;
        RECT 432.400 407.600 433.000 408.000 ;
        RECT 420.400 402.200 421.200 407.000 ;
        RECT 423.600 402.200 424.400 407.000 ;
        RECT 428.800 406.800 433.000 407.600 ;
        RECT 434.800 407.400 435.600 413.000 ;
        RECT 433.600 406.800 435.600 407.400 ;
        RECT 425.200 402.200 426.000 405.000 ;
        RECT 426.800 402.200 427.600 405.000 ;
        RECT 430.000 402.200 430.800 406.800 ;
        RECT 433.600 406.200 434.200 406.800 ;
        RECT 433.200 405.600 434.200 406.200 ;
        RECT 433.200 402.200 434.000 405.600 ;
        RECT 438.000 402.200 438.800 413.700 ;
        RECT 446.000 415.800 446.800 419.800 ;
        RECT 449.200 417.800 450.000 419.800 ;
        RECT 446.000 412.400 446.600 415.800 ;
        RECT 449.200 415.600 449.800 417.800 ;
        RECT 450.800 415.600 451.600 417.200 ;
        RECT 447.400 415.000 449.800 415.600 ;
        RECT 441.200 412.300 442.000 412.400 ;
        RECT 446.000 412.300 446.800 412.400 ;
        RECT 441.200 411.700 446.800 412.300 ;
        RECT 441.200 411.600 442.000 411.700 ;
        RECT 446.000 411.600 446.800 411.700 ;
        RECT 447.400 412.000 448.000 415.000 ;
        RECT 452.400 412.400 453.200 419.800 ;
        RECT 455.600 415.200 456.400 419.800 ;
        RECT 454.200 414.600 456.400 415.200 ;
        RECT 457.200 415.200 458.000 419.800 ;
        RECT 463.600 416.000 464.400 419.800 ;
        RECT 463.400 415.200 464.400 416.000 ;
        RECT 457.200 414.600 459.400 415.200 ;
        RECT 446.000 410.200 446.600 411.600 ;
        RECT 447.400 411.400 448.200 412.000 ;
        RECT 447.400 411.200 451.600 411.400 ;
        RECT 447.600 410.800 451.600 411.200 ;
        RECT 446.000 409.600 447.400 410.200 ;
        RECT 446.600 402.200 447.400 409.600 ;
        RECT 450.800 402.200 451.600 410.800 ;
        RECT 452.400 410.200 453.000 412.400 ;
        RECT 454.200 411.600 454.800 414.600 ;
        RECT 457.200 411.600 458.000 413.200 ;
        RECT 458.800 411.600 459.400 414.600 ;
        RECT 453.600 410.800 454.800 411.600 ;
        RECT 454.200 410.200 454.800 410.800 ;
        RECT 458.800 410.800 460.000 411.600 ;
        RECT 463.400 410.800 464.200 415.200 ;
        RECT 465.200 414.600 466.000 419.800 ;
        RECT 471.600 416.600 472.400 419.800 ;
        RECT 473.200 417.000 474.000 419.800 ;
        RECT 474.800 417.000 475.600 419.800 ;
        RECT 476.400 417.000 477.200 419.800 ;
        RECT 478.000 417.000 478.800 419.800 ;
        RECT 481.200 417.000 482.000 419.800 ;
        RECT 484.400 417.000 485.200 419.800 ;
        RECT 486.000 417.000 486.800 419.800 ;
        RECT 487.600 417.000 488.400 419.800 ;
        RECT 470.000 415.800 472.400 416.600 ;
        RECT 489.200 416.600 490.000 419.800 ;
        RECT 470.000 415.200 470.800 415.800 ;
        RECT 464.800 414.000 466.000 414.600 ;
        RECT 469.000 414.600 470.800 415.200 ;
        RECT 474.800 415.600 475.800 416.400 ;
        RECT 478.800 415.600 480.400 416.400 ;
        RECT 481.200 415.800 485.800 416.400 ;
        RECT 489.200 415.800 491.800 416.600 ;
        RECT 481.200 415.600 482.000 415.800 ;
        RECT 464.800 412.000 465.400 414.000 ;
        RECT 469.000 413.400 469.800 414.600 ;
        RECT 466.000 412.600 469.800 413.400 ;
        RECT 474.800 412.800 475.600 415.600 ;
        RECT 481.200 414.800 482.000 415.000 ;
        RECT 477.600 414.200 482.000 414.800 ;
        RECT 477.600 414.000 478.400 414.200 ;
        RECT 485.000 413.400 485.800 415.800 ;
        RECT 491.000 415.200 491.800 415.800 ;
        RECT 491.000 414.400 494.000 415.200 ;
        RECT 495.600 413.800 496.400 419.800 ;
        RECT 497.800 416.400 498.600 419.800 ;
        RECT 497.800 415.800 499.600 416.400 ;
        RECT 478.000 412.600 481.200 413.400 ;
        RECT 485.000 412.600 487.000 413.400 ;
        RECT 487.600 413.000 496.400 413.800 ;
        RECT 497.200 414.300 498.000 414.400 ;
        RECT 498.800 414.300 499.600 415.800 ;
        RECT 497.200 413.700 499.600 414.300 ;
        RECT 497.200 413.600 498.000 413.700 ;
        RECT 471.600 412.000 472.400 412.600 ;
        RECT 489.200 412.000 490.000 412.400 ;
        RECT 492.400 412.000 493.200 412.400 ;
        RECT 494.200 412.000 495.000 412.200 ;
        RECT 464.800 411.400 465.600 412.000 ;
        RECT 471.600 411.400 495.000 412.000 ;
        RECT 458.800 410.200 459.400 410.800 ;
        RECT 452.400 402.200 453.200 410.200 ;
        RECT 454.200 409.600 456.400 410.200 ;
        RECT 455.600 402.200 456.400 409.600 ;
        RECT 457.200 409.600 459.400 410.200 ;
        RECT 463.400 410.000 464.400 410.800 ;
        RECT 457.200 402.200 458.000 409.600 ;
        RECT 463.600 402.200 464.400 410.000 ;
        RECT 465.000 409.600 465.600 411.400 ;
        RECT 466.200 410.800 467.000 411.000 ;
        RECT 466.200 410.300 493.200 410.800 ;
        RECT 494.000 410.300 494.800 410.400 ;
        RECT 466.200 410.200 494.800 410.300 ;
        RECT 489.000 410.000 489.800 410.200 ;
        RECT 492.400 409.700 494.800 410.200 ;
        RECT 492.400 409.600 493.200 409.700 ;
        RECT 494.000 409.600 494.800 409.700 ;
        RECT 465.000 409.000 474.000 409.600 ;
        RECT 465.000 407.400 465.600 409.000 ;
        RECT 473.200 408.800 474.000 409.000 ;
        RECT 476.400 409.000 485.000 409.600 ;
        RECT 476.400 408.800 477.200 409.000 ;
        RECT 468.200 407.600 470.800 408.400 ;
        RECT 465.000 406.800 467.600 407.400 ;
        RECT 466.800 402.200 467.600 406.800 ;
        RECT 470.000 402.200 470.800 407.600 ;
        RECT 471.400 406.800 475.600 407.600 ;
        RECT 473.200 402.200 474.000 405.000 ;
        RECT 474.800 402.200 475.600 405.000 ;
        RECT 476.400 402.200 477.200 405.000 ;
        RECT 478.000 402.200 478.800 408.400 ;
        RECT 481.200 407.600 483.800 408.400 ;
        RECT 484.400 408.200 485.000 409.000 ;
        RECT 486.000 409.400 486.800 409.600 ;
        RECT 486.000 409.000 491.400 409.400 ;
        RECT 486.000 408.800 492.200 409.000 ;
        RECT 490.800 408.200 492.200 408.800 ;
        RECT 484.400 407.600 490.200 408.200 ;
        RECT 493.200 408.000 494.800 408.800 ;
        RECT 493.200 407.600 493.800 408.000 ;
        RECT 481.200 402.200 482.000 407.000 ;
        RECT 484.400 402.200 485.200 407.000 ;
        RECT 489.600 406.800 493.800 407.600 ;
        RECT 495.600 407.400 496.400 413.000 ;
        RECT 494.400 406.800 496.400 407.400 ;
        RECT 486.000 402.200 486.800 405.000 ;
        RECT 487.600 402.200 488.400 405.000 ;
        RECT 490.800 402.200 491.600 406.800 ;
        RECT 494.400 406.200 495.000 406.800 ;
        RECT 494.000 405.600 495.000 406.200 ;
        RECT 494.000 402.200 494.800 405.600 ;
        RECT 498.800 402.200 499.600 413.700 ;
        RECT 502.000 415.800 502.800 419.800 ;
        RECT 505.200 417.800 506.000 419.800 ;
        RECT 502.000 412.400 502.600 415.800 ;
        RECT 505.200 415.600 505.800 417.800 ;
        RECT 506.800 415.600 507.600 417.200 ;
        RECT 503.400 415.000 505.800 415.600 ;
        RECT 508.400 415.200 509.200 419.800 ;
        RECT 502.000 411.600 502.800 412.400 ;
        RECT 503.400 412.000 504.000 415.000 ;
        RECT 508.400 414.600 510.600 415.200 ;
        RECT 502.000 410.200 502.600 411.600 ;
        RECT 503.400 411.400 504.200 412.000 ;
        RECT 510.000 411.600 510.600 414.600 ;
        RECT 511.600 412.400 512.400 419.800 ;
        RECT 503.400 411.200 507.600 411.400 ;
        RECT 503.600 410.800 507.600 411.200 ;
        RECT 502.000 409.600 503.400 410.200 ;
        RECT 502.600 402.200 503.400 409.600 ;
        RECT 506.800 402.200 507.600 410.800 ;
        RECT 510.000 410.800 511.200 411.600 ;
        RECT 510.000 410.200 510.600 410.800 ;
        RECT 511.800 410.200 512.400 412.400 ;
        RECT 508.400 409.600 510.600 410.200 ;
        RECT 508.400 402.200 509.200 409.600 ;
        RECT 511.600 402.200 512.400 410.200 ;
        RECT 513.200 413.800 514.000 419.800 ;
        RECT 519.600 416.600 520.400 419.800 ;
        RECT 521.200 417.000 522.000 419.800 ;
        RECT 522.800 417.000 523.600 419.800 ;
        RECT 524.400 417.000 525.200 419.800 ;
        RECT 527.600 417.000 528.400 419.800 ;
        RECT 530.800 417.000 531.600 419.800 ;
        RECT 532.400 417.000 533.200 419.800 ;
        RECT 534.000 417.000 534.800 419.800 ;
        RECT 535.600 417.000 536.400 419.800 ;
        RECT 517.800 415.800 520.400 416.600 ;
        RECT 537.200 416.600 538.000 419.800 ;
        RECT 523.800 415.800 528.400 416.400 ;
        RECT 517.800 415.200 518.600 415.800 ;
        RECT 515.600 414.400 518.600 415.200 ;
        RECT 513.200 413.000 522.000 413.800 ;
        RECT 523.800 413.400 524.600 415.800 ;
        RECT 527.600 415.600 528.400 415.800 ;
        RECT 529.200 415.600 530.800 416.400 ;
        RECT 533.800 415.600 534.800 416.400 ;
        RECT 537.200 415.800 539.600 416.600 ;
        RECT 526.000 413.600 526.800 415.200 ;
        RECT 527.600 414.800 528.400 415.000 ;
        RECT 527.600 414.200 532.000 414.800 ;
        RECT 531.200 414.000 532.000 414.200 ;
        RECT 513.200 407.400 514.000 413.000 ;
        RECT 522.600 412.600 524.600 413.400 ;
        RECT 528.400 412.600 531.600 413.400 ;
        RECT 534.000 412.800 534.800 415.600 ;
        RECT 538.800 415.200 539.600 415.800 ;
        RECT 538.800 414.600 540.600 415.200 ;
        RECT 539.800 413.400 540.600 414.600 ;
        RECT 543.600 414.600 544.400 419.800 ;
        RECT 545.200 416.000 546.000 419.800 ;
        RECT 550.000 416.000 550.800 419.800 ;
        RECT 545.200 415.200 546.200 416.000 ;
        RECT 543.600 414.000 544.800 414.600 ;
        RECT 539.800 412.600 543.600 413.400 ;
        RECT 514.800 412.200 515.600 412.400 ;
        RECT 514.600 412.000 515.600 412.200 ;
        RECT 519.600 412.000 520.400 412.400 ;
        RECT 537.200 412.000 538.000 412.600 ;
        RECT 544.200 412.000 544.800 414.000 ;
        RECT 514.600 411.400 538.000 412.000 ;
        RECT 544.000 411.400 544.800 412.000 ;
        RECT 544.000 409.600 544.600 411.400 ;
        RECT 545.400 410.800 546.200 415.200 ;
        RECT 522.800 409.400 523.600 409.600 ;
        RECT 518.200 409.000 523.600 409.400 ;
        RECT 517.400 408.800 523.600 409.000 ;
        RECT 524.600 409.000 533.200 409.600 ;
        RECT 514.800 408.000 516.400 408.800 ;
        RECT 517.400 408.200 518.800 408.800 ;
        RECT 524.600 408.200 525.200 409.000 ;
        RECT 532.400 408.800 533.200 409.000 ;
        RECT 535.600 409.000 544.600 409.600 ;
        RECT 535.600 408.800 536.400 409.000 ;
        RECT 515.800 407.600 516.400 408.000 ;
        RECT 519.400 407.600 525.200 408.200 ;
        RECT 525.800 407.600 528.400 408.400 ;
        RECT 513.200 406.800 515.200 407.400 ;
        RECT 515.800 406.800 520.000 407.600 ;
        RECT 514.600 406.200 515.200 406.800 ;
        RECT 514.600 405.600 515.600 406.200 ;
        RECT 514.800 402.200 515.600 405.600 ;
        RECT 518.000 402.200 518.800 406.800 ;
        RECT 521.200 402.200 522.000 405.000 ;
        RECT 522.800 402.200 523.600 405.000 ;
        RECT 524.400 402.200 525.200 407.000 ;
        RECT 527.600 402.200 528.400 407.000 ;
        RECT 530.800 402.200 531.600 408.400 ;
        RECT 538.800 407.600 541.400 408.400 ;
        RECT 534.000 406.800 538.200 407.600 ;
        RECT 532.400 402.200 533.200 405.000 ;
        RECT 534.000 402.200 534.800 405.000 ;
        RECT 535.600 402.200 536.400 405.000 ;
        RECT 538.800 402.200 539.600 407.600 ;
        RECT 544.000 407.400 544.600 409.000 ;
        RECT 542.000 406.800 544.600 407.400 ;
        RECT 545.200 410.000 546.200 410.800 ;
        RECT 549.800 415.200 550.800 416.000 ;
        RECT 549.800 410.800 550.600 415.200 ;
        RECT 551.600 414.600 552.400 419.800 ;
        RECT 558.000 416.600 558.800 419.800 ;
        RECT 559.600 417.000 560.400 419.800 ;
        RECT 561.200 417.000 562.000 419.800 ;
        RECT 562.800 417.000 563.600 419.800 ;
        RECT 564.400 417.000 565.200 419.800 ;
        RECT 567.600 417.000 568.400 419.800 ;
        RECT 570.800 417.000 571.600 419.800 ;
        RECT 572.400 417.000 573.200 419.800 ;
        RECT 574.000 417.000 574.800 419.800 ;
        RECT 556.400 415.800 558.800 416.600 ;
        RECT 575.600 416.600 576.400 419.800 ;
        RECT 556.400 415.200 557.200 415.800 ;
        RECT 551.200 414.000 552.400 414.600 ;
        RECT 555.400 414.600 557.200 415.200 ;
        RECT 561.200 415.600 562.200 416.400 ;
        RECT 565.200 415.600 566.800 416.400 ;
        RECT 567.600 415.800 572.200 416.400 ;
        RECT 575.600 415.800 578.200 416.600 ;
        RECT 567.600 415.600 568.400 415.800 ;
        RECT 551.200 412.000 551.800 414.000 ;
        RECT 555.400 413.400 556.200 414.600 ;
        RECT 552.400 412.600 556.200 413.400 ;
        RECT 561.200 412.800 562.000 415.600 ;
        RECT 567.600 414.800 568.400 415.000 ;
        RECT 564.000 414.200 568.400 414.800 ;
        RECT 564.000 414.000 564.800 414.200 ;
        RECT 569.200 413.600 570.000 415.200 ;
        RECT 571.400 413.400 572.200 415.800 ;
        RECT 577.400 415.200 578.200 415.800 ;
        RECT 577.400 414.400 580.400 415.200 ;
        RECT 582.000 413.800 582.800 419.800 ;
        RECT 564.400 412.600 567.600 413.400 ;
        RECT 571.400 412.600 573.400 413.400 ;
        RECT 574.000 413.000 582.800 413.800 ;
        RECT 558.000 412.000 558.800 412.600 ;
        RECT 575.600 412.000 576.400 412.400 ;
        RECT 580.600 412.000 581.400 412.200 ;
        RECT 551.200 411.400 552.000 412.000 ;
        RECT 558.000 411.400 581.400 412.000 ;
        RECT 549.800 410.000 550.800 410.800 ;
        RECT 542.000 402.200 542.800 406.800 ;
        RECT 545.200 402.200 546.000 410.000 ;
        RECT 550.000 402.200 550.800 410.000 ;
        RECT 551.400 409.600 552.000 411.400 ;
        RECT 551.400 409.000 560.400 409.600 ;
        RECT 551.400 407.400 552.000 409.000 ;
        RECT 559.600 408.800 560.400 409.000 ;
        RECT 562.800 409.000 571.400 409.600 ;
        RECT 562.800 408.800 563.600 409.000 ;
        RECT 554.600 407.600 557.200 408.400 ;
        RECT 551.400 406.800 554.000 407.400 ;
        RECT 553.200 402.200 554.000 406.800 ;
        RECT 556.400 402.200 557.200 407.600 ;
        RECT 557.800 406.800 562.000 407.600 ;
        RECT 559.600 402.200 560.400 405.000 ;
        RECT 561.200 402.200 562.000 405.000 ;
        RECT 562.800 402.200 563.600 405.000 ;
        RECT 564.400 402.200 565.200 408.400 ;
        RECT 567.600 407.600 570.200 408.400 ;
        RECT 570.800 408.200 571.400 409.000 ;
        RECT 572.400 409.400 573.200 409.600 ;
        RECT 572.400 409.000 577.800 409.400 ;
        RECT 572.400 408.800 578.600 409.000 ;
        RECT 577.200 408.200 578.600 408.800 ;
        RECT 570.800 407.600 576.600 408.200 ;
        RECT 579.600 408.000 581.200 408.800 ;
        RECT 579.600 407.600 580.200 408.000 ;
        RECT 567.600 402.200 568.400 407.000 ;
        RECT 570.800 402.200 571.600 407.000 ;
        RECT 576.000 406.800 580.200 407.600 ;
        RECT 582.000 407.400 582.800 413.000 ;
        RECT 580.800 406.800 582.800 407.400 ;
        RECT 572.400 402.200 573.200 405.000 ;
        RECT 574.000 402.200 574.800 405.000 ;
        RECT 577.200 402.200 578.000 406.800 ;
        RECT 580.800 406.200 581.400 406.800 ;
        RECT 580.400 405.600 581.400 406.200 ;
        RECT 580.400 402.200 581.200 405.600 ;
        RECT 3.800 392.400 4.600 399.800 ;
        RECT 5.200 393.600 6.000 394.400 ;
        RECT 5.400 392.400 6.000 393.600 ;
        RECT 3.800 391.800 4.800 392.400 ;
        RECT 5.400 392.300 6.800 392.400 ;
        RECT 9.200 392.300 10.000 399.800 ;
        RECT 5.400 391.800 10.000 392.300 ;
        RECT 2.800 388.800 3.600 390.400 ;
        RECT 4.200 388.400 4.800 391.800 ;
        RECT 6.000 391.700 10.000 391.800 ;
        RECT 6.000 391.600 6.800 391.700 ;
        RECT 1.200 388.200 2.000 388.400 ;
        RECT 1.200 387.600 2.800 388.200 ;
        RECT 4.200 387.600 6.800 388.400 ;
        RECT 2.000 387.200 2.800 387.600 ;
        RECT 1.400 386.200 5.000 386.600 ;
        RECT 6.000 386.200 6.600 387.600 ;
        RECT 7.600 386.800 8.400 388.400 ;
        RECT 9.200 386.200 10.000 391.700 ;
        RECT 10.800 391.600 11.600 393.200 ;
        RECT 12.400 391.600 13.200 393.200 ;
        RECT 14.000 392.300 14.800 399.800 ;
        RECT 17.200 392.300 18.000 393.200 ;
        RECT 14.000 391.700 18.000 392.300 ;
        RECT 14.000 386.200 14.800 391.700 ;
        RECT 17.200 391.600 18.000 391.700 ;
        RECT 18.800 392.300 19.600 399.800 ;
        RECT 22.000 392.300 22.800 392.400 ;
        RECT 18.800 391.700 22.800 392.300 ;
        RECT 15.600 386.800 16.400 388.400 ;
        RECT 18.800 386.200 19.600 391.700 ;
        RECT 22.000 391.600 22.800 391.700 ;
        RECT 20.400 386.800 21.200 388.400 ;
        RECT 22.000 386.800 22.800 388.400 ;
        RECT 1.200 386.000 5.200 386.200 ;
        RECT 1.200 382.200 2.000 386.000 ;
        RECT 4.400 382.200 5.200 386.000 ;
        RECT 6.000 382.200 6.800 386.200 ;
        RECT 9.200 385.600 11.000 386.200 ;
        RECT 10.200 382.200 11.000 385.600 ;
        RECT 13.000 385.600 14.800 386.200 ;
        RECT 17.800 385.600 19.600 386.200 ;
        RECT 23.600 386.200 24.400 399.800 ;
        RECT 25.200 391.600 26.000 393.200 ;
        RECT 27.400 392.600 28.200 399.800 ;
        RECT 27.400 391.800 29.200 392.600 ;
        RECT 31.600 392.400 32.400 399.800 ;
        RECT 34.800 392.400 35.600 399.800 ;
        RECT 31.600 391.800 35.600 392.400 ;
        RECT 36.400 391.800 37.200 399.800 ;
        RECT 38.800 393.600 39.600 394.400 ;
        RECT 38.800 392.400 39.400 393.600 ;
        RECT 40.200 392.400 41.000 399.800 ;
        RECT 38.000 391.800 39.400 392.400 ;
        RECT 25.300 390.300 25.900 391.600 ;
        RECT 26.800 390.300 27.600 391.200 ;
        RECT 25.300 389.700 27.600 390.300 ;
        RECT 26.800 389.600 27.600 389.700 ;
        RECT 28.400 390.300 29.000 391.800 ;
        RECT 32.400 390.400 33.200 390.800 ;
        RECT 36.400 390.400 37.000 391.800 ;
        RECT 38.000 391.600 38.800 391.800 ;
        RECT 40.000 391.600 42.000 392.400 ;
        RECT 44.400 391.600 45.200 393.200 ;
        RECT 31.600 390.300 33.200 390.400 ;
        RECT 28.400 389.800 33.200 390.300 ;
        RECT 34.800 389.800 37.200 390.400 ;
        RECT 28.400 389.700 32.400 389.800 ;
        RECT 28.400 388.400 29.000 389.700 ;
        RECT 31.600 389.600 32.400 389.700 ;
        RECT 28.400 387.600 29.200 388.400 ;
        RECT 33.200 387.600 34.000 389.200 ;
        RECT 23.600 385.600 25.400 386.200 ;
        RECT 13.000 382.200 13.800 385.600 ;
        RECT 17.800 382.200 18.600 385.600 ;
        RECT 24.600 384.400 25.400 385.600 ;
        RECT 23.600 383.600 25.400 384.400 ;
        RECT 24.600 382.200 25.400 383.600 ;
        RECT 28.400 384.200 29.000 387.600 ;
        RECT 30.000 384.800 30.800 386.400 ;
        RECT 34.800 386.200 35.400 389.800 ;
        RECT 36.400 389.600 37.200 389.800 ;
        RECT 40.000 388.400 40.600 391.600 ;
        RECT 41.200 388.800 42.000 390.400 ;
        RECT 38.000 387.600 40.600 388.400 ;
        RECT 42.800 388.200 43.600 388.400 ;
        RECT 42.000 387.600 43.600 388.200 ;
        RECT 28.400 382.200 29.200 384.200 ;
        RECT 34.800 382.200 35.600 386.200 ;
        RECT 36.400 385.600 37.200 386.400 ;
        RECT 38.200 386.200 38.800 387.600 ;
        RECT 42.000 387.200 42.800 387.600 ;
        RECT 39.800 386.200 43.400 386.600 ;
        RECT 46.000 386.200 46.800 399.800 ;
        RECT 47.600 386.800 48.400 388.400 ;
        RECT 49.200 386.800 50.000 388.400 ;
        RECT 50.800 388.300 51.600 399.800 ;
        RECT 52.400 391.600 53.200 393.200 ;
        RECT 54.600 392.600 55.400 399.800 ;
        RECT 54.600 391.800 56.400 392.600 ;
        RECT 58.800 391.800 59.600 399.800 ;
        RECT 60.400 392.400 61.200 399.800 ;
        RECT 63.600 392.400 64.400 399.800 ;
        RECT 60.400 391.800 64.400 392.400 ;
        RECT 65.200 392.400 66.000 399.800 ;
        RECT 66.800 392.400 67.600 392.600 ;
        RECT 65.200 391.800 67.600 392.400 ;
        RECT 69.600 391.800 71.200 399.800 ;
        RECT 73.000 392.400 73.800 392.600 ;
        RECT 74.800 392.400 75.600 399.800 ;
        RECT 73.000 391.800 75.600 392.400 ;
        RECT 54.000 389.600 54.800 391.200 ;
        RECT 55.600 388.400 56.200 391.800 ;
        RECT 59.000 390.400 59.600 391.800 ;
        RECT 62.800 390.400 63.600 390.800 ;
        RECT 70.000 390.400 70.600 391.800 ;
        RECT 71.800 390.400 72.600 390.600 ;
        RECT 58.800 389.800 61.200 390.400 ;
        RECT 62.800 389.800 64.400 390.400 ;
        RECT 58.800 389.600 59.600 389.800 ;
        RECT 54.000 388.300 54.800 388.400 ;
        RECT 50.800 387.700 54.800 388.300 ;
        RECT 36.200 384.800 37.000 385.600 ;
        RECT 38.000 382.200 38.800 386.200 ;
        RECT 39.600 386.000 43.600 386.200 ;
        RECT 39.600 382.200 40.400 386.000 ;
        RECT 42.800 382.200 43.600 386.000 ;
        RECT 45.000 385.600 46.800 386.200 ;
        RECT 50.800 386.200 51.600 387.700 ;
        RECT 54.000 387.600 54.800 387.700 ;
        RECT 55.600 388.300 56.400 388.400 ;
        RECT 55.600 387.700 59.500 388.300 ;
        RECT 55.600 387.600 56.400 387.700 ;
        RECT 50.800 385.600 52.600 386.200 ;
        RECT 45.000 384.400 45.800 385.600 ;
        RECT 44.400 383.600 45.800 384.400 ;
        RECT 45.000 382.200 45.800 383.600 ;
        RECT 51.800 382.200 52.600 385.600 ;
        RECT 55.600 384.200 56.200 387.600 ;
        RECT 58.900 386.400 59.500 387.700 ;
        RECT 57.200 384.800 58.000 386.400 ;
        RECT 58.800 385.600 59.600 386.400 ;
        RECT 60.600 386.200 61.200 389.800 ;
        RECT 63.600 389.600 64.400 389.800 ;
        RECT 70.000 389.600 70.800 390.400 ;
        RECT 71.800 389.800 73.400 390.400 ;
        RECT 72.600 389.600 73.400 389.800 ;
        RECT 78.000 390.300 78.800 399.800 ;
        RECT 82.200 392.400 83.000 399.800 ;
        RECT 83.600 393.600 84.400 394.400 ;
        RECT 83.800 392.400 84.400 393.600 ;
        RECT 86.800 393.600 87.600 394.400 ;
        RECT 86.800 392.400 87.400 393.600 ;
        RECT 88.200 392.400 89.000 399.800 ;
        RECT 82.200 391.800 83.200 392.400 ;
        RECT 83.800 391.800 85.200 392.400 ;
        RECT 81.200 390.300 82.000 390.400 ;
        RECT 78.000 389.700 82.000 390.300 ;
        RECT 62.000 387.600 62.800 389.200 ;
        RECT 70.000 388.400 70.600 389.600 ;
        RECT 63.600 388.300 64.400 388.400 ;
        RECT 65.200 388.300 66.800 388.400 ;
        RECT 63.600 387.700 66.800 388.300 ;
        RECT 63.600 387.600 64.400 387.700 ;
        RECT 65.200 387.600 66.800 387.700 ;
        RECT 68.000 387.600 68.800 388.400 ;
        RECT 68.200 387.200 68.800 387.600 ;
        RECT 69.600 387.800 70.600 388.400 ;
        RECT 71.200 388.600 72.000 388.800 ;
        RECT 71.200 388.400 74.000 388.600 ;
        RECT 71.200 388.000 75.600 388.400 ;
        RECT 73.400 387.800 75.600 388.000 ;
        RECT 66.800 386.800 67.600 387.000 ;
        RECT 59.000 384.800 59.800 385.600 ;
        RECT 55.600 382.200 56.400 384.200 ;
        RECT 60.400 382.200 61.200 386.200 ;
        RECT 65.200 386.200 67.600 386.800 ;
        RECT 68.200 386.400 69.000 387.200 ;
        RECT 65.200 382.200 66.000 386.200 ;
        RECT 69.600 385.800 70.200 387.800 ;
        RECT 74.000 387.600 75.600 387.800 ;
        RECT 70.800 386.400 72.400 387.200 ;
        RECT 73.000 386.800 73.800 387.000 ;
        RECT 73.000 386.200 75.600 386.800 ;
        RECT 69.600 382.200 71.200 385.800 ;
        RECT 74.800 382.200 75.600 386.200 ;
        RECT 76.400 384.800 77.200 386.400 ;
        RECT 78.000 382.200 78.800 389.700 ;
        RECT 81.200 388.800 82.000 389.700 ;
        RECT 82.600 388.400 83.200 391.800 ;
        RECT 84.400 391.600 85.200 391.800 ;
        RECT 86.000 391.800 87.400 392.400 ;
        RECT 88.000 391.800 89.000 392.400 ;
        RECT 86.000 391.600 86.800 391.800 ;
        RECT 84.500 390.300 85.100 391.600 ;
        RECT 88.000 390.300 88.600 391.800 ;
        RECT 92.400 391.600 93.200 393.200 ;
        RECT 84.500 389.700 88.600 390.300 ;
        RECT 88.000 388.400 88.600 389.700 ;
        RECT 89.200 388.800 90.000 390.400 ;
        RECT 79.600 388.200 80.400 388.400 ;
        RECT 79.600 387.600 81.200 388.200 ;
        RECT 82.600 387.600 85.200 388.400 ;
        RECT 86.000 387.600 88.600 388.400 ;
        RECT 90.800 388.300 91.600 388.400 ;
        RECT 92.400 388.300 93.200 388.400 ;
        RECT 90.800 388.200 93.200 388.300 ;
        RECT 90.000 387.700 93.200 388.200 ;
        RECT 90.000 387.600 91.600 387.700 ;
        RECT 92.400 387.600 93.200 387.700 ;
        RECT 80.400 387.200 81.200 387.600 ;
        RECT 79.800 386.200 83.400 386.600 ;
        RECT 84.400 386.200 85.000 387.600 ;
        RECT 86.200 386.200 86.800 387.600 ;
        RECT 90.000 387.200 90.800 387.600 ;
        RECT 87.800 386.200 91.400 386.600 ;
        RECT 94.000 386.200 94.800 399.800 ;
        RECT 97.200 391.600 98.000 393.200 ;
        RECT 95.600 388.300 96.400 388.400 ;
        RECT 98.800 388.300 99.600 399.800 ;
        RECT 103.600 392.300 104.400 399.800 ;
        RECT 105.200 392.300 106.000 393.200 ;
        RECT 103.600 391.700 106.000 392.300 ;
        RECT 95.600 387.700 99.600 388.300 ;
        RECT 95.600 386.800 96.400 387.700 ;
        RECT 98.800 386.200 99.600 387.700 ;
        RECT 100.400 388.300 101.200 388.400 ;
        RECT 100.400 387.700 102.700 388.300 ;
        RECT 100.400 386.800 101.200 387.700 ;
        RECT 102.100 386.400 102.700 387.700 ;
        RECT 79.600 386.000 83.600 386.200 ;
        RECT 79.600 382.200 80.400 386.000 ;
        RECT 82.800 382.200 83.600 386.000 ;
        RECT 84.400 382.200 85.200 386.200 ;
        RECT 86.000 382.200 86.800 386.200 ;
        RECT 87.600 386.000 91.600 386.200 ;
        RECT 87.600 382.200 88.400 386.000 ;
        RECT 90.800 382.200 91.600 386.000 ;
        RECT 93.000 385.600 94.800 386.200 ;
        RECT 97.800 385.600 99.600 386.200 ;
        RECT 93.000 384.400 93.800 385.600 ;
        RECT 93.000 383.600 94.800 384.400 ;
        RECT 93.000 382.200 93.800 383.600 ;
        RECT 97.800 382.200 98.600 385.600 ;
        RECT 102.000 384.800 102.800 386.400 ;
        RECT 103.600 382.200 104.400 391.700 ;
        RECT 105.200 391.600 106.000 391.700 ;
        RECT 105.200 390.300 106.000 390.400 ;
        RECT 106.800 390.300 107.600 399.800 ;
        RECT 108.400 392.300 109.200 392.400 ;
        RECT 110.000 392.300 110.800 399.800 ;
        RECT 108.400 391.700 110.800 392.300 ;
        RECT 108.400 391.600 109.200 391.700 ;
        RECT 105.200 389.700 107.600 390.300 ;
        RECT 105.200 389.600 106.000 389.700 ;
        RECT 106.800 386.200 107.600 389.700 ;
        RECT 108.400 386.800 109.200 388.400 ;
        RECT 105.800 385.600 107.600 386.200 ;
        RECT 105.800 382.200 106.600 385.600 ;
        RECT 110.000 382.200 110.800 391.700 ;
        RECT 113.200 391.200 114.000 399.800 ;
        RECT 117.400 395.800 118.600 399.800 ;
        RECT 122.000 395.800 122.800 399.800 ;
        RECT 126.400 396.400 127.200 399.800 ;
        RECT 126.400 395.800 128.400 396.400 ;
        RECT 118.000 395.000 118.800 395.800 ;
        RECT 122.200 395.200 122.800 395.800 ;
        RECT 121.400 394.600 125.000 395.200 ;
        RECT 127.600 395.000 128.400 395.800 ;
        RECT 121.400 394.400 122.200 394.600 ;
        RECT 124.200 394.400 125.000 394.600 ;
        RECT 117.200 393.200 118.600 394.000 ;
        RECT 118.000 392.200 118.600 393.200 ;
        RECT 120.200 393.000 122.400 393.600 ;
        RECT 120.200 392.800 121.000 393.000 ;
        RECT 118.000 391.600 120.400 392.200 ;
        RECT 113.200 390.600 117.400 391.200 ;
        RECT 113.200 387.200 114.000 390.600 ;
        RECT 116.600 390.400 117.400 390.600 ;
        RECT 119.800 390.400 120.400 391.600 ;
        RECT 121.800 391.800 122.400 393.000 ;
        RECT 123.000 393.000 123.800 393.200 ;
        RECT 127.600 393.000 128.400 393.200 ;
        RECT 123.000 392.400 128.400 393.000 ;
        RECT 121.800 391.400 126.600 391.800 ;
        RECT 130.800 391.400 131.600 399.800 ;
        RECT 137.200 392.400 138.000 399.800 ;
        RECT 141.600 394.400 143.200 399.800 ;
        RECT 140.400 393.600 143.200 394.400 ;
        RECT 138.600 392.400 139.400 392.600 ;
        RECT 137.200 391.800 139.400 392.400 ;
        RECT 141.600 392.400 143.200 393.600 ;
        RECT 145.200 392.400 146.000 392.600 ;
        RECT 146.800 392.400 147.600 399.800 ;
        RECT 141.600 391.800 143.600 392.400 ;
        RECT 145.200 391.800 147.600 392.400 ;
        RECT 148.400 392.400 149.200 399.800 ;
        RECT 149.800 392.400 150.600 392.600 ;
        RECT 148.400 391.800 150.600 392.400 ;
        RECT 152.800 392.400 154.400 399.800 ;
        RECT 156.400 392.400 157.200 392.600 ;
        RECT 158.000 392.400 158.800 399.800 ;
        RECT 152.800 391.800 154.800 392.400 ;
        RECT 156.400 391.800 158.800 392.400 ;
        RECT 162.200 392.400 163.000 399.800 ;
        RECT 163.600 393.600 164.400 394.400 ;
        RECT 163.800 392.400 164.400 393.600 ;
        RECT 166.800 393.600 167.600 394.400 ;
        RECT 166.800 392.400 167.400 393.600 ;
        RECT 168.200 392.400 169.000 399.800 ;
        RECT 162.200 391.800 163.200 392.400 ;
        RECT 163.800 391.800 165.200 392.400 ;
        RECT 121.800 391.200 131.600 391.400 ;
        RECT 125.800 391.000 131.600 391.200 ;
        RECT 126.000 390.800 131.600 391.000 ;
        RECT 138.800 391.200 139.400 391.800 ;
        RECT 138.800 390.600 142.200 391.200 ;
        RECT 141.400 390.400 142.200 390.600 ;
        RECT 143.000 390.400 143.600 391.800 ;
        RECT 150.000 391.200 150.600 391.800 ;
        RECT 150.000 390.600 153.400 391.200 ;
        RECT 152.600 390.400 153.400 390.600 ;
        RECT 154.200 390.400 154.800 391.800 ;
        RECT 115.000 389.800 115.800 390.000 ;
        RECT 115.000 389.200 118.800 389.800 ;
        RECT 119.600 389.600 120.400 390.400 ;
        RECT 124.400 390.200 125.200 390.400 ;
        RECT 124.400 389.600 129.400 390.200 ;
        RECT 118.000 389.000 118.800 389.200 ;
        RECT 119.800 388.400 120.400 389.600 ;
        RECT 126.000 389.400 126.800 389.600 ;
        RECT 128.600 389.400 129.400 389.600 ;
        RECT 139.200 389.800 140.000 390.000 ;
        RECT 143.000 389.800 144.400 390.400 ;
        RECT 139.200 389.200 141.800 389.800 ;
        RECT 141.200 388.600 141.800 389.200 ;
        RECT 142.600 389.600 144.400 389.800 ;
        RECT 150.400 389.800 151.200 390.000 ;
        RECT 154.200 389.800 155.600 390.400 ;
        RECT 142.600 389.200 143.600 389.600 ;
        RECT 150.400 389.200 153.000 389.800 ;
        RECT 127.000 388.400 127.800 388.600 ;
        RECT 119.800 387.800 130.800 388.400 ;
        RECT 120.200 387.600 121.000 387.800 ;
        RECT 113.200 386.600 117.000 387.200 ;
        RECT 111.600 384.800 112.400 386.400 ;
        RECT 113.200 382.200 114.000 386.600 ;
        RECT 116.200 386.400 117.000 386.600 ;
        RECT 126.000 385.600 126.600 387.800 ;
        RECT 129.200 387.600 130.800 387.800 ;
        RECT 137.200 388.200 138.800 388.400 ;
        RECT 137.200 387.600 140.600 388.200 ;
        RECT 141.200 387.800 142.000 388.600 ;
        RECT 140.000 387.200 140.600 387.600 ;
        RECT 124.200 385.400 125.000 385.600 ;
        RECT 118.000 384.200 118.800 385.000 ;
        RECT 122.200 384.800 125.000 385.400 ;
        RECT 126.000 384.800 126.800 385.600 ;
        RECT 122.200 384.200 122.800 384.800 ;
        RECT 127.600 384.200 128.400 385.000 ;
        RECT 117.400 383.600 118.800 384.200 ;
        RECT 117.400 382.200 118.600 383.600 ;
        RECT 122.000 382.200 122.800 384.200 ;
        RECT 126.400 383.600 128.400 384.200 ;
        RECT 126.400 382.200 127.200 383.600 ;
        RECT 130.800 382.200 131.600 387.000 ;
        RECT 138.600 386.800 139.400 387.000 ;
        RECT 137.200 386.200 139.400 386.800 ;
        RECT 140.000 386.600 142.000 387.200 ;
        RECT 140.400 386.400 142.000 386.600 ;
        RECT 137.200 382.200 138.000 386.200 ;
        RECT 142.600 385.800 143.200 389.200 ;
        RECT 152.400 388.600 153.000 389.200 ;
        RECT 153.800 389.600 155.600 389.800 ;
        RECT 153.800 389.200 154.800 389.600 ;
        RECT 144.000 387.600 144.800 388.400 ;
        RECT 146.000 387.600 147.600 388.400 ;
        RECT 148.400 388.200 150.000 388.400 ;
        RECT 148.400 387.600 151.800 388.200 ;
        RECT 152.400 387.800 153.200 388.600 ;
        RECT 144.000 387.200 144.600 387.600 ;
        RECT 143.800 386.400 144.600 387.200 ;
        RECT 151.200 387.200 151.800 387.600 ;
        RECT 145.200 386.800 146.000 387.000 ;
        RECT 149.800 386.800 150.600 387.000 ;
        RECT 145.200 386.200 147.600 386.800 ;
        RECT 141.600 382.200 143.200 385.800 ;
        RECT 146.800 382.200 147.600 386.200 ;
        RECT 148.400 386.200 150.600 386.800 ;
        RECT 151.200 386.600 153.200 387.200 ;
        RECT 151.600 386.400 153.200 386.600 ;
        RECT 148.400 382.200 149.200 386.200 ;
        RECT 153.800 385.800 154.400 389.200 ;
        RECT 161.200 388.800 162.000 390.400 ;
        RECT 162.600 388.400 163.200 391.800 ;
        RECT 164.400 391.600 165.200 391.800 ;
        RECT 166.000 391.800 167.400 392.400 ;
        RECT 168.000 391.800 169.000 392.400 ;
        RECT 166.000 391.600 166.800 391.800 ;
        RECT 168.000 388.400 168.600 391.800 ;
        RECT 172.400 391.600 173.200 393.200 ;
        RECT 169.200 388.800 170.000 390.400 ;
        RECT 172.400 390.300 173.200 390.400 ;
        RECT 174.000 390.300 174.800 399.800 ;
        RECT 179.800 396.400 180.600 399.800 ;
        RECT 178.800 395.600 180.600 396.400 ;
        RECT 179.800 392.400 180.600 395.600 ;
        RECT 181.200 393.600 182.000 394.400 ;
        RECT 181.400 392.400 182.000 393.600 ;
        RECT 184.400 393.600 185.200 394.400 ;
        RECT 184.400 392.400 185.000 393.600 ;
        RECT 185.800 392.400 186.600 399.800 ;
        RECT 179.800 391.800 180.800 392.400 ;
        RECT 181.400 391.800 182.800 392.400 ;
        RECT 172.400 389.700 174.800 390.300 ;
        RECT 172.400 389.600 173.200 389.700 ;
        RECT 155.200 387.600 156.000 388.400 ;
        RECT 157.200 387.600 158.800 388.400 ;
        RECT 159.600 388.200 160.400 388.400 ;
        RECT 159.600 387.600 161.200 388.200 ;
        RECT 162.600 387.600 165.200 388.400 ;
        RECT 166.000 387.600 168.600 388.400 ;
        RECT 170.800 388.200 171.600 388.400 ;
        RECT 170.000 387.600 171.600 388.200 ;
        RECT 155.200 387.200 155.800 387.600 ;
        RECT 160.400 387.200 161.200 387.600 ;
        RECT 155.000 386.400 155.800 387.200 ;
        RECT 156.400 386.800 157.200 387.000 ;
        RECT 156.400 386.200 158.800 386.800 ;
        RECT 159.800 386.200 163.400 386.600 ;
        RECT 164.400 386.200 165.000 387.600 ;
        RECT 166.200 386.200 166.800 387.600 ;
        RECT 170.000 387.200 170.800 387.600 ;
        RECT 167.800 386.200 171.400 386.600 ;
        RECT 174.000 386.200 174.800 389.700 ;
        RECT 178.800 388.800 179.600 390.400 ;
        RECT 180.200 388.400 180.800 391.800 ;
        RECT 182.000 391.600 182.800 391.800 ;
        RECT 183.600 391.800 185.000 392.400 ;
        RECT 185.600 391.800 186.600 392.400 ;
        RECT 183.600 391.600 184.400 391.800 ;
        RECT 182.100 390.300 182.700 391.600 ;
        RECT 185.600 390.300 186.200 391.800 ;
        RECT 182.100 389.700 186.200 390.300 ;
        RECT 185.600 388.400 186.200 389.700 ;
        RECT 186.800 388.800 187.600 390.400 ;
        RECT 175.600 386.800 176.400 388.400 ;
        RECT 177.200 388.200 178.000 388.400 ;
        RECT 177.200 387.600 178.800 388.200 ;
        RECT 180.200 387.600 182.800 388.400 ;
        RECT 183.600 387.600 186.200 388.400 ;
        RECT 188.400 388.200 189.200 388.400 ;
        RECT 187.600 387.600 189.200 388.200 ;
        RECT 178.000 387.200 178.800 387.600 ;
        RECT 177.400 386.200 181.000 386.600 ;
        RECT 182.000 386.200 182.600 387.600 ;
        RECT 183.800 386.200 184.400 387.600 ;
        RECT 187.600 387.200 188.400 387.600 ;
        RECT 190.000 386.800 190.800 388.400 ;
        RECT 185.400 386.200 189.000 386.600 ;
        RECT 191.600 386.200 192.400 399.800 ;
        RECT 193.200 392.300 194.000 393.200 ;
        RECT 194.800 392.300 195.600 399.800 ;
        RECT 193.200 391.700 195.600 392.300 ;
        RECT 200.600 392.400 201.400 399.800 ;
        RECT 202.000 393.600 202.800 394.400 ;
        RECT 202.200 392.400 202.800 393.600 ;
        RECT 207.000 392.600 207.800 399.800 ;
        RECT 200.600 391.800 201.600 392.400 ;
        RECT 202.200 391.800 203.600 392.400 ;
        RECT 206.000 391.800 207.800 392.600 ;
        RECT 209.200 392.400 210.000 399.800 ;
        RECT 212.400 392.400 213.200 399.800 ;
        RECT 209.200 391.800 213.200 392.400 ;
        RECT 214.000 391.800 214.800 399.800 ;
        RECT 216.200 392.600 217.000 399.800 ;
        RECT 216.200 391.800 218.000 392.600 ;
        RECT 193.200 391.600 194.000 391.700 ;
        RECT 152.800 384.400 154.400 385.800 ;
        RECT 151.600 383.600 154.400 384.400 ;
        RECT 152.800 382.200 154.400 383.600 ;
        RECT 158.000 382.200 158.800 386.200 ;
        RECT 159.600 386.000 163.600 386.200 ;
        RECT 159.600 382.200 160.400 386.000 ;
        RECT 162.800 382.200 163.600 386.000 ;
        RECT 164.400 382.200 165.200 386.200 ;
        RECT 166.000 382.200 166.800 386.200 ;
        RECT 167.600 386.000 171.600 386.200 ;
        RECT 167.600 382.200 168.400 386.000 ;
        RECT 170.800 382.200 171.600 386.000 ;
        RECT 173.000 385.600 174.800 386.200 ;
        RECT 177.200 386.000 181.200 386.200 ;
        RECT 173.000 382.200 173.800 385.600 ;
        RECT 177.200 382.200 178.000 386.000 ;
        RECT 180.400 382.200 181.200 386.000 ;
        RECT 182.000 382.200 182.800 386.200 ;
        RECT 183.600 382.200 184.400 386.200 ;
        RECT 185.200 386.000 189.200 386.200 ;
        RECT 185.200 382.200 186.000 386.000 ;
        RECT 188.400 382.200 189.200 386.000 ;
        RECT 191.600 385.600 193.400 386.200 ;
        RECT 192.600 384.400 193.400 385.600 ;
        RECT 191.600 383.600 193.400 384.400 ;
        RECT 192.600 382.200 193.400 383.600 ;
        RECT 194.800 382.200 195.600 391.700 ;
        RECT 199.600 388.800 200.400 390.400 ;
        RECT 201.000 388.400 201.600 391.800 ;
        RECT 202.800 391.600 203.600 391.800 ;
        RECT 206.200 388.400 206.800 391.800 ;
        RECT 207.600 389.600 208.400 391.200 ;
        RECT 210.000 390.400 210.800 390.800 ;
        RECT 214.000 390.400 214.600 391.800 ;
        RECT 209.200 389.800 210.800 390.400 ;
        RECT 212.400 389.800 214.800 390.400 ;
        RECT 209.200 389.600 210.000 389.800 ;
        RECT 196.400 386.800 197.200 388.400 ;
        RECT 198.000 388.200 198.800 388.400 ;
        RECT 198.000 387.600 199.600 388.200 ;
        RECT 201.000 387.600 203.600 388.400 ;
        RECT 206.000 388.300 206.800 388.400 ;
        RECT 210.800 388.300 211.600 389.200 ;
        RECT 206.000 387.700 211.600 388.300 ;
        RECT 206.000 387.600 206.800 387.700 ;
        RECT 210.800 387.600 211.600 387.700 ;
        RECT 212.400 388.400 213.000 389.800 ;
        RECT 214.000 389.600 214.800 389.800 ;
        RECT 215.600 389.600 216.400 391.200 ;
        RECT 217.200 388.400 217.800 391.800 ;
        RECT 220.400 391.600 221.200 393.200 ;
        RECT 222.000 392.300 222.800 399.800 ;
        RECT 225.200 392.300 226.000 393.200 ;
        RECT 222.000 391.700 226.000 392.300 ;
        RECT 212.400 387.600 213.200 388.400 ;
        RECT 217.200 387.600 218.000 388.400 ;
        RECT 198.800 387.200 199.600 387.600 ;
        RECT 198.200 386.200 201.800 386.600 ;
        RECT 202.800 386.200 203.400 387.600 ;
        RECT 198.000 386.000 202.000 386.200 ;
        RECT 198.000 382.200 198.800 386.000 ;
        RECT 201.200 382.200 202.000 386.000 ;
        RECT 202.800 382.200 203.600 386.200 ;
        RECT 204.400 384.800 205.200 386.400 ;
        RECT 206.200 384.200 206.800 387.600 ;
        RECT 206.000 382.200 206.800 384.200 ;
        RECT 212.400 386.200 213.000 387.600 ;
        RECT 214.000 386.300 214.800 386.400 ;
        RECT 217.200 386.300 217.800 387.600 ;
        RECT 212.400 382.200 213.200 386.200 ;
        RECT 214.000 385.700 217.900 386.300 ;
        RECT 214.000 385.600 214.800 385.700 ;
        RECT 213.800 384.800 214.600 385.600 ;
        RECT 217.200 384.200 217.800 385.700 ;
        RECT 218.800 384.800 219.600 386.400 ;
        RECT 222.000 386.200 222.800 391.700 ;
        RECT 225.200 391.600 226.000 391.700 ;
        RECT 223.600 386.800 224.400 388.400 ;
        RECT 226.800 386.200 227.600 399.800 ;
        RECT 228.400 386.800 229.200 388.400 ;
        RECT 231.600 388.300 232.400 399.800 ;
        RECT 235.800 396.400 236.600 399.800 ;
        RECT 234.800 395.600 236.600 396.400 ;
        RECT 235.800 392.400 236.600 395.600 ;
        RECT 237.200 393.600 238.000 394.400 ;
        RECT 237.400 392.400 238.000 393.600 ;
        RECT 235.800 391.800 236.800 392.400 ;
        RECT 237.400 391.800 238.800 392.400 ;
        RECT 233.200 390.300 234.000 390.400 ;
        RECT 234.800 390.300 235.600 390.400 ;
        RECT 233.200 389.700 235.600 390.300 ;
        RECT 233.200 389.600 234.000 389.700 ;
        RECT 234.800 388.800 235.600 389.700 ;
        RECT 236.200 388.400 236.800 391.800 ;
        RECT 238.000 391.600 238.800 391.800 ;
        RECT 239.600 391.600 240.400 393.200 ;
        RECT 238.100 390.400 238.700 391.600 ;
        RECT 238.000 390.300 238.800 390.400 ;
        RECT 241.200 390.300 242.000 399.800 ;
        RECT 244.400 391.800 245.200 399.800 ;
        RECT 246.000 392.400 246.800 399.800 ;
        RECT 249.200 392.400 250.000 399.800 ;
        RECT 253.400 392.600 254.200 399.800 ;
        RECT 246.000 391.800 250.000 392.400 ;
        RECT 252.400 391.800 254.200 392.600 ;
        RECT 255.600 392.400 256.400 399.800 ;
        RECT 257.000 392.400 257.800 392.600 ;
        RECT 255.600 391.800 257.800 392.400 ;
        RECT 260.000 392.400 261.600 399.800 ;
        RECT 263.600 392.400 264.400 392.600 ;
        RECT 265.200 392.400 266.000 399.800 ;
        RECT 260.000 391.800 262.000 392.400 ;
        RECT 263.600 391.800 266.000 392.400 ;
        RECT 244.600 390.400 245.200 391.800 ;
        RECT 248.400 390.400 249.200 390.800 ;
        RECT 238.000 389.700 242.000 390.300 ;
        RECT 238.000 389.600 238.800 389.700 ;
        RECT 233.200 388.300 234.000 388.400 ;
        RECT 231.600 388.200 234.000 388.300 ;
        RECT 231.600 387.700 234.800 388.200 ;
        RECT 221.000 385.600 222.800 386.200 ;
        RECT 225.800 385.600 227.600 386.200 ;
        RECT 217.200 382.200 218.000 384.200 ;
        RECT 221.000 382.200 221.800 385.600 ;
        RECT 225.800 382.200 226.600 385.600 ;
        RECT 230.000 384.800 230.800 386.400 ;
        RECT 231.600 382.200 232.400 387.700 ;
        RECT 233.200 387.600 234.800 387.700 ;
        RECT 236.200 387.600 238.800 388.400 ;
        RECT 234.000 387.200 234.800 387.600 ;
        RECT 233.400 386.200 237.000 386.600 ;
        RECT 238.000 386.200 238.600 387.600 ;
        RECT 241.200 386.200 242.000 389.700 ;
        RECT 244.400 389.800 246.800 390.400 ;
        RECT 248.400 389.800 250.000 390.400 ;
        RECT 244.400 389.600 245.200 389.800 ;
        RECT 242.800 386.800 243.600 388.400 ;
        RECT 233.200 386.000 237.200 386.200 ;
        RECT 233.200 382.200 234.000 386.000 ;
        RECT 236.400 382.200 237.200 386.000 ;
        RECT 238.000 382.200 238.800 386.200 ;
        RECT 240.200 385.600 242.000 386.200 ;
        RECT 244.400 385.600 245.200 386.400 ;
        RECT 246.200 386.200 246.800 389.800 ;
        RECT 249.200 389.600 250.000 389.800 ;
        RECT 247.600 388.300 248.400 389.200 ;
        RECT 252.600 388.400 253.200 391.800 ;
        RECT 257.200 391.200 257.800 391.800 ;
        RECT 254.000 389.600 254.800 391.200 ;
        RECT 257.200 390.600 260.600 391.200 ;
        RECT 259.800 390.400 260.600 390.600 ;
        RECT 261.400 390.400 262.000 391.800 ;
        RECT 266.800 391.600 267.600 393.200 ;
        RECT 257.600 389.800 258.400 390.000 ;
        RECT 261.400 389.800 262.800 390.400 ;
        RECT 257.600 389.200 260.200 389.800 ;
        RECT 259.600 388.600 260.200 389.200 ;
        RECT 261.000 389.600 262.800 389.800 ;
        RECT 261.000 389.200 262.000 389.600 ;
        RECT 247.600 387.700 251.500 388.300 ;
        RECT 247.600 387.600 248.400 387.700 ;
        RECT 250.900 386.400 251.500 387.700 ;
        RECT 252.400 387.600 253.200 388.400 ;
        RECT 255.600 388.200 257.200 388.400 ;
        RECT 255.600 387.600 259.000 388.200 ;
        RECT 259.600 387.800 260.400 388.600 ;
        RECT 240.200 382.200 241.000 385.600 ;
        RECT 244.600 384.800 245.400 385.600 ;
        RECT 246.000 382.200 246.800 386.200 ;
        RECT 250.800 384.800 251.600 386.400 ;
        RECT 252.600 384.400 253.200 387.600 ;
        RECT 258.400 387.200 259.000 387.600 ;
        RECT 257.000 386.800 257.800 387.000 ;
        RECT 252.400 382.200 253.200 384.400 ;
        RECT 255.600 386.200 257.800 386.800 ;
        RECT 258.400 386.600 260.400 387.200 ;
        RECT 258.800 386.400 260.400 386.600 ;
        RECT 255.600 382.200 256.400 386.200 ;
        RECT 261.000 385.800 261.600 389.200 ;
        RECT 262.400 387.600 263.200 388.400 ;
        RECT 264.400 388.300 266.000 388.400 ;
        RECT 268.400 388.300 269.200 399.800 ;
        RECT 271.600 391.600 272.400 393.200 ;
        RECT 264.400 387.700 269.200 388.300 ;
        RECT 264.400 387.600 266.000 387.700 ;
        RECT 262.400 387.200 263.000 387.600 ;
        RECT 262.200 386.400 263.000 387.200 ;
        RECT 263.600 386.800 264.400 387.000 ;
        RECT 263.600 386.200 266.000 386.800 ;
        RECT 268.400 386.200 269.200 387.700 ;
        RECT 270.000 386.800 270.800 388.400 ;
        RECT 273.200 386.200 274.000 399.800 ;
        RECT 279.000 392.400 279.800 399.800 ;
        RECT 280.400 393.600 281.200 394.400 ;
        RECT 280.600 392.400 281.200 393.600 ;
        RECT 282.800 392.400 283.600 399.800 ;
        RECT 284.200 392.400 285.000 392.600 ;
        RECT 279.000 391.800 280.000 392.400 ;
        RECT 280.600 391.800 282.000 392.400 ;
        RECT 282.800 391.800 285.000 392.400 ;
        RECT 287.200 392.400 288.800 399.800 ;
        RECT 290.800 392.400 291.600 392.600 ;
        RECT 292.400 392.400 293.200 399.800 ;
        RECT 301.400 398.400 302.200 399.800 ;
        RECT 300.400 397.600 302.200 398.400 ;
        RECT 301.400 392.600 302.200 397.600 ;
        RECT 287.200 391.800 289.200 392.400 ;
        RECT 290.800 391.800 293.200 392.400 ;
        RECT 300.400 391.800 302.200 392.600 ;
        RECT 274.800 390.300 275.600 390.400 ;
        RECT 278.000 390.300 278.800 390.400 ;
        RECT 274.800 389.700 278.800 390.300 ;
        RECT 274.800 389.600 275.600 389.700 ;
        RECT 278.000 388.800 278.800 389.700 ;
        RECT 279.400 388.400 280.000 391.800 ;
        RECT 281.200 391.600 282.000 391.800 ;
        RECT 284.400 391.200 285.000 391.800 ;
        RECT 284.400 390.600 287.800 391.200 ;
        RECT 287.000 390.400 287.800 390.600 ;
        RECT 288.600 390.400 289.200 391.800 ;
        RECT 284.800 389.800 285.600 390.000 ;
        RECT 288.600 389.800 290.000 390.400 ;
        RECT 284.800 389.200 287.400 389.800 ;
        RECT 286.800 388.600 287.400 389.200 ;
        RECT 288.200 389.600 290.000 389.800 ;
        RECT 288.200 389.200 289.200 389.600 ;
        RECT 274.800 386.800 275.600 388.400 ;
        RECT 276.400 388.200 277.200 388.400 ;
        RECT 276.400 387.600 278.000 388.200 ;
        RECT 279.400 387.600 282.000 388.400 ;
        RECT 282.800 388.200 284.400 388.400 ;
        RECT 282.800 387.600 286.200 388.200 ;
        RECT 286.800 387.800 287.600 388.600 ;
        RECT 277.200 387.200 278.000 387.600 ;
        RECT 276.600 386.200 280.200 386.600 ;
        RECT 281.200 386.200 281.800 387.600 ;
        RECT 285.600 387.200 286.200 387.600 ;
        RECT 284.200 386.800 285.000 387.000 ;
        RECT 282.800 386.200 285.000 386.800 ;
        RECT 285.600 386.600 287.600 387.200 ;
        RECT 286.000 386.400 287.600 386.600 ;
        RECT 260.000 384.400 261.600 385.800 ;
        RECT 258.800 383.600 261.600 384.400 ;
        RECT 260.000 382.200 261.600 383.600 ;
        RECT 265.200 382.200 266.000 386.200 ;
        RECT 267.400 385.600 269.200 386.200 ;
        RECT 272.200 385.600 274.000 386.200 ;
        RECT 276.400 386.000 280.400 386.200 ;
        RECT 267.400 382.200 268.200 385.600 ;
        RECT 272.200 384.400 273.000 385.600 ;
        RECT 272.200 383.600 274.000 384.400 ;
        RECT 272.200 382.200 273.000 383.600 ;
        RECT 276.400 382.200 277.200 386.000 ;
        RECT 279.600 382.200 280.400 386.000 ;
        RECT 281.200 382.200 282.000 386.200 ;
        RECT 282.800 382.200 283.600 386.200 ;
        RECT 288.200 385.800 288.800 389.200 ;
        RECT 300.600 388.400 301.200 391.800 ;
        RECT 302.000 389.600 302.800 391.200 ;
        RECT 289.600 387.600 290.400 388.400 ;
        RECT 291.600 387.600 293.200 388.400 ;
        RECT 300.400 387.600 301.200 388.400 ;
        RECT 289.600 387.200 290.200 387.600 ;
        RECT 289.400 386.400 290.200 387.200 ;
        RECT 290.800 386.800 291.600 387.000 ;
        RECT 290.800 386.200 293.200 386.800 ;
        RECT 287.200 382.200 288.800 385.800 ;
        RECT 292.400 382.200 293.200 386.200 ;
        RECT 298.800 384.800 299.600 386.400 ;
        RECT 300.600 384.200 301.200 387.600 ;
        RECT 303.600 386.800 304.400 388.400 ;
        RECT 305.200 386.200 306.000 399.800 ;
        RECT 306.800 392.300 307.600 393.200 ;
        RECT 308.400 392.300 309.200 393.200 ;
        RECT 306.800 391.700 309.200 392.300 ;
        RECT 306.800 391.600 307.600 391.700 ;
        RECT 308.400 391.600 309.200 391.700 ;
        RECT 310.000 386.200 310.800 399.800 ;
        RECT 314.000 393.600 314.800 394.400 ;
        RECT 314.000 392.400 314.600 393.600 ;
        RECT 315.400 392.400 316.200 399.800 ;
        RECT 313.200 391.800 314.600 392.400 ;
        RECT 315.200 391.800 316.200 392.400 ;
        RECT 322.200 392.400 323.000 399.800 ;
        RECT 323.600 393.600 324.400 394.400 ;
        RECT 323.800 392.400 324.400 393.600 ;
        RECT 322.200 391.800 323.200 392.400 ;
        RECT 323.800 391.800 325.200 392.400 ;
        RECT 313.200 391.600 314.000 391.800 ;
        RECT 311.600 390.300 312.400 390.400 ;
        RECT 315.200 390.300 315.800 391.800 ;
        RECT 311.600 389.700 315.800 390.300 ;
        RECT 311.600 389.600 312.400 389.700 ;
        RECT 315.200 388.400 315.800 389.700 ;
        RECT 316.400 388.800 317.200 390.400 ;
        RECT 321.200 388.800 322.000 390.400 ;
        RECT 322.600 388.400 323.200 391.800 ;
        RECT 324.400 391.600 325.200 391.800 ;
        RECT 311.600 386.800 312.400 388.400 ;
        RECT 313.200 387.600 315.800 388.400 ;
        RECT 318.000 388.300 318.800 388.400 ;
        RECT 319.600 388.300 320.400 388.400 ;
        RECT 318.000 388.200 320.400 388.300 ;
        RECT 317.200 387.700 321.200 388.200 ;
        RECT 317.200 387.600 318.800 387.700 ;
        RECT 319.600 387.600 321.200 387.700 ;
        RECT 322.600 387.600 325.200 388.400 ;
        RECT 313.400 386.200 314.000 387.600 ;
        RECT 317.200 387.200 318.000 387.600 ;
        RECT 320.400 387.200 321.200 387.600 ;
        RECT 315.000 386.200 318.600 386.600 ;
        RECT 319.800 386.200 323.400 386.600 ;
        RECT 324.400 386.200 325.000 387.600 ;
        RECT 305.200 385.600 307.000 386.200 ;
        RECT 300.400 382.200 301.200 384.200 ;
        RECT 306.200 382.200 307.000 385.600 ;
        RECT 309.000 385.600 310.800 386.200 ;
        RECT 309.000 384.400 309.800 385.600 ;
        RECT 309.000 383.600 310.800 384.400 ;
        RECT 309.000 382.200 309.800 383.600 ;
        RECT 313.200 382.200 314.000 386.200 ;
        RECT 314.800 386.000 318.800 386.200 ;
        RECT 314.800 382.200 315.600 386.000 ;
        RECT 318.000 382.200 318.800 386.000 ;
        RECT 319.600 386.000 323.600 386.200 ;
        RECT 319.600 382.200 320.400 386.000 ;
        RECT 322.800 382.200 323.600 386.000 ;
        RECT 324.400 382.200 325.200 386.200 ;
        RECT 326.000 382.200 326.800 399.800 ;
        RECT 327.600 394.300 328.400 394.400 ;
        RECT 329.200 394.300 330.000 399.800 ;
        RECT 333.400 395.800 334.600 399.800 ;
        RECT 338.000 395.800 338.800 399.800 ;
        RECT 342.400 396.400 343.200 399.800 ;
        RECT 342.400 395.800 344.400 396.400 ;
        RECT 334.000 395.000 334.800 395.800 ;
        RECT 338.200 395.200 338.800 395.800 ;
        RECT 337.400 394.600 341.000 395.200 ;
        RECT 343.600 395.000 344.400 395.800 ;
        RECT 337.400 394.400 338.200 394.600 ;
        RECT 340.200 394.400 341.000 394.600 ;
        RECT 327.600 393.700 330.000 394.300 ;
        RECT 327.600 393.600 328.400 393.700 ;
        RECT 329.200 391.200 330.000 393.700 ;
        RECT 333.200 393.200 334.600 394.000 ;
        RECT 334.000 392.200 334.600 393.200 ;
        RECT 336.200 393.000 338.400 393.600 ;
        RECT 336.200 392.800 337.000 393.000 ;
        RECT 334.000 391.600 336.400 392.200 ;
        RECT 329.200 390.600 333.400 391.200 ;
        RECT 329.200 387.200 330.000 390.600 ;
        RECT 332.600 390.400 333.400 390.600 ;
        RECT 331.000 389.800 331.800 390.000 ;
        RECT 331.000 389.200 334.800 389.800 ;
        RECT 334.000 389.000 334.800 389.200 ;
        RECT 335.800 388.400 336.400 391.600 ;
        RECT 337.800 391.800 338.400 393.000 ;
        RECT 339.000 393.000 339.800 393.200 ;
        RECT 343.600 393.000 344.400 393.200 ;
        RECT 339.000 392.400 344.400 393.000 ;
        RECT 337.800 391.400 342.600 391.800 ;
        RECT 346.800 391.400 347.600 399.800 ;
        RECT 349.000 392.600 349.800 399.800 ;
        RECT 349.000 391.800 350.800 392.600 ;
        RECT 353.200 392.400 354.000 399.800 ;
        RECT 353.200 391.800 355.400 392.400 ;
        RECT 356.400 391.800 357.200 399.800 ;
        RECT 337.800 391.200 347.600 391.400 ;
        RECT 341.800 391.000 347.600 391.200 ;
        RECT 342.000 390.800 347.600 391.000 ;
        RECT 340.400 390.200 341.200 390.400 ;
        RECT 340.400 389.600 345.400 390.200 ;
        RECT 348.400 389.600 349.200 391.200 ;
        RECT 342.000 389.400 342.800 389.600 ;
        RECT 344.600 389.400 345.400 389.600 ;
        RECT 343.000 388.400 343.800 388.600 ;
        RECT 350.000 388.400 350.600 391.800 ;
        RECT 354.800 391.200 355.400 391.800 ;
        RECT 354.800 390.400 356.000 391.200 ;
        RECT 353.200 388.800 354.000 390.400 ;
        RECT 335.800 387.800 346.800 388.400 ;
        RECT 336.200 387.600 337.000 387.800 ;
        RECT 338.800 387.600 339.600 387.800 ;
        RECT 329.200 386.600 333.000 387.200 ;
        RECT 327.600 384.800 328.400 386.400 ;
        RECT 329.200 382.200 330.000 386.600 ;
        RECT 332.200 386.400 333.000 386.600 ;
        RECT 342.000 385.600 342.600 387.800 ;
        RECT 345.200 387.600 346.800 387.800 ;
        RECT 348.400 388.300 349.200 388.400 ;
        RECT 350.000 388.300 350.800 388.400 ;
        RECT 348.400 387.700 350.800 388.300 ;
        RECT 348.400 387.600 349.200 387.700 ;
        RECT 350.000 387.600 350.800 387.700 ;
        RECT 340.200 385.400 341.000 385.600 ;
        RECT 334.000 384.200 334.800 385.000 ;
        RECT 338.200 384.800 341.000 385.400 ;
        RECT 342.000 384.800 342.800 385.600 ;
        RECT 338.200 384.200 338.800 384.800 ;
        RECT 343.600 384.200 344.400 385.000 ;
        RECT 333.400 383.600 334.800 384.200 ;
        RECT 333.400 382.200 334.600 383.600 ;
        RECT 338.000 382.200 338.800 384.200 ;
        RECT 342.400 383.600 344.400 384.200 ;
        RECT 342.400 382.200 343.200 383.600 ;
        RECT 346.800 382.200 347.600 387.000 ;
        RECT 350.000 384.200 350.600 387.600 ;
        RECT 354.800 387.400 355.400 390.400 ;
        RECT 356.600 389.600 357.200 391.800 ;
        RECT 353.200 386.800 355.400 387.400 ;
        RECT 351.600 384.800 352.400 386.400 ;
        RECT 350.000 382.200 350.800 384.200 ;
        RECT 353.200 382.200 354.000 386.800 ;
        RECT 356.400 382.200 357.200 389.600 ;
        RECT 359.600 390.300 360.400 399.800 ;
        RECT 361.800 392.600 362.600 399.800 ;
        RECT 361.800 391.800 363.600 392.600 ;
        RECT 366.000 391.800 366.800 399.800 ;
        RECT 369.200 392.400 370.000 399.800 ;
        RECT 367.800 391.800 370.000 392.400 ;
        RECT 370.800 391.800 371.600 399.800 ;
        RECT 374.000 392.400 374.800 399.800 ;
        RECT 372.600 391.800 374.800 392.400 ;
        RECT 361.200 390.300 362.000 391.200 ;
        RECT 359.600 389.700 362.000 390.300 ;
        RECT 358.000 386.800 358.800 388.400 ;
        RECT 359.600 386.300 360.400 389.700 ;
        RECT 361.200 389.600 362.000 389.700 ;
        RECT 362.800 388.400 363.400 391.800 ;
        RECT 366.000 389.600 366.600 391.800 ;
        RECT 367.800 391.200 368.400 391.800 ;
        RECT 367.200 390.400 368.400 391.200 ;
        RECT 362.800 387.600 363.600 388.400 ;
        RECT 361.200 386.300 362.000 386.400 ;
        RECT 359.600 385.700 362.000 386.300 ;
        RECT 359.600 382.200 360.400 385.700 ;
        RECT 361.200 385.600 362.000 385.700 ;
        RECT 362.800 384.400 363.400 387.600 ;
        RECT 364.400 384.800 365.200 386.400 ;
        RECT 362.800 382.200 363.600 384.400 ;
        RECT 366.000 382.200 366.800 389.600 ;
        RECT 367.800 387.400 368.400 390.400 ;
        RECT 369.200 388.800 370.000 390.400 ;
        RECT 370.800 389.600 371.400 391.800 ;
        RECT 372.600 391.200 373.200 391.800 ;
        RECT 377.200 391.200 378.000 399.800 ;
        RECT 380.400 391.200 381.200 399.800 ;
        RECT 383.600 391.200 384.400 399.800 ;
        RECT 386.800 391.200 387.600 399.800 ;
        RECT 372.000 390.400 373.200 391.200 ;
        RECT 375.600 390.400 378.000 391.200 ;
        RECT 367.800 386.800 370.000 387.400 ;
        RECT 369.200 382.200 370.000 386.800 ;
        RECT 370.800 382.200 371.600 389.600 ;
        RECT 372.600 387.400 373.200 390.400 ;
        RECT 374.000 388.800 374.800 390.400 ;
        RECT 375.600 387.600 376.400 390.400 ;
        RECT 377.200 389.600 378.000 390.400 ;
        RECT 379.000 390.400 381.200 391.200 ;
        RECT 382.200 390.400 384.400 391.200 ;
        RECT 385.800 390.400 387.600 391.200 ;
        RECT 390.000 391.200 390.800 399.800 ;
        RECT 394.200 395.800 395.400 399.800 ;
        RECT 398.800 395.800 399.600 399.800 ;
        RECT 403.200 396.400 404.000 399.800 ;
        RECT 403.200 395.800 405.200 396.400 ;
        RECT 394.800 395.000 395.600 395.800 ;
        RECT 399.000 395.200 399.600 395.800 ;
        RECT 398.200 394.600 401.800 395.200 ;
        RECT 404.400 395.000 405.200 395.800 ;
        RECT 398.200 394.400 399.000 394.600 ;
        RECT 401.000 394.400 401.800 394.600 ;
        RECT 394.000 393.200 395.400 394.000 ;
        RECT 394.800 392.200 395.400 393.200 ;
        RECT 397.000 393.000 399.200 393.600 ;
        RECT 397.000 392.800 397.800 393.000 ;
        RECT 394.800 391.600 397.200 392.200 ;
        RECT 390.000 390.600 394.200 391.200 ;
        RECT 379.000 389.000 379.800 390.400 ;
        RECT 382.200 389.000 383.000 390.400 ;
        RECT 385.800 389.000 386.600 390.400 ;
        RECT 377.200 388.200 379.800 389.000 ;
        RECT 380.600 388.200 383.000 389.000 ;
        RECT 384.000 388.200 386.600 389.000 ;
        RECT 379.000 387.600 379.800 388.200 ;
        RECT 382.200 387.600 383.000 388.200 ;
        RECT 385.800 387.600 386.600 388.200 ;
        RECT 372.600 386.800 374.800 387.400 ;
        RECT 375.600 386.800 378.000 387.600 ;
        RECT 379.000 386.800 381.200 387.600 ;
        RECT 382.200 386.800 384.400 387.600 ;
        RECT 385.800 386.800 387.600 387.600 ;
        RECT 374.000 382.200 374.800 386.800 ;
        RECT 377.200 382.200 378.000 386.800 ;
        RECT 380.400 382.200 381.200 386.800 ;
        RECT 383.600 382.200 384.400 386.800 ;
        RECT 386.800 382.200 387.600 386.800 ;
        RECT 390.000 387.200 390.800 390.600 ;
        RECT 393.400 390.400 394.200 390.600 ;
        RECT 396.600 390.400 397.200 391.600 ;
        RECT 398.600 391.800 399.200 393.000 ;
        RECT 399.800 393.000 400.600 393.200 ;
        RECT 404.400 393.000 405.200 393.200 ;
        RECT 399.800 392.400 405.200 393.000 ;
        RECT 398.600 391.400 403.400 391.800 ;
        RECT 407.600 391.400 408.400 399.800 ;
        RECT 398.600 391.200 408.400 391.400 ;
        RECT 402.600 391.000 408.400 391.200 ;
        RECT 402.800 390.800 408.400 391.000 ;
        RECT 409.200 391.800 410.000 399.800 ;
        RECT 412.400 392.400 413.200 399.800 ;
        RECT 411.000 391.800 413.200 392.400 ;
        RECT 414.000 392.400 414.800 399.800 ;
        RECT 414.000 391.800 416.200 392.400 ;
        RECT 417.200 391.800 418.000 399.800 ;
        RECT 418.800 392.400 419.600 399.800 ;
        RECT 418.800 391.800 421.000 392.400 ;
        RECT 422.000 391.800 422.800 399.800 ;
        RECT 423.600 392.400 424.400 399.800 ;
        RECT 423.600 391.800 425.800 392.400 ;
        RECT 426.800 391.800 427.600 399.800 ;
        RECT 428.400 392.400 429.200 399.800 ;
        RECT 428.400 391.800 430.600 392.400 ;
        RECT 431.600 391.800 432.400 399.800 ;
        RECT 391.800 389.800 392.600 390.000 ;
        RECT 391.800 389.200 395.600 389.800 ;
        RECT 396.400 389.600 397.200 390.400 ;
        RECT 401.200 390.200 402.000 390.400 ;
        RECT 401.200 389.600 406.200 390.200 ;
        RECT 394.800 389.000 395.600 389.200 ;
        RECT 396.600 388.400 397.200 389.600 ;
        RECT 402.800 389.400 403.600 389.600 ;
        RECT 405.400 389.400 406.200 389.600 ;
        RECT 409.200 389.600 409.800 391.800 ;
        RECT 411.000 391.200 411.600 391.800 ;
        RECT 410.400 390.400 411.600 391.200 ;
        RECT 415.600 391.200 416.200 391.800 ;
        RECT 415.600 390.400 416.800 391.200 ;
        RECT 403.800 388.400 404.600 388.600 ;
        RECT 396.600 387.800 407.600 388.400 ;
        RECT 397.000 387.600 397.800 387.800 ;
        RECT 390.000 386.600 393.800 387.200 ;
        RECT 390.000 382.200 390.800 386.600 ;
        RECT 393.000 386.400 393.800 386.600 ;
        RECT 402.800 386.400 403.400 387.800 ;
        RECT 406.000 387.600 407.600 387.800 ;
        RECT 401.000 385.400 401.800 385.600 ;
        RECT 394.800 384.200 395.600 385.000 ;
        RECT 399.000 384.800 401.800 385.400 ;
        RECT 402.800 384.800 403.600 386.400 ;
        RECT 399.000 384.200 399.600 384.800 ;
        RECT 404.400 384.200 405.200 385.000 ;
        RECT 394.200 383.600 395.600 384.200 ;
        RECT 394.200 382.200 395.400 383.600 ;
        RECT 398.800 382.200 399.600 384.200 ;
        RECT 403.200 383.600 405.200 384.200 ;
        RECT 403.200 382.200 404.000 383.600 ;
        RECT 407.600 382.200 408.400 387.000 ;
        RECT 409.200 382.200 410.000 389.600 ;
        RECT 411.000 387.400 411.600 390.400 ;
        RECT 412.400 390.300 413.200 390.400 ;
        RECT 414.000 390.300 414.800 390.400 ;
        RECT 412.400 389.700 414.800 390.300 ;
        RECT 412.400 388.800 413.200 389.700 ;
        RECT 414.000 388.800 414.800 389.700 ;
        RECT 415.600 387.400 416.200 390.400 ;
        RECT 417.400 389.600 418.000 391.800 ;
        RECT 420.400 391.200 421.000 391.800 ;
        RECT 420.400 390.400 421.600 391.200 ;
        RECT 411.000 386.800 413.200 387.400 ;
        RECT 412.400 382.200 413.200 386.800 ;
        RECT 414.000 386.800 416.200 387.400 ;
        RECT 414.000 382.200 414.800 386.800 ;
        RECT 417.200 382.200 418.000 389.600 ;
        RECT 418.800 388.800 419.600 390.400 ;
        RECT 420.400 387.400 421.000 390.400 ;
        RECT 422.200 389.600 422.800 391.800 ;
        RECT 425.200 391.200 425.800 391.800 ;
        RECT 425.200 390.400 426.400 391.200 ;
        RECT 418.800 386.800 421.000 387.400 ;
        RECT 418.800 382.200 419.600 386.800 ;
        RECT 422.000 382.200 422.800 389.600 ;
        RECT 423.600 388.800 424.400 390.400 ;
        RECT 425.200 387.400 425.800 390.400 ;
        RECT 427.000 389.600 427.600 391.800 ;
        RECT 430.000 391.200 430.600 391.800 ;
        RECT 430.000 390.400 431.200 391.200 ;
        RECT 423.600 386.800 425.800 387.400 ;
        RECT 423.600 382.200 424.400 386.800 ;
        RECT 426.800 382.200 427.600 389.600 ;
        RECT 428.400 388.800 429.200 390.400 ;
        RECT 430.000 387.400 430.600 390.400 ;
        RECT 431.800 389.600 432.400 391.800 ;
        RECT 428.400 386.800 430.600 387.400 ;
        RECT 428.400 382.200 429.200 386.800 ;
        RECT 431.600 382.200 432.400 389.600 ;
        RECT 434.800 386.200 435.600 399.800 ;
        RECT 444.400 392.000 445.200 399.800 ;
        RECT 447.600 395.200 448.400 399.800 ;
        RECT 444.200 391.200 445.200 392.000 ;
        RECT 445.800 394.600 448.400 395.200 ;
        RECT 445.800 393.000 446.400 394.600 ;
        RECT 450.800 394.400 451.600 399.800 ;
        RECT 454.000 397.000 454.800 399.800 ;
        RECT 455.600 397.000 456.400 399.800 ;
        RECT 457.200 397.000 458.000 399.800 ;
        RECT 452.200 394.400 456.400 395.200 ;
        RECT 449.000 393.600 451.600 394.400 ;
        RECT 458.800 393.600 459.600 399.800 ;
        RECT 462.000 395.000 462.800 399.800 ;
        RECT 465.200 395.000 466.000 399.800 ;
        RECT 466.800 397.000 467.600 399.800 ;
        RECT 468.400 397.000 469.200 399.800 ;
        RECT 471.600 395.200 472.400 399.800 ;
        RECT 474.800 396.400 475.600 399.800 ;
        RECT 474.800 395.800 475.800 396.400 ;
        RECT 475.200 395.200 475.800 395.800 ;
        RECT 470.400 394.400 474.600 395.200 ;
        RECT 475.200 394.600 477.200 395.200 ;
        RECT 462.000 393.600 464.600 394.400 ;
        RECT 465.200 393.800 471.000 394.400 ;
        RECT 474.000 394.000 474.600 394.400 ;
        RECT 454.000 393.000 454.800 393.200 ;
        RECT 445.800 392.400 454.800 393.000 ;
        RECT 457.200 393.000 458.000 393.200 ;
        RECT 465.200 393.000 465.800 393.800 ;
        RECT 471.600 393.200 473.000 393.800 ;
        RECT 474.000 393.200 475.600 394.000 ;
        RECT 457.200 392.400 465.800 393.000 ;
        RECT 466.800 393.000 473.000 393.200 ;
        RECT 466.800 392.600 472.200 393.000 ;
        RECT 466.800 392.400 467.600 392.600 ;
        RECT 444.200 386.800 445.000 391.200 ;
        RECT 445.800 390.600 446.400 392.400 ;
        RECT 473.200 392.300 474.000 392.400 ;
        RECT 474.800 392.300 475.600 392.400 ;
        RECT 469.800 391.800 470.600 392.000 ;
        RECT 473.200 391.800 475.600 392.300 ;
        RECT 447.000 391.700 475.600 391.800 ;
        RECT 447.000 391.200 474.000 391.700 ;
        RECT 474.800 391.600 475.600 391.700 ;
        RECT 447.000 391.000 447.800 391.200 ;
        RECT 445.600 390.000 446.400 390.600 ;
        RECT 452.400 390.000 475.800 390.600 ;
        RECT 445.600 388.000 446.200 390.000 ;
        RECT 452.400 389.400 453.200 390.000 ;
        RECT 470.000 389.600 470.800 390.000 ;
        RECT 473.200 389.600 474.000 390.000 ;
        RECT 475.000 389.800 475.800 390.000 ;
        RECT 446.800 388.600 450.600 389.400 ;
        RECT 445.600 387.400 446.800 388.000 ;
        RECT 434.800 385.600 436.600 386.200 ;
        RECT 444.200 386.000 445.200 386.800 ;
        RECT 435.800 384.400 436.600 385.600 ;
        RECT 434.800 383.600 436.600 384.400 ;
        RECT 435.800 382.200 436.600 383.600 ;
        RECT 444.400 382.200 445.200 386.000 ;
        RECT 446.000 382.200 446.800 387.400 ;
        RECT 449.800 387.400 450.600 388.600 ;
        RECT 449.800 386.800 451.600 387.400 ;
        RECT 450.800 386.200 451.600 386.800 ;
        RECT 455.600 386.400 456.400 389.200 ;
        RECT 458.800 388.600 462.000 389.400 ;
        RECT 465.800 388.600 467.800 389.400 ;
        RECT 476.400 389.000 477.200 394.600 ;
        RECT 458.400 387.800 459.200 388.000 ;
        RECT 458.400 387.200 462.800 387.800 ;
        RECT 462.000 387.000 462.800 387.200 ;
        RECT 450.800 385.400 453.200 386.200 ;
        RECT 455.600 385.600 456.600 386.400 ;
        RECT 459.600 385.600 461.200 386.400 ;
        RECT 462.000 386.200 462.800 386.400 ;
        RECT 465.800 386.200 466.600 388.600 ;
        RECT 468.400 388.200 477.200 389.000 ;
        RECT 471.800 386.800 474.800 387.600 ;
        RECT 471.800 386.200 472.600 386.800 ;
        RECT 462.000 385.600 466.600 386.200 ;
        RECT 452.400 382.200 453.200 385.400 ;
        RECT 470.000 385.400 472.600 386.200 ;
        RECT 454.000 382.200 454.800 385.000 ;
        RECT 455.600 382.200 456.400 385.000 ;
        RECT 457.200 382.200 458.000 385.000 ;
        RECT 458.800 382.200 459.600 385.000 ;
        RECT 462.000 382.200 462.800 385.000 ;
        RECT 465.200 382.200 466.000 385.000 ;
        RECT 466.800 382.200 467.600 385.000 ;
        RECT 468.400 382.200 469.200 385.000 ;
        RECT 470.000 382.200 470.800 385.400 ;
        RECT 476.400 382.200 477.200 388.200 ;
        RECT 478.000 388.300 478.800 388.400 ;
        RECT 479.600 388.300 480.400 399.800 ;
        RECT 483.400 392.400 484.200 399.800 ;
        RECT 482.800 391.800 484.200 392.400 ;
        RECT 482.800 390.400 483.400 391.800 ;
        RECT 487.600 391.200 488.400 399.800 ;
        RECT 484.400 390.800 488.400 391.200 ;
        RECT 484.200 390.600 488.400 390.800 ;
        RECT 481.200 390.300 482.000 390.400 ;
        RECT 482.800 390.300 483.600 390.400 ;
        RECT 481.200 389.700 483.600 390.300 ;
        RECT 481.200 389.600 482.000 389.700 ;
        RECT 482.800 389.600 483.600 389.700 ;
        RECT 484.200 390.000 485.000 390.600 ;
        RECT 478.000 387.700 480.400 388.300 ;
        RECT 478.000 387.600 478.800 387.700 ;
        RECT 479.600 386.200 480.400 387.700 ;
        RECT 478.600 385.600 480.400 386.200 ;
        RECT 482.800 386.200 483.400 389.600 ;
        RECT 484.200 387.000 484.800 390.000 ;
        RECT 484.200 386.400 486.600 387.000 ;
        RECT 478.600 382.200 479.400 385.600 ;
        RECT 482.800 382.200 483.600 386.200 ;
        RECT 486.000 384.200 486.600 386.400 ;
        RECT 487.600 384.800 488.400 386.400 ;
        RECT 490.800 386.200 491.600 399.800 ;
        RECT 495.600 392.800 496.400 399.800 ;
        RECT 489.800 385.600 491.600 386.200 ;
        RECT 495.400 391.800 496.400 392.800 ;
        RECT 498.800 392.400 499.600 399.800 ;
        RECT 502.000 392.800 502.800 399.800 ;
        RECT 497.000 391.800 499.600 392.400 ;
        RECT 501.800 391.800 502.800 392.800 ;
        RECT 505.200 392.400 506.000 399.800 ;
        RECT 510.000 392.400 510.800 399.800 ;
        RECT 513.200 396.400 514.000 399.800 ;
        RECT 513.000 395.800 514.000 396.400 ;
        RECT 513.000 395.200 513.600 395.800 ;
        RECT 516.400 395.200 517.200 399.800 ;
        RECT 519.600 397.000 520.400 399.800 ;
        RECT 521.200 397.000 522.000 399.800 ;
        RECT 503.400 391.800 506.000 392.400 ;
        RECT 508.600 391.800 510.800 392.400 ;
        RECT 511.600 394.600 513.600 395.200 ;
        RECT 495.400 388.400 496.000 391.800 ;
        RECT 497.000 389.800 497.600 391.800 ;
        RECT 496.600 389.000 497.600 389.800 ;
        RECT 495.400 387.600 496.400 388.400 ;
        RECT 495.400 386.400 496.000 387.600 ;
        RECT 497.000 387.400 497.600 389.000 ;
        RECT 498.600 389.600 499.600 390.400 ;
        RECT 498.600 388.800 499.400 389.600 ;
        RECT 501.800 388.400 502.400 391.800 ;
        RECT 503.400 389.800 504.000 391.800 ;
        RECT 508.600 391.200 509.200 391.800 ;
        RECT 508.000 390.400 509.200 391.200 ;
        RECT 503.000 389.000 504.000 389.800 ;
        RECT 501.800 387.600 502.800 388.400 ;
        RECT 497.000 386.800 499.600 387.400 ;
        RECT 495.400 385.600 496.400 386.400 ;
        RECT 489.800 384.400 490.600 385.600 ;
        RECT 486.000 382.200 486.800 384.200 ;
        RECT 489.800 383.600 491.600 384.400 ;
        RECT 489.800 382.200 490.600 383.600 ;
        RECT 495.600 382.200 496.400 385.600 ;
        RECT 498.800 382.200 499.600 386.800 ;
        RECT 501.800 386.200 502.400 387.600 ;
        RECT 503.400 387.400 504.000 389.000 ;
        RECT 505.000 389.600 506.000 390.400 ;
        RECT 505.000 388.800 505.800 389.600 ;
        RECT 508.600 387.400 509.200 390.400 ;
        RECT 510.000 388.800 510.800 390.400 ;
        RECT 511.600 389.000 512.400 394.600 ;
        RECT 514.200 394.400 518.400 395.200 ;
        RECT 522.800 395.000 523.600 399.800 ;
        RECT 526.000 395.000 526.800 399.800 ;
        RECT 514.200 394.000 514.800 394.400 ;
        RECT 513.200 393.200 514.800 394.000 ;
        RECT 517.800 393.800 523.600 394.400 ;
        RECT 515.800 393.200 517.200 393.800 ;
        RECT 515.800 393.000 522.000 393.200 ;
        RECT 516.600 392.600 522.000 393.000 ;
        RECT 521.200 392.400 522.000 392.600 ;
        RECT 523.000 393.000 523.600 393.800 ;
        RECT 524.200 393.600 526.800 394.400 ;
        RECT 529.200 393.600 530.000 399.800 ;
        RECT 530.800 397.000 531.600 399.800 ;
        RECT 532.400 397.000 533.200 399.800 ;
        RECT 534.000 397.000 534.800 399.800 ;
        RECT 532.400 394.400 536.600 395.200 ;
        RECT 537.200 394.400 538.000 399.800 ;
        RECT 540.400 395.200 541.200 399.800 ;
        RECT 540.400 394.600 543.000 395.200 ;
        RECT 537.200 393.600 539.800 394.400 ;
        RECT 530.800 393.000 531.600 393.200 ;
        RECT 523.000 392.400 531.600 393.000 ;
        RECT 534.000 393.000 534.800 393.200 ;
        RECT 542.400 393.000 543.000 394.600 ;
        RECT 534.000 392.400 543.000 393.000 ;
        RECT 542.400 390.600 543.000 392.400 ;
        RECT 543.600 392.000 544.400 399.800 ;
        RECT 548.400 396.400 549.200 399.800 ;
        RECT 548.200 395.800 549.200 396.400 ;
        RECT 548.200 395.200 548.800 395.800 ;
        RECT 551.600 395.200 552.400 399.800 ;
        RECT 554.800 397.000 555.600 399.800 ;
        RECT 556.400 397.000 557.200 399.800 ;
        RECT 546.800 394.600 548.800 395.200 ;
        RECT 543.600 391.200 544.600 392.000 ;
        RECT 513.000 390.000 536.400 390.600 ;
        RECT 542.400 390.000 543.200 390.600 ;
        RECT 513.000 389.800 513.800 390.000 ;
        RECT 514.800 389.600 515.600 390.000 ;
        RECT 518.000 389.600 518.800 390.000 ;
        RECT 535.600 389.400 536.400 390.000 ;
        RECT 511.600 388.200 520.400 389.000 ;
        RECT 521.000 388.600 523.000 389.400 ;
        RECT 526.800 388.600 530.000 389.400 ;
        RECT 503.400 386.800 506.000 387.400 ;
        RECT 508.600 386.800 510.800 387.400 ;
        RECT 501.800 385.600 502.800 386.200 ;
        RECT 502.000 382.200 502.800 385.600 ;
        RECT 505.200 382.200 506.000 386.800 ;
        RECT 510.000 382.200 510.800 386.800 ;
        RECT 511.600 382.200 512.400 388.200 ;
        RECT 514.000 386.800 517.000 387.600 ;
        RECT 516.200 386.200 517.000 386.800 ;
        RECT 522.200 386.200 523.000 388.600 ;
        RECT 524.400 386.800 525.200 388.400 ;
        RECT 529.600 387.800 530.400 388.000 ;
        RECT 526.000 387.200 530.400 387.800 ;
        RECT 526.000 387.000 526.800 387.200 ;
        RECT 532.400 386.400 533.200 389.200 ;
        RECT 538.200 388.600 542.000 389.400 ;
        RECT 538.200 387.400 539.000 388.600 ;
        RECT 542.600 388.000 543.200 390.000 ;
        RECT 526.000 386.200 526.800 386.400 ;
        RECT 516.200 385.400 518.800 386.200 ;
        RECT 522.200 385.600 526.800 386.200 ;
        RECT 527.600 385.600 529.200 386.400 ;
        RECT 532.200 385.600 533.200 386.400 ;
        RECT 537.200 386.800 539.000 387.400 ;
        RECT 542.000 387.400 543.200 388.000 ;
        RECT 537.200 386.200 538.000 386.800 ;
        RECT 518.000 382.200 518.800 385.400 ;
        RECT 535.600 385.400 538.000 386.200 ;
        RECT 519.600 382.200 520.400 385.000 ;
        RECT 521.200 382.200 522.000 385.000 ;
        RECT 522.800 382.200 523.600 385.000 ;
        RECT 526.000 382.200 526.800 385.000 ;
        RECT 529.200 382.200 530.000 385.000 ;
        RECT 530.800 382.200 531.600 385.000 ;
        RECT 532.400 382.200 533.200 385.000 ;
        RECT 534.000 382.200 534.800 385.000 ;
        RECT 535.600 382.200 536.400 385.400 ;
        RECT 542.000 382.200 542.800 387.400 ;
        RECT 543.800 386.800 544.600 391.200 ;
        RECT 543.600 386.000 544.600 386.800 ;
        RECT 546.800 389.000 547.600 394.600 ;
        RECT 549.400 394.400 553.600 395.200 ;
        RECT 558.000 395.000 558.800 399.800 ;
        RECT 561.200 395.000 562.000 399.800 ;
        RECT 549.400 394.000 550.000 394.400 ;
        RECT 548.400 393.200 550.000 394.000 ;
        RECT 553.000 393.800 558.800 394.400 ;
        RECT 551.000 393.200 552.400 393.800 ;
        RECT 551.000 393.000 557.200 393.200 ;
        RECT 551.800 392.600 557.200 393.000 ;
        RECT 556.400 392.400 557.200 392.600 ;
        RECT 558.200 393.000 558.800 393.800 ;
        RECT 559.400 393.600 562.000 394.400 ;
        RECT 564.400 393.600 565.200 399.800 ;
        RECT 566.000 397.000 566.800 399.800 ;
        RECT 567.600 397.000 568.400 399.800 ;
        RECT 569.200 397.000 570.000 399.800 ;
        RECT 567.600 394.400 571.800 395.200 ;
        RECT 572.400 394.400 573.200 399.800 ;
        RECT 575.600 395.200 576.400 399.800 ;
        RECT 575.600 394.600 578.200 395.200 ;
        RECT 572.400 393.600 575.000 394.400 ;
        RECT 566.000 393.000 566.800 393.200 ;
        RECT 558.200 392.400 566.800 393.000 ;
        RECT 569.200 393.000 570.000 393.200 ;
        RECT 577.600 393.000 578.200 394.600 ;
        RECT 569.200 392.400 578.200 393.000 ;
        RECT 577.600 390.600 578.200 392.400 ;
        RECT 578.800 392.000 579.600 399.800 ;
        RECT 578.800 391.200 579.800 392.000 ;
        RECT 548.200 390.000 571.600 390.600 ;
        RECT 577.600 390.000 578.400 390.600 ;
        RECT 548.200 389.800 549.000 390.000 ;
        RECT 551.600 389.600 552.400 390.000 ;
        RECT 553.200 389.600 554.000 390.000 ;
        RECT 570.800 389.400 571.600 390.000 ;
        RECT 546.800 388.200 555.600 389.000 ;
        RECT 556.200 388.600 558.200 389.400 ;
        RECT 562.000 388.600 565.200 389.400 ;
        RECT 543.600 382.200 544.400 386.000 ;
        RECT 546.800 382.200 547.600 388.200 ;
        RECT 549.200 386.800 552.200 387.600 ;
        RECT 551.400 386.200 552.200 386.800 ;
        RECT 557.400 386.200 558.200 388.600 ;
        RECT 559.600 386.800 560.400 388.400 ;
        RECT 564.800 387.800 565.600 388.000 ;
        RECT 561.200 387.200 565.600 387.800 ;
        RECT 561.200 387.000 562.000 387.200 ;
        RECT 567.600 386.400 568.400 389.200 ;
        RECT 573.400 388.600 577.200 389.400 ;
        RECT 573.400 387.400 574.200 388.600 ;
        RECT 577.800 388.000 578.400 390.000 ;
        RECT 561.200 386.200 562.000 386.400 ;
        RECT 551.400 385.400 554.000 386.200 ;
        RECT 557.400 385.600 562.000 386.200 ;
        RECT 562.800 385.600 564.400 386.400 ;
        RECT 567.400 385.600 568.400 386.400 ;
        RECT 572.400 386.800 574.200 387.400 ;
        RECT 577.200 387.400 578.400 388.000 ;
        RECT 572.400 386.200 573.200 386.800 ;
        RECT 553.200 382.200 554.000 385.400 ;
        RECT 570.800 385.400 573.200 386.200 ;
        RECT 554.800 382.200 555.600 385.000 ;
        RECT 556.400 382.200 557.200 385.000 ;
        RECT 558.000 382.200 558.800 385.000 ;
        RECT 561.200 382.200 562.000 385.000 ;
        RECT 564.400 382.200 565.200 385.000 ;
        RECT 566.000 382.200 566.800 385.000 ;
        RECT 567.600 382.200 568.400 385.000 ;
        RECT 569.200 382.200 570.000 385.000 ;
        RECT 570.800 382.200 571.600 385.400 ;
        RECT 577.200 382.200 578.000 387.400 ;
        RECT 579.000 386.800 579.800 391.200 ;
        RECT 578.800 386.000 579.800 386.800 ;
        RECT 578.800 382.200 579.600 386.000 ;
        RECT 3.800 376.400 4.600 379.800 ;
        RECT 2.800 375.800 4.600 376.400 ;
        RECT 6.000 375.800 6.800 379.800 ;
        RECT 7.600 376.000 8.400 379.800 ;
        RECT 10.800 376.000 11.600 379.800 ;
        RECT 7.600 375.800 11.600 376.000 ;
        RECT 14.000 377.800 14.800 379.800 ;
        RECT 1.200 373.600 2.000 375.200 ;
        RECT 1.200 368.300 2.000 368.400 ;
        RECT 2.800 368.300 3.600 375.800 ;
        RECT 6.200 374.400 6.800 375.800 ;
        RECT 7.800 375.400 11.400 375.800 ;
        RECT 10.000 374.400 10.800 374.800 ;
        RECT 14.000 374.400 14.600 377.800 ;
        RECT 15.600 375.600 16.400 377.200 ;
        RECT 6.000 373.600 8.600 374.400 ;
        RECT 10.000 373.800 11.600 374.400 ;
        RECT 10.800 373.600 11.600 373.800 ;
        RECT 14.000 373.600 14.800 374.400 ;
        RECT 8.000 372.300 8.600 373.600 ;
        RECT 4.500 371.700 8.600 372.300 ;
        RECT 4.500 370.400 5.100 371.700 ;
        RECT 4.400 368.800 5.200 370.400 ;
        RECT 6.000 370.200 6.800 370.400 ;
        RECT 8.000 370.200 8.600 371.700 ;
        RECT 9.200 371.600 10.000 373.200 ;
        RECT 10.900 372.300 11.500 373.600 ;
        RECT 12.400 372.300 13.200 372.400 ;
        RECT 10.900 371.700 13.200 372.300 ;
        RECT 12.400 370.800 13.200 371.700 ;
        RECT 14.000 370.200 14.600 373.600 ;
        RECT 6.000 369.600 7.400 370.200 ;
        RECT 8.000 369.600 9.000 370.200 ;
        RECT 1.200 367.700 3.600 368.300 ;
        RECT 1.200 367.600 2.000 367.700 ;
        RECT 2.800 362.200 3.600 367.700 ;
        RECT 6.800 368.400 7.400 369.600 ;
        RECT 6.800 367.600 7.600 368.400 ;
        RECT 8.200 362.200 9.000 369.600 ;
        RECT 13.000 369.400 14.800 370.200 ;
        RECT 13.000 368.400 13.800 369.400 ;
        RECT 13.000 367.600 14.800 368.400 ;
        RECT 13.000 362.200 13.800 367.600 ;
        RECT 17.200 362.200 18.000 379.800 ;
        RECT 18.800 375.600 19.600 377.200 ;
        RECT 20.400 375.800 21.200 379.800 ;
        RECT 22.000 376.000 22.800 379.800 ;
        RECT 25.200 376.000 26.000 379.800 ;
        RECT 22.000 375.800 26.000 376.000 ;
        RECT 27.400 376.400 28.200 379.800 ;
        RECT 33.200 377.600 34.000 379.800 ;
        RECT 27.400 375.800 29.200 376.400 ;
        RECT 20.600 374.400 21.200 375.800 ;
        RECT 22.200 375.400 25.800 375.800 ;
        RECT 24.400 374.400 25.200 374.800 ;
        RECT 20.400 373.600 23.000 374.400 ;
        RECT 24.400 373.800 26.000 374.400 ;
        RECT 25.200 373.600 26.000 373.800 ;
        RECT 22.400 372.400 23.000 373.600 ;
        RECT 22.000 371.600 23.000 372.400 ;
        RECT 23.600 372.300 24.400 373.200 ;
        RECT 25.200 372.300 26.000 372.400 ;
        RECT 23.600 371.700 26.000 372.300 ;
        RECT 23.600 371.600 24.400 371.700 ;
        RECT 25.200 371.600 26.000 371.700 ;
        RECT 20.400 370.200 21.200 370.400 ;
        RECT 22.400 370.200 23.000 371.600 ;
        RECT 20.400 369.600 21.800 370.200 ;
        RECT 22.400 369.600 23.400 370.200 ;
        RECT 21.200 368.400 21.800 369.600 ;
        RECT 21.200 367.600 22.000 368.400 ;
        RECT 22.600 362.200 23.400 369.600 ;
        RECT 26.800 368.800 27.600 370.400 ;
        RECT 28.400 362.200 29.200 375.800 ;
        RECT 31.600 375.600 32.400 377.200 ;
        RECT 30.000 373.600 30.800 375.200 ;
        RECT 33.400 374.400 34.000 377.600 ;
        RECT 36.400 376.000 37.200 379.800 ;
        RECT 39.600 376.000 40.400 379.800 ;
        RECT 36.400 375.800 40.400 376.000 ;
        RECT 41.200 375.800 42.000 379.800 ;
        RECT 42.800 375.800 43.600 379.800 ;
        RECT 44.400 376.000 45.200 379.800 ;
        RECT 47.600 376.000 48.400 379.800 ;
        RECT 44.400 375.800 48.400 376.000 ;
        RECT 36.600 375.400 40.200 375.800 ;
        RECT 37.200 374.400 38.000 374.800 ;
        RECT 41.200 374.400 41.800 375.800 ;
        RECT 43.000 374.400 43.600 375.800 ;
        RECT 44.600 375.400 48.200 375.800 ;
        RECT 49.200 375.400 50.000 379.800 ;
        RECT 53.400 378.400 54.600 379.800 ;
        RECT 53.400 377.800 54.800 378.400 ;
        RECT 58.000 377.800 58.800 379.800 ;
        RECT 62.400 378.400 63.200 379.800 ;
        RECT 62.400 377.800 64.400 378.400 ;
        RECT 54.000 377.000 54.800 377.800 ;
        RECT 58.200 377.200 58.800 377.800 ;
        RECT 58.200 376.600 61.000 377.200 ;
        RECT 60.200 376.400 61.000 376.600 ;
        RECT 62.000 376.400 62.800 377.200 ;
        RECT 63.600 377.000 64.400 377.800 ;
        RECT 52.200 375.400 53.000 375.600 ;
        RECT 49.200 374.800 53.000 375.400 ;
        RECT 46.800 374.400 47.600 374.800 ;
        RECT 33.200 373.600 34.000 374.400 ;
        RECT 36.400 373.800 38.000 374.400 ;
        RECT 36.400 373.600 37.200 373.800 ;
        RECT 39.400 373.600 42.000 374.400 ;
        RECT 42.800 373.600 45.400 374.400 ;
        RECT 46.800 373.800 48.400 374.400 ;
        RECT 47.600 373.600 48.400 373.800 ;
        RECT 33.400 370.200 34.000 373.600 ;
        RECT 34.800 370.800 35.600 372.400 ;
        RECT 38.000 371.600 38.800 373.200 ;
        RECT 39.400 370.200 40.000 373.600 ;
        RECT 44.800 372.300 45.400 373.600 ;
        RECT 41.300 371.700 45.400 372.300 ;
        RECT 41.300 370.400 41.900 371.700 ;
        RECT 41.200 370.200 42.000 370.400 ;
        RECT 33.200 369.400 35.000 370.200 ;
        RECT 34.200 362.200 35.000 369.400 ;
        RECT 39.000 369.600 40.000 370.200 ;
        RECT 40.600 369.600 42.000 370.200 ;
        RECT 42.800 370.200 43.600 370.400 ;
        RECT 44.800 370.200 45.400 371.700 ;
        RECT 46.000 371.600 46.800 373.200 ;
        RECT 49.200 371.400 50.000 374.800 ;
        RECT 56.200 374.200 57.000 374.400 ;
        RECT 62.000 374.200 62.600 376.400 ;
        RECT 66.800 375.000 67.600 379.800 ;
        RECT 69.000 376.800 69.800 379.800 ;
        RECT 68.400 375.800 69.800 376.800 ;
        RECT 73.200 375.800 74.000 379.800 ;
        RECT 65.200 374.200 66.800 374.400 ;
        RECT 55.800 373.600 66.800 374.200 ;
        RECT 54.000 372.800 54.800 373.000 ;
        RECT 51.000 372.200 54.800 372.800 ;
        RECT 51.000 372.000 51.800 372.200 ;
        RECT 52.600 371.400 53.400 371.600 ;
        RECT 49.200 370.800 53.400 371.400 ;
        RECT 42.800 369.600 44.200 370.200 ;
        RECT 44.800 369.600 45.800 370.200 ;
        RECT 39.000 362.200 39.800 369.600 ;
        RECT 40.600 368.400 41.200 369.600 ;
        RECT 40.400 367.600 41.200 368.400 ;
        RECT 43.600 368.400 44.200 369.600 ;
        RECT 43.600 367.600 44.400 368.400 ;
        RECT 45.000 362.200 45.800 369.600 ;
        RECT 49.200 362.200 50.000 370.800 ;
        RECT 55.800 370.400 56.400 373.600 ;
        RECT 63.000 373.400 63.800 373.600 ;
        RECT 62.000 372.400 62.800 372.600 ;
        RECT 64.600 372.400 65.400 372.600 ;
        RECT 60.400 371.800 65.400 372.400 ;
        RECT 68.400 372.400 69.000 375.800 ;
        RECT 73.200 375.600 73.800 375.800 ;
        RECT 72.000 375.200 73.800 375.600 ;
        RECT 69.600 375.000 73.800 375.200 ;
        RECT 69.600 374.600 72.600 375.000 ;
        RECT 69.600 374.400 70.400 374.600 ;
        RECT 60.400 371.600 61.200 371.800 ;
        RECT 68.400 371.600 69.200 372.400 ;
        RECT 62.000 371.000 67.600 371.200 ;
        RECT 61.800 370.800 67.600 371.000 ;
        RECT 54.000 369.800 56.400 370.400 ;
        RECT 57.800 370.600 67.600 370.800 ;
        RECT 57.800 370.200 62.600 370.600 ;
        RECT 54.000 368.800 54.600 369.800 ;
        RECT 53.200 368.000 54.600 368.800 ;
        RECT 56.200 369.000 57.000 369.200 ;
        RECT 57.800 369.000 58.400 370.200 ;
        RECT 56.200 368.400 58.400 369.000 ;
        RECT 59.000 369.000 64.400 369.600 ;
        RECT 59.000 368.800 59.800 369.000 ;
        RECT 63.600 368.800 64.400 369.000 ;
        RECT 57.400 367.400 58.200 367.600 ;
        RECT 60.200 367.400 61.000 367.600 ;
        RECT 54.000 366.200 54.800 367.000 ;
        RECT 57.400 366.800 61.000 367.400 ;
        RECT 58.200 366.200 58.800 366.800 ;
        RECT 63.600 366.200 64.400 367.000 ;
        RECT 53.400 362.200 54.600 366.200 ;
        RECT 58.000 362.200 58.800 366.200 ;
        RECT 62.400 365.600 64.400 366.200 ;
        RECT 62.400 362.200 63.200 365.600 ;
        RECT 66.800 362.200 67.600 370.600 ;
        RECT 68.400 370.400 69.000 371.600 ;
        RECT 69.800 371.000 70.400 374.400 ;
        RECT 71.200 373.800 72.000 374.000 ;
        RECT 71.200 373.200 72.200 373.800 ;
        RECT 71.600 372.400 72.200 373.200 ;
        RECT 73.200 372.800 74.000 374.400 ;
        RECT 71.600 371.600 72.400 372.400 ;
        RECT 69.800 370.400 72.200 371.000 ;
        RECT 68.400 362.200 69.200 370.400 ;
        RECT 71.600 366.200 72.200 370.400 ;
        RECT 71.600 362.200 72.400 366.200 ;
        RECT 74.800 362.200 75.600 379.800 ;
        RECT 78.000 375.400 78.800 379.800 ;
        RECT 82.200 378.400 83.400 379.800 ;
        RECT 82.200 377.800 83.600 378.400 ;
        RECT 86.800 377.800 87.600 379.800 ;
        RECT 91.200 378.400 92.000 379.800 ;
        RECT 91.200 377.800 93.200 378.400 ;
        RECT 82.800 377.000 83.600 377.800 ;
        RECT 87.000 377.200 87.600 377.800 ;
        RECT 87.000 376.600 89.800 377.200 ;
        RECT 89.000 376.400 89.800 376.600 ;
        RECT 90.800 376.400 91.600 377.200 ;
        RECT 92.400 377.000 93.200 377.800 ;
        RECT 81.000 375.400 81.800 375.600 ;
        RECT 76.400 373.600 77.200 375.200 ;
        RECT 78.000 374.800 81.800 375.400 ;
        RECT 78.000 371.400 78.800 374.800 ;
        RECT 85.000 374.200 85.800 374.400 ;
        RECT 90.800 374.200 91.400 376.400 ;
        RECT 95.600 375.000 96.400 379.800 ;
        RECT 97.200 375.400 98.000 379.800 ;
        RECT 101.400 378.400 102.600 379.800 ;
        RECT 101.400 377.800 102.800 378.400 ;
        RECT 106.000 377.800 106.800 379.800 ;
        RECT 110.400 378.400 111.200 379.800 ;
        RECT 110.400 377.800 112.400 378.400 ;
        RECT 102.000 377.000 102.800 377.800 ;
        RECT 106.200 377.200 106.800 377.800 ;
        RECT 106.200 376.600 109.000 377.200 ;
        RECT 108.200 376.400 109.000 376.600 ;
        RECT 110.000 375.600 110.800 377.200 ;
        RECT 111.600 377.000 112.400 377.800 ;
        RECT 100.200 375.400 101.000 375.600 ;
        RECT 97.200 374.800 101.000 375.400 ;
        RECT 94.000 374.200 95.600 374.400 ;
        RECT 84.600 373.600 95.600 374.200 ;
        RECT 82.800 372.800 83.600 373.000 ;
        RECT 79.800 372.200 83.600 372.800 ;
        RECT 84.600 372.400 85.200 373.600 ;
        RECT 91.800 373.400 92.600 373.600 ;
        RECT 90.800 372.400 91.600 372.600 ;
        RECT 93.400 372.400 94.200 372.600 ;
        RECT 79.800 372.000 80.600 372.200 ;
        RECT 84.400 371.600 85.200 372.400 ;
        RECT 89.200 371.800 94.200 372.400 ;
        RECT 89.200 371.600 90.000 371.800 ;
        RECT 81.400 371.400 82.200 371.600 ;
        RECT 78.000 370.800 82.200 371.400 ;
        RECT 78.000 362.200 78.800 370.800 ;
        RECT 84.600 370.400 85.200 371.600 ;
        RECT 97.200 371.400 98.000 374.800 ;
        RECT 104.200 374.200 105.000 374.400 ;
        RECT 110.000 374.200 110.600 375.600 ;
        RECT 114.800 375.000 115.600 379.800 ;
        RECT 116.400 375.400 117.200 379.800 ;
        RECT 120.600 378.400 121.800 379.800 ;
        RECT 120.600 377.800 122.000 378.400 ;
        RECT 125.200 377.800 126.000 379.800 ;
        RECT 129.600 378.400 130.400 379.800 ;
        RECT 129.600 377.800 131.600 378.400 ;
        RECT 121.200 377.000 122.000 377.800 ;
        RECT 125.400 377.200 126.000 377.800 ;
        RECT 125.400 376.600 128.200 377.200 ;
        RECT 127.400 376.400 128.200 376.600 ;
        RECT 129.200 375.600 130.000 377.200 ;
        RECT 130.800 377.000 131.600 377.800 ;
        RECT 119.400 375.400 120.200 375.600 ;
        RECT 116.400 374.800 120.200 375.400 ;
        RECT 113.200 374.200 114.800 374.400 ;
        RECT 103.800 373.600 114.800 374.200 ;
        RECT 102.000 372.800 102.800 373.000 ;
        RECT 99.000 372.200 102.800 372.800 ;
        RECT 99.000 372.000 99.800 372.200 ;
        RECT 100.600 371.400 101.400 371.600 ;
        RECT 90.800 371.000 96.400 371.200 ;
        RECT 90.600 370.800 96.400 371.000 ;
        RECT 82.800 369.800 85.200 370.400 ;
        RECT 86.600 370.600 96.400 370.800 ;
        RECT 86.600 370.200 91.400 370.600 ;
        RECT 82.800 368.800 83.400 369.800 ;
        RECT 82.000 368.000 83.400 368.800 ;
        RECT 85.000 369.000 85.800 369.200 ;
        RECT 86.600 369.000 87.200 370.200 ;
        RECT 85.000 368.400 87.200 369.000 ;
        RECT 87.800 369.000 93.200 369.600 ;
        RECT 87.800 368.800 88.600 369.000 ;
        RECT 92.400 368.800 93.200 369.000 ;
        RECT 86.200 367.400 87.000 367.600 ;
        RECT 89.000 367.400 89.800 367.600 ;
        RECT 82.800 366.200 83.600 367.000 ;
        RECT 86.200 366.800 89.800 367.400 ;
        RECT 87.000 366.200 87.600 366.800 ;
        RECT 92.400 366.200 93.200 367.000 ;
        RECT 82.200 362.200 83.400 366.200 ;
        RECT 86.800 362.200 87.600 366.200 ;
        RECT 91.200 365.600 93.200 366.200 ;
        RECT 91.200 362.200 92.000 365.600 ;
        RECT 95.600 362.200 96.400 370.600 ;
        RECT 97.200 370.800 101.400 371.400 ;
        RECT 97.200 362.200 98.000 370.800 ;
        RECT 103.800 370.400 104.400 373.600 ;
        RECT 111.000 373.400 111.800 373.600 ;
        RECT 110.000 372.400 110.800 372.600 ;
        RECT 112.600 372.400 113.400 372.600 ;
        RECT 108.400 371.800 113.400 372.400 ;
        RECT 108.400 371.600 109.200 371.800 ;
        RECT 116.400 371.400 117.200 374.800 ;
        RECT 123.400 374.200 124.200 374.400 ;
        RECT 129.200 374.200 129.800 375.600 ;
        RECT 134.000 375.000 134.800 379.800 ;
        RECT 140.400 375.400 141.200 379.800 ;
        RECT 144.600 378.400 145.800 379.800 ;
        RECT 144.600 377.800 146.000 378.400 ;
        RECT 149.200 377.800 150.000 379.800 ;
        RECT 153.600 378.400 154.400 379.800 ;
        RECT 153.600 377.800 155.600 378.400 ;
        RECT 145.200 377.000 146.000 377.800 ;
        RECT 149.400 377.200 150.000 377.800 ;
        RECT 149.400 376.600 152.200 377.200 ;
        RECT 151.400 376.400 152.200 376.600 ;
        RECT 153.200 376.400 154.000 377.200 ;
        RECT 154.800 377.000 155.600 377.800 ;
        RECT 143.400 375.400 144.200 375.600 ;
        RECT 140.400 374.800 144.200 375.400 ;
        RECT 132.400 374.200 134.000 374.400 ;
        RECT 123.000 373.600 134.000 374.200 ;
        RECT 121.200 372.800 122.000 373.000 ;
        RECT 118.200 372.200 122.000 372.800 ;
        RECT 118.200 372.000 119.000 372.200 ;
        RECT 119.800 371.400 120.600 371.600 ;
        RECT 110.000 371.000 115.600 371.200 ;
        RECT 109.800 370.800 115.600 371.000 ;
        RECT 102.000 369.800 104.400 370.400 ;
        RECT 105.800 370.600 115.600 370.800 ;
        RECT 105.800 370.200 110.600 370.600 ;
        RECT 102.000 368.800 102.600 369.800 ;
        RECT 101.200 368.400 102.600 368.800 ;
        RECT 104.200 369.000 105.000 369.200 ;
        RECT 105.800 369.000 106.400 370.200 ;
        RECT 104.200 368.400 106.400 369.000 ;
        RECT 107.000 369.000 112.400 369.600 ;
        RECT 107.000 368.800 107.800 369.000 ;
        RECT 111.600 368.800 112.400 369.000 ;
        RECT 100.400 368.000 102.600 368.400 ;
        RECT 100.400 367.600 101.800 368.000 ;
        RECT 105.400 367.400 106.200 367.600 ;
        RECT 108.200 367.400 109.000 367.600 ;
        RECT 102.000 366.200 102.800 367.000 ;
        RECT 105.400 366.800 109.000 367.400 ;
        RECT 106.200 366.200 106.800 366.800 ;
        RECT 111.600 366.200 112.400 367.000 ;
        RECT 101.400 362.200 102.600 366.200 ;
        RECT 106.000 362.200 106.800 366.200 ;
        RECT 110.400 365.600 112.400 366.200 ;
        RECT 110.400 362.200 111.200 365.600 ;
        RECT 114.800 362.200 115.600 370.600 ;
        RECT 116.400 370.800 120.600 371.400 ;
        RECT 116.400 362.200 117.200 370.800 ;
        RECT 123.000 370.400 123.600 373.600 ;
        RECT 130.200 373.400 131.000 373.600 ;
        RECT 131.800 372.400 132.600 372.600 ;
        RECT 127.600 371.800 132.600 372.400 ;
        RECT 127.600 371.600 128.400 371.800 ;
        RECT 140.400 371.400 141.200 374.800 ;
        RECT 147.400 374.200 148.200 374.400 ;
        RECT 150.000 374.200 150.800 374.400 ;
        RECT 153.200 374.200 153.800 376.400 ;
        RECT 158.000 375.000 158.800 379.800 ;
        RECT 159.600 375.800 160.400 379.800 ;
        RECT 164.000 376.200 165.600 379.800 ;
        RECT 159.600 375.200 162.000 375.800 ;
        RECT 161.200 375.000 162.000 375.200 ;
        RECT 162.600 374.800 163.400 375.600 ;
        RECT 162.600 374.400 163.200 374.800 ;
        RECT 156.400 374.200 158.000 374.400 ;
        RECT 147.000 373.600 158.000 374.200 ;
        RECT 159.600 373.600 161.200 374.400 ;
        RECT 162.400 373.600 163.200 374.400 ;
        RECT 145.200 372.800 146.000 373.000 ;
        RECT 142.200 372.200 146.000 372.800 ;
        RECT 142.200 372.000 143.000 372.200 ;
        RECT 143.800 371.400 144.600 371.600 ;
        RECT 129.200 371.000 134.800 371.200 ;
        RECT 129.000 370.800 134.800 371.000 ;
        RECT 121.200 369.800 123.600 370.400 ;
        RECT 125.000 370.600 134.800 370.800 ;
        RECT 125.000 370.200 129.800 370.600 ;
        RECT 121.200 368.800 121.800 369.800 ;
        RECT 120.400 368.000 121.800 368.800 ;
        RECT 123.400 369.000 124.200 369.200 ;
        RECT 125.000 369.000 125.600 370.200 ;
        RECT 123.400 368.400 125.600 369.000 ;
        RECT 126.200 369.000 131.600 369.600 ;
        RECT 126.200 368.800 127.000 369.000 ;
        RECT 130.800 368.800 131.600 369.000 ;
        RECT 124.600 367.400 125.400 367.600 ;
        RECT 127.400 367.400 128.200 367.600 ;
        RECT 121.200 366.200 122.000 367.000 ;
        RECT 124.600 366.800 128.200 367.400 ;
        RECT 125.400 366.200 126.000 366.800 ;
        RECT 130.800 366.200 131.600 367.000 ;
        RECT 120.600 362.200 121.800 366.200 ;
        RECT 125.200 362.200 126.000 366.200 ;
        RECT 129.600 365.600 131.600 366.200 ;
        RECT 129.600 362.200 130.400 365.600 ;
        RECT 134.000 362.200 134.800 370.600 ;
        RECT 140.400 370.800 144.600 371.400 ;
        RECT 140.400 362.200 141.200 370.800 ;
        RECT 147.000 370.400 147.600 373.600 ;
        RECT 154.200 373.400 155.000 373.600 ;
        RECT 164.000 372.800 164.600 376.200 ;
        RECT 169.200 375.800 170.000 379.800 ;
        RECT 174.600 376.000 175.400 379.000 ;
        RECT 178.800 377.000 179.600 379.000 ;
        RECT 182.000 377.800 182.800 379.800 ;
        RECT 165.200 375.400 166.800 375.600 ;
        RECT 165.200 374.800 167.200 375.400 ;
        RECT 167.800 375.200 170.000 375.800 ;
        RECT 173.800 375.400 175.400 376.000 ;
        RECT 167.800 375.000 168.600 375.200 ;
        RECT 173.800 375.000 174.600 375.400 ;
        RECT 166.600 374.400 167.200 374.800 ;
        RECT 173.800 374.400 174.400 375.000 ;
        RECT 179.000 374.800 179.600 377.000 ;
        RECT 180.400 375.600 181.200 377.200 ;
        RECT 166.600 374.300 170.000 374.400 ;
        RECT 172.400 374.300 174.400 374.400 ;
        RECT 165.200 373.400 166.000 374.200 ;
        RECT 166.600 373.800 174.400 374.300 ;
        RECT 175.400 374.200 179.600 374.800 ;
        RECT 182.200 374.400 182.800 377.800 ;
        RECT 188.400 375.800 189.200 379.800 ;
        RECT 189.800 376.400 190.600 377.200 ;
        RECT 192.200 376.400 193.000 379.800 ;
        RECT 199.000 378.400 199.800 379.800 ;
        RECT 198.000 377.600 199.800 378.400 ;
        RECT 199.000 376.400 199.800 377.600 ;
        RECT 203.800 376.400 204.600 379.800 ;
        RECT 182.000 374.300 182.800 374.400 ;
        RECT 186.800 374.300 187.600 374.400 ;
        RECT 175.400 373.800 176.400 374.200 ;
        RECT 168.400 373.700 174.400 373.800 ;
        RECT 168.400 373.600 170.000 373.700 ;
        RECT 172.400 373.600 174.400 373.700 ;
        RECT 153.200 372.400 154.000 372.600 ;
        RECT 155.800 372.400 156.600 372.600 ;
        RECT 163.600 372.400 164.600 372.800 ;
        RECT 151.600 371.800 156.600 372.400 ;
        RECT 162.800 372.200 164.600 372.400 ;
        RECT 165.400 372.800 166.000 373.400 ;
        RECT 165.400 372.200 168.000 372.800 ;
        RECT 151.600 371.600 152.400 371.800 ;
        RECT 162.800 371.600 164.200 372.200 ;
        RECT 167.200 372.000 168.000 372.200 ;
        RECT 153.200 371.000 158.800 371.200 ;
        RECT 153.000 370.800 158.800 371.000 ;
        RECT 145.200 369.800 147.600 370.400 ;
        RECT 149.000 370.600 158.800 370.800 ;
        RECT 149.000 370.200 153.800 370.600 ;
        RECT 145.200 368.800 145.800 369.800 ;
        RECT 144.400 368.000 145.800 368.800 ;
        RECT 147.400 369.000 148.200 369.200 ;
        RECT 149.000 369.000 149.600 370.200 ;
        RECT 147.400 368.400 149.600 369.000 ;
        RECT 150.200 369.000 155.600 369.600 ;
        RECT 150.200 368.800 151.000 369.000 ;
        RECT 154.800 368.800 155.600 369.000 ;
        RECT 148.600 367.400 149.400 367.600 ;
        RECT 151.400 367.400 152.200 367.600 ;
        RECT 145.200 366.200 146.000 367.000 ;
        RECT 148.600 366.800 152.200 367.400 ;
        RECT 149.400 366.200 150.000 366.800 ;
        RECT 154.800 366.200 155.600 367.000 ;
        RECT 144.600 362.200 145.800 366.200 ;
        RECT 149.200 362.200 150.000 366.200 ;
        RECT 153.600 365.600 155.600 366.200 ;
        RECT 153.600 362.200 154.400 365.600 ;
        RECT 158.000 362.200 158.800 370.600 ;
        RECT 163.600 370.400 164.200 371.600 ;
        RECT 165.000 371.400 165.800 371.600 ;
        RECT 165.000 370.800 168.400 371.400 ;
        RECT 172.400 370.800 173.200 372.400 ;
        RECT 162.800 370.200 164.200 370.400 ;
        RECT 167.800 370.200 168.400 370.800 ;
        RECT 159.600 369.600 162.000 370.200 ;
        RECT 162.800 369.600 165.600 370.200 ;
        RECT 159.600 362.200 160.400 369.600 ;
        RECT 161.200 369.400 162.000 369.600 ;
        RECT 164.000 362.200 165.600 369.600 ;
        RECT 167.800 369.600 170.000 370.200 ;
        RECT 167.800 369.400 168.600 369.600 ;
        RECT 169.200 362.200 170.000 369.600 ;
        RECT 173.800 369.800 174.400 373.600 ;
        RECT 175.000 373.000 176.400 373.800 ;
        RECT 182.000 373.700 187.600 374.300 ;
        RECT 182.000 373.600 182.800 373.700 ;
        RECT 175.800 371.000 176.400 373.000 ;
        RECT 177.200 371.600 178.000 373.200 ;
        RECT 178.800 371.600 179.600 373.200 ;
        RECT 175.800 370.400 179.600 371.000 ;
        RECT 173.800 369.200 175.400 369.800 ;
        RECT 174.600 362.200 175.400 369.200 ;
        RECT 179.000 367.000 179.600 370.400 ;
        RECT 182.200 370.200 182.800 373.600 ;
        RECT 186.800 372.800 187.600 373.700 ;
        RECT 183.600 370.800 184.400 372.400 ;
        RECT 185.200 372.200 186.000 372.400 ;
        RECT 188.400 372.200 189.000 375.800 ;
        RECT 190.000 375.600 190.800 376.400 ;
        RECT 191.600 375.600 194.000 376.400 ;
        RECT 190.100 374.300 190.700 375.600 ;
        RECT 191.600 374.300 192.400 374.400 ;
        RECT 190.100 373.700 192.400 374.300 ;
        RECT 191.600 373.600 192.400 373.700 ;
        RECT 190.000 372.200 190.800 372.400 ;
        RECT 185.200 371.600 186.800 372.200 ;
        RECT 188.400 371.600 190.800 372.200 ;
        RECT 193.200 372.300 194.000 375.600 ;
        RECT 198.000 375.800 199.800 376.400 ;
        RECT 202.800 375.800 204.600 376.400 ;
        RECT 206.000 376.000 206.800 379.800 ;
        RECT 209.200 376.000 210.000 379.800 ;
        RECT 206.000 375.800 210.000 376.000 ;
        RECT 210.800 375.800 211.600 379.800 ;
        RECT 215.000 376.400 215.800 379.800 ;
        RECT 214.000 375.800 215.800 376.400 ;
        RECT 217.800 376.400 218.600 379.800 ;
        RECT 217.800 375.800 219.600 376.400 ;
        RECT 194.800 373.600 195.600 375.200 ;
        RECT 196.400 373.600 197.200 375.200 ;
        RECT 196.500 372.300 197.100 373.600 ;
        RECT 193.200 371.700 197.100 372.300 ;
        RECT 186.000 371.200 186.800 371.600 ;
        RECT 190.000 370.200 190.600 371.600 ;
        RECT 182.000 369.400 183.800 370.200 ;
        RECT 178.800 363.000 179.600 367.000 ;
        RECT 183.000 362.200 183.800 369.400 ;
        RECT 185.200 369.600 189.200 370.200 ;
        RECT 185.200 362.200 186.000 369.600 ;
        RECT 188.400 362.200 189.200 369.600 ;
        RECT 190.000 362.200 190.800 370.200 ;
        RECT 191.600 368.800 192.400 370.400 ;
        RECT 193.200 362.200 194.000 371.700 ;
        RECT 198.000 362.200 198.800 375.800 ;
        RECT 199.600 374.300 200.400 374.400 ;
        RECT 201.200 374.300 202.000 375.200 ;
        RECT 199.600 373.700 202.000 374.300 ;
        RECT 199.600 373.600 200.400 373.700 ;
        RECT 201.200 373.600 202.000 373.700 ;
        RECT 202.800 374.300 203.600 375.800 ;
        RECT 206.200 375.400 209.800 375.800 ;
        RECT 206.800 374.400 207.600 374.800 ;
        RECT 210.800 374.400 211.400 375.800 ;
        RECT 206.000 374.300 207.600 374.400 ;
        RECT 202.800 373.800 207.600 374.300 ;
        RECT 202.800 373.700 206.800 373.800 ;
        RECT 199.600 368.800 200.400 370.400 ;
        RECT 202.800 362.200 203.600 373.700 ;
        RECT 206.000 373.600 206.800 373.700 ;
        RECT 209.000 373.600 211.600 374.400 ;
        RECT 212.400 373.600 213.200 375.200 ;
        RECT 207.600 371.600 208.400 373.200 ;
        RECT 204.400 368.800 205.200 370.400 ;
        RECT 209.000 370.200 209.600 373.600 ;
        RECT 210.800 372.300 211.600 372.400 ;
        RECT 214.000 372.300 214.800 375.800 ;
        RECT 218.800 372.300 219.600 375.800 ;
        RECT 220.400 373.600 221.200 375.200 ;
        RECT 210.800 371.700 214.800 372.300 ;
        RECT 210.800 371.600 211.600 371.700 ;
        RECT 210.800 370.300 211.600 370.400 ;
        RECT 212.400 370.300 213.200 370.400 ;
        RECT 210.800 370.200 213.200 370.300 ;
        RECT 208.600 369.600 209.600 370.200 ;
        RECT 210.200 369.700 213.200 370.200 ;
        RECT 210.200 369.600 211.600 369.700 ;
        RECT 212.400 369.600 213.200 369.700 ;
        RECT 208.600 368.400 209.400 369.600 ;
        RECT 210.200 368.400 210.800 369.600 ;
        RECT 207.600 367.600 209.400 368.400 ;
        RECT 210.000 367.600 210.800 368.400 ;
        RECT 208.600 362.200 209.400 367.600 ;
        RECT 214.000 362.200 214.800 371.700 ;
        RECT 215.700 371.700 219.600 372.300 ;
        RECT 215.700 370.400 216.300 371.700 ;
        RECT 215.600 368.800 216.400 370.400 ;
        RECT 217.200 368.800 218.000 370.400 ;
        RECT 218.800 362.200 219.600 371.700 ;
        RECT 222.000 362.200 222.800 379.800 ;
        RECT 225.800 376.400 226.600 379.800 ;
        RECT 225.800 375.800 227.600 376.400 ;
        RECT 223.600 373.600 224.400 375.200 ;
        RECT 225.200 374.300 226.000 374.400 ;
        RECT 226.800 374.300 227.600 375.800 ;
        RECT 230.000 375.800 230.800 379.800 ;
        RECT 234.400 378.400 236.000 379.800 ;
        RECT 233.200 377.600 236.000 378.400 ;
        RECT 234.400 376.200 236.000 377.600 ;
        RECT 230.000 375.200 232.600 375.800 ;
        RECT 225.200 373.700 227.600 374.300 ;
        RECT 225.200 373.600 226.000 373.700 ;
        RECT 225.200 368.800 226.000 370.400 ;
        RECT 226.800 362.200 227.600 373.700 ;
        RECT 228.400 373.600 229.200 375.200 ;
        RECT 231.800 375.000 232.600 375.200 ;
        RECT 233.200 374.800 234.800 375.600 ;
        RECT 230.000 374.200 231.600 374.400 ;
        RECT 235.400 374.200 236.000 376.200 ;
        RECT 239.600 375.800 240.400 379.800 ;
        RECT 236.600 374.800 237.400 375.600 ;
        RECT 238.000 375.200 240.400 375.800 ;
        RECT 238.000 375.000 238.800 375.200 ;
        RECT 230.000 374.000 232.200 374.200 ;
        RECT 230.000 373.600 234.400 374.000 ;
        RECT 231.600 373.400 234.400 373.600 ;
        RECT 233.600 373.200 234.400 373.400 ;
        RECT 235.000 373.600 236.000 374.200 ;
        RECT 236.800 374.400 237.400 374.800 ;
        RECT 236.800 373.600 237.600 374.400 ;
        RECT 238.800 373.600 240.400 374.400 ;
        RECT 235.000 372.400 235.600 373.600 ;
        RECT 232.200 372.200 233.000 372.400 ;
        RECT 232.200 371.600 233.800 372.200 ;
        RECT 234.800 371.600 235.600 372.400 ;
        RECT 233.000 371.400 233.800 371.600 ;
        RECT 235.000 370.200 235.600 371.600 ;
        RECT 241.200 372.300 242.000 379.800 ;
        RECT 242.800 375.600 243.600 377.200 ;
        RECT 246.000 376.400 246.800 379.800 ;
        RECT 245.800 375.800 246.800 376.400 ;
        RECT 245.800 374.400 246.400 375.800 ;
        RECT 249.200 375.200 250.000 379.800 ;
        RECT 250.800 379.200 254.800 379.800 ;
        RECT 250.800 375.800 251.600 379.200 ;
        RECT 252.400 375.800 253.200 378.600 ;
        RECT 254.000 376.000 254.800 379.200 ;
        RECT 257.200 376.000 258.000 379.800 ;
        RECT 261.400 378.400 262.200 379.800 ;
        RECT 261.400 377.600 262.800 378.400 ;
        RECT 261.400 376.400 262.200 377.600 ;
        RECT 254.000 375.800 258.000 376.000 ;
        RECT 260.400 375.800 262.200 376.400 ;
        RECT 263.600 375.800 264.400 379.800 ;
        RECT 265.200 376.000 266.000 379.800 ;
        RECT 268.400 376.000 269.200 379.800 ;
        RECT 270.200 376.400 271.000 377.200 ;
        RECT 265.200 375.800 269.200 376.000 ;
        RECT 247.400 374.600 250.000 375.200 ;
        RECT 245.800 373.600 246.800 374.400 ;
        RECT 244.400 372.300 245.200 372.400 ;
        RECT 241.200 371.700 245.200 372.300 ;
        RECT 230.000 369.600 232.600 370.200 ;
        RECT 230.000 362.200 230.800 369.600 ;
        RECT 231.800 369.400 232.600 369.600 ;
        RECT 234.400 362.200 236.000 370.200 ;
        RECT 238.000 369.600 240.400 370.200 ;
        RECT 238.000 369.400 238.800 369.600 ;
        RECT 239.600 362.200 240.400 369.600 ;
        RECT 241.200 362.200 242.000 371.700 ;
        RECT 244.400 371.600 245.200 371.700 ;
        RECT 245.800 370.200 246.400 373.600 ;
        RECT 247.400 373.000 248.000 374.600 ;
        RECT 252.400 374.400 253.000 375.800 ;
        RECT 254.200 375.400 257.800 375.800 ;
        RECT 256.400 374.400 257.200 374.800 ;
        RECT 247.000 372.200 248.000 373.000 ;
        RECT 247.400 370.200 248.000 372.200 ;
        RECT 249.000 372.400 249.800 373.200 ;
        RECT 250.800 372.800 251.600 374.400 ;
        RECT 252.400 373.800 254.800 374.400 ;
        RECT 256.400 374.300 258.000 374.400 ;
        RECT 258.800 374.300 259.600 375.200 ;
        RECT 256.400 373.800 259.600 374.300 ;
        RECT 254.000 373.600 254.800 373.800 ;
        RECT 257.200 373.700 259.600 373.800 ;
        RECT 257.200 373.600 258.000 373.700 ;
        RECT 258.800 373.600 259.600 373.700 ;
        RECT 249.000 371.600 250.000 372.400 ;
        RECT 252.400 371.600 253.200 373.200 ;
        RECT 254.200 370.200 254.800 373.600 ;
        RECT 255.600 371.600 256.400 373.200 ;
        RECT 245.800 369.200 246.800 370.200 ;
        RECT 247.400 369.600 250.000 370.200 ;
        RECT 246.000 362.200 246.800 369.200 ;
        RECT 249.200 362.200 250.000 369.600 ;
        RECT 253.400 368.400 255.400 370.200 ;
        RECT 253.400 367.600 256.400 368.400 ;
        RECT 253.400 362.200 255.400 367.600 ;
        RECT 260.400 362.200 261.200 375.800 ;
        RECT 263.800 374.400 264.400 375.800 ;
        RECT 265.400 375.400 269.000 375.800 ;
        RECT 270.000 375.600 270.800 376.400 ;
        RECT 271.600 375.800 272.400 379.800 ;
        RECT 267.600 374.400 268.400 374.800 ;
        RECT 263.600 373.600 266.200 374.400 ;
        RECT 267.600 373.800 269.200 374.400 ;
        RECT 268.400 373.600 269.200 373.800 ;
        RECT 262.000 368.800 262.800 370.400 ;
        RECT 263.600 370.200 264.400 370.400 ;
        RECT 265.600 370.200 266.200 373.600 ;
        RECT 266.800 371.600 267.600 373.200 ;
        RECT 270.000 372.200 270.800 372.400 ;
        RECT 271.800 372.200 272.400 375.800 ;
        RECT 273.200 372.800 274.000 374.400 ;
        RECT 274.800 372.200 275.600 372.400 ;
        RECT 270.000 371.600 272.400 372.200 ;
        RECT 274.000 371.600 275.600 372.200 ;
        RECT 276.400 372.300 277.200 379.800 ;
        RECT 278.000 375.600 278.800 377.200 ;
        RECT 279.600 376.000 280.400 379.800 ;
        RECT 282.800 376.000 283.600 379.800 ;
        RECT 279.600 375.800 283.600 376.000 ;
        RECT 284.400 375.800 285.200 379.800 ;
        RECT 286.600 376.400 287.400 379.800 ;
        RECT 286.600 375.800 288.400 376.400 ;
        RECT 279.800 375.400 283.400 375.800 ;
        RECT 280.400 374.400 281.200 374.800 ;
        RECT 284.400 374.400 285.000 375.800 ;
        RECT 279.600 373.800 281.200 374.400 ;
        RECT 279.600 373.600 280.400 373.800 ;
        RECT 282.600 373.600 285.200 374.400 ;
        RECT 281.200 372.300 282.000 373.200 ;
        RECT 276.400 371.700 282.000 372.300 ;
        RECT 270.200 370.200 270.800 371.600 ;
        RECT 274.000 371.200 274.800 371.600 ;
        RECT 263.600 369.600 265.000 370.200 ;
        RECT 265.600 369.600 266.600 370.200 ;
        RECT 264.400 368.400 265.000 369.600 ;
        RECT 264.400 367.600 265.200 368.400 ;
        RECT 265.800 364.400 266.600 369.600 ;
        RECT 265.800 363.600 267.600 364.400 ;
        RECT 265.800 362.200 266.600 363.600 ;
        RECT 270.000 362.200 270.800 370.200 ;
        RECT 271.600 369.600 275.600 370.200 ;
        RECT 271.600 362.200 272.400 369.600 ;
        RECT 274.800 362.200 275.600 369.600 ;
        RECT 276.400 362.200 277.200 371.700 ;
        RECT 281.200 371.600 282.000 371.700 ;
        RECT 282.600 370.200 283.200 373.600 ;
        RECT 287.600 372.300 288.400 375.800 ;
        RECT 295.600 375.200 296.400 379.800 ;
        RECT 298.800 376.400 299.600 379.800 ;
        RECT 298.800 375.800 299.800 376.400 ;
        RECT 289.200 373.600 290.000 375.200 ;
        RECT 295.600 374.600 298.200 375.200 ;
        RECT 295.800 372.400 296.600 373.200 ;
        RECT 284.500 371.700 288.400 372.300 ;
        RECT 284.500 370.400 285.100 371.700 ;
        RECT 284.400 370.200 285.200 370.400 ;
        RECT 282.200 369.600 283.200 370.200 ;
        RECT 283.800 369.600 285.200 370.200 ;
        RECT 282.200 362.200 283.000 369.600 ;
        RECT 283.800 368.400 284.400 369.600 ;
        RECT 286.000 368.800 286.800 370.400 ;
        RECT 283.600 367.600 284.400 368.400 ;
        RECT 287.600 362.200 288.400 371.700 ;
        RECT 289.200 372.300 290.000 372.400 ;
        RECT 295.600 372.300 296.600 372.400 ;
        RECT 289.200 371.700 296.600 372.300 ;
        RECT 289.200 371.600 290.000 371.700 ;
        RECT 295.600 371.600 296.600 371.700 ;
        RECT 297.600 373.000 298.200 374.600 ;
        RECT 299.200 374.400 299.800 375.800 ;
        RECT 302.000 375.600 302.800 377.200 ;
        RECT 298.800 374.300 299.800 374.400 ;
        RECT 302.000 374.300 302.800 374.400 ;
        RECT 298.800 373.700 302.800 374.300 ;
        RECT 298.800 373.600 299.800 373.700 ;
        RECT 302.000 373.600 302.800 373.700 ;
        RECT 297.600 372.200 298.600 373.000 ;
        RECT 297.600 370.200 298.200 372.200 ;
        RECT 299.200 370.200 299.800 373.600 ;
        RECT 295.600 369.600 298.200 370.200 ;
        RECT 295.600 362.200 296.400 369.600 ;
        RECT 298.800 369.200 299.800 370.200 ;
        RECT 303.600 372.300 304.400 379.800 ;
        RECT 305.200 376.000 306.000 379.800 ;
        RECT 308.400 376.000 309.200 379.800 ;
        RECT 305.200 375.800 309.200 376.000 ;
        RECT 310.000 375.800 310.800 379.800 ;
        RECT 305.400 375.400 309.000 375.800 ;
        RECT 306.000 374.400 306.800 374.800 ;
        RECT 310.000 374.400 310.600 375.800 ;
        RECT 311.600 375.400 312.400 379.800 ;
        RECT 315.800 378.400 317.000 379.800 ;
        RECT 315.800 377.800 317.200 378.400 ;
        RECT 320.400 377.800 321.200 379.800 ;
        RECT 324.800 378.400 325.600 379.800 ;
        RECT 324.800 377.800 326.800 378.400 ;
        RECT 316.400 377.000 317.200 377.800 ;
        RECT 320.600 377.200 321.200 377.800 ;
        RECT 320.600 376.600 323.400 377.200 ;
        RECT 322.600 376.400 323.400 376.600 ;
        RECT 324.400 376.400 325.200 377.200 ;
        RECT 326.000 377.000 326.800 377.800 ;
        RECT 314.600 375.400 315.400 375.600 ;
        RECT 311.600 374.800 315.400 375.400 ;
        RECT 305.200 373.800 306.800 374.400 ;
        RECT 305.200 373.600 306.000 373.800 ;
        RECT 308.200 373.600 310.800 374.400 ;
        RECT 306.800 372.300 307.600 373.200 ;
        RECT 303.600 371.700 307.600 372.300 ;
        RECT 298.800 362.200 299.600 369.200 ;
        RECT 303.600 362.200 304.400 371.700 ;
        RECT 306.800 371.600 307.600 371.700 ;
        RECT 308.200 370.200 308.800 373.600 ;
        RECT 311.600 371.400 312.400 374.800 ;
        RECT 318.600 374.200 319.400 374.400 ;
        RECT 324.400 374.200 325.000 376.400 ;
        RECT 329.200 375.000 330.000 379.800 ;
        RECT 330.800 375.400 331.600 379.800 ;
        RECT 335.000 378.400 336.200 379.800 ;
        RECT 335.000 377.800 336.400 378.400 ;
        RECT 339.600 377.800 340.400 379.800 ;
        RECT 344.000 378.400 344.800 379.800 ;
        RECT 344.000 377.800 346.000 378.400 ;
        RECT 335.600 377.000 336.400 377.800 ;
        RECT 339.800 377.200 340.400 377.800 ;
        RECT 339.800 376.600 342.600 377.200 ;
        RECT 341.800 376.400 342.600 376.600 ;
        RECT 343.600 376.400 344.400 377.200 ;
        RECT 345.200 377.000 346.000 377.800 ;
        RECT 333.800 375.400 334.600 375.600 ;
        RECT 330.800 374.800 334.600 375.400 ;
        RECT 327.600 374.200 329.200 374.400 ;
        RECT 318.200 373.600 329.200 374.200 ;
        RECT 316.400 372.800 317.200 373.000 ;
        RECT 313.400 372.200 317.200 372.800 ;
        RECT 318.200 372.300 318.800 373.600 ;
        RECT 325.400 373.400 326.200 373.600 ;
        RECT 324.400 372.400 325.200 372.600 ;
        RECT 327.000 372.400 327.800 372.600 ;
        RECT 319.600 372.300 320.400 372.400 ;
        RECT 313.400 372.000 314.200 372.200 ;
        RECT 318.100 371.700 320.400 372.300 ;
        RECT 315.000 371.400 315.800 371.600 ;
        RECT 311.600 370.800 315.800 371.400 ;
        RECT 310.000 370.200 310.800 370.400 ;
        RECT 307.800 369.600 308.800 370.200 ;
        RECT 309.400 369.600 310.800 370.200 ;
        RECT 307.800 364.400 308.600 369.600 ;
        RECT 309.400 368.400 310.000 369.600 ;
        RECT 309.200 367.600 310.000 368.400 ;
        RECT 306.800 363.600 308.600 364.400 ;
        RECT 307.800 362.200 308.600 363.600 ;
        RECT 311.600 362.200 312.400 370.800 ;
        RECT 318.200 370.400 318.800 371.700 ;
        RECT 319.600 371.600 320.400 371.700 ;
        RECT 322.800 371.800 327.800 372.400 ;
        RECT 322.800 371.600 323.600 371.800 ;
        RECT 330.800 371.400 331.600 374.800 ;
        RECT 337.800 374.200 338.600 374.400 ;
        RECT 343.600 374.200 344.200 376.400 ;
        RECT 348.400 375.000 349.200 379.800 ;
        RECT 350.000 376.000 350.800 379.800 ;
        RECT 353.200 376.000 354.000 379.800 ;
        RECT 350.000 375.800 354.000 376.000 ;
        RECT 354.800 375.800 355.600 379.800 ;
        RECT 350.200 375.400 353.800 375.800 ;
        RECT 350.800 374.400 351.600 374.800 ;
        RECT 354.800 374.400 355.400 375.800 ;
        RECT 346.800 374.200 348.400 374.400 ;
        RECT 337.400 373.600 348.400 374.200 ;
        RECT 350.000 373.800 351.600 374.400 ;
        RECT 350.000 373.600 350.800 373.800 ;
        RECT 353.000 373.600 355.600 374.400 ;
        RECT 335.600 372.800 336.400 373.000 ;
        RECT 332.600 372.200 336.400 372.800 ;
        RECT 337.400 372.300 338.000 373.600 ;
        RECT 344.600 373.400 345.400 373.600 ;
        RECT 343.600 372.400 344.400 372.600 ;
        RECT 346.200 372.400 347.000 372.600 ;
        RECT 338.800 372.300 339.600 372.400 ;
        RECT 332.600 372.000 333.400 372.200 ;
        RECT 337.300 371.700 339.600 372.300 ;
        RECT 334.200 371.400 335.000 371.600 ;
        RECT 324.400 371.000 330.000 371.200 ;
        RECT 324.200 370.800 330.000 371.000 ;
        RECT 316.400 369.800 318.800 370.400 ;
        RECT 320.200 370.600 330.000 370.800 ;
        RECT 320.200 370.200 325.000 370.600 ;
        RECT 316.400 368.800 317.000 369.800 ;
        RECT 315.600 368.000 317.000 368.800 ;
        RECT 318.600 369.000 319.400 369.200 ;
        RECT 320.200 369.000 320.800 370.200 ;
        RECT 318.600 368.400 320.800 369.000 ;
        RECT 321.400 369.000 326.800 369.600 ;
        RECT 321.400 368.800 322.200 369.000 ;
        RECT 326.000 368.800 326.800 369.000 ;
        RECT 319.800 367.400 320.600 367.600 ;
        RECT 322.600 367.400 323.400 367.600 ;
        RECT 316.400 366.200 317.200 367.000 ;
        RECT 319.800 366.800 323.400 367.400 ;
        RECT 320.600 366.200 321.200 366.800 ;
        RECT 326.000 366.200 326.800 367.000 ;
        RECT 315.800 362.200 317.000 366.200 ;
        RECT 320.400 362.200 321.200 366.200 ;
        RECT 324.800 365.600 326.800 366.200 ;
        RECT 324.800 362.200 325.600 365.600 ;
        RECT 329.200 362.200 330.000 370.600 ;
        RECT 330.800 370.800 335.000 371.400 ;
        RECT 330.800 362.200 331.600 370.800 ;
        RECT 337.400 370.400 338.000 371.700 ;
        RECT 338.800 371.600 339.600 371.700 ;
        RECT 342.000 371.800 347.000 372.400 ;
        RECT 342.000 371.600 342.800 371.800 ;
        RECT 351.600 371.600 352.400 373.200 ;
        RECT 353.000 372.400 353.600 373.600 ;
        RECT 356.400 372.400 357.200 379.800 ;
        RECT 359.600 375.200 360.400 379.800 ;
        RECT 361.200 376.000 362.000 379.800 ;
        RECT 364.400 376.000 365.200 379.800 ;
        RECT 361.200 375.800 365.200 376.000 ;
        RECT 366.000 375.800 366.800 379.800 ;
        RECT 369.200 377.600 370.000 379.800 ;
        RECT 374.000 377.800 374.800 379.800 ;
        RECT 361.400 375.400 365.000 375.800 ;
        RECT 358.200 374.600 360.400 375.200 ;
        RECT 353.000 371.600 354.000 372.400 ;
        RECT 343.600 371.000 349.200 371.200 ;
        RECT 343.400 370.800 349.200 371.000 ;
        RECT 335.600 369.800 338.000 370.400 ;
        RECT 339.400 370.600 349.200 370.800 ;
        RECT 339.400 370.200 344.200 370.600 ;
        RECT 335.600 368.800 336.200 369.800 ;
        RECT 334.800 368.000 336.200 368.800 ;
        RECT 337.800 369.000 338.600 369.200 ;
        RECT 339.400 369.000 340.000 370.200 ;
        RECT 337.800 368.400 340.000 369.000 ;
        RECT 340.600 369.000 346.000 369.600 ;
        RECT 340.600 368.800 341.400 369.000 ;
        RECT 345.200 368.800 346.000 369.000 ;
        RECT 339.000 367.400 339.800 367.600 ;
        RECT 341.800 367.400 342.600 367.600 ;
        RECT 335.600 366.200 336.400 367.000 ;
        RECT 339.000 366.800 342.600 367.400 ;
        RECT 339.800 366.200 340.400 366.800 ;
        RECT 345.200 366.200 346.000 367.000 ;
        RECT 335.000 362.200 336.200 366.200 ;
        RECT 339.600 362.200 340.400 366.200 ;
        RECT 344.000 365.600 346.000 366.200 ;
        RECT 344.000 362.200 344.800 365.600 ;
        RECT 348.400 362.200 349.200 370.600 ;
        RECT 353.000 370.200 353.600 371.600 ;
        RECT 354.800 370.200 355.600 370.400 ;
        RECT 352.600 369.600 353.600 370.200 ;
        RECT 354.200 369.600 355.600 370.200 ;
        RECT 356.400 370.200 357.000 372.400 ;
        RECT 358.200 371.600 358.800 374.600 ;
        RECT 362.000 374.400 362.800 374.800 ;
        RECT 366.000 374.400 366.600 375.800 ;
        RECT 369.200 374.400 369.800 377.600 ;
        RECT 370.800 375.600 371.600 377.200 ;
        RECT 372.400 375.600 373.200 377.200 ;
        RECT 361.200 373.800 362.800 374.400 ;
        RECT 361.200 373.600 362.000 373.800 ;
        RECT 364.200 373.600 366.800 374.400 ;
        RECT 369.200 373.600 370.000 374.400 ;
        RECT 370.900 374.300 371.500 375.600 ;
        RECT 374.200 374.400 374.800 377.800 ;
        RECT 377.200 375.800 378.000 379.800 ;
        RECT 378.800 376.000 379.600 379.800 ;
        RECT 382.000 376.000 382.800 379.800 ;
        RECT 378.800 375.800 382.800 376.000 ;
        RECT 377.400 374.400 378.000 375.800 ;
        RECT 379.000 375.400 382.600 375.800 ;
        RECT 381.200 374.400 382.000 374.800 ;
        RECT 374.000 374.300 374.800 374.400 ;
        RECT 370.900 373.700 374.800 374.300 ;
        RECT 374.000 373.600 374.800 373.700 ;
        RECT 377.200 373.600 379.800 374.400 ;
        RECT 381.200 373.800 382.800 374.400 ;
        RECT 382.000 373.600 382.800 373.800 ;
        RECT 359.600 372.300 360.400 373.200 ;
        RECT 362.800 372.300 363.600 373.200 ;
        RECT 359.600 371.700 363.600 372.300 ;
        RECT 359.600 371.600 360.400 371.700 ;
        RECT 362.800 371.600 363.600 371.700 ;
        RECT 364.200 372.400 364.800 373.600 ;
        RECT 364.200 371.600 365.200 372.400 ;
        RECT 357.600 370.800 358.800 371.600 ;
        RECT 358.200 370.200 358.800 370.800 ;
        RECT 364.200 370.200 364.800 371.600 ;
        RECT 367.600 370.800 368.400 372.400 ;
        RECT 366.000 370.200 366.800 370.400 ;
        RECT 369.200 370.200 369.800 373.600 ;
        RECT 374.200 370.200 374.800 373.600 ;
        RECT 375.600 370.800 376.400 372.400 ;
        RECT 377.200 370.200 378.000 370.400 ;
        RECT 379.200 370.200 379.800 373.600 ;
        RECT 380.400 372.300 381.200 373.200 ;
        RECT 383.600 372.300 384.400 379.800 ;
        RECT 385.200 375.600 386.000 377.200 ;
        RECT 380.400 371.700 384.400 372.300 ;
        RECT 380.400 371.600 381.200 371.700 ;
        RECT 352.600 362.200 353.400 369.600 ;
        RECT 354.200 368.400 354.800 369.600 ;
        RECT 354.000 367.600 354.800 368.400 ;
        RECT 356.400 362.200 357.200 370.200 ;
        RECT 358.200 369.600 360.400 370.200 ;
        RECT 359.600 362.200 360.400 369.600 ;
        RECT 363.800 369.600 364.800 370.200 ;
        RECT 365.400 369.600 366.800 370.200 ;
        RECT 363.800 362.200 364.600 369.600 ;
        RECT 365.400 368.400 366.000 369.600 ;
        RECT 365.200 367.600 366.000 368.400 ;
        RECT 368.200 369.400 370.000 370.200 ;
        RECT 374.000 369.400 375.800 370.200 ;
        RECT 377.200 369.600 378.600 370.200 ;
        RECT 379.200 369.600 380.200 370.200 ;
        RECT 368.200 364.400 369.000 369.400 ;
        RECT 368.200 363.600 370.000 364.400 ;
        RECT 368.200 362.200 369.000 363.600 ;
        RECT 375.000 362.200 375.800 369.400 ;
        RECT 378.000 368.400 378.600 369.600 ;
        RECT 379.400 368.400 380.200 369.600 ;
        RECT 378.000 367.600 378.800 368.400 ;
        RECT 379.400 367.600 381.200 368.400 ;
        RECT 379.400 362.200 380.200 367.600 ;
        RECT 383.600 362.200 384.400 371.700 ;
        RECT 386.800 375.400 387.600 379.800 ;
        RECT 391.000 378.400 392.200 379.800 ;
        RECT 391.000 377.800 392.400 378.400 ;
        RECT 395.600 377.800 396.400 379.800 ;
        RECT 400.000 378.400 400.800 379.800 ;
        RECT 400.000 377.800 402.000 378.400 ;
        RECT 391.600 377.000 392.400 377.800 ;
        RECT 395.800 377.200 396.400 377.800 ;
        RECT 395.800 376.600 398.600 377.200 ;
        RECT 397.800 376.400 398.600 376.600 ;
        RECT 399.600 376.400 400.400 377.200 ;
        RECT 401.200 377.000 402.000 377.800 ;
        RECT 389.800 375.400 390.600 375.600 ;
        RECT 386.800 374.800 390.600 375.400 ;
        RECT 386.800 371.400 387.600 374.800 ;
        RECT 393.800 374.200 394.600 374.400 ;
        RECT 399.600 374.200 400.200 376.400 ;
        RECT 404.400 375.000 405.200 379.800 ;
        RECT 402.800 374.200 404.400 374.400 ;
        RECT 393.400 373.600 404.400 374.200 ;
        RECT 391.600 372.800 392.400 373.000 ;
        RECT 388.600 372.200 392.400 372.800 ;
        RECT 393.400 372.400 394.000 373.600 ;
        RECT 400.600 373.400 401.400 373.600 ;
        RECT 399.600 372.400 400.400 372.600 ;
        RECT 402.200 372.400 403.000 372.600 ;
        RECT 388.600 372.000 389.400 372.200 ;
        RECT 393.200 371.600 394.000 372.400 ;
        RECT 398.000 371.800 403.000 372.400 ;
        RECT 406.000 372.300 406.800 372.400 ;
        RECT 407.600 372.300 408.400 379.800 ;
        RECT 412.400 376.000 413.200 379.800 ;
        RECT 412.200 375.200 413.200 376.000 ;
        RECT 409.200 374.300 410.000 375.200 ;
        RECT 410.800 374.300 411.600 374.400 ;
        RECT 409.200 373.700 411.600 374.300 ;
        RECT 409.200 373.600 410.000 373.700 ;
        RECT 410.800 373.600 411.600 373.700 ;
        RECT 398.000 371.600 398.800 371.800 ;
        RECT 406.000 371.700 408.400 372.300 ;
        RECT 406.000 371.600 406.800 371.700 ;
        RECT 390.200 371.400 391.000 371.600 ;
        RECT 386.800 370.800 391.000 371.400 ;
        RECT 386.800 362.200 387.600 370.800 ;
        RECT 393.400 370.400 394.000 371.600 ;
        RECT 399.600 371.000 405.200 371.200 ;
        RECT 399.400 370.800 405.200 371.000 ;
        RECT 391.600 369.800 394.000 370.400 ;
        RECT 395.400 370.600 405.200 370.800 ;
        RECT 395.400 370.200 400.200 370.600 ;
        RECT 391.600 368.800 392.200 369.800 ;
        RECT 390.800 368.000 392.200 368.800 ;
        RECT 393.800 369.000 394.600 369.200 ;
        RECT 395.400 369.000 396.000 370.200 ;
        RECT 393.800 368.400 396.000 369.000 ;
        RECT 396.600 369.000 402.000 369.600 ;
        RECT 396.600 368.800 397.400 369.000 ;
        RECT 401.200 368.800 402.000 369.000 ;
        RECT 395.000 367.400 395.800 367.600 ;
        RECT 397.800 367.400 398.600 367.600 ;
        RECT 391.600 366.200 392.400 367.000 ;
        RECT 395.000 366.800 398.600 367.400 ;
        RECT 395.800 366.200 396.400 366.800 ;
        RECT 401.200 366.200 402.000 367.000 ;
        RECT 391.000 362.200 392.200 366.200 ;
        RECT 395.600 362.200 396.400 366.200 ;
        RECT 400.000 365.600 402.000 366.200 ;
        RECT 400.000 362.200 400.800 365.600 ;
        RECT 404.400 362.200 405.200 370.600 ;
        RECT 407.600 362.200 408.400 371.700 ;
        RECT 412.200 370.800 413.000 375.200 ;
        RECT 414.000 374.600 414.800 379.800 ;
        RECT 420.400 376.600 421.200 379.800 ;
        RECT 422.000 377.000 422.800 379.800 ;
        RECT 423.600 377.000 424.400 379.800 ;
        RECT 425.200 377.000 426.000 379.800 ;
        RECT 426.800 377.000 427.600 379.800 ;
        RECT 430.000 377.000 430.800 379.800 ;
        RECT 433.200 377.000 434.000 379.800 ;
        RECT 434.800 377.000 435.600 379.800 ;
        RECT 436.400 377.000 437.200 379.800 ;
        RECT 418.800 375.800 421.200 376.600 ;
        RECT 438.000 376.600 438.800 379.800 ;
        RECT 418.800 375.200 419.600 375.800 ;
        RECT 413.600 374.000 414.800 374.600 ;
        RECT 417.800 374.600 419.600 375.200 ;
        RECT 423.600 375.600 424.600 376.400 ;
        RECT 427.600 375.600 429.200 376.400 ;
        RECT 430.000 375.800 434.600 376.400 ;
        RECT 438.000 375.800 440.600 376.600 ;
        RECT 430.000 375.600 430.800 375.800 ;
        RECT 413.600 372.000 414.200 374.000 ;
        RECT 417.800 373.400 418.600 374.600 ;
        RECT 414.800 372.600 418.600 373.400 ;
        RECT 423.600 372.800 424.400 375.600 ;
        RECT 430.000 374.800 430.800 375.000 ;
        RECT 426.400 374.200 430.800 374.800 ;
        RECT 426.400 374.000 427.200 374.200 ;
        RECT 433.800 373.400 434.600 375.800 ;
        RECT 439.800 375.200 440.600 375.800 ;
        RECT 439.800 374.400 442.800 375.200 ;
        RECT 444.400 373.800 445.200 379.800 ;
        RECT 426.800 372.600 430.000 373.400 ;
        RECT 433.800 372.600 435.800 373.400 ;
        RECT 436.400 373.000 445.200 373.800 ;
        RECT 420.400 372.000 421.200 372.600 ;
        RECT 438.000 372.000 438.800 372.400 ;
        RECT 441.200 372.000 442.000 372.400 ;
        RECT 443.000 372.000 443.800 372.200 ;
        RECT 413.600 371.400 414.400 372.000 ;
        RECT 420.400 371.400 443.800 372.000 ;
        RECT 412.200 370.000 413.200 370.800 ;
        RECT 412.400 362.200 413.200 370.000 ;
        RECT 413.800 369.600 414.400 371.400 ;
        RECT 415.000 370.800 415.800 371.000 ;
        RECT 415.000 370.200 442.000 370.800 ;
        RECT 437.800 370.000 438.800 370.200 ;
        RECT 441.200 369.600 442.000 370.200 ;
        RECT 413.800 369.000 422.800 369.600 ;
        RECT 413.800 367.400 414.400 369.000 ;
        RECT 422.000 368.800 422.800 369.000 ;
        RECT 425.200 369.000 433.800 369.600 ;
        RECT 425.200 368.800 426.000 369.000 ;
        RECT 417.000 367.600 419.600 368.400 ;
        RECT 413.800 366.800 416.400 367.400 ;
        RECT 415.600 362.200 416.400 366.800 ;
        RECT 418.800 362.200 419.600 367.600 ;
        RECT 420.200 366.800 424.400 367.600 ;
        RECT 422.000 362.200 422.800 365.000 ;
        RECT 423.600 362.200 424.400 365.000 ;
        RECT 425.200 362.200 426.000 365.000 ;
        RECT 426.800 362.200 427.600 368.400 ;
        RECT 430.000 367.600 432.600 368.400 ;
        RECT 433.200 368.200 433.800 369.000 ;
        RECT 434.800 369.400 435.600 369.600 ;
        RECT 434.800 369.000 440.200 369.400 ;
        RECT 434.800 368.800 441.000 369.000 ;
        RECT 439.600 368.200 441.000 368.800 ;
        RECT 433.200 367.600 439.000 368.200 ;
        RECT 442.000 368.000 443.600 368.800 ;
        RECT 442.000 367.600 442.600 368.000 ;
        RECT 430.000 362.200 430.800 367.000 ;
        RECT 433.200 362.200 434.000 367.000 ;
        RECT 438.400 366.800 442.600 367.600 ;
        RECT 444.400 367.400 445.200 373.000 ;
        RECT 450.800 375.800 451.600 379.800 ;
        RECT 454.000 377.800 454.800 379.800 ;
        RECT 450.800 372.400 451.400 375.800 ;
        RECT 454.000 375.600 454.600 377.800 ;
        RECT 455.600 375.600 456.400 377.200 ;
        RECT 458.800 376.000 459.600 379.800 ;
        RECT 452.200 375.000 454.600 375.600 ;
        RECT 458.600 375.200 459.600 376.000 ;
        RECT 446.000 372.300 446.800 372.400 ;
        RECT 450.800 372.300 451.600 372.400 ;
        RECT 446.000 371.700 451.600 372.300 ;
        RECT 446.000 371.600 446.800 371.700 ;
        RECT 450.800 371.600 451.600 371.700 ;
        RECT 452.200 372.000 452.800 375.000 ;
        RECT 450.800 370.200 451.400 371.600 ;
        RECT 452.200 371.400 453.000 372.000 ;
        RECT 452.200 371.200 456.400 371.400 ;
        RECT 452.400 370.800 456.400 371.200 ;
        RECT 450.800 369.600 452.200 370.200 ;
        RECT 443.200 366.800 445.200 367.400 ;
        RECT 434.800 362.200 435.600 365.000 ;
        RECT 436.400 362.200 437.200 365.000 ;
        RECT 439.600 362.200 440.400 366.800 ;
        RECT 443.200 366.200 443.800 366.800 ;
        RECT 442.800 365.600 443.800 366.200 ;
        RECT 442.800 362.200 443.600 365.600 ;
        RECT 451.400 362.200 452.200 369.600 ;
        RECT 455.600 362.200 456.400 370.800 ;
        RECT 458.600 370.800 459.400 375.200 ;
        RECT 460.400 374.600 461.200 379.800 ;
        RECT 466.800 376.600 467.600 379.800 ;
        RECT 468.400 377.000 469.200 379.800 ;
        RECT 470.000 377.000 470.800 379.800 ;
        RECT 471.600 377.000 472.400 379.800 ;
        RECT 473.200 377.000 474.000 379.800 ;
        RECT 476.400 377.000 477.200 379.800 ;
        RECT 479.600 377.000 480.400 379.800 ;
        RECT 481.200 377.000 482.000 379.800 ;
        RECT 482.800 377.000 483.600 379.800 ;
        RECT 465.200 375.800 467.600 376.600 ;
        RECT 484.400 376.600 485.200 379.800 ;
        RECT 465.200 375.200 466.000 375.800 ;
        RECT 460.000 374.000 461.200 374.600 ;
        RECT 464.200 374.600 466.000 375.200 ;
        RECT 470.000 375.600 471.000 376.400 ;
        RECT 474.000 375.600 475.600 376.400 ;
        RECT 476.400 375.800 481.000 376.400 ;
        RECT 484.400 375.800 487.000 376.600 ;
        RECT 476.400 375.600 477.200 375.800 ;
        RECT 460.000 372.000 460.600 374.000 ;
        RECT 464.200 373.400 465.000 374.600 ;
        RECT 461.200 372.600 465.000 373.400 ;
        RECT 470.000 372.800 470.800 375.600 ;
        RECT 476.400 374.800 477.200 375.000 ;
        RECT 472.800 374.200 477.200 374.800 ;
        RECT 472.800 374.000 473.600 374.200 ;
        RECT 480.200 373.400 481.000 375.800 ;
        RECT 486.200 375.200 487.000 375.800 ;
        RECT 486.200 374.400 489.200 375.200 ;
        RECT 490.800 373.800 491.600 379.800 ;
        RECT 473.200 372.600 476.400 373.400 ;
        RECT 480.200 372.600 482.200 373.400 ;
        RECT 482.800 373.000 491.600 373.800 ;
        RECT 466.800 372.000 467.600 372.600 ;
        RECT 484.400 372.000 485.200 372.400 ;
        RECT 487.600 372.000 488.400 372.400 ;
        RECT 489.400 372.000 490.200 372.200 ;
        RECT 460.000 371.400 460.800 372.000 ;
        RECT 466.800 371.400 490.200 372.000 ;
        RECT 458.600 370.000 459.600 370.800 ;
        RECT 458.800 362.200 459.600 370.000 ;
        RECT 460.200 369.600 460.800 371.400 ;
        RECT 461.400 370.800 462.200 371.000 ;
        RECT 461.400 370.300 488.400 370.800 ;
        RECT 489.200 370.300 490.000 370.400 ;
        RECT 461.400 370.200 490.000 370.300 ;
        RECT 484.200 370.000 485.000 370.200 ;
        RECT 487.600 369.700 490.000 370.200 ;
        RECT 487.600 369.600 488.400 369.700 ;
        RECT 489.200 369.600 490.000 369.700 ;
        RECT 460.200 369.000 469.200 369.600 ;
        RECT 460.200 367.400 460.800 369.000 ;
        RECT 468.400 368.800 469.200 369.000 ;
        RECT 471.600 369.000 480.200 369.600 ;
        RECT 471.600 368.800 472.400 369.000 ;
        RECT 463.400 367.600 466.000 368.400 ;
        RECT 460.200 366.800 462.800 367.400 ;
        RECT 462.000 362.200 462.800 366.800 ;
        RECT 465.200 362.200 466.000 367.600 ;
        RECT 466.600 366.800 470.800 367.600 ;
        RECT 468.400 362.200 469.200 365.000 ;
        RECT 470.000 362.200 470.800 365.000 ;
        RECT 471.600 362.200 472.400 365.000 ;
        RECT 473.200 362.200 474.000 368.400 ;
        RECT 476.400 367.600 479.000 368.400 ;
        RECT 479.600 368.200 480.200 369.000 ;
        RECT 481.200 369.400 482.000 369.600 ;
        RECT 481.200 369.000 486.600 369.400 ;
        RECT 481.200 368.800 487.400 369.000 ;
        RECT 486.000 368.200 487.400 368.800 ;
        RECT 479.600 367.600 485.400 368.200 ;
        RECT 488.400 368.000 490.000 368.800 ;
        RECT 488.400 367.600 489.000 368.000 ;
        RECT 476.400 362.200 477.200 367.000 ;
        RECT 479.600 362.200 480.400 367.000 ;
        RECT 484.800 366.800 489.000 367.600 ;
        RECT 490.800 367.400 491.600 373.000 ;
        RECT 492.400 375.800 493.200 379.800 ;
        RECT 495.600 377.800 496.400 379.800 ;
        RECT 492.400 372.400 493.000 375.800 ;
        RECT 495.600 375.600 496.200 377.800 ;
        RECT 497.200 375.600 498.000 377.200 ;
        RECT 493.800 375.000 496.200 375.600 ;
        RECT 492.400 371.600 493.200 372.400 ;
        RECT 493.800 372.000 494.400 375.000 ;
        RECT 498.800 373.800 499.600 379.800 ;
        RECT 505.200 376.600 506.000 379.800 ;
        RECT 506.800 377.000 507.600 379.800 ;
        RECT 508.400 377.000 509.200 379.800 ;
        RECT 510.000 377.000 510.800 379.800 ;
        RECT 513.200 377.000 514.000 379.800 ;
        RECT 516.400 377.000 517.200 379.800 ;
        RECT 518.000 377.000 518.800 379.800 ;
        RECT 519.600 377.000 520.400 379.800 ;
        RECT 521.200 377.000 522.000 379.800 ;
        RECT 503.400 375.800 506.000 376.600 ;
        RECT 522.800 376.600 523.600 379.800 ;
        RECT 509.400 375.800 514.000 376.400 ;
        RECT 503.400 375.200 504.200 375.800 ;
        RECT 501.200 374.400 504.200 375.200 ;
        RECT 498.800 373.000 507.600 373.800 ;
        RECT 509.400 373.400 510.200 375.800 ;
        RECT 513.200 375.600 514.000 375.800 ;
        RECT 514.800 375.600 516.400 376.400 ;
        RECT 519.400 375.600 520.400 376.400 ;
        RECT 522.800 375.800 525.200 376.600 ;
        RECT 513.200 374.800 514.000 375.000 ;
        RECT 513.200 374.200 517.600 374.800 ;
        RECT 516.800 374.000 517.600 374.200 ;
        RECT 492.400 370.200 493.000 371.600 ;
        RECT 493.800 371.400 494.600 372.000 ;
        RECT 493.800 371.200 498.000 371.400 ;
        RECT 494.000 370.800 498.000 371.200 ;
        RECT 492.400 369.600 493.800 370.200 ;
        RECT 489.600 366.800 491.600 367.400 ;
        RECT 481.200 362.200 482.000 365.000 ;
        RECT 482.800 362.200 483.600 365.000 ;
        RECT 486.000 362.200 486.800 366.800 ;
        RECT 489.600 366.200 490.200 366.800 ;
        RECT 489.200 365.600 490.200 366.200 ;
        RECT 489.200 362.200 490.000 365.600 ;
        RECT 493.000 362.200 493.800 369.600 ;
        RECT 497.200 362.200 498.000 370.800 ;
        RECT 498.800 367.400 499.600 373.000 ;
        RECT 508.200 372.600 510.200 373.400 ;
        RECT 514.000 372.600 517.200 373.400 ;
        RECT 519.600 372.800 520.400 375.600 ;
        RECT 524.400 375.200 525.200 375.800 ;
        RECT 524.400 374.600 526.200 375.200 ;
        RECT 525.400 373.400 526.200 374.600 ;
        RECT 529.200 374.600 530.000 379.800 ;
        RECT 530.800 376.000 531.600 379.800 ;
        RECT 530.800 375.200 531.800 376.000 ;
        RECT 529.200 374.000 530.400 374.600 ;
        RECT 525.400 372.600 529.200 373.400 ;
        RECT 500.200 372.000 501.000 372.200 ;
        RECT 502.000 372.000 502.800 372.400 ;
        RECT 505.200 372.000 506.000 372.400 ;
        RECT 522.800 372.000 523.600 372.600 ;
        RECT 529.800 372.000 530.400 374.000 ;
        RECT 500.200 371.400 523.600 372.000 ;
        RECT 529.600 371.400 530.400 372.000 ;
        RECT 529.600 369.600 530.200 371.400 ;
        RECT 531.000 370.800 531.800 375.200 ;
        RECT 535.600 375.200 536.400 379.800 ;
        RECT 538.800 375.200 539.600 379.800 ;
        RECT 535.600 374.400 539.600 375.200 ;
        RECT 542.000 375.200 542.800 379.800 ;
        RECT 545.200 376.400 546.000 379.800 ;
        RECT 545.200 375.800 546.200 376.400 ;
        RECT 542.000 374.600 544.600 375.200 ;
        RECT 538.800 371.600 539.600 374.400 ;
        RECT 542.200 372.400 543.000 373.200 ;
        RECT 542.000 371.600 543.000 372.400 ;
        RECT 544.000 373.000 544.600 374.600 ;
        RECT 545.600 374.400 546.200 375.800 ;
        RECT 545.200 374.300 546.200 374.400 ;
        RECT 546.800 374.300 547.600 374.400 ;
        RECT 545.200 373.700 547.600 374.300 ;
        RECT 545.200 373.600 546.200 373.700 ;
        RECT 546.800 373.600 547.600 373.700 ;
        RECT 548.400 373.800 549.200 379.800 ;
        RECT 554.800 376.600 555.600 379.800 ;
        RECT 556.400 377.000 557.200 379.800 ;
        RECT 558.000 377.000 558.800 379.800 ;
        RECT 559.600 377.000 560.400 379.800 ;
        RECT 562.800 377.000 563.600 379.800 ;
        RECT 566.000 377.000 566.800 379.800 ;
        RECT 567.600 377.000 568.400 379.800 ;
        RECT 569.200 377.000 570.000 379.800 ;
        RECT 570.800 377.000 571.600 379.800 ;
        RECT 553.000 375.800 555.600 376.600 ;
        RECT 572.400 376.600 573.200 379.800 ;
        RECT 559.000 375.800 563.600 376.400 ;
        RECT 553.000 375.200 553.800 375.800 ;
        RECT 550.800 374.400 553.800 375.200 ;
        RECT 544.000 372.200 545.000 373.000 ;
        RECT 508.400 369.400 509.200 369.600 ;
        RECT 503.800 369.000 509.200 369.400 ;
        RECT 503.000 368.800 509.200 369.000 ;
        RECT 510.200 369.000 518.800 369.600 ;
        RECT 500.400 368.000 502.000 368.800 ;
        RECT 503.000 368.200 504.400 368.800 ;
        RECT 510.200 368.200 510.800 369.000 ;
        RECT 518.000 368.800 518.800 369.000 ;
        RECT 521.200 369.000 530.200 369.600 ;
        RECT 521.200 368.800 522.000 369.000 ;
        RECT 501.400 367.600 502.000 368.000 ;
        RECT 505.000 367.600 510.800 368.200 ;
        RECT 511.400 367.600 514.000 368.400 ;
        RECT 498.800 366.800 500.800 367.400 ;
        RECT 501.400 366.800 505.600 367.600 ;
        RECT 500.200 366.200 500.800 366.800 ;
        RECT 500.200 365.600 501.200 366.200 ;
        RECT 500.400 362.200 501.200 365.600 ;
        RECT 503.600 362.200 504.400 366.800 ;
        RECT 506.800 362.200 507.600 365.000 ;
        RECT 508.400 362.200 509.200 365.000 ;
        RECT 510.000 362.200 510.800 367.000 ;
        RECT 513.200 362.200 514.000 367.000 ;
        RECT 516.400 362.200 517.200 368.400 ;
        RECT 524.400 367.600 527.000 368.400 ;
        RECT 519.600 366.800 523.800 367.600 ;
        RECT 518.000 362.200 518.800 365.000 ;
        RECT 519.600 362.200 520.400 365.000 ;
        RECT 521.200 362.200 522.000 365.000 ;
        RECT 524.400 362.200 525.200 367.600 ;
        RECT 529.600 367.400 530.200 369.000 ;
        RECT 527.600 366.800 530.200 367.400 ;
        RECT 530.800 370.000 531.800 370.800 ;
        RECT 535.600 370.800 539.600 371.600 ;
        RECT 527.600 362.200 528.400 366.800 ;
        RECT 530.800 362.200 531.600 370.000 ;
        RECT 535.600 362.200 536.400 370.800 ;
        RECT 538.800 362.200 539.600 370.800 ;
        RECT 544.000 370.200 544.600 372.200 ;
        RECT 545.600 370.200 546.200 373.600 ;
        RECT 542.000 369.600 544.600 370.200 ;
        RECT 542.000 362.200 542.800 369.600 ;
        RECT 545.200 369.200 546.200 370.200 ;
        RECT 548.400 373.000 557.200 373.800 ;
        RECT 559.000 373.400 559.800 375.800 ;
        RECT 562.800 375.600 563.600 375.800 ;
        RECT 564.400 375.600 566.000 376.400 ;
        RECT 569.000 375.600 570.000 376.400 ;
        RECT 572.400 375.800 574.800 376.600 ;
        RECT 561.200 373.600 562.000 375.200 ;
        RECT 562.800 374.800 563.600 375.000 ;
        RECT 562.800 374.200 567.200 374.800 ;
        RECT 566.400 374.000 567.200 374.200 ;
        RECT 545.200 362.200 546.000 369.200 ;
        RECT 548.400 367.400 549.200 373.000 ;
        RECT 557.800 372.600 559.800 373.400 ;
        RECT 563.600 372.600 566.800 373.400 ;
        RECT 569.200 372.800 570.000 375.600 ;
        RECT 574.000 375.200 574.800 375.800 ;
        RECT 574.000 374.600 575.800 375.200 ;
        RECT 575.000 373.400 575.800 374.600 ;
        RECT 578.800 374.600 579.600 379.800 ;
        RECT 580.400 376.000 581.200 379.800 ;
        RECT 580.400 375.200 581.400 376.000 ;
        RECT 578.800 374.000 580.000 374.600 ;
        RECT 575.000 372.600 578.800 373.400 ;
        RECT 549.800 372.000 550.600 372.200 ;
        RECT 551.600 372.000 552.400 372.400 ;
        RECT 554.800 372.000 555.600 372.400 ;
        RECT 572.400 372.000 573.200 372.600 ;
        RECT 579.400 372.000 580.000 374.000 ;
        RECT 549.800 371.400 573.200 372.000 ;
        RECT 579.200 371.400 580.000 372.000 ;
        RECT 579.200 369.600 579.800 371.400 ;
        RECT 580.600 370.800 581.400 375.200 ;
        RECT 558.000 369.400 558.800 369.600 ;
        RECT 553.400 369.000 558.800 369.400 ;
        RECT 552.600 368.800 558.800 369.000 ;
        RECT 559.800 369.000 568.400 369.600 ;
        RECT 550.000 368.000 551.600 368.800 ;
        RECT 552.600 368.200 554.000 368.800 ;
        RECT 559.800 368.200 560.400 369.000 ;
        RECT 567.600 368.800 568.400 369.000 ;
        RECT 570.800 369.000 579.800 369.600 ;
        RECT 570.800 368.800 571.600 369.000 ;
        RECT 551.000 367.600 551.600 368.000 ;
        RECT 554.600 367.600 560.400 368.200 ;
        RECT 561.000 367.600 563.600 368.400 ;
        RECT 548.400 366.800 550.400 367.400 ;
        RECT 551.000 366.800 555.200 367.600 ;
        RECT 549.800 366.200 550.400 366.800 ;
        RECT 549.800 365.600 550.800 366.200 ;
        RECT 550.000 362.200 550.800 365.600 ;
        RECT 553.200 362.200 554.000 366.800 ;
        RECT 556.400 362.200 557.200 365.000 ;
        RECT 558.000 362.200 558.800 365.000 ;
        RECT 559.600 362.200 560.400 367.000 ;
        RECT 562.800 362.200 563.600 367.000 ;
        RECT 566.000 362.200 566.800 368.400 ;
        RECT 574.000 367.600 576.600 368.400 ;
        RECT 569.200 366.800 573.400 367.600 ;
        RECT 567.600 362.200 568.400 365.000 ;
        RECT 569.200 362.200 570.000 365.000 ;
        RECT 570.800 362.200 571.600 365.000 ;
        RECT 574.000 362.200 574.800 367.600 ;
        RECT 579.200 367.400 579.800 369.000 ;
        RECT 577.200 366.800 579.800 367.400 ;
        RECT 580.400 370.000 581.400 370.800 ;
        RECT 577.200 362.200 578.000 366.800 ;
        RECT 580.400 362.200 581.200 370.000 ;
        RECT 2.000 353.600 2.800 354.400 ;
        RECT 2.000 352.400 2.600 353.600 ;
        RECT 3.400 352.400 4.200 359.800 ;
        RECT 7.600 352.400 8.400 359.800 ;
        RECT 9.000 352.400 9.800 352.600 ;
        RECT 1.200 351.800 2.600 352.400 ;
        RECT 1.200 351.600 2.000 351.800 ;
        RECT 3.200 351.600 5.200 352.400 ;
        RECT 7.600 351.800 9.800 352.400 ;
        RECT 12.000 352.400 13.600 359.800 ;
        RECT 15.600 352.400 16.400 352.600 ;
        RECT 17.200 352.400 18.000 359.800 ;
        RECT 12.000 351.800 14.000 352.400 ;
        RECT 15.600 351.800 18.000 352.400 ;
        RECT 3.200 348.400 3.800 351.600 ;
        RECT 9.200 351.200 9.800 351.800 ;
        RECT 9.200 350.600 12.600 351.200 ;
        RECT 11.800 350.400 12.600 350.600 ;
        RECT 13.400 350.400 14.000 351.800 ;
        RECT 4.400 348.800 5.200 350.400 ;
        RECT 6.000 350.300 6.800 350.400 ;
        RECT 6.000 349.700 8.300 350.300 ;
        RECT 6.000 349.600 6.800 349.700 ;
        RECT 7.700 348.400 8.300 349.700 ;
        RECT 9.600 349.800 10.400 350.000 ;
        RECT 13.400 349.800 14.800 350.400 ;
        RECT 9.600 349.200 12.200 349.800 ;
        RECT 11.600 348.600 12.200 349.200 ;
        RECT 13.000 349.600 14.800 349.800 ;
        RECT 13.000 349.200 14.000 349.600 ;
        RECT 1.200 347.600 3.800 348.400 ;
        RECT 6.000 348.200 6.800 348.400 ;
        RECT 5.200 347.600 6.800 348.200 ;
        RECT 7.600 348.200 9.200 348.400 ;
        RECT 7.600 347.600 11.000 348.200 ;
        RECT 11.600 347.800 12.400 348.600 ;
        RECT 1.400 346.200 2.000 347.600 ;
        RECT 5.200 347.200 6.000 347.600 ;
        RECT 10.400 347.200 11.000 347.600 ;
        RECT 9.000 346.800 9.800 347.000 ;
        RECT 3.000 346.200 6.600 346.600 ;
        RECT 7.600 346.200 9.800 346.800 ;
        RECT 10.400 346.600 12.400 347.200 ;
        RECT 10.800 346.400 12.400 346.600 ;
        RECT 1.200 342.200 2.000 346.200 ;
        RECT 2.800 346.000 6.800 346.200 ;
        RECT 2.800 342.200 3.600 346.000 ;
        RECT 6.000 342.200 6.800 346.000 ;
        RECT 7.600 342.200 8.400 346.200 ;
        RECT 13.000 345.800 13.600 349.200 ;
        RECT 14.400 347.600 15.200 348.400 ;
        RECT 16.400 347.600 18.000 348.400 ;
        RECT 14.400 347.200 15.000 347.600 ;
        RECT 14.200 346.400 15.000 347.200 ;
        RECT 15.600 346.800 16.400 347.000 ;
        RECT 15.600 346.200 18.000 346.800 ;
        RECT 12.000 342.200 13.600 345.800 ;
        RECT 17.200 342.200 18.000 346.200 ;
        RECT 18.800 344.800 19.600 346.400 ;
        RECT 20.400 342.200 21.200 359.800 ;
        RECT 22.000 352.400 22.800 359.800 ;
        RECT 23.400 352.400 24.200 352.600 ;
        RECT 22.000 351.800 24.200 352.400 ;
        RECT 26.400 352.400 28.000 359.800 ;
        RECT 30.000 352.400 30.800 352.600 ;
        RECT 31.600 352.400 32.400 359.800 ;
        RECT 26.400 351.800 29.200 352.400 ;
        RECT 30.000 351.800 32.400 352.400 ;
        RECT 23.600 351.200 24.200 351.800 ;
        RECT 27.800 351.600 29.200 351.800 ;
        RECT 23.600 350.600 27.000 351.200 ;
        RECT 26.200 350.400 27.000 350.600 ;
        RECT 27.800 350.400 28.400 351.600 ;
        RECT 24.000 349.800 24.800 350.000 ;
        RECT 27.800 349.800 29.200 350.400 ;
        RECT 24.000 349.200 26.600 349.800 ;
        RECT 26.000 348.600 26.600 349.200 ;
        RECT 27.400 349.600 29.200 349.800 ;
        RECT 27.400 349.200 28.400 349.600 ;
        RECT 22.000 348.200 23.600 348.400 ;
        RECT 22.000 347.600 25.400 348.200 ;
        RECT 26.000 347.800 26.800 348.600 ;
        RECT 24.800 347.200 25.400 347.600 ;
        RECT 23.400 346.800 24.200 347.000 ;
        RECT 22.000 346.200 24.200 346.800 ;
        RECT 24.800 346.600 26.800 347.200 ;
        RECT 25.200 346.400 26.800 346.600 ;
        RECT 22.000 342.200 22.800 346.200 ;
        RECT 27.400 345.800 28.000 349.200 ;
        RECT 28.800 347.600 29.600 348.400 ;
        RECT 30.800 348.300 32.400 348.400 ;
        RECT 33.200 348.300 34.000 348.400 ;
        RECT 30.800 347.700 34.000 348.300 ;
        RECT 30.800 347.600 32.400 347.700 ;
        RECT 33.200 347.600 34.000 347.700 ;
        RECT 28.800 347.200 29.400 347.600 ;
        RECT 28.600 346.400 29.400 347.200 ;
        RECT 30.000 346.800 30.800 347.000 ;
        RECT 30.000 346.200 32.400 346.800 ;
        RECT 26.400 344.400 28.000 345.800 ;
        RECT 25.200 343.600 28.000 344.400 ;
        RECT 26.400 342.200 28.000 343.600 ;
        RECT 31.600 342.200 32.400 346.200 ;
        RECT 33.200 344.800 34.000 346.400 ;
        RECT 34.800 342.200 35.600 359.800 ;
        RECT 36.400 351.200 37.200 359.800 ;
        RECT 40.600 352.400 41.400 359.800 ;
        RECT 40.600 351.800 42.000 352.400 ;
        RECT 42.800 351.800 43.600 359.800 ;
        RECT 44.400 352.400 45.200 359.800 ;
        RECT 47.600 352.400 48.400 359.800 ;
        RECT 50.000 353.600 50.800 354.400 ;
        RECT 50.000 352.400 50.600 353.600 ;
        RECT 51.400 352.400 52.200 359.800 ;
        RECT 44.400 351.800 48.400 352.400 ;
        RECT 49.200 351.800 50.600 352.400 ;
        RECT 51.200 351.800 52.200 352.400 ;
        RECT 58.200 352.400 59.000 359.800 ;
        RECT 59.600 353.600 60.400 354.400 ;
        RECT 59.800 352.400 60.400 353.600 ;
        RECT 62.000 352.400 62.800 359.800 ;
        RECT 65.200 352.400 66.000 359.800 ;
        RECT 58.200 351.800 59.200 352.400 ;
        RECT 59.800 351.800 61.200 352.400 ;
        RECT 62.000 351.800 66.000 352.400 ;
        RECT 66.800 351.800 67.600 359.800 ;
        RECT 69.000 352.600 69.800 359.800 ;
        RECT 75.800 352.600 76.600 359.800 ;
        RECT 69.000 351.800 70.800 352.600 ;
        RECT 74.800 351.800 76.600 352.600 ;
        RECT 78.000 352.400 78.800 359.800 ;
        RECT 81.200 352.400 82.000 359.800 ;
        RECT 78.000 351.800 82.000 352.400 ;
        RECT 82.800 351.800 83.600 359.800 ;
        RECT 87.000 352.600 87.800 359.800 ;
        RECT 86.000 351.800 87.800 352.600 ;
        RECT 36.400 350.800 40.400 351.200 ;
        RECT 36.400 350.600 40.600 350.800 ;
        RECT 39.800 350.000 40.600 350.600 ;
        RECT 41.400 350.400 42.000 351.800 ;
        RECT 43.000 350.400 43.600 351.800 ;
        RECT 49.200 351.600 50.000 351.800 ;
        RECT 46.800 350.400 47.600 350.800 ;
        RECT 38.400 348.400 39.200 349.200 ;
        RECT 38.000 347.600 39.000 348.400 ;
        RECT 40.000 347.000 40.600 350.000 ;
        RECT 41.200 349.600 42.000 350.400 ;
        RECT 42.800 349.800 45.200 350.400 ;
        RECT 46.800 349.800 48.400 350.400 ;
        RECT 42.800 349.600 43.600 349.800 ;
        RECT 38.200 346.400 40.600 347.000 ;
        RECT 36.400 344.800 37.200 346.400 ;
        RECT 38.200 344.200 38.800 346.400 ;
        RECT 41.400 346.200 42.000 349.600 ;
        RECT 38.000 342.200 38.800 344.200 ;
        RECT 41.200 342.200 42.000 346.200 ;
        RECT 42.800 345.600 43.600 346.400 ;
        RECT 44.600 346.200 45.200 349.800 ;
        RECT 47.600 349.600 48.400 349.800 ;
        RECT 46.000 347.600 46.800 349.200 ;
        RECT 51.200 348.400 51.800 351.800 ;
        RECT 52.400 348.800 53.200 350.400 ;
        RECT 57.200 348.800 58.000 350.400 ;
        RECT 58.600 348.400 59.200 351.800 ;
        RECT 60.400 351.600 61.200 351.800 ;
        RECT 62.800 350.400 63.600 350.800 ;
        RECT 66.800 350.400 67.400 351.800 ;
        RECT 62.000 349.800 63.600 350.400 ;
        RECT 65.200 349.800 67.600 350.400 ;
        RECT 62.000 349.600 62.800 349.800 ;
        RECT 65.200 349.600 66.000 349.800 ;
        RECT 66.800 349.600 67.600 349.800 ;
        RECT 68.400 349.600 69.200 351.200 ;
        RECT 49.200 347.600 51.800 348.400 ;
        RECT 54.000 348.200 54.800 348.400 ;
        RECT 53.200 347.600 54.800 348.200 ;
        RECT 55.600 348.200 56.400 348.400 ;
        RECT 58.600 348.300 61.200 348.400 ;
        RECT 62.000 348.300 62.800 348.400 ;
        RECT 55.600 347.600 57.200 348.200 ;
        RECT 58.600 347.700 62.800 348.300 ;
        RECT 58.600 347.600 61.200 347.700 ;
        RECT 62.000 347.600 62.800 347.700 ;
        RECT 63.600 347.600 64.400 349.200 ;
        RECT 49.400 346.200 50.000 347.600 ;
        RECT 53.200 347.200 54.000 347.600 ;
        RECT 56.400 347.200 57.200 347.600 ;
        RECT 51.000 346.200 54.600 346.600 ;
        RECT 55.800 346.200 59.400 346.600 ;
        RECT 60.400 346.200 61.000 347.600 ;
        RECT 65.200 346.200 65.800 349.600 ;
        RECT 70.000 348.400 70.600 351.800 ;
        RECT 75.000 348.400 75.600 351.800 ;
        RECT 76.400 349.600 77.200 351.200 ;
        RECT 78.800 350.400 79.600 350.800 ;
        RECT 82.800 350.400 83.400 351.800 ;
        RECT 78.000 349.800 79.600 350.400 ;
        RECT 81.200 349.800 83.600 350.400 ;
        RECT 78.000 349.600 78.800 349.800 ;
        RECT 70.000 347.600 70.800 348.400 ;
        RECT 74.800 347.600 75.600 348.400 ;
        RECT 76.400 348.300 77.200 348.400 ;
        RECT 79.600 348.300 80.400 349.200 ;
        RECT 76.400 347.700 80.400 348.300 ;
        RECT 76.400 347.600 77.200 347.700 ;
        RECT 79.600 347.600 80.400 347.700 ;
        RECT 66.800 346.300 67.600 346.400 ;
        RECT 70.000 346.300 70.600 347.600 ;
        RECT 71.600 346.300 72.400 346.400 ;
        RECT 73.200 346.300 74.000 346.400 ;
        RECT 43.000 344.800 43.800 345.600 ;
        RECT 44.400 342.200 45.200 346.200 ;
        RECT 49.200 342.200 50.000 346.200 ;
        RECT 50.800 346.000 54.800 346.200 ;
        RECT 50.800 342.200 51.600 346.000 ;
        RECT 54.000 342.200 54.800 346.000 ;
        RECT 55.600 346.000 59.600 346.200 ;
        RECT 55.600 342.200 56.400 346.000 ;
        RECT 58.800 342.200 59.600 346.000 ;
        RECT 60.400 342.200 61.200 346.200 ;
        RECT 65.200 342.200 66.000 346.200 ;
        RECT 66.800 345.700 70.700 346.300 ;
        RECT 71.600 345.700 74.000 346.300 ;
        RECT 66.800 345.600 67.600 345.700 ;
        RECT 66.600 344.800 67.400 345.600 ;
        RECT 70.000 344.200 70.600 345.700 ;
        RECT 71.600 344.800 72.400 345.700 ;
        RECT 73.200 344.800 74.000 345.700 ;
        RECT 75.000 344.400 75.600 347.600 ;
        RECT 70.000 342.200 70.800 344.200 ;
        RECT 74.800 342.200 75.600 344.400 ;
        RECT 81.200 346.200 81.800 349.800 ;
        RECT 82.800 349.600 83.600 349.800 ;
        RECT 86.200 348.400 86.800 351.800 ;
        RECT 89.200 351.600 90.000 353.200 ;
        RECT 87.600 349.600 88.400 351.200 ;
        RECT 86.000 348.300 86.800 348.400 ;
        RECT 82.900 347.700 86.800 348.300 ;
        RECT 82.900 346.400 83.500 347.700 ;
        RECT 86.000 347.600 86.800 347.700 ;
        RECT 81.200 342.200 82.000 346.200 ;
        RECT 82.800 345.600 83.600 346.400 ;
        RECT 82.600 344.800 83.400 345.600 ;
        RECT 84.400 344.800 85.200 346.400 ;
        RECT 86.200 344.200 86.800 347.600 ;
        RECT 90.800 346.200 91.600 359.800 ;
        RECT 94.000 351.200 94.800 359.800 ;
        RECT 98.200 355.800 99.400 359.800 ;
        RECT 102.800 355.800 103.600 359.800 ;
        RECT 107.200 356.400 108.000 359.800 ;
        RECT 107.200 355.800 109.200 356.400 ;
        RECT 98.800 355.000 99.600 355.800 ;
        RECT 103.000 355.200 103.600 355.800 ;
        RECT 102.200 354.600 105.800 355.200 ;
        RECT 108.400 355.000 109.200 355.800 ;
        RECT 102.200 354.400 103.000 354.600 ;
        RECT 105.000 354.400 105.800 354.600 ;
        RECT 98.000 353.200 99.400 354.000 ;
        RECT 98.800 352.200 99.400 353.200 ;
        RECT 101.000 353.000 103.200 353.600 ;
        RECT 101.000 352.800 101.800 353.000 ;
        RECT 98.800 351.600 101.200 352.200 ;
        RECT 94.000 350.600 98.200 351.200 ;
        RECT 92.400 348.300 93.200 348.400 ;
        RECT 94.000 348.300 94.800 350.600 ;
        RECT 97.400 350.400 98.200 350.600 ;
        RECT 100.600 350.400 101.200 351.600 ;
        RECT 102.600 351.800 103.200 353.000 ;
        RECT 103.800 353.000 104.600 353.200 ;
        RECT 108.400 353.000 109.200 353.200 ;
        RECT 103.800 352.400 109.200 353.000 ;
        RECT 102.600 351.400 107.400 351.800 ;
        RECT 111.600 351.400 112.400 359.800 ;
        RECT 113.200 351.600 114.000 353.200 ;
        RECT 102.600 351.200 112.400 351.400 ;
        RECT 106.600 351.000 112.400 351.200 ;
        RECT 106.800 350.800 112.400 351.000 ;
        RECT 95.800 349.800 96.600 350.000 ;
        RECT 95.800 349.200 99.600 349.800 ;
        RECT 100.400 349.600 101.200 350.400 ;
        RECT 105.200 350.200 106.000 350.400 ;
        RECT 105.200 349.600 110.200 350.200 ;
        RECT 98.800 349.000 99.600 349.200 ;
        RECT 92.400 347.700 94.800 348.300 ;
        RECT 100.600 348.400 101.200 349.600 ;
        RECT 106.800 349.400 107.600 349.600 ;
        RECT 109.400 349.400 110.200 349.600 ;
        RECT 107.800 348.400 108.600 348.600 ;
        RECT 100.600 347.800 111.600 348.400 ;
        RECT 92.400 346.800 93.200 347.700 ;
        RECT 94.000 347.200 94.800 347.700 ;
        RECT 101.000 347.600 101.800 347.800 ;
        RECT 89.800 345.600 91.600 346.200 ;
        RECT 94.000 346.600 97.800 347.200 ;
        RECT 89.800 344.400 90.600 345.600 ;
        RECT 86.000 342.200 86.800 344.200 ;
        RECT 89.200 343.600 90.600 344.400 ;
        RECT 89.800 342.200 90.600 343.600 ;
        RECT 94.000 342.200 94.800 346.600 ;
        RECT 97.000 346.400 97.800 346.600 ;
        RECT 106.800 345.600 107.400 347.800 ;
        RECT 110.000 347.600 111.600 347.800 ;
        RECT 105.000 345.400 105.800 345.600 ;
        RECT 98.800 344.200 99.600 345.000 ;
        RECT 103.000 344.800 105.800 345.400 ;
        RECT 106.800 344.800 107.600 345.600 ;
        RECT 103.000 344.200 103.600 344.800 ;
        RECT 108.400 344.200 109.200 345.000 ;
        RECT 98.200 343.600 99.600 344.200 ;
        RECT 98.200 342.200 99.400 343.600 ;
        RECT 102.800 342.200 103.600 344.200 ;
        RECT 107.200 343.600 109.200 344.200 ;
        RECT 107.200 342.200 108.000 343.600 ;
        RECT 111.600 342.200 112.400 347.000 ;
        RECT 114.800 346.200 115.600 359.800 ;
        RECT 116.400 346.800 117.200 348.400 ;
        RECT 113.800 345.600 115.600 346.200 ;
        RECT 113.800 344.400 114.600 345.600 ;
        RECT 113.200 343.600 114.600 344.400 ;
        RECT 113.800 342.200 114.600 343.600 ;
        RECT 118.000 342.200 118.800 359.800 ;
        RECT 121.200 352.400 122.000 359.800 ;
        RECT 123.000 352.400 123.800 352.600 ;
        RECT 121.200 351.800 123.800 352.400 ;
        RECT 125.600 351.800 127.200 359.800 ;
        RECT 129.200 352.400 130.000 352.600 ;
        RECT 130.800 352.400 131.600 359.800 ;
        RECT 129.200 351.800 131.600 352.400 ;
        RECT 124.200 350.400 125.000 350.600 ;
        RECT 126.200 350.400 126.800 351.800 ;
        RECT 123.400 349.800 125.000 350.400 ;
        RECT 123.400 349.600 124.200 349.800 ;
        RECT 126.000 349.600 126.800 350.400 ;
        RECT 124.800 348.600 125.600 348.800 ;
        RECT 122.800 348.400 125.600 348.600 ;
        RECT 119.600 346.800 120.400 348.400 ;
        RECT 121.200 348.000 125.600 348.400 ;
        RECT 126.200 348.400 126.800 349.600 ;
        RECT 121.200 347.800 123.400 348.000 ;
        RECT 126.200 347.800 127.200 348.400 ;
        RECT 121.200 347.600 122.800 347.800 ;
        RECT 123.000 346.800 123.800 347.000 ;
        RECT 121.200 346.200 123.800 346.800 ;
        RECT 124.400 346.400 126.000 347.200 ;
        RECT 121.200 342.200 122.000 346.200 ;
        RECT 126.600 345.800 127.200 347.800 ;
        RECT 128.000 347.600 128.800 348.400 ;
        RECT 130.000 347.600 131.600 348.400 ;
        RECT 128.000 347.200 128.600 347.600 ;
        RECT 127.800 346.400 128.600 347.200 ;
        RECT 129.200 346.800 130.000 347.000 ;
        RECT 132.400 346.800 133.200 348.400 ;
        RECT 129.200 346.200 131.600 346.800 ;
        RECT 125.600 344.400 127.200 345.800 ;
        RECT 125.600 343.600 128.400 344.400 ;
        RECT 125.600 342.200 127.200 343.600 ;
        RECT 130.800 342.200 131.600 346.200 ;
        RECT 134.000 346.200 134.800 359.800 ;
        RECT 135.600 351.600 136.400 353.200 ;
        RECT 142.000 352.400 142.800 359.800 ;
        RECT 143.800 352.400 144.600 352.600 ;
        RECT 142.000 351.800 144.600 352.400 ;
        RECT 146.400 351.800 148.000 359.800 ;
        RECT 150.000 352.400 150.800 352.600 ;
        RECT 151.600 352.400 152.400 359.800 ;
        RECT 150.000 351.800 152.400 352.400 ;
        RECT 145.000 350.400 145.800 350.600 ;
        RECT 147.000 350.400 147.600 351.800 ;
        RECT 144.200 349.800 145.800 350.400 ;
        RECT 144.200 349.600 145.000 349.800 ;
        RECT 146.800 349.600 147.600 350.400 ;
        RECT 145.600 348.600 146.400 348.800 ;
        RECT 143.600 348.400 146.400 348.600 ;
        RECT 142.000 348.000 146.400 348.400 ;
        RECT 147.000 348.400 147.600 349.600 ;
        RECT 153.200 351.200 154.000 359.800 ;
        RECT 157.400 355.800 158.600 359.800 ;
        RECT 162.000 355.800 162.800 359.800 ;
        RECT 166.400 356.400 167.200 359.800 ;
        RECT 166.400 355.800 168.400 356.400 ;
        RECT 158.000 355.000 158.800 355.800 ;
        RECT 162.200 355.200 162.800 355.800 ;
        RECT 161.400 354.600 165.000 355.200 ;
        RECT 167.600 355.000 168.400 355.800 ;
        RECT 161.400 354.400 162.200 354.600 ;
        RECT 164.200 354.400 165.000 354.600 ;
        RECT 157.200 353.200 158.600 354.000 ;
        RECT 158.000 352.200 158.600 353.200 ;
        RECT 160.200 353.000 162.400 353.600 ;
        RECT 160.200 352.800 161.000 353.000 ;
        RECT 158.000 351.600 160.400 352.200 ;
        RECT 153.200 350.600 157.400 351.200 ;
        RECT 142.000 347.800 144.200 348.000 ;
        RECT 147.000 347.800 148.000 348.400 ;
        RECT 142.000 347.600 143.600 347.800 ;
        RECT 143.800 346.800 144.600 347.000 ;
        RECT 142.000 346.200 144.600 346.800 ;
        RECT 145.200 346.400 146.800 347.200 ;
        RECT 134.000 345.600 135.800 346.200 ;
        RECT 135.000 344.300 135.800 345.600 ;
        RECT 140.400 344.300 141.200 344.400 ;
        RECT 135.000 343.700 141.200 344.300 ;
        RECT 135.000 342.200 135.800 343.700 ;
        RECT 140.400 343.600 141.200 343.700 ;
        RECT 142.000 342.200 142.800 346.200 ;
        RECT 147.400 345.800 148.000 347.800 ;
        RECT 148.800 347.600 149.600 348.400 ;
        RECT 150.800 347.600 152.400 348.400 ;
        RECT 148.800 347.200 149.400 347.600 ;
        RECT 148.600 346.400 149.400 347.200 ;
        RECT 153.200 347.200 154.000 350.600 ;
        RECT 156.600 350.400 157.400 350.600 ;
        RECT 159.800 350.400 160.400 351.600 ;
        RECT 161.800 351.800 162.400 353.000 ;
        RECT 163.000 353.000 163.800 353.200 ;
        RECT 167.600 353.000 168.400 353.200 ;
        RECT 163.000 352.400 168.400 353.000 ;
        RECT 161.800 351.400 166.600 351.800 ;
        RECT 170.800 351.400 171.600 359.800 ;
        RECT 161.800 351.200 171.600 351.400 ;
        RECT 165.800 351.000 171.600 351.200 ;
        RECT 166.000 350.800 171.600 351.000 ;
        RECT 172.400 351.200 173.200 359.800 ;
        RECT 176.600 355.800 177.800 359.800 ;
        RECT 181.200 355.800 182.000 359.800 ;
        RECT 185.600 356.400 186.400 359.800 ;
        RECT 185.600 355.800 187.600 356.400 ;
        RECT 177.200 355.000 178.000 355.800 ;
        RECT 181.400 355.200 182.000 355.800 ;
        RECT 180.600 354.600 184.200 355.200 ;
        RECT 186.800 355.000 187.600 355.800 ;
        RECT 180.600 354.400 181.400 354.600 ;
        RECT 183.400 354.400 184.200 354.600 ;
        RECT 176.400 353.200 177.800 354.000 ;
        RECT 177.200 352.200 177.800 353.200 ;
        RECT 179.400 353.000 181.600 353.600 ;
        RECT 179.400 352.800 180.200 353.000 ;
        RECT 177.200 351.600 179.600 352.200 ;
        RECT 172.400 350.600 176.600 351.200 ;
        RECT 155.000 349.800 155.800 350.000 ;
        RECT 155.000 349.200 158.800 349.800 ;
        RECT 159.600 349.600 160.400 350.400 ;
        RECT 164.400 350.200 165.200 350.400 ;
        RECT 164.400 349.600 169.400 350.200 ;
        RECT 158.000 349.000 158.800 349.200 ;
        RECT 159.800 348.400 160.400 349.600 ;
        RECT 166.000 349.400 166.800 349.600 ;
        RECT 168.600 349.400 169.400 349.600 ;
        RECT 167.000 348.400 167.800 348.600 ;
        RECT 159.800 347.800 170.800 348.400 ;
        RECT 160.200 347.600 161.000 347.800 ;
        RECT 150.000 346.800 150.800 347.000 ;
        RECT 150.000 346.200 152.400 346.800 ;
        RECT 146.400 344.400 148.000 345.800 ;
        RECT 146.400 343.600 149.200 344.400 ;
        RECT 146.400 342.200 148.000 343.600 ;
        RECT 151.600 342.200 152.400 346.200 ;
        RECT 153.200 346.600 157.000 347.200 ;
        RECT 153.200 342.200 154.000 346.600 ;
        RECT 156.200 346.400 157.000 346.600 ;
        RECT 166.000 345.600 166.600 347.800 ;
        RECT 169.200 347.600 170.800 347.800 ;
        RECT 172.400 347.200 173.200 350.600 ;
        RECT 175.800 350.400 176.600 350.600 ;
        RECT 179.000 350.400 179.600 351.600 ;
        RECT 181.000 351.800 181.600 353.000 ;
        RECT 182.200 353.000 183.000 353.200 ;
        RECT 186.800 353.000 187.600 353.200 ;
        RECT 182.200 352.400 187.600 353.000 ;
        RECT 181.000 351.400 185.800 351.800 ;
        RECT 190.000 351.400 190.800 359.800 ;
        RECT 192.200 352.600 193.000 359.800 ;
        RECT 192.200 351.800 194.000 352.600 ;
        RECT 196.400 352.400 197.200 359.800 ;
        RECT 198.200 352.400 199.000 352.600 ;
        RECT 200.800 352.400 202.400 359.800 ;
        RECT 196.400 351.800 199.000 352.400 ;
        RECT 199.600 351.800 202.400 352.400 ;
        RECT 204.400 352.400 205.200 352.600 ;
        RECT 206.000 352.400 206.800 359.800 ;
        RECT 204.400 351.800 206.800 352.400 ;
        RECT 210.200 351.800 212.200 359.800 ;
        RECT 215.600 351.800 216.400 359.800 ;
        RECT 217.200 352.400 218.000 359.800 ;
        RECT 220.400 352.400 221.200 359.800 ;
        RECT 217.200 351.800 221.200 352.400 ;
        RECT 222.000 352.400 222.800 359.800 ;
        RECT 223.800 352.400 224.600 352.600 ;
        RECT 222.000 351.800 224.600 352.400 ;
        RECT 226.400 351.800 228.000 359.800 ;
        RECT 230.000 352.400 230.800 352.600 ;
        RECT 231.600 352.400 232.400 359.800 ;
        RECT 234.000 353.600 234.800 354.400 ;
        RECT 234.000 352.400 234.600 353.600 ;
        RECT 235.400 352.400 236.200 359.800 ;
        RECT 230.000 351.800 232.400 352.400 ;
        RECT 233.200 351.800 234.600 352.400 ;
        RECT 235.200 351.800 236.200 352.400 ;
        RECT 181.000 351.200 190.800 351.400 ;
        RECT 185.000 351.000 190.800 351.200 ;
        RECT 185.200 350.800 190.800 351.000 ;
        RECT 174.200 349.800 175.000 350.000 ;
        RECT 174.200 349.200 178.000 349.800 ;
        RECT 178.800 349.600 179.600 350.400 ;
        RECT 183.600 350.200 184.400 350.400 ;
        RECT 183.600 349.600 188.600 350.200 ;
        RECT 191.600 349.600 192.400 351.200 ;
        RECT 193.200 350.300 193.800 351.800 ;
        RECT 199.600 351.600 202.000 351.800 ;
        RECT 199.400 350.400 200.200 350.600 ;
        RECT 201.400 350.400 202.000 351.600 ;
        RECT 196.400 350.300 197.200 350.400 ;
        RECT 193.200 349.700 197.200 350.300 ;
        RECT 177.200 349.000 178.000 349.200 ;
        RECT 179.000 348.400 179.600 349.600 ;
        RECT 185.200 349.400 186.000 349.600 ;
        RECT 187.800 349.400 188.600 349.600 ;
        RECT 186.200 348.400 187.000 348.600 ;
        RECT 193.200 348.400 193.800 349.700 ;
        RECT 196.400 349.600 197.200 349.700 ;
        RECT 198.600 349.800 200.200 350.400 ;
        RECT 198.600 349.600 199.400 349.800 ;
        RECT 201.200 349.600 202.000 350.400 ;
        RECT 200.000 348.600 200.800 348.800 ;
        RECT 198.000 348.400 200.800 348.600 ;
        RECT 179.000 347.800 190.000 348.400 ;
        RECT 179.400 347.600 180.200 347.800 ;
        RECT 164.200 345.400 165.000 345.600 ;
        RECT 158.000 344.200 158.800 345.000 ;
        RECT 162.200 344.800 165.000 345.400 ;
        RECT 166.000 344.800 166.800 345.600 ;
        RECT 162.200 344.200 162.800 344.800 ;
        RECT 167.600 344.200 168.400 345.000 ;
        RECT 157.400 343.600 158.800 344.200 ;
        RECT 157.400 342.200 158.600 343.600 ;
        RECT 162.000 342.200 162.800 344.200 ;
        RECT 166.400 343.600 168.400 344.200 ;
        RECT 166.400 342.200 167.200 343.600 ;
        RECT 170.800 342.200 171.600 347.000 ;
        RECT 172.400 346.600 176.200 347.200 ;
        RECT 172.400 342.200 173.200 346.600 ;
        RECT 175.400 346.400 176.200 346.600 ;
        RECT 185.200 345.600 185.800 347.800 ;
        RECT 188.400 347.600 190.000 347.800 ;
        RECT 193.200 347.600 194.000 348.400 ;
        RECT 196.400 348.000 200.800 348.400 ;
        RECT 201.400 348.400 202.000 349.600 ;
        RECT 196.400 347.800 198.600 348.000 ;
        RECT 201.400 347.800 202.400 348.400 ;
        RECT 196.400 347.600 198.000 347.800 ;
        RECT 183.400 345.400 184.200 345.600 ;
        RECT 177.200 344.200 178.000 345.000 ;
        RECT 181.400 344.800 184.200 345.400 ;
        RECT 185.200 344.800 186.000 345.600 ;
        RECT 181.400 344.200 182.000 344.800 ;
        RECT 186.800 344.200 187.600 345.000 ;
        RECT 176.600 343.600 178.000 344.200 ;
        RECT 176.600 342.200 177.800 343.600 ;
        RECT 181.200 342.200 182.000 344.200 ;
        RECT 185.600 343.600 187.600 344.200 ;
        RECT 185.600 342.200 186.400 343.600 ;
        RECT 190.000 342.200 190.800 347.000 ;
        RECT 193.200 344.200 193.800 347.600 ;
        RECT 198.200 346.800 199.000 347.000 ;
        RECT 194.800 344.800 195.600 346.400 ;
        RECT 196.400 346.200 199.000 346.800 ;
        RECT 199.600 346.400 201.200 347.200 ;
        RECT 193.200 342.200 194.000 344.200 ;
        RECT 196.400 342.200 197.200 346.200 ;
        RECT 201.800 345.800 202.400 347.800 ;
        RECT 203.200 347.600 204.000 348.400 ;
        RECT 205.200 347.600 206.800 348.400 ;
        RECT 207.600 347.600 208.400 349.200 ;
        RECT 209.200 348.800 210.000 350.400 ;
        RECT 211.000 348.400 211.600 351.800 ;
        RECT 215.800 350.400 216.400 351.800 ;
        RECT 219.600 350.400 220.400 350.800 ;
        RECT 225.000 350.400 225.800 350.600 ;
        RECT 227.000 350.400 227.600 351.800 ;
        RECT 233.200 351.600 234.000 351.800 ;
        RECT 212.400 350.300 213.200 350.400 ;
        RECT 215.600 350.300 218.000 350.400 ;
        RECT 212.400 349.800 218.000 350.300 ;
        RECT 219.600 350.300 221.200 350.400 ;
        RECT 219.600 349.800 222.700 350.300 ;
        RECT 212.400 349.700 216.400 349.800 ;
        RECT 212.400 348.800 213.200 349.700 ;
        RECT 215.600 349.600 216.400 349.700 ;
        RECT 210.800 348.200 211.600 348.400 ;
        RECT 214.000 348.200 214.800 348.400 ;
        RECT 209.200 347.600 211.600 348.200 ;
        RECT 213.200 347.600 214.800 348.200 ;
        RECT 203.200 347.200 203.800 347.600 ;
        RECT 203.000 346.400 203.800 347.200 ;
        RECT 204.400 346.800 205.200 347.000 ;
        RECT 204.400 346.200 206.800 346.800 ;
        RECT 209.200 346.400 209.800 347.600 ;
        RECT 213.200 347.200 214.000 347.600 ;
        RECT 200.800 342.200 202.400 345.800 ;
        RECT 206.000 342.200 206.800 346.200 ;
        RECT 207.600 342.800 208.400 346.200 ;
        RECT 209.200 343.400 210.000 346.400 ;
        RECT 211.000 346.200 214.600 346.600 ;
        RECT 210.800 346.000 214.800 346.200 ;
        RECT 210.800 342.800 211.600 346.000 ;
        RECT 207.600 342.200 211.600 342.800 ;
        RECT 214.000 342.200 214.800 346.000 ;
        RECT 215.600 345.600 216.400 346.400 ;
        RECT 217.400 346.200 218.000 349.800 ;
        RECT 220.400 349.700 222.700 349.800 ;
        RECT 220.400 349.600 221.200 349.700 ;
        RECT 218.800 347.600 219.600 349.200 ;
        RECT 222.100 348.400 222.700 349.700 ;
        RECT 224.200 349.800 225.800 350.400 ;
        RECT 224.200 349.600 225.000 349.800 ;
        RECT 226.800 349.600 227.600 350.400 ;
        RECT 228.400 350.300 229.200 350.400 ;
        RECT 235.200 350.300 235.800 351.800 ;
        RECT 239.600 351.600 240.400 353.200 ;
        RECT 228.400 349.700 235.800 350.300 ;
        RECT 228.400 349.600 229.200 349.700 ;
        RECT 225.600 348.600 226.400 348.800 ;
        RECT 223.600 348.400 226.400 348.600 ;
        RECT 222.000 348.000 226.400 348.400 ;
        RECT 227.000 348.400 227.600 349.600 ;
        RECT 235.200 348.400 235.800 349.700 ;
        RECT 236.400 348.800 237.200 350.400 ;
        RECT 222.000 347.800 224.200 348.000 ;
        RECT 227.000 347.800 228.000 348.400 ;
        RECT 222.000 347.600 223.600 347.800 ;
        RECT 223.800 346.800 224.600 347.000 ;
        RECT 215.800 344.800 216.600 345.600 ;
        RECT 217.200 342.200 218.000 346.200 ;
        RECT 222.000 346.200 224.600 346.800 ;
        RECT 225.200 346.400 226.800 347.200 ;
        RECT 222.000 342.200 222.800 346.200 ;
        RECT 227.400 345.800 228.000 347.800 ;
        RECT 228.800 347.600 229.600 348.400 ;
        RECT 230.800 347.600 232.400 348.400 ;
        RECT 233.200 347.600 235.800 348.400 ;
        RECT 238.000 348.200 238.800 348.400 ;
        RECT 237.200 347.600 238.800 348.200 ;
        RECT 228.800 347.200 229.400 347.600 ;
        RECT 228.600 346.400 229.400 347.200 ;
        RECT 230.000 346.800 230.800 347.000 ;
        RECT 230.000 346.200 232.400 346.800 ;
        RECT 233.400 346.200 234.000 347.600 ;
        RECT 237.200 347.200 238.000 347.600 ;
        RECT 235.000 346.200 238.600 346.600 ;
        RECT 241.200 346.200 242.000 359.800 ;
        RECT 242.800 346.800 243.600 348.400 ;
        RECT 244.400 346.800 245.200 348.400 ;
        RECT 226.400 344.400 228.000 345.800 ;
        RECT 225.200 343.600 228.000 344.400 ;
        RECT 226.400 342.200 228.000 343.600 ;
        RECT 231.600 342.200 232.400 346.200 ;
        RECT 233.200 342.200 234.000 346.200 ;
        RECT 234.800 346.000 238.800 346.200 ;
        RECT 234.800 342.200 235.600 346.000 ;
        RECT 238.000 342.200 238.800 346.000 ;
        RECT 240.200 345.600 242.000 346.200 ;
        RECT 246.000 346.200 246.800 359.800 ;
        RECT 247.600 351.600 248.400 353.200 ;
        RECT 247.600 350.300 248.400 350.400 ;
        RECT 250.800 350.300 251.600 359.800 ;
        RECT 247.600 349.700 251.600 350.300 ;
        RECT 247.600 349.600 248.400 349.700 ;
        RECT 249.200 346.800 250.000 348.400 ;
        RECT 246.000 345.600 247.800 346.200 ;
        RECT 240.200 344.400 241.000 345.600 ;
        RECT 247.000 344.400 247.800 345.600 ;
        RECT 240.200 343.600 242.000 344.400 ;
        RECT 247.000 343.600 248.400 344.400 ;
        RECT 240.200 342.200 241.000 343.600 ;
        RECT 247.000 342.200 247.800 343.600 ;
        RECT 250.800 342.200 251.600 349.700 ;
        RECT 254.000 346.800 254.800 348.400 ;
        RECT 255.600 342.200 256.400 359.800 ;
        RECT 258.800 351.200 259.600 359.800 ;
        RECT 262.000 351.200 262.800 359.800 ;
        RECT 265.200 352.400 266.000 359.800 ;
        RECT 269.600 356.400 271.200 359.800 ;
        RECT 268.400 355.600 271.200 356.400 ;
        RECT 266.600 352.400 267.400 352.600 ;
        RECT 265.200 351.800 267.400 352.400 ;
        RECT 269.600 352.400 271.200 355.600 ;
        RECT 273.200 352.400 274.000 352.600 ;
        RECT 274.800 352.400 275.600 359.800 ;
        RECT 279.000 352.400 279.800 359.800 ;
        RECT 280.400 353.600 281.200 354.400 ;
        RECT 280.600 352.400 281.200 353.600 ;
        RECT 269.600 351.800 271.600 352.400 ;
        RECT 273.200 351.800 275.600 352.400 ;
        RECT 258.800 350.400 262.800 351.200 ;
        RECT 266.800 351.200 267.400 351.800 ;
        RECT 266.800 350.600 270.200 351.200 ;
        RECT 269.400 350.400 270.200 350.600 ;
        RECT 271.000 350.400 271.600 351.800 ;
        RECT 278.000 351.600 280.000 352.400 ;
        RECT 280.600 351.800 282.000 352.400 ;
        RECT 281.200 351.600 282.000 351.800 ;
        RECT 282.800 351.600 283.600 353.200 ;
        RECT 258.800 347.600 259.600 350.400 ;
        RECT 267.200 349.800 268.000 350.000 ;
        RECT 271.000 349.800 272.400 350.400 ;
        RECT 267.200 349.200 269.800 349.800 ;
        RECT 269.200 348.600 269.800 349.200 ;
        RECT 270.600 349.600 272.400 349.800 ;
        RECT 276.400 350.300 277.200 350.400 ;
        RECT 278.000 350.300 278.800 350.400 ;
        RECT 276.400 349.700 278.800 350.300 ;
        RECT 276.400 349.600 277.200 349.700 ;
        RECT 270.600 349.200 271.600 349.600 ;
        RECT 258.800 346.800 262.800 347.600 ;
        RECT 263.600 346.800 264.400 348.400 ;
        RECT 265.200 348.200 266.800 348.400 ;
        RECT 265.200 347.600 268.600 348.200 ;
        RECT 269.200 347.800 270.000 348.600 ;
        RECT 268.000 347.200 268.600 347.600 ;
        RECT 266.600 346.800 267.400 347.000 ;
        RECT 258.800 342.200 259.600 346.800 ;
        RECT 262.000 342.200 262.800 346.800 ;
        RECT 265.200 346.200 267.400 346.800 ;
        RECT 268.000 346.600 270.000 347.200 ;
        RECT 268.400 346.400 270.000 346.600 ;
        RECT 265.200 342.200 266.000 346.200 ;
        RECT 270.600 345.800 271.200 349.200 ;
        RECT 278.000 348.800 278.800 349.700 ;
        RECT 279.400 348.400 280.000 351.600 ;
        RECT 281.300 350.300 281.900 351.600 ;
        RECT 284.400 350.300 285.200 359.800 ;
        RECT 292.400 352.400 293.200 359.800 ;
        RECT 295.600 352.400 296.400 359.800 ;
        RECT 292.400 351.800 296.400 352.400 ;
        RECT 297.200 351.800 298.000 359.800 ;
        RECT 299.400 352.600 300.200 359.800 ;
        RECT 299.400 351.800 301.200 352.600 ;
        RECT 304.200 352.400 305.000 359.800 ;
        RECT 303.600 351.800 305.000 352.400 ;
        RECT 293.200 350.400 294.000 350.800 ;
        RECT 297.200 350.400 297.800 351.800 ;
        RECT 281.300 349.700 285.200 350.300 ;
        RECT 272.000 347.600 272.800 348.400 ;
        RECT 274.000 347.600 275.600 348.400 ;
        RECT 276.400 348.200 277.200 348.400 ;
        RECT 276.400 347.600 278.000 348.200 ;
        RECT 279.400 347.600 282.000 348.400 ;
        RECT 272.000 347.200 272.600 347.600 ;
        RECT 277.200 347.200 278.000 347.600 ;
        RECT 271.800 346.400 272.600 347.200 ;
        RECT 273.200 346.800 274.000 347.000 ;
        RECT 273.200 346.200 275.600 346.800 ;
        RECT 276.600 346.200 280.200 346.600 ;
        RECT 281.200 346.200 281.800 347.600 ;
        RECT 284.400 346.200 285.200 349.700 ;
        RECT 292.400 349.800 294.000 350.400 ;
        RECT 295.600 349.800 298.000 350.400 ;
        RECT 292.400 349.600 293.200 349.800 ;
        RECT 286.000 346.800 286.800 348.400 ;
        RECT 294.000 347.600 294.800 349.200 ;
        RECT 269.600 342.200 271.200 345.800 ;
        RECT 274.800 342.200 275.600 346.200 ;
        RECT 276.400 346.000 280.400 346.200 ;
        RECT 276.400 342.200 277.200 346.000 ;
        RECT 279.600 342.200 280.400 346.000 ;
        RECT 281.200 342.200 282.000 346.200 ;
        RECT 283.400 345.600 285.200 346.200 ;
        RECT 295.600 346.400 296.200 349.800 ;
        RECT 297.200 349.600 298.000 349.800 ;
        RECT 298.800 349.600 299.600 351.200 ;
        RECT 300.400 348.400 301.000 351.800 ;
        RECT 303.600 351.600 304.400 351.800 ;
        RECT 303.600 350.400 304.200 351.600 ;
        RECT 308.400 351.200 309.200 359.800 ;
        RECT 312.600 352.600 313.400 359.800 ;
        RECT 311.600 351.800 313.400 352.600 ;
        RECT 305.200 350.800 309.200 351.200 ;
        RECT 305.000 350.600 309.200 350.800 ;
        RECT 303.600 349.600 304.400 350.400 ;
        RECT 305.000 350.000 305.800 350.600 ;
        RECT 300.400 347.600 301.200 348.400 ;
        RECT 283.400 342.200 284.200 345.600 ;
        RECT 295.600 342.200 296.400 346.400 ;
        RECT 297.200 346.300 298.000 346.400 ;
        RECT 300.400 346.300 301.000 347.600 ;
        RECT 297.200 345.700 301.100 346.300 ;
        RECT 297.200 345.600 298.000 345.700 ;
        RECT 297.000 344.800 297.800 345.600 ;
        RECT 300.400 344.200 301.000 345.700 ;
        RECT 302.000 344.800 302.800 346.400 ;
        RECT 303.600 346.200 304.200 349.600 ;
        RECT 305.000 347.000 305.600 350.000 ;
        RECT 306.400 348.400 307.200 349.200 ;
        RECT 311.800 348.400 312.400 351.800 ;
        RECT 313.200 349.600 314.000 351.200 ;
        RECT 314.800 350.300 315.600 350.400 ;
        RECT 316.400 350.300 317.200 359.800 ;
        RECT 318.600 352.600 319.400 359.800 ;
        RECT 325.000 356.400 325.800 359.800 ;
        RECT 325.000 355.600 326.800 356.400 ;
        RECT 323.600 353.600 324.400 354.400 ;
        RECT 318.600 351.800 320.400 352.600 ;
        RECT 323.600 352.400 324.200 353.600 ;
        RECT 325.000 352.400 325.800 355.600 ;
        RECT 322.800 351.800 324.200 352.400 ;
        RECT 324.800 351.800 325.800 352.400 ;
        RECT 318.000 350.300 318.800 351.200 ;
        RECT 314.800 349.700 318.800 350.300 ;
        RECT 314.800 349.600 315.600 349.700 ;
        RECT 306.600 348.300 307.600 348.400 ;
        RECT 311.600 348.300 312.400 348.400 ;
        RECT 306.600 347.700 312.400 348.300 ;
        RECT 306.600 347.600 307.600 347.700 ;
        RECT 311.600 347.600 312.400 347.700 ;
        RECT 305.000 346.400 307.400 347.000 ;
        RECT 300.400 342.200 301.200 344.200 ;
        RECT 303.600 342.200 304.400 346.200 ;
        RECT 306.800 344.200 307.400 346.400 ;
        RECT 308.400 344.800 309.200 346.400 ;
        RECT 310.000 344.800 310.800 346.400 ;
        RECT 311.800 344.400 312.400 347.600 ;
        RECT 313.200 346.300 314.000 346.400 ;
        RECT 314.800 346.300 315.600 346.400 ;
        RECT 313.200 345.700 315.600 346.300 ;
        RECT 313.200 345.600 314.000 345.700 ;
        RECT 314.800 344.800 315.600 345.700 ;
        RECT 306.800 342.200 307.600 344.200 ;
        RECT 311.600 342.200 312.400 344.400 ;
        RECT 316.400 342.200 317.200 349.700 ;
        RECT 318.000 349.600 318.800 349.700 ;
        RECT 319.600 348.400 320.200 351.800 ;
        RECT 322.800 351.600 323.600 351.800 ;
        RECT 324.800 348.400 325.400 351.800 ;
        RECT 326.000 350.300 326.800 350.400 ;
        RECT 329.200 350.300 330.000 359.800 ;
        RECT 330.800 354.300 331.600 354.400 ;
        RECT 332.400 354.300 333.200 359.800 ;
        RECT 336.600 355.800 337.800 359.800 ;
        RECT 341.200 355.800 342.000 359.800 ;
        RECT 345.600 356.400 346.400 359.800 ;
        RECT 345.600 355.800 347.600 356.400 ;
        RECT 337.200 355.000 338.000 355.800 ;
        RECT 341.400 355.200 342.000 355.800 ;
        RECT 340.600 354.600 344.200 355.200 ;
        RECT 346.800 355.000 347.600 355.800 ;
        RECT 340.600 354.400 341.400 354.600 ;
        RECT 343.400 354.400 344.200 354.600 ;
        RECT 330.800 353.700 333.200 354.300 ;
        RECT 330.800 353.600 331.600 353.700 ;
        RECT 326.000 349.700 330.000 350.300 ;
        RECT 326.000 348.800 326.800 349.700 ;
        RECT 319.600 347.600 320.400 348.400 ;
        RECT 322.800 347.600 325.400 348.400 ;
        RECT 327.600 348.200 328.400 348.400 ;
        RECT 326.800 347.600 328.400 348.200 ;
        RECT 319.600 344.400 320.200 347.600 ;
        RECT 321.200 344.800 322.000 346.400 ;
        RECT 323.000 346.200 323.600 347.600 ;
        RECT 326.800 347.200 327.600 347.600 ;
        RECT 324.600 346.200 328.200 346.600 ;
        RECT 319.600 342.200 320.400 344.400 ;
        RECT 322.800 342.200 323.600 346.200 ;
        RECT 324.400 346.000 328.400 346.200 ;
        RECT 324.400 342.200 325.200 346.000 ;
        RECT 327.600 342.200 328.400 346.000 ;
        RECT 329.200 342.200 330.000 349.700 ;
        RECT 332.400 351.200 333.200 353.700 ;
        RECT 336.400 353.200 337.800 354.000 ;
        RECT 337.200 352.200 337.800 353.200 ;
        RECT 339.400 353.000 341.600 353.600 ;
        RECT 339.400 352.800 340.200 353.000 ;
        RECT 337.200 351.600 339.600 352.200 ;
        RECT 332.400 350.600 336.600 351.200 ;
        RECT 332.400 347.200 333.200 350.600 ;
        RECT 335.800 350.400 336.600 350.600 ;
        RECT 339.000 350.400 339.600 351.600 ;
        RECT 341.000 351.800 341.600 353.000 ;
        RECT 342.200 353.000 343.000 353.200 ;
        RECT 346.800 353.000 347.600 353.200 ;
        RECT 342.200 352.400 347.600 353.000 ;
        RECT 341.000 351.400 345.800 351.800 ;
        RECT 350.000 351.400 350.800 359.800 ;
        RECT 341.000 351.200 350.800 351.400 ;
        RECT 345.000 351.000 350.800 351.200 ;
        RECT 345.200 350.800 350.800 351.000 ;
        RECT 334.200 349.800 335.000 350.000 ;
        RECT 334.200 349.200 338.000 349.800 ;
        RECT 338.800 349.600 339.600 350.400 ;
        RECT 343.600 350.200 344.400 350.400 ;
        RECT 343.600 349.600 348.600 350.200 ;
        RECT 337.200 349.000 338.000 349.200 ;
        RECT 339.000 348.400 339.600 349.600 ;
        RECT 345.200 349.400 346.000 349.600 ;
        RECT 347.800 349.400 348.600 349.600 ;
        RECT 346.200 348.400 347.000 348.600 ;
        RECT 339.000 347.800 350.000 348.400 ;
        RECT 339.400 347.600 340.200 347.800 ;
        RECT 332.400 346.600 336.200 347.200 ;
        RECT 330.800 344.800 331.600 346.400 ;
        RECT 332.400 342.200 333.200 346.600 ;
        RECT 335.400 346.400 336.200 346.600 ;
        RECT 345.200 346.400 345.800 347.800 ;
        RECT 348.400 347.600 350.000 347.800 ;
        RECT 343.400 345.400 344.200 345.600 ;
        RECT 337.200 344.200 338.000 345.000 ;
        RECT 341.400 344.800 344.200 345.400 ;
        RECT 345.200 344.800 346.000 346.400 ;
        RECT 341.400 344.200 342.000 344.800 ;
        RECT 346.800 344.200 347.600 345.000 ;
        RECT 336.600 343.600 338.000 344.200 ;
        RECT 336.600 342.200 337.800 343.600 ;
        RECT 341.200 342.200 342.000 344.200 ;
        RECT 345.600 343.600 347.600 344.200 ;
        RECT 345.600 342.200 346.400 343.600 ;
        RECT 350.000 342.200 350.800 347.000 ;
        RECT 351.600 342.200 352.400 359.800 ;
        RECT 354.800 351.200 355.600 359.800 ;
        RECT 359.000 355.800 360.200 359.800 ;
        RECT 363.600 355.800 364.400 359.800 ;
        RECT 368.000 356.400 368.800 359.800 ;
        RECT 368.000 355.800 370.000 356.400 ;
        RECT 359.600 355.000 360.400 355.800 ;
        RECT 363.800 355.200 364.400 355.800 ;
        RECT 363.000 354.600 366.600 355.200 ;
        RECT 369.200 355.000 370.000 355.800 ;
        RECT 363.000 354.400 363.800 354.600 ;
        RECT 365.800 354.400 366.600 354.600 ;
        RECT 358.800 353.200 360.200 354.000 ;
        RECT 359.600 352.200 360.200 353.200 ;
        RECT 361.800 353.000 364.000 353.600 ;
        RECT 361.800 352.800 362.600 353.000 ;
        RECT 359.600 351.600 362.000 352.200 ;
        RECT 354.800 350.600 359.000 351.200 ;
        RECT 354.800 347.200 355.600 350.600 ;
        RECT 358.200 350.400 359.000 350.600 ;
        RECT 356.600 349.800 357.400 350.000 ;
        RECT 356.600 349.200 360.400 349.800 ;
        RECT 359.600 349.000 360.400 349.200 ;
        RECT 361.400 348.400 362.000 351.600 ;
        RECT 363.400 351.800 364.000 353.000 ;
        RECT 364.600 353.000 365.400 353.200 ;
        RECT 369.200 353.000 370.000 353.200 ;
        RECT 364.600 352.400 370.000 353.000 ;
        RECT 363.400 351.400 368.200 351.800 ;
        RECT 372.400 351.400 373.200 359.800 ;
        RECT 374.000 352.400 374.800 359.800 ;
        RECT 374.000 351.800 376.200 352.400 ;
        RECT 377.200 351.800 378.000 359.800 ;
        RECT 378.800 352.400 379.600 359.800 ;
        RECT 380.200 352.400 381.000 352.600 ;
        RECT 378.800 351.800 381.000 352.400 ;
        RECT 383.200 352.400 384.800 359.800 ;
        RECT 386.800 352.400 387.600 352.600 ;
        RECT 388.400 352.400 389.200 359.800 ;
        RECT 383.200 351.800 385.200 352.400 ;
        RECT 386.800 351.800 389.200 352.400 ;
        RECT 363.400 351.200 373.200 351.400 ;
        RECT 367.400 351.000 373.200 351.200 ;
        RECT 367.600 350.800 373.200 351.000 ;
        RECT 375.600 351.200 376.200 351.800 ;
        RECT 375.600 350.400 376.800 351.200 ;
        RECT 364.400 350.300 365.200 350.400 ;
        RECT 366.000 350.300 366.800 350.400 ;
        RECT 364.400 350.200 366.800 350.300 ;
        RECT 364.400 349.700 371.000 350.200 ;
        RECT 364.400 349.600 365.200 349.700 ;
        RECT 366.000 349.600 371.000 349.700 ;
        RECT 370.200 349.400 371.000 349.600 ;
        RECT 374.000 348.800 374.800 350.400 ;
        RECT 368.600 348.400 369.400 348.600 ;
        RECT 361.400 347.800 372.400 348.400 ;
        RECT 361.800 347.600 362.600 347.800 ;
        RECT 354.800 346.600 358.600 347.200 ;
        RECT 353.200 344.800 354.000 346.400 ;
        RECT 354.800 342.200 355.600 346.600 ;
        RECT 357.800 346.400 358.600 346.600 ;
        RECT 367.600 346.400 368.200 347.800 ;
        RECT 370.800 347.600 372.400 347.800 ;
        RECT 375.600 347.400 376.200 350.400 ;
        RECT 377.400 349.600 378.000 351.800 ;
        RECT 380.400 351.200 381.000 351.800 ;
        RECT 380.400 350.600 383.800 351.200 ;
        RECT 383.000 350.400 383.800 350.600 ;
        RECT 384.600 350.400 385.200 351.800 ;
        RECT 365.800 345.400 366.600 345.600 ;
        RECT 359.600 344.200 360.400 345.000 ;
        RECT 363.800 344.800 366.600 345.400 ;
        RECT 367.600 344.800 368.400 346.400 ;
        RECT 363.800 344.200 364.400 344.800 ;
        RECT 369.200 344.200 370.000 345.000 ;
        RECT 359.000 343.600 360.400 344.200 ;
        RECT 359.000 342.200 360.200 343.600 ;
        RECT 363.600 342.200 364.400 344.200 ;
        RECT 368.000 343.600 370.000 344.200 ;
        RECT 368.000 342.200 368.800 343.600 ;
        RECT 372.400 342.200 373.200 347.000 ;
        RECT 374.000 346.800 376.200 347.400 ;
        RECT 374.000 342.200 374.800 346.800 ;
        RECT 377.200 342.200 378.000 349.600 ;
        RECT 380.800 349.800 381.600 350.000 ;
        RECT 384.600 349.800 386.000 350.400 ;
        RECT 380.800 349.200 383.400 349.800 ;
        RECT 382.800 348.600 383.400 349.200 ;
        RECT 384.200 349.600 386.000 349.800 ;
        RECT 384.200 349.200 385.200 349.600 ;
        RECT 378.800 348.200 380.400 348.400 ;
        RECT 378.800 347.600 382.200 348.200 ;
        RECT 382.800 347.800 383.600 348.600 ;
        RECT 381.600 347.200 382.200 347.600 ;
        RECT 380.200 346.800 381.000 347.000 ;
        RECT 378.800 346.200 381.000 346.800 ;
        RECT 381.600 346.600 383.600 347.200 ;
        RECT 382.000 346.400 383.600 346.600 ;
        RECT 378.800 342.200 379.600 346.200 ;
        RECT 384.200 345.800 384.800 349.200 ;
        RECT 385.600 347.600 386.400 348.400 ;
        RECT 387.600 348.300 389.200 348.400 ;
        RECT 390.000 348.300 390.800 359.800 ;
        RECT 393.200 351.200 394.000 359.800 ;
        RECT 397.400 355.800 398.600 359.800 ;
        RECT 402.000 355.800 402.800 359.800 ;
        RECT 406.400 356.400 407.200 359.800 ;
        RECT 406.400 355.800 408.400 356.400 ;
        RECT 398.000 355.000 398.800 355.800 ;
        RECT 402.200 355.200 402.800 355.800 ;
        RECT 401.400 354.600 405.000 355.200 ;
        RECT 407.600 355.000 408.400 355.800 ;
        RECT 401.400 354.400 402.200 354.600 ;
        RECT 404.200 354.400 405.000 354.600 ;
        RECT 397.200 353.200 398.600 354.000 ;
        RECT 398.000 352.200 398.600 353.200 ;
        RECT 400.200 353.000 402.400 353.600 ;
        RECT 400.200 352.800 401.000 353.000 ;
        RECT 398.000 351.600 400.400 352.200 ;
        RECT 393.200 350.600 397.400 351.200 ;
        RECT 387.600 347.700 390.800 348.300 ;
        RECT 387.600 347.600 389.200 347.700 ;
        RECT 385.600 347.200 386.200 347.600 ;
        RECT 385.400 346.400 386.200 347.200 ;
        RECT 386.800 346.800 387.600 347.000 ;
        RECT 386.800 346.200 389.200 346.800 ;
        RECT 383.200 342.200 384.800 345.800 ;
        RECT 388.400 342.200 389.200 346.200 ;
        RECT 390.000 342.200 390.800 347.700 ;
        RECT 391.600 346.800 392.400 348.400 ;
        RECT 393.200 347.200 394.000 350.600 ;
        RECT 396.600 350.400 397.400 350.600 ;
        RECT 395.000 349.800 395.800 350.000 ;
        RECT 395.000 349.200 398.800 349.800 ;
        RECT 398.000 349.000 398.800 349.200 ;
        RECT 399.800 348.400 400.400 351.600 ;
        RECT 401.800 351.800 402.400 353.000 ;
        RECT 403.000 353.000 403.800 353.200 ;
        RECT 407.600 353.000 408.400 353.200 ;
        RECT 403.000 352.400 408.400 353.000 ;
        RECT 401.800 351.400 406.600 351.800 ;
        RECT 410.800 351.400 411.600 359.800 ;
        RECT 413.200 353.600 414.000 354.400 ;
        RECT 413.200 352.400 413.800 353.600 ;
        RECT 414.600 352.400 415.400 359.800 ;
        RECT 419.600 353.600 420.400 354.400 ;
        RECT 419.600 352.400 420.200 353.600 ;
        RECT 421.000 352.400 421.800 359.800 ;
        RECT 412.400 351.800 413.800 352.400 ;
        RECT 414.400 351.800 415.400 352.400 ;
        RECT 418.800 351.800 420.200 352.400 ;
        RECT 420.800 351.800 421.800 352.400 ;
        RECT 427.800 352.400 428.600 359.800 ;
        RECT 429.200 353.600 430.000 354.400 ;
        RECT 429.400 352.400 430.000 353.600 ;
        RECT 432.400 353.600 433.200 354.400 ;
        RECT 432.400 352.400 433.000 353.600 ;
        RECT 433.800 352.400 434.600 359.800 ;
        RECT 427.800 351.800 428.800 352.400 ;
        RECT 429.400 351.800 430.800 352.400 ;
        RECT 412.400 351.600 413.200 351.800 ;
        RECT 401.800 351.200 411.600 351.400 ;
        RECT 405.800 351.000 411.600 351.200 ;
        RECT 406.000 350.800 411.600 351.000 ;
        RECT 404.400 350.200 405.200 350.400 ;
        RECT 412.400 350.300 413.200 350.400 ;
        RECT 414.400 350.300 415.000 351.800 ;
        RECT 418.800 351.600 419.600 351.800 ;
        RECT 404.400 349.600 409.400 350.200 ;
        RECT 412.400 349.700 415.000 350.300 ;
        RECT 412.400 349.600 413.200 349.700 ;
        RECT 406.000 349.400 406.800 349.600 ;
        RECT 408.600 349.400 409.400 349.600 ;
        RECT 407.000 348.400 407.800 348.600 ;
        RECT 414.400 348.400 415.000 349.700 ;
        RECT 415.600 348.800 416.400 350.400 ;
        RECT 417.200 350.300 418.000 350.400 ;
        RECT 420.800 350.300 421.400 351.800 ;
        RECT 417.200 349.700 421.400 350.300 ;
        RECT 417.200 349.600 418.000 349.700 ;
        RECT 420.800 348.400 421.400 349.700 ;
        RECT 422.000 350.300 422.800 350.400 ;
        RECT 426.800 350.300 427.600 350.400 ;
        RECT 422.000 349.700 427.600 350.300 ;
        RECT 422.000 348.800 422.800 349.700 ;
        RECT 426.800 348.800 427.600 349.700 ;
        RECT 428.200 348.400 428.800 351.800 ;
        RECT 430.000 351.600 430.800 351.800 ;
        RECT 431.600 351.800 433.000 352.400 ;
        RECT 433.600 351.800 434.600 352.400 ;
        RECT 431.600 351.600 432.400 351.800 ;
        RECT 430.100 350.400 430.700 351.600 ;
        RECT 430.000 350.300 430.800 350.400 ;
        RECT 433.600 350.300 434.200 351.800 ;
        RECT 430.000 349.700 434.200 350.300 ;
        RECT 430.000 349.600 430.800 349.700 ;
        RECT 433.600 348.400 434.200 349.700 ;
        RECT 434.800 348.800 435.600 350.400 ;
        RECT 399.800 347.800 410.800 348.400 ;
        RECT 400.200 347.600 401.000 347.800 ;
        RECT 402.800 347.600 403.600 347.800 ;
        RECT 393.200 346.600 397.000 347.200 ;
        RECT 393.200 342.200 394.000 346.600 ;
        RECT 396.200 346.400 397.000 346.600 ;
        RECT 406.000 345.600 406.600 347.800 ;
        RECT 409.200 347.600 410.800 347.800 ;
        RECT 412.400 347.600 415.000 348.400 ;
        RECT 417.200 348.200 418.000 348.400 ;
        RECT 416.400 347.600 418.000 348.200 ;
        RECT 418.800 347.600 421.400 348.400 ;
        RECT 423.600 348.200 424.400 348.400 ;
        RECT 422.800 347.600 424.400 348.200 ;
        RECT 425.200 348.200 426.000 348.400 ;
        RECT 425.200 347.600 426.800 348.200 ;
        RECT 428.200 347.600 430.800 348.400 ;
        RECT 431.600 347.600 434.200 348.400 ;
        RECT 436.400 348.300 437.200 348.400 ;
        RECT 438.000 348.300 438.800 359.800 ;
        RECT 436.400 348.200 438.800 348.300 ;
        RECT 435.600 347.700 438.800 348.200 ;
        RECT 435.600 347.600 437.200 347.700 ;
        RECT 404.200 345.400 405.000 345.600 ;
        RECT 398.000 344.200 398.800 345.000 ;
        RECT 402.200 344.800 405.000 345.400 ;
        RECT 406.000 344.800 406.800 345.600 ;
        RECT 402.200 344.200 402.800 344.800 ;
        RECT 407.600 344.200 408.400 345.000 ;
        RECT 397.400 343.600 398.800 344.200 ;
        RECT 397.400 342.200 398.600 343.600 ;
        RECT 402.000 342.200 402.800 344.200 ;
        RECT 406.400 343.600 408.400 344.200 ;
        RECT 406.400 342.200 407.200 343.600 ;
        RECT 410.800 342.200 411.600 347.000 ;
        RECT 412.600 346.200 413.200 347.600 ;
        RECT 416.400 347.200 417.200 347.600 ;
        RECT 414.200 346.200 417.800 346.600 ;
        RECT 419.000 346.200 419.600 347.600 ;
        RECT 422.800 347.200 423.600 347.600 ;
        RECT 426.000 347.200 426.800 347.600 ;
        RECT 420.600 346.200 424.200 346.600 ;
        RECT 425.400 346.200 429.000 346.600 ;
        RECT 430.000 346.200 430.600 347.600 ;
        RECT 431.800 346.200 432.400 347.600 ;
        RECT 435.600 347.200 436.400 347.600 ;
        RECT 433.400 346.200 437.000 346.600 ;
        RECT 412.400 342.200 413.200 346.200 ;
        RECT 414.000 346.000 418.000 346.200 ;
        RECT 414.000 342.200 414.800 346.000 ;
        RECT 417.200 342.200 418.000 346.000 ;
        RECT 418.800 342.200 419.600 346.200 ;
        RECT 420.400 346.000 424.400 346.200 ;
        RECT 420.400 342.200 421.200 346.000 ;
        RECT 423.600 342.200 424.400 346.000 ;
        RECT 425.200 346.000 429.200 346.200 ;
        RECT 425.200 342.200 426.000 346.000 ;
        RECT 428.400 342.200 429.200 346.000 ;
        RECT 430.000 342.200 430.800 346.200 ;
        RECT 431.600 342.200 432.400 346.200 ;
        RECT 433.200 346.000 437.200 346.200 ;
        RECT 433.200 342.200 434.000 346.000 ;
        RECT 436.400 342.200 437.200 346.000 ;
        RECT 438.000 342.200 438.800 347.700 ;
        RECT 439.600 344.800 440.400 346.400 ;
        RECT 441.200 342.200 442.000 359.800 ;
        RECT 451.800 352.600 452.600 359.800 ;
        RECT 450.800 351.800 452.600 352.600 ;
        RECT 450.800 351.600 451.600 351.800 ;
        RECT 451.000 348.400 451.600 351.600 ;
        RECT 452.400 349.600 453.200 351.200 ;
        RECT 450.800 347.600 451.600 348.400 ;
        RECT 442.800 344.800 443.600 346.400 ;
        RECT 449.200 344.800 450.000 346.400 ;
        RECT 451.000 344.200 451.600 347.600 ;
        RECT 454.000 346.800 454.800 348.400 ;
        RECT 455.600 346.200 456.400 359.800 ;
        RECT 457.200 351.600 458.000 353.200 ;
        RECT 458.800 351.800 459.600 359.800 ;
        RECT 460.400 352.400 461.200 359.800 ;
        RECT 463.600 352.400 464.400 359.800 ;
        RECT 460.400 351.800 464.400 352.400 ;
        RECT 459.000 350.400 459.600 351.800 ;
        RECT 462.800 350.400 463.600 350.800 ;
        RECT 458.800 349.800 461.200 350.400 ;
        RECT 462.800 349.800 464.400 350.400 ;
        RECT 458.800 349.600 459.600 349.800 ;
        RECT 455.600 345.600 457.400 346.200 ;
        RECT 458.800 345.600 459.600 346.400 ;
        RECT 460.600 346.200 461.200 349.800 ;
        RECT 463.600 349.600 464.400 349.800 ;
        RECT 462.000 348.300 462.800 349.200 ;
        RECT 463.600 348.300 464.400 348.400 ;
        RECT 465.200 348.300 466.000 348.400 ;
        RECT 462.000 347.700 466.000 348.300 ;
        RECT 462.000 347.600 462.800 347.700 ;
        RECT 463.600 347.600 464.400 347.700 ;
        RECT 465.200 346.800 466.000 347.700 ;
        RECT 456.600 344.400 457.400 345.600 ;
        RECT 459.000 344.800 459.800 345.600 ;
        RECT 450.800 342.200 451.600 344.200 ;
        RECT 455.600 343.600 457.400 344.400 ;
        RECT 456.600 342.200 457.400 343.600 ;
        RECT 460.400 342.200 461.200 346.200 ;
        RECT 466.800 346.200 467.600 359.800 ;
        RECT 468.400 351.600 469.200 353.200 ;
        RECT 470.000 352.400 470.800 359.800 ;
        RECT 471.600 352.400 472.400 352.600 ;
        RECT 474.400 352.400 476.000 359.800 ;
        RECT 470.000 351.800 472.400 352.400 ;
        RECT 474.000 351.800 476.000 352.400 ;
        RECT 478.200 352.400 479.000 352.600 ;
        RECT 479.600 352.400 480.400 359.800 ;
        RECT 478.200 351.800 480.400 352.400 ;
        RECT 474.000 350.400 474.600 351.800 ;
        RECT 478.200 351.200 478.800 351.800 ;
        RECT 475.400 350.600 478.800 351.200 ;
        RECT 481.200 351.200 482.000 359.800 ;
        RECT 485.400 355.800 486.600 359.800 ;
        RECT 490.000 355.800 490.800 359.800 ;
        RECT 494.400 356.400 495.200 359.800 ;
        RECT 494.400 355.800 496.400 356.400 ;
        RECT 486.000 355.000 486.800 355.800 ;
        RECT 490.200 355.200 490.800 355.800 ;
        RECT 489.400 354.600 493.000 355.200 ;
        RECT 495.600 355.000 496.400 355.800 ;
        RECT 489.400 354.400 490.200 354.600 ;
        RECT 492.200 354.400 493.000 354.600 ;
        RECT 484.400 354.000 485.800 354.400 ;
        RECT 484.400 353.600 486.600 354.000 ;
        RECT 485.200 353.200 486.600 353.600 ;
        RECT 486.000 352.200 486.600 353.200 ;
        RECT 488.200 353.000 490.400 353.600 ;
        RECT 488.200 352.800 489.000 353.000 ;
        RECT 486.000 351.600 488.400 352.200 ;
        RECT 481.200 350.600 485.400 351.200 ;
        RECT 475.400 350.400 476.200 350.600 ;
        RECT 473.200 349.800 474.600 350.400 ;
        RECT 477.600 349.800 478.400 350.000 ;
        RECT 473.200 349.600 475.000 349.800 ;
        RECT 474.000 349.200 475.000 349.600 ;
        RECT 468.400 348.300 469.200 348.400 ;
        RECT 470.000 348.300 471.600 348.400 ;
        RECT 468.400 347.700 471.600 348.300 ;
        RECT 468.400 347.600 469.200 347.700 ;
        RECT 470.000 347.600 471.600 347.700 ;
        RECT 472.800 347.600 473.600 348.400 ;
        RECT 473.000 347.200 473.600 347.600 ;
        RECT 471.600 346.800 472.400 347.000 ;
        RECT 470.000 346.200 472.400 346.800 ;
        RECT 473.000 346.400 473.800 347.200 ;
        RECT 466.800 345.600 468.600 346.200 ;
        RECT 467.800 344.400 468.600 345.600 ;
        RECT 467.800 343.600 469.200 344.400 ;
        RECT 467.800 342.200 468.600 343.600 ;
        RECT 470.000 342.200 470.800 346.200 ;
        RECT 474.400 345.800 475.000 349.200 ;
        RECT 475.800 349.200 478.400 349.800 ;
        RECT 475.800 348.600 476.400 349.200 ;
        RECT 475.600 347.800 476.400 348.600 ;
        RECT 478.800 348.200 480.400 348.400 ;
        RECT 477.000 347.600 480.400 348.200 ;
        RECT 477.000 347.200 477.600 347.600 ;
        RECT 475.600 346.600 477.600 347.200 ;
        RECT 481.200 347.200 482.000 350.600 ;
        RECT 484.600 350.400 485.400 350.600 ;
        RECT 483.000 349.800 483.800 350.000 ;
        RECT 483.000 349.200 486.800 349.800 ;
        RECT 486.000 349.000 486.800 349.200 ;
        RECT 487.800 348.400 488.400 351.600 ;
        RECT 489.800 351.800 490.400 353.000 ;
        RECT 491.000 353.000 491.800 353.200 ;
        RECT 495.600 353.000 496.400 353.200 ;
        RECT 491.000 352.400 496.400 353.000 ;
        RECT 489.800 351.400 494.600 351.800 ;
        RECT 498.800 351.400 499.600 359.800 ;
        RECT 489.800 351.200 499.600 351.400 ;
        RECT 493.800 351.000 499.600 351.200 ;
        RECT 494.000 350.800 499.600 351.000 ;
        RECT 502.000 351.200 502.800 359.800 ;
        RECT 505.200 351.200 506.000 359.800 ;
        RECT 508.400 351.200 509.200 359.800 ;
        RECT 511.600 351.200 512.400 359.800 ;
        RECT 516.400 356.400 517.200 359.800 ;
        RECT 516.200 355.800 517.200 356.400 ;
        RECT 516.200 355.200 516.800 355.800 ;
        RECT 519.600 355.200 520.400 359.800 ;
        RECT 522.800 357.000 523.600 359.800 ;
        RECT 524.400 357.000 525.200 359.800 ;
        RECT 514.800 354.600 516.800 355.200 ;
        RECT 502.000 350.400 503.800 351.200 ;
        RECT 505.200 350.400 507.400 351.200 ;
        RECT 508.400 350.400 510.600 351.200 ;
        RECT 511.600 350.400 514.000 351.200 ;
        RECT 492.400 350.200 493.200 350.400 ;
        RECT 492.400 349.600 497.400 350.200 ;
        RECT 494.000 349.400 494.800 349.600 ;
        RECT 496.600 349.400 497.400 349.600 ;
        RECT 503.000 349.000 503.800 350.400 ;
        RECT 506.600 349.000 507.400 350.400 ;
        RECT 509.800 349.000 510.600 350.400 ;
        RECT 495.000 348.400 495.800 348.600 ;
        RECT 487.600 347.800 498.800 348.400 ;
        RECT 487.600 347.600 489.000 347.800 ;
        RECT 478.200 346.800 479.000 347.000 ;
        RECT 475.600 346.400 477.200 346.600 ;
        RECT 478.200 346.200 480.400 346.800 ;
        RECT 474.400 344.400 476.000 345.800 ;
        RECT 473.200 343.600 476.000 344.400 ;
        RECT 474.400 342.200 476.000 343.600 ;
        RECT 479.600 342.200 480.400 346.200 ;
        RECT 481.200 346.600 485.000 347.200 ;
        RECT 481.200 342.200 482.000 346.600 ;
        RECT 484.200 346.400 485.000 346.600 ;
        RECT 494.000 345.600 494.600 347.800 ;
        RECT 497.200 347.600 498.800 347.800 ;
        RECT 503.000 348.200 505.600 349.000 ;
        RECT 506.600 348.200 509.000 349.000 ;
        RECT 509.800 348.200 512.400 349.000 ;
        RECT 503.000 347.600 503.800 348.200 ;
        RECT 506.600 347.600 507.400 348.200 ;
        RECT 509.800 347.600 510.600 348.200 ;
        RECT 513.200 347.600 514.000 350.400 ;
        RECT 492.200 345.400 493.000 345.600 ;
        RECT 486.000 344.200 486.800 345.000 ;
        RECT 490.200 344.800 493.000 345.400 ;
        RECT 494.000 344.800 494.800 345.600 ;
        RECT 490.200 344.200 490.800 344.800 ;
        RECT 495.600 344.200 496.400 345.000 ;
        RECT 485.400 343.600 486.800 344.200 ;
        RECT 485.400 342.200 486.600 343.600 ;
        RECT 490.000 342.200 490.800 344.200 ;
        RECT 494.400 343.600 496.400 344.200 ;
        RECT 494.400 342.200 495.200 343.600 ;
        RECT 498.800 342.200 499.600 347.000 ;
        RECT 502.000 346.800 503.800 347.600 ;
        RECT 505.200 346.800 507.400 347.600 ;
        RECT 508.400 346.800 510.600 347.600 ;
        RECT 511.600 346.800 514.000 347.600 ;
        RECT 514.800 349.000 515.600 354.600 ;
        RECT 517.400 354.400 521.600 355.200 ;
        RECT 526.000 355.000 526.800 359.800 ;
        RECT 529.200 355.000 530.000 359.800 ;
        RECT 517.400 354.000 518.000 354.400 ;
        RECT 516.400 353.200 518.000 354.000 ;
        RECT 521.000 353.800 526.800 354.400 ;
        RECT 519.000 353.200 520.400 353.800 ;
        RECT 519.000 353.000 525.200 353.200 ;
        RECT 519.800 352.600 525.200 353.000 ;
        RECT 524.400 352.400 525.200 352.600 ;
        RECT 526.200 353.000 526.800 353.800 ;
        RECT 527.400 353.600 530.000 354.400 ;
        RECT 532.400 353.600 533.200 359.800 ;
        RECT 534.000 357.000 534.800 359.800 ;
        RECT 535.600 357.000 536.400 359.800 ;
        RECT 537.200 357.000 538.000 359.800 ;
        RECT 535.600 354.400 539.800 355.200 ;
        RECT 540.400 354.400 541.200 359.800 ;
        RECT 543.600 355.200 544.400 359.800 ;
        RECT 543.600 354.600 546.200 355.200 ;
        RECT 540.400 353.600 543.000 354.400 ;
        RECT 534.000 353.000 534.800 353.200 ;
        RECT 526.200 352.400 534.800 353.000 ;
        RECT 537.200 353.000 538.000 353.200 ;
        RECT 545.600 353.000 546.200 354.600 ;
        RECT 537.200 352.400 546.200 353.000 ;
        RECT 545.600 350.600 546.200 352.400 ;
        RECT 546.800 352.000 547.600 359.800 ;
        RECT 551.600 356.400 552.400 359.800 ;
        RECT 551.400 355.800 552.400 356.400 ;
        RECT 551.400 355.200 552.000 355.800 ;
        RECT 554.800 355.200 555.600 359.800 ;
        RECT 558.000 357.000 558.800 359.800 ;
        RECT 559.600 357.000 560.400 359.800 ;
        RECT 550.000 354.600 552.000 355.200 ;
        RECT 546.800 351.200 547.800 352.000 ;
        RECT 516.200 350.000 539.600 350.600 ;
        RECT 545.600 350.000 546.400 350.600 ;
        RECT 516.200 349.800 517.000 350.000 ;
        RECT 518.000 349.600 518.800 350.000 ;
        RECT 521.200 349.600 522.000 350.000 ;
        RECT 538.800 349.400 539.600 350.000 ;
        RECT 514.800 348.200 523.600 349.000 ;
        RECT 524.200 348.600 526.200 349.400 ;
        RECT 530.000 348.600 533.200 349.400 ;
        RECT 502.000 342.200 502.800 346.800 ;
        RECT 505.200 342.200 506.000 346.800 ;
        RECT 508.400 342.200 509.200 346.800 ;
        RECT 511.600 342.200 512.400 346.800 ;
        RECT 514.800 342.200 515.600 348.200 ;
        RECT 517.200 346.800 520.200 347.600 ;
        RECT 519.400 346.200 520.200 346.800 ;
        RECT 525.400 346.200 526.200 348.600 ;
        RECT 527.600 346.800 528.400 348.400 ;
        RECT 532.800 347.800 533.600 348.000 ;
        RECT 529.200 347.200 533.600 347.800 ;
        RECT 529.200 347.000 530.000 347.200 ;
        RECT 535.600 346.400 536.400 349.200 ;
        RECT 541.400 348.600 545.200 349.400 ;
        RECT 541.400 347.400 542.200 348.600 ;
        RECT 545.800 348.000 546.400 350.000 ;
        RECT 529.200 346.200 530.000 346.400 ;
        RECT 519.400 345.400 522.000 346.200 ;
        RECT 525.400 345.600 530.000 346.200 ;
        RECT 530.800 345.600 532.400 346.400 ;
        RECT 535.400 345.600 536.400 346.400 ;
        RECT 540.400 346.800 542.200 347.400 ;
        RECT 545.200 347.400 546.400 348.000 ;
        RECT 540.400 346.200 541.200 346.800 ;
        RECT 521.200 342.200 522.000 345.400 ;
        RECT 538.800 345.400 541.200 346.200 ;
        RECT 522.800 342.200 523.600 345.000 ;
        RECT 524.400 342.200 525.200 345.000 ;
        RECT 526.000 342.200 526.800 345.000 ;
        RECT 529.200 342.200 530.000 345.000 ;
        RECT 532.400 342.200 533.200 345.000 ;
        RECT 534.000 342.200 534.800 345.000 ;
        RECT 535.600 342.200 536.400 345.000 ;
        RECT 537.200 342.200 538.000 345.000 ;
        RECT 538.800 342.200 539.600 345.400 ;
        RECT 545.200 342.200 546.000 347.400 ;
        RECT 547.000 346.800 547.800 351.200 ;
        RECT 546.800 346.000 547.800 346.800 ;
        RECT 550.000 349.000 550.800 354.600 ;
        RECT 552.600 354.400 556.800 355.200 ;
        RECT 561.200 355.000 562.000 359.800 ;
        RECT 564.400 355.000 565.200 359.800 ;
        RECT 552.600 354.000 553.200 354.400 ;
        RECT 551.600 353.200 553.200 354.000 ;
        RECT 556.200 353.800 562.000 354.400 ;
        RECT 554.200 353.200 555.600 353.800 ;
        RECT 554.200 353.000 560.400 353.200 ;
        RECT 555.000 352.600 560.400 353.000 ;
        RECT 559.600 352.400 560.400 352.600 ;
        RECT 561.400 353.000 562.000 353.800 ;
        RECT 562.600 353.600 565.200 354.400 ;
        RECT 567.600 353.600 568.400 359.800 ;
        RECT 569.200 357.000 570.000 359.800 ;
        RECT 570.800 357.000 571.600 359.800 ;
        RECT 572.400 357.000 573.200 359.800 ;
        RECT 570.800 354.400 575.000 355.200 ;
        RECT 575.600 354.400 576.400 359.800 ;
        RECT 578.800 355.200 579.600 359.800 ;
        RECT 578.800 354.600 581.400 355.200 ;
        RECT 575.600 353.600 578.200 354.400 ;
        RECT 569.200 353.000 570.000 353.200 ;
        RECT 561.400 352.400 570.000 353.000 ;
        RECT 572.400 353.000 573.200 353.200 ;
        RECT 580.800 353.000 581.400 354.600 ;
        RECT 572.400 352.400 581.400 353.000 ;
        RECT 580.800 350.600 581.400 352.400 ;
        RECT 582.000 352.000 582.800 359.800 ;
        RECT 582.000 351.200 583.000 352.000 ;
        RECT 551.400 350.000 574.800 350.600 ;
        RECT 580.800 350.000 581.600 350.600 ;
        RECT 551.400 349.800 552.400 350.000 ;
        RECT 551.600 349.600 552.400 349.800 ;
        RECT 553.200 349.600 554.000 350.000 ;
        RECT 556.400 349.600 557.200 350.000 ;
        RECT 574.000 349.400 574.800 350.000 ;
        RECT 550.000 348.200 558.800 349.000 ;
        RECT 559.400 348.600 561.400 349.400 ;
        RECT 565.200 348.600 568.400 349.400 ;
        RECT 546.800 342.200 547.600 346.000 ;
        RECT 550.000 342.200 550.800 348.200 ;
        RECT 552.400 346.800 555.400 347.600 ;
        RECT 554.600 346.200 555.400 346.800 ;
        RECT 560.600 346.200 561.400 348.600 ;
        RECT 562.800 346.800 563.600 348.400 ;
        RECT 568.000 347.800 568.800 348.000 ;
        RECT 564.400 347.200 568.800 347.800 ;
        RECT 564.400 347.000 565.200 347.200 ;
        RECT 570.800 346.400 571.600 349.200 ;
        RECT 576.600 348.600 580.400 349.400 ;
        RECT 576.600 347.400 577.400 348.600 ;
        RECT 581.000 348.000 581.600 350.000 ;
        RECT 564.400 346.200 565.200 346.400 ;
        RECT 554.600 345.400 557.200 346.200 ;
        RECT 560.600 345.600 565.200 346.200 ;
        RECT 566.000 345.600 567.600 346.400 ;
        RECT 570.600 345.600 571.600 346.400 ;
        RECT 575.600 346.800 577.400 347.400 ;
        RECT 580.400 347.400 581.600 348.000 ;
        RECT 575.600 346.200 576.400 346.800 ;
        RECT 556.400 342.200 557.200 345.400 ;
        RECT 574.000 345.400 576.400 346.200 ;
        RECT 558.000 342.200 558.800 345.000 ;
        RECT 559.600 342.200 560.400 345.000 ;
        RECT 561.200 342.200 562.000 345.000 ;
        RECT 564.400 342.200 565.200 345.000 ;
        RECT 567.600 342.200 568.400 345.000 ;
        RECT 569.200 342.200 570.000 345.000 ;
        RECT 570.800 342.200 571.600 345.000 ;
        RECT 572.400 342.200 573.200 345.000 ;
        RECT 574.000 342.200 574.800 345.400 ;
        RECT 580.400 342.200 581.200 347.400 ;
        RECT 582.200 346.800 583.000 351.200 ;
        RECT 582.000 346.000 583.000 346.800 ;
        RECT 582.000 342.200 582.800 346.000 ;
        RECT 1.200 335.800 2.000 339.800 ;
        RECT 5.600 336.200 7.200 339.800 ;
        RECT 1.200 335.200 3.400 335.800 ;
        RECT 4.400 335.400 6.000 335.600 ;
        RECT 2.600 335.000 3.400 335.200 ;
        RECT 4.000 334.800 6.000 335.400 ;
        RECT 4.000 334.400 4.600 334.800 ;
        RECT 1.200 333.800 4.600 334.400 ;
        RECT 1.200 333.600 2.800 333.800 ;
        RECT 5.200 333.400 6.000 334.200 ;
        RECT 5.200 332.800 5.800 333.400 ;
        RECT 3.200 332.200 5.800 332.800 ;
        RECT 6.600 332.800 7.200 336.200 ;
        RECT 10.800 335.800 11.600 339.800 ;
        RECT 7.800 334.800 8.600 335.600 ;
        RECT 9.200 335.200 11.600 335.800 ;
        RECT 14.000 335.200 14.800 339.800 ;
        RECT 17.200 335.200 18.000 339.800 ;
        RECT 22.000 336.400 22.800 339.800 ;
        RECT 21.800 335.800 22.800 336.400 ;
        RECT 9.200 335.000 10.000 335.200 ;
        RECT 8.000 334.400 8.600 334.800 ;
        RECT 14.000 334.400 18.000 335.200 ;
        RECT 8.000 333.600 8.800 334.400 ;
        RECT 10.000 333.600 11.600 334.400 ;
        RECT 6.600 332.400 7.600 332.800 ;
        RECT 6.600 332.200 8.400 332.400 ;
        RECT 3.200 332.000 4.000 332.200 ;
        RECT 7.000 331.600 8.400 332.200 ;
        RECT 14.000 331.600 14.800 334.400 ;
        RECT 18.800 333.600 19.600 335.200 ;
        RECT 21.800 334.400 22.400 335.800 ;
        RECT 25.200 335.200 26.000 339.800 ;
        RECT 26.800 335.600 27.600 337.200 ;
        RECT 23.400 334.600 26.000 335.200 ;
        RECT 21.800 333.600 22.800 334.400 ;
        RECT 5.400 331.400 6.200 331.600 ;
        RECT 2.800 330.800 6.200 331.400 ;
        RECT 2.800 330.200 3.400 330.800 ;
        RECT 7.000 330.200 7.600 331.600 ;
        RECT 14.000 330.800 18.000 331.600 ;
        RECT 1.200 329.600 3.400 330.200 ;
        RECT 1.200 322.200 2.000 329.600 ;
        RECT 2.600 329.400 3.400 329.600 ;
        RECT 5.600 329.600 7.600 330.200 ;
        RECT 9.200 329.600 11.600 330.200 ;
        RECT 5.600 322.200 7.200 329.600 ;
        RECT 9.200 329.400 10.000 329.600 ;
        RECT 10.800 322.200 11.600 329.600 ;
        RECT 14.000 322.200 14.800 330.800 ;
        RECT 17.200 322.200 18.000 330.800 ;
        RECT 21.800 330.200 22.400 333.600 ;
        RECT 23.400 333.000 24.000 334.600 ;
        RECT 23.000 332.200 24.000 333.000 ;
        RECT 23.400 330.200 24.000 332.200 ;
        RECT 25.000 332.400 25.800 333.200 ;
        RECT 25.000 331.600 26.000 332.400 ;
        RECT 21.800 329.200 22.800 330.200 ;
        RECT 23.400 329.600 26.000 330.200 ;
        RECT 22.000 322.200 22.800 329.200 ;
        RECT 25.200 322.200 26.000 329.600 ;
        RECT 28.400 322.200 29.200 339.800 ;
        RECT 30.000 335.200 30.800 339.800 ;
        RECT 33.200 336.400 34.000 339.800 ;
        RECT 33.200 335.800 34.200 336.400 ;
        RECT 39.400 335.800 41.000 339.800 ;
        RECT 44.400 335.800 45.200 339.800 ;
        RECT 46.000 336.000 46.800 339.800 ;
        RECT 49.200 336.000 50.000 339.800 ;
        RECT 46.000 335.800 50.000 336.000 ;
        RECT 30.000 334.600 32.600 335.200 ;
        RECT 30.200 332.400 31.000 333.200 ;
        RECT 30.000 331.600 31.000 332.400 ;
        RECT 32.000 333.000 32.600 334.600 ;
        RECT 33.600 334.400 34.200 335.800 ;
        RECT 33.200 333.600 34.200 334.400 ;
        RECT 32.000 332.200 33.000 333.000 ;
        RECT 32.000 330.200 32.600 332.200 ;
        RECT 33.600 330.200 34.200 333.600 ;
        RECT 38.000 332.800 38.800 334.400 ;
        RECT 39.800 332.400 40.400 335.800 ;
        RECT 44.600 334.400 45.200 335.800 ;
        RECT 46.200 335.400 49.800 335.800 ;
        RECT 48.400 334.400 49.200 334.800 ;
        RECT 41.200 333.600 42.000 334.400 ;
        RECT 44.400 333.600 47.000 334.400 ;
        RECT 48.400 333.800 50.000 334.400 ;
        RECT 52.000 334.200 52.800 339.800 ;
        RECT 49.200 333.600 50.000 333.800 ;
        RECT 51.000 333.800 52.800 334.200 ;
        RECT 51.000 333.600 52.600 333.800 ;
        RECT 41.200 333.200 41.800 333.600 ;
        RECT 41.000 332.400 41.800 333.200 ;
        RECT 36.400 332.200 37.200 332.400 ;
        RECT 36.400 331.600 38.000 332.200 ;
        RECT 39.600 331.600 40.400 332.400 ;
        RECT 37.200 331.200 38.000 331.600 ;
        RECT 39.800 331.400 40.400 331.600 ;
        RECT 42.800 332.300 43.600 332.400 ;
        RECT 44.400 332.300 45.200 332.400 ;
        RECT 42.800 331.700 45.200 332.300 ;
        RECT 39.800 330.800 41.800 331.400 ;
        RECT 42.800 330.800 43.600 331.700 ;
        RECT 44.400 331.600 45.200 331.700 ;
        RECT 41.200 330.200 41.800 330.800 ;
        RECT 44.400 330.200 45.200 330.400 ;
        RECT 46.400 330.200 47.000 333.600 ;
        RECT 47.600 331.600 48.400 333.200 ;
        RECT 51.000 330.400 51.600 333.600 ;
        RECT 53.200 331.600 54.800 332.400 ;
        RECT 30.000 329.600 32.600 330.200 ;
        RECT 30.000 322.200 30.800 329.600 ;
        RECT 33.200 329.200 34.200 330.200 ;
        RECT 36.400 329.600 40.400 330.200 ;
        RECT 33.200 322.200 34.000 329.200 ;
        RECT 36.400 322.200 37.200 329.600 ;
        RECT 39.600 322.800 40.400 329.600 ;
        RECT 41.200 323.400 42.000 330.200 ;
        RECT 42.800 322.800 43.600 330.200 ;
        RECT 44.400 329.600 45.800 330.200 ;
        RECT 46.400 329.600 47.400 330.200 ;
        RECT 50.800 329.600 51.600 330.400 ;
        RECT 55.600 330.300 56.400 331.200 ;
        RECT 57.200 330.300 58.000 339.800 ;
        RECT 58.800 335.600 59.600 337.200 ;
        RECT 60.400 335.600 61.200 337.200 ;
        RECT 55.600 329.700 58.000 330.300 ;
        RECT 55.600 329.600 56.400 329.700 ;
        RECT 45.200 328.400 45.800 329.600 ;
        RECT 46.600 328.400 47.400 329.600 ;
        RECT 45.200 327.600 46.000 328.400 ;
        RECT 46.600 327.600 48.400 328.400 ;
        RECT 39.600 322.200 43.600 322.800 ;
        RECT 46.600 322.200 47.400 327.600 ;
        RECT 51.000 327.000 51.600 329.600 ;
        RECT 52.400 327.600 53.200 329.200 ;
        RECT 51.000 326.400 54.600 327.000 ;
        RECT 51.000 326.200 51.600 326.400 ;
        RECT 50.800 322.200 51.600 326.200 ;
        RECT 54.000 326.200 54.600 326.400 ;
        RECT 54.000 322.200 54.800 326.200 ;
        RECT 57.200 322.200 58.000 329.700 ;
        RECT 62.000 334.300 62.800 339.800 ;
        RECT 66.200 336.400 67.000 339.800 ;
        RECT 65.200 335.800 67.000 336.400 ;
        RECT 63.600 334.300 64.400 335.200 ;
        RECT 62.000 333.700 64.400 334.300 ;
        RECT 62.000 322.200 62.800 333.700 ;
        RECT 63.600 333.600 64.400 333.700 ;
        RECT 65.200 322.200 66.000 335.800 ;
        RECT 69.600 334.200 70.400 339.800 ;
        RECT 74.800 335.800 75.600 339.800 ;
        RECT 76.400 336.000 77.200 339.800 ;
        RECT 79.600 336.000 80.400 339.800 ;
        RECT 83.800 338.400 84.600 339.800 ;
        RECT 82.800 337.600 84.600 338.400 ;
        RECT 83.800 336.400 84.600 337.600 ;
        RECT 76.400 335.800 80.400 336.000 ;
        RECT 82.800 335.800 84.600 336.400 ;
        RECT 86.600 336.400 87.400 339.800 ;
        RECT 86.600 335.800 88.400 336.400 ;
        RECT 90.800 335.800 91.600 339.800 ;
        RECT 92.400 336.000 93.200 339.800 ;
        RECT 95.600 336.000 96.400 339.800 ;
        RECT 92.400 335.800 96.400 336.000 ;
        RECT 97.200 335.800 98.000 339.800 ;
        RECT 98.800 336.000 99.600 339.800 ;
        RECT 102.000 336.000 102.800 339.800 ;
        RECT 105.200 337.800 106.000 339.800 ;
        RECT 98.800 335.800 102.800 336.000 ;
        RECT 75.000 334.400 75.600 335.800 ;
        RECT 76.600 335.400 80.200 335.800 ;
        RECT 78.800 334.400 79.600 334.800 ;
        RECT 68.600 333.800 70.400 334.200 ;
        RECT 68.600 333.600 70.200 333.800 ;
        RECT 74.800 333.600 77.400 334.400 ;
        RECT 78.800 333.800 80.400 334.400 ;
        RECT 79.600 333.600 80.400 333.800 ;
        RECT 81.200 333.600 82.000 335.200 ;
        RECT 68.600 330.400 69.200 333.600 ;
        RECT 70.800 331.600 72.400 332.400 ;
        RECT 66.800 328.800 67.600 330.400 ;
        RECT 68.400 329.600 69.200 330.400 ;
        RECT 73.200 329.600 74.000 331.200 ;
        RECT 74.800 330.200 75.600 330.400 ;
        RECT 76.800 330.200 77.400 333.600 ;
        RECT 78.000 331.600 78.800 333.200 ;
        RECT 74.800 329.600 76.200 330.200 ;
        RECT 76.800 329.600 77.800 330.200 ;
        RECT 68.600 327.000 69.200 329.600 ;
        RECT 70.000 327.600 70.800 329.200 ;
        RECT 75.600 328.400 76.200 329.600 ;
        RECT 75.600 327.600 76.400 328.400 ;
        RECT 68.600 326.400 72.200 327.000 ;
        RECT 68.600 326.200 69.200 326.400 ;
        RECT 68.400 322.200 69.200 326.200 ;
        RECT 71.600 322.200 72.400 326.400 ;
        RECT 77.000 324.400 77.800 329.600 ;
        RECT 77.000 323.600 78.800 324.400 ;
        RECT 77.000 322.200 77.800 323.600 ;
        RECT 82.800 322.200 83.600 335.800 ;
        RECT 87.600 332.300 88.400 335.800 ;
        RECT 89.200 333.600 90.000 335.200 ;
        RECT 91.000 334.400 91.600 335.800 ;
        RECT 92.600 335.400 96.200 335.800 ;
        RECT 94.800 334.400 95.600 334.800 ;
        RECT 97.400 334.400 98.000 335.800 ;
        RECT 99.000 335.400 102.600 335.800 ;
        RECT 103.600 335.600 104.400 337.200 ;
        RECT 101.200 334.400 102.000 334.800 ;
        RECT 105.400 334.400 106.000 337.800 ;
        RECT 108.400 336.000 109.200 339.800 ;
        RECT 111.600 336.000 112.400 339.800 ;
        RECT 108.400 335.800 112.400 336.000 ;
        RECT 113.200 335.800 114.000 339.800 ;
        RECT 108.600 335.400 112.200 335.800 ;
        RECT 109.200 334.400 110.000 334.800 ;
        RECT 113.200 334.400 113.800 335.800 ;
        RECT 90.800 333.600 93.400 334.400 ;
        RECT 94.800 333.800 96.400 334.400 ;
        RECT 95.600 333.600 96.400 333.800 ;
        RECT 97.200 333.600 99.800 334.400 ;
        RECT 101.200 333.800 102.800 334.400 ;
        RECT 102.000 333.600 102.800 333.800 ;
        RECT 105.200 334.300 106.000 334.400 ;
        RECT 106.800 334.300 107.600 334.400 ;
        RECT 105.200 333.700 107.600 334.300 ;
        RECT 105.200 333.600 106.000 333.700 ;
        RECT 106.800 333.600 107.600 333.700 ;
        RECT 108.400 333.800 110.000 334.400 ;
        RECT 108.400 333.600 109.200 333.800 ;
        RECT 111.400 333.600 114.000 334.400 ;
        RECT 84.500 331.700 88.400 332.300 ;
        RECT 84.500 330.400 85.100 331.700 ;
        RECT 84.400 328.800 85.200 330.400 ;
        RECT 86.000 328.800 86.800 330.400 ;
        RECT 87.600 322.200 88.400 331.700 ;
        RECT 90.800 332.300 91.600 332.400 ;
        RECT 92.800 332.300 93.400 333.600 ;
        RECT 90.800 331.700 93.400 332.300 ;
        RECT 90.800 331.600 91.600 331.700 ;
        RECT 89.200 330.300 90.000 330.400 ;
        RECT 90.800 330.300 91.600 330.400 ;
        RECT 89.200 330.200 91.600 330.300 ;
        RECT 92.800 330.200 93.400 331.700 ;
        RECT 94.000 332.300 94.800 333.200 ;
        RECT 95.600 332.300 96.400 332.400 ;
        RECT 94.000 331.700 96.400 332.300 ;
        RECT 94.000 331.600 94.800 331.700 ;
        RECT 95.600 331.600 96.400 331.700 ;
        RECT 97.200 330.200 98.000 330.400 ;
        RECT 99.200 330.200 99.800 333.600 ;
        RECT 100.400 332.300 101.200 333.200 ;
        RECT 102.000 332.300 102.800 332.400 ;
        RECT 100.400 331.700 102.800 332.300 ;
        RECT 100.400 331.600 101.200 331.700 ;
        RECT 102.000 331.600 102.800 331.700 ;
        RECT 105.400 330.200 106.000 333.600 ;
        RECT 106.800 332.300 107.600 332.400 ;
        RECT 110.000 332.300 110.800 333.200 ;
        RECT 106.800 331.700 110.800 332.300 ;
        RECT 106.800 330.800 107.600 331.700 ;
        RECT 110.000 331.600 110.800 331.700 ;
        RECT 111.400 330.200 112.000 333.600 ;
        RECT 113.200 332.300 114.000 332.400 ;
        RECT 114.800 332.300 115.600 339.800 ;
        RECT 118.000 339.200 122.000 339.800 ;
        RECT 116.400 335.600 117.200 337.200 ;
        RECT 118.000 335.800 118.800 339.200 ;
        RECT 119.600 335.800 120.400 338.600 ;
        RECT 121.200 336.000 122.000 339.200 ;
        RECT 124.400 336.000 125.200 339.800 ;
        RECT 121.200 335.800 125.200 336.000 ;
        RECT 126.000 336.000 126.800 339.800 ;
        RECT 129.200 336.000 130.000 339.800 ;
        RECT 126.000 335.800 130.000 336.000 ;
        RECT 130.800 335.800 131.600 339.800 ;
        RECT 132.400 335.800 133.200 339.800 ;
        RECT 134.000 336.000 134.800 339.800 ;
        RECT 137.200 336.000 138.000 339.800 ;
        RECT 134.000 335.800 138.000 336.000 ;
        RECT 143.600 335.800 144.400 339.800 ;
        RECT 148.000 336.200 149.600 339.800 ;
        RECT 119.600 334.400 120.200 335.800 ;
        RECT 121.400 335.400 125.000 335.800 ;
        RECT 126.200 335.400 129.800 335.800 ;
        RECT 123.600 334.400 124.400 334.800 ;
        RECT 126.800 334.400 127.600 334.800 ;
        RECT 130.800 334.400 131.400 335.800 ;
        RECT 132.600 334.400 133.200 335.800 ;
        RECT 134.200 335.400 137.800 335.800 ;
        RECT 143.600 335.200 145.800 335.800 ;
        RECT 146.800 335.400 148.400 335.600 ;
        RECT 145.000 335.000 145.800 335.200 ;
        RECT 146.400 334.800 148.400 335.400 ;
        RECT 136.400 334.400 137.200 334.800 ;
        RECT 146.400 334.400 147.000 334.800 ;
        RECT 118.000 332.800 118.800 334.400 ;
        RECT 119.600 333.800 122.000 334.400 ;
        RECT 123.600 334.300 125.200 334.400 ;
        RECT 126.000 334.300 127.600 334.400 ;
        RECT 123.600 333.800 127.600 334.300 ;
        RECT 121.200 333.600 122.000 333.800 ;
        RECT 124.400 333.700 126.800 333.800 ;
        RECT 124.400 333.600 125.200 333.700 ;
        RECT 126.000 333.600 126.800 333.700 ;
        RECT 129.000 333.600 131.600 334.400 ;
        RECT 132.400 333.600 135.000 334.400 ;
        RECT 136.400 333.800 138.000 334.400 ;
        RECT 137.200 333.600 138.000 333.800 ;
        RECT 143.600 333.800 147.000 334.400 ;
        RECT 143.600 333.600 145.200 333.800 ;
        RECT 113.200 331.700 115.600 332.300 ;
        RECT 113.200 331.600 114.000 331.700 ;
        RECT 113.200 330.200 114.000 330.400 ;
        RECT 89.200 329.700 92.200 330.200 ;
        RECT 89.200 329.600 90.000 329.700 ;
        RECT 90.800 329.600 92.200 329.700 ;
        RECT 92.800 329.600 93.800 330.200 ;
        RECT 97.200 329.600 98.600 330.200 ;
        RECT 99.200 329.600 100.200 330.200 ;
        RECT 91.600 328.400 92.200 329.600 ;
        RECT 91.600 327.600 92.400 328.400 ;
        RECT 93.000 322.200 93.800 329.600 ;
        RECT 98.000 328.400 98.600 329.600 ;
        RECT 98.000 327.600 98.800 328.400 ;
        RECT 99.400 324.400 100.200 329.600 ;
        RECT 105.200 329.400 107.000 330.200 ;
        RECT 99.400 323.600 101.200 324.400 ;
        RECT 99.400 322.200 100.200 323.600 ;
        RECT 106.200 322.200 107.000 329.400 ;
        RECT 111.000 329.600 112.000 330.200 ;
        RECT 112.600 329.600 114.000 330.200 ;
        RECT 111.000 322.200 111.800 329.600 ;
        RECT 112.600 328.400 113.200 329.600 ;
        RECT 112.400 327.600 113.200 328.400 ;
        RECT 114.800 322.200 115.600 331.700 ;
        RECT 119.600 331.600 120.400 333.200 ;
        RECT 121.400 330.400 122.000 333.600 ;
        RECT 122.800 332.300 123.600 333.200 ;
        RECT 127.600 332.300 128.400 333.200 ;
        RECT 122.800 331.700 128.400 332.300 ;
        RECT 122.800 331.600 123.600 331.700 ;
        RECT 127.600 331.600 128.400 331.700 ;
        RECT 129.000 332.300 129.600 333.600 ;
        RECT 129.000 331.700 133.100 332.300 ;
        RECT 119.600 330.200 122.000 330.400 ;
        RECT 129.000 330.200 129.600 331.700 ;
        RECT 132.500 330.400 133.100 331.700 ;
        RECT 130.800 330.200 131.600 330.400 ;
        RECT 119.600 329.600 122.600 330.200 ;
        RECT 120.600 322.200 122.600 329.600 ;
        RECT 128.600 329.600 129.600 330.200 ;
        RECT 130.200 329.600 131.600 330.200 ;
        RECT 132.400 330.200 133.200 330.400 ;
        RECT 134.400 330.200 135.000 333.600 ;
        RECT 147.600 333.400 148.400 334.200 ;
        RECT 135.600 332.300 136.400 333.200 ;
        RECT 147.600 332.800 148.200 333.400 ;
        RECT 138.800 332.300 139.600 332.400 ;
        RECT 135.600 331.700 139.600 332.300 ;
        RECT 145.600 332.200 148.200 332.800 ;
        RECT 149.000 332.800 149.600 336.200 ;
        RECT 153.200 335.800 154.000 339.800 ;
        RECT 150.200 334.800 151.000 335.600 ;
        RECT 151.600 335.200 154.000 335.800 ;
        RECT 158.000 335.800 158.800 339.800 ;
        RECT 159.400 336.400 160.200 337.200 ;
        RECT 151.600 335.000 152.400 335.200 ;
        RECT 150.400 334.400 151.000 334.800 ;
        RECT 150.400 333.600 151.200 334.400 ;
        RECT 152.400 334.300 154.000 334.400 ;
        RECT 154.800 334.300 155.600 334.400 ;
        RECT 152.400 333.700 155.600 334.300 ;
        RECT 152.400 333.600 154.000 333.700 ;
        RECT 154.800 333.600 155.600 333.700 ;
        RECT 156.400 332.800 157.200 334.400 ;
        RECT 149.000 332.400 150.000 332.800 ;
        RECT 158.000 332.400 158.600 335.800 ;
        RECT 159.600 335.600 160.400 336.400 ;
        RECT 159.600 334.300 160.400 334.400 ;
        RECT 161.200 334.300 162.000 339.800 ;
        RECT 162.800 335.600 163.600 337.200 ;
        RECT 164.400 335.600 165.200 337.200 ;
        RECT 159.600 333.700 162.000 334.300 ;
        RECT 159.600 333.600 160.400 333.700 ;
        RECT 149.000 332.200 150.800 332.400 ;
        RECT 145.600 332.000 146.400 332.200 ;
        RECT 135.600 331.600 136.400 331.700 ;
        RECT 138.800 331.600 139.600 331.700 ;
        RECT 149.400 331.600 150.800 332.200 ;
        RECT 154.800 332.200 155.600 332.400 ;
        RECT 158.000 332.200 158.800 332.400 ;
        RECT 159.600 332.200 160.400 332.400 ;
        RECT 154.800 331.600 156.400 332.200 ;
        RECT 158.000 331.600 160.400 332.200 ;
        RECT 147.800 331.400 148.600 331.600 ;
        RECT 145.200 330.800 148.600 331.400 ;
        RECT 145.200 330.200 145.800 330.800 ;
        RECT 149.400 330.200 150.000 331.600 ;
        RECT 155.600 331.200 156.400 331.600 ;
        RECT 159.600 330.200 160.200 331.600 ;
        RECT 132.400 329.600 133.800 330.200 ;
        RECT 134.400 329.600 135.400 330.200 ;
        RECT 128.600 322.200 129.400 329.600 ;
        RECT 130.200 328.400 130.800 329.600 ;
        RECT 130.000 327.600 130.800 328.400 ;
        RECT 133.200 328.400 133.800 329.600 ;
        RECT 133.200 327.600 134.000 328.400 ;
        RECT 134.600 322.200 135.400 329.600 ;
        RECT 143.600 329.600 145.800 330.200 ;
        RECT 143.600 322.200 144.400 329.600 ;
        RECT 145.000 329.400 145.800 329.600 ;
        RECT 148.000 329.600 150.000 330.200 ;
        RECT 151.600 329.600 154.000 330.200 ;
        RECT 148.000 324.400 149.600 329.600 ;
        RECT 151.600 329.400 152.400 329.600 ;
        RECT 146.800 323.600 149.600 324.400 ;
        RECT 148.000 322.200 149.600 323.600 ;
        RECT 153.200 322.200 154.000 329.600 ;
        RECT 154.800 329.600 158.800 330.200 ;
        RECT 154.800 322.200 155.600 329.600 ;
        RECT 158.000 322.200 158.800 329.600 ;
        RECT 159.600 322.200 160.400 330.200 ;
        RECT 161.200 322.200 162.000 333.700 ;
        RECT 166.000 330.300 166.800 339.800 ;
        RECT 167.600 335.800 168.400 339.800 ;
        RECT 169.200 336.000 170.000 339.800 ;
        RECT 172.400 336.000 173.200 339.800 ;
        RECT 169.200 335.800 173.200 336.000 ;
        RECT 174.000 335.800 174.800 339.800 ;
        RECT 178.400 336.200 180.000 339.800 ;
        RECT 167.800 334.400 168.400 335.800 ;
        RECT 169.400 335.400 173.000 335.800 ;
        RECT 174.000 335.200 176.400 335.800 ;
        RECT 175.600 335.000 176.400 335.200 ;
        RECT 177.000 334.800 177.800 335.600 ;
        RECT 171.600 334.400 172.400 334.800 ;
        RECT 177.000 334.400 177.600 334.800 ;
        RECT 167.600 333.600 170.200 334.400 ;
        RECT 171.600 333.800 173.200 334.400 ;
        RECT 172.400 333.600 173.200 333.800 ;
        RECT 174.000 333.600 175.600 334.400 ;
        RECT 176.800 333.600 177.600 334.400 ;
        RECT 167.600 332.300 168.400 332.400 ;
        RECT 169.600 332.300 170.200 333.600 ;
        RECT 167.600 331.700 170.200 332.300 ;
        RECT 167.600 331.600 168.400 331.700 ;
        RECT 167.600 330.300 168.400 330.400 ;
        RECT 166.000 330.200 168.400 330.300 ;
        RECT 169.600 330.200 170.200 331.700 ;
        RECT 170.800 332.300 171.600 333.200 ;
        RECT 178.400 332.800 179.000 336.200 ;
        RECT 183.600 335.800 184.400 339.800 ;
        RECT 179.600 335.400 181.200 335.600 ;
        RECT 179.600 334.800 181.600 335.400 ;
        RECT 182.200 335.200 184.400 335.800 ;
        RECT 186.800 335.200 187.600 339.800 ;
        RECT 190.000 335.200 190.800 339.800 ;
        RECT 193.200 335.200 194.000 339.800 ;
        RECT 196.400 335.200 197.200 339.800 ;
        RECT 182.200 335.000 183.000 335.200 ;
        RECT 181.000 334.400 181.600 334.800 ;
        RECT 185.200 334.400 187.600 335.200 ;
        RECT 188.600 334.400 190.800 335.200 ;
        RECT 191.800 334.400 194.000 335.200 ;
        RECT 195.400 334.400 197.200 335.200 ;
        RECT 199.600 335.400 200.400 339.800 ;
        RECT 203.800 338.400 205.000 339.800 ;
        RECT 203.800 337.800 205.200 338.400 ;
        RECT 208.400 337.800 209.200 339.800 ;
        RECT 212.800 338.400 213.600 339.800 ;
        RECT 212.800 337.800 214.800 338.400 ;
        RECT 204.400 337.000 205.200 337.800 ;
        RECT 208.600 337.200 209.200 337.800 ;
        RECT 208.600 336.600 211.400 337.200 ;
        RECT 210.600 336.400 211.400 336.600 ;
        RECT 212.400 336.400 213.200 337.200 ;
        RECT 214.000 337.000 214.800 337.800 ;
        RECT 202.600 335.400 203.400 335.600 ;
        RECT 199.600 334.800 203.400 335.400 ;
        RECT 179.600 333.400 180.400 334.200 ;
        RECT 181.000 333.800 184.400 334.400 ;
        RECT 182.800 333.600 184.400 333.800 ;
        RECT 178.000 332.400 179.000 332.800 ;
        RECT 177.200 332.300 179.000 332.400 ;
        RECT 170.800 332.200 179.000 332.300 ;
        RECT 179.800 332.800 180.400 333.400 ;
        RECT 179.800 332.200 182.400 332.800 ;
        RECT 170.800 331.700 178.600 332.200 ;
        RECT 181.600 332.000 182.400 332.200 ;
        RECT 170.800 331.600 171.600 331.700 ;
        RECT 177.200 331.600 178.600 331.700 ;
        RECT 185.200 331.600 186.000 334.400 ;
        RECT 188.600 333.800 189.400 334.400 ;
        RECT 191.800 333.800 192.600 334.400 ;
        RECT 195.400 333.800 196.200 334.400 ;
        RECT 186.800 333.000 189.400 333.800 ;
        RECT 190.200 333.000 192.600 333.800 ;
        RECT 193.600 333.000 196.200 333.800 ;
        RECT 188.600 331.600 189.400 333.000 ;
        RECT 191.800 331.600 192.600 333.000 ;
        RECT 195.400 331.600 196.200 333.000 ;
        RECT 178.000 330.200 178.600 331.600 ;
        RECT 179.400 331.400 180.200 331.600 ;
        RECT 179.400 330.800 182.800 331.400 ;
        RECT 185.200 330.800 187.600 331.600 ;
        RECT 188.600 330.800 190.800 331.600 ;
        RECT 191.800 330.800 194.000 331.600 ;
        RECT 195.400 330.800 197.200 331.600 ;
        RECT 182.200 330.200 182.800 330.800 ;
        RECT 166.000 329.700 169.000 330.200 ;
        RECT 166.000 322.200 166.800 329.700 ;
        RECT 167.600 329.600 169.000 329.700 ;
        RECT 169.600 329.600 170.600 330.200 ;
        RECT 168.400 328.400 169.000 329.600 ;
        RECT 168.400 327.600 169.200 328.400 ;
        RECT 169.800 322.200 170.600 329.600 ;
        RECT 174.000 329.600 176.400 330.200 ;
        RECT 178.000 329.600 180.000 330.200 ;
        RECT 174.000 322.200 174.800 329.600 ;
        RECT 175.600 329.400 176.400 329.600 ;
        RECT 178.400 322.200 180.000 329.600 ;
        RECT 182.200 329.600 184.400 330.200 ;
        RECT 182.200 329.400 183.000 329.600 ;
        RECT 183.600 322.200 184.400 329.600 ;
        RECT 186.800 322.200 187.600 330.800 ;
        RECT 190.000 322.200 190.800 330.800 ;
        RECT 193.200 322.200 194.000 330.800 ;
        RECT 196.400 322.200 197.200 330.800 ;
        RECT 199.600 331.400 200.400 334.800 ;
        RECT 206.600 334.200 207.400 334.400 ;
        RECT 210.800 334.200 211.600 334.400 ;
        RECT 212.400 334.200 213.000 336.400 ;
        RECT 217.200 335.000 218.000 339.800 ;
        RECT 218.800 335.800 219.600 339.800 ;
        RECT 223.200 336.200 224.800 339.800 ;
        RECT 218.800 335.200 221.200 335.800 ;
        RECT 220.400 335.000 221.200 335.200 ;
        RECT 221.800 334.800 222.600 335.600 ;
        RECT 221.800 334.400 222.400 334.800 ;
        RECT 215.600 334.200 217.200 334.400 ;
        RECT 206.200 333.600 217.200 334.200 ;
        RECT 218.800 333.600 220.400 334.400 ;
        RECT 221.600 333.600 222.400 334.400 ;
        RECT 204.400 332.800 205.200 333.000 ;
        RECT 201.400 332.200 205.200 332.800 ;
        RECT 201.400 332.000 202.200 332.200 ;
        RECT 203.000 331.400 203.800 331.600 ;
        RECT 199.600 330.800 203.800 331.400 ;
        RECT 199.600 322.200 200.400 330.800 ;
        RECT 206.200 330.400 206.800 333.600 ;
        RECT 213.400 333.400 214.200 333.600 ;
        RECT 223.200 332.800 223.800 336.200 ;
        RECT 228.400 335.800 229.200 339.800 ;
        RECT 224.400 335.400 226.000 335.600 ;
        RECT 224.400 334.800 226.400 335.400 ;
        RECT 227.000 335.200 229.200 335.800 ;
        RECT 230.000 335.800 230.800 339.800 ;
        RECT 234.400 338.400 236.000 339.800 ;
        RECT 233.200 337.600 236.000 338.400 ;
        RECT 234.400 336.200 236.000 337.600 ;
        RECT 230.000 335.200 232.400 335.800 ;
        RECT 227.000 335.000 227.800 335.200 ;
        RECT 231.600 335.000 232.400 335.200 ;
        RECT 225.800 334.400 226.400 334.800 ;
        RECT 233.000 334.800 233.800 335.600 ;
        RECT 233.000 334.400 233.600 334.800 ;
        RECT 224.400 333.400 225.200 334.200 ;
        RECT 225.800 333.800 229.200 334.400 ;
        RECT 227.600 333.600 229.200 333.800 ;
        RECT 230.000 333.600 231.600 334.400 ;
        RECT 232.800 333.600 233.600 334.400 ;
        RECT 234.400 334.200 235.000 336.200 ;
        RECT 239.600 335.800 240.400 339.800 ;
        RECT 241.200 335.800 242.000 339.800 ;
        RECT 242.800 336.000 243.600 339.800 ;
        RECT 246.000 336.000 246.800 339.800 ;
        RECT 242.800 335.800 246.800 336.000 ;
        RECT 248.200 336.400 249.000 339.800 ;
        RECT 248.200 335.800 250.000 336.400 ;
        RECT 235.600 334.800 237.200 335.600 ;
        RECT 237.800 335.200 240.400 335.800 ;
        RECT 237.800 335.000 238.600 335.200 ;
        RECT 241.400 334.400 242.000 335.800 ;
        RECT 243.000 335.400 246.600 335.800 ;
        RECT 245.200 334.400 246.000 334.800 ;
        RECT 238.800 334.200 240.400 334.400 ;
        RECT 234.400 333.600 235.400 334.200 ;
        RECT 238.200 334.000 240.400 334.200 ;
        RECT 212.400 332.400 213.200 332.600 ;
        RECT 215.000 332.400 215.800 332.600 ;
        RECT 222.800 332.400 223.800 332.800 ;
        RECT 210.800 331.800 215.800 332.400 ;
        RECT 218.800 332.300 219.600 332.400 ;
        RECT 222.000 332.300 223.800 332.400 ;
        RECT 218.800 332.200 223.800 332.300 ;
        RECT 224.600 332.800 225.200 333.400 ;
        RECT 224.600 332.200 227.200 332.800 ;
        RECT 210.800 331.600 211.600 331.800 ;
        RECT 218.800 331.700 223.400 332.200 ;
        RECT 226.400 332.000 227.200 332.200 ;
        RECT 234.800 332.400 235.400 333.600 ;
        RECT 236.000 333.600 240.400 334.000 ;
        RECT 241.200 333.600 243.800 334.400 ;
        RECT 245.200 333.800 246.800 334.400 ;
        RECT 246.000 333.600 246.800 333.800 ;
        RECT 236.000 333.400 238.800 333.600 ;
        RECT 236.000 333.200 236.800 333.400 ;
        RECT 218.800 331.600 219.600 331.700 ;
        RECT 222.000 331.600 223.400 331.700 ;
        RECT 234.800 331.600 235.600 332.400 ;
        RECT 237.400 332.200 238.200 332.400 ;
        RECT 236.600 331.600 238.200 332.200 ;
        RECT 212.400 331.000 218.000 331.200 ;
        RECT 212.200 330.800 218.000 331.000 ;
        RECT 204.400 329.800 206.800 330.400 ;
        RECT 208.200 330.600 218.000 330.800 ;
        RECT 208.200 330.200 213.000 330.600 ;
        RECT 204.400 328.800 205.000 329.800 ;
        RECT 203.600 328.000 205.000 328.800 ;
        RECT 206.600 329.000 207.400 329.200 ;
        RECT 208.200 329.000 208.800 330.200 ;
        RECT 206.600 328.400 208.800 329.000 ;
        RECT 209.400 329.000 214.800 329.600 ;
        RECT 209.400 328.800 210.200 329.000 ;
        RECT 214.000 328.800 214.800 329.000 ;
        RECT 207.800 327.400 208.600 327.600 ;
        RECT 210.600 327.400 211.400 327.600 ;
        RECT 204.400 326.200 205.200 327.000 ;
        RECT 207.800 326.800 211.400 327.400 ;
        RECT 208.600 326.200 209.200 326.800 ;
        RECT 214.000 326.200 214.800 327.000 ;
        RECT 203.800 322.200 205.000 326.200 ;
        RECT 208.400 322.200 209.200 326.200 ;
        RECT 212.800 325.600 214.800 326.200 ;
        RECT 212.800 322.200 213.600 325.600 ;
        RECT 217.200 322.200 218.000 330.600 ;
        RECT 222.800 330.200 223.400 331.600 ;
        RECT 224.200 331.400 225.000 331.600 ;
        RECT 224.200 330.800 227.600 331.400 ;
        RECT 227.000 330.200 227.600 330.800 ;
        RECT 234.800 330.200 235.400 331.600 ;
        RECT 236.600 331.400 237.400 331.600 ;
        RECT 241.200 330.200 242.000 330.400 ;
        RECT 243.200 330.200 243.800 333.600 ;
        RECT 244.400 331.600 245.200 333.200 ;
        RECT 218.800 329.600 221.200 330.200 ;
        RECT 222.800 329.600 224.800 330.200 ;
        RECT 218.800 322.200 219.600 329.600 ;
        RECT 220.400 329.400 221.200 329.600 ;
        RECT 223.200 322.200 224.800 329.600 ;
        RECT 227.000 329.600 229.200 330.200 ;
        RECT 227.000 329.400 227.800 329.600 ;
        RECT 228.400 322.200 229.200 329.600 ;
        RECT 230.000 329.600 232.400 330.200 ;
        RECT 230.000 322.200 230.800 329.600 ;
        RECT 231.600 329.400 232.400 329.600 ;
        RECT 234.400 322.200 236.000 330.200 ;
        RECT 237.800 329.600 240.400 330.200 ;
        RECT 241.200 329.600 242.600 330.200 ;
        RECT 243.200 329.600 244.200 330.200 ;
        RECT 237.800 329.400 238.600 329.600 ;
        RECT 239.600 322.200 240.400 329.600 ;
        RECT 242.000 328.400 242.600 329.600 ;
        RECT 242.000 327.600 242.800 328.400 ;
        RECT 243.400 324.400 244.200 329.600 ;
        RECT 247.600 328.800 248.400 330.400 ;
        RECT 249.200 328.300 250.000 335.800 ;
        RECT 250.800 333.600 251.600 335.200 ;
        RECT 256.000 334.200 256.800 339.800 ;
        RECT 259.400 336.400 260.200 339.800 ;
        RECT 259.400 335.800 261.200 336.400 ;
        RECT 256.000 333.800 257.800 334.200 ;
        RECT 256.200 333.600 257.800 333.800 ;
        RECT 254.000 331.600 255.600 332.400 ;
        RECT 250.800 330.300 251.600 330.400 ;
        RECT 252.400 330.300 253.200 331.200 ;
        RECT 250.800 329.700 253.200 330.300 ;
        RECT 250.800 329.600 251.600 329.700 ;
        RECT 252.400 329.600 253.200 329.700 ;
        RECT 257.200 330.400 257.800 333.600 ;
        RECT 257.200 330.300 258.000 330.400 ;
        RECT 258.800 330.300 259.600 330.400 ;
        RECT 257.200 329.700 259.600 330.300 ;
        RECT 257.200 329.600 258.000 329.700 ;
        RECT 254.000 328.300 254.800 328.400 ;
        RECT 249.200 327.700 254.800 328.300 ;
        RECT 243.400 323.600 245.200 324.400 ;
        RECT 243.400 322.200 244.200 323.600 ;
        RECT 249.200 322.200 250.000 327.700 ;
        RECT 254.000 327.600 254.800 327.700 ;
        RECT 255.600 327.600 256.400 329.200 ;
        RECT 257.200 327.000 257.800 329.600 ;
        RECT 258.800 328.800 259.600 329.700 ;
        RECT 254.200 326.400 257.800 327.000 ;
        RECT 254.200 326.200 254.800 326.400 ;
        RECT 254.000 322.200 254.800 326.200 ;
        RECT 257.200 326.200 257.800 326.400 ;
        RECT 257.200 322.200 258.000 326.200 ;
        RECT 260.400 322.200 261.200 335.800 ;
        RECT 266.800 335.800 267.600 339.800 ;
        RECT 271.600 337.800 272.400 339.800 ;
        RECT 268.200 336.400 269.000 337.200 ;
        RECT 262.000 333.600 262.800 335.200 ;
        RECT 265.200 332.800 266.000 334.400 ;
        RECT 263.600 332.200 264.400 332.400 ;
        RECT 266.800 332.200 267.400 335.800 ;
        RECT 268.400 335.600 269.200 336.400 ;
        RECT 270.000 335.600 270.800 337.200 ;
        RECT 271.800 336.300 272.400 337.800 ;
        RECT 273.200 336.300 274.000 336.400 ;
        RECT 271.700 335.700 274.000 336.300 ;
        RECT 274.800 336.000 275.600 339.800 ;
        RECT 278.000 336.000 278.800 339.800 ;
        RECT 274.800 335.800 278.800 336.000 ;
        RECT 279.600 335.800 280.400 339.800 ;
        RECT 271.800 334.400 272.400 335.700 ;
        RECT 273.200 335.600 274.000 335.700 ;
        RECT 275.000 335.400 278.600 335.800 ;
        RECT 275.600 334.400 276.400 334.800 ;
        RECT 279.600 334.400 280.200 335.800 ;
        RECT 281.200 335.600 282.000 337.200 ;
        RECT 271.600 333.600 272.400 334.400 ;
        RECT 274.800 333.800 276.400 334.400 ;
        RECT 274.800 333.600 275.600 333.800 ;
        RECT 277.800 333.600 280.400 334.400 ;
        RECT 282.800 334.300 283.600 339.800 ;
        RECT 287.600 335.800 288.400 339.800 ;
        RECT 297.200 337.800 298.000 339.800 ;
        RECT 289.000 336.400 289.800 337.200 ;
        RECT 289.200 336.300 290.000 336.400 ;
        RECT 297.200 336.300 297.800 337.800 ;
        RECT 286.000 334.300 286.800 334.400 ;
        RECT 282.800 333.700 286.800 334.300 ;
        RECT 268.400 332.200 269.200 332.400 ;
        RECT 263.600 331.600 265.200 332.200 ;
        RECT 266.800 331.600 269.200 332.200 ;
        RECT 264.400 331.200 265.200 331.600 ;
        RECT 268.400 330.200 269.000 331.600 ;
        RECT 271.800 330.200 272.400 333.600 ;
        RECT 273.200 332.300 274.000 332.400 ;
        RECT 276.400 332.300 277.200 333.200 ;
        RECT 273.200 331.700 277.200 332.300 ;
        RECT 273.200 330.800 274.000 331.700 ;
        RECT 276.400 331.600 277.200 331.700 ;
        RECT 277.800 330.200 278.400 333.600 ;
        RECT 279.600 330.200 280.400 330.400 ;
        RECT 263.600 329.600 267.600 330.200 ;
        RECT 263.600 322.200 264.400 329.600 ;
        RECT 266.800 322.200 267.600 329.600 ;
        RECT 268.400 322.200 269.200 330.200 ;
        RECT 271.600 329.400 273.400 330.200 ;
        RECT 272.600 322.200 273.400 329.400 ;
        RECT 277.400 329.600 278.400 330.200 ;
        RECT 279.000 329.600 280.400 330.200 ;
        RECT 277.400 326.400 278.200 329.600 ;
        RECT 279.000 328.400 279.600 329.600 ;
        RECT 278.800 327.600 279.600 328.400 ;
        RECT 276.400 325.600 278.200 326.400 ;
        RECT 277.400 322.200 278.200 325.600 ;
        RECT 282.800 322.200 283.600 333.700 ;
        RECT 286.000 332.800 286.800 333.700 ;
        RECT 284.400 332.200 285.200 332.400 ;
        RECT 287.600 332.200 288.200 335.800 ;
        RECT 289.200 335.700 297.900 336.300 ;
        RECT 289.200 335.600 290.000 335.700 ;
        RECT 297.200 334.400 297.800 335.700 ;
        RECT 298.800 335.600 299.600 337.200 ;
        RECT 300.400 336.000 301.200 339.800 ;
        RECT 303.600 336.000 304.400 339.800 ;
        RECT 300.400 335.800 304.400 336.000 ;
        RECT 305.200 335.800 306.000 339.800 ;
        RECT 309.400 336.400 310.200 339.800 ;
        RECT 311.800 336.400 312.600 337.200 ;
        RECT 308.400 335.800 310.200 336.400 ;
        RECT 300.600 335.400 304.200 335.800 ;
        RECT 301.200 334.400 302.000 334.800 ;
        RECT 305.200 334.400 305.800 335.800 ;
        RECT 297.200 333.600 298.000 334.400 ;
        RECT 300.400 333.800 302.000 334.400 ;
        RECT 300.400 333.600 301.200 333.800 ;
        RECT 303.400 333.600 306.000 334.400 ;
        RECT 306.800 333.600 307.600 335.200 ;
        RECT 289.200 332.200 290.000 332.400 ;
        RECT 284.400 331.600 286.000 332.200 ;
        RECT 287.600 331.600 290.000 332.200 ;
        RECT 285.200 331.200 286.000 331.600 ;
        RECT 289.200 330.200 289.800 331.600 ;
        RECT 295.600 330.800 296.400 332.400 ;
        RECT 297.200 330.200 297.800 333.600 ;
        RECT 302.000 331.600 302.800 333.200 ;
        RECT 303.400 330.200 304.000 333.600 ;
        RECT 305.200 330.300 306.000 330.400 ;
        RECT 308.400 330.300 309.200 335.800 ;
        RECT 311.600 335.600 312.400 336.400 ;
        RECT 313.200 335.800 314.000 339.800 ;
        RECT 319.600 337.800 320.400 339.800 ;
        RECT 311.600 332.200 312.400 332.400 ;
        RECT 313.400 332.200 314.000 335.800 ;
        RECT 318.000 335.600 318.800 337.200 ;
        RECT 319.800 334.400 320.400 337.800 ;
        RECT 322.800 335.800 323.600 339.800 ;
        RECT 327.200 336.200 328.800 339.800 ;
        RECT 322.800 335.200 325.000 335.800 ;
        RECT 326.000 335.400 327.600 335.600 ;
        RECT 324.200 335.000 325.000 335.200 ;
        RECT 325.600 334.800 327.600 335.400 ;
        RECT 325.600 334.400 326.200 334.800 ;
        RECT 314.800 332.800 315.600 334.400 ;
        RECT 319.600 333.600 320.400 334.400 ;
        RECT 322.800 333.800 326.200 334.400 ;
        RECT 322.800 333.600 324.400 333.800 ;
        RECT 316.400 332.300 317.200 332.400 ;
        RECT 319.800 332.300 320.400 333.600 ;
        RECT 326.800 333.400 327.600 334.200 ;
        RECT 326.800 332.800 327.400 333.400 ;
        RECT 316.400 332.200 320.400 332.300 ;
        RECT 311.600 331.600 314.000 332.200 ;
        RECT 315.600 331.700 320.400 332.200 ;
        RECT 315.600 331.600 317.200 331.700 ;
        RECT 305.200 330.200 309.200 330.300 ;
        RECT 284.400 329.600 288.400 330.200 ;
        RECT 284.400 322.200 285.200 329.600 ;
        RECT 287.600 322.200 288.400 329.600 ;
        RECT 289.200 322.200 290.000 330.200 ;
        RECT 296.200 329.400 298.000 330.200 ;
        RECT 303.000 329.600 304.000 330.200 ;
        RECT 304.600 329.700 309.200 330.200 ;
        RECT 304.600 329.600 306.000 329.700 ;
        RECT 296.200 322.200 297.000 329.400 ;
        RECT 303.000 328.400 303.800 329.600 ;
        RECT 304.600 328.400 305.200 329.600 ;
        RECT 302.000 327.600 303.800 328.400 ;
        RECT 304.400 327.600 305.200 328.400 ;
        RECT 303.000 322.200 303.800 327.600 ;
        RECT 308.400 322.200 309.200 329.700 ;
        RECT 310.000 330.300 310.800 330.400 ;
        RECT 311.800 330.300 312.400 331.600 ;
        RECT 315.600 331.200 316.400 331.600 ;
        RECT 310.000 329.700 312.400 330.300 ;
        RECT 319.800 330.200 320.400 331.700 ;
        RECT 321.200 330.800 322.000 332.400 ;
        RECT 324.800 332.200 327.400 332.800 ;
        RECT 328.200 332.800 328.800 336.200 ;
        RECT 332.400 335.800 333.200 339.800 ;
        RECT 329.400 334.800 330.200 335.600 ;
        RECT 330.800 335.200 333.200 335.800 ;
        RECT 334.000 335.400 334.800 339.800 ;
        RECT 338.200 338.400 339.400 339.800 ;
        RECT 338.200 337.800 339.600 338.400 ;
        RECT 342.800 337.800 343.600 339.800 ;
        RECT 347.200 338.400 348.000 339.800 ;
        RECT 347.200 337.800 349.200 338.400 ;
        RECT 338.800 337.000 339.600 337.800 ;
        RECT 343.000 337.200 343.600 337.800 ;
        RECT 343.000 336.600 345.800 337.200 ;
        RECT 345.000 336.400 345.800 336.600 ;
        RECT 346.800 336.400 347.600 337.200 ;
        RECT 348.400 337.000 349.200 337.800 ;
        RECT 337.000 335.400 337.800 335.600 ;
        RECT 330.800 335.000 331.600 335.200 ;
        RECT 329.600 334.400 330.200 334.800 ;
        RECT 334.000 334.800 337.800 335.400 ;
        RECT 329.600 333.600 330.400 334.400 ;
        RECT 331.600 333.600 333.200 334.400 ;
        RECT 328.200 332.400 329.200 332.800 ;
        RECT 328.200 332.200 330.000 332.400 ;
        RECT 324.800 332.000 325.600 332.200 ;
        RECT 328.600 331.600 330.000 332.200 ;
        RECT 327.000 331.400 327.800 331.600 ;
        RECT 324.400 330.800 327.800 331.400 ;
        RECT 324.400 330.200 325.000 330.800 ;
        RECT 328.600 330.200 329.200 331.600 ;
        RECT 334.000 331.400 334.800 334.800 ;
        RECT 341.000 334.200 341.800 334.400 ;
        RECT 345.200 334.200 346.000 334.400 ;
        RECT 346.800 334.200 347.400 336.400 ;
        RECT 351.600 335.000 352.400 339.800 ;
        RECT 350.000 334.200 351.600 334.400 ;
        RECT 340.600 333.600 351.600 334.200 ;
        RECT 338.800 332.800 339.600 333.000 ;
        RECT 335.800 332.200 339.600 332.800 ;
        RECT 340.600 332.400 341.200 333.600 ;
        RECT 347.800 333.400 348.600 333.600 ;
        RECT 346.800 332.400 347.600 332.600 ;
        RECT 349.400 332.400 350.200 332.600 ;
        RECT 335.800 332.000 336.600 332.200 ;
        RECT 340.400 331.600 341.200 332.400 ;
        RECT 345.200 331.800 350.200 332.400 ;
        RECT 345.200 331.600 346.000 331.800 ;
        RECT 337.400 331.400 338.200 331.600 ;
        RECT 334.000 330.800 338.200 331.400 ;
        RECT 310.000 328.800 310.800 329.700 ;
        RECT 311.600 322.200 312.400 329.700 ;
        RECT 313.200 329.600 317.200 330.200 ;
        RECT 313.200 322.200 314.000 329.600 ;
        RECT 316.400 322.200 317.200 329.600 ;
        RECT 319.600 329.400 321.400 330.200 ;
        RECT 320.600 322.200 321.400 329.400 ;
        RECT 322.800 329.600 325.000 330.200 ;
        RECT 322.800 322.200 323.600 329.600 ;
        RECT 324.200 329.400 325.000 329.600 ;
        RECT 327.200 329.600 329.200 330.200 ;
        RECT 330.800 329.600 333.200 330.200 ;
        RECT 327.200 324.400 328.800 329.600 ;
        RECT 330.800 329.400 331.600 329.600 ;
        RECT 326.000 323.600 328.800 324.400 ;
        RECT 327.200 322.200 328.800 323.600 ;
        RECT 332.400 322.200 333.200 329.600 ;
        RECT 334.000 322.200 334.800 330.800 ;
        RECT 340.600 330.400 341.200 331.600 ;
        RECT 346.800 331.000 352.400 331.200 ;
        RECT 346.600 330.800 352.400 331.000 ;
        RECT 338.800 329.800 341.200 330.400 ;
        RECT 342.600 330.600 352.400 330.800 ;
        RECT 342.600 330.200 347.400 330.600 ;
        RECT 338.800 328.800 339.400 329.800 ;
        RECT 338.000 328.000 339.400 328.800 ;
        RECT 341.000 329.000 341.800 329.200 ;
        RECT 342.600 329.000 343.200 330.200 ;
        RECT 341.000 328.400 343.200 329.000 ;
        RECT 343.800 329.000 349.200 329.600 ;
        RECT 343.800 328.800 344.600 329.000 ;
        RECT 348.400 328.800 349.200 329.000 ;
        RECT 342.200 327.400 343.000 327.600 ;
        RECT 345.000 327.400 345.800 327.600 ;
        RECT 338.800 326.200 339.600 327.000 ;
        RECT 342.200 326.800 345.800 327.400 ;
        RECT 343.000 326.200 343.600 326.800 ;
        RECT 348.400 326.200 349.200 327.000 ;
        RECT 338.200 322.200 339.400 326.200 ;
        RECT 342.800 322.200 343.600 326.200 ;
        RECT 347.200 325.600 349.200 326.200 ;
        RECT 347.200 322.200 348.000 325.600 ;
        RECT 351.600 322.200 352.400 330.600 ;
        RECT 353.200 322.200 354.000 339.800 ;
        RECT 354.800 335.600 355.600 337.200 ;
        RECT 356.400 335.400 357.200 339.800 ;
        RECT 360.600 338.400 361.800 339.800 ;
        RECT 360.600 337.800 362.000 338.400 ;
        RECT 365.200 337.800 366.000 339.800 ;
        RECT 369.600 338.400 370.400 339.800 ;
        RECT 369.600 337.800 371.600 338.400 ;
        RECT 361.200 337.000 362.000 337.800 ;
        RECT 365.400 337.200 366.000 337.800 ;
        RECT 365.400 336.600 368.200 337.200 ;
        RECT 367.400 336.400 368.200 336.600 ;
        RECT 369.200 336.400 370.000 337.200 ;
        RECT 370.800 337.000 371.600 337.800 ;
        RECT 359.400 335.400 360.200 335.600 ;
        RECT 356.400 334.800 360.200 335.400 ;
        RECT 356.400 331.400 357.200 334.800 ;
        RECT 363.400 334.200 364.200 334.400 ;
        RECT 367.600 334.200 368.400 334.400 ;
        RECT 369.200 334.200 369.800 336.400 ;
        RECT 374.000 335.000 374.800 339.800 ;
        RECT 375.600 336.000 376.400 339.800 ;
        RECT 378.800 339.200 382.800 339.800 ;
        RECT 378.800 336.000 379.600 339.200 ;
        RECT 375.600 335.800 379.600 336.000 ;
        RECT 380.400 335.800 381.200 338.600 ;
        RECT 382.000 335.800 382.800 339.200 ;
        RECT 383.600 335.800 384.400 339.800 ;
        RECT 385.200 336.000 386.000 339.800 ;
        RECT 388.400 336.000 389.200 339.800 ;
        RECT 392.600 336.400 393.400 339.800 ;
        RECT 385.200 335.800 389.200 336.000 ;
        RECT 391.600 335.800 393.400 336.400 ;
        RECT 375.800 335.400 379.400 335.800 ;
        RECT 376.400 334.400 377.200 334.800 ;
        RECT 380.600 334.400 381.200 335.800 ;
        RECT 383.800 334.400 384.400 335.800 ;
        RECT 385.400 335.400 389.000 335.800 ;
        RECT 387.600 334.400 388.400 334.800 ;
        RECT 372.400 334.200 374.000 334.400 ;
        RECT 363.000 333.600 374.000 334.200 ;
        RECT 375.600 333.800 377.200 334.400 ;
        RECT 378.800 333.800 381.200 334.400 ;
        RECT 375.600 333.600 376.400 333.800 ;
        RECT 378.800 333.600 379.600 333.800 ;
        RECT 361.200 332.800 362.000 333.000 ;
        RECT 358.200 332.200 362.000 332.800 ;
        RECT 358.200 332.000 359.000 332.200 ;
        RECT 359.800 331.400 360.600 331.600 ;
        RECT 356.400 330.800 360.600 331.400 ;
        RECT 356.400 322.200 357.200 330.800 ;
        RECT 363.000 330.400 363.600 333.600 ;
        RECT 370.200 333.400 371.000 333.600 ;
        RECT 369.200 332.400 370.000 332.600 ;
        RECT 371.800 332.400 372.600 332.600 ;
        RECT 367.600 331.800 372.600 332.400 ;
        RECT 367.600 331.600 368.400 331.800 ;
        RECT 377.200 331.600 378.000 333.200 ;
        RECT 369.200 331.000 374.800 331.200 ;
        RECT 369.000 330.800 374.800 331.000 ;
        RECT 361.200 329.800 363.600 330.400 ;
        RECT 365.000 330.600 374.800 330.800 ;
        RECT 365.000 330.200 369.800 330.600 ;
        RECT 361.200 328.800 361.800 329.800 ;
        RECT 360.400 328.000 361.800 328.800 ;
        RECT 363.400 329.000 364.200 329.200 ;
        RECT 365.000 329.000 365.600 330.200 ;
        RECT 363.400 328.400 365.600 329.000 ;
        RECT 366.200 329.000 371.600 329.600 ;
        RECT 366.200 328.800 367.000 329.000 ;
        RECT 370.800 328.800 371.600 329.000 ;
        RECT 364.600 327.400 365.400 327.600 ;
        RECT 367.400 327.400 368.200 327.600 ;
        RECT 361.200 326.200 362.000 327.000 ;
        RECT 364.600 326.800 368.200 327.400 ;
        RECT 365.400 326.200 366.000 326.800 ;
        RECT 370.800 326.200 371.600 327.000 ;
        RECT 360.600 322.200 361.800 326.200 ;
        RECT 365.200 322.200 366.000 326.200 ;
        RECT 369.600 325.600 371.600 326.200 ;
        RECT 369.600 322.200 370.400 325.600 ;
        RECT 374.000 322.200 374.800 330.600 ;
        RECT 378.800 330.200 379.400 333.600 ;
        RECT 380.400 331.600 381.200 333.200 ;
        RECT 382.000 332.800 382.800 334.400 ;
        RECT 383.600 333.600 386.200 334.400 ;
        RECT 387.600 333.800 389.200 334.400 ;
        RECT 388.400 333.600 389.200 333.800 ;
        RECT 390.000 333.600 390.800 335.200 ;
        RECT 385.600 332.400 386.200 333.600 ;
        RECT 385.200 331.600 386.200 332.400 ;
        RECT 386.800 332.300 387.600 333.200 ;
        RECT 391.600 332.300 392.400 335.800 ;
        RECT 386.800 331.700 392.400 332.300 ;
        RECT 386.800 331.600 387.600 331.700 ;
        RECT 383.600 330.200 384.400 330.400 ;
        RECT 385.600 330.200 386.200 331.600 ;
        RECT 378.200 324.400 380.200 330.200 ;
        RECT 383.600 329.600 385.000 330.200 ;
        RECT 385.600 329.600 386.600 330.200 ;
        RECT 384.400 328.400 385.000 329.600 ;
        RECT 384.400 327.600 385.200 328.400 ;
        RECT 377.200 323.600 380.200 324.400 ;
        RECT 378.200 322.200 380.200 323.600 ;
        RECT 385.800 322.200 386.600 329.600 ;
        RECT 391.600 322.200 392.400 331.700 ;
        RECT 394.800 335.400 395.600 339.800 ;
        RECT 399.000 338.400 400.200 339.800 ;
        RECT 399.000 337.800 400.400 338.400 ;
        RECT 403.600 337.800 404.400 339.800 ;
        RECT 408.000 338.400 408.800 339.800 ;
        RECT 408.000 337.800 410.000 338.400 ;
        RECT 399.600 337.000 400.400 337.800 ;
        RECT 403.800 337.200 404.400 337.800 ;
        RECT 403.800 336.600 406.600 337.200 ;
        RECT 405.800 336.400 406.600 336.600 ;
        RECT 407.600 336.400 408.400 337.200 ;
        RECT 409.200 337.000 410.000 337.800 ;
        RECT 397.800 335.400 398.600 335.600 ;
        RECT 394.800 334.800 398.600 335.400 ;
        RECT 394.800 331.400 395.600 334.800 ;
        RECT 401.800 334.200 402.600 334.400 ;
        RECT 407.600 334.200 408.200 336.400 ;
        RECT 412.400 335.000 413.200 339.800 ;
        RECT 414.000 335.400 414.800 339.800 ;
        RECT 418.200 338.400 419.400 339.800 ;
        RECT 418.200 337.800 419.600 338.400 ;
        RECT 422.800 337.800 423.600 339.800 ;
        RECT 427.200 338.400 428.000 339.800 ;
        RECT 427.200 337.800 429.200 338.400 ;
        RECT 418.800 337.000 419.600 337.800 ;
        RECT 423.000 337.200 423.600 337.800 ;
        RECT 423.000 336.600 425.800 337.200 ;
        RECT 425.000 336.400 425.800 336.600 ;
        RECT 426.800 336.400 427.600 337.200 ;
        RECT 428.400 337.000 429.200 337.800 ;
        RECT 417.000 335.400 417.800 335.600 ;
        RECT 414.000 334.800 417.800 335.400 ;
        RECT 410.800 334.200 412.400 334.400 ;
        RECT 401.400 333.600 412.400 334.200 ;
        RECT 399.600 332.800 400.400 333.000 ;
        RECT 396.600 332.200 400.400 332.800 ;
        RECT 401.400 332.300 402.000 333.600 ;
        RECT 408.600 333.400 409.400 333.600 ;
        RECT 407.600 332.400 408.400 332.600 ;
        RECT 410.200 332.400 411.000 332.600 ;
        RECT 402.800 332.300 403.600 332.400 ;
        RECT 396.600 332.000 397.400 332.200 ;
        RECT 401.300 331.700 403.600 332.300 ;
        RECT 398.200 331.400 399.000 331.600 ;
        RECT 394.800 330.800 399.000 331.400 ;
        RECT 393.200 328.800 394.000 330.400 ;
        RECT 394.800 322.200 395.600 330.800 ;
        RECT 401.400 330.400 402.000 331.700 ;
        RECT 402.800 331.600 403.600 331.700 ;
        RECT 406.000 331.800 411.000 332.400 ;
        RECT 406.000 331.600 406.800 331.800 ;
        RECT 414.000 331.400 414.800 334.800 ;
        RECT 421.000 334.200 421.800 334.400 ;
        RECT 423.600 334.200 424.400 334.400 ;
        RECT 426.800 334.200 427.400 336.400 ;
        RECT 431.600 335.000 432.400 339.800 ;
        RECT 433.200 335.800 434.000 339.800 ;
        RECT 437.600 336.200 439.200 339.800 ;
        RECT 433.200 335.200 435.400 335.800 ;
        RECT 436.400 335.400 438.000 335.600 ;
        RECT 434.600 335.000 435.400 335.200 ;
        RECT 436.000 334.800 438.000 335.400 ;
        RECT 436.000 334.400 436.600 334.800 ;
        RECT 430.000 334.200 431.600 334.400 ;
        RECT 420.600 333.600 431.600 334.200 ;
        RECT 433.200 333.800 436.600 334.400 ;
        RECT 433.200 333.600 434.800 333.800 ;
        RECT 418.800 332.800 419.600 333.000 ;
        RECT 415.800 332.200 419.600 332.800 ;
        RECT 415.800 332.000 416.600 332.200 ;
        RECT 417.400 331.400 418.200 331.600 ;
        RECT 407.600 331.000 413.200 331.200 ;
        RECT 407.400 330.800 413.200 331.000 ;
        RECT 399.600 329.800 402.000 330.400 ;
        RECT 403.400 330.600 413.200 330.800 ;
        RECT 403.400 330.200 408.200 330.600 ;
        RECT 399.600 328.800 400.200 329.800 ;
        RECT 398.800 328.000 400.200 328.800 ;
        RECT 401.800 329.000 402.600 329.200 ;
        RECT 403.400 329.000 404.000 330.200 ;
        RECT 401.800 328.400 404.000 329.000 ;
        RECT 404.600 329.000 410.000 329.600 ;
        RECT 404.600 328.800 405.400 329.000 ;
        RECT 409.200 328.800 410.000 329.000 ;
        RECT 403.000 327.400 403.800 327.600 ;
        RECT 405.800 327.400 406.600 327.600 ;
        RECT 399.600 326.200 400.400 327.000 ;
        RECT 403.000 326.800 406.600 327.400 ;
        RECT 403.800 326.200 404.400 326.800 ;
        RECT 409.200 326.200 410.000 327.000 ;
        RECT 399.000 322.200 400.200 326.200 ;
        RECT 403.600 322.200 404.400 326.200 ;
        RECT 408.000 325.600 410.000 326.200 ;
        RECT 408.000 322.200 408.800 325.600 ;
        RECT 412.400 322.200 413.200 330.600 ;
        RECT 414.000 330.800 418.200 331.400 ;
        RECT 414.000 322.200 414.800 330.800 ;
        RECT 420.600 330.400 421.200 333.600 ;
        RECT 427.800 333.400 428.600 333.600 ;
        RECT 437.200 333.400 438.000 334.200 ;
        RECT 437.200 332.800 437.800 333.400 ;
        RECT 426.800 332.400 427.600 332.600 ;
        RECT 429.400 332.400 430.200 332.600 ;
        RECT 425.200 331.800 430.200 332.400 ;
        RECT 435.200 332.200 437.800 332.800 ;
        RECT 438.600 332.800 439.200 336.200 ;
        RECT 442.800 335.800 443.600 339.800 ;
        RECT 439.800 334.800 440.600 335.600 ;
        RECT 441.200 335.200 443.600 335.800 ;
        RECT 449.200 335.200 450.000 339.800 ;
        RECT 441.200 335.000 442.000 335.200 ;
        RECT 440.000 334.400 440.600 334.800 ;
        RECT 449.200 334.600 451.400 335.200 ;
        RECT 440.000 333.600 440.800 334.400 ;
        RECT 442.000 334.300 443.600 334.400 ;
        RECT 447.600 334.300 448.400 334.400 ;
        RECT 442.000 333.700 448.400 334.300 ;
        RECT 442.000 333.600 443.600 333.700 ;
        RECT 447.600 333.600 448.400 333.700 ;
        RECT 438.600 332.400 439.600 332.800 ;
        RECT 438.600 332.200 440.400 332.400 ;
        RECT 435.200 332.000 436.000 332.200 ;
        RECT 425.200 331.600 426.000 331.800 ;
        RECT 439.000 331.600 440.400 332.200 ;
        RECT 449.200 331.600 450.000 333.200 ;
        RECT 450.800 331.600 451.400 334.600 ;
        RECT 452.400 332.400 453.200 339.800 ;
        RECT 454.000 336.000 454.800 339.800 ;
        RECT 457.200 336.000 458.000 339.800 ;
        RECT 454.000 335.800 458.000 336.000 ;
        RECT 458.800 335.800 459.600 339.800 ;
        RECT 462.000 337.800 462.800 339.800 ;
        RECT 454.200 335.400 457.800 335.800 ;
        RECT 454.800 334.400 455.600 334.800 ;
        RECT 458.800 334.400 459.400 335.800 ;
        RECT 462.000 334.400 462.600 337.800 ;
        RECT 463.600 335.600 464.400 337.200 ;
        RECT 465.800 336.400 466.600 339.800 ;
        RECT 465.800 335.800 467.600 336.400 ;
        RECT 470.000 336.000 470.800 339.800 ;
        RECT 473.200 336.000 474.000 339.800 ;
        RECT 470.000 335.800 474.000 336.000 ;
        RECT 474.800 335.800 475.600 339.800 ;
        RECT 454.000 333.800 455.600 334.400 ;
        RECT 454.000 333.600 454.800 333.800 ;
        RECT 457.000 333.600 459.600 334.400 ;
        RECT 462.000 333.600 462.800 334.400 ;
        RECT 437.400 331.400 438.200 331.600 ;
        RECT 426.800 331.000 432.400 331.200 ;
        RECT 426.600 330.800 432.400 331.000 ;
        RECT 418.800 329.800 421.200 330.400 ;
        RECT 422.600 330.600 432.400 330.800 ;
        RECT 422.600 330.200 427.400 330.600 ;
        RECT 418.800 328.800 419.400 329.800 ;
        RECT 418.000 328.000 419.400 328.800 ;
        RECT 421.000 329.000 421.800 329.200 ;
        RECT 422.600 329.000 423.200 330.200 ;
        RECT 421.000 328.400 423.200 329.000 ;
        RECT 423.800 329.000 429.200 329.600 ;
        RECT 423.800 328.800 424.600 329.000 ;
        RECT 428.400 328.800 429.200 329.000 ;
        RECT 422.200 327.400 423.000 327.600 ;
        RECT 425.000 327.400 425.800 327.600 ;
        RECT 418.800 326.200 419.600 327.000 ;
        RECT 422.200 326.800 425.800 327.400 ;
        RECT 423.000 326.200 423.600 326.800 ;
        RECT 428.400 326.200 429.200 327.000 ;
        RECT 418.200 322.200 419.400 326.200 ;
        RECT 422.800 322.200 423.600 326.200 ;
        RECT 427.200 325.600 429.200 326.200 ;
        RECT 427.200 322.200 428.000 325.600 ;
        RECT 431.600 322.200 432.400 330.600 ;
        RECT 434.800 330.800 438.200 331.400 ;
        RECT 434.800 330.200 435.400 330.800 ;
        RECT 439.000 330.200 439.600 331.600 ;
        RECT 450.800 330.800 452.000 331.600 ;
        RECT 450.800 330.200 451.400 330.800 ;
        RECT 452.600 330.200 453.200 332.400 ;
        RECT 455.600 331.600 456.400 333.200 ;
        RECT 457.000 330.200 457.600 333.600 ;
        RECT 460.400 330.800 461.200 332.400 ;
        RECT 462.000 332.300 462.600 333.600 ;
        RECT 462.000 331.700 465.900 332.300 ;
        RECT 458.800 330.200 459.600 330.400 ;
        RECT 462.000 330.200 462.600 331.700 ;
        RECT 465.300 330.400 465.900 331.700 ;
        RECT 433.200 329.600 435.400 330.200 ;
        RECT 433.200 322.200 434.000 329.600 ;
        RECT 434.600 329.400 435.400 329.600 ;
        RECT 437.600 329.600 439.600 330.200 ;
        RECT 441.200 329.600 443.600 330.200 ;
        RECT 437.600 328.400 439.200 329.600 ;
        RECT 441.200 329.400 442.000 329.600 ;
        RECT 436.400 327.600 439.200 328.400 ;
        RECT 437.600 322.200 439.200 327.600 ;
        RECT 442.800 322.200 443.600 329.600 ;
        RECT 449.200 329.600 451.400 330.200 ;
        RECT 449.200 322.200 450.000 329.600 ;
        RECT 452.400 322.200 453.200 330.200 ;
        RECT 456.600 329.600 457.600 330.200 ;
        RECT 458.200 329.600 459.600 330.200 ;
        RECT 456.600 324.400 457.400 329.600 ;
        RECT 458.200 328.400 458.800 329.600 ;
        RECT 458.000 327.600 458.800 328.400 ;
        RECT 461.000 329.400 462.800 330.200 ;
        RECT 455.600 323.600 457.400 324.400 ;
        RECT 456.600 322.200 457.400 323.600 ;
        RECT 461.000 322.200 461.800 329.400 ;
        RECT 465.200 328.800 466.000 330.400 ;
        RECT 466.800 330.300 467.600 335.800 ;
        RECT 470.200 335.400 473.800 335.800 ;
        RECT 468.400 334.300 469.200 335.200 ;
        RECT 470.800 334.400 471.600 334.800 ;
        RECT 474.800 334.400 475.400 335.800 ;
        RECT 476.400 335.000 477.200 339.800 ;
        RECT 480.800 338.400 481.600 339.800 ;
        RECT 479.600 337.800 481.600 338.400 ;
        RECT 485.200 337.800 486.000 339.800 ;
        RECT 489.400 338.400 490.600 339.800 ;
        RECT 489.200 337.800 490.600 338.400 ;
        RECT 479.600 337.000 480.400 337.800 ;
        RECT 485.200 337.200 485.800 337.800 ;
        RECT 481.200 336.400 482.000 337.200 ;
        RECT 483.000 336.600 485.800 337.200 ;
        RECT 489.200 337.000 490.000 337.800 ;
        RECT 483.000 336.400 483.800 336.600 ;
        RECT 470.000 334.300 471.600 334.400 ;
        RECT 468.400 333.800 471.600 334.300 ;
        RECT 468.400 333.700 470.800 333.800 ;
        RECT 468.400 333.600 469.200 333.700 ;
        RECT 470.000 333.600 470.800 333.700 ;
        RECT 473.000 333.600 475.600 334.400 ;
        RECT 477.200 334.200 478.800 334.400 ;
        RECT 481.400 334.200 482.000 336.400 ;
        RECT 491.000 335.400 491.800 335.600 ;
        RECT 494.000 335.400 494.800 339.800 ;
        RECT 491.000 334.800 494.800 335.400 ;
        RECT 495.600 335.000 496.400 339.800 ;
        RECT 500.000 338.400 500.800 339.800 ;
        RECT 498.800 337.800 500.800 338.400 ;
        RECT 504.400 337.800 505.200 339.800 ;
        RECT 508.600 338.400 509.800 339.800 ;
        RECT 508.400 337.800 509.800 338.400 ;
        RECT 498.800 337.000 499.600 337.800 ;
        RECT 504.400 337.200 505.000 337.800 ;
        RECT 500.400 336.400 501.200 337.200 ;
        RECT 502.200 336.600 505.000 337.200 ;
        RECT 508.400 337.000 509.200 337.800 ;
        RECT 502.200 336.400 503.000 336.600 ;
        RECT 487.000 334.200 487.800 334.400 ;
        RECT 477.200 333.600 488.200 334.200 ;
        RECT 468.400 332.300 469.200 332.400 ;
        RECT 471.600 332.300 472.400 333.200 ;
        RECT 468.400 331.700 472.400 332.300 ;
        RECT 468.400 331.600 469.200 331.700 ;
        RECT 471.600 331.600 472.400 331.700 ;
        RECT 468.400 330.300 469.200 330.400 ;
        RECT 466.800 329.700 469.200 330.300 ;
        RECT 473.000 330.200 473.600 333.600 ;
        RECT 480.200 333.400 481.000 333.600 ;
        RECT 478.600 332.400 479.400 332.600 ;
        RECT 487.600 332.400 488.200 333.600 ;
        RECT 489.200 332.800 490.000 333.000 ;
        RECT 478.600 332.300 483.600 332.400 ;
        RECT 486.000 332.300 486.800 332.400 ;
        RECT 478.600 331.800 486.800 332.300 ;
        RECT 482.800 331.700 486.800 331.800 ;
        RECT 482.800 331.600 483.600 331.700 ;
        RECT 486.000 331.600 486.800 331.700 ;
        RECT 487.600 331.600 488.400 332.400 ;
        RECT 489.200 332.200 493.000 332.800 ;
        RECT 492.200 332.000 493.000 332.200 ;
        RECT 476.400 331.000 482.000 331.200 ;
        RECT 476.400 330.800 482.200 331.000 ;
        RECT 476.400 330.600 486.200 330.800 ;
        RECT 474.800 330.200 475.600 330.400 ;
        RECT 466.800 322.200 467.600 329.700 ;
        RECT 468.400 329.600 469.200 329.700 ;
        RECT 472.600 329.600 473.600 330.200 ;
        RECT 474.200 329.600 475.600 330.200 ;
        RECT 472.600 322.200 473.400 329.600 ;
        RECT 474.200 328.400 474.800 329.600 ;
        RECT 474.000 327.600 474.800 328.400 ;
        RECT 476.400 322.200 477.200 330.600 ;
        RECT 481.400 330.200 486.200 330.600 ;
        RECT 479.600 329.000 485.000 329.600 ;
        RECT 479.600 328.800 480.400 329.000 ;
        RECT 484.200 328.800 485.000 329.000 ;
        RECT 485.600 329.000 486.200 330.200 ;
        RECT 487.600 330.400 488.200 331.600 ;
        RECT 490.600 331.400 491.400 331.600 ;
        RECT 494.000 331.400 494.800 334.800 ;
        RECT 496.400 334.200 498.000 334.400 ;
        RECT 500.600 334.200 501.200 336.400 ;
        RECT 510.200 335.400 511.000 335.600 ;
        RECT 513.200 335.400 514.000 339.800 ;
        RECT 510.200 334.800 514.000 335.400 ;
        RECT 506.200 334.200 507.000 334.400 ;
        RECT 496.400 333.600 507.400 334.200 ;
        RECT 499.400 333.400 500.200 333.600 ;
        RECT 497.800 332.400 498.600 332.600 ;
        RECT 500.400 332.400 501.200 332.600 ;
        RECT 506.800 332.400 507.400 333.600 ;
        RECT 508.400 332.800 509.200 333.000 ;
        RECT 497.800 331.800 502.800 332.400 ;
        RECT 502.000 331.600 502.800 331.800 ;
        RECT 506.800 331.600 507.600 332.400 ;
        RECT 508.400 332.200 512.200 332.800 ;
        RECT 511.400 332.000 512.200 332.200 ;
        RECT 490.600 330.800 494.800 331.400 ;
        RECT 487.600 329.800 490.000 330.400 ;
        RECT 487.000 329.000 487.800 329.200 ;
        RECT 485.600 328.400 487.800 329.000 ;
        RECT 489.400 328.800 490.000 329.800 ;
        RECT 489.400 328.000 490.800 328.800 ;
        RECT 483.000 327.400 483.800 327.600 ;
        RECT 485.800 327.400 486.600 327.600 ;
        RECT 479.600 326.200 480.400 327.000 ;
        RECT 483.000 326.800 486.600 327.400 ;
        RECT 485.200 326.200 485.800 326.800 ;
        RECT 489.200 326.200 490.000 327.000 ;
        RECT 479.600 325.600 481.600 326.200 ;
        RECT 480.800 322.200 481.600 325.600 ;
        RECT 485.200 322.200 486.000 326.200 ;
        RECT 489.400 322.200 490.600 326.200 ;
        RECT 494.000 322.200 494.800 330.800 ;
        RECT 495.600 331.000 501.200 331.200 ;
        RECT 495.600 330.800 501.400 331.000 ;
        RECT 495.600 330.600 505.400 330.800 ;
        RECT 495.600 322.200 496.400 330.600 ;
        RECT 500.600 330.200 505.400 330.600 ;
        RECT 498.800 329.000 504.200 329.600 ;
        RECT 498.800 328.800 499.600 329.000 ;
        RECT 503.400 328.800 504.200 329.000 ;
        RECT 504.800 329.000 505.400 330.200 ;
        RECT 506.800 330.400 507.400 331.600 ;
        RECT 509.800 331.400 510.600 331.600 ;
        RECT 513.200 331.400 514.000 334.800 ;
        RECT 514.800 335.200 515.600 339.800 ;
        RECT 514.800 334.600 517.000 335.200 ;
        RECT 509.800 330.800 514.000 331.400 ;
        RECT 506.800 329.800 509.200 330.400 ;
        RECT 506.200 329.000 507.000 329.200 ;
        RECT 504.800 328.400 507.000 329.000 ;
        RECT 508.600 328.800 509.200 329.800 ;
        RECT 508.600 328.000 510.000 328.800 ;
        RECT 502.200 327.400 503.000 327.600 ;
        RECT 505.000 327.400 505.800 327.600 ;
        RECT 498.800 326.200 499.600 327.000 ;
        RECT 502.200 326.800 505.800 327.400 ;
        RECT 504.400 326.200 505.000 326.800 ;
        RECT 508.400 326.200 509.200 327.000 ;
        RECT 498.800 325.600 500.800 326.200 ;
        RECT 500.000 322.200 500.800 325.600 ;
        RECT 504.400 322.200 505.200 326.200 ;
        RECT 508.600 322.200 509.800 326.200 ;
        RECT 513.200 322.200 514.000 330.800 ;
        RECT 516.400 331.600 517.000 334.600 ;
        RECT 518.000 332.400 518.800 339.800 ;
        RECT 521.200 336.000 522.000 339.800 ;
        RECT 516.400 330.800 517.600 331.600 ;
        RECT 516.400 330.200 517.000 330.800 ;
        RECT 518.200 330.200 518.800 332.400 ;
        RECT 514.800 329.600 517.000 330.200 ;
        RECT 514.800 322.200 515.600 329.600 ;
        RECT 518.000 322.200 518.800 330.200 ;
        RECT 521.000 335.200 522.000 336.000 ;
        RECT 521.000 330.800 521.800 335.200 ;
        RECT 522.800 334.600 523.600 339.800 ;
        RECT 529.200 336.600 530.000 339.800 ;
        RECT 530.800 337.000 531.600 339.800 ;
        RECT 532.400 337.000 533.200 339.800 ;
        RECT 534.000 337.000 534.800 339.800 ;
        RECT 535.600 337.000 536.400 339.800 ;
        RECT 538.800 337.000 539.600 339.800 ;
        RECT 542.000 337.000 542.800 339.800 ;
        RECT 543.600 337.000 544.400 339.800 ;
        RECT 545.200 337.000 546.000 339.800 ;
        RECT 527.600 335.800 530.000 336.600 ;
        RECT 546.800 336.600 547.600 339.800 ;
        RECT 527.600 335.200 528.400 335.800 ;
        RECT 522.400 334.000 523.600 334.600 ;
        RECT 526.600 334.600 528.400 335.200 ;
        RECT 532.400 335.600 533.400 336.400 ;
        RECT 536.400 335.600 538.000 336.400 ;
        RECT 538.800 335.800 543.400 336.400 ;
        RECT 546.800 335.800 549.400 336.600 ;
        RECT 538.800 335.600 539.600 335.800 ;
        RECT 522.400 332.000 523.000 334.000 ;
        RECT 526.600 333.400 527.400 334.600 ;
        RECT 523.600 332.600 527.400 333.400 ;
        RECT 532.400 332.800 533.200 335.600 ;
        RECT 538.800 334.800 539.600 335.000 ;
        RECT 535.200 334.200 539.600 334.800 ;
        RECT 535.200 334.000 536.000 334.200 ;
        RECT 540.400 333.600 541.200 335.200 ;
        RECT 542.600 333.400 543.400 335.800 ;
        RECT 548.600 335.200 549.400 335.800 ;
        RECT 548.600 334.400 551.600 335.200 ;
        RECT 553.200 333.800 554.000 339.800 ;
        RECT 535.600 332.600 538.800 333.400 ;
        RECT 542.600 332.600 544.600 333.400 ;
        RECT 545.200 333.000 554.000 333.800 ;
        RECT 529.200 332.000 530.000 332.600 ;
        RECT 546.800 332.000 547.600 332.400 ;
        RECT 551.800 332.000 552.600 332.200 ;
        RECT 522.400 331.400 523.200 332.000 ;
        RECT 529.200 331.400 552.600 332.000 ;
        RECT 521.000 330.000 522.000 330.800 ;
        RECT 521.200 322.200 522.000 330.000 ;
        RECT 522.600 329.600 523.200 331.400 ;
        RECT 522.600 329.000 531.600 329.600 ;
        RECT 522.600 327.400 523.200 329.000 ;
        RECT 530.800 328.800 531.600 329.000 ;
        RECT 534.000 329.000 542.600 329.600 ;
        RECT 534.000 328.800 534.800 329.000 ;
        RECT 525.800 327.600 528.400 328.400 ;
        RECT 522.600 326.800 525.200 327.400 ;
        RECT 524.400 322.200 525.200 326.800 ;
        RECT 527.600 322.200 528.400 327.600 ;
        RECT 529.000 326.800 533.200 327.600 ;
        RECT 530.800 322.200 531.600 325.000 ;
        RECT 532.400 322.200 533.200 325.000 ;
        RECT 534.000 322.200 534.800 325.000 ;
        RECT 535.600 322.200 536.400 328.400 ;
        RECT 538.800 327.600 541.400 328.400 ;
        RECT 542.000 328.200 542.600 329.000 ;
        RECT 543.600 329.400 544.400 329.600 ;
        RECT 543.600 329.000 549.000 329.400 ;
        RECT 543.600 328.800 549.800 329.000 ;
        RECT 548.400 328.200 549.800 328.800 ;
        RECT 542.000 327.600 547.800 328.200 ;
        RECT 550.800 328.000 552.400 328.800 ;
        RECT 550.800 327.600 551.400 328.000 ;
        RECT 538.800 322.200 539.600 327.000 ;
        RECT 542.000 322.200 542.800 327.000 ;
        RECT 547.200 326.800 551.400 327.600 ;
        RECT 553.200 327.400 554.000 333.000 ;
        RECT 552.000 326.800 554.000 327.400 ;
        RECT 554.800 335.400 555.600 339.800 ;
        RECT 559.000 338.400 560.200 339.800 ;
        RECT 559.000 337.800 560.400 338.400 ;
        RECT 563.600 337.800 564.400 339.800 ;
        RECT 568.000 338.400 568.800 339.800 ;
        RECT 568.000 337.800 570.000 338.400 ;
        RECT 559.600 337.000 560.400 337.800 ;
        RECT 563.800 337.200 564.400 337.800 ;
        RECT 563.800 336.600 566.600 337.200 ;
        RECT 565.800 336.400 566.600 336.600 ;
        RECT 567.600 336.400 568.400 337.200 ;
        RECT 569.200 337.000 570.000 337.800 ;
        RECT 557.800 335.400 558.600 335.600 ;
        RECT 554.800 334.800 558.600 335.400 ;
        RECT 554.800 331.400 555.600 334.800 ;
        RECT 561.800 334.200 562.600 334.400 ;
        RECT 567.600 334.200 568.200 336.400 ;
        RECT 572.400 335.000 573.200 339.800 ;
        RECT 574.000 335.200 574.800 339.800 ;
        RECT 578.800 335.200 579.600 339.800 ;
        RECT 574.000 334.600 576.200 335.200 ;
        RECT 578.800 334.600 581.000 335.200 ;
        RECT 570.800 334.200 572.400 334.400 ;
        RECT 561.400 333.600 572.400 334.200 ;
        RECT 559.600 332.800 560.400 333.000 ;
        RECT 556.600 332.200 560.400 332.800 ;
        RECT 561.400 332.400 562.000 333.600 ;
        RECT 568.600 333.400 569.400 333.600 ;
        RECT 570.200 332.400 571.000 332.600 ;
        RECT 556.600 332.000 557.400 332.200 ;
        RECT 561.200 331.600 562.000 332.400 ;
        RECT 566.000 331.800 571.000 332.400 ;
        RECT 566.000 331.600 566.800 331.800 ;
        RECT 574.000 331.600 574.800 333.200 ;
        RECT 575.600 331.600 576.200 334.600 ;
        RECT 578.800 331.600 579.600 333.200 ;
        RECT 580.400 331.600 581.000 334.600 ;
        RECT 558.200 331.400 559.000 331.600 ;
        RECT 554.800 330.800 559.000 331.400 ;
        RECT 543.600 322.200 544.400 325.000 ;
        RECT 545.200 322.200 546.000 325.000 ;
        RECT 548.400 322.200 549.200 326.800 ;
        RECT 552.000 326.200 552.600 326.800 ;
        RECT 551.600 325.600 552.600 326.200 ;
        RECT 551.600 322.200 552.400 325.600 ;
        RECT 554.800 322.200 555.600 330.800 ;
        RECT 561.400 330.400 562.000 331.600 ;
        RECT 567.600 331.000 573.200 331.200 ;
        RECT 567.400 330.800 573.200 331.000 ;
        RECT 559.600 329.800 562.000 330.400 ;
        RECT 563.400 330.600 573.200 330.800 ;
        RECT 563.400 330.200 568.200 330.600 ;
        RECT 559.600 328.800 560.200 329.800 ;
        RECT 558.800 328.000 560.200 328.800 ;
        RECT 561.800 329.000 562.600 329.200 ;
        RECT 563.400 329.000 564.000 330.200 ;
        RECT 561.800 328.400 564.000 329.000 ;
        RECT 564.600 329.000 570.000 329.600 ;
        RECT 564.600 328.800 565.400 329.000 ;
        RECT 569.200 328.800 570.000 329.000 ;
        RECT 563.000 327.400 563.800 327.600 ;
        RECT 565.800 327.400 566.600 327.600 ;
        RECT 559.600 326.200 560.400 327.000 ;
        RECT 563.000 326.800 566.600 327.400 ;
        RECT 563.800 326.200 564.400 326.800 ;
        RECT 569.200 326.200 570.000 327.000 ;
        RECT 559.000 322.200 560.200 326.200 ;
        RECT 563.600 322.200 564.400 326.200 ;
        RECT 568.000 325.600 570.000 326.200 ;
        RECT 568.000 322.200 568.800 325.600 ;
        RECT 572.400 322.200 573.200 330.600 ;
        RECT 575.600 330.800 576.800 331.600 ;
        RECT 580.400 330.800 581.600 331.600 ;
        RECT 575.600 330.200 576.200 330.800 ;
        RECT 580.400 330.200 581.000 330.800 ;
        RECT 574.000 329.600 576.200 330.200 ;
        RECT 578.800 329.600 581.000 330.200 ;
        RECT 574.000 322.200 574.800 329.600 ;
        RECT 578.800 322.200 579.600 329.600 ;
        RECT 2.000 313.600 2.800 314.400 ;
        RECT 2.000 312.400 2.600 313.600 ;
        RECT 3.400 312.400 4.200 319.800 ;
        RECT 10.200 312.600 11.000 319.800 ;
        RECT 15.000 312.600 15.800 319.800 ;
        RECT 1.200 311.800 2.600 312.400 ;
        RECT 3.200 311.800 4.200 312.400 ;
        RECT 9.200 311.800 11.000 312.600 ;
        RECT 14.000 311.800 15.800 312.600 ;
        RECT 1.200 311.600 2.000 311.800 ;
        RECT 3.200 308.400 3.800 311.800 ;
        RECT 4.400 308.800 5.200 310.400 ;
        RECT 9.400 308.400 10.000 311.800 ;
        RECT 10.800 309.600 11.600 311.200 ;
        RECT 14.200 308.400 14.800 311.800 ;
        RECT 15.600 309.600 16.400 311.200 ;
        RECT 18.800 310.300 19.600 319.800 ;
        RECT 21.000 312.600 21.800 319.800 ;
        RECT 26.000 313.600 26.800 314.400 ;
        RECT 21.000 311.800 22.800 312.600 ;
        RECT 26.000 312.400 26.600 313.600 ;
        RECT 27.400 312.400 28.200 319.800 ;
        RECT 25.200 311.800 26.600 312.400 ;
        RECT 27.200 311.800 28.200 312.400 ;
        RECT 20.400 310.300 21.200 311.200 ;
        RECT 18.800 309.700 21.200 310.300 ;
        RECT 1.200 307.600 3.800 308.400 ;
        RECT 6.000 308.300 6.800 308.400 ;
        RECT 7.600 308.300 8.400 308.400 ;
        RECT 6.000 308.200 8.400 308.300 ;
        RECT 5.200 307.700 8.400 308.200 ;
        RECT 5.200 307.600 6.800 307.700 ;
        RECT 7.600 307.600 8.400 307.700 ;
        RECT 9.200 307.600 10.000 308.400 ;
        RECT 14.000 307.600 14.800 308.400 ;
        RECT 1.400 306.200 2.000 307.600 ;
        RECT 5.200 307.200 6.000 307.600 ;
        RECT 3.000 306.200 6.600 306.600 ;
        RECT 7.700 306.400 8.300 307.600 ;
        RECT 1.200 302.200 2.000 306.200 ;
        RECT 2.800 306.000 6.800 306.200 ;
        RECT 2.800 302.200 3.600 306.000 ;
        RECT 6.000 302.200 6.800 306.000 ;
        RECT 7.600 304.800 8.400 306.400 ;
        RECT 9.400 306.300 10.000 307.600 ;
        RECT 12.400 306.300 13.200 306.400 ;
        RECT 9.300 305.700 13.200 306.300 ;
        RECT 9.400 304.200 10.000 305.700 ;
        RECT 12.400 304.800 13.200 305.700 ;
        RECT 14.200 304.400 14.800 307.600 ;
        RECT 17.200 306.800 18.000 308.400 ;
        RECT 9.200 302.200 10.000 304.200 ;
        RECT 14.000 302.200 14.800 304.400 ;
        RECT 18.800 302.200 19.600 309.700 ;
        RECT 20.400 309.600 21.200 309.700 ;
        RECT 22.000 308.400 22.600 311.800 ;
        RECT 25.200 311.600 26.000 311.800 ;
        RECT 27.200 308.400 27.800 311.800 ;
        RECT 31.600 311.600 32.400 313.200 ;
        RECT 28.400 308.800 29.200 310.400 ;
        RECT 22.000 307.600 22.800 308.400 ;
        RECT 25.200 307.600 27.800 308.400 ;
        RECT 30.000 308.200 30.800 308.400 ;
        RECT 29.200 307.600 30.800 308.200 ;
        RECT 20.400 306.300 21.200 306.400 ;
        RECT 22.000 306.300 22.600 307.600 ;
        RECT 20.400 305.700 22.700 306.300 ;
        RECT 20.400 305.600 21.200 305.700 ;
        RECT 22.000 304.200 22.600 305.700 ;
        RECT 23.600 304.800 24.400 306.400 ;
        RECT 25.400 306.200 26.000 307.600 ;
        RECT 29.200 307.200 30.000 307.600 ;
        RECT 27.000 306.200 30.600 306.600 ;
        RECT 33.200 306.200 34.000 319.800 ;
        RECT 37.000 312.600 37.800 319.800 ;
        RECT 37.000 311.800 38.800 312.600 ;
        RECT 36.400 309.600 37.200 311.200 ;
        RECT 38.000 308.400 38.600 311.800 ;
        RECT 42.800 310.300 43.600 319.800 ;
        RECT 46.800 313.600 47.600 314.400 ;
        RECT 44.400 311.600 45.200 313.200 ;
        RECT 46.800 312.400 47.400 313.600 ;
        RECT 48.200 312.400 49.000 319.800 ;
        RECT 52.400 312.400 53.200 319.800 ;
        RECT 53.800 312.400 54.600 312.600 ;
        RECT 46.000 311.800 47.400 312.400 ;
        RECT 46.000 311.600 46.800 311.800 ;
        RECT 48.000 311.600 50.000 312.400 ;
        RECT 52.400 311.800 54.600 312.400 ;
        RECT 56.800 312.400 58.400 319.800 ;
        RECT 60.400 312.400 61.200 312.600 ;
        RECT 62.000 312.400 62.800 319.800 ;
        RECT 56.800 311.800 58.800 312.400 ;
        RECT 60.400 311.800 62.800 312.400 ;
        RECT 46.100 310.300 46.700 311.600 ;
        RECT 42.800 309.700 46.700 310.300 ;
        RECT 34.800 306.800 35.600 308.400 ;
        RECT 38.000 307.600 38.800 308.400 ;
        RECT 22.000 302.200 22.800 304.200 ;
        RECT 25.200 302.200 26.000 306.200 ;
        RECT 26.800 306.000 30.800 306.200 ;
        RECT 26.800 302.200 27.600 306.000 ;
        RECT 30.000 302.200 30.800 306.000 ;
        RECT 32.200 305.600 34.000 306.200 ;
        RECT 32.200 304.400 33.000 305.600 ;
        RECT 38.000 304.400 38.600 307.600 ;
        RECT 41.200 306.800 42.000 308.400 ;
        RECT 39.600 304.800 40.400 306.400 ;
        RECT 42.800 306.200 43.600 309.700 ;
        RECT 48.000 308.400 48.600 311.600 ;
        RECT 54.000 311.200 54.600 311.800 ;
        RECT 54.000 310.600 57.400 311.200 ;
        RECT 56.600 310.400 57.400 310.600 ;
        RECT 58.200 310.400 58.800 311.800 ;
        RECT 63.600 311.600 64.400 313.200 ;
        RECT 49.200 308.800 50.000 310.400 ;
        RECT 50.800 310.300 51.600 310.400 ;
        RECT 50.800 309.700 53.100 310.300 ;
        RECT 50.800 309.600 51.600 309.700 ;
        RECT 52.500 308.400 53.100 309.700 ;
        RECT 54.400 309.800 55.200 310.000 ;
        RECT 58.200 309.800 59.600 310.400 ;
        RECT 54.400 309.200 57.000 309.800 ;
        RECT 56.400 308.600 57.000 309.200 ;
        RECT 57.800 309.600 59.600 309.800 ;
        RECT 57.800 309.200 58.800 309.600 ;
        RECT 46.000 307.600 48.600 308.400 ;
        RECT 50.800 308.200 51.600 308.400 ;
        RECT 50.000 307.600 51.600 308.200 ;
        RECT 52.400 308.200 54.000 308.400 ;
        RECT 52.400 307.600 55.800 308.200 ;
        RECT 56.400 307.800 57.200 308.600 ;
        RECT 46.200 306.200 46.800 307.600 ;
        RECT 50.000 307.200 50.800 307.600 ;
        RECT 55.200 307.200 55.800 307.600 ;
        RECT 53.800 306.800 54.600 307.000 ;
        RECT 47.800 306.200 51.400 306.600 ;
        RECT 52.400 306.200 54.600 306.800 ;
        RECT 55.200 306.600 57.200 307.200 ;
        RECT 55.600 306.400 57.200 306.600 ;
        RECT 42.800 305.600 44.600 306.200 ;
        RECT 32.200 303.600 34.000 304.400 ;
        RECT 32.200 302.200 33.000 303.600 ;
        RECT 38.000 302.200 38.800 304.400 ;
        RECT 43.800 302.200 44.600 305.600 ;
        RECT 46.000 302.200 46.800 306.200 ;
        RECT 47.600 306.000 51.600 306.200 ;
        RECT 47.600 302.200 48.400 306.000 ;
        RECT 50.800 302.200 51.600 306.000 ;
        RECT 52.400 302.200 53.200 306.200 ;
        RECT 57.800 305.800 58.400 309.200 ;
        RECT 59.200 307.600 60.000 308.400 ;
        RECT 61.200 307.600 62.800 308.400 ;
        RECT 59.200 307.200 59.800 307.600 ;
        RECT 59.000 306.400 59.800 307.200 ;
        RECT 60.400 306.800 61.200 307.000 ;
        RECT 60.400 306.200 62.800 306.800 ;
        RECT 65.200 306.200 66.000 319.800 ;
        RECT 66.800 308.300 67.600 308.400 ;
        RECT 68.400 308.300 69.200 308.400 ;
        RECT 66.800 307.700 69.200 308.300 ;
        RECT 66.800 306.800 67.600 307.700 ;
        RECT 68.400 307.600 69.200 307.700 ;
        RECT 56.800 304.400 58.400 305.800 ;
        RECT 55.600 303.600 58.400 304.400 ;
        RECT 56.800 302.200 58.400 303.600 ;
        RECT 62.000 302.200 62.800 306.200 ;
        RECT 64.200 305.600 66.000 306.200 ;
        RECT 64.200 304.400 65.000 305.600 ;
        RECT 68.400 304.800 69.200 306.400 ;
        RECT 64.200 303.600 66.000 304.400 ;
        RECT 64.200 302.200 65.000 303.600 ;
        RECT 70.000 302.200 70.800 319.800 ;
        RECT 71.600 312.400 72.400 319.800 ;
        RECT 74.800 312.800 75.600 319.800 ;
        RECT 78.000 319.200 82.000 319.800 ;
        RECT 71.600 311.800 74.200 312.400 ;
        RECT 74.800 311.800 75.800 312.800 ;
        RECT 78.000 311.800 78.800 319.200 ;
        RECT 79.600 311.800 80.400 318.600 ;
        RECT 81.200 312.400 82.000 319.200 ;
        RECT 84.400 312.400 85.200 319.800 ;
        RECT 81.200 311.800 85.200 312.400 ;
        RECT 71.600 309.600 72.600 310.400 ;
        RECT 71.800 308.800 72.600 309.600 ;
        RECT 73.600 309.800 74.200 311.800 ;
        RECT 73.600 309.000 74.600 309.800 ;
        RECT 73.600 307.400 74.200 309.000 ;
        RECT 75.200 308.400 75.800 311.800 ;
        RECT 79.800 311.200 80.400 311.800 ;
        RECT 76.400 310.300 77.200 310.400 ;
        RECT 78.000 310.300 78.800 311.200 ;
        RECT 79.800 310.600 81.800 311.200 ;
        RECT 76.400 309.700 78.800 310.300 ;
        RECT 76.400 309.600 77.200 309.700 ;
        RECT 78.000 309.600 78.800 309.700 ;
        RECT 81.200 310.400 81.800 310.600 ;
        RECT 83.600 310.400 84.400 310.800 ;
        RECT 81.200 309.600 82.000 310.400 ;
        RECT 83.600 309.800 85.200 310.400 ;
        RECT 84.400 309.600 85.200 309.800 ;
        RECT 79.800 308.800 80.600 309.600 ;
        RECT 79.800 308.400 80.400 308.800 ;
        RECT 74.800 307.600 75.800 308.400 ;
        RECT 79.600 307.600 80.400 308.400 ;
        RECT 71.600 306.800 74.200 307.400 ;
        RECT 71.600 302.200 72.400 306.800 ;
        RECT 75.200 306.200 75.800 307.600 ;
        RECT 81.200 306.200 81.800 309.600 ;
        RECT 82.800 307.600 83.600 309.200 ;
        RECT 86.000 306.800 86.800 308.400 ;
        RECT 87.600 306.200 88.400 319.800 ;
        RECT 89.200 312.300 90.000 313.200 ;
        RECT 90.800 312.300 91.600 319.800 ;
        RECT 89.200 311.700 91.600 312.300 ;
        RECT 96.600 312.400 97.400 319.800 ;
        RECT 98.000 313.600 98.800 314.400 ;
        RECT 98.200 312.400 98.800 313.600 ;
        RECT 103.000 312.600 103.800 319.800 ;
        RECT 96.600 311.800 97.600 312.400 ;
        RECT 98.200 311.800 99.600 312.400 ;
        RECT 102.000 311.800 103.800 312.600 ;
        RECT 107.800 312.400 108.600 319.800 ;
        RECT 109.200 313.600 110.000 314.400 ;
        RECT 109.400 312.400 110.000 313.600 ;
        RECT 111.600 312.400 112.400 319.800 ;
        RECT 114.800 312.400 115.600 319.800 ;
        RECT 107.800 311.800 108.800 312.400 ;
        RECT 109.400 311.800 110.800 312.400 ;
        RECT 111.600 311.800 115.600 312.400 ;
        RECT 116.400 311.800 117.200 319.800 ;
        RECT 120.600 314.400 121.400 319.800 ;
        RECT 119.600 313.600 121.400 314.400 ;
        RECT 122.000 313.600 122.800 314.400 ;
        RECT 120.600 312.400 121.400 313.600 ;
        RECT 122.200 312.400 122.800 313.600 ;
        RECT 120.600 311.800 121.600 312.400 ;
        RECT 122.200 311.800 123.600 312.400 ;
        RECT 89.200 311.600 90.000 311.700 ;
        RECT 74.800 305.600 75.800 306.200 ;
        RECT 74.800 302.200 75.600 305.600 ;
        RECT 80.600 302.200 82.200 306.200 ;
        RECT 87.600 305.600 89.400 306.200 ;
        RECT 88.600 302.200 89.400 305.600 ;
        RECT 90.800 302.200 91.600 311.700 ;
        RECT 95.600 308.800 96.400 310.400 ;
        RECT 97.000 308.400 97.600 311.800 ;
        RECT 98.800 311.600 99.600 311.800 ;
        RECT 102.200 308.400 102.800 311.800 ;
        RECT 103.600 310.300 104.400 311.200 ;
        RECT 106.800 310.300 107.600 310.400 ;
        RECT 103.600 309.700 107.600 310.300 ;
        RECT 103.600 309.600 104.400 309.700 ;
        RECT 106.800 308.800 107.600 309.700 ;
        RECT 108.200 308.400 108.800 311.800 ;
        RECT 110.000 311.600 110.800 311.800 ;
        RECT 112.400 310.400 113.200 310.800 ;
        RECT 116.400 310.400 117.000 311.800 ;
        RECT 111.600 309.800 113.200 310.400 ;
        RECT 114.800 310.300 117.200 310.400 ;
        RECT 119.600 310.300 120.400 310.400 ;
        RECT 114.800 309.800 120.400 310.300 ;
        RECT 111.600 309.600 112.400 309.800 ;
        RECT 92.400 308.300 93.200 308.400 ;
        RECT 94.000 308.300 94.800 308.400 ;
        RECT 92.400 308.200 94.800 308.300 ;
        RECT 92.400 307.700 95.600 308.200 ;
        RECT 92.400 307.600 93.200 307.700 ;
        RECT 94.000 307.600 95.600 307.700 ;
        RECT 97.000 307.600 99.600 308.400 ;
        RECT 102.000 307.600 102.800 308.400 ;
        RECT 105.200 308.200 106.000 308.400 ;
        RECT 105.200 307.600 106.800 308.200 ;
        RECT 108.200 307.600 110.800 308.400 ;
        RECT 113.200 307.600 114.000 309.200 ;
        RECT 94.800 307.200 95.600 307.600 ;
        RECT 92.400 304.800 93.200 306.400 ;
        RECT 94.200 306.200 97.800 306.600 ;
        RECT 98.800 306.200 99.400 307.600 ;
        RECT 94.000 306.000 98.000 306.200 ;
        RECT 94.000 302.200 94.800 306.000 ;
        RECT 97.200 302.200 98.000 306.000 ;
        RECT 98.800 302.200 99.600 306.200 ;
        RECT 100.400 304.800 101.200 306.400 ;
        RECT 102.200 304.400 102.800 307.600 ;
        RECT 106.000 307.200 106.800 307.600 ;
        RECT 105.400 306.200 109.000 306.600 ;
        RECT 110.000 306.200 110.600 307.600 ;
        RECT 114.800 306.200 115.400 309.800 ;
        RECT 116.400 309.700 120.400 309.800 ;
        RECT 116.400 309.600 117.200 309.700 ;
        RECT 119.600 308.800 120.400 309.700 ;
        RECT 121.000 308.400 121.600 311.800 ;
        RECT 122.800 311.600 123.600 311.800 ;
        RECT 118.000 308.200 118.800 308.400 ;
        RECT 118.000 307.600 119.600 308.200 ;
        RECT 121.000 307.600 123.600 308.400 ;
        RECT 118.800 307.200 119.600 307.600 ;
        RECT 102.000 302.200 102.800 304.400 ;
        RECT 105.200 306.000 109.200 306.200 ;
        RECT 105.200 302.200 106.000 306.000 ;
        RECT 108.400 302.200 109.200 306.000 ;
        RECT 110.000 302.200 110.800 306.200 ;
        RECT 114.800 302.200 115.600 306.200 ;
        RECT 116.400 305.600 117.200 306.400 ;
        RECT 118.200 306.200 121.800 306.600 ;
        RECT 122.800 306.200 123.400 307.600 ;
        RECT 118.000 306.000 122.000 306.200 ;
        RECT 116.200 304.800 117.000 305.600 ;
        RECT 118.000 302.200 118.800 306.000 ;
        RECT 121.200 302.200 122.000 306.000 ;
        RECT 122.800 302.200 123.600 306.200 ;
        RECT 124.400 304.800 125.200 306.400 ;
        RECT 126.000 302.200 126.800 319.800 ;
        RECT 127.600 311.600 128.400 313.200 ;
        RECT 129.200 306.200 130.000 319.800 ;
        RECT 130.800 306.800 131.600 308.400 ;
        RECT 128.200 305.600 130.000 306.200 ;
        RECT 128.200 304.400 129.000 305.600 ;
        RECT 128.200 303.600 130.000 304.400 ;
        RECT 128.200 302.200 129.000 303.600 ;
        RECT 132.400 302.200 133.200 319.800 ;
        RECT 141.200 313.600 142.000 314.400 ;
        RECT 141.200 312.400 141.800 313.600 ;
        RECT 142.600 312.400 143.400 319.800 ;
        RECT 137.200 312.300 138.000 312.400 ;
        RECT 140.400 312.300 141.800 312.400 ;
        RECT 137.200 311.800 141.800 312.300 ;
        RECT 142.400 311.800 143.400 312.400 ;
        RECT 137.200 311.700 141.200 311.800 ;
        RECT 137.200 311.600 138.000 311.700 ;
        RECT 140.400 311.600 141.200 311.700 ;
        RECT 142.400 308.400 143.000 311.800 ;
        RECT 143.600 308.800 144.400 310.400 ;
        RECT 148.400 310.300 149.200 319.800 ;
        RECT 152.400 313.600 153.200 314.400 ;
        RECT 150.000 311.600 150.800 313.200 ;
        RECT 152.400 312.400 153.000 313.600 ;
        RECT 153.800 312.400 154.600 319.800 ;
        RECT 151.600 311.800 153.000 312.400 ;
        RECT 153.600 311.800 154.600 312.400 ;
        RECT 158.600 312.600 159.400 319.800 ;
        RECT 158.600 311.800 160.400 312.600 ;
        RECT 163.400 312.400 164.200 319.800 ;
        RECT 162.800 311.800 164.200 312.400 ;
        RECT 151.600 311.600 152.400 311.800 ;
        RECT 151.700 310.300 152.300 311.600 ;
        RECT 148.400 309.700 152.300 310.300 ;
        RECT 140.400 307.600 143.000 308.400 ;
        RECT 145.200 308.200 146.000 308.400 ;
        RECT 144.400 307.600 146.000 308.200 ;
        RECT 134.000 304.800 134.800 306.400 ;
        RECT 140.600 306.200 141.200 307.600 ;
        RECT 144.400 307.200 145.200 307.600 ;
        RECT 146.800 306.800 147.600 308.400 ;
        RECT 142.200 306.200 145.800 306.600 ;
        RECT 148.400 306.200 149.200 309.700 ;
        RECT 153.600 308.400 154.200 311.800 ;
        RECT 154.800 310.300 155.600 310.400 ;
        RECT 156.400 310.300 157.200 310.400 ;
        RECT 154.800 309.700 157.200 310.300 ;
        RECT 154.800 308.800 155.600 309.700 ;
        RECT 156.400 309.600 157.200 309.700 ;
        RECT 158.000 309.600 158.800 311.200 ;
        RECT 159.600 308.400 160.200 311.800 ;
        RECT 162.800 310.400 163.400 311.800 ;
        RECT 167.600 311.200 168.400 319.800 ;
        RECT 169.800 312.600 170.600 319.800 ;
        RECT 175.600 315.800 176.400 319.800 ;
        RECT 169.800 311.800 171.600 312.600 ;
        RECT 164.400 310.800 168.400 311.200 ;
        RECT 164.200 310.600 168.400 310.800 ;
        RECT 162.800 309.600 163.600 310.400 ;
        RECT 164.200 310.000 165.000 310.600 ;
        RECT 151.600 307.600 154.200 308.400 ;
        RECT 156.400 308.300 157.200 308.400 ;
        RECT 158.000 308.300 158.800 308.400 ;
        RECT 156.400 308.200 158.800 308.300 ;
        RECT 155.600 307.700 158.800 308.200 ;
        RECT 155.600 307.600 157.200 307.700 ;
        RECT 158.000 307.600 158.800 307.700 ;
        RECT 159.600 307.600 160.400 308.400 ;
        RECT 161.200 308.300 162.000 308.400 ;
        RECT 162.800 308.300 163.400 309.600 ;
        RECT 161.200 307.700 163.500 308.300 ;
        RECT 161.200 307.600 162.000 307.700 ;
        RECT 151.800 306.200 152.400 307.600 ;
        RECT 155.600 307.200 156.400 307.600 ;
        RECT 153.400 306.200 157.000 306.600 ;
        RECT 140.400 302.200 141.200 306.200 ;
        RECT 142.000 306.000 146.000 306.200 ;
        RECT 142.000 302.200 142.800 306.000 ;
        RECT 145.200 302.200 146.000 306.000 ;
        RECT 148.400 305.600 150.200 306.200 ;
        RECT 149.400 304.400 150.200 305.600 ;
        RECT 149.400 303.600 150.800 304.400 ;
        RECT 149.400 302.200 150.200 303.600 ;
        RECT 151.600 302.200 152.400 306.200 ;
        RECT 153.200 306.000 157.200 306.200 ;
        RECT 153.200 302.200 154.000 306.000 ;
        RECT 156.400 302.200 157.200 306.000 ;
        RECT 159.600 304.400 160.200 307.600 ;
        RECT 161.200 304.800 162.000 306.400 ;
        RECT 162.800 306.200 163.400 307.700 ;
        RECT 164.200 307.000 164.800 310.000 ;
        RECT 169.200 309.600 170.000 311.200 ;
        RECT 165.600 308.400 166.400 309.200 ;
        RECT 170.800 308.400 171.400 311.800 ;
        RECT 175.800 311.600 176.400 315.800 ;
        RECT 178.800 311.800 179.600 319.800 ;
        RECT 175.800 311.000 178.200 311.600 ;
        RECT 175.600 309.600 176.400 310.400 ;
        RECT 165.800 308.300 166.800 308.400 ;
        RECT 170.800 308.300 171.600 308.400 ;
        RECT 174.000 308.300 174.800 309.200 ;
        RECT 165.800 307.700 171.600 308.300 ;
        RECT 165.800 307.600 166.800 307.700 ;
        RECT 170.800 307.600 171.600 307.700 ;
        RECT 172.500 307.700 174.800 308.300 ;
        RECT 175.800 308.800 176.400 309.600 ;
        RECT 175.800 308.200 176.800 308.800 ;
        RECT 176.000 308.000 176.800 308.200 ;
        RECT 164.200 306.400 166.600 307.000 ;
        RECT 159.600 302.200 160.400 304.400 ;
        RECT 162.800 302.200 163.600 306.200 ;
        RECT 166.000 304.200 166.600 306.400 ;
        RECT 167.600 306.300 168.400 306.400 ;
        RECT 169.200 306.300 170.000 306.400 ;
        RECT 167.600 305.700 170.000 306.300 ;
        RECT 167.600 304.800 168.400 305.700 ;
        RECT 169.200 305.600 170.000 305.700 ;
        RECT 170.800 304.400 171.400 307.600 ;
        RECT 172.500 306.400 173.100 307.700 ;
        RECT 174.000 307.600 174.800 307.700 ;
        RECT 177.600 307.600 178.200 311.000 ;
        RECT 179.000 310.400 179.600 311.800 ;
        RECT 178.800 309.600 179.600 310.400 ;
        RECT 177.600 307.400 178.400 307.600 ;
        RECT 175.400 307.000 178.400 307.400 ;
        RECT 174.200 306.800 178.400 307.000 ;
        RECT 174.200 306.400 176.000 306.800 ;
        RECT 172.400 304.800 173.200 306.400 ;
        RECT 174.200 306.200 174.800 306.400 ;
        RECT 179.000 306.200 179.600 309.600 ;
        RECT 166.000 302.200 166.800 304.200 ;
        RECT 170.800 302.200 171.600 304.400 ;
        RECT 174.000 302.200 174.800 306.200 ;
        RECT 178.200 305.200 179.600 306.200 ;
        RECT 180.400 311.200 181.200 319.800 ;
        RECT 184.600 315.800 185.800 319.800 ;
        RECT 189.200 315.800 190.000 319.800 ;
        RECT 193.600 316.400 194.400 319.800 ;
        RECT 193.600 315.800 195.600 316.400 ;
        RECT 185.200 315.000 186.000 315.800 ;
        RECT 189.400 315.200 190.000 315.800 ;
        RECT 188.600 314.600 192.200 315.200 ;
        RECT 194.800 315.000 195.600 315.800 ;
        RECT 188.600 314.400 189.400 314.600 ;
        RECT 191.400 314.400 192.200 314.600 ;
        RECT 184.400 313.200 185.800 314.000 ;
        RECT 185.200 312.200 185.800 313.200 ;
        RECT 187.400 313.000 189.600 313.600 ;
        RECT 187.400 312.800 188.200 313.000 ;
        RECT 185.200 311.600 187.600 312.200 ;
        RECT 180.400 310.600 184.600 311.200 ;
        RECT 180.400 307.200 181.200 310.600 ;
        RECT 183.800 310.400 184.600 310.600 ;
        RECT 187.000 310.400 187.600 311.600 ;
        RECT 189.000 311.800 189.600 313.000 ;
        RECT 190.200 313.000 191.000 313.200 ;
        RECT 194.800 313.000 195.600 313.200 ;
        RECT 190.200 312.400 195.600 313.000 ;
        RECT 189.000 311.400 193.800 311.800 ;
        RECT 198.000 311.400 198.800 319.800 ;
        RECT 189.000 311.200 198.800 311.400 ;
        RECT 193.000 311.000 198.800 311.200 ;
        RECT 193.200 310.800 198.800 311.000 ;
        RECT 199.600 311.200 200.400 319.800 ;
        RECT 203.800 315.800 205.000 319.800 ;
        RECT 208.400 315.800 209.200 319.800 ;
        RECT 212.800 316.400 213.600 319.800 ;
        RECT 212.800 315.800 214.800 316.400 ;
        RECT 204.400 315.000 205.200 315.800 ;
        RECT 208.600 315.200 209.200 315.800 ;
        RECT 207.800 314.600 211.400 315.200 ;
        RECT 214.000 315.000 214.800 315.800 ;
        RECT 207.800 314.400 208.600 314.600 ;
        RECT 210.600 314.400 211.400 314.600 ;
        RECT 203.600 313.200 205.000 314.000 ;
        RECT 204.400 312.200 205.000 313.200 ;
        RECT 206.600 313.000 208.800 313.600 ;
        RECT 206.600 312.800 207.400 313.000 ;
        RECT 204.400 311.600 206.800 312.200 ;
        RECT 199.600 310.600 203.800 311.200 ;
        RECT 182.200 309.800 183.000 310.000 ;
        RECT 182.200 309.200 186.000 309.800 ;
        RECT 186.800 309.600 187.600 310.400 ;
        RECT 191.600 310.200 192.400 310.400 ;
        RECT 191.600 309.600 196.600 310.200 ;
        RECT 185.200 309.000 186.000 309.200 ;
        RECT 187.000 308.400 187.600 309.600 ;
        RECT 193.200 309.400 194.000 309.600 ;
        RECT 195.800 309.400 196.600 309.600 ;
        RECT 194.200 308.400 195.000 308.600 ;
        RECT 187.000 307.800 198.000 308.400 ;
        RECT 187.400 307.600 188.200 307.800 ;
        RECT 180.400 306.600 184.200 307.200 ;
        RECT 178.200 304.400 179.000 305.200 ;
        RECT 178.200 303.600 179.600 304.400 ;
        RECT 178.200 302.200 179.000 303.600 ;
        RECT 180.400 302.200 181.200 306.600 ;
        RECT 183.400 306.400 184.200 306.600 ;
        RECT 193.200 305.600 193.800 307.800 ;
        RECT 196.400 307.600 198.000 307.800 ;
        RECT 199.600 307.200 200.400 310.600 ;
        RECT 203.000 310.400 203.800 310.600 ;
        RECT 201.400 309.800 202.200 310.000 ;
        RECT 201.400 309.200 205.200 309.800 ;
        RECT 204.400 309.000 205.200 309.200 ;
        RECT 206.200 308.400 206.800 311.600 ;
        RECT 208.200 311.800 208.800 313.000 ;
        RECT 209.400 313.000 210.200 313.200 ;
        RECT 214.000 313.000 214.800 313.200 ;
        RECT 209.400 312.400 214.800 313.000 ;
        RECT 208.200 311.400 213.000 311.800 ;
        RECT 217.200 311.400 218.000 319.800 ;
        RECT 208.200 311.200 218.000 311.400 ;
        RECT 212.200 311.000 218.000 311.200 ;
        RECT 212.400 310.800 218.000 311.000 ;
        RECT 218.800 311.800 219.600 319.800 ;
        RECT 222.000 312.400 222.800 319.800 ;
        RECT 220.600 311.800 222.800 312.400 ;
        RECT 223.600 311.800 224.400 319.800 ;
        RECT 226.800 312.400 227.600 319.800 ;
        RECT 229.200 313.600 230.000 314.400 ;
        RECT 229.200 312.400 229.800 313.600 ;
        RECT 230.600 312.400 231.400 319.800 ;
        RECT 235.600 313.600 236.400 314.400 ;
        RECT 235.600 312.400 236.200 313.600 ;
        RECT 237.000 312.400 237.800 319.800 ;
        RECT 225.400 311.800 227.600 312.400 ;
        RECT 228.400 311.800 229.800 312.400 ;
        RECT 210.800 310.200 211.600 310.400 ;
        RECT 210.800 309.600 215.800 310.200 ;
        RECT 212.400 309.400 213.200 309.600 ;
        RECT 215.000 309.400 215.800 309.600 ;
        RECT 218.800 309.600 219.400 311.800 ;
        RECT 220.600 311.200 221.200 311.800 ;
        RECT 220.000 310.400 221.200 311.200 ;
        RECT 213.400 308.400 214.200 308.600 ;
        RECT 206.200 307.800 217.200 308.400 ;
        RECT 206.600 307.600 207.400 307.800 ;
        RECT 210.800 307.600 211.600 307.800 ;
        RECT 191.400 305.400 192.200 305.600 ;
        RECT 185.200 304.200 186.000 305.000 ;
        RECT 189.400 304.800 192.200 305.400 ;
        RECT 193.200 304.800 194.000 305.600 ;
        RECT 189.400 304.200 190.000 304.800 ;
        RECT 194.800 304.200 195.600 305.000 ;
        RECT 184.600 303.600 186.000 304.200 ;
        RECT 184.600 302.200 185.800 303.600 ;
        RECT 189.200 302.200 190.000 304.200 ;
        RECT 193.600 303.600 195.600 304.200 ;
        RECT 193.600 302.200 194.400 303.600 ;
        RECT 198.000 302.200 198.800 307.000 ;
        RECT 199.600 306.600 203.400 307.200 ;
        RECT 199.600 302.200 200.400 306.600 ;
        RECT 202.600 306.400 203.400 306.600 ;
        RECT 212.400 305.600 213.000 307.800 ;
        RECT 215.600 307.600 217.200 307.800 ;
        RECT 210.600 305.400 211.400 305.600 ;
        RECT 204.400 304.200 205.200 305.000 ;
        RECT 208.600 304.800 211.400 305.400 ;
        RECT 212.400 304.800 213.200 305.600 ;
        RECT 208.600 304.200 209.200 304.800 ;
        RECT 214.000 304.200 214.800 305.000 ;
        RECT 203.800 303.600 205.200 304.200 ;
        RECT 203.800 302.200 205.000 303.600 ;
        RECT 208.400 302.200 209.200 304.200 ;
        RECT 212.800 303.600 214.800 304.200 ;
        RECT 212.800 302.200 213.600 303.600 ;
        RECT 217.200 302.200 218.000 307.000 ;
        RECT 218.800 302.200 219.600 309.600 ;
        RECT 220.600 307.400 221.200 310.400 ;
        RECT 223.600 309.600 224.200 311.800 ;
        RECT 225.400 311.200 226.000 311.800 ;
        RECT 228.400 311.600 229.200 311.800 ;
        RECT 230.400 311.600 232.400 312.400 ;
        RECT 234.800 311.800 236.200 312.400 ;
        RECT 236.800 311.800 237.800 312.400 ;
        RECT 241.200 311.800 242.000 319.800 ;
        RECT 242.800 312.400 243.600 319.800 ;
        RECT 246.000 312.400 246.800 319.800 ;
        RECT 242.800 311.800 246.800 312.400 ;
        RECT 234.800 311.600 235.600 311.800 ;
        RECT 224.800 310.400 226.000 311.200 ;
        RECT 220.600 306.800 222.800 307.400 ;
        RECT 222.000 302.200 222.800 306.800 ;
        RECT 223.600 302.200 224.400 309.600 ;
        RECT 225.400 307.400 226.000 310.400 ;
        RECT 226.800 310.300 227.600 310.400 ;
        RECT 228.400 310.300 229.200 310.400 ;
        RECT 226.800 309.700 229.200 310.300 ;
        RECT 226.800 308.800 227.600 309.700 ;
        RECT 228.400 309.600 229.200 309.700 ;
        RECT 230.400 308.400 231.000 311.600 ;
        RECT 231.600 308.800 232.400 310.400 ;
        RECT 236.800 308.400 237.400 311.800 ;
        RECT 241.400 310.400 242.000 311.800 ;
        RECT 245.200 310.400 246.000 310.800 ;
        RECT 238.000 310.300 238.800 310.400 ;
        RECT 239.600 310.300 240.400 310.400 ;
        RECT 238.000 309.700 240.400 310.300 ;
        RECT 238.000 308.800 238.800 309.700 ;
        RECT 239.600 309.600 240.400 309.700 ;
        RECT 241.200 309.800 243.600 310.400 ;
        RECT 245.200 310.300 246.800 310.400 ;
        RECT 247.600 310.300 248.400 319.800 ;
        RECT 253.400 312.400 254.200 319.800 ;
        RECT 254.800 313.600 255.600 314.400 ;
        RECT 255.000 312.400 255.600 313.600 ;
        RECT 261.000 312.800 261.800 319.800 ;
        RECT 265.200 315.000 266.000 319.000 ;
        RECT 253.400 311.800 254.400 312.400 ;
        RECT 255.000 311.800 256.400 312.400 ;
        RECT 245.200 309.800 248.400 310.300 ;
        RECT 241.200 309.600 242.000 309.800 ;
        RECT 242.800 309.600 243.600 309.800 ;
        RECT 246.000 309.700 248.400 309.800 ;
        RECT 246.000 309.600 246.800 309.700 ;
        RECT 228.400 307.600 231.000 308.400 ;
        RECT 233.200 308.300 234.000 308.400 ;
        RECT 234.800 308.300 237.400 308.400 ;
        RECT 233.200 308.200 237.400 308.300 ;
        RECT 239.600 308.200 240.400 308.400 ;
        RECT 232.400 307.700 237.400 308.200 ;
        RECT 232.400 307.600 234.000 307.700 ;
        RECT 234.800 307.600 237.400 307.700 ;
        RECT 238.800 307.600 240.400 308.200 ;
        RECT 225.400 306.800 227.600 307.400 ;
        RECT 226.800 302.200 227.600 306.800 ;
        RECT 228.600 306.200 229.200 307.600 ;
        RECT 232.400 307.200 233.200 307.600 ;
        RECT 230.200 306.200 233.800 306.600 ;
        RECT 235.000 306.200 235.600 307.600 ;
        RECT 238.800 307.200 239.600 307.600 ;
        RECT 236.600 306.200 240.200 306.600 ;
        RECT 228.400 302.200 229.200 306.200 ;
        RECT 230.000 306.000 234.000 306.200 ;
        RECT 230.000 302.200 230.800 306.000 ;
        RECT 233.200 302.200 234.000 306.000 ;
        RECT 234.800 302.200 235.600 306.200 ;
        RECT 236.400 306.000 240.400 306.200 ;
        RECT 236.400 302.200 237.200 306.000 ;
        RECT 239.600 302.200 240.400 306.000 ;
        RECT 241.200 305.600 242.000 306.400 ;
        RECT 243.000 306.200 243.600 309.600 ;
        RECT 244.400 307.600 245.200 309.200 ;
        RECT 241.400 304.800 242.200 305.600 ;
        RECT 242.800 302.200 243.600 306.200 ;
        RECT 247.600 302.200 248.400 309.700 ;
        RECT 252.400 308.800 253.200 310.400 ;
        RECT 253.800 310.300 254.400 311.800 ;
        RECT 255.600 311.600 256.400 311.800 ;
        RECT 260.200 312.200 261.800 312.800 ;
        RECT 258.800 310.300 259.600 311.200 ;
        RECT 253.800 309.700 259.600 310.300 ;
        RECT 253.800 308.400 254.400 309.700 ;
        RECT 258.800 309.600 259.600 309.700 ;
        RECT 260.200 308.400 260.800 312.200 ;
        RECT 265.400 311.600 266.000 315.000 ;
        RECT 268.400 312.800 269.200 319.800 ;
        RECT 262.200 311.000 266.000 311.600 ;
        RECT 268.200 311.800 269.200 312.800 ;
        RECT 271.600 312.400 272.400 319.800 ;
        RECT 269.800 311.800 272.400 312.400 ;
        RECT 262.200 309.000 262.800 311.000 ;
        RECT 250.800 308.200 251.600 308.400 ;
        RECT 250.800 307.600 252.400 308.200 ;
        RECT 253.800 307.600 256.400 308.400 ;
        RECT 257.200 308.300 258.000 308.400 ;
        RECT 258.800 308.300 260.800 308.400 ;
        RECT 257.200 307.700 260.800 308.300 ;
        RECT 261.400 308.200 262.800 309.000 ;
        RECT 263.600 308.800 264.400 310.400 ;
        RECT 265.200 310.300 266.000 310.400 ;
        RECT 266.800 310.300 267.600 310.400 ;
        RECT 265.200 309.700 267.600 310.300 ;
        RECT 265.200 308.800 266.000 309.700 ;
        RECT 266.800 309.600 267.600 309.700 ;
        RECT 257.200 307.600 258.000 307.700 ;
        RECT 258.800 307.600 260.800 307.700 ;
        RECT 251.600 307.200 252.400 307.600 ;
        RECT 249.200 304.800 250.000 306.400 ;
        RECT 251.000 306.200 254.600 306.600 ;
        RECT 255.600 306.200 256.200 307.600 ;
        RECT 260.200 307.000 260.800 307.600 ;
        RECT 261.800 307.800 262.800 308.200 ;
        RECT 266.900 308.300 267.500 309.600 ;
        RECT 268.200 308.400 268.800 311.800 ;
        RECT 269.800 309.800 270.400 311.800 ;
        RECT 273.200 311.200 274.000 319.800 ;
        RECT 277.400 315.800 278.600 319.800 ;
        RECT 282.000 315.800 282.800 319.800 ;
        RECT 286.400 316.400 287.200 319.800 ;
        RECT 286.400 315.800 288.400 316.400 ;
        RECT 278.000 315.000 278.800 315.800 ;
        RECT 282.200 315.200 282.800 315.800 ;
        RECT 281.400 314.600 285.000 315.200 ;
        RECT 287.600 315.000 288.400 315.800 ;
        RECT 281.400 314.400 282.200 314.600 ;
        RECT 284.200 314.400 285.000 314.600 ;
        RECT 277.200 313.200 278.600 314.000 ;
        RECT 278.000 312.200 278.600 313.200 ;
        RECT 280.200 313.000 282.400 313.600 ;
        RECT 280.200 312.800 281.000 313.000 ;
        RECT 278.000 311.600 280.400 312.200 ;
        RECT 273.200 310.600 277.400 311.200 ;
        RECT 269.400 309.000 270.400 309.800 ;
        RECT 268.200 308.300 269.200 308.400 ;
        RECT 261.800 307.200 266.000 307.800 ;
        RECT 266.900 307.700 269.200 308.300 ;
        RECT 260.200 306.600 261.000 307.000 ;
        RECT 250.800 306.000 254.800 306.200 ;
        RECT 250.800 302.200 251.600 306.000 ;
        RECT 254.000 302.200 254.800 306.000 ;
        RECT 255.600 302.200 256.400 306.200 ;
        RECT 260.200 306.000 261.800 306.600 ;
        RECT 261.000 303.000 261.800 306.000 ;
        RECT 265.400 305.000 266.000 307.200 ;
        RECT 268.200 307.600 269.200 307.700 ;
        RECT 268.200 306.200 268.800 307.600 ;
        RECT 269.800 307.400 270.400 309.000 ;
        RECT 271.400 309.600 272.400 310.400 ;
        RECT 271.400 308.800 272.200 309.600 ;
        RECT 269.800 306.800 272.400 307.400 ;
        RECT 268.200 305.600 269.200 306.200 ;
        RECT 265.200 303.000 266.000 305.000 ;
        RECT 268.400 302.200 269.200 305.600 ;
        RECT 271.600 302.200 272.400 306.800 ;
        RECT 273.200 307.200 274.000 310.600 ;
        RECT 276.600 310.400 277.400 310.600 ;
        RECT 275.000 309.800 275.800 310.000 ;
        RECT 275.000 309.200 278.800 309.800 ;
        RECT 278.000 309.000 278.800 309.200 ;
        RECT 279.800 308.400 280.400 311.600 ;
        RECT 281.800 311.800 282.400 313.000 ;
        RECT 283.000 313.000 283.800 313.200 ;
        RECT 287.600 313.000 288.400 313.200 ;
        RECT 283.000 312.400 288.400 313.000 ;
        RECT 281.800 311.400 286.600 311.800 ;
        RECT 290.800 311.400 291.600 319.800 ;
        RECT 281.800 311.200 291.600 311.400 ;
        RECT 285.800 311.000 291.600 311.200 ;
        RECT 286.000 310.800 291.600 311.000 ;
        RECT 297.200 311.200 298.000 319.800 ;
        RECT 301.400 315.800 302.600 319.800 ;
        RECT 306.000 315.800 306.800 319.800 ;
        RECT 310.400 316.400 311.200 319.800 ;
        RECT 310.400 315.800 312.400 316.400 ;
        RECT 302.000 315.000 302.800 315.800 ;
        RECT 306.200 315.200 306.800 315.800 ;
        RECT 305.400 314.600 309.000 315.200 ;
        RECT 311.600 315.000 312.400 315.800 ;
        RECT 305.400 314.400 306.200 314.600 ;
        RECT 308.200 314.400 309.000 314.600 ;
        RECT 301.200 313.200 302.600 314.000 ;
        RECT 302.000 312.200 302.600 313.200 ;
        RECT 304.200 313.000 306.400 313.600 ;
        RECT 304.200 312.800 305.000 313.000 ;
        RECT 302.000 311.600 304.400 312.200 ;
        RECT 297.200 310.600 301.400 311.200 ;
        RECT 284.400 310.200 285.200 310.400 ;
        RECT 284.400 309.600 289.400 310.200 ;
        RECT 286.000 309.400 286.800 309.600 ;
        RECT 288.600 309.400 289.400 309.600 ;
        RECT 287.000 308.400 287.800 308.600 ;
        RECT 279.800 308.300 290.800 308.400 ;
        RECT 292.400 308.300 293.200 308.400 ;
        RECT 279.800 307.800 293.200 308.300 ;
        RECT 280.200 307.600 281.000 307.800 ;
        RECT 282.800 307.600 283.600 307.800 ;
        RECT 273.200 306.600 277.000 307.200 ;
        RECT 273.200 302.200 274.000 306.600 ;
        RECT 276.200 306.400 277.000 306.600 ;
        RECT 286.000 305.600 286.600 307.800 ;
        RECT 289.200 307.700 293.200 307.800 ;
        RECT 289.200 307.600 290.800 307.700 ;
        RECT 292.400 307.600 293.200 307.700 ;
        RECT 297.200 307.200 298.000 310.600 ;
        RECT 300.600 310.400 301.400 310.600 ;
        RECT 303.800 310.400 304.400 311.600 ;
        RECT 305.800 311.800 306.400 313.000 ;
        RECT 307.000 313.000 307.800 313.200 ;
        RECT 311.600 313.000 312.400 313.200 ;
        RECT 307.000 312.400 312.400 313.000 ;
        RECT 305.800 311.400 310.600 311.800 ;
        RECT 314.800 311.400 315.600 319.800 ;
        RECT 316.400 312.400 317.200 319.800 ;
        RECT 319.600 312.800 320.400 319.800 ;
        RECT 316.400 311.800 319.000 312.400 ;
        RECT 319.600 311.800 320.600 312.800 ;
        RECT 305.800 311.200 315.600 311.400 ;
        RECT 309.800 311.000 315.600 311.200 ;
        RECT 310.000 310.800 315.600 311.000 ;
        RECT 299.000 309.800 299.800 310.000 ;
        RECT 299.000 309.200 302.800 309.800 ;
        RECT 303.600 309.600 304.400 310.400 ;
        RECT 308.400 310.200 309.200 310.400 ;
        RECT 308.400 309.600 313.400 310.200 ;
        RECT 316.400 309.600 317.400 310.400 ;
        RECT 302.000 309.000 302.800 309.200 ;
        RECT 303.800 308.400 304.400 309.600 ;
        RECT 310.000 309.400 310.800 309.600 ;
        RECT 312.600 309.400 313.400 309.600 ;
        RECT 316.600 308.800 317.400 309.600 ;
        RECT 318.400 309.800 319.000 311.800 ;
        RECT 318.400 309.000 319.400 309.800 ;
        RECT 311.000 308.400 311.800 308.600 ;
        RECT 303.800 307.800 314.800 308.400 ;
        RECT 304.200 307.600 305.000 307.800 ;
        RECT 284.200 305.400 285.000 305.600 ;
        RECT 278.000 304.200 278.800 305.000 ;
        RECT 282.200 304.800 285.000 305.400 ;
        RECT 286.000 304.800 286.800 305.600 ;
        RECT 282.200 304.200 282.800 304.800 ;
        RECT 287.600 304.200 288.400 305.000 ;
        RECT 277.400 303.600 278.800 304.200 ;
        RECT 277.400 302.200 278.600 303.600 ;
        RECT 282.000 302.200 282.800 304.200 ;
        RECT 286.400 303.600 288.400 304.200 ;
        RECT 286.400 302.200 287.200 303.600 ;
        RECT 290.800 302.200 291.600 307.000 ;
        RECT 297.200 306.600 301.000 307.200 ;
        RECT 297.200 302.200 298.000 306.600 ;
        RECT 300.200 306.400 301.000 306.600 ;
        RECT 310.000 305.600 310.600 307.800 ;
        RECT 313.200 307.600 314.800 307.800 ;
        RECT 318.400 307.400 319.000 309.000 ;
        RECT 320.000 308.400 320.600 311.800 ;
        RECT 322.800 311.600 323.600 313.200 ;
        RECT 319.600 308.300 320.600 308.400 ;
        RECT 321.200 308.300 322.000 308.400 ;
        RECT 319.600 307.700 322.000 308.300 ;
        RECT 319.600 307.600 320.600 307.700 ;
        RECT 321.200 307.600 322.000 307.700 ;
        RECT 308.200 305.400 309.000 305.600 ;
        RECT 302.000 304.200 302.800 305.000 ;
        RECT 306.200 304.800 309.000 305.400 ;
        RECT 310.000 304.800 310.800 305.600 ;
        RECT 306.200 304.200 306.800 304.800 ;
        RECT 311.600 304.200 312.400 305.000 ;
        RECT 301.400 303.600 302.800 304.200 ;
        RECT 301.400 302.200 302.600 303.600 ;
        RECT 306.000 302.200 306.800 304.200 ;
        RECT 310.400 303.600 312.400 304.200 ;
        RECT 310.400 302.200 311.200 303.600 ;
        RECT 314.800 302.200 315.600 307.000 ;
        RECT 316.400 306.800 319.000 307.400 ;
        RECT 316.400 302.200 317.200 306.800 ;
        RECT 320.000 306.200 320.600 307.600 ;
        RECT 324.400 306.200 325.200 319.800 ;
        RECT 327.600 311.600 328.400 313.200 ;
        RECT 326.000 308.300 326.800 308.400 ;
        RECT 329.200 308.300 330.000 319.800 ;
        RECT 333.200 313.600 334.000 314.400 ;
        RECT 333.200 312.400 333.800 313.600 ;
        RECT 334.600 312.400 335.400 319.800 ;
        RECT 339.600 313.600 340.400 314.400 ;
        RECT 339.600 312.400 340.200 313.600 ;
        RECT 341.000 312.400 341.800 319.800 ;
        RECT 346.000 313.600 346.800 314.400 ;
        RECT 346.000 312.400 346.600 313.600 ;
        RECT 347.400 312.400 348.200 319.800 ;
        RECT 332.400 311.800 333.800 312.400 ;
        RECT 334.400 311.800 335.400 312.400 ;
        RECT 338.800 311.800 340.200 312.400 ;
        RECT 340.800 311.800 341.800 312.400 ;
        RECT 345.200 311.800 346.600 312.400 ;
        RECT 347.200 311.800 348.200 312.400 ;
        RECT 332.400 311.600 333.200 311.800 ;
        RECT 330.800 310.300 331.600 310.400 ;
        RECT 334.400 310.300 335.000 311.800 ;
        RECT 338.800 311.600 339.600 311.800 ;
        RECT 330.800 309.700 335.000 310.300 ;
        RECT 330.800 309.600 331.600 309.700 ;
        RECT 334.400 308.400 335.000 309.700 ;
        RECT 335.600 310.300 336.400 310.400 ;
        RECT 340.800 310.300 341.400 311.800 ;
        RECT 345.200 311.600 346.000 311.800 ;
        RECT 335.600 309.700 341.400 310.300 ;
        RECT 335.600 308.800 336.400 309.700 ;
        RECT 340.800 308.400 341.400 309.700 ;
        RECT 342.000 308.800 342.800 310.400 ;
        RECT 343.600 310.300 344.400 310.400 ;
        RECT 347.200 310.300 347.800 311.800 ;
        RECT 343.600 309.700 347.800 310.300 ;
        RECT 343.600 309.600 344.400 309.700 ;
        RECT 347.200 308.400 347.800 309.700 ;
        RECT 348.400 308.800 349.200 310.400 ;
        RECT 326.000 307.700 330.000 308.300 ;
        RECT 326.000 306.800 326.800 307.700 ;
        RECT 329.200 306.200 330.000 307.700 ;
        RECT 330.800 306.800 331.600 308.400 ;
        RECT 332.400 307.600 335.000 308.400 ;
        RECT 337.200 308.200 338.000 308.400 ;
        RECT 336.400 307.600 338.000 308.200 ;
        RECT 338.800 307.600 341.400 308.400 ;
        RECT 343.600 308.200 344.400 308.400 ;
        RECT 342.800 307.600 344.400 308.200 ;
        RECT 345.200 307.600 347.800 308.400 ;
        RECT 350.000 308.300 350.800 308.400 ;
        RECT 351.600 308.300 352.400 319.800 ;
        RECT 354.800 312.400 355.600 319.800 ;
        RECT 356.400 312.400 357.200 312.600 ;
        RECT 359.200 312.400 360.800 319.800 ;
        RECT 354.800 311.800 357.200 312.400 ;
        RECT 358.800 311.800 360.800 312.400 ;
        RECT 363.000 312.400 363.800 312.600 ;
        RECT 364.400 312.400 365.200 319.800 ;
        RECT 363.000 311.800 365.200 312.400 ;
        RECT 366.000 312.400 366.800 319.800 ;
        RECT 367.800 312.400 368.600 312.600 ;
        RECT 366.000 311.800 368.600 312.400 ;
        RECT 370.400 311.800 372.000 319.800 ;
        RECT 374.000 312.400 374.800 312.600 ;
        RECT 375.600 312.400 376.400 319.800 ;
        RECT 374.000 311.800 376.400 312.400 ;
        RECT 358.800 310.400 359.400 311.800 ;
        RECT 363.000 311.200 363.600 311.800 ;
        RECT 360.200 310.600 363.600 311.200 ;
        RECT 360.200 310.400 361.000 310.600 ;
        RECT 369.000 310.400 369.800 310.600 ;
        RECT 371.000 310.400 371.600 311.800 ;
        RECT 353.200 310.300 354.000 310.400 ;
        RECT 358.000 310.300 359.400 310.400 ;
        RECT 353.200 309.800 359.400 310.300 ;
        RECT 362.400 309.800 363.200 310.000 ;
        RECT 353.200 309.700 359.800 309.800 ;
        RECT 353.200 309.600 354.000 309.700 ;
        RECT 358.000 309.600 359.800 309.700 ;
        RECT 358.800 309.200 359.800 309.600 ;
        RECT 354.800 308.300 356.400 308.400 ;
        RECT 350.000 308.200 352.400 308.300 ;
        RECT 349.200 307.700 352.400 308.200 ;
        RECT 349.200 307.600 350.800 307.700 ;
        RECT 332.600 306.200 333.200 307.600 ;
        RECT 336.400 307.200 337.200 307.600 ;
        RECT 334.200 306.200 337.800 306.600 ;
        RECT 339.000 306.200 339.600 307.600 ;
        RECT 342.800 307.200 343.600 307.600 ;
        RECT 340.600 306.200 344.200 306.600 ;
        RECT 345.400 306.200 346.000 307.600 ;
        RECT 349.200 307.200 350.000 307.600 ;
        RECT 347.000 306.200 350.600 306.600 ;
        RECT 319.600 305.600 320.600 306.200 ;
        RECT 323.400 305.600 325.200 306.200 ;
        RECT 328.200 305.600 330.000 306.200 ;
        RECT 319.600 302.200 320.400 305.600 ;
        RECT 323.400 304.400 324.200 305.600 ;
        RECT 322.800 303.600 324.200 304.400 ;
        RECT 323.400 302.200 324.200 303.600 ;
        RECT 328.200 302.200 329.000 305.600 ;
        RECT 332.400 302.200 333.200 306.200 ;
        RECT 334.000 306.000 338.000 306.200 ;
        RECT 334.000 302.200 334.800 306.000 ;
        RECT 337.200 302.200 338.000 306.000 ;
        RECT 338.800 302.200 339.600 306.200 ;
        RECT 340.400 306.000 344.400 306.200 ;
        RECT 340.400 302.200 341.200 306.000 ;
        RECT 343.600 302.200 344.400 306.000 ;
        RECT 345.200 302.200 346.000 306.200 ;
        RECT 346.800 306.000 350.800 306.200 ;
        RECT 346.800 302.200 347.600 306.000 ;
        RECT 350.000 302.200 350.800 306.000 ;
        RECT 351.600 302.200 352.400 307.700 ;
        RECT 353.300 307.700 356.400 308.300 ;
        RECT 353.300 306.400 353.900 307.700 ;
        RECT 354.800 307.600 356.400 307.700 ;
        RECT 357.600 307.600 358.400 308.400 ;
        RECT 357.800 307.200 358.400 307.600 ;
        RECT 356.400 306.800 357.200 307.000 ;
        RECT 353.200 304.800 354.000 306.400 ;
        RECT 354.800 306.200 357.200 306.800 ;
        RECT 357.800 306.400 358.600 307.200 ;
        RECT 354.800 302.200 355.600 306.200 ;
        RECT 359.200 305.800 359.800 309.200 ;
        RECT 360.600 309.200 363.200 309.800 ;
        RECT 368.200 309.800 369.800 310.400 ;
        RECT 368.200 309.600 369.000 309.800 ;
        RECT 370.800 309.600 371.600 310.400 ;
        RECT 375.600 310.300 376.400 310.400 ;
        RECT 375.600 309.700 377.900 310.300 ;
        RECT 375.600 309.600 376.400 309.700 ;
        RECT 360.600 308.600 361.200 309.200 ;
        RECT 369.600 308.600 370.400 308.800 ;
        RECT 360.400 307.800 361.200 308.600 ;
        RECT 367.600 308.400 370.400 308.600 ;
        RECT 363.600 308.200 365.200 308.400 ;
        RECT 361.800 307.600 365.200 308.200 ;
        RECT 366.000 308.000 370.400 308.400 ;
        RECT 371.000 308.400 371.600 309.600 ;
        RECT 377.300 308.400 377.900 309.700 ;
        RECT 366.000 307.800 368.200 308.000 ;
        RECT 371.000 307.800 372.000 308.400 ;
        RECT 366.000 307.600 367.600 307.800 ;
        RECT 361.800 307.200 362.400 307.600 ;
        RECT 360.400 306.600 362.400 307.200 ;
        RECT 363.000 306.800 363.800 307.000 ;
        RECT 367.800 306.800 368.600 307.000 ;
        RECT 360.400 306.400 362.000 306.600 ;
        RECT 363.000 306.200 365.200 306.800 ;
        RECT 359.200 302.200 360.800 305.800 ;
        RECT 364.400 302.200 365.200 306.200 ;
        RECT 366.000 306.200 368.600 306.800 ;
        RECT 369.200 306.400 370.800 307.200 ;
        RECT 366.000 302.200 366.800 306.200 ;
        RECT 371.400 305.800 372.000 307.800 ;
        RECT 372.800 307.600 373.600 308.400 ;
        RECT 374.800 307.600 376.400 308.400 ;
        RECT 372.800 307.200 373.400 307.600 ;
        RECT 372.600 306.400 373.400 307.200 ;
        RECT 374.000 306.800 374.800 307.000 ;
        RECT 377.200 306.800 378.000 308.400 ;
        RECT 374.000 306.200 376.400 306.800 ;
        RECT 370.400 304.400 372.000 305.800 ;
        RECT 369.200 303.600 372.000 304.400 ;
        RECT 370.400 302.200 372.000 303.600 ;
        RECT 375.600 302.200 376.400 306.200 ;
        RECT 378.800 306.200 379.600 319.800 ;
        RECT 380.400 311.600 381.200 313.200 ;
        RECT 384.600 312.600 385.400 319.800 ;
        RECT 383.600 311.800 385.400 312.600 ;
        RECT 389.400 311.800 391.400 319.800 ;
        RECT 380.500 310.400 381.100 311.600 ;
        RECT 380.400 310.300 381.200 310.400 ;
        RECT 383.800 310.300 384.400 311.800 ;
        RECT 380.400 309.700 384.400 310.300 ;
        RECT 380.400 309.600 381.200 309.700 ;
        RECT 383.800 308.400 384.400 309.700 ;
        RECT 385.200 309.600 386.000 311.200 ;
        RECT 383.600 307.600 384.400 308.400 ;
        RECT 386.800 307.600 387.600 309.200 ;
        RECT 388.400 308.800 389.200 310.400 ;
        RECT 390.200 308.400 390.800 311.800 ;
        RECT 391.600 308.800 392.400 310.400 ;
        RECT 390.000 308.200 390.800 308.400 ;
        RECT 393.200 308.300 394.000 308.400 ;
        RECT 394.800 308.300 395.600 319.800 ;
        RECT 398.600 312.400 399.400 319.800 ;
        RECT 398.000 311.800 399.400 312.400 ;
        RECT 398.000 310.400 398.600 311.800 ;
        RECT 402.800 311.200 403.600 319.800 ;
        RECT 399.600 310.800 403.600 311.200 ;
        RECT 399.400 310.600 403.600 310.800 ;
        RECT 404.400 311.200 405.200 319.800 ;
        RECT 408.600 315.800 409.800 319.800 ;
        RECT 413.200 315.800 414.000 319.800 ;
        RECT 417.600 316.400 418.400 319.800 ;
        RECT 417.600 315.800 419.600 316.400 ;
        RECT 409.200 315.000 410.000 315.800 ;
        RECT 413.400 315.200 414.000 315.800 ;
        RECT 412.600 314.600 416.200 315.200 ;
        RECT 418.800 315.000 419.600 315.800 ;
        RECT 412.600 314.400 413.400 314.600 ;
        RECT 415.400 314.400 416.200 314.600 ;
        RECT 408.400 313.200 409.800 314.000 ;
        RECT 409.200 312.200 409.800 313.200 ;
        RECT 411.400 313.000 413.600 313.600 ;
        RECT 411.400 312.800 412.200 313.000 ;
        RECT 409.200 311.600 411.600 312.200 ;
        RECT 404.400 310.600 408.600 311.200 ;
        RECT 396.400 310.300 397.200 310.400 ;
        RECT 398.000 310.300 398.800 310.400 ;
        RECT 396.400 309.700 398.800 310.300 ;
        RECT 396.400 309.600 397.200 309.700 ;
        RECT 398.000 309.600 398.800 309.700 ;
        RECT 399.400 310.000 400.200 310.600 ;
        RECT 393.200 308.200 395.600 308.300 ;
        RECT 388.400 307.600 390.800 308.200 ;
        RECT 392.400 307.700 395.600 308.200 ;
        RECT 392.400 307.600 394.000 307.700 ;
        RECT 378.800 305.600 380.600 306.200 ;
        RECT 379.800 302.200 380.600 305.600 ;
        RECT 382.000 304.800 382.800 306.400 ;
        RECT 383.800 304.200 384.400 307.600 ;
        RECT 388.400 306.400 389.000 307.600 ;
        RECT 392.400 307.200 393.200 307.600 ;
        RECT 383.600 302.200 384.400 304.200 ;
        RECT 386.800 302.800 387.600 306.200 ;
        RECT 388.400 303.400 389.200 306.400 ;
        RECT 390.200 306.200 393.800 306.600 ;
        RECT 390.000 306.000 394.000 306.200 ;
        RECT 390.000 302.800 390.800 306.000 ;
        RECT 386.800 302.200 390.800 302.800 ;
        RECT 393.200 302.200 394.000 306.000 ;
        RECT 394.800 302.200 395.600 307.700 ;
        RECT 396.400 304.800 397.200 306.400 ;
        RECT 398.000 306.200 398.600 309.600 ;
        RECT 399.400 307.000 400.000 310.000 ;
        RECT 400.800 308.400 401.600 309.200 ;
        RECT 401.000 307.600 402.000 308.400 ;
        RECT 404.400 307.200 405.200 310.600 ;
        RECT 407.800 310.400 408.600 310.600 ;
        RECT 411.000 310.400 411.600 311.600 ;
        RECT 413.000 311.800 413.600 313.000 ;
        RECT 414.200 313.000 415.000 313.200 ;
        RECT 418.800 313.000 419.600 313.200 ;
        RECT 414.200 312.400 419.600 313.000 ;
        RECT 413.000 311.400 417.800 311.800 ;
        RECT 422.000 311.400 422.800 319.800 ;
        RECT 423.600 319.200 427.600 319.800 ;
        RECT 423.600 311.800 424.400 319.200 ;
        RECT 425.200 311.800 426.000 318.600 ;
        RECT 426.800 312.400 427.600 319.200 ;
        RECT 430.000 312.400 430.800 319.800 ;
        RECT 426.800 311.800 430.800 312.400 ;
        RECT 433.200 312.300 434.000 319.800 ;
        RECT 435.600 313.600 436.400 314.400 ;
        RECT 435.600 312.400 436.200 313.600 ;
        RECT 437.000 312.400 437.800 319.800 ;
        RECT 434.800 312.300 436.200 312.400 ;
        RECT 433.200 311.800 436.200 312.300 ;
        RECT 436.800 311.800 437.800 312.400 ;
        RECT 413.000 311.200 422.800 311.400 ;
        RECT 425.400 311.200 426.000 311.800 ;
        RECT 433.200 311.700 435.600 311.800 ;
        RECT 417.000 311.000 422.800 311.200 ;
        RECT 417.200 310.800 422.800 311.000 ;
        RECT 406.200 309.800 407.000 310.000 ;
        RECT 406.200 309.200 410.000 309.800 ;
        RECT 410.800 309.600 411.600 310.400 ;
        RECT 415.600 310.200 416.400 310.400 ;
        RECT 415.600 309.600 420.600 310.200 ;
        RECT 423.600 309.600 424.400 311.200 ;
        RECT 425.400 310.600 427.400 311.200 ;
        RECT 426.800 310.400 427.400 310.600 ;
        RECT 429.200 310.400 430.000 310.800 ;
        RECT 426.800 309.600 427.600 310.400 ;
        RECT 429.200 309.800 430.800 310.400 ;
        RECT 430.000 309.600 430.800 309.800 ;
        RECT 409.200 309.000 410.000 309.200 ;
        RECT 411.000 308.400 411.600 309.600 ;
        RECT 417.200 309.400 418.000 309.600 ;
        RECT 419.800 309.400 420.600 309.600 ;
        RECT 425.400 308.800 426.200 309.600 ;
        RECT 418.200 308.400 419.000 308.600 ;
        RECT 425.400 308.400 426.000 308.800 ;
        RECT 411.000 307.800 422.000 308.400 ;
        RECT 411.400 307.600 412.200 307.800 ;
        RECT 399.400 306.400 401.800 307.000 ;
        RECT 404.400 306.600 408.200 307.200 ;
        RECT 398.000 302.200 398.800 306.200 ;
        RECT 401.200 304.200 401.800 306.400 ;
        RECT 402.800 304.800 403.600 306.400 ;
        RECT 401.200 302.200 402.000 304.200 ;
        RECT 404.400 302.200 405.200 306.600 ;
        RECT 407.400 306.400 408.200 306.600 ;
        RECT 417.200 305.600 417.800 307.800 ;
        RECT 420.400 307.600 422.000 307.800 ;
        RECT 425.200 307.600 426.000 308.400 ;
        RECT 415.400 305.400 416.200 305.600 ;
        RECT 409.200 304.200 410.000 305.000 ;
        RECT 413.400 304.800 416.200 305.400 ;
        RECT 417.200 304.800 418.000 305.600 ;
        RECT 413.400 304.200 414.000 304.800 ;
        RECT 418.800 304.200 419.600 305.000 ;
        RECT 408.600 303.600 410.000 304.200 ;
        RECT 408.600 302.200 409.800 303.600 ;
        RECT 413.200 302.200 414.000 304.200 ;
        RECT 417.600 303.600 419.600 304.200 ;
        RECT 417.600 302.200 418.400 303.600 ;
        RECT 422.000 302.200 422.800 307.000 ;
        RECT 426.800 306.200 427.400 309.600 ;
        RECT 428.400 308.300 429.200 309.200 ;
        RECT 428.400 307.700 432.300 308.300 ;
        RECT 428.400 307.600 429.200 307.700 ;
        RECT 431.700 306.400 432.300 307.700 ;
        RECT 426.200 304.400 427.800 306.200 ;
        RECT 431.600 304.800 432.400 306.400 ;
        RECT 425.200 303.600 427.800 304.400 ;
        RECT 426.200 302.200 427.800 303.600 ;
        RECT 433.200 302.200 434.000 311.700 ;
        RECT 434.800 311.600 435.600 311.700 ;
        RECT 434.800 310.300 435.600 310.400 ;
        RECT 436.800 310.300 437.400 311.800 ;
        RECT 434.800 309.700 437.400 310.300 ;
        RECT 434.800 309.600 435.600 309.700 ;
        RECT 436.800 308.400 437.400 309.700 ;
        RECT 438.000 308.800 438.800 310.400 ;
        RECT 439.600 310.300 440.400 310.400 ;
        RECT 442.800 310.300 443.600 319.800 ;
        RECT 444.400 311.600 445.200 313.200 ;
        RECT 439.600 309.700 443.600 310.300 ;
        RECT 439.600 309.600 440.400 309.700 ;
        RECT 434.800 307.600 437.400 308.400 ;
        RECT 439.600 308.300 440.400 308.400 ;
        RECT 441.200 308.300 442.000 308.400 ;
        RECT 439.600 308.200 442.000 308.300 ;
        RECT 438.800 307.700 442.000 308.200 ;
        RECT 438.800 307.600 440.400 307.700 ;
        RECT 435.000 306.200 435.600 307.600 ;
        RECT 438.800 307.200 439.600 307.600 ;
        RECT 441.200 306.800 442.000 307.700 ;
        RECT 436.600 306.200 440.200 306.600 ;
        RECT 442.800 306.200 443.600 309.700 ;
        RECT 452.400 310.300 453.200 319.800 ;
        RECT 456.400 313.600 457.200 314.400 ;
        RECT 454.000 311.600 454.800 313.200 ;
        RECT 456.400 312.400 457.000 313.600 ;
        RECT 457.800 312.400 458.600 319.800 ;
        RECT 455.600 311.800 457.000 312.400 ;
        RECT 457.600 311.800 458.600 312.400 ;
        RECT 455.600 311.600 456.400 311.800 ;
        RECT 455.700 310.300 456.300 311.600 ;
        RECT 457.600 310.400 458.200 311.800 ;
        RECT 452.400 309.700 456.300 310.300 ;
        RECT 450.800 306.800 451.600 308.400 ;
        RECT 452.400 306.200 453.200 309.700 ;
        RECT 457.200 309.600 458.200 310.400 ;
        RECT 457.600 308.400 458.200 309.600 ;
        RECT 458.800 308.800 459.600 310.400 ;
        RECT 455.600 307.600 458.200 308.400 ;
        RECT 460.400 308.200 461.200 308.400 ;
        RECT 459.600 307.600 461.200 308.200 ;
        RECT 455.800 306.200 456.400 307.600 ;
        RECT 459.600 307.200 460.400 307.600 ;
        RECT 457.400 306.200 461.000 306.600 ;
        RECT 434.800 302.200 435.600 306.200 ;
        RECT 436.400 306.000 440.400 306.200 ;
        RECT 436.400 302.200 437.200 306.000 ;
        RECT 439.600 302.200 440.400 306.000 ;
        RECT 442.800 305.600 444.600 306.200 ;
        RECT 452.400 305.600 454.200 306.200 ;
        RECT 443.800 304.300 444.600 305.600 ;
        RECT 449.200 304.300 450.000 304.400 ;
        RECT 443.800 303.700 450.000 304.300 ;
        RECT 443.800 302.200 444.600 303.700 ;
        RECT 449.200 303.600 450.000 303.700 ;
        RECT 453.400 302.200 454.200 305.600 ;
        RECT 455.600 302.200 456.400 306.200 ;
        RECT 457.200 306.000 461.200 306.200 ;
        RECT 457.200 302.200 458.000 306.000 ;
        RECT 460.400 302.200 461.200 306.000 ;
        RECT 462.000 302.200 462.800 319.800 ;
        RECT 465.200 312.400 466.000 319.800 ;
        RECT 469.600 318.400 471.200 319.800 ;
        RECT 468.400 317.600 471.200 318.400 ;
        RECT 466.800 312.400 467.600 312.600 ;
        RECT 469.600 312.400 471.200 317.600 ;
        RECT 465.200 311.800 467.600 312.400 ;
        RECT 469.200 311.800 471.200 312.400 ;
        RECT 473.400 312.400 474.200 312.600 ;
        RECT 474.800 312.400 475.600 319.800 ;
        RECT 473.400 311.800 475.600 312.400 ;
        RECT 469.200 310.400 469.800 311.800 ;
        RECT 473.400 311.200 474.000 311.800 ;
        RECT 470.600 310.600 474.000 311.200 ;
        RECT 470.600 310.400 471.400 310.600 ;
        RECT 468.400 309.800 469.800 310.400 ;
        RECT 472.800 309.800 473.600 310.000 ;
        RECT 468.400 309.600 470.200 309.800 ;
        RECT 469.200 309.200 470.200 309.600 ;
        RECT 463.600 308.300 464.400 308.400 ;
        RECT 465.200 308.300 466.800 308.400 ;
        RECT 463.600 307.700 466.800 308.300 ;
        RECT 463.600 307.600 464.400 307.700 ;
        RECT 465.200 307.600 466.800 307.700 ;
        RECT 468.000 307.600 468.800 308.400 ;
        RECT 463.700 306.400 464.300 307.600 ;
        RECT 468.200 307.200 468.800 307.600 ;
        RECT 466.800 306.800 467.600 307.000 ;
        RECT 463.600 304.800 464.400 306.400 ;
        RECT 465.200 306.200 467.600 306.800 ;
        RECT 468.200 306.400 469.000 307.200 ;
        RECT 465.200 302.200 466.000 306.200 ;
        RECT 469.600 305.800 470.200 309.200 ;
        RECT 471.000 309.200 473.600 309.800 ;
        RECT 471.000 308.600 471.600 309.200 ;
        RECT 470.800 307.800 471.600 308.600 ;
        RECT 474.000 308.200 475.600 308.400 ;
        RECT 472.200 307.600 475.600 308.200 ;
        RECT 472.200 307.200 472.800 307.600 ;
        RECT 470.800 306.600 472.800 307.200 ;
        RECT 473.400 306.800 474.200 307.000 ;
        RECT 470.800 306.400 472.400 306.600 ;
        RECT 473.400 306.200 475.600 306.800 ;
        RECT 469.600 302.200 471.200 305.800 ;
        RECT 474.800 302.200 475.600 306.200 ;
        RECT 476.400 302.200 477.200 319.800 ;
        RECT 479.600 311.400 480.400 319.800 ;
        RECT 484.000 316.400 484.800 319.800 ;
        RECT 482.800 315.800 484.800 316.400 ;
        RECT 488.400 315.800 489.200 319.800 ;
        RECT 492.600 315.800 493.800 319.800 ;
        RECT 482.800 315.000 483.600 315.800 ;
        RECT 488.400 315.200 489.000 315.800 ;
        RECT 486.200 314.600 489.800 315.200 ;
        RECT 492.400 315.000 493.200 315.800 ;
        RECT 486.200 314.400 487.000 314.600 ;
        RECT 489.000 314.400 489.800 314.600 ;
        RECT 482.800 313.000 483.600 313.200 ;
        RECT 487.400 313.000 488.200 313.200 ;
        RECT 482.800 312.400 488.200 313.000 ;
        RECT 488.800 313.000 491.000 313.600 ;
        RECT 488.800 311.800 489.400 313.000 ;
        RECT 490.200 312.800 491.000 313.000 ;
        RECT 492.600 313.200 494.000 314.000 ;
        RECT 492.600 312.200 493.200 313.200 ;
        RECT 484.600 311.400 489.400 311.800 ;
        RECT 479.600 311.200 489.400 311.400 ;
        RECT 490.800 311.600 493.200 312.200 ;
        RECT 479.600 311.000 485.400 311.200 ;
        RECT 479.600 310.800 485.200 311.000 ;
        RECT 486.000 310.200 486.800 310.400 ;
        RECT 481.800 309.600 486.800 310.200 ;
        RECT 481.800 309.400 482.600 309.600 ;
        RECT 484.400 309.400 485.200 309.600 ;
        RECT 483.400 308.400 484.200 308.600 ;
        RECT 490.800 308.400 491.400 311.600 ;
        RECT 497.200 311.200 498.000 319.800 ;
        RECT 500.400 312.000 501.200 319.800 ;
        RECT 503.600 315.200 504.400 319.800 ;
        RECT 493.800 310.600 498.000 311.200 ;
        RECT 493.800 310.400 494.600 310.600 ;
        RECT 495.400 309.800 496.200 310.000 ;
        RECT 492.400 309.200 496.200 309.800 ;
        RECT 492.400 309.000 493.200 309.200 ;
        RECT 480.400 307.800 491.400 308.400 ;
        RECT 480.400 307.600 482.000 307.800 ;
        RECT 478.000 304.800 478.800 306.400 ;
        RECT 479.600 302.200 480.400 307.000 ;
        RECT 484.600 305.600 485.200 307.800 ;
        RECT 487.600 307.600 488.400 307.800 ;
        RECT 490.200 307.600 491.000 307.800 ;
        RECT 497.200 307.200 498.000 310.600 ;
        RECT 494.200 306.600 498.000 307.200 ;
        RECT 494.200 306.400 495.000 306.600 ;
        RECT 482.800 304.200 483.600 305.000 ;
        RECT 484.400 304.800 485.200 305.600 ;
        RECT 486.200 305.400 487.000 305.600 ;
        RECT 486.200 304.800 489.000 305.400 ;
        RECT 488.400 304.200 489.000 304.800 ;
        RECT 492.400 304.200 493.200 305.000 ;
        RECT 482.800 303.600 484.800 304.200 ;
        RECT 484.000 302.200 484.800 303.600 ;
        RECT 488.400 302.200 489.200 304.200 ;
        RECT 492.400 303.600 493.800 304.200 ;
        RECT 492.600 302.200 493.800 303.600 ;
        RECT 497.200 302.200 498.000 306.600 ;
        RECT 500.200 311.200 501.200 312.000 ;
        RECT 501.800 314.600 504.400 315.200 ;
        RECT 501.800 313.000 502.400 314.600 ;
        RECT 506.800 314.400 507.600 319.800 ;
        RECT 510.000 317.000 510.800 319.800 ;
        RECT 511.600 317.000 512.400 319.800 ;
        RECT 513.200 317.000 514.000 319.800 ;
        RECT 508.200 314.400 512.400 315.200 ;
        RECT 505.000 313.600 507.600 314.400 ;
        RECT 514.800 313.600 515.600 319.800 ;
        RECT 518.000 315.000 518.800 319.800 ;
        RECT 521.200 315.000 522.000 319.800 ;
        RECT 522.800 317.000 523.600 319.800 ;
        RECT 524.400 317.000 525.200 319.800 ;
        RECT 527.600 315.200 528.400 319.800 ;
        RECT 530.800 316.400 531.600 319.800 ;
        RECT 530.800 315.800 531.800 316.400 ;
        RECT 531.200 315.200 531.800 315.800 ;
        RECT 526.400 314.400 530.600 315.200 ;
        RECT 531.200 314.600 533.200 315.200 ;
        RECT 518.000 313.600 520.600 314.400 ;
        RECT 521.200 313.800 527.000 314.400 ;
        RECT 530.000 314.000 530.600 314.400 ;
        RECT 510.000 313.000 510.800 313.200 ;
        RECT 501.800 312.400 510.800 313.000 ;
        RECT 513.200 313.000 514.000 313.200 ;
        RECT 521.200 313.000 521.800 313.800 ;
        RECT 527.600 313.200 529.000 313.800 ;
        RECT 530.000 313.200 531.600 314.000 ;
        RECT 513.200 312.400 521.800 313.000 ;
        RECT 522.800 313.000 529.000 313.200 ;
        RECT 522.800 312.600 528.200 313.000 ;
        RECT 522.800 312.400 523.600 312.600 ;
        RECT 500.200 306.800 501.000 311.200 ;
        RECT 501.800 310.600 502.400 312.400 ;
        RECT 525.800 311.800 526.600 312.000 ;
        RECT 529.200 311.800 530.000 312.400 ;
        RECT 503.000 311.200 530.000 311.800 ;
        RECT 503.000 311.000 503.800 311.200 ;
        RECT 501.600 310.000 502.400 310.600 ;
        RECT 508.400 310.000 531.800 310.600 ;
        RECT 501.600 308.000 502.200 310.000 ;
        RECT 508.400 309.400 509.200 310.000 ;
        RECT 526.000 309.600 526.800 310.000 ;
        RECT 529.200 309.600 530.000 310.000 ;
        RECT 531.000 309.800 531.800 310.000 ;
        RECT 502.800 308.600 506.600 309.400 ;
        RECT 501.600 307.400 502.800 308.000 ;
        RECT 500.200 306.000 501.200 306.800 ;
        RECT 500.400 302.200 501.200 306.000 ;
        RECT 502.000 302.200 502.800 307.400 ;
        RECT 505.800 307.400 506.600 308.600 ;
        RECT 505.800 306.800 507.600 307.400 ;
        RECT 506.800 306.200 507.600 306.800 ;
        RECT 511.600 306.400 512.400 309.200 ;
        RECT 514.800 308.600 518.000 309.400 ;
        RECT 521.800 308.600 523.800 309.400 ;
        RECT 532.400 309.000 533.200 314.600 ;
        RECT 514.400 307.800 515.200 308.000 ;
        RECT 514.400 307.200 518.800 307.800 ;
        RECT 518.000 307.000 518.800 307.200 ;
        RECT 506.800 305.400 509.200 306.200 ;
        RECT 511.600 305.600 512.600 306.400 ;
        RECT 515.600 305.600 517.200 306.400 ;
        RECT 518.000 306.200 518.800 306.400 ;
        RECT 521.800 306.200 522.600 308.600 ;
        RECT 524.400 308.200 533.200 309.000 ;
        RECT 527.800 306.800 530.800 307.600 ;
        RECT 527.800 306.200 528.600 306.800 ;
        RECT 518.000 305.600 522.600 306.200 ;
        RECT 508.400 302.200 509.200 305.400 ;
        RECT 526.000 305.400 528.600 306.200 ;
        RECT 510.000 302.200 510.800 305.000 ;
        RECT 511.600 302.200 512.400 305.000 ;
        RECT 513.200 302.200 514.000 305.000 ;
        RECT 514.800 302.200 515.600 305.000 ;
        RECT 518.000 302.200 518.800 305.000 ;
        RECT 521.200 302.200 522.000 305.000 ;
        RECT 522.800 302.200 523.600 305.000 ;
        RECT 524.400 302.200 525.200 305.000 ;
        RECT 526.000 302.200 526.800 305.400 ;
        RECT 532.400 302.200 533.200 308.200 ;
        RECT 535.600 306.200 536.400 319.800 ;
        RECT 539.400 312.400 540.200 319.800 ;
        RECT 538.800 311.800 540.200 312.400 ;
        RECT 538.800 310.400 539.400 311.800 ;
        RECT 543.600 311.200 544.400 319.800 ;
        RECT 540.400 310.800 544.400 311.200 ;
        RECT 545.200 311.400 546.000 319.800 ;
        RECT 549.600 316.400 550.400 319.800 ;
        RECT 548.400 315.800 550.400 316.400 ;
        RECT 554.000 315.800 554.800 319.800 ;
        RECT 558.200 315.800 559.400 319.800 ;
        RECT 548.400 315.000 549.200 315.800 ;
        RECT 554.000 315.200 554.600 315.800 ;
        RECT 551.800 314.600 555.400 315.200 ;
        RECT 558.000 315.000 558.800 315.800 ;
        RECT 551.800 314.400 552.600 314.600 ;
        RECT 554.600 314.400 555.400 314.600 ;
        RECT 548.400 313.000 549.200 313.200 ;
        RECT 553.000 313.000 553.800 313.200 ;
        RECT 548.400 312.400 553.800 313.000 ;
        RECT 554.400 313.000 556.600 313.600 ;
        RECT 554.400 311.800 555.000 313.000 ;
        RECT 555.800 312.800 556.600 313.000 ;
        RECT 558.200 313.200 559.600 314.000 ;
        RECT 558.200 312.200 558.800 313.200 ;
        RECT 550.200 311.400 555.000 311.800 ;
        RECT 545.200 311.200 555.000 311.400 ;
        RECT 556.400 311.600 558.800 312.200 ;
        RECT 545.200 311.000 551.000 311.200 ;
        RECT 545.200 310.800 550.800 311.000 ;
        RECT 540.200 310.600 544.400 310.800 ;
        RECT 537.200 310.300 538.000 310.400 ;
        RECT 538.800 310.300 539.600 310.400 ;
        RECT 537.200 309.700 539.600 310.300 ;
        RECT 537.200 309.600 538.000 309.700 ;
        RECT 538.800 309.600 539.600 309.700 ;
        RECT 540.200 310.000 541.000 310.600 ;
        RECT 551.600 310.200 552.400 310.400 ;
        RECT 534.600 305.600 536.400 306.200 ;
        RECT 538.800 306.200 539.400 309.600 ;
        RECT 540.200 307.000 540.800 310.000 ;
        RECT 547.400 309.600 552.400 310.200 ;
        RECT 547.400 309.400 548.200 309.600 ;
        RECT 550.000 309.400 550.800 309.600 ;
        RECT 549.000 308.400 549.800 308.600 ;
        RECT 556.400 308.400 557.000 311.600 ;
        RECT 562.800 311.200 563.600 319.800 ;
        RECT 559.400 310.600 563.600 311.200 ;
        RECT 564.400 311.400 565.200 319.800 ;
        RECT 568.800 316.400 569.600 319.800 ;
        RECT 567.600 315.800 569.600 316.400 ;
        RECT 573.200 315.800 574.000 319.800 ;
        RECT 577.400 315.800 578.600 319.800 ;
        RECT 567.600 315.000 568.400 315.800 ;
        RECT 573.200 315.200 573.800 315.800 ;
        RECT 571.000 314.600 574.600 315.200 ;
        RECT 577.200 315.000 578.000 315.800 ;
        RECT 571.000 314.400 571.800 314.600 ;
        RECT 573.800 314.400 574.600 314.600 ;
        RECT 567.600 313.000 568.400 313.200 ;
        RECT 572.200 313.000 573.000 313.200 ;
        RECT 567.600 312.400 573.000 313.000 ;
        RECT 573.600 313.000 575.800 313.600 ;
        RECT 573.600 311.800 574.200 313.000 ;
        RECT 575.000 312.800 575.800 313.000 ;
        RECT 577.400 313.200 578.800 314.000 ;
        RECT 577.400 312.200 578.000 313.200 ;
        RECT 569.400 311.400 574.200 311.800 ;
        RECT 564.400 311.200 574.200 311.400 ;
        RECT 575.600 311.600 578.000 312.200 ;
        RECT 564.400 311.000 570.200 311.200 ;
        RECT 564.400 310.800 570.000 311.000 ;
        RECT 559.400 310.400 560.200 310.600 ;
        RECT 561.000 309.800 561.800 310.000 ;
        RECT 558.000 309.200 561.800 309.800 ;
        RECT 558.000 309.000 558.800 309.200 ;
        RECT 546.000 307.800 557.000 308.400 ;
        RECT 546.000 307.600 547.600 307.800 ;
        RECT 540.200 306.400 542.600 307.000 ;
        RECT 534.600 302.200 535.400 305.600 ;
        RECT 538.800 302.200 539.600 306.200 ;
        RECT 542.000 304.200 542.600 306.400 ;
        RECT 543.600 304.800 544.400 306.400 ;
        RECT 542.000 302.200 542.800 304.200 ;
        RECT 545.200 302.200 546.000 307.000 ;
        RECT 550.200 305.600 550.800 307.800 ;
        RECT 551.600 307.600 552.400 307.800 ;
        RECT 555.800 307.600 556.600 307.800 ;
        RECT 562.800 307.200 563.600 310.600 ;
        RECT 570.800 310.200 571.600 310.400 ;
        RECT 566.600 309.600 571.600 310.200 ;
        RECT 566.600 309.400 567.400 309.600 ;
        RECT 569.200 309.400 570.000 309.600 ;
        RECT 568.200 308.400 569.000 308.600 ;
        RECT 575.600 308.400 576.200 311.600 ;
        RECT 582.000 311.200 582.800 319.800 ;
        RECT 578.600 310.600 582.800 311.200 ;
        RECT 578.600 310.400 579.400 310.600 ;
        RECT 580.200 309.800 581.000 310.000 ;
        RECT 577.200 309.200 581.000 309.800 ;
        RECT 577.200 309.000 578.000 309.200 ;
        RECT 565.200 307.800 576.200 308.400 ;
        RECT 565.200 307.600 566.800 307.800 ;
        RECT 559.800 306.600 563.600 307.200 ;
        RECT 559.800 306.400 560.600 306.600 ;
        RECT 548.400 304.200 549.200 305.000 ;
        RECT 550.000 304.800 550.800 305.600 ;
        RECT 551.800 305.400 552.600 305.600 ;
        RECT 551.800 304.800 554.600 305.400 ;
        RECT 554.000 304.200 554.600 304.800 ;
        RECT 558.000 304.200 558.800 305.000 ;
        RECT 548.400 303.600 550.400 304.200 ;
        RECT 549.600 302.200 550.400 303.600 ;
        RECT 554.000 302.200 554.800 304.200 ;
        RECT 558.000 303.600 559.400 304.200 ;
        RECT 558.200 302.200 559.400 303.600 ;
        RECT 562.800 302.200 563.600 306.600 ;
        RECT 564.400 302.200 565.200 307.000 ;
        RECT 569.400 305.600 570.000 307.800 ;
        RECT 575.000 307.600 575.800 307.800 ;
        RECT 582.000 307.200 582.800 310.600 ;
        RECT 579.000 306.600 582.800 307.200 ;
        RECT 579.000 306.400 579.800 306.600 ;
        RECT 567.600 304.200 568.400 305.000 ;
        RECT 569.200 304.800 570.000 305.600 ;
        RECT 571.000 305.400 571.800 305.600 ;
        RECT 571.000 304.800 573.800 305.400 ;
        RECT 573.200 304.200 573.800 304.800 ;
        RECT 577.200 304.200 578.000 305.000 ;
        RECT 567.600 303.600 569.600 304.200 ;
        RECT 568.800 302.200 569.600 303.600 ;
        RECT 573.200 302.200 574.000 304.200 ;
        RECT 577.200 303.600 578.600 304.200 ;
        RECT 577.400 302.200 578.600 303.600 ;
        RECT 582.000 302.200 582.800 306.600 ;
        RECT 1.200 295.600 2.000 297.200 ;
        RECT 2.800 282.200 3.600 299.800 ;
        RECT 4.400 282.200 5.200 299.800 ;
        RECT 6.000 295.600 6.800 297.200 ;
        RECT 7.600 295.800 8.400 299.800 ;
        RECT 9.200 296.000 10.000 299.800 ;
        RECT 12.400 296.000 13.200 299.800 ;
        RECT 9.200 295.800 13.200 296.000 ;
        RECT 7.800 294.400 8.400 295.800 ;
        RECT 9.400 295.400 13.000 295.800 ;
        RECT 11.600 294.400 12.400 294.800 ;
        RECT 7.600 293.600 10.200 294.400 ;
        RECT 11.600 293.800 13.200 294.400 ;
        RECT 15.200 294.200 16.000 299.800 ;
        RECT 20.400 296.000 21.200 299.800 ;
        RECT 23.600 296.000 24.400 299.800 ;
        RECT 20.400 295.800 24.400 296.000 ;
        RECT 25.200 295.800 26.000 299.800 ;
        RECT 20.600 295.400 24.200 295.800 ;
        RECT 21.200 294.400 22.000 294.800 ;
        RECT 25.200 294.400 25.800 295.800 ;
        RECT 12.400 293.600 13.200 293.800 ;
        RECT 14.200 293.800 16.000 294.200 ;
        RECT 20.400 293.800 22.000 294.400 ;
        RECT 14.200 293.600 15.800 293.800 ;
        RECT 20.400 293.600 21.200 293.800 ;
        RECT 23.400 293.600 26.000 294.400 ;
        RECT 7.600 290.200 8.400 290.400 ;
        RECT 9.600 290.200 10.200 293.600 ;
        RECT 10.800 292.300 11.600 293.200 ;
        RECT 12.400 292.300 13.200 292.400 ;
        RECT 10.800 291.700 13.200 292.300 ;
        RECT 10.800 291.600 11.600 291.700 ;
        RECT 12.400 291.600 13.200 291.700 ;
        RECT 14.200 290.400 14.800 293.600 ;
        RECT 16.400 291.600 18.000 292.400 ;
        RECT 22.000 291.600 22.800 293.200 ;
        RECT 23.400 292.400 24.000 293.600 ;
        RECT 23.400 291.600 24.400 292.400 ;
        RECT 7.600 289.600 9.000 290.200 ;
        RECT 9.600 289.600 10.600 290.200 ;
        RECT 14.000 289.600 14.800 290.400 ;
        RECT 18.800 289.600 19.600 291.200 ;
        RECT 23.400 290.200 24.000 291.600 ;
        RECT 25.200 290.300 26.000 290.400 ;
        RECT 26.800 290.300 27.600 299.800 ;
        RECT 28.400 295.600 29.200 297.200 ;
        RECT 30.000 295.800 30.800 299.800 ;
        RECT 31.600 296.000 32.400 299.800 ;
        RECT 34.800 296.000 35.600 299.800 ;
        RECT 36.600 296.400 37.400 297.200 ;
        RECT 31.600 295.800 35.600 296.000 ;
        RECT 30.200 294.400 30.800 295.800 ;
        RECT 31.800 295.400 35.400 295.800 ;
        RECT 36.400 295.600 37.200 296.400 ;
        RECT 38.000 295.800 38.800 299.800 ;
        RECT 45.800 295.800 47.400 299.800 ;
        RECT 50.800 296.000 51.600 299.800 ;
        RECT 54.000 296.000 54.800 299.800 ;
        RECT 50.800 295.800 54.800 296.000 ;
        RECT 55.600 295.800 56.400 299.800 ;
        RECT 57.200 295.800 58.000 299.800 ;
        RECT 58.800 296.000 59.600 299.800 ;
        RECT 62.000 296.000 62.800 299.800 ;
        RECT 58.800 295.800 62.800 296.000 ;
        RECT 63.600 296.000 64.400 299.800 ;
        RECT 66.800 296.000 67.600 299.800 ;
        RECT 63.600 295.800 67.600 296.000 ;
        RECT 68.400 295.800 69.200 299.800 ;
        RECT 70.600 296.400 71.400 299.800 ;
        RECT 76.400 297.600 77.200 299.800 ;
        RECT 70.600 295.800 72.400 296.400 ;
        RECT 34.000 294.400 34.800 294.800 ;
        RECT 30.000 293.600 32.600 294.400 ;
        RECT 34.000 293.800 35.600 294.400 ;
        RECT 34.800 293.600 35.600 293.800 ;
        RECT 28.400 292.300 29.200 292.400 ;
        RECT 32.000 292.300 32.600 293.600 ;
        RECT 28.400 291.700 32.600 292.300 ;
        RECT 28.400 291.600 29.200 291.700 ;
        RECT 25.200 290.200 27.600 290.300 ;
        RECT 23.000 289.600 24.000 290.200 ;
        RECT 24.600 289.700 27.600 290.200 ;
        RECT 24.600 289.600 26.000 289.700 ;
        RECT 8.400 288.400 9.000 289.600 ;
        RECT 8.400 287.600 9.200 288.400 ;
        RECT 9.800 284.400 10.600 289.600 ;
        RECT 14.200 287.000 14.800 289.600 ;
        RECT 15.600 287.600 16.400 289.200 ;
        RECT 14.200 286.400 17.800 287.000 ;
        RECT 14.200 286.200 14.800 286.400 ;
        RECT 9.800 283.600 11.600 284.400 ;
        RECT 9.800 282.200 10.600 283.600 ;
        RECT 14.000 282.200 14.800 286.200 ;
        RECT 17.200 286.200 17.800 286.400 ;
        RECT 17.200 282.200 18.000 286.200 ;
        RECT 23.000 282.200 23.800 289.600 ;
        RECT 24.600 288.400 25.200 289.600 ;
        RECT 24.400 287.600 25.200 288.400 ;
        RECT 26.800 282.200 27.600 289.700 ;
        RECT 30.000 290.200 30.800 290.400 ;
        RECT 32.000 290.200 32.600 291.700 ;
        RECT 33.200 291.600 34.000 293.200 ;
        RECT 36.400 292.200 37.200 292.400 ;
        RECT 38.200 292.200 38.800 295.800 ;
        RECT 39.600 292.800 40.400 294.400 ;
        RECT 44.400 292.800 45.200 294.400 ;
        RECT 46.200 292.400 46.800 295.800 ;
        RECT 51.000 295.400 54.600 295.800 ;
        RECT 51.600 294.400 52.400 294.800 ;
        RECT 55.600 294.400 56.200 295.800 ;
        RECT 57.400 294.400 58.000 295.800 ;
        RECT 59.000 295.400 62.600 295.800 ;
        RECT 63.800 295.400 67.400 295.800 ;
        RECT 61.200 294.400 62.000 294.800 ;
        RECT 64.400 294.400 65.200 294.800 ;
        RECT 68.400 294.400 69.000 295.800 ;
        RECT 47.600 293.600 48.400 294.400 ;
        RECT 50.800 293.800 52.400 294.400 ;
        RECT 50.800 293.600 51.600 293.800 ;
        RECT 53.800 293.600 56.400 294.400 ;
        RECT 57.200 293.600 59.800 294.400 ;
        RECT 61.200 293.800 62.800 294.400 ;
        RECT 62.000 293.600 62.800 293.800 ;
        RECT 63.600 293.800 65.200 294.400 ;
        RECT 63.600 293.600 64.400 293.800 ;
        RECT 66.600 293.600 69.200 294.400 ;
        RECT 47.600 293.200 48.200 293.600 ;
        RECT 47.400 292.400 48.200 293.200 ;
        RECT 41.200 292.300 42.000 292.400 ;
        RECT 42.800 292.300 43.600 292.400 ;
        RECT 41.200 292.200 43.600 292.300 ;
        RECT 36.400 291.600 38.800 292.200 ;
        RECT 40.400 291.700 44.400 292.200 ;
        RECT 40.400 291.600 42.000 291.700 ;
        RECT 42.800 291.600 44.400 291.700 ;
        RECT 46.000 291.600 46.800 292.400 ;
        RECT 36.600 290.200 37.200 291.600 ;
        RECT 40.400 291.200 41.200 291.600 ;
        RECT 43.600 291.200 44.400 291.600 ;
        RECT 46.200 291.400 46.800 291.600 ;
        RECT 46.200 290.800 48.200 291.400 ;
        RECT 49.200 290.800 50.000 292.400 ;
        RECT 52.400 291.600 53.200 293.200 ;
        RECT 53.800 292.300 54.400 293.600 ;
        RECT 53.800 291.700 57.900 292.300 ;
        RECT 47.600 290.200 48.200 290.800 ;
        RECT 53.800 290.200 54.400 291.700 ;
        RECT 57.300 290.400 57.900 291.700 ;
        RECT 55.600 290.200 56.400 290.400 ;
        RECT 30.000 289.600 31.400 290.200 ;
        RECT 32.000 289.600 33.000 290.200 ;
        RECT 30.800 288.400 31.400 289.600 ;
        RECT 30.800 287.600 31.600 288.400 ;
        RECT 32.200 282.200 33.000 289.600 ;
        RECT 36.400 282.200 37.200 290.200 ;
        RECT 38.000 289.600 42.000 290.200 ;
        RECT 38.000 282.200 38.800 289.600 ;
        RECT 41.200 282.200 42.000 289.600 ;
        RECT 42.800 289.600 46.800 290.200 ;
        RECT 42.800 282.200 43.600 289.600 ;
        RECT 46.000 282.800 46.800 289.600 ;
        RECT 47.600 283.400 48.400 290.200 ;
        RECT 49.200 282.800 50.000 290.200 ;
        RECT 46.000 282.200 50.000 282.800 ;
        RECT 53.400 289.600 54.400 290.200 ;
        RECT 55.000 289.600 56.400 290.200 ;
        RECT 57.200 290.200 58.000 290.400 ;
        RECT 59.200 290.200 59.800 293.600 ;
        RECT 60.400 292.300 61.200 293.200 ;
        RECT 65.200 292.300 66.000 293.200 ;
        RECT 60.400 291.700 66.000 292.300 ;
        RECT 60.400 291.600 61.200 291.700 ;
        RECT 65.200 291.600 66.000 291.700 ;
        RECT 66.600 290.200 67.200 293.600 ;
        RECT 71.600 292.300 72.400 295.800 ;
        RECT 73.200 293.600 74.000 295.200 ;
        RECT 76.400 294.400 77.000 297.600 ;
        RECT 78.000 295.600 78.800 297.200 ;
        RECT 82.200 295.800 83.800 299.800 ;
        RECT 90.200 298.400 91.000 299.800 ;
        RECT 90.200 297.600 91.600 298.400 ;
        RECT 90.200 296.400 91.000 297.600 ;
        RECT 89.200 295.800 91.000 296.400 ;
        RECT 92.400 295.800 93.200 299.800 ;
        RECT 96.800 296.200 98.400 299.800 ;
        RECT 76.400 293.600 77.200 294.400 ;
        RECT 79.600 294.300 80.400 294.400 ;
        RECT 81.200 294.300 82.000 294.400 ;
        RECT 79.600 293.700 82.000 294.300 ;
        RECT 79.600 293.600 80.400 293.700 ;
        RECT 81.200 293.600 82.000 293.700 ;
        RECT 68.500 291.700 72.400 292.300 ;
        RECT 68.500 290.400 69.100 291.700 ;
        RECT 68.400 290.200 69.200 290.400 ;
        RECT 57.200 289.600 58.600 290.200 ;
        RECT 59.200 289.600 60.200 290.200 ;
        RECT 53.400 282.200 54.200 289.600 ;
        RECT 55.000 288.400 55.600 289.600 ;
        RECT 54.800 287.600 55.600 288.400 ;
        RECT 58.000 288.400 58.600 289.600 ;
        RECT 58.000 287.600 58.800 288.400 ;
        RECT 59.400 286.400 60.200 289.600 ;
        RECT 66.200 289.600 67.200 290.200 ;
        RECT 67.800 289.600 69.200 290.200 ;
        RECT 59.400 285.600 61.200 286.400 ;
        RECT 59.400 282.200 60.200 285.600 ;
        RECT 66.200 284.400 67.000 289.600 ;
        RECT 67.800 288.400 68.400 289.600 ;
        RECT 70.000 288.800 70.800 290.400 ;
        RECT 67.600 287.600 68.400 288.400 ;
        RECT 65.200 283.600 67.000 284.400 ;
        RECT 66.200 282.200 67.000 283.600 ;
        RECT 71.600 282.200 72.400 291.700 ;
        RECT 74.800 290.800 75.600 292.400 ;
        RECT 76.400 292.300 77.000 293.600 ;
        RECT 81.400 293.200 82.000 293.600 ;
        RECT 81.400 292.400 82.200 293.200 ;
        RECT 82.800 292.400 83.400 295.800 ;
        RECT 84.400 292.800 85.200 294.400 ;
        RECT 87.600 293.600 88.400 295.200 ;
        RECT 79.600 292.300 80.400 292.400 ;
        RECT 76.400 291.700 80.400 292.300 ;
        RECT 76.400 290.200 77.000 291.700 ;
        RECT 79.600 290.800 80.400 291.700 ;
        RECT 82.800 291.600 83.600 292.400 ;
        RECT 86.000 292.200 86.800 292.400 ;
        RECT 85.200 291.600 86.800 292.200 ;
        RECT 82.800 291.400 83.400 291.600 ;
        RECT 81.400 290.800 83.400 291.400 ;
        RECT 85.200 291.200 86.000 291.600 ;
        RECT 81.400 290.200 82.000 290.800 ;
        RECT 75.400 289.400 77.200 290.200 ;
        RECT 75.400 282.200 76.200 289.400 ;
        RECT 79.600 282.800 80.400 290.200 ;
        RECT 81.200 283.400 82.000 290.200 ;
        RECT 82.800 289.600 86.800 290.200 ;
        RECT 82.800 282.800 83.600 289.600 ;
        RECT 79.600 282.200 83.600 282.800 ;
        RECT 86.000 282.200 86.800 289.600 ;
        RECT 89.200 282.200 90.000 295.800 ;
        RECT 92.400 295.200 94.800 295.800 ;
        RECT 94.000 295.000 94.800 295.200 ;
        RECT 95.400 294.800 96.200 295.600 ;
        RECT 95.400 294.400 96.000 294.800 ;
        RECT 92.400 293.600 94.000 294.400 ;
        RECT 95.200 293.600 96.000 294.400 ;
        RECT 96.800 292.800 97.400 296.200 ;
        RECT 102.000 295.800 102.800 299.800 ;
        RECT 98.000 295.400 99.600 295.600 ;
        RECT 98.000 294.800 100.000 295.400 ;
        RECT 100.600 295.200 102.800 295.800 ;
        RECT 100.600 295.000 101.400 295.200 ;
        RECT 99.400 294.400 100.000 294.800 ;
        RECT 98.000 293.400 98.800 294.200 ;
        RECT 99.400 293.800 102.800 294.400 ;
        RECT 101.200 293.600 102.800 293.800 ;
        RECT 96.400 292.400 97.400 292.800 ;
        RECT 90.800 292.300 91.600 292.400 ;
        RECT 95.600 292.300 97.400 292.400 ;
        RECT 90.800 292.200 97.400 292.300 ;
        RECT 98.200 292.800 98.800 293.400 ;
        RECT 98.200 292.200 100.800 292.800 ;
        RECT 90.800 291.700 97.000 292.200 ;
        RECT 100.000 292.000 100.800 292.200 ;
        RECT 103.600 292.300 104.400 299.800 ;
        RECT 106.800 296.000 107.600 299.800 ;
        RECT 110.000 296.000 110.800 299.800 ;
        RECT 106.800 295.800 110.800 296.000 ;
        RECT 111.600 295.800 112.400 299.800 ;
        RECT 107.000 295.400 110.600 295.800 ;
        RECT 105.200 293.600 106.000 295.200 ;
        RECT 107.600 294.400 108.400 294.800 ;
        RECT 111.600 294.400 112.200 295.800 ;
        RECT 113.200 295.600 114.000 297.200 ;
        RECT 114.800 296.300 115.600 299.800 ;
        RECT 116.600 296.400 117.400 297.200 ;
        RECT 116.400 296.300 117.200 296.400 ;
        RECT 114.800 295.700 117.200 296.300 ;
        RECT 118.000 295.800 118.800 299.800 ;
        RECT 122.800 295.800 123.600 299.800 ;
        RECT 124.400 296.000 125.200 299.800 ;
        RECT 127.600 296.000 128.400 299.800 ;
        RECT 131.800 296.400 132.600 299.800 ;
        RECT 136.600 296.400 137.400 299.800 ;
        RECT 124.400 295.800 128.400 296.000 ;
        RECT 130.800 295.800 132.600 296.400 ;
        RECT 135.600 295.800 137.400 296.400 ;
        RECT 144.200 296.400 145.000 299.800 ;
        RECT 150.000 297.600 150.800 299.800 ;
        RECT 144.200 295.800 146.000 296.400 ;
        RECT 106.800 293.800 108.400 294.400 ;
        RECT 106.800 293.600 107.600 293.800 ;
        RECT 109.800 293.600 112.400 294.400 ;
        RECT 106.800 292.300 107.600 292.400 ;
        RECT 90.800 291.600 91.600 291.700 ;
        RECT 95.600 291.600 97.000 291.700 ;
        RECT 103.600 291.700 107.600 292.300 ;
        RECT 90.800 288.800 91.600 290.400 ;
        RECT 96.400 290.200 97.000 291.600 ;
        RECT 97.800 291.400 98.600 291.600 ;
        RECT 97.800 290.800 101.200 291.400 ;
        RECT 100.600 290.200 101.200 290.800 ;
        RECT 92.400 289.600 94.800 290.200 ;
        RECT 96.400 289.600 98.400 290.200 ;
        RECT 92.400 282.200 93.200 289.600 ;
        RECT 94.000 289.400 94.800 289.600 ;
        RECT 96.800 282.200 98.400 289.600 ;
        RECT 100.600 289.600 102.800 290.200 ;
        RECT 100.600 289.400 101.400 289.600 ;
        RECT 102.000 282.200 102.800 289.600 ;
        RECT 103.600 282.200 104.400 291.700 ;
        RECT 106.800 291.600 107.600 291.700 ;
        RECT 108.400 291.600 109.200 293.200 ;
        RECT 109.800 290.200 110.400 293.600 ;
        RECT 111.600 290.300 112.400 290.400 ;
        RECT 113.200 290.300 114.000 290.400 ;
        RECT 111.600 290.200 114.000 290.300 ;
        RECT 109.400 289.600 110.400 290.200 ;
        RECT 111.000 289.700 114.000 290.200 ;
        RECT 111.000 289.600 112.400 289.700 ;
        RECT 113.200 289.600 114.000 289.700 ;
        RECT 109.400 286.400 110.200 289.600 ;
        RECT 111.000 288.400 111.600 289.600 ;
        RECT 110.800 287.600 111.600 288.400 ;
        RECT 108.400 285.600 110.200 286.400 ;
        RECT 109.400 282.200 110.200 285.600 ;
        RECT 114.800 282.200 115.600 295.700 ;
        RECT 116.400 295.600 117.200 295.700 ;
        RECT 116.400 292.200 117.200 292.400 ;
        RECT 118.200 292.200 118.800 295.800 ;
        RECT 123.000 294.400 123.600 295.800 ;
        RECT 124.600 295.400 128.200 295.800 ;
        RECT 126.800 294.400 127.600 294.800 ;
        RECT 119.600 292.800 120.400 294.400 ;
        RECT 122.800 293.600 125.400 294.400 ;
        RECT 126.800 293.800 128.400 294.400 ;
        RECT 127.600 293.600 128.400 293.800 ;
        RECT 129.200 293.600 130.000 295.200 ;
        RECT 130.800 294.300 131.600 295.800 ;
        RECT 134.000 294.300 134.800 295.200 ;
        RECT 130.800 293.700 134.800 294.300 ;
        RECT 121.200 292.200 122.000 292.400 ;
        RECT 116.400 291.600 118.800 292.200 ;
        RECT 120.400 291.600 122.000 292.200 ;
        RECT 116.600 290.200 117.200 291.600 ;
        RECT 120.400 291.200 121.200 291.600 ;
        RECT 122.800 290.200 123.600 290.400 ;
        RECT 124.800 290.200 125.400 293.600 ;
        RECT 126.000 291.600 126.800 293.200 ;
        RECT 116.400 282.200 117.200 290.200 ;
        RECT 118.000 289.600 122.000 290.200 ;
        RECT 122.800 289.600 124.200 290.200 ;
        RECT 124.800 289.600 125.800 290.200 ;
        RECT 118.000 282.200 118.800 289.600 ;
        RECT 121.200 282.200 122.000 289.600 ;
        RECT 123.600 288.400 124.200 289.600 ;
        RECT 123.600 287.600 124.400 288.400 ;
        RECT 125.000 282.200 125.800 289.600 ;
        RECT 130.800 282.200 131.600 293.700 ;
        RECT 134.000 293.600 134.800 293.700 ;
        RECT 132.400 288.800 133.200 290.400 ;
        RECT 135.600 282.200 136.400 295.800 ;
        RECT 137.200 292.300 138.000 292.400 ;
        RECT 145.200 292.300 146.000 295.800 ;
        RECT 146.800 293.600 147.600 295.200 ;
        RECT 150.000 294.400 150.600 297.600 ;
        RECT 151.600 295.600 152.400 297.200 ;
        RECT 156.400 295.800 157.200 299.800 ;
        RECT 157.800 296.400 158.600 297.200 ;
        RECT 150.000 293.600 150.800 294.400 ;
        RECT 153.200 294.300 154.000 294.400 ;
        RECT 154.800 294.300 155.600 294.400 ;
        RECT 153.200 293.700 155.600 294.300 ;
        RECT 153.200 293.600 154.000 293.700 ;
        RECT 137.200 291.700 146.000 292.300 ;
        RECT 137.200 291.600 138.000 291.700 ;
        RECT 137.300 290.400 137.900 291.600 ;
        RECT 137.200 288.800 138.000 290.400 ;
        RECT 143.600 288.800 144.400 290.400 ;
        RECT 145.200 282.200 146.000 291.700 ;
        RECT 148.400 290.800 149.200 292.400 ;
        RECT 150.000 290.200 150.600 293.600 ;
        RECT 154.800 292.800 155.600 293.700 ;
        RECT 153.200 292.200 154.000 292.400 ;
        RECT 156.400 292.200 157.000 295.800 ;
        RECT 158.000 295.600 158.800 296.400 ;
        RECT 159.600 296.000 160.400 299.800 ;
        RECT 162.800 296.000 163.600 299.800 ;
        RECT 159.600 295.800 163.600 296.000 ;
        RECT 164.400 295.800 165.200 299.800 ;
        RECT 159.800 295.400 163.400 295.800 ;
        RECT 160.400 294.400 161.200 294.800 ;
        RECT 164.400 294.400 165.000 295.800 ;
        RECT 159.600 293.800 161.200 294.400 ;
        RECT 159.600 293.600 160.400 293.800 ;
        RECT 162.600 293.600 165.200 294.400 ;
        RECT 158.000 292.200 158.800 292.400 ;
        RECT 153.200 291.600 154.800 292.200 ;
        RECT 156.400 291.600 158.800 292.200 ;
        RECT 161.200 291.600 162.000 293.200 ;
        RECT 154.000 291.200 154.800 291.600 ;
        RECT 158.000 290.200 158.600 291.600 ;
        RECT 162.600 290.400 163.200 293.600 ;
        RECT 149.000 289.400 150.800 290.200 ;
        RECT 153.200 289.600 157.200 290.200 ;
        RECT 149.000 282.200 149.800 289.400 ;
        RECT 153.200 282.200 154.000 289.600 ;
        RECT 156.400 282.200 157.200 289.600 ;
        RECT 158.000 282.200 158.800 290.200 ;
        RECT 161.200 289.600 163.200 290.400 ;
        RECT 164.400 290.300 165.200 290.400 ;
        RECT 166.000 290.300 166.800 299.800 ;
        RECT 167.600 296.300 168.400 297.200 ;
        RECT 169.400 296.400 170.200 297.200 ;
        RECT 169.200 296.300 170.000 296.400 ;
        RECT 167.600 295.700 170.000 296.300 ;
        RECT 170.800 295.800 171.600 299.800 ;
        RECT 167.600 295.600 168.400 295.700 ;
        RECT 169.200 295.600 170.000 295.700 ;
        RECT 169.200 292.200 170.000 292.400 ;
        RECT 171.000 292.200 171.600 295.800 ;
        RECT 177.200 297.800 178.000 299.800 ;
        RECT 177.200 294.400 177.800 297.800 ;
        RECT 178.800 295.600 179.600 297.200 ;
        RECT 180.400 296.000 181.200 299.800 ;
        RECT 183.600 296.000 184.400 299.800 ;
        RECT 180.400 295.800 184.400 296.000 ;
        RECT 185.200 295.800 186.000 299.800 ;
        RECT 186.800 295.800 187.600 299.800 ;
        RECT 191.200 296.200 192.800 299.800 ;
        RECT 172.400 294.300 173.200 294.400 ;
        RECT 175.600 294.300 176.400 294.400 ;
        RECT 172.400 293.700 176.400 294.300 ;
        RECT 172.400 292.800 173.200 293.700 ;
        RECT 175.600 293.600 176.400 293.700 ;
        RECT 177.200 293.600 178.000 294.400 ;
        RECT 178.900 294.300 179.500 295.600 ;
        RECT 180.600 295.400 184.200 295.800 ;
        RECT 181.200 294.400 182.000 294.800 ;
        RECT 185.200 294.400 185.800 295.800 ;
        RECT 186.800 295.200 189.000 295.800 ;
        RECT 190.000 295.400 191.600 295.600 ;
        RECT 188.200 295.000 189.000 295.200 ;
        RECT 189.600 294.800 191.600 295.400 ;
        RECT 189.600 294.400 190.200 294.800 ;
        RECT 180.400 294.300 182.000 294.400 ;
        RECT 178.900 293.800 182.000 294.300 ;
        RECT 178.900 293.700 181.200 293.800 ;
        RECT 180.400 293.600 181.200 293.700 ;
        RECT 183.400 293.600 186.000 294.400 ;
        RECT 186.800 293.800 190.200 294.400 ;
        RECT 186.800 293.600 188.400 293.800 ;
        RECT 174.000 292.200 174.800 292.400 ;
        RECT 169.200 291.600 171.600 292.200 ;
        RECT 173.200 291.600 174.800 292.200 ;
        RECT 164.400 290.200 166.800 290.300 ;
        RECT 169.400 290.200 170.000 291.600 ;
        RECT 173.200 291.200 174.000 291.600 ;
        RECT 175.600 290.800 176.400 292.400 ;
        RECT 177.200 290.200 177.800 293.600 ;
        RECT 182.000 291.600 182.800 293.200 ;
        RECT 183.400 290.200 184.000 293.600 ;
        RECT 185.200 292.300 186.000 292.400 ;
        RECT 186.900 292.300 187.500 293.600 ;
        RECT 190.800 293.400 191.600 294.200 ;
        RECT 190.800 292.800 191.400 293.400 ;
        RECT 185.200 291.700 187.500 292.300 ;
        RECT 188.800 292.200 191.400 292.800 ;
        RECT 192.200 292.800 192.800 296.200 ;
        RECT 196.400 295.800 197.200 299.800 ;
        RECT 193.400 294.800 194.200 295.600 ;
        RECT 194.800 295.200 197.200 295.800 ;
        RECT 198.000 295.400 198.800 299.800 ;
        RECT 202.200 298.400 203.400 299.800 ;
        RECT 202.200 297.800 203.600 298.400 ;
        RECT 206.800 297.800 207.600 299.800 ;
        RECT 211.200 298.400 212.000 299.800 ;
        RECT 211.200 297.800 213.200 298.400 ;
        RECT 202.800 297.000 203.600 297.800 ;
        RECT 207.000 297.200 207.600 297.800 ;
        RECT 207.000 296.600 209.800 297.200 ;
        RECT 209.000 296.400 209.800 296.600 ;
        RECT 210.800 295.600 211.600 297.200 ;
        RECT 212.400 297.000 213.200 297.800 ;
        RECT 201.000 295.400 201.800 295.600 ;
        RECT 194.800 295.000 195.600 295.200 ;
        RECT 193.600 294.400 194.200 294.800 ;
        RECT 198.000 294.800 201.800 295.400 ;
        RECT 193.600 293.600 194.400 294.400 ;
        RECT 195.600 294.300 197.200 294.400 ;
        RECT 198.000 294.300 198.800 294.800 ;
        RECT 195.600 293.700 198.800 294.300 ;
        RECT 205.000 294.200 205.800 294.400 ;
        RECT 210.800 294.200 211.400 295.600 ;
        RECT 215.600 295.000 216.400 299.800 ;
        RECT 214.000 294.200 215.600 294.400 ;
        RECT 195.600 293.600 197.200 293.700 ;
        RECT 192.200 292.400 193.200 292.800 ;
        RECT 192.200 292.200 194.000 292.400 ;
        RECT 188.800 292.000 189.600 292.200 ;
        RECT 185.200 291.600 186.000 291.700 ;
        RECT 192.600 291.600 194.000 292.200 ;
        RECT 191.000 291.400 191.800 291.600 ;
        RECT 188.400 290.800 191.800 291.400 ;
        RECT 185.200 290.200 186.000 290.400 ;
        RECT 188.400 290.200 189.000 290.800 ;
        RECT 192.600 290.200 193.200 291.600 ;
        RECT 198.000 291.400 198.800 293.700 ;
        RECT 204.600 293.600 215.600 294.200 ;
        RECT 202.800 292.800 203.600 293.000 ;
        RECT 199.800 292.200 203.600 292.800 ;
        RECT 204.600 292.400 205.200 293.600 ;
        RECT 211.800 293.400 212.600 293.600 ;
        RECT 210.800 292.400 211.600 292.600 ;
        RECT 213.400 292.400 214.200 292.600 ;
        RECT 199.800 292.000 200.600 292.200 ;
        RECT 204.400 291.600 205.200 292.400 ;
        RECT 209.200 291.800 214.200 292.400 ;
        RECT 217.200 292.400 218.000 299.800 ;
        RECT 220.400 295.200 221.200 299.800 ;
        RECT 219.000 294.600 221.200 295.200 ;
        RECT 222.000 295.200 222.800 299.800 ;
        RECT 222.000 294.600 224.200 295.200 ;
        RECT 209.200 291.600 210.000 291.800 ;
        RECT 201.400 291.400 202.200 291.600 ;
        RECT 198.000 290.800 202.200 291.400 ;
        RECT 163.800 289.700 166.800 290.200 ;
        RECT 163.800 289.600 165.200 289.700 ;
        RECT 162.200 282.200 163.000 289.600 ;
        RECT 163.800 288.400 164.400 289.600 ;
        RECT 163.600 287.600 164.400 288.400 ;
        RECT 166.000 282.200 166.800 289.700 ;
        RECT 169.200 282.200 170.000 290.200 ;
        RECT 170.800 289.600 174.800 290.200 ;
        RECT 170.800 282.200 171.600 289.600 ;
        RECT 174.000 282.200 174.800 289.600 ;
        RECT 176.200 289.400 178.000 290.200 ;
        RECT 183.000 289.600 184.000 290.200 ;
        RECT 184.600 289.600 186.000 290.200 ;
        RECT 186.800 289.600 189.000 290.200 ;
        RECT 176.200 284.400 177.000 289.400 ;
        RECT 175.600 283.600 177.000 284.400 ;
        RECT 176.200 282.200 177.000 283.600 ;
        RECT 183.000 282.200 183.800 289.600 ;
        RECT 184.600 288.400 185.200 289.600 ;
        RECT 184.400 287.600 185.200 288.400 ;
        RECT 186.800 282.200 187.600 289.600 ;
        RECT 188.200 289.400 189.000 289.600 ;
        RECT 191.200 289.600 193.200 290.200 ;
        RECT 194.800 289.600 197.200 290.200 ;
        RECT 191.200 288.400 192.800 289.600 ;
        RECT 194.800 289.400 195.600 289.600 ;
        RECT 190.000 287.600 192.800 288.400 ;
        RECT 191.200 282.200 192.800 287.600 ;
        RECT 196.400 282.200 197.200 289.600 ;
        RECT 198.000 282.200 198.800 290.800 ;
        RECT 204.600 290.400 205.200 291.600 ;
        RECT 210.800 291.000 216.400 291.200 ;
        RECT 210.600 290.800 216.400 291.000 ;
        RECT 202.800 289.800 205.200 290.400 ;
        RECT 206.600 290.600 216.400 290.800 ;
        RECT 206.600 290.200 211.400 290.600 ;
        RECT 202.800 288.800 203.400 289.800 ;
        RECT 202.000 288.000 203.400 288.800 ;
        RECT 205.000 289.000 205.800 289.200 ;
        RECT 206.600 289.000 207.200 290.200 ;
        RECT 205.000 288.400 207.200 289.000 ;
        RECT 207.800 289.000 213.200 289.600 ;
        RECT 207.800 288.800 208.600 289.000 ;
        RECT 212.400 288.800 213.200 289.000 ;
        RECT 206.200 287.400 207.000 287.600 ;
        RECT 209.000 287.400 209.800 287.600 ;
        RECT 202.800 286.200 203.600 287.000 ;
        RECT 206.200 286.800 209.800 287.400 ;
        RECT 207.000 286.200 207.600 286.800 ;
        RECT 212.400 286.200 213.200 287.000 ;
        RECT 202.200 282.200 203.400 286.200 ;
        RECT 206.800 282.200 207.600 286.200 ;
        RECT 211.200 285.600 213.200 286.200 ;
        RECT 211.200 282.200 212.000 285.600 ;
        RECT 215.600 282.200 216.400 290.600 ;
        RECT 217.200 290.200 217.800 292.400 ;
        RECT 219.000 291.600 219.600 294.600 ;
        RECT 218.400 290.800 219.600 291.600 ;
        RECT 219.000 290.200 219.600 290.800 ;
        RECT 223.600 291.600 224.200 294.600 ;
        RECT 225.200 292.400 226.000 299.800 ;
        RECT 226.800 295.000 227.600 299.800 ;
        RECT 231.200 298.400 232.000 299.800 ;
        RECT 230.000 297.800 232.000 298.400 ;
        RECT 235.600 297.800 236.400 299.800 ;
        RECT 239.800 298.400 241.000 299.800 ;
        RECT 239.600 297.800 241.000 298.400 ;
        RECT 230.000 297.000 230.800 297.800 ;
        RECT 235.600 297.200 236.200 297.800 ;
        RECT 231.600 296.400 232.400 297.200 ;
        RECT 233.400 296.600 236.200 297.200 ;
        RECT 239.600 297.000 240.400 297.800 ;
        RECT 233.400 296.400 234.200 296.600 ;
        RECT 231.800 294.400 232.400 296.400 ;
        RECT 241.400 295.400 242.200 295.600 ;
        RECT 244.400 295.400 245.200 299.800 ;
        RECT 241.400 294.800 245.200 295.400 ;
        RECT 246.000 295.800 246.800 299.800 ;
        RECT 250.400 296.200 252.000 299.800 ;
        RECT 246.000 295.200 248.400 295.800 ;
        RECT 247.600 295.000 248.400 295.200 ;
        RECT 227.600 294.200 229.200 294.400 ;
        RECT 231.600 294.200 232.400 294.400 ;
        RECT 237.400 294.200 238.200 294.400 ;
        RECT 227.600 293.600 238.600 294.200 ;
        RECT 230.600 293.400 231.400 293.600 ;
        RECT 223.600 290.800 224.800 291.600 ;
        RECT 223.600 290.200 224.200 290.800 ;
        RECT 225.400 290.200 226.000 292.400 ;
        RECT 217.200 282.200 218.000 290.200 ;
        RECT 219.000 289.600 221.200 290.200 ;
        RECT 220.400 282.200 221.200 289.600 ;
        RECT 222.000 289.600 224.200 290.200 ;
        RECT 222.000 282.200 222.800 289.600 ;
        RECT 225.200 282.200 226.000 290.200 ;
        RECT 226.800 291.000 232.400 291.200 ;
        RECT 226.800 290.800 232.600 291.000 ;
        RECT 226.800 290.600 236.600 290.800 ;
        RECT 226.800 282.200 227.600 290.600 ;
        RECT 231.800 290.200 236.600 290.600 ;
        RECT 230.000 289.000 235.400 289.600 ;
        RECT 230.000 288.800 230.800 289.000 ;
        RECT 234.600 288.800 235.400 289.000 ;
        RECT 236.000 289.000 236.600 290.200 ;
        RECT 238.000 290.400 238.600 293.600 ;
        RECT 239.600 292.800 240.400 293.000 ;
        RECT 239.600 292.200 243.400 292.800 ;
        RECT 242.600 292.000 243.400 292.200 ;
        RECT 241.000 291.400 241.800 291.600 ;
        RECT 244.400 291.400 245.200 294.800 ;
        RECT 249.000 294.800 249.800 295.600 ;
        RECT 249.000 294.400 249.600 294.800 ;
        RECT 246.000 293.600 247.600 294.400 ;
        RECT 248.800 293.600 249.600 294.400 ;
        RECT 250.400 294.200 251.000 296.200 ;
        RECT 255.600 295.800 256.400 299.800 ;
        RECT 251.600 294.800 253.200 295.600 ;
        RECT 253.800 295.200 256.400 295.800 ;
        RECT 257.200 295.400 258.000 299.800 ;
        RECT 261.400 298.400 262.600 299.800 ;
        RECT 261.400 297.800 262.800 298.400 ;
        RECT 266.000 297.800 266.800 299.800 ;
        RECT 270.400 298.400 271.200 299.800 ;
        RECT 270.400 297.800 272.400 298.400 ;
        RECT 262.000 297.000 262.800 297.800 ;
        RECT 266.200 297.200 266.800 297.800 ;
        RECT 266.200 296.600 269.000 297.200 ;
        RECT 268.200 296.400 269.000 296.600 ;
        RECT 270.000 296.400 270.800 297.200 ;
        RECT 271.600 297.000 272.400 297.800 ;
        RECT 260.200 295.400 261.000 295.600 ;
        RECT 253.800 295.000 254.600 295.200 ;
        RECT 257.200 294.800 261.000 295.400 ;
        RECT 254.800 294.200 256.400 294.400 ;
        RECT 250.400 293.600 251.400 294.200 ;
        RECT 254.200 294.000 256.400 294.200 ;
        RECT 250.800 292.400 251.400 293.600 ;
        RECT 252.000 293.600 256.400 294.000 ;
        RECT 252.000 293.400 254.800 293.600 ;
        RECT 252.000 293.200 252.800 293.400 ;
        RECT 246.000 292.300 246.800 292.400 ;
        RECT 250.800 292.300 251.600 292.400 ;
        RECT 246.000 291.700 251.600 292.300 ;
        RECT 253.400 292.200 254.200 292.400 ;
        RECT 246.000 291.600 246.800 291.700 ;
        RECT 250.800 291.600 251.600 291.700 ;
        RECT 252.600 291.600 254.200 292.200 ;
        RECT 241.000 290.800 245.200 291.400 ;
        RECT 238.000 289.800 240.400 290.400 ;
        RECT 237.400 289.000 238.200 289.200 ;
        RECT 236.000 288.400 238.200 289.000 ;
        RECT 239.800 288.800 240.400 289.800 ;
        RECT 239.800 288.000 241.200 288.800 ;
        RECT 233.400 287.400 234.200 287.600 ;
        RECT 236.200 287.400 237.000 287.600 ;
        RECT 230.000 286.200 230.800 287.000 ;
        RECT 233.400 286.800 237.000 287.400 ;
        RECT 235.600 286.200 236.200 286.800 ;
        RECT 239.600 286.200 240.400 287.000 ;
        RECT 230.000 285.600 232.000 286.200 ;
        RECT 231.200 282.200 232.000 285.600 ;
        RECT 235.600 282.200 236.400 286.200 ;
        RECT 239.800 282.200 241.000 286.200 ;
        RECT 244.400 282.200 245.200 290.800 ;
        RECT 250.800 290.200 251.400 291.600 ;
        RECT 252.600 291.400 253.400 291.600 ;
        RECT 257.200 291.400 258.000 294.800 ;
        RECT 264.200 294.200 265.000 294.400 ;
        RECT 270.000 294.200 270.600 296.400 ;
        RECT 274.800 295.000 275.600 299.800 ;
        RECT 276.400 295.400 277.200 299.800 ;
        RECT 280.600 298.400 281.800 299.800 ;
        RECT 280.600 297.800 282.000 298.400 ;
        RECT 285.200 297.800 286.000 299.800 ;
        RECT 289.600 298.400 290.400 299.800 ;
        RECT 289.600 297.800 291.600 298.400 ;
        RECT 281.200 297.000 282.000 297.800 ;
        RECT 285.400 297.200 286.000 297.800 ;
        RECT 285.400 296.600 288.200 297.200 ;
        RECT 287.400 296.400 288.200 296.600 ;
        RECT 289.200 296.400 290.000 297.200 ;
        RECT 290.800 297.000 291.600 297.800 ;
        RECT 279.400 295.400 280.200 295.600 ;
        RECT 276.400 294.800 280.200 295.400 ;
        RECT 273.200 294.200 274.800 294.400 ;
        RECT 263.800 293.600 274.800 294.200 ;
        RECT 262.000 292.800 262.800 293.000 ;
        RECT 259.000 292.200 262.800 292.800 ;
        RECT 263.800 292.400 264.400 293.600 ;
        RECT 271.000 293.400 271.800 293.600 ;
        RECT 270.000 292.400 270.800 292.600 ;
        RECT 272.600 292.400 273.400 292.600 ;
        RECT 259.000 292.000 259.800 292.200 ;
        RECT 263.600 291.600 264.400 292.400 ;
        RECT 268.400 291.800 273.400 292.400 ;
        RECT 268.400 291.600 269.200 291.800 ;
        RECT 260.600 291.400 261.400 291.600 ;
        RECT 257.200 290.800 261.400 291.400 ;
        RECT 246.000 289.600 248.400 290.200 ;
        RECT 246.000 282.200 246.800 289.600 ;
        RECT 247.600 289.400 248.400 289.600 ;
        RECT 250.400 282.200 252.000 290.200 ;
        RECT 253.800 289.600 256.400 290.200 ;
        RECT 253.800 289.400 254.600 289.600 ;
        RECT 255.600 282.200 256.400 289.600 ;
        RECT 257.200 282.200 258.000 290.800 ;
        RECT 263.800 290.400 264.400 291.600 ;
        RECT 276.400 291.400 277.200 294.800 ;
        RECT 283.400 294.200 284.200 294.400 ;
        RECT 289.200 294.200 289.800 296.400 ;
        RECT 294.000 295.000 294.800 299.800 ;
        RECT 303.000 296.400 303.800 299.800 ;
        RECT 302.000 295.800 303.800 296.400 ;
        RECT 305.200 295.800 306.000 299.800 ;
        RECT 309.600 296.200 311.200 299.800 ;
        RECT 292.400 294.200 294.000 294.400 ;
        RECT 283.000 293.600 294.000 294.200 ;
        RECT 300.400 293.600 301.200 295.200 ;
        RECT 281.200 292.800 282.000 293.000 ;
        RECT 278.200 292.200 282.000 292.800 ;
        RECT 283.000 292.400 283.600 293.600 ;
        RECT 290.200 293.400 291.000 293.600 ;
        RECT 289.200 292.400 290.000 292.600 ;
        RECT 291.800 292.400 292.600 292.600 ;
        RECT 278.200 292.000 279.000 292.200 ;
        RECT 282.800 291.600 283.600 292.400 ;
        RECT 287.600 291.800 292.600 292.400 ;
        RECT 287.600 291.600 288.400 291.800 ;
        RECT 279.800 291.400 280.600 291.600 ;
        RECT 270.000 291.000 275.600 291.200 ;
        RECT 269.800 290.800 275.600 291.000 ;
        RECT 262.000 289.800 264.400 290.400 ;
        RECT 265.800 290.600 275.600 290.800 ;
        RECT 265.800 290.200 270.600 290.600 ;
        RECT 262.000 288.800 262.600 289.800 ;
        RECT 261.200 288.000 262.600 288.800 ;
        RECT 264.200 289.000 265.000 289.200 ;
        RECT 265.800 289.000 266.400 290.200 ;
        RECT 264.200 288.400 266.400 289.000 ;
        RECT 267.000 289.000 272.400 289.600 ;
        RECT 267.000 288.800 267.800 289.000 ;
        RECT 271.600 288.800 272.400 289.000 ;
        RECT 265.400 287.400 266.200 287.600 ;
        RECT 268.200 287.400 269.000 287.600 ;
        RECT 262.000 286.200 262.800 287.000 ;
        RECT 265.400 286.800 269.000 287.400 ;
        RECT 266.200 286.200 266.800 286.800 ;
        RECT 271.600 286.200 272.400 287.000 ;
        RECT 261.400 282.200 262.600 286.200 ;
        RECT 266.000 282.200 266.800 286.200 ;
        RECT 270.400 285.600 272.400 286.200 ;
        RECT 270.400 282.200 271.200 285.600 ;
        RECT 274.800 282.200 275.600 290.600 ;
        RECT 276.400 290.800 280.600 291.400 ;
        RECT 276.400 282.200 277.200 290.800 ;
        RECT 283.000 290.400 283.600 291.600 ;
        RECT 289.200 291.000 294.800 291.200 ;
        RECT 289.000 290.800 294.800 291.000 ;
        RECT 281.200 289.800 283.600 290.400 ;
        RECT 285.000 290.600 294.800 290.800 ;
        RECT 285.000 290.200 289.800 290.600 ;
        RECT 281.200 288.800 281.800 289.800 ;
        RECT 280.400 288.000 281.800 288.800 ;
        RECT 283.400 289.000 284.200 289.200 ;
        RECT 285.000 289.000 285.600 290.200 ;
        RECT 283.400 288.400 285.600 289.000 ;
        RECT 286.200 289.000 291.600 289.600 ;
        RECT 286.200 288.800 287.000 289.000 ;
        RECT 290.800 288.800 291.600 289.000 ;
        RECT 284.600 287.400 285.400 287.600 ;
        RECT 287.400 287.400 288.200 287.600 ;
        RECT 281.200 286.200 282.000 287.000 ;
        RECT 284.600 286.800 288.200 287.400 ;
        RECT 285.400 286.200 286.000 286.800 ;
        RECT 290.800 286.200 291.600 287.000 ;
        RECT 280.600 282.200 281.800 286.200 ;
        RECT 285.200 282.200 286.000 286.200 ;
        RECT 289.600 285.600 291.600 286.200 ;
        RECT 289.600 282.200 290.400 285.600 ;
        RECT 294.000 282.200 294.800 290.600 ;
        RECT 302.000 282.200 302.800 295.800 ;
        RECT 305.200 295.200 307.600 295.800 ;
        RECT 306.800 295.000 307.600 295.200 ;
        RECT 308.200 294.800 309.000 295.600 ;
        RECT 308.200 294.400 308.800 294.800 ;
        RECT 305.200 293.600 306.800 294.400 ;
        RECT 308.000 293.600 308.800 294.400 ;
        RECT 309.600 292.800 310.200 296.200 ;
        RECT 314.800 295.800 315.600 299.800 ;
        RECT 316.400 295.800 317.200 299.800 ;
        RECT 318.000 296.000 318.800 299.800 ;
        RECT 321.200 296.000 322.000 299.800 ;
        RECT 318.000 295.800 322.000 296.000 ;
        RECT 322.800 295.800 323.600 299.800 ;
        RECT 326.000 297.800 326.800 299.800 ;
        RECT 310.800 295.400 312.400 295.600 ;
        RECT 310.800 294.800 312.800 295.400 ;
        RECT 313.400 295.200 315.600 295.800 ;
        RECT 313.400 295.000 314.200 295.200 ;
        RECT 312.200 294.400 312.800 294.800 ;
        RECT 316.600 294.400 317.200 295.800 ;
        RECT 318.200 295.400 321.800 295.800 ;
        RECT 320.400 294.400 321.200 294.800 ;
        RECT 312.200 294.300 315.600 294.400 ;
        RECT 316.400 294.300 319.000 294.400 ;
        RECT 310.800 293.400 311.600 294.200 ;
        RECT 312.200 293.800 319.000 294.300 ;
        RECT 320.400 293.800 322.000 294.400 ;
        RECT 314.000 293.700 319.000 293.800 ;
        RECT 314.000 293.600 315.600 293.700 ;
        RECT 316.400 293.600 319.000 293.700 ;
        RECT 321.200 293.600 322.000 293.800 ;
        RECT 309.200 292.400 310.200 292.800 ;
        RECT 303.600 292.300 304.400 292.400 ;
        RECT 308.400 292.300 310.200 292.400 ;
        RECT 303.600 292.200 310.200 292.300 ;
        RECT 311.000 292.800 311.600 293.400 ;
        RECT 311.000 292.200 313.600 292.800 ;
        RECT 303.600 291.700 309.800 292.200 ;
        RECT 312.800 292.000 313.600 292.200 ;
        RECT 303.600 291.600 304.400 291.700 ;
        RECT 308.400 291.600 309.800 291.700 ;
        RECT 303.600 288.800 304.400 290.400 ;
        RECT 309.200 290.200 309.800 291.600 ;
        RECT 310.600 291.400 311.400 291.600 ;
        RECT 310.600 290.800 314.000 291.400 ;
        RECT 313.400 290.200 314.000 290.800 ;
        RECT 316.400 290.200 317.200 290.400 ;
        RECT 318.400 290.200 319.000 293.600 ;
        RECT 319.600 292.300 320.400 293.200 ;
        RECT 322.800 292.400 323.400 295.800 ;
        RECT 326.000 295.600 326.600 297.800 ;
        RECT 327.600 295.600 328.400 297.200 ;
        RECT 324.200 295.000 326.600 295.600 ;
        RECT 329.200 295.400 330.000 299.800 ;
        RECT 333.400 298.400 334.600 299.800 ;
        RECT 333.400 297.800 334.800 298.400 ;
        RECT 338.000 297.800 338.800 299.800 ;
        RECT 342.400 298.400 343.200 299.800 ;
        RECT 342.400 297.800 344.400 298.400 ;
        RECT 334.000 297.000 334.800 297.800 ;
        RECT 338.200 297.200 338.800 297.800 ;
        RECT 338.200 296.600 341.000 297.200 ;
        RECT 340.200 296.400 341.000 296.600 ;
        RECT 342.000 296.400 342.800 297.200 ;
        RECT 343.600 297.000 344.400 297.800 ;
        RECT 332.200 295.400 333.000 295.600 ;
        RECT 322.800 292.300 323.600 292.400 ;
        RECT 319.600 291.700 323.600 292.300 ;
        RECT 319.600 291.600 320.400 291.700 ;
        RECT 322.800 291.600 323.600 291.700 ;
        RECT 324.200 292.000 324.800 295.000 ;
        RECT 329.200 294.800 333.000 295.400 ;
        RECT 325.800 294.300 326.800 294.400 ;
        RECT 329.200 294.300 330.000 294.800 ;
        RECT 325.800 293.700 330.000 294.300 ;
        RECT 336.200 294.200 337.000 294.400 ;
        RECT 340.400 294.200 341.200 294.400 ;
        RECT 342.000 294.200 342.600 296.400 ;
        RECT 346.800 295.000 347.600 299.800 ;
        RECT 348.400 295.400 349.200 299.800 ;
        RECT 352.600 298.400 353.800 299.800 ;
        RECT 352.600 297.800 354.000 298.400 ;
        RECT 357.200 297.800 358.000 299.800 ;
        RECT 361.600 298.400 362.400 299.800 ;
        RECT 361.600 297.800 363.600 298.400 ;
        RECT 353.200 297.000 354.000 297.800 ;
        RECT 357.400 297.200 358.000 297.800 ;
        RECT 357.400 296.600 360.200 297.200 ;
        RECT 359.400 296.400 360.200 296.600 ;
        RECT 361.200 296.400 362.000 297.200 ;
        RECT 362.800 297.000 363.600 297.800 ;
        RECT 351.400 295.400 352.200 295.600 ;
        RECT 348.400 294.800 352.200 295.400 ;
        RECT 345.200 294.200 346.800 294.400 ;
        RECT 325.800 293.600 326.800 293.700 ;
        RECT 325.600 292.800 326.400 293.600 ;
        RECT 322.800 290.200 323.400 291.600 ;
        RECT 324.200 291.400 325.000 292.000 ;
        RECT 329.200 291.400 330.000 293.700 ;
        RECT 335.800 293.600 346.800 294.200 ;
        RECT 334.000 292.800 334.800 293.000 ;
        RECT 331.000 292.200 334.800 292.800 ;
        RECT 331.000 292.000 331.800 292.200 ;
        RECT 332.600 291.400 333.400 291.600 ;
        RECT 324.200 291.200 328.400 291.400 ;
        RECT 324.400 290.800 328.400 291.200 ;
        RECT 305.200 289.600 307.600 290.200 ;
        RECT 309.200 289.600 311.200 290.200 ;
        RECT 305.200 282.200 306.000 289.600 ;
        RECT 306.800 289.400 307.600 289.600 ;
        RECT 309.600 282.200 311.200 289.600 ;
        RECT 313.400 289.600 315.600 290.200 ;
        RECT 316.400 289.600 317.800 290.200 ;
        RECT 318.400 289.600 319.400 290.200 ;
        RECT 322.800 289.600 324.200 290.200 ;
        RECT 313.400 289.400 314.200 289.600 ;
        RECT 314.800 282.200 315.600 289.600 ;
        RECT 317.200 288.400 317.800 289.600 ;
        RECT 317.200 287.600 318.000 288.400 ;
        RECT 318.600 282.200 319.400 289.600 ;
        RECT 323.400 282.200 324.200 289.600 ;
        RECT 327.600 282.200 328.400 290.800 ;
        RECT 329.200 290.800 333.400 291.400 ;
        RECT 329.200 282.200 330.000 290.800 ;
        RECT 335.800 290.400 336.400 293.600 ;
        RECT 343.000 293.400 343.800 293.600 ;
        RECT 342.000 292.400 342.800 292.600 ;
        RECT 344.600 292.400 345.400 292.600 ;
        RECT 340.400 291.800 345.400 292.400 ;
        RECT 340.400 291.600 341.200 291.800 ;
        RECT 348.400 291.400 349.200 294.800 ;
        RECT 355.400 294.200 356.200 294.400 ;
        RECT 361.200 294.200 361.800 296.400 ;
        RECT 366.000 295.000 366.800 299.800 ;
        RECT 367.600 295.400 368.400 299.800 ;
        RECT 371.800 298.400 373.000 299.800 ;
        RECT 371.800 297.800 373.200 298.400 ;
        RECT 376.400 297.800 377.200 299.800 ;
        RECT 380.800 298.400 381.600 299.800 ;
        RECT 380.800 297.800 382.800 298.400 ;
        RECT 372.400 297.000 373.200 297.800 ;
        RECT 376.600 297.200 377.200 297.800 ;
        RECT 376.600 296.600 379.400 297.200 ;
        RECT 378.600 296.400 379.400 296.600 ;
        RECT 380.400 296.400 381.200 297.200 ;
        RECT 382.000 297.000 382.800 297.800 ;
        RECT 370.600 295.400 371.400 295.600 ;
        RECT 367.600 294.800 371.400 295.400 ;
        RECT 364.400 294.200 366.000 294.400 ;
        RECT 355.000 293.600 366.000 294.200 ;
        RECT 353.200 292.800 354.000 293.000 ;
        RECT 350.200 292.200 354.000 292.800 ;
        RECT 355.000 292.400 355.600 293.600 ;
        RECT 362.200 293.400 363.000 293.600 ;
        RECT 361.200 292.400 362.000 292.600 ;
        RECT 363.800 292.400 364.600 292.600 ;
        RECT 350.200 292.000 351.000 292.200 ;
        RECT 354.800 291.600 355.600 292.400 ;
        RECT 359.600 291.800 364.600 292.400 ;
        RECT 359.600 291.600 360.400 291.800 ;
        RECT 351.800 291.400 352.600 291.600 ;
        RECT 342.000 291.000 347.600 291.200 ;
        RECT 341.800 290.800 347.600 291.000 ;
        RECT 334.000 289.800 336.400 290.400 ;
        RECT 337.800 290.600 347.600 290.800 ;
        RECT 337.800 290.200 342.600 290.600 ;
        RECT 334.000 288.800 334.600 289.800 ;
        RECT 333.200 288.000 334.600 288.800 ;
        RECT 336.200 289.000 337.000 289.200 ;
        RECT 337.800 289.000 338.400 290.200 ;
        RECT 336.200 288.400 338.400 289.000 ;
        RECT 339.000 289.000 344.400 289.600 ;
        RECT 339.000 288.800 339.800 289.000 ;
        RECT 343.600 288.800 344.400 289.000 ;
        RECT 337.400 287.400 338.200 287.600 ;
        RECT 340.200 287.400 341.000 287.600 ;
        RECT 334.000 286.200 334.800 287.000 ;
        RECT 337.400 286.800 341.000 287.400 ;
        RECT 338.200 286.200 338.800 286.800 ;
        RECT 343.600 286.200 344.400 287.000 ;
        RECT 333.400 282.200 334.600 286.200 ;
        RECT 338.000 282.200 338.800 286.200 ;
        RECT 342.400 285.600 344.400 286.200 ;
        RECT 342.400 282.200 343.200 285.600 ;
        RECT 346.800 282.200 347.600 290.600 ;
        RECT 348.400 290.800 352.600 291.400 ;
        RECT 348.400 282.200 349.200 290.800 ;
        RECT 355.000 290.400 355.600 291.600 ;
        RECT 367.600 291.400 368.400 294.800 ;
        RECT 374.600 294.200 375.400 294.400 ;
        RECT 380.400 294.200 381.000 296.400 ;
        RECT 385.200 295.000 386.000 299.800 ;
        RECT 386.800 295.800 387.600 299.800 ;
        RECT 391.200 296.200 392.800 299.800 ;
        RECT 386.800 295.200 389.200 295.800 ;
        RECT 388.400 295.000 389.200 295.200 ;
        RECT 389.800 294.800 390.600 295.600 ;
        RECT 389.800 294.400 390.400 294.800 ;
        RECT 383.600 294.200 385.200 294.400 ;
        RECT 374.200 293.600 385.200 294.200 ;
        RECT 386.800 293.600 388.400 294.400 ;
        RECT 389.600 293.600 390.400 294.400 ;
        RECT 372.400 292.800 373.200 293.000 ;
        RECT 369.400 292.200 373.200 292.800 ;
        RECT 374.200 292.400 374.800 293.600 ;
        RECT 381.400 293.400 382.200 293.600 ;
        RECT 391.200 292.800 391.800 296.200 ;
        RECT 396.400 295.800 397.200 299.800 ;
        RECT 398.000 295.800 398.800 299.800 ;
        RECT 399.600 296.000 400.400 299.800 ;
        RECT 402.800 296.000 403.600 299.800 ;
        RECT 399.600 295.800 403.600 296.000 ;
        RECT 392.400 295.400 394.000 295.600 ;
        RECT 392.400 294.800 394.400 295.400 ;
        RECT 395.000 295.200 397.200 295.800 ;
        RECT 395.000 295.000 395.800 295.200 ;
        RECT 393.800 294.400 394.400 294.800 ;
        RECT 398.200 294.400 398.800 295.800 ;
        RECT 399.800 295.400 403.400 295.800 ;
        RECT 404.400 295.600 405.200 297.200 ;
        RECT 402.000 294.400 402.800 294.800 ;
        RECT 393.800 294.300 397.200 294.400 ;
        RECT 398.000 294.300 400.600 294.400 ;
        RECT 392.400 293.400 393.200 294.200 ;
        RECT 393.800 293.800 400.600 294.300 ;
        RECT 402.000 293.800 403.600 294.400 ;
        RECT 395.600 293.700 400.600 293.800 ;
        RECT 395.600 293.600 397.200 293.700 ;
        RECT 398.000 293.600 400.600 293.700 ;
        RECT 402.800 293.600 403.600 293.800 ;
        RECT 380.400 292.400 381.200 292.600 ;
        RECT 383.000 292.400 383.800 292.600 ;
        RECT 390.800 292.400 391.800 292.800 ;
        RECT 369.400 292.000 370.200 292.200 ;
        RECT 374.000 291.600 374.800 292.400 ;
        RECT 378.800 291.800 383.800 292.400 ;
        RECT 390.000 292.200 391.800 292.400 ;
        RECT 392.600 292.800 393.200 293.400 ;
        RECT 392.600 292.200 395.200 292.800 ;
        RECT 378.800 291.600 379.600 291.800 ;
        RECT 390.000 291.600 391.400 292.200 ;
        RECT 394.400 292.000 395.200 292.200 ;
        RECT 371.000 291.400 371.800 291.600 ;
        RECT 361.200 291.000 366.800 291.200 ;
        RECT 361.000 290.800 366.800 291.000 ;
        RECT 353.200 289.800 355.600 290.400 ;
        RECT 357.000 290.600 366.800 290.800 ;
        RECT 357.000 290.200 361.800 290.600 ;
        RECT 353.200 288.800 353.800 289.800 ;
        RECT 352.400 288.000 353.800 288.800 ;
        RECT 355.400 289.000 356.200 289.200 ;
        RECT 357.000 289.000 357.600 290.200 ;
        RECT 355.400 288.400 357.600 289.000 ;
        RECT 358.200 289.000 363.600 289.600 ;
        RECT 358.200 288.800 359.000 289.000 ;
        RECT 362.800 288.800 363.600 289.000 ;
        RECT 356.600 287.400 357.400 287.600 ;
        RECT 359.400 287.400 360.200 287.600 ;
        RECT 353.200 286.200 354.000 287.000 ;
        RECT 356.600 286.800 360.200 287.400 ;
        RECT 357.400 286.200 358.000 286.800 ;
        RECT 362.800 286.200 363.600 287.000 ;
        RECT 352.600 282.200 353.800 286.200 ;
        RECT 357.200 282.200 358.000 286.200 ;
        RECT 361.600 285.600 363.600 286.200 ;
        RECT 361.600 282.200 362.400 285.600 ;
        RECT 366.000 282.200 366.800 290.600 ;
        RECT 367.600 290.800 371.800 291.400 ;
        RECT 367.600 282.200 368.400 290.800 ;
        RECT 374.200 290.400 374.800 291.600 ;
        RECT 380.400 291.000 386.000 291.200 ;
        RECT 380.200 290.800 386.000 291.000 ;
        RECT 372.400 289.800 374.800 290.400 ;
        RECT 376.200 290.600 386.000 290.800 ;
        RECT 376.200 290.200 381.000 290.600 ;
        RECT 372.400 288.800 373.000 289.800 ;
        RECT 371.600 288.000 373.000 288.800 ;
        RECT 374.600 289.000 375.400 289.200 ;
        RECT 376.200 289.000 376.800 290.200 ;
        RECT 374.600 288.400 376.800 289.000 ;
        RECT 377.400 289.000 382.800 289.600 ;
        RECT 377.400 288.800 378.200 289.000 ;
        RECT 382.000 288.800 382.800 289.000 ;
        RECT 375.800 287.400 376.600 287.600 ;
        RECT 378.600 287.400 379.400 287.600 ;
        RECT 372.400 286.200 373.200 287.000 ;
        RECT 375.800 286.800 379.400 287.400 ;
        RECT 376.600 286.200 377.200 286.800 ;
        RECT 382.000 286.200 382.800 287.000 ;
        RECT 371.800 282.200 373.000 286.200 ;
        RECT 376.400 282.200 377.200 286.200 ;
        RECT 380.800 285.600 382.800 286.200 ;
        RECT 380.800 282.200 381.600 285.600 ;
        RECT 385.200 282.200 386.000 290.600 ;
        RECT 390.800 290.200 391.400 291.600 ;
        RECT 392.200 291.400 393.000 291.600 ;
        RECT 392.200 290.800 395.600 291.400 ;
        RECT 395.000 290.200 395.600 290.800 ;
        RECT 398.000 290.200 398.800 290.400 ;
        RECT 400.000 290.200 400.600 293.600 ;
        RECT 401.200 291.600 402.000 293.200 ;
        RECT 406.000 290.300 406.800 299.800 ;
        RECT 407.600 295.800 408.400 299.800 ;
        RECT 409.200 296.000 410.000 299.800 ;
        RECT 412.400 296.000 413.200 299.800 ;
        RECT 409.200 295.800 413.200 296.000 ;
        RECT 407.800 294.400 408.400 295.800 ;
        RECT 409.400 295.400 413.000 295.800 ;
        RECT 414.000 295.400 414.800 299.800 ;
        RECT 418.200 298.400 419.400 299.800 ;
        RECT 418.200 297.800 419.600 298.400 ;
        RECT 422.800 297.800 423.600 299.800 ;
        RECT 427.200 298.400 428.000 299.800 ;
        RECT 427.200 297.800 429.200 298.400 ;
        RECT 418.800 297.000 419.600 297.800 ;
        RECT 423.000 297.200 423.600 297.800 ;
        RECT 423.000 296.600 425.800 297.200 ;
        RECT 425.000 296.400 425.800 296.600 ;
        RECT 426.800 296.400 427.600 297.200 ;
        RECT 428.400 297.000 429.200 297.800 ;
        RECT 417.000 295.400 417.800 295.600 ;
        RECT 414.000 294.800 417.800 295.400 ;
        RECT 411.600 294.400 412.400 294.800 ;
        RECT 407.600 293.600 410.200 294.400 ;
        RECT 411.600 293.800 413.200 294.400 ;
        RECT 412.400 293.600 413.200 293.800 ;
        RECT 407.600 292.300 408.400 292.400 ;
        RECT 409.600 292.300 410.200 293.600 ;
        RECT 407.600 291.700 410.200 292.300 ;
        RECT 407.600 291.600 408.400 291.700 ;
        RECT 407.600 290.300 408.400 290.400 ;
        RECT 406.000 290.200 408.400 290.300 ;
        RECT 409.600 290.200 410.200 291.700 ;
        RECT 410.800 291.600 411.600 293.200 ;
        RECT 414.000 291.400 414.800 294.800 ;
        RECT 421.000 294.200 421.800 294.400 ;
        RECT 426.800 294.200 427.400 296.400 ;
        RECT 431.600 295.000 432.400 299.800 ;
        RECT 433.200 295.800 434.000 299.800 ;
        RECT 437.600 296.200 439.200 299.800 ;
        RECT 433.200 295.200 435.600 295.800 ;
        RECT 434.800 295.000 435.600 295.200 ;
        RECT 436.200 294.800 437.000 295.600 ;
        RECT 436.200 294.400 436.800 294.800 ;
        RECT 430.000 294.200 431.600 294.400 ;
        RECT 420.600 293.600 431.600 294.200 ;
        RECT 433.200 293.600 434.800 294.400 ;
        RECT 436.000 293.600 436.800 294.400 ;
        RECT 418.800 292.800 419.600 293.000 ;
        RECT 415.800 292.200 419.600 292.800 ;
        RECT 420.600 292.400 421.200 293.600 ;
        RECT 427.800 293.400 428.600 293.600 ;
        RECT 437.600 292.800 438.200 296.200 ;
        RECT 442.800 295.800 443.600 299.800 ;
        RECT 438.800 295.400 440.400 295.600 ;
        RECT 438.800 294.800 440.800 295.400 ;
        RECT 441.400 295.200 443.600 295.800 ;
        RECT 449.200 295.600 450.000 297.200 ;
        RECT 441.400 295.000 442.200 295.200 ;
        RECT 440.200 294.400 440.800 294.800 ;
        RECT 438.800 293.400 439.600 294.200 ;
        RECT 440.200 293.800 443.600 294.400 ;
        RECT 442.000 293.600 443.600 293.800 ;
        RECT 429.400 292.400 430.200 292.600 ;
        RECT 437.200 292.400 438.200 292.800 ;
        RECT 415.800 292.000 416.600 292.200 ;
        RECT 420.400 291.600 421.200 292.400 ;
        RECT 425.200 291.800 430.200 292.400 ;
        RECT 436.400 292.200 438.200 292.400 ;
        RECT 439.000 292.800 439.600 293.400 ;
        RECT 439.000 292.200 441.600 292.800 ;
        RECT 425.200 291.600 426.000 291.800 ;
        RECT 436.400 291.600 437.800 292.200 ;
        RECT 440.800 292.000 441.600 292.200 ;
        RECT 450.800 292.300 451.600 299.800 ;
        RECT 452.400 296.000 453.200 299.800 ;
        RECT 455.600 296.000 456.400 299.800 ;
        RECT 452.400 295.800 456.400 296.000 ;
        RECT 457.200 295.800 458.000 299.800 ;
        RECT 458.800 296.000 459.600 299.800 ;
        RECT 462.000 296.000 462.800 299.800 ;
        RECT 458.800 295.800 462.800 296.000 ;
        RECT 463.600 295.800 464.400 299.800 ;
        RECT 452.600 295.400 456.200 295.800 ;
        RECT 453.200 294.400 454.000 294.800 ;
        RECT 457.200 294.400 457.800 295.800 ;
        RECT 459.000 295.400 462.600 295.800 ;
        RECT 459.600 294.400 460.400 294.800 ;
        RECT 463.600 294.400 464.200 295.800 ;
        RECT 465.200 295.000 466.000 299.800 ;
        RECT 469.600 298.400 470.400 299.800 ;
        RECT 468.400 297.800 470.400 298.400 ;
        RECT 474.000 297.800 474.800 299.800 ;
        RECT 478.200 298.400 479.400 299.800 ;
        RECT 478.000 297.800 479.400 298.400 ;
        RECT 468.400 297.000 469.200 297.800 ;
        RECT 474.000 297.200 474.600 297.800 ;
        RECT 470.000 296.400 470.800 297.200 ;
        RECT 471.800 296.600 474.600 297.200 ;
        RECT 478.000 297.000 478.800 297.800 ;
        RECT 471.800 296.400 472.600 296.600 ;
        RECT 452.400 293.800 454.000 294.400 ;
        RECT 452.400 293.600 453.200 293.800 ;
        RECT 455.400 293.600 458.000 294.400 ;
        RECT 458.800 293.800 460.400 294.400 ;
        RECT 458.800 293.600 459.600 293.800 ;
        RECT 461.800 293.600 464.400 294.400 ;
        RECT 466.000 294.200 467.600 294.400 ;
        RECT 470.200 294.200 470.800 296.400 ;
        RECT 479.800 295.400 480.600 295.600 ;
        RECT 482.800 295.400 483.600 299.800 ;
        RECT 479.800 294.800 483.600 295.400 ;
        RECT 484.400 295.800 485.200 299.800 ;
        RECT 488.800 298.400 490.400 299.800 ;
        RECT 487.600 297.600 490.400 298.400 ;
        RECT 488.800 296.200 490.400 297.600 ;
        RECT 484.400 295.200 486.800 295.800 ;
        RECT 486.000 295.000 486.800 295.200 ;
        RECT 475.800 294.200 476.600 294.400 ;
        RECT 466.000 293.600 477.000 294.200 ;
        RECT 454.000 292.300 454.800 293.200 ;
        RECT 450.800 291.700 454.800 292.300 ;
        RECT 417.400 291.400 418.200 291.600 ;
        RECT 414.000 290.800 418.200 291.400 ;
        RECT 386.800 289.600 389.200 290.200 ;
        RECT 390.800 289.600 392.800 290.200 ;
        RECT 386.800 282.200 387.600 289.600 ;
        RECT 388.400 289.400 389.200 289.600 ;
        RECT 391.200 288.400 392.800 289.600 ;
        RECT 395.000 289.600 397.200 290.200 ;
        RECT 398.000 289.600 399.400 290.200 ;
        RECT 400.000 289.600 401.000 290.200 ;
        RECT 395.000 289.400 395.800 289.600 ;
        RECT 390.000 287.600 392.800 288.400 ;
        RECT 391.200 282.200 392.800 287.600 ;
        RECT 396.400 282.200 397.200 289.600 ;
        RECT 398.800 288.400 399.400 289.600 ;
        RECT 398.800 287.600 399.600 288.400 ;
        RECT 400.200 282.200 401.000 289.600 ;
        RECT 406.000 289.700 409.000 290.200 ;
        RECT 406.000 282.200 406.800 289.700 ;
        RECT 407.600 289.600 409.000 289.700 ;
        RECT 409.600 289.600 410.600 290.200 ;
        RECT 408.400 288.400 409.000 289.600 ;
        RECT 408.400 287.600 409.200 288.400 ;
        RECT 409.800 282.200 410.600 289.600 ;
        RECT 414.000 282.200 414.800 290.800 ;
        RECT 420.600 290.400 421.200 291.600 ;
        RECT 426.800 291.000 432.400 291.200 ;
        RECT 426.600 290.800 432.400 291.000 ;
        RECT 418.800 289.800 421.200 290.400 ;
        RECT 422.600 290.600 432.400 290.800 ;
        RECT 422.600 290.200 427.400 290.600 ;
        RECT 418.800 288.800 419.400 289.800 ;
        RECT 418.000 288.000 419.400 288.800 ;
        RECT 421.000 289.000 421.800 289.200 ;
        RECT 422.600 289.000 423.200 290.200 ;
        RECT 421.000 288.400 423.200 289.000 ;
        RECT 423.800 289.000 429.200 289.600 ;
        RECT 423.800 288.800 424.600 289.000 ;
        RECT 428.400 288.800 429.200 289.000 ;
        RECT 422.200 287.400 423.000 287.600 ;
        RECT 425.000 287.400 425.800 287.600 ;
        RECT 418.800 286.200 419.600 287.000 ;
        RECT 422.200 286.800 425.800 287.400 ;
        RECT 423.000 286.200 423.600 286.800 ;
        RECT 428.400 286.200 429.200 287.000 ;
        RECT 418.200 282.200 419.400 286.200 ;
        RECT 422.800 282.200 423.600 286.200 ;
        RECT 427.200 285.600 429.200 286.200 ;
        RECT 427.200 282.200 428.000 285.600 ;
        RECT 431.600 282.200 432.400 290.600 ;
        RECT 437.200 290.200 437.800 291.600 ;
        RECT 438.600 291.400 439.400 291.600 ;
        RECT 438.600 290.800 442.000 291.400 ;
        RECT 441.400 290.200 442.000 290.800 ;
        RECT 433.200 289.600 435.600 290.200 ;
        RECT 437.200 289.600 439.200 290.200 ;
        RECT 433.200 282.200 434.000 289.600 ;
        RECT 434.800 289.400 435.600 289.600 ;
        RECT 437.600 286.400 439.200 289.600 ;
        RECT 441.400 289.600 443.600 290.200 ;
        RECT 441.400 289.400 442.200 289.600 ;
        RECT 436.400 285.600 439.200 286.400 ;
        RECT 437.600 282.200 439.200 285.600 ;
        RECT 442.800 282.200 443.600 289.600 ;
        RECT 450.800 282.200 451.600 291.700 ;
        RECT 454.000 291.600 454.800 291.700 ;
        RECT 455.400 290.200 456.000 293.600 ;
        RECT 460.400 291.600 461.200 293.200 ;
        RECT 457.200 290.200 458.000 290.400 ;
        RECT 461.800 290.200 462.400 293.600 ;
        RECT 469.000 293.400 469.800 293.600 ;
        RECT 467.400 292.400 468.200 292.600 ;
        RECT 470.000 292.400 470.800 292.600 ;
        RECT 467.400 291.800 472.400 292.400 ;
        RECT 471.600 291.600 472.400 291.800 ;
        RECT 465.200 291.000 470.800 291.200 ;
        RECT 465.200 290.800 471.000 291.000 ;
        RECT 465.200 290.600 475.000 290.800 ;
        RECT 463.600 290.200 464.400 290.400 ;
        RECT 455.000 289.600 456.000 290.200 ;
        RECT 456.600 289.600 458.000 290.200 ;
        RECT 461.400 289.600 462.400 290.200 ;
        RECT 463.000 289.600 464.400 290.200 ;
        RECT 455.000 282.200 455.800 289.600 ;
        RECT 456.600 288.400 457.200 289.600 ;
        RECT 461.400 288.400 462.200 289.600 ;
        RECT 463.000 288.400 463.600 289.600 ;
        RECT 456.400 287.600 457.200 288.400 ;
        RECT 460.400 287.600 462.200 288.400 ;
        RECT 462.800 287.600 463.600 288.400 ;
        RECT 461.400 282.200 462.200 287.600 ;
        RECT 465.200 282.200 466.000 290.600 ;
        RECT 470.200 290.200 475.000 290.600 ;
        RECT 468.400 289.000 473.800 289.600 ;
        RECT 468.400 288.800 469.200 289.000 ;
        RECT 473.000 288.800 473.800 289.000 ;
        RECT 474.400 289.000 475.000 290.200 ;
        RECT 476.400 290.400 477.000 293.600 ;
        RECT 478.000 292.800 478.800 293.000 ;
        RECT 478.000 292.200 481.800 292.800 ;
        RECT 481.000 292.000 481.800 292.200 ;
        RECT 479.400 291.400 480.200 291.600 ;
        RECT 482.800 291.400 483.600 294.800 ;
        RECT 487.400 294.800 488.200 295.600 ;
        RECT 487.400 294.400 488.000 294.800 ;
        RECT 484.400 293.600 486.000 294.400 ;
        RECT 487.200 293.600 488.000 294.400 ;
        RECT 488.800 292.800 489.400 296.200 ;
        RECT 494.000 295.800 494.800 299.800 ;
        RECT 490.000 295.400 491.600 295.600 ;
        RECT 490.000 294.800 492.000 295.400 ;
        RECT 492.600 295.200 494.800 295.800 ;
        RECT 497.200 295.200 498.000 299.800 ;
        RECT 500.400 295.200 501.200 299.800 ;
        RECT 503.600 295.200 504.400 299.800 ;
        RECT 506.800 295.200 507.600 299.800 ;
        RECT 492.600 295.000 493.400 295.200 ;
        RECT 491.400 294.400 492.000 294.800 ;
        RECT 497.200 294.400 499.000 295.200 ;
        RECT 500.400 294.400 502.600 295.200 ;
        RECT 503.600 294.400 505.800 295.200 ;
        RECT 506.800 294.400 509.200 295.200 ;
        RECT 510.000 295.000 510.800 299.800 ;
        RECT 514.400 298.400 515.200 299.800 ;
        RECT 513.200 297.800 515.200 298.400 ;
        RECT 518.800 297.800 519.600 299.800 ;
        RECT 523.000 298.400 524.200 299.800 ;
        RECT 522.800 297.800 524.200 298.400 ;
        RECT 513.200 297.000 514.000 297.800 ;
        RECT 518.800 297.200 519.400 297.800 ;
        RECT 514.800 296.400 515.600 297.200 ;
        RECT 516.600 296.600 519.400 297.200 ;
        RECT 522.800 297.000 523.600 297.800 ;
        RECT 516.600 296.400 517.400 296.600 ;
        RECT 490.000 293.400 490.800 294.200 ;
        RECT 491.400 293.800 494.800 294.400 ;
        RECT 493.200 293.600 494.800 293.800 ;
        RECT 498.200 293.800 499.000 294.400 ;
        RECT 501.800 293.800 502.600 294.400 ;
        RECT 505.000 293.800 505.800 294.400 ;
        RECT 488.400 292.400 489.400 292.800 ;
        RECT 487.600 292.200 489.400 292.400 ;
        RECT 490.200 292.800 490.800 293.400 ;
        RECT 498.200 293.000 500.800 293.800 ;
        RECT 501.800 293.000 504.200 293.800 ;
        RECT 505.000 293.000 507.600 293.800 ;
        RECT 490.200 292.200 492.800 292.800 ;
        RECT 487.600 291.600 489.000 292.200 ;
        RECT 492.000 292.000 492.800 292.200 ;
        RECT 498.200 291.600 499.000 293.000 ;
        RECT 501.800 291.600 502.600 293.000 ;
        RECT 505.000 291.600 505.800 293.000 ;
        RECT 508.400 291.600 509.200 294.400 ;
        RECT 510.800 294.200 512.400 294.400 ;
        RECT 515.000 294.200 515.600 296.400 ;
        RECT 524.600 295.400 525.400 295.600 ;
        RECT 527.600 295.400 528.400 299.800 ;
        RECT 524.600 294.800 528.400 295.400 ;
        RECT 516.400 294.200 517.200 294.400 ;
        RECT 520.600 294.200 521.400 294.400 ;
        RECT 510.800 293.600 521.800 294.200 ;
        RECT 513.800 293.400 514.600 293.600 ;
        RECT 512.200 292.400 513.000 292.600 ;
        RECT 514.800 292.400 515.600 292.600 ;
        RECT 512.200 291.800 517.200 292.400 ;
        RECT 516.400 291.600 517.200 291.800 ;
        RECT 479.400 290.800 483.600 291.400 ;
        RECT 476.400 289.800 478.800 290.400 ;
        RECT 475.800 289.000 476.600 289.200 ;
        RECT 474.400 288.400 476.600 289.000 ;
        RECT 478.200 288.800 478.800 289.800 ;
        RECT 478.200 288.000 479.600 288.800 ;
        RECT 471.800 287.400 472.600 287.600 ;
        RECT 474.600 287.400 475.400 287.600 ;
        RECT 468.400 286.200 469.200 287.000 ;
        RECT 471.800 286.800 475.400 287.400 ;
        RECT 474.000 286.200 474.600 286.800 ;
        RECT 478.000 286.200 478.800 287.000 ;
        RECT 468.400 285.600 470.400 286.200 ;
        RECT 469.600 282.200 470.400 285.600 ;
        RECT 474.000 282.200 474.800 286.200 ;
        RECT 478.200 282.200 479.400 286.200 ;
        RECT 482.800 282.200 483.600 290.800 ;
        RECT 488.400 290.200 489.000 291.600 ;
        RECT 489.800 291.400 490.600 291.600 ;
        RECT 489.800 290.800 493.200 291.400 ;
        RECT 492.600 290.200 493.200 290.800 ;
        RECT 497.200 290.800 499.000 291.600 ;
        RECT 500.400 290.800 502.600 291.600 ;
        RECT 503.600 290.800 505.800 291.600 ;
        RECT 506.800 290.800 509.200 291.600 ;
        RECT 510.000 291.000 515.600 291.200 ;
        RECT 510.000 290.800 515.800 291.000 ;
        RECT 484.400 289.600 486.800 290.200 ;
        RECT 488.400 289.600 490.400 290.200 ;
        RECT 484.400 282.200 485.200 289.600 ;
        RECT 486.000 289.400 486.800 289.600 ;
        RECT 488.800 282.200 490.400 289.600 ;
        RECT 492.600 289.600 494.800 290.200 ;
        RECT 492.600 289.400 493.400 289.600 ;
        RECT 494.000 282.200 494.800 289.600 ;
        RECT 497.200 282.200 498.000 290.800 ;
        RECT 500.400 282.200 501.200 290.800 ;
        RECT 503.600 282.200 504.400 290.800 ;
        RECT 506.800 282.200 507.600 290.800 ;
        RECT 510.000 290.600 519.800 290.800 ;
        RECT 510.000 282.200 510.800 290.600 ;
        RECT 515.000 290.200 519.800 290.600 ;
        RECT 513.200 289.000 518.600 289.600 ;
        RECT 513.200 288.800 514.000 289.000 ;
        RECT 517.800 288.800 518.600 289.000 ;
        RECT 519.200 289.000 519.800 290.200 ;
        RECT 521.200 290.400 521.800 293.600 ;
        RECT 522.800 292.800 523.600 293.000 ;
        RECT 522.800 292.200 526.600 292.800 ;
        RECT 525.800 292.000 526.600 292.200 ;
        RECT 524.200 291.400 525.000 291.600 ;
        RECT 527.600 291.400 528.400 294.800 ;
        RECT 524.200 290.800 528.400 291.400 ;
        RECT 521.200 289.800 523.600 290.400 ;
        RECT 520.600 289.000 521.400 289.200 ;
        RECT 519.200 288.400 521.400 289.000 ;
        RECT 523.000 288.800 523.600 289.800 ;
        RECT 523.000 288.400 524.400 288.800 ;
        RECT 523.000 288.000 525.200 288.400 ;
        RECT 523.800 287.600 525.200 288.000 ;
        RECT 516.600 287.400 517.400 287.600 ;
        RECT 519.400 287.400 520.200 287.600 ;
        RECT 513.200 286.200 514.000 287.000 ;
        RECT 516.600 286.800 520.200 287.400 ;
        RECT 518.800 286.200 519.400 286.800 ;
        RECT 522.800 286.200 523.600 287.000 ;
        RECT 513.200 285.600 515.200 286.200 ;
        RECT 514.400 282.200 515.200 285.600 ;
        RECT 518.800 282.200 519.600 286.200 ;
        RECT 523.000 282.200 524.200 286.200 ;
        RECT 527.600 282.200 528.400 290.800 ;
        RECT 529.200 292.400 530.000 299.800 ;
        RECT 532.400 295.200 533.200 299.800 ;
        RECT 535.600 296.000 536.400 299.800 ;
        RECT 531.000 294.600 533.200 295.200 ;
        RECT 535.400 295.200 536.400 296.000 ;
        RECT 529.200 290.200 529.800 292.400 ;
        RECT 531.000 291.600 531.600 294.600 ;
        RECT 532.400 292.300 533.200 293.200 ;
        RECT 535.400 292.300 536.200 295.200 ;
        RECT 537.200 294.600 538.000 299.800 ;
        RECT 543.600 296.600 544.400 299.800 ;
        RECT 545.200 297.000 546.000 299.800 ;
        RECT 546.800 297.000 547.600 299.800 ;
        RECT 548.400 297.000 549.200 299.800 ;
        RECT 550.000 297.000 550.800 299.800 ;
        RECT 553.200 297.000 554.000 299.800 ;
        RECT 556.400 297.000 557.200 299.800 ;
        RECT 558.000 297.000 558.800 299.800 ;
        RECT 559.600 297.000 560.400 299.800 ;
        RECT 542.000 295.800 544.400 296.600 ;
        RECT 561.200 296.600 562.000 299.800 ;
        RECT 542.000 295.200 542.800 295.800 ;
        RECT 532.400 291.700 536.200 292.300 ;
        RECT 532.400 291.600 533.200 291.700 ;
        RECT 530.400 290.800 531.600 291.600 ;
        RECT 531.000 290.200 531.600 290.800 ;
        RECT 535.400 290.800 536.200 291.700 ;
        RECT 536.800 294.000 538.000 294.600 ;
        RECT 541.000 294.600 542.800 295.200 ;
        RECT 546.800 295.600 547.800 296.400 ;
        RECT 550.800 295.600 552.400 296.400 ;
        RECT 553.200 295.800 557.800 296.400 ;
        RECT 561.200 295.800 563.800 296.600 ;
        RECT 553.200 295.600 554.000 295.800 ;
        RECT 536.800 292.000 537.400 294.000 ;
        RECT 541.000 293.400 541.800 294.600 ;
        RECT 538.000 292.600 541.800 293.400 ;
        RECT 546.800 292.800 547.600 295.600 ;
        RECT 553.200 294.800 554.000 295.000 ;
        RECT 549.600 294.200 554.000 294.800 ;
        RECT 549.600 294.000 550.400 294.200 ;
        RECT 557.000 293.400 557.800 295.800 ;
        RECT 563.000 295.200 563.800 295.800 ;
        RECT 563.000 294.400 566.000 295.200 ;
        RECT 567.600 293.800 568.400 299.800 ;
        RECT 571.800 296.400 572.600 299.800 ;
        RECT 550.000 292.600 553.200 293.400 ;
        RECT 557.000 292.600 559.000 293.400 ;
        RECT 559.600 293.000 568.400 293.800 ;
        RECT 543.600 292.000 544.400 292.600 ;
        RECT 561.200 292.000 562.000 292.400 ;
        RECT 564.400 292.000 565.200 292.400 ;
        RECT 566.200 292.000 567.000 292.200 ;
        RECT 536.800 291.400 537.600 292.000 ;
        RECT 543.600 291.400 567.000 292.000 ;
        RECT 529.200 282.200 530.000 290.200 ;
        RECT 531.000 289.600 533.200 290.200 ;
        RECT 535.400 290.000 536.400 290.800 ;
        RECT 532.400 282.200 533.200 289.600 ;
        RECT 535.600 282.200 536.400 290.000 ;
        RECT 537.000 289.600 537.600 291.400 ;
        RECT 538.200 290.800 539.000 291.000 ;
        RECT 538.200 290.200 565.200 290.800 ;
        RECT 561.000 290.000 561.800 290.200 ;
        RECT 564.400 289.600 565.200 290.200 ;
        RECT 537.000 289.000 546.000 289.600 ;
        RECT 537.000 287.400 537.600 289.000 ;
        RECT 545.200 288.800 546.000 289.000 ;
        RECT 548.400 289.000 557.000 289.600 ;
        RECT 548.400 288.800 549.200 289.000 ;
        RECT 540.200 287.600 542.800 288.400 ;
        RECT 537.000 286.800 539.600 287.400 ;
        RECT 538.800 282.200 539.600 286.800 ;
        RECT 542.000 282.200 542.800 287.600 ;
        RECT 543.400 286.800 547.600 287.600 ;
        RECT 545.200 282.200 546.000 285.000 ;
        RECT 546.800 282.200 547.600 285.000 ;
        RECT 548.400 282.200 549.200 285.000 ;
        RECT 550.000 282.200 550.800 288.400 ;
        RECT 553.200 287.600 555.800 288.400 ;
        RECT 556.400 288.200 557.000 289.000 ;
        RECT 558.000 289.400 558.800 289.600 ;
        RECT 558.000 289.000 563.400 289.400 ;
        RECT 558.000 288.800 564.200 289.000 ;
        RECT 562.800 288.200 564.200 288.800 ;
        RECT 556.400 287.600 562.200 288.200 ;
        RECT 565.200 288.000 566.800 288.800 ;
        RECT 565.200 287.600 565.800 288.000 ;
        RECT 553.200 282.200 554.000 287.000 ;
        RECT 556.400 282.200 557.200 287.000 ;
        RECT 561.600 286.800 565.800 287.600 ;
        RECT 567.600 287.400 568.400 293.000 ;
        RECT 570.800 295.800 572.600 296.400 ;
        RECT 574.000 295.800 574.800 299.800 ;
        RECT 577.200 297.800 578.000 299.800 ;
        RECT 569.200 290.300 570.000 290.400 ;
        RECT 570.800 290.300 571.600 295.800 ;
        RECT 569.200 289.700 571.600 290.300 ;
        RECT 569.200 289.600 570.000 289.700 ;
        RECT 566.400 286.800 568.400 287.400 ;
        RECT 558.000 282.200 558.800 285.000 ;
        RECT 559.600 282.200 560.400 285.000 ;
        RECT 562.800 282.200 563.600 286.800 ;
        RECT 566.400 286.200 567.000 286.800 ;
        RECT 566.000 285.600 567.000 286.200 ;
        RECT 566.000 282.200 566.800 285.600 ;
        RECT 570.800 282.200 571.600 289.700 ;
        RECT 574.000 292.400 574.600 295.800 ;
        RECT 577.200 295.600 577.800 297.800 ;
        RECT 578.800 295.600 579.600 297.200 ;
        RECT 575.400 295.000 577.800 295.600 ;
        RECT 580.400 295.200 581.200 299.800 ;
        RECT 574.000 291.600 574.800 292.400 ;
        RECT 575.400 292.000 576.000 295.000 ;
        RECT 580.400 294.600 582.600 295.200 ;
        RECT 574.000 290.200 574.600 291.600 ;
        RECT 575.400 291.400 576.200 292.000 ;
        RECT 580.400 291.600 581.200 293.200 ;
        RECT 582.000 291.600 582.600 294.600 ;
        RECT 575.400 291.200 579.600 291.400 ;
        RECT 575.600 290.800 579.600 291.200 ;
        RECT 574.000 289.600 575.400 290.200 ;
        RECT 574.600 282.200 575.400 289.600 ;
        RECT 578.800 282.200 579.600 290.800 ;
        RECT 582.000 290.800 583.200 291.600 ;
        RECT 582.000 290.200 582.600 290.800 ;
        RECT 580.400 289.600 582.600 290.200 ;
        RECT 580.400 282.200 581.200 289.600 ;
        RECT 1.200 271.800 2.000 279.800 ;
        RECT 2.800 272.400 3.600 279.800 ;
        RECT 6.000 272.400 6.800 279.800 ;
        RECT 2.800 271.800 6.800 272.400 ;
        RECT 7.600 272.400 8.400 279.800 ;
        RECT 9.200 272.400 10.000 272.600 ;
        RECT 7.600 271.800 10.000 272.400 ;
        RECT 12.000 271.800 13.600 279.800 ;
        RECT 15.400 272.400 16.200 272.600 ;
        RECT 17.200 272.400 18.000 279.800 ;
        RECT 18.800 274.300 19.600 274.400 ;
        RECT 20.400 274.300 21.200 279.800 ;
        RECT 18.800 273.700 21.200 274.300 ;
        RECT 18.800 273.600 19.600 273.700 ;
        RECT 15.400 271.800 18.000 272.400 ;
        RECT 1.400 270.400 2.000 271.800 ;
        RECT 5.200 270.400 6.000 270.800 ;
        RECT 12.400 270.400 13.000 271.800 ;
        RECT 14.200 270.400 15.000 270.600 ;
        RECT 1.200 269.800 3.600 270.400 ;
        RECT 5.200 269.800 6.800 270.400 ;
        RECT 1.200 269.600 2.000 269.800 ;
        RECT 1.200 265.600 2.000 266.400 ;
        RECT 3.000 266.200 3.600 269.800 ;
        RECT 6.000 269.600 6.800 269.800 ;
        RECT 12.400 269.600 13.200 270.400 ;
        RECT 14.200 269.800 15.800 270.400 ;
        RECT 15.000 269.600 15.800 269.800 ;
        RECT 4.400 267.600 5.200 269.200 ;
        RECT 12.400 268.400 13.000 269.600 ;
        RECT 7.600 267.600 9.200 268.400 ;
        RECT 10.400 267.600 11.200 268.400 ;
        RECT 10.600 267.200 11.200 267.600 ;
        RECT 12.000 267.800 13.000 268.400 ;
        RECT 13.600 268.600 14.400 268.800 ;
        RECT 13.600 268.400 16.400 268.600 ;
        RECT 13.600 268.000 18.000 268.400 ;
        RECT 15.800 267.800 18.000 268.000 ;
        RECT 9.200 266.800 10.000 267.000 ;
        RECT 1.400 264.800 2.200 265.600 ;
        RECT 2.800 262.200 3.600 266.200 ;
        RECT 7.600 266.200 10.000 266.800 ;
        RECT 10.600 266.400 11.400 267.200 ;
        RECT 7.600 262.200 8.400 266.200 ;
        RECT 12.000 265.800 12.600 267.800 ;
        RECT 16.400 267.600 18.000 267.800 ;
        RECT 13.200 266.400 14.800 267.200 ;
        RECT 15.400 266.800 16.200 267.000 ;
        RECT 15.400 266.200 18.000 266.800 ;
        RECT 12.000 262.200 13.600 265.800 ;
        RECT 17.200 262.200 18.000 266.200 ;
        RECT 18.800 264.800 19.600 266.400 ;
        RECT 20.400 262.200 21.200 273.700 ;
        RECT 22.800 273.600 23.600 274.400 ;
        RECT 22.800 272.400 23.400 273.600 ;
        RECT 24.200 272.400 25.000 279.800 ;
        RECT 22.000 271.800 23.400 272.400 ;
        RECT 24.000 271.800 25.000 272.400 ;
        RECT 22.000 271.600 22.800 271.800 ;
        RECT 24.000 268.400 24.600 271.800 ;
        RECT 25.200 270.300 26.000 270.400 ;
        RECT 26.800 270.300 27.600 270.400 ;
        RECT 25.200 269.700 27.600 270.300 ;
        RECT 25.200 268.800 26.000 269.700 ;
        RECT 26.800 269.600 27.600 269.700 ;
        RECT 22.000 267.600 24.600 268.400 ;
        RECT 26.800 268.300 27.600 268.400 ;
        RECT 26.800 268.200 29.100 268.300 ;
        RECT 26.000 267.700 29.100 268.200 ;
        RECT 26.000 267.600 27.600 267.700 ;
        RECT 22.200 266.200 22.800 267.600 ;
        RECT 26.000 267.200 26.800 267.600 ;
        RECT 23.800 266.200 27.400 266.600 ;
        RECT 28.500 266.400 29.100 267.700 ;
        RECT 22.000 262.200 22.800 266.200 ;
        RECT 23.600 266.000 27.600 266.200 ;
        RECT 23.600 262.200 24.400 266.000 ;
        RECT 26.800 262.200 27.600 266.000 ;
        RECT 28.400 264.800 29.200 266.400 ;
        RECT 30.000 262.200 30.800 279.800 ;
        RECT 32.400 273.600 33.200 274.400 ;
        RECT 32.400 272.400 33.000 273.600 ;
        RECT 33.800 272.400 34.600 279.800 ;
        RECT 31.600 271.800 33.000 272.400 ;
        RECT 33.600 271.800 34.600 272.400 ;
        RECT 38.000 271.800 38.800 279.800 ;
        RECT 39.600 272.400 40.400 279.800 ;
        RECT 42.800 272.400 43.600 279.800 ;
        RECT 39.600 271.800 43.600 272.400 ;
        RECT 31.600 271.600 32.400 271.800 ;
        RECT 33.600 268.400 34.200 271.800 ;
        RECT 38.200 270.400 38.800 271.800 ;
        RECT 42.000 270.400 42.800 270.800 ;
        RECT 34.800 268.800 35.600 270.400 ;
        RECT 38.000 269.800 40.400 270.400 ;
        RECT 42.000 269.800 43.600 270.400 ;
        RECT 38.000 269.600 38.800 269.800 ;
        RECT 31.600 267.600 34.200 268.400 ;
        RECT 36.400 268.200 37.200 268.400 ;
        RECT 35.600 267.600 37.200 268.200 ;
        RECT 31.800 266.200 32.400 267.600 ;
        RECT 35.600 267.200 36.400 267.600 ;
        RECT 33.400 266.200 37.000 266.600 ;
        RECT 31.600 262.200 32.400 266.200 ;
        RECT 33.200 266.000 37.200 266.200 ;
        RECT 33.200 262.200 34.000 266.000 ;
        RECT 36.400 262.200 37.200 266.000 ;
        RECT 38.000 265.600 38.800 266.400 ;
        RECT 39.800 266.200 40.400 269.800 ;
        RECT 42.800 269.600 43.600 269.800 ;
        RECT 41.200 268.300 42.000 269.200 ;
        RECT 44.400 268.300 45.200 279.800 ;
        RECT 47.600 272.400 48.400 279.800 ;
        RECT 50.800 279.200 54.800 279.800 ;
        RECT 50.800 272.400 51.600 279.200 ;
        RECT 47.600 271.800 51.600 272.400 ;
        RECT 52.400 271.800 53.200 278.600 ;
        RECT 54.000 271.800 54.800 279.200 ;
        RECT 52.400 271.200 53.000 271.800 ;
        RECT 48.400 270.400 49.200 270.800 ;
        RECT 51.000 270.600 53.000 271.200 ;
        RECT 51.000 270.400 51.600 270.600 ;
        RECT 47.600 269.800 49.200 270.400 ;
        RECT 47.600 269.600 48.400 269.800 ;
        RECT 50.800 269.600 51.600 270.400 ;
        RECT 54.000 270.300 54.800 271.200 ;
        RECT 55.600 270.300 56.400 270.400 ;
        RECT 54.000 269.700 56.400 270.300 ;
        RECT 54.000 269.600 54.800 269.700 ;
        RECT 55.600 269.600 56.400 269.700 ;
        RECT 41.200 267.700 45.200 268.300 ;
        RECT 41.200 267.600 42.000 267.700 ;
        RECT 38.200 264.800 39.000 265.600 ;
        RECT 39.600 262.200 40.400 266.200 ;
        RECT 44.400 262.200 45.200 267.700 ;
        RECT 46.000 268.300 46.800 268.400 ;
        RECT 49.200 268.300 50.000 269.200 ;
        RECT 46.000 267.700 50.000 268.300 ;
        RECT 46.000 267.600 46.800 267.700 ;
        RECT 49.200 267.600 50.000 267.700 ;
        RECT 46.000 264.800 46.800 266.400 ;
        RECT 51.000 266.200 51.600 269.600 ;
        RECT 52.200 268.800 53.000 269.600 ;
        RECT 52.400 268.400 53.000 268.800 ;
        RECT 52.400 267.600 53.200 268.400 ;
        RECT 50.600 262.200 52.200 266.200 ;
        RECT 55.600 264.800 56.400 266.400 ;
        RECT 57.200 262.200 58.000 279.800 ;
        RECT 58.800 272.400 59.600 279.800 ;
        RECT 60.400 272.400 61.200 272.600 ;
        RECT 63.200 272.400 64.800 279.800 ;
        RECT 58.800 271.800 61.200 272.400 ;
        RECT 62.800 271.800 64.800 272.400 ;
        RECT 67.000 272.400 67.800 272.600 ;
        RECT 68.400 272.400 69.200 279.800 ;
        RECT 67.000 271.800 69.200 272.400 ;
        RECT 70.000 275.000 70.800 279.000 ;
        RECT 62.800 270.400 63.400 271.800 ;
        RECT 67.000 271.200 67.600 271.800 ;
        RECT 64.200 270.600 67.600 271.200 ;
        RECT 70.000 271.600 70.600 275.000 ;
        RECT 74.200 272.800 75.000 279.800 ;
        RECT 80.400 273.600 81.200 274.400 ;
        RECT 74.200 272.200 75.800 272.800 ;
        RECT 80.400 272.400 81.000 273.600 ;
        RECT 81.800 272.400 82.600 279.800 ;
        RECT 70.000 271.000 73.800 271.600 ;
        RECT 64.200 270.400 65.000 270.600 ;
        RECT 62.000 269.800 63.400 270.400 ;
        RECT 68.400 270.300 69.200 270.400 ;
        RECT 70.000 270.300 70.800 270.400 ;
        RECT 66.400 269.800 67.200 270.000 ;
        RECT 62.000 269.600 63.800 269.800 ;
        RECT 62.800 269.200 63.800 269.600 ;
        RECT 58.800 267.600 60.400 268.400 ;
        RECT 61.600 267.600 62.400 268.400 ;
        RECT 61.800 267.200 62.400 267.600 ;
        RECT 60.400 266.800 61.200 267.000 ;
        RECT 58.800 266.200 61.200 266.800 ;
        RECT 61.800 266.400 62.600 267.200 ;
        RECT 58.800 262.200 59.600 266.200 ;
        RECT 63.200 265.800 63.800 269.200 ;
        RECT 64.600 269.200 67.200 269.800 ;
        RECT 68.400 269.700 70.800 270.300 ;
        RECT 68.400 269.600 69.200 269.700 ;
        RECT 64.600 268.600 65.200 269.200 ;
        RECT 70.000 268.800 70.800 269.700 ;
        RECT 71.600 268.800 72.400 270.400 ;
        RECT 73.200 269.000 73.800 271.000 ;
        RECT 64.400 267.800 65.200 268.600 ;
        RECT 67.600 268.200 69.200 268.400 ;
        RECT 65.800 267.600 69.200 268.200 ;
        RECT 73.200 268.200 74.600 269.000 ;
        RECT 75.200 268.400 75.800 272.200 ;
        RECT 79.600 271.800 81.000 272.400 ;
        RECT 81.600 271.800 82.600 272.400 ;
        RECT 86.000 272.400 86.800 279.800 ;
        RECT 87.400 272.400 88.200 272.600 ;
        RECT 86.000 271.800 88.200 272.400 ;
        RECT 90.400 272.400 92.000 279.800 ;
        RECT 94.000 272.400 94.800 272.600 ;
        RECT 95.600 272.400 96.400 279.800 ;
        RECT 90.400 271.800 92.400 272.400 ;
        RECT 94.000 271.800 96.400 272.400 ;
        RECT 97.200 272.400 98.000 279.800 ;
        RECT 100.400 272.400 101.200 279.800 ;
        RECT 97.200 271.800 101.200 272.400 ;
        RECT 102.000 271.800 102.800 279.800 ;
        RECT 79.600 271.600 80.400 271.800 ;
        RECT 76.400 269.600 77.200 271.200 ;
        RECT 81.600 268.400 82.200 271.800 ;
        RECT 87.600 271.200 88.200 271.800 ;
        RECT 87.600 270.600 91.000 271.200 ;
        RECT 90.200 270.400 91.000 270.600 ;
        RECT 91.800 270.400 92.400 271.800 ;
        RECT 98.000 270.400 98.800 270.800 ;
        RECT 102.000 270.400 102.600 271.800 ;
        RECT 82.800 268.800 83.600 270.400 ;
        RECT 88.000 269.800 88.800 270.000 ;
        RECT 91.800 269.800 93.200 270.400 ;
        RECT 88.000 269.200 90.600 269.800 ;
        RECT 90.000 268.600 90.600 269.200 ;
        RECT 91.400 269.600 93.200 269.800 ;
        RECT 97.200 269.800 98.800 270.400 ;
        RECT 100.400 269.800 102.800 270.400 ;
        RECT 97.200 269.600 98.000 269.800 ;
        RECT 91.400 269.200 92.400 269.600 ;
        RECT 73.200 267.800 74.200 268.200 ;
        RECT 65.800 267.200 66.400 267.600 ;
        RECT 64.400 266.600 66.400 267.200 ;
        RECT 70.000 267.200 74.200 267.800 ;
        RECT 75.200 267.600 77.200 268.400 ;
        RECT 79.600 267.600 82.200 268.400 ;
        RECT 84.400 268.200 85.200 268.400 ;
        RECT 83.600 267.600 85.200 268.200 ;
        RECT 86.000 268.200 87.600 268.400 ;
        RECT 86.000 267.600 89.400 268.200 ;
        RECT 90.000 267.800 90.800 268.600 ;
        RECT 67.000 266.800 67.800 267.000 ;
        RECT 64.400 266.400 66.000 266.600 ;
        RECT 67.000 266.200 69.200 266.800 ;
        RECT 63.200 264.400 64.800 265.800 ;
        RECT 62.000 263.600 64.800 264.400 ;
        RECT 63.200 262.200 64.800 263.600 ;
        RECT 68.400 262.200 69.200 266.200 ;
        RECT 70.000 265.000 70.600 267.200 ;
        RECT 75.200 267.000 75.800 267.600 ;
        RECT 75.000 266.600 75.800 267.000 ;
        RECT 74.200 266.000 75.800 266.600 ;
        RECT 79.800 266.200 80.400 267.600 ;
        RECT 83.600 267.200 84.400 267.600 ;
        RECT 88.800 267.200 89.400 267.600 ;
        RECT 87.400 266.800 88.200 267.000 ;
        RECT 81.400 266.200 85.000 266.600 ;
        RECT 86.000 266.200 88.200 266.800 ;
        RECT 88.800 266.600 90.800 267.200 ;
        RECT 89.200 266.400 90.800 266.600 ;
        RECT 70.000 263.000 70.800 265.000 ;
        RECT 74.200 264.400 75.000 266.000 ;
        RECT 73.200 263.600 75.000 264.400 ;
        RECT 74.200 263.000 75.000 263.600 ;
        RECT 79.600 262.200 80.400 266.200 ;
        RECT 81.200 266.000 85.200 266.200 ;
        RECT 81.200 262.200 82.000 266.000 ;
        RECT 84.400 262.200 85.200 266.000 ;
        RECT 86.000 262.200 86.800 266.200 ;
        RECT 91.400 265.800 92.000 269.200 ;
        RECT 92.800 267.600 93.600 268.400 ;
        RECT 94.800 267.600 96.400 268.400 ;
        RECT 98.800 267.600 99.600 269.200 ;
        RECT 92.800 267.200 93.400 267.600 ;
        RECT 92.600 266.400 93.400 267.200 ;
        RECT 94.000 266.800 94.800 267.000 ;
        RECT 94.000 266.200 96.400 266.800 ;
        RECT 90.400 264.400 92.000 265.800 ;
        RECT 90.400 263.600 93.200 264.400 ;
        RECT 90.400 262.200 92.000 263.600 ;
        RECT 95.600 262.200 96.400 266.200 ;
        RECT 100.400 266.400 101.000 269.800 ;
        RECT 102.000 269.600 102.800 269.800 ;
        RECT 102.000 268.300 102.800 268.400 ;
        RECT 103.600 268.300 104.400 279.800 ;
        RECT 109.400 272.600 110.200 279.800 ;
        RECT 108.400 271.800 110.200 272.600 ;
        RECT 111.600 272.400 112.400 279.800 ;
        RECT 114.800 272.800 115.600 279.800 ;
        RECT 118.800 273.600 119.600 274.400 ;
        RECT 111.600 271.800 114.200 272.400 ;
        RECT 114.800 271.800 115.800 272.800 ;
        RECT 118.800 272.400 119.400 273.600 ;
        RECT 120.200 272.400 121.000 279.800 ;
        RECT 108.600 268.400 109.200 271.800 ;
        RECT 110.000 269.600 110.800 271.200 ;
        RECT 111.600 269.600 112.600 270.400 ;
        RECT 111.800 268.800 112.600 269.600 ;
        RECT 113.600 269.800 114.200 271.800 ;
        RECT 113.600 269.000 114.600 269.800 ;
        RECT 108.400 268.300 109.200 268.400 ;
        RECT 102.000 267.700 104.400 268.300 ;
        RECT 102.000 267.600 102.800 267.700 ;
        RECT 100.400 262.200 101.200 266.400 ;
        RECT 102.000 265.600 102.800 266.400 ;
        RECT 101.800 264.800 102.600 265.600 ;
        RECT 103.600 262.200 104.400 267.700 ;
        RECT 105.300 267.700 109.200 268.300 ;
        RECT 105.300 266.400 105.900 267.700 ;
        RECT 108.400 267.600 109.200 267.700 ;
        RECT 105.200 264.800 106.000 266.400 ;
        RECT 106.800 264.800 107.600 266.400 ;
        RECT 108.600 264.200 109.200 267.600 ;
        RECT 113.600 267.400 114.200 269.000 ;
        RECT 115.200 268.400 115.800 271.800 ;
        RECT 118.000 271.800 119.400 272.400 ;
        RECT 120.000 271.800 121.000 272.400 ;
        RECT 118.000 271.600 118.800 271.800 ;
        RECT 120.000 268.400 120.600 271.800 ;
        RECT 121.200 268.800 122.000 270.400 ;
        RECT 122.800 270.300 123.600 270.400 ;
        RECT 126.000 270.300 126.800 279.800 ;
        RECT 128.400 273.600 129.200 274.400 ;
        RECT 128.400 272.400 129.000 273.600 ;
        RECT 129.800 272.400 130.600 279.800 ;
        RECT 127.600 271.800 129.000 272.400 ;
        RECT 129.600 271.800 130.600 272.400 ;
        RECT 127.600 271.600 128.400 271.800 ;
        RECT 122.800 269.700 126.800 270.300 ;
        RECT 122.800 269.600 123.600 269.700 ;
        RECT 114.800 268.300 115.800 268.400 ;
        RECT 116.400 268.300 117.200 268.400 ;
        RECT 114.800 267.700 117.200 268.300 ;
        RECT 114.800 267.600 115.800 267.700 ;
        RECT 116.400 267.600 117.200 267.700 ;
        RECT 118.000 267.600 120.600 268.400 ;
        RECT 122.800 268.300 123.600 268.400 ;
        RECT 124.400 268.300 125.200 268.400 ;
        RECT 122.800 268.200 125.200 268.300 ;
        RECT 122.000 267.700 125.200 268.200 ;
        RECT 122.000 267.600 123.600 267.700 ;
        RECT 108.400 262.200 109.200 264.200 ;
        RECT 111.600 266.800 114.200 267.400 ;
        RECT 111.600 262.200 112.400 266.800 ;
        RECT 115.200 266.200 115.800 267.600 ;
        RECT 118.200 266.200 118.800 267.600 ;
        RECT 122.000 267.200 122.800 267.600 ;
        RECT 124.400 266.800 125.200 267.700 ;
        RECT 119.800 266.200 123.400 266.600 ;
        RECT 114.800 265.600 115.800 266.200 ;
        RECT 114.800 262.200 115.600 265.600 ;
        RECT 118.000 262.200 118.800 266.200 ;
        RECT 119.600 266.000 123.600 266.200 ;
        RECT 119.600 262.200 120.400 266.000 ;
        RECT 122.800 262.200 123.600 266.000 ;
        RECT 126.000 262.200 126.800 269.700 ;
        RECT 129.600 268.400 130.200 271.800 ;
        RECT 130.800 268.800 131.600 270.400 ;
        RECT 127.600 267.600 130.200 268.400 ;
        RECT 132.400 268.200 133.200 268.400 ;
        RECT 131.600 267.600 133.200 268.200 ;
        RECT 127.800 266.200 128.400 267.600 ;
        RECT 131.600 267.200 132.400 267.600 ;
        RECT 134.000 266.800 134.800 268.400 ;
        RECT 135.600 268.300 136.400 279.800 ;
        RECT 137.200 271.600 138.000 273.200 ;
        RECT 146.200 272.400 147.000 279.800 ;
        RECT 147.600 273.600 148.400 274.400 ;
        RECT 147.800 272.400 148.400 273.600 ;
        RECT 150.800 273.600 151.600 274.400 ;
        RECT 150.800 272.400 151.400 273.600 ;
        RECT 152.200 272.400 153.000 279.800 ;
        RECT 146.200 271.800 147.200 272.400 ;
        RECT 147.800 271.800 149.200 272.400 ;
        RECT 146.600 270.400 147.200 271.800 ;
        RECT 148.400 271.600 149.200 271.800 ;
        RECT 150.000 271.800 151.400 272.400 ;
        RECT 150.000 271.600 150.800 271.800 ;
        RECT 152.000 271.600 154.000 272.400 ;
        RECT 145.200 268.800 146.000 270.400 ;
        RECT 146.600 269.600 147.600 270.400 ;
        RECT 146.600 268.400 147.200 269.600 ;
        RECT 152.000 268.400 152.600 271.600 ;
        RECT 153.200 270.300 154.000 270.400 ;
        RECT 156.400 270.300 157.200 279.800 ;
        RECT 162.200 271.800 164.200 279.800 ;
        RECT 170.200 272.400 171.000 279.800 ;
        RECT 171.600 273.600 172.400 274.400 ;
        RECT 171.800 272.400 172.400 273.600 ;
        RECT 170.200 271.800 171.200 272.400 ;
        RECT 171.800 271.800 173.200 272.400 ;
        RECT 163.000 270.400 163.600 271.800 ;
        RECT 158.000 270.300 158.800 270.400 ;
        RECT 153.200 269.700 158.800 270.300 ;
        RECT 153.200 268.800 154.000 269.700 ;
        RECT 143.600 268.300 144.400 268.400 ;
        RECT 135.600 268.200 144.400 268.300 ;
        RECT 135.600 267.700 145.200 268.200 ;
        RECT 129.400 266.200 133.000 266.600 ;
        RECT 135.600 266.200 136.400 267.700 ;
        RECT 143.600 267.600 145.200 267.700 ;
        RECT 146.600 267.600 149.200 268.400 ;
        RECT 150.000 267.600 152.600 268.400 ;
        RECT 154.800 268.200 155.600 268.400 ;
        RECT 154.000 267.600 155.600 268.200 ;
        RECT 144.400 267.200 145.200 267.600 ;
        RECT 143.800 266.200 147.400 266.600 ;
        RECT 148.400 266.200 149.000 267.600 ;
        RECT 150.200 266.200 150.800 267.600 ;
        RECT 154.000 267.200 154.800 267.600 ;
        RECT 151.800 266.200 155.400 266.600 ;
        RECT 127.600 262.200 128.400 266.200 ;
        RECT 129.200 266.000 133.200 266.200 ;
        RECT 129.200 262.200 130.000 266.000 ;
        RECT 132.400 262.200 133.200 266.000 ;
        RECT 135.600 265.600 137.400 266.200 ;
        RECT 136.600 262.200 137.400 265.600 ;
        RECT 143.600 266.000 147.600 266.200 ;
        RECT 143.600 262.200 144.400 266.000 ;
        RECT 146.800 262.200 147.600 266.000 ;
        RECT 148.400 262.200 149.200 266.200 ;
        RECT 150.000 262.200 150.800 266.200 ;
        RECT 151.600 266.000 155.600 266.200 ;
        RECT 151.600 262.200 152.400 266.000 ;
        RECT 154.800 262.200 155.600 266.000 ;
        RECT 156.400 262.200 157.200 269.700 ;
        RECT 158.000 269.600 158.800 269.700 ;
        RECT 159.600 267.600 160.400 269.200 ;
        RECT 161.200 268.800 162.000 270.400 ;
        RECT 162.800 269.600 163.600 270.400 ;
        RECT 163.000 268.400 163.600 269.600 ;
        RECT 164.400 270.300 165.200 270.400 ;
        RECT 164.400 269.700 168.300 270.300 ;
        RECT 164.400 268.800 165.200 269.700 ;
        RECT 167.700 268.400 168.300 269.700 ;
        RECT 169.200 268.800 170.000 270.400 ;
        RECT 170.600 270.300 171.200 271.800 ;
        RECT 172.400 271.600 173.200 271.800 ;
        RECT 174.000 271.600 174.800 273.200 ;
        RECT 174.100 270.300 174.700 271.600 ;
        RECT 170.600 269.700 174.700 270.300 ;
        RECT 170.600 268.400 171.200 269.700 ;
        RECT 162.800 268.200 163.600 268.400 ;
        RECT 166.000 268.200 166.800 268.400 ;
        RECT 161.200 267.600 163.600 268.200 ;
        RECT 165.200 267.600 166.800 268.200 ;
        RECT 167.600 268.200 168.400 268.400 ;
        RECT 167.600 267.600 169.200 268.200 ;
        RECT 170.600 267.600 173.200 268.400 ;
        RECT 158.000 264.800 158.800 266.400 ;
        RECT 161.200 266.200 161.800 267.600 ;
        RECT 165.200 267.200 166.000 267.600 ;
        RECT 168.400 267.200 169.200 267.600 ;
        RECT 163.000 266.200 166.600 266.600 ;
        RECT 167.800 266.200 171.400 266.600 ;
        RECT 172.400 266.200 173.000 267.600 ;
        RECT 175.600 266.200 176.400 279.800 ;
        RECT 178.800 271.200 179.600 279.800 ;
        RECT 183.000 275.800 184.200 279.800 ;
        RECT 187.600 275.800 188.400 279.800 ;
        RECT 192.000 276.400 192.800 279.800 ;
        RECT 192.000 275.800 194.000 276.400 ;
        RECT 183.600 275.000 184.400 275.800 ;
        RECT 187.800 275.200 188.400 275.800 ;
        RECT 187.000 274.600 190.600 275.200 ;
        RECT 193.200 275.000 194.000 275.800 ;
        RECT 187.000 274.400 187.800 274.600 ;
        RECT 189.800 274.400 190.600 274.600 ;
        RECT 182.800 273.200 184.200 274.000 ;
        RECT 183.600 272.200 184.200 273.200 ;
        RECT 185.800 273.000 188.000 273.600 ;
        RECT 185.800 272.800 186.600 273.000 ;
        RECT 183.600 271.600 186.000 272.200 ;
        RECT 178.800 270.600 183.000 271.200 ;
        RECT 177.200 266.800 178.000 268.400 ;
        RECT 178.800 267.200 179.600 270.600 ;
        RECT 182.200 270.400 183.000 270.600 ;
        RECT 185.400 270.300 186.000 271.600 ;
        RECT 187.400 271.800 188.000 273.000 ;
        RECT 188.600 273.000 189.400 273.200 ;
        RECT 193.200 273.000 194.000 273.200 ;
        RECT 188.600 272.400 194.000 273.000 ;
        RECT 187.400 271.400 192.200 271.800 ;
        RECT 196.400 271.400 197.200 279.800 ;
        RECT 187.400 271.200 197.200 271.400 ;
        RECT 191.400 271.000 197.200 271.200 ;
        RECT 191.600 270.800 197.200 271.000 ;
        RECT 198.000 271.200 198.800 279.800 ;
        RECT 202.200 275.800 203.400 279.800 ;
        RECT 206.800 275.800 207.600 279.800 ;
        RECT 211.200 276.400 212.000 279.800 ;
        RECT 211.200 275.800 213.200 276.400 ;
        RECT 202.800 275.000 203.600 275.800 ;
        RECT 207.000 275.200 207.600 275.800 ;
        RECT 206.200 274.600 209.800 275.200 ;
        RECT 212.400 275.000 213.200 275.800 ;
        RECT 206.200 274.400 207.000 274.600 ;
        RECT 209.000 274.400 209.800 274.600 ;
        RECT 202.000 273.200 203.400 274.000 ;
        RECT 202.800 272.200 203.400 273.200 ;
        RECT 205.000 273.000 207.200 273.600 ;
        RECT 205.000 272.800 205.800 273.000 ;
        RECT 202.800 271.600 205.200 272.200 ;
        RECT 198.000 270.600 202.200 271.200 ;
        RECT 186.800 270.300 187.600 270.400 ;
        RECT 180.600 269.800 181.400 270.000 ;
        RECT 180.600 269.200 184.400 269.800 ;
        RECT 185.300 269.700 187.600 270.300 ;
        RECT 183.600 269.000 184.400 269.200 ;
        RECT 185.400 268.400 186.000 269.700 ;
        RECT 186.800 269.600 187.600 269.700 ;
        RECT 190.000 270.200 190.800 270.400 ;
        RECT 190.000 269.600 195.000 270.200 ;
        RECT 191.600 269.400 192.400 269.600 ;
        RECT 194.200 269.400 195.000 269.600 ;
        RECT 192.600 268.400 193.400 268.600 ;
        RECT 185.200 267.800 196.400 268.400 ;
        RECT 185.200 267.600 186.600 267.800 ;
        RECT 159.600 262.800 160.400 266.200 ;
        RECT 161.200 263.400 162.000 266.200 ;
        RECT 162.800 266.000 166.800 266.200 ;
        RECT 162.800 262.800 163.600 266.000 ;
        RECT 159.600 262.200 163.600 262.800 ;
        RECT 166.000 262.200 166.800 266.000 ;
        RECT 167.600 266.000 171.600 266.200 ;
        RECT 167.600 262.200 168.400 266.000 ;
        RECT 170.800 262.200 171.600 266.000 ;
        RECT 172.400 262.200 173.200 266.200 ;
        RECT 174.600 265.600 176.400 266.200 ;
        RECT 178.800 266.600 182.600 267.200 ;
        RECT 174.600 264.400 175.400 265.600 ;
        RECT 174.000 263.600 175.400 264.400 ;
        RECT 174.600 262.200 175.400 263.600 ;
        RECT 178.800 262.200 179.600 266.600 ;
        RECT 181.800 266.400 182.600 266.600 ;
        RECT 191.600 265.600 192.200 267.800 ;
        RECT 194.800 267.600 196.400 267.800 ;
        RECT 198.000 267.200 198.800 270.600 ;
        RECT 201.400 270.400 202.200 270.600 ;
        RECT 204.600 270.300 205.200 271.600 ;
        RECT 206.600 271.800 207.200 273.000 ;
        RECT 207.800 273.000 208.600 273.200 ;
        RECT 212.400 273.000 213.200 273.200 ;
        RECT 207.800 272.400 213.200 273.000 ;
        RECT 206.600 271.400 211.400 271.800 ;
        RECT 215.600 271.400 216.400 279.800 ;
        RECT 217.200 272.400 218.000 279.800 ;
        RECT 221.600 274.400 223.200 279.800 ;
        RECT 220.400 273.600 223.200 274.400 ;
        RECT 218.600 272.400 219.400 272.600 ;
        RECT 217.200 271.800 219.400 272.400 ;
        RECT 221.600 272.400 223.200 273.600 ;
        RECT 225.200 272.400 226.000 272.600 ;
        RECT 226.800 272.400 227.600 279.800 ;
        RECT 221.600 271.800 223.600 272.400 ;
        RECT 225.200 271.800 227.600 272.400 ;
        RECT 228.400 272.400 229.200 279.800 ;
        RECT 231.600 272.400 232.400 279.800 ;
        RECT 228.400 271.800 232.400 272.400 ;
        RECT 233.200 271.800 234.000 279.800 ;
        RECT 237.400 272.600 238.200 279.800 ;
        RECT 236.400 271.800 238.200 272.600 ;
        RECT 240.400 273.600 241.200 274.400 ;
        RECT 240.400 272.400 241.000 273.600 ;
        RECT 241.800 272.400 242.600 279.800 ;
        RECT 246.800 273.600 247.600 274.400 ;
        RECT 246.800 272.400 247.400 273.600 ;
        RECT 248.200 272.400 249.000 279.800 ;
        RECT 239.600 271.800 241.000 272.400 ;
        RECT 241.600 271.800 242.600 272.400 ;
        RECT 246.000 271.800 247.400 272.400 ;
        RECT 248.000 271.800 249.000 272.400 ;
        RECT 252.400 271.800 253.200 279.800 ;
        RECT 255.600 275.800 256.400 279.800 ;
        RECT 206.600 271.200 216.400 271.400 ;
        RECT 210.600 271.000 216.400 271.200 ;
        RECT 210.800 270.800 216.400 271.000 ;
        RECT 218.800 271.200 219.400 271.800 ;
        RECT 218.800 270.600 222.200 271.200 ;
        RECT 221.400 270.400 222.200 270.600 ;
        RECT 223.000 270.400 223.600 271.800 ;
        RECT 229.200 270.400 230.000 270.800 ;
        RECT 233.200 270.400 233.800 271.800 ;
        RECT 206.000 270.300 206.800 270.400 ;
        RECT 199.800 269.800 200.600 270.000 ;
        RECT 199.800 269.200 203.600 269.800 ;
        RECT 204.500 269.700 206.800 270.300 ;
        RECT 202.800 269.000 203.600 269.200 ;
        RECT 204.600 268.400 205.200 269.700 ;
        RECT 206.000 269.600 206.800 269.700 ;
        RECT 209.200 270.200 210.000 270.400 ;
        RECT 209.200 269.600 214.200 270.200 ;
        RECT 210.800 269.400 211.600 269.600 ;
        RECT 213.400 269.400 214.200 269.600 ;
        RECT 219.200 269.800 220.000 270.000 ;
        RECT 223.000 269.800 224.400 270.400 ;
        RECT 219.200 269.200 221.800 269.800 ;
        RECT 221.200 268.600 221.800 269.200 ;
        RECT 222.600 269.600 224.400 269.800 ;
        RECT 228.400 269.800 230.000 270.400 ;
        RECT 231.600 269.800 234.000 270.400 ;
        RECT 228.400 269.600 229.200 269.800 ;
        RECT 222.600 269.200 223.600 269.600 ;
        RECT 211.800 268.400 212.600 268.600 ;
        RECT 204.600 267.800 215.600 268.400 ;
        RECT 205.000 267.600 205.800 267.800 ;
        RECT 189.800 265.400 190.600 265.600 ;
        RECT 183.600 264.200 184.400 265.000 ;
        RECT 187.800 264.800 190.600 265.400 ;
        RECT 191.600 264.800 192.400 265.600 ;
        RECT 187.800 264.200 188.400 264.800 ;
        RECT 193.200 264.200 194.000 265.000 ;
        RECT 183.000 263.600 184.400 264.200 ;
        RECT 183.000 262.200 184.200 263.600 ;
        RECT 187.600 262.200 188.400 264.200 ;
        RECT 192.000 263.600 194.000 264.200 ;
        RECT 192.000 262.200 192.800 263.600 ;
        RECT 196.400 262.200 197.200 267.000 ;
        RECT 198.000 266.600 201.800 267.200 ;
        RECT 198.000 262.200 198.800 266.600 ;
        RECT 201.000 266.400 201.800 266.600 ;
        RECT 210.800 265.600 211.400 267.800 ;
        RECT 214.000 267.600 215.600 267.800 ;
        RECT 217.200 268.200 218.800 268.400 ;
        RECT 217.200 267.600 220.600 268.200 ;
        RECT 221.200 267.800 222.000 268.600 ;
        RECT 220.000 267.200 220.600 267.600 ;
        RECT 209.000 265.400 209.800 265.600 ;
        RECT 202.800 264.200 203.600 265.000 ;
        RECT 207.000 264.800 209.800 265.400 ;
        RECT 210.800 264.800 211.600 265.600 ;
        RECT 207.000 264.200 207.600 264.800 ;
        RECT 212.400 264.200 213.200 265.000 ;
        RECT 202.200 263.600 203.600 264.200 ;
        RECT 202.200 262.200 203.400 263.600 ;
        RECT 206.800 262.200 207.600 264.200 ;
        RECT 211.200 263.600 213.200 264.200 ;
        RECT 211.200 262.200 212.000 263.600 ;
        RECT 215.600 262.200 216.400 267.000 ;
        RECT 218.600 266.800 219.400 267.000 ;
        RECT 217.200 266.200 219.400 266.800 ;
        RECT 220.000 266.600 222.000 267.200 ;
        RECT 220.400 266.400 222.000 266.600 ;
        RECT 217.200 262.200 218.000 266.200 ;
        RECT 222.600 265.800 223.200 269.200 ;
        RECT 224.000 267.600 224.800 268.400 ;
        RECT 226.000 268.300 227.600 268.400 ;
        RECT 228.500 268.300 229.100 269.600 ;
        RECT 226.000 267.700 229.100 268.300 ;
        RECT 226.000 267.600 227.600 267.700 ;
        RECT 230.000 267.600 230.800 269.200 ;
        RECT 224.000 267.200 224.600 267.600 ;
        RECT 223.800 266.400 224.600 267.200 ;
        RECT 225.200 266.800 226.000 267.000 ;
        RECT 225.200 266.200 227.600 266.800 ;
        RECT 221.600 262.200 223.200 265.800 ;
        RECT 226.800 262.200 227.600 266.200 ;
        RECT 231.600 266.200 232.200 269.800 ;
        RECT 233.200 269.600 234.000 269.800 ;
        RECT 236.600 268.400 237.200 271.800 ;
        RECT 239.600 271.600 240.400 271.800 ;
        RECT 238.000 269.600 238.800 271.200 ;
        RECT 241.600 270.400 242.200 271.800 ;
        RECT 246.000 271.600 246.800 271.800 ;
        RECT 241.200 269.600 242.200 270.400 ;
        RECT 241.600 268.400 242.200 269.600 ;
        RECT 242.800 268.800 243.600 270.400 ;
        RECT 246.100 270.300 246.700 271.600 ;
        RECT 244.500 269.700 246.700 270.300 ;
        RECT 244.500 268.400 245.100 269.700 ;
        RECT 248.000 268.400 248.600 271.800 ;
        RECT 252.400 270.400 253.000 271.800 ;
        RECT 255.600 271.600 256.200 275.800 ;
        RECT 260.400 274.300 261.200 279.800 ;
        RECT 262.000 274.300 262.800 274.400 ;
        RECT 260.400 273.700 262.800 274.300 ;
        RECT 258.800 271.600 259.600 273.200 ;
        RECT 253.800 271.000 256.200 271.600 ;
        RECT 249.200 268.800 250.000 270.400 ;
        RECT 250.800 270.300 251.600 270.400 ;
        RECT 252.400 270.300 253.200 270.400 ;
        RECT 250.800 269.700 253.200 270.300 ;
        RECT 250.800 269.600 251.600 269.700 ;
        RECT 252.400 269.600 253.200 269.700 ;
        RECT 236.400 268.300 237.200 268.400 ;
        RECT 233.300 267.700 237.200 268.300 ;
        RECT 233.300 266.400 233.900 267.700 ;
        RECT 236.400 267.600 237.200 267.700 ;
        RECT 239.600 267.600 242.200 268.400 ;
        RECT 244.400 268.200 245.200 268.400 ;
        RECT 243.600 267.600 245.200 268.200 ;
        RECT 246.000 267.600 248.600 268.400 ;
        RECT 250.800 268.200 251.600 268.400 ;
        RECT 250.000 267.600 251.600 268.200 ;
        RECT 231.600 262.200 232.400 266.200 ;
        RECT 233.200 265.600 234.000 266.400 ;
        RECT 233.000 264.800 233.800 265.600 ;
        RECT 234.800 264.800 235.600 266.400 ;
        RECT 236.600 264.200 237.200 267.600 ;
        RECT 239.800 266.200 240.400 267.600 ;
        RECT 243.600 267.200 244.400 267.600 ;
        RECT 241.400 266.200 245.000 266.600 ;
        RECT 246.200 266.200 246.800 267.600 ;
        RECT 250.000 267.200 250.800 267.600 ;
        RECT 247.800 266.200 251.400 266.600 ;
        RECT 252.400 266.200 253.000 269.600 ;
        RECT 253.800 267.600 254.400 271.000 ;
        RECT 255.600 269.600 256.400 270.400 ;
        RECT 255.600 268.800 256.200 269.600 ;
        RECT 255.200 268.000 256.400 268.800 ;
        RECT 257.200 267.600 258.000 269.200 ;
        RECT 253.600 267.400 254.400 267.600 ;
        RECT 253.600 267.000 256.600 267.400 ;
        RECT 253.600 266.800 257.800 267.000 ;
        RECT 256.000 266.400 257.800 266.800 ;
        RECT 257.200 266.200 257.800 266.400 ;
        RECT 260.400 266.200 261.200 273.700 ;
        RECT 262.000 273.600 262.800 273.700 ;
        RECT 266.200 272.400 267.000 279.800 ;
        RECT 267.600 273.600 268.400 274.400 ;
        RECT 267.800 272.400 268.400 273.600 ;
        RECT 270.000 272.400 270.800 279.800 ;
        RECT 271.400 272.400 272.200 272.600 ;
        RECT 266.200 271.800 267.200 272.400 ;
        RECT 267.800 271.800 269.200 272.400 ;
        RECT 270.000 271.800 272.200 272.400 ;
        RECT 274.400 272.400 276.000 279.800 ;
        RECT 278.000 272.400 278.800 272.600 ;
        RECT 279.600 272.400 280.400 279.800 ;
        RECT 274.400 271.800 276.400 272.400 ;
        RECT 278.000 271.800 280.400 272.400 ;
        RECT 265.200 268.800 266.000 270.400 ;
        RECT 266.600 268.400 267.200 271.800 ;
        RECT 268.400 271.600 269.200 271.800 ;
        RECT 271.600 271.200 272.200 271.800 ;
        RECT 271.600 270.600 275.000 271.200 ;
        RECT 274.200 270.400 275.000 270.600 ;
        RECT 275.800 270.400 276.400 271.800 ;
        RECT 272.000 269.800 272.800 270.000 ;
        RECT 275.800 269.800 277.200 270.400 ;
        RECT 272.000 269.200 274.600 269.800 ;
        RECT 274.000 268.600 274.600 269.200 ;
        RECT 275.400 269.600 277.200 269.800 ;
        RECT 275.400 269.200 276.400 269.600 ;
        RECT 262.000 268.300 262.800 268.400 ;
        RECT 263.600 268.300 264.400 268.400 ;
        RECT 262.000 268.200 264.400 268.300 ;
        RECT 266.600 268.300 269.200 268.400 ;
        RECT 270.000 268.300 271.600 268.400 ;
        RECT 266.600 268.200 271.600 268.300 ;
        RECT 262.000 267.700 265.200 268.200 ;
        RECT 262.000 266.800 262.800 267.700 ;
        RECT 263.600 267.600 265.200 267.700 ;
        RECT 266.600 267.700 273.400 268.200 ;
        RECT 274.000 267.800 274.800 268.600 ;
        RECT 266.600 267.600 269.200 267.700 ;
        RECT 270.000 267.600 273.400 267.700 ;
        RECT 264.400 267.200 265.200 267.600 ;
        RECT 263.800 266.200 267.400 266.600 ;
        RECT 268.400 266.200 269.000 267.600 ;
        RECT 272.800 267.200 273.400 267.600 ;
        RECT 271.400 266.800 272.200 267.000 ;
        RECT 270.000 266.200 272.200 266.800 ;
        RECT 272.800 266.600 274.800 267.200 ;
        RECT 273.200 266.400 274.800 266.600 ;
        RECT 236.400 262.200 237.200 264.200 ;
        RECT 239.600 262.200 240.400 266.200 ;
        RECT 241.200 266.000 245.200 266.200 ;
        RECT 241.200 262.200 242.000 266.000 ;
        RECT 244.400 262.200 245.200 266.000 ;
        RECT 246.000 262.200 246.800 266.200 ;
        RECT 247.600 266.000 251.600 266.200 ;
        RECT 247.600 262.200 248.400 266.000 ;
        RECT 250.800 262.200 251.600 266.000 ;
        RECT 252.400 265.200 253.800 266.200 ;
        RECT 253.000 262.200 253.800 265.200 ;
        RECT 257.200 262.200 258.000 266.200 ;
        RECT 259.400 265.600 261.200 266.200 ;
        RECT 263.600 266.000 267.600 266.200 ;
        RECT 259.400 262.200 260.200 265.600 ;
        RECT 263.600 262.200 264.400 266.000 ;
        RECT 266.800 262.200 267.600 266.000 ;
        RECT 268.400 262.200 269.200 266.200 ;
        RECT 270.000 262.200 270.800 266.200 ;
        RECT 275.400 265.800 276.000 269.200 ;
        RECT 276.800 267.600 277.600 268.400 ;
        RECT 278.800 267.600 280.400 268.400 ;
        RECT 276.800 267.200 277.400 267.600 ;
        RECT 276.600 266.400 277.400 267.200 ;
        RECT 278.000 266.800 278.800 267.000 ;
        RECT 278.000 266.200 280.400 266.800 ;
        RECT 274.400 264.400 276.000 265.800 ;
        RECT 273.200 263.600 276.000 264.400 ;
        RECT 274.400 262.200 276.000 263.600 ;
        RECT 279.600 262.200 280.400 266.200 ;
        RECT 281.200 262.200 282.000 279.800 ;
        RECT 284.400 272.400 285.200 279.800 ;
        RECT 285.800 272.400 286.600 272.600 ;
        RECT 284.400 271.800 286.600 272.400 ;
        RECT 288.800 272.400 290.400 279.800 ;
        RECT 292.400 272.400 293.200 272.600 ;
        RECT 294.000 272.400 294.800 279.800 ;
        RECT 288.800 271.800 290.800 272.400 ;
        RECT 292.400 271.800 294.800 272.400 ;
        RECT 301.000 272.600 301.800 279.800 ;
        RECT 307.800 272.600 308.600 279.800 ;
        RECT 301.000 271.800 302.800 272.600 ;
        RECT 306.800 271.800 308.600 272.600 ;
        RECT 286.000 271.200 286.600 271.800 ;
        RECT 286.000 270.600 289.400 271.200 ;
        RECT 288.600 270.400 289.400 270.600 ;
        RECT 290.200 270.400 290.800 271.800 ;
        RECT 286.400 269.800 287.200 270.000 ;
        RECT 290.200 269.800 291.600 270.400 ;
        RECT 286.400 269.200 289.000 269.800 ;
        RECT 288.400 268.600 289.000 269.200 ;
        RECT 289.800 269.600 291.600 269.800 ;
        RECT 300.400 269.600 301.200 271.200 ;
        RECT 289.800 269.200 290.800 269.600 ;
        RECT 284.400 268.200 286.000 268.400 ;
        RECT 284.400 267.600 287.800 268.200 ;
        RECT 288.400 267.800 289.200 268.600 ;
        RECT 287.200 267.200 287.800 267.600 ;
        RECT 285.800 266.800 286.600 267.000 ;
        RECT 282.800 264.800 283.600 266.400 ;
        RECT 284.400 266.200 286.600 266.800 ;
        RECT 287.200 266.600 289.200 267.200 ;
        RECT 287.600 266.400 289.200 266.600 ;
        RECT 284.400 262.200 285.200 266.200 ;
        RECT 289.800 265.800 290.400 269.200 ;
        RECT 302.000 268.400 302.600 271.800 ;
        RECT 303.600 270.300 304.400 270.400 ;
        RECT 307.000 270.300 307.600 271.800 ;
        RECT 303.600 269.700 307.600 270.300 ;
        RECT 303.600 269.600 304.400 269.700 ;
        RECT 307.000 268.400 307.600 269.700 ;
        RECT 308.400 269.600 309.200 271.200 ;
        RECT 291.200 267.600 292.000 268.400 ;
        RECT 293.200 267.600 294.800 268.400 ;
        RECT 295.600 268.300 296.400 268.400 ;
        RECT 302.000 268.300 302.800 268.400 ;
        RECT 305.200 268.300 306.000 268.400 ;
        RECT 295.600 267.700 302.800 268.300 ;
        RECT 295.600 267.600 296.400 267.700 ;
        RECT 302.000 267.600 302.800 267.700 ;
        RECT 303.700 267.700 306.000 268.300 ;
        RECT 291.200 267.200 291.800 267.600 ;
        RECT 291.000 266.400 291.800 267.200 ;
        RECT 292.400 266.800 293.200 267.000 ;
        RECT 292.400 266.200 294.800 266.800 ;
        RECT 288.800 264.400 290.400 265.800 ;
        RECT 287.600 263.600 290.400 264.400 ;
        RECT 288.800 262.200 290.400 263.600 ;
        RECT 294.000 262.200 294.800 266.200 ;
        RECT 302.000 264.200 302.600 267.600 ;
        RECT 303.700 266.400 304.300 267.700 ;
        RECT 305.200 267.600 306.000 267.700 ;
        RECT 306.800 267.600 307.600 268.400 ;
        RECT 308.400 268.300 309.200 268.400 ;
        RECT 310.000 268.300 310.800 279.800 ;
        RECT 314.000 273.600 314.800 274.400 ;
        RECT 314.000 272.400 314.600 273.600 ;
        RECT 315.400 272.400 316.200 279.800 ;
        RECT 313.200 271.800 314.600 272.400 ;
        RECT 315.200 271.800 316.200 272.400 ;
        RECT 322.200 271.800 324.200 279.800 ;
        RECT 313.200 271.600 314.000 271.800 ;
        RECT 311.600 270.300 312.400 270.400 ;
        RECT 315.200 270.300 315.800 271.800 ;
        RECT 311.600 269.700 315.800 270.300 ;
        RECT 311.600 269.600 312.400 269.700 ;
        RECT 315.200 268.400 315.800 269.700 ;
        RECT 316.400 268.800 317.200 270.400 ;
        RECT 308.400 267.700 310.800 268.300 ;
        RECT 308.400 267.600 309.200 267.700 ;
        RECT 303.600 264.800 304.400 266.400 ;
        RECT 305.200 264.800 306.000 266.400 ;
        RECT 307.000 264.200 307.600 267.600 ;
        RECT 302.000 262.200 302.800 264.200 ;
        RECT 306.800 262.200 307.600 264.200 ;
        RECT 310.000 262.200 310.800 267.700 ;
        RECT 313.200 267.600 315.800 268.400 ;
        RECT 318.000 268.200 318.800 268.400 ;
        RECT 317.200 267.600 318.800 268.200 ;
        RECT 319.600 267.600 320.400 269.200 ;
        RECT 321.200 268.800 322.000 270.400 ;
        RECT 323.000 268.400 323.600 271.800 ;
        RECT 324.400 268.800 325.200 270.400 ;
        RECT 322.800 268.200 323.600 268.400 ;
        RECT 326.000 268.300 326.800 268.400 ;
        RECT 327.600 268.300 328.400 279.800 ;
        RECT 330.800 271.600 331.600 273.200 ;
        RECT 326.000 268.200 328.400 268.300 ;
        RECT 321.200 267.600 323.600 268.200 ;
        RECT 325.200 267.700 328.400 268.200 ;
        RECT 325.200 267.600 326.800 267.700 ;
        RECT 311.600 264.800 312.400 266.400 ;
        RECT 313.400 266.200 314.000 267.600 ;
        RECT 317.200 267.200 318.000 267.600 ;
        RECT 315.000 266.200 318.600 266.600 ;
        RECT 321.200 266.400 321.800 267.600 ;
        RECT 325.200 267.200 326.000 267.600 ;
        RECT 313.200 262.200 314.000 266.200 ;
        RECT 314.800 266.000 318.800 266.200 ;
        RECT 314.800 262.200 315.600 266.000 ;
        RECT 318.000 262.200 318.800 266.000 ;
        RECT 319.600 262.800 320.400 266.200 ;
        RECT 321.200 263.400 322.000 266.400 ;
        RECT 323.000 266.200 326.600 266.600 ;
        RECT 322.800 266.000 326.800 266.200 ;
        RECT 322.800 262.800 323.600 266.000 ;
        RECT 319.600 262.200 323.600 262.800 ;
        RECT 326.000 262.200 326.800 266.000 ;
        RECT 327.600 262.200 328.400 267.700 ;
        RECT 329.200 264.800 330.000 266.400 ;
        RECT 332.400 266.200 333.200 279.800 ;
        RECT 336.200 272.400 337.000 279.800 ;
        RECT 335.600 271.800 337.000 272.400 ;
        RECT 335.600 270.400 336.200 271.800 ;
        RECT 340.400 271.200 341.200 279.800 ;
        RECT 337.200 270.800 341.200 271.200 ;
        RECT 337.000 270.600 341.200 270.800 ;
        RECT 342.000 271.200 342.800 279.800 ;
        RECT 346.200 275.800 347.400 279.800 ;
        RECT 350.800 275.800 351.600 279.800 ;
        RECT 355.200 276.400 356.000 279.800 ;
        RECT 355.200 275.800 357.200 276.400 ;
        RECT 346.800 275.000 347.600 275.800 ;
        RECT 351.000 275.200 351.600 275.800 ;
        RECT 350.200 274.600 353.800 275.200 ;
        RECT 356.400 275.000 357.200 275.800 ;
        RECT 350.200 274.400 351.000 274.600 ;
        RECT 353.000 274.400 353.800 274.600 ;
        RECT 346.000 273.200 347.400 274.000 ;
        RECT 346.800 272.200 347.400 273.200 ;
        RECT 349.000 273.000 351.200 273.600 ;
        RECT 349.000 272.800 349.800 273.000 ;
        RECT 346.800 271.600 349.200 272.200 ;
        RECT 342.000 270.600 346.200 271.200 ;
        RECT 334.000 270.300 334.800 270.400 ;
        RECT 335.600 270.300 336.400 270.400 ;
        RECT 334.000 269.700 336.400 270.300 ;
        RECT 334.000 269.600 334.800 269.700 ;
        RECT 335.600 269.600 336.400 269.700 ;
        RECT 337.000 270.000 337.800 270.600 ;
        RECT 334.000 266.800 334.800 268.400 ;
        RECT 331.400 265.600 333.200 266.200 ;
        RECT 335.600 266.200 336.200 269.600 ;
        RECT 337.000 267.000 337.600 270.000 ;
        RECT 338.400 268.400 339.200 269.200 ;
        RECT 338.600 267.600 339.600 268.400 ;
        RECT 342.000 267.200 342.800 270.600 ;
        RECT 345.400 270.400 346.200 270.600 ;
        RECT 343.800 269.800 344.600 270.000 ;
        RECT 343.800 269.200 347.600 269.800 ;
        RECT 346.800 269.000 347.600 269.200 ;
        RECT 348.600 268.400 349.200 271.600 ;
        RECT 350.600 271.800 351.200 273.000 ;
        RECT 351.800 273.000 352.600 273.200 ;
        RECT 356.400 273.000 357.200 273.200 ;
        RECT 351.800 272.400 357.200 273.000 ;
        RECT 350.600 271.400 355.400 271.800 ;
        RECT 359.600 271.400 360.400 279.800 ;
        RECT 361.200 272.400 362.000 279.800 ;
        RECT 365.600 274.400 367.200 279.800 ;
        RECT 364.400 273.600 367.200 274.400 ;
        RECT 362.600 272.400 363.400 272.600 ;
        RECT 361.200 271.800 363.400 272.400 ;
        RECT 365.600 272.400 367.200 273.600 ;
        RECT 369.200 272.400 370.000 272.600 ;
        RECT 370.800 272.400 371.600 279.800 ;
        RECT 373.200 273.600 374.000 274.400 ;
        RECT 373.200 272.400 373.800 273.600 ;
        RECT 374.600 272.400 375.400 279.800 ;
        RECT 365.600 271.800 367.600 272.400 ;
        RECT 369.200 271.800 371.600 272.400 ;
        RECT 372.400 271.800 373.800 272.400 ;
        RECT 374.400 271.800 375.400 272.400 ;
        RECT 350.600 271.200 360.400 271.400 ;
        RECT 354.600 271.000 360.400 271.200 ;
        RECT 354.800 270.800 360.400 271.000 ;
        RECT 362.800 271.200 363.400 271.800 ;
        RECT 362.800 270.600 366.200 271.200 ;
        RECT 365.400 270.400 366.200 270.600 ;
        RECT 367.000 270.400 367.600 271.800 ;
        RECT 372.400 271.600 373.200 271.800 ;
        RECT 353.200 270.200 354.000 270.400 ;
        RECT 353.200 269.600 358.200 270.200 ;
        RECT 354.800 269.400 355.600 269.600 ;
        RECT 357.400 269.400 358.200 269.600 ;
        RECT 363.200 269.800 364.000 270.000 ;
        RECT 367.000 269.800 368.400 270.400 ;
        RECT 363.200 269.200 365.800 269.800 ;
        RECT 365.200 268.600 365.800 269.200 ;
        RECT 366.600 269.600 368.400 269.800 ;
        RECT 370.800 270.300 371.600 270.400 ;
        RECT 374.400 270.300 375.000 271.800 ;
        RECT 370.800 269.700 375.000 270.300 ;
        RECT 370.800 269.600 371.600 269.700 ;
        RECT 366.600 269.200 367.600 269.600 ;
        RECT 355.800 268.400 356.600 268.600 ;
        RECT 348.600 267.800 359.600 268.400 ;
        RECT 349.000 267.600 349.800 267.800 ;
        RECT 351.600 267.600 352.400 267.800 ;
        RECT 337.000 266.400 339.400 267.000 ;
        RECT 342.000 266.600 345.800 267.200 ;
        RECT 331.400 264.400 332.200 265.600 ;
        RECT 331.400 263.600 333.200 264.400 ;
        RECT 331.400 262.200 332.200 263.600 ;
        RECT 335.600 262.200 336.400 266.200 ;
        RECT 338.800 264.200 339.400 266.400 ;
        RECT 340.400 264.800 341.200 266.400 ;
        RECT 338.800 262.200 339.600 264.200 ;
        RECT 342.000 262.200 342.800 266.600 ;
        RECT 345.000 266.400 345.800 266.600 ;
        RECT 354.800 265.600 355.400 267.800 ;
        RECT 358.000 267.600 359.600 267.800 ;
        RECT 361.200 268.200 362.800 268.400 ;
        RECT 361.200 267.600 364.600 268.200 ;
        RECT 365.200 267.800 366.000 268.600 ;
        RECT 364.000 267.200 364.600 267.600 ;
        RECT 353.000 265.400 353.800 265.600 ;
        RECT 346.800 264.200 347.600 265.000 ;
        RECT 351.000 264.800 353.800 265.400 ;
        RECT 354.800 264.800 355.600 265.600 ;
        RECT 351.000 264.200 351.600 264.800 ;
        RECT 356.400 264.200 357.200 265.000 ;
        RECT 346.200 263.600 347.600 264.200 ;
        RECT 346.200 262.200 347.400 263.600 ;
        RECT 350.800 262.200 351.600 264.200 ;
        RECT 355.200 263.600 357.200 264.200 ;
        RECT 355.200 262.200 356.000 263.600 ;
        RECT 359.600 262.200 360.400 267.000 ;
        RECT 362.600 266.800 363.400 267.000 ;
        RECT 361.200 266.200 363.400 266.800 ;
        RECT 364.000 266.600 366.000 267.200 ;
        RECT 364.400 266.400 366.000 266.600 ;
        RECT 361.200 262.200 362.000 266.200 ;
        RECT 366.600 265.800 367.200 269.200 ;
        RECT 374.400 268.400 375.000 269.700 ;
        RECT 375.600 270.300 376.400 270.400 ;
        RECT 378.800 270.300 379.600 279.800 ;
        RECT 383.600 275.800 384.400 279.800 ;
        RECT 383.800 275.600 384.400 275.800 ;
        RECT 386.800 275.800 387.600 279.800 ;
        RECT 386.800 275.600 387.400 275.800 ;
        RECT 383.800 275.000 387.400 275.600 ;
        RECT 385.200 272.800 386.000 274.400 ;
        RECT 386.800 272.400 387.400 275.000 ;
        RECT 388.400 272.400 389.200 279.800 ;
        RECT 391.600 272.400 392.400 279.800 ;
        RECT 382.000 270.800 382.800 272.400 ;
        RECT 386.800 271.600 387.600 272.400 ;
        RECT 388.400 271.800 392.400 272.400 ;
        RECT 393.200 271.800 394.000 279.800 ;
        RECT 375.600 269.700 379.600 270.300 ;
        RECT 375.600 268.800 376.400 269.700 ;
        RECT 368.000 267.600 368.800 268.400 ;
        RECT 370.000 267.600 371.600 268.400 ;
        RECT 372.400 267.600 375.000 268.400 ;
        RECT 377.200 268.200 378.000 268.400 ;
        RECT 376.400 267.600 378.000 268.200 ;
        RECT 368.000 267.200 368.600 267.600 ;
        RECT 367.800 266.400 368.600 267.200 ;
        RECT 369.200 266.800 370.000 267.000 ;
        RECT 369.200 266.200 371.600 266.800 ;
        RECT 372.600 266.200 373.200 267.600 ;
        RECT 376.400 267.200 377.200 267.600 ;
        RECT 374.200 266.200 377.800 266.600 ;
        RECT 365.600 262.200 367.200 265.800 ;
        RECT 370.800 262.200 371.600 266.200 ;
        RECT 372.400 262.200 373.200 266.200 ;
        RECT 374.000 266.000 378.000 266.200 ;
        RECT 374.000 262.200 374.800 266.000 ;
        RECT 377.200 262.200 378.000 266.000 ;
        RECT 378.800 262.200 379.600 269.700 ;
        RECT 383.600 269.600 385.200 270.400 ;
        RECT 386.800 268.400 387.400 271.600 ;
        RECT 389.200 270.400 390.000 270.800 ;
        RECT 393.200 270.400 393.800 271.800 ;
        RECT 388.400 269.800 390.000 270.400 ;
        RECT 391.600 269.800 394.000 270.400 ;
        RECT 388.400 269.600 389.200 269.800 ;
        RECT 385.800 268.200 387.400 268.400 ;
        RECT 385.600 267.800 387.400 268.200 ;
        RECT 380.400 264.800 381.200 266.400 ;
        RECT 385.600 262.200 386.400 267.800 ;
        RECT 390.000 267.600 390.800 269.200 ;
        RECT 391.600 266.200 392.200 269.800 ;
        RECT 393.200 269.600 394.000 269.800 ;
        RECT 391.600 262.200 392.400 266.200 ;
        RECT 393.200 265.600 394.000 266.400 ;
        RECT 393.000 264.800 393.800 265.600 ;
        RECT 394.800 262.200 395.600 279.800 ;
        RECT 398.000 271.600 398.800 273.200 ;
        RECT 396.400 264.800 397.200 266.400 ;
        RECT 399.600 266.200 400.400 279.800 ;
        RECT 405.400 272.600 406.200 279.800 ;
        RECT 404.400 271.800 406.200 272.600 ;
        RECT 404.400 271.600 405.200 271.800 ;
        RECT 404.600 268.400 405.200 271.600 ;
        RECT 406.000 269.600 406.800 271.200 ;
        RECT 401.200 268.300 402.000 268.400 ;
        RECT 402.800 268.300 403.600 268.400 ;
        RECT 401.200 267.700 403.600 268.300 ;
        RECT 401.200 266.800 402.000 267.700 ;
        RECT 402.800 267.600 403.600 267.700 ;
        RECT 404.400 267.600 405.200 268.400 ;
        RECT 398.600 265.600 400.400 266.200 ;
        RECT 398.600 264.400 399.400 265.600 ;
        RECT 402.800 264.800 403.600 266.400 ;
        RECT 398.000 263.600 399.400 264.400 ;
        RECT 404.600 264.200 405.200 267.600 ;
        RECT 406.000 266.300 406.800 266.400 ;
        RECT 407.600 266.300 408.400 266.400 ;
        RECT 406.000 265.700 408.400 266.300 ;
        RECT 406.000 265.600 406.800 265.700 ;
        RECT 407.600 264.800 408.400 265.700 ;
        RECT 398.600 262.200 399.400 263.600 ;
        RECT 404.400 262.200 405.200 264.200 ;
        RECT 409.200 262.200 410.000 279.800 ;
        RECT 410.800 262.200 411.600 279.800 ;
        RECT 412.400 274.300 413.200 274.400 ;
        RECT 414.000 274.300 414.800 279.800 ;
        RECT 418.200 275.800 419.400 279.800 ;
        RECT 422.800 275.800 423.600 279.800 ;
        RECT 427.200 276.400 428.000 279.800 ;
        RECT 427.200 275.800 429.200 276.400 ;
        RECT 418.800 275.000 419.600 275.800 ;
        RECT 423.000 275.200 423.600 275.800 ;
        RECT 422.200 274.600 425.800 275.200 ;
        RECT 428.400 275.000 429.200 275.800 ;
        RECT 422.200 274.400 423.000 274.600 ;
        RECT 425.000 274.400 425.800 274.600 ;
        RECT 412.400 273.700 414.800 274.300 ;
        RECT 412.400 273.600 413.200 273.700 ;
        RECT 414.000 271.200 414.800 273.700 ;
        RECT 418.000 273.200 419.400 274.000 ;
        RECT 418.800 272.200 419.400 273.200 ;
        RECT 421.000 273.000 423.200 273.600 ;
        RECT 421.000 272.800 421.800 273.000 ;
        RECT 418.800 271.600 421.200 272.200 ;
        RECT 414.000 270.600 418.200 271.200 ;
        RECT 414.000 267.200 414.800 270.600 ;
        RECT 417.400 270.400 418.200 270.600 ;
        RECT 420.600 270.400 421.200 271.600 ;
        RECT 422.600 271.800 423.200 273.000 ;
        RECT 423.800 273.000 424.600 273.200 ;
        RECT 428.400 273.000 429.200 273.200 ;
        RECT 423.800 272.400 429.200 273.000 ;
        RECT 422.600 271.400 427.400 271.800 ;
        RECT 431.600 271.400 432.400 279.800 ;
        RECT 433.800 272.600 434.600 279.800 ;
        RECT 438.800 273.600 439.600 274.400 ;
        RECT 433.800 271.800 435.600 272.600 ;
        RECT 438.800 272.400 439.400 273.600 ;
        RECT 440.200 272.400 441.000 279.800 ;
        RECT 438.000 271.800 439.400 272.400 ;
        RECT 440.000 271.800 441.000 272.400 ;
        RECT 449.200 272.400 450.000 279.800 ;
        RECT 453.600 278.400 455.200 279.800 ;
        RECT 453.600 277.600 456.400 278.400 ;
        RECT 451.000 272.400 451.800 272.600 ;
        RECT 449.200 271.800 451.800 272.400 ;
        RECT 453.600 271.800 455.200 277.600 ;
        RECT 457.200 272.400 458.000 272.600 ;
        RECT 458.800 272.400 459.600 279.800 ;
        RECT 457.200 271.800 459.600 272.400 ;
        RECT 422.600 271.200 432.400 271.400 ;
        RECT 426.600 271.000 432.400 271.200 ;
        RECT 426.800 270.800 432.400 271.000 ;
        RECT 415.800 269.800 416.600 270.000 ;
        RECT 415.800 269.200 419.600 269.800 ;
        RECT 420.400 269.600 421.200 270.400 ;
        RECT 425.200 270.200 426.000 270.400 ;
        RECT 425.200 269.600 430.200 270.200 ;
        RECT 433.200 269.600 434.000 271.200 ;
        RECT 418.800 269.000 419.600 269.200 ;
        RECT 420.600 268.400 421.200 269.600 ;
        RECT 426.800 269.400 427.600 269.600 ;
        RECT 429.400 269.400 430.200 269.600 ;
        RECT 427.800 268.400 428.600 268.600 ;
        RECT 434.800 268.400 435.400 271.800 ;
        RECT 438.000 271.600 438.800 271.800 ;
        RECT 440.000 270.400 440.600 271.800 ;
        RECT 452.200 270.400 453.000 270.600 ;
        RECT 454.200 270.400 454.800 271.800 ;
        RECT 439.600 269.600 440.600 270.400 ;
        RECT 440.000 268.400 440.600 269.600 ;
        RECT 441.200 270.300 442.000 270.400 ;
        RECT 444.400 270.300 445.200 270.400 ;
        RECT 441.200 269.700 445.200 270.300 ;
        RECT 441.200 268.800 442.000 269.700 ;
        RECT 444.400 269.600 445.200 269.700 ;
        RECT 451.400 269.800 453.000 270.400 ;
        RECT 451.400 269.600 452.200 269.800 ;
        RECT 454.000 269.600 454.800 270.400 ;
        RECT 452.800 268.600 453.600 268.800 ;
        RECT 450.800 268.400 453.600 268.600 ;
        RECT 420.600 267.800 431.600 268.400 ;
        RECT 421.000 267.600 421.800 267.800 ;
        RECT 414.000 266.600 417.800 267.200 ;
        RECT 412.400 264.800 413.200 266.400 ;
        RECT 414.000 262.200 414.800 266.600 ;
        RECT 417.000 266.400 417.800 266.600 ;
        RECT 426.800 265.600 427.400 267.800 ;
        RECT 430.000 267.600 431.600 267.800 ;
        RECT 434.800 267.600 435.600 268.400 ;
        RECT 438.000 267.600 440.600 268.400 ;
        RECT 442.800 268.200 443.600 268.400 ;
        RECT 442.000 267.600 443.600 268.200 ;
        RECT 449.200 268.000 453.600 268.400 ;
        RECT 454.200 268.400 454.800 269.600 ;
        RECT 449.200 267.800 451.400 268.000 ;
        RECT 454.200 267.800 455.200 268.400 ;
        RECT 449.200 267.600 450.800 267.800 ;
        RECT 425.000 265.400 425.800 265.600 ;
        RECT 418.800 264.200 419.600 265.000 ;
        RECT 423.000 264.800 425.800 265.400 ;
        RECT 426.800 264.800 427.600 265.600 ;
        RECT 423.000 264.200 423.600 264.800 ;
        RECT 428.400 264.200 429.200 265.000 ;
        RECT 418.200 263.600 419.600 264.200 ;
        RECT 418.200 262.200 419.400 263.600 ;
        RECT 422.800 262.200 423.600 264.200 ;
        RECT 427.200 263.600 429.200 264.200 ;
        RECT 427.200 262.200 428.000 263.600 ;
        RECT 431.600 262.200 432.400 267.000 ;
        RECT 434.800 264.400 435.400 267.600 ;
        RECT 436.400 264.800 437.200 266.400 ;
        RECT 438.200 266.200 438.800 267.600 ;
        RECT 442.000 267.200 442.800 267.600 ;
        RECT 451.000 266.800 451.800 267.000 ;
        RECT 439.800 266.200 443.400 266.600 ;
        RECT 449.200 266.200 451.800 266.800 ;
        RECT 452.400 266.400 454.000 267.200 ;
        RECT 434.800 262.200 435.600 264.400 ;
        RECT 438.000 262.200 438.800 266.200 ;
        RECT 439.600 266.000 443.600 266.200 ;
        RECT 439.600 262.200 440.400 266.000 ;
        RECT 442.800 262.200 443.600 266.000 ;
        RECT 449.200 262.200 450.000 266.200 ;
        RECT 454.600 265.800 455.200 267.800 ;
        RECT 456.000 267.600 456.800 268.400 ;
        RECT 458.000 267.600 459.600 268.400 ;
        RECT 456.000 267.200 456.600 267.600 ;
        RECT 455.800 266.400 456.600 267.200 ;
        RECT 457.200 266.800 458.000 267.000 ;
        RECT 460.400 266.800 461.200 268.400 ;
        RECT 457.200 266.200 459.600 266.800 ;
        RECT 453.600 262.200 455.200 265.800 ;
        RECT 458.800 262.200 459.600 266.200 ;
        RECT 462.000 266.200 462.800 279.800 ;
        RECT 463.600 271.600 464.400 273.200 ;
        RECT 465.200 271.400 466.000 279.800 ;
        RECT 469.600 276.400 470.400 279.800 ;
        RECT 468.400 275.800 470.400 276.400 ;
        RECT 474.000 275.800 474.800 279.800 ;
        RECT 478.200 275.800 479.400 279.800 ;
        RECT 468.400 275.000 469.200 275.800 ;
        RECT 474.000 275.200 474.600 275.800 ;
        RECT 471.800 274.600 475.400 275.200 ;
        RECT 478.000 275.000 478.800 275.800 ;
        RECT 471.800 274.400 472.600 274.600 ;
        RECT 474.600 274.400 475.400 274.600 ;
        RECT 468.400 273.000 469.200 273.200 ;
        RECT 473.000 273.000 473.800 273.200 ;
        RECT 468.400 272.400 473.800 273.000 ;
        RECT 474.400 273.000 476.600 273.600 ;
        RECT 474.400 271.800 475.000 273.000 ;
        RECT 475.800 272.800 476.600 273.000 ;
        RECT 478.200 273.200 479.600 274.000 ;
        RECT 478.200 272.200 478.800 273.200 ;
        RECT 470.200 271.400 475.000 271.800 ;
        RECT 465.200 271.200 475.000 271.400 ;
        RECT 476.400 271.600 478.800 272.200 ;
        RECT 465.200 271.000 471.000 271.200 ;
        RECT 465.200 270.800 470.800 271.000 ;
        RECT 471.600 270.200 472.400 270.400 ;
        RECT 467.400 269.600 472.400 270.200 ;
        RECT 467.400 269.400 468.200 269.600 ;
        RECT 470.000 269.400 470.800 269.600 ;
        RECT 469.000 268.400 469.800 268.600 ;
        RECT 476.400 268.400 477.000 271.600 ;
        RECT 482.800 271.200 483.600 279.800 ;
        RECT 479.400 270.600 483.600 271.200 ;
        RECT 484.400 271.400 485.200 279.800 ;
        RECT 488.800 276.400 489.600 279.800 ;
        RECT 487.600 275.800 489.600 276.400 ;
        RECT 493.200 275.800 494.000 279.800 ;
        RECT 497.400 275.800 498.600 279.800 ;
        RECT 487.600 275.000 488.400 275.800 ;
        RECT 493.200 275.200 493.800 275.800 ;
        RECT 491.000 274.600 494.600 275.200 ;
        RECT 497.200 275.000 498.000 275.800 ;
        RECT 491.000 274.400 491.800 274.600 ;
        RECT 493.800 274.400 494.600 274.600 ;
        RECT 487.600 273.000 488.400 273.200 ;
        RECT 492.200 273.000 493.000 273.200 ;
        RECT 487.600 272.400 493.000 273.000 ;
        RECT 493.600 273.000 495.800 273.600 ;
        RECT 493.600 271.800 494.200 273.000 ;
        RECT 495.000 272.800 495.800 273.000 ;
        RECT 497.400 273.200 498.800 274.000 ;
        RECT 497.400 272.200 498.000 273.200 ;
        RECT 489.400 271.400 494.200 271.800 ;
        RECT 484.400 271.200 494.200 271.400 ;
        RECT 495.600 271.600 498.000 272.200 ;
        RECT 484.400 271.000 490.200 271.200 ;
        RECT 484.400 270.800 490.000 271.000 ;
        RECT 479.400 270.400 480.200 270.600 ;
        RECT 481.000 269.800 481.800 270.000 ;
        RECT 478.000 269.200 481.800 269.800 ;
        RECT 478.000 269.000 478.800 269.200 ;
        RECT 466.000 267.800 477.000 268.400 ;
        RECT 466.000 267.600 467.600 267.800 ;
        RECT 462.000 265.600 463.800 266.200 ;
        RECT 463.000 262.200 463.800 265.600 ;
        RECT 465.200 262.200 466.000 267.000 ;
        RECT 470.200 265.600 470.800 267.800 ;
        RECT 475.800 267.600 476.600 267.800 ;
        RECT 482.800 267.200 483.600 270.600 ;
        RECT 495.600 270.400 496.200 271.600 ;
        RECT 502.000 271.200 502.800 279.800 ;
        RECT 498.600 270.600 502.800 271.200 ;
        RECT 503.600 271.400 504.400 279.800 ;
        RECT 508.000 276.400 508.800 279.800 ;
        RECT 506.800 275.800 508.800 276.400 ;
        RECT 512.400 275.800 513.200 279.800 ;
        RECT 516.600 275.800 517.800 279.800 ;
        RECT 506.800 275.000 507.600 275.800 ;
        RECT 512.400 275.200 513.000 275.800 ;
        RECT 510.200 274.600 513.800 275.200 ;
        RECT 516.400 275.000 517.200 275.800 ;
        RECT 510.200 274.400 511.000 274.600 ;
        RECT 513.000 274.400 513.800 274.600 ;
        RECT 506.800 273.000 507.600 273.200 ;
        RECT 511.400 273.000 512.200 273.200 ;
        RECT 506.800 272.400 512.200 273.000 ;
        RECT 512.800 273.000 515.000 273.600 ;
        RECT 512.800 271.800 513.400 273.000 ;
        RECT 514.200 272.800 515.000 273.000 ;
        RECT 516.600 273.200 518.000 274.000 ;
        RECT 516.600 272.200 517.200 273.200 ;
        RECT 508.600 271.400 513.400 271.800 ;
        RECT 503.600 271.200 513.400 271.400 ;
        RECT 514.800 271.600 517.200 272.200 ;
        RECT 503.600 271.000 509.400 271.200 ;
        RECT 503.600 270.800 509.200 271.000 ;
        RECT 498.600 270.400 499.400 270.600 ;
        RECT 490.800 270.200 491.600 270.400 ;
        RECT 486.600 269.600 491.600 270.200 ;
        RECT 495.600 269.600 496.400 270.400 ;
        RECT 500.200 269.800 501.000 270.000 ;
        RECT 486.600 269.400 487.400 269.600 ;
        RECT 489.200 269.400 490.000 269.600 ;
        RECT 488.200 268.400 489.000 268.600 ;
        RECT 495.600 268.400 496.200 269.600 ;
        RECT 497.200 269.200 501.000 269.800 ;
        RECT 497.200 269.000 498.000 269.200 ;
        RECT 485.200 267.800 496.200 268.400 ;
        RECT 485.200 267.600 486.800 267.800 ;
        RECT 479.800 266.600 483.600 267.200 ;
        RECT 479.800 266.400 480.600 266.600 ;
        RECT 468.400 264.200 469.200 265.000 ;
        RECT 470.000 264.800 470.800 265.600 ;
        RECT 471.800 265.400 472.600 265.600 ;
        RECT 471.800 264.800 474.600 265.400 ;
        RECT 474.000 264.200 474.600 264.800 ;
        RECT 478.000 264.200 478.800 265.000 ;
        RECT 468.400 263.600 470.400 264.200 ;
        RECT 469.600 262.200 470.400 263.600 ;
        RECT 474.000 262.200 474.800 264.200 ;
        RECT 478.000 263.600 479.400 264.200 ;
        RECT 478.200 262.200 479.400 263.600 ;
        RECT 482.800 262.200 483.600 266.600 ;
        RECT 484.400 262.200 485.200 267.000 ;
        RECT 489.400 265.600 490.000 267.800 ;
        RECT 492.400 267.600 493.200 267.800 ;
        RECT 495.000 267.600 495.800 267.800 ;
        RECT 502.000 267.200 502.800 270.600 ;
        RECT 510.000 270.200 510.800 270.400 ;
        RECT 505.800 269.600 510.800 270.200 ;
        RECT 505.800 269.400 506.600 269.600 ;
        RECT 507.400 268.400 508.200 268.600 ;
        RECT 514.800 268.400 515.400 271.600 ;
        RECT 521.200 271.200 522.000 279.800 ;
        RECT 517.800 270.600 522.000 271.200 ;
        RECT 522.800 271.400 523.600 279.800 ;
        RECT 527.200 276.400 528.000 279.800 ;
        RECT 526.000 275.800 528.000 276.400 ;
        RECT 531.600 275.800 532.400 279.800 ;
        RECT 535.800 275.800 537.000 279.800 ;
        RECT 526.000 275.000 526.800 275.800 ;
        RECT 531.600 275.200 532.200 275.800 ;
        RECT 529.400 274.600 533.000 275.200 ;
        RECT 535.600 275.000 536.400 275.800 ;
        RECT 529.400 274.400 530.200 274.600 ;
        RECT 532.200 274.400 533.000 274.600 ;
        RECT 526.000 273.000 526.800 273.200 ;
        RECT 530.600 273.000 531.400 273.200 ;
        RECT 526.000 272.400 531.400 273.000 ;
        RECT 532.000 273.000 534.200 273.600 ;
        RECT 532.000 271.800 532.600 273.000 ;
        RECT 533.400 272.800 534.200 273.000 ;
        RECT 535.800 273.200 537.200 274.000 ;
        RECT 535.800 272.200 536.400 273.200 ;
        RECT 527.800 271.400 532.600 271.800 ;
        RECT 522.800 271.200 532.600 271.400 ;
        RECT 534.000 271.600 536.400 272.200 ;
        RECT 522.800 271.000 528.600 271.200 ;
        RECT 522.800 270.800 528.400 271.000 ;
        RECT 517.800 270.400 518.600 270.600 ;
        RECT 519.400 269.800 520.200 270.000 ;
        RECT 516.400 269.200 520.200 269.800 ;
        RECT 516.400 269.000 517.200 269.200 ;
        RECT 504.400 267.800 515.400 268.400 ;
        RECT 504.400 267.600 506.000 267.800 ;
        RECT 499.000 266.600 502.800 267.200 ;
        RECT 499.000 266.400 499.800 266.600 ;
        RECT 487.600 264.200 488.400 265.000 ;
        RECT 489.200 264.800 490.000 265.600 ;
        RECT 491.000 265.400 491.800 265.600 ;
        RECT 491.000 264.800 493.800 265.400 ;
        RECT 493.200 264.200 493.800 264.800 ;
        RECT 497.200 264.200 498.000 265.000 ;
        RECT 487.600 263.600 489.600 264.200 ;
        RECT 488.800 262.200 489.600 263.600 ;
        RECT 493.200 262.200 494.000 264.200 ;
        RECT 497.200 263.600 498.600 264.200 ;
        RECT 497.400 262.200 498.600 263.600 ;
        RECT 502.000 262.200 502.800 266.600 ;
        RECT 503.600 262.200 504.400 267.000 ;
        RECT 508.600 265.600 509.200 267.800 ;
        RECT 511.600 267.600 512.400 267.800 ;
        RECT 514.200 267.600 515.000 267.800 ;
        RECT 521.200 267.200 522.000 270.600 ;
        RECT 529.200 270.200 530.000 270.400 ;
        RECT 525.000 269.600 530.000 270.200 ;
        RECT 525.000 269.400 525.800 269.600 ;
        RECT 527.600 269.400 528.400 269.600 ;
        RECT 526.600 268.400 527.400 268.600 ;
        RECT 534.000 268.400 534.600 271.600 ;
        RECT 540.400 271.200 541.200 279.800 ;
        RECT 537.000 270.600 541.200 271.200 ;
        RECT 542.000 271.400 542.800 279.800 ;
        RECT 546.400 276.400 547.200 279.800 ;
        RECT 545.200 275.800 547.200 276.400 ;
        RECT 550.800 275.800 551.600 279.800 ;
        RECT 555.000 275.800 556.200 279.800 ;
        RECT 545.200 275.000 546.000 275.800 ;
        RECT 550.800 275.200 551.400 275.800 ;
        RECT 548.600 274.600 552.200 275.200 ;
        RECT 554.800 275.000 555.600 275.800 ;
        RECT 548.600 274.400 549.400 274.600 ;
        RECT 551.400 274.400 552.200 274.600 ;
        RECT 545.200 273.000 546.000 273.200 ;
        RECT 549.800 273.000 550.600 273.200 ;
        RECT 545.200 272.400 550.600 273.000 ;
        RECT 551.200 273.000 553.400 273.600 ;
        RECT 551.200 271.800 551.800 273.000 ;
        RECT 552.600 272.800 553.400 273.000 ;
        RECT 555.000 273.200 556.400 274.000 ;
        RECT 555.000 272.200 555.600 273.200 ;
        RECT 547.000 271.400 551.800 271.800 ;
        RECT 542.000 271.200 551.800 271.400 ;
        RECT 553.200 271.600 555.600 272.200 ;
        RECT 542.000 271.000 547.800 271.200 ;
        RECT 542.000 270.800 547.600 271.000 ;
        RECT 537.000 270.400 537.800 270.600 ;
        RECT 538.600 269.800 539.400 270.000 ;
        RECT 535.600 269.200 539.400 269.800 ;
        RECT 535.600 269.000 536.400 269.200 ;
        RECT 523.600 267.800 534.800 268.400 ;
        RECT 523.600 267.600 525.200 267.800 ;
        RECT 518.200 266.600 522.000 267.200 ;
        RECT 518.200 266.400 519.000 266.600 ;
        RECT 506.800 264.200 507.600 265.000 ;
        RECT 508.400 264.800 509.200 265.600 ;
        RECT 510.200 265.400 511.000 265.600 ;
        RECT 510.200 264.800 513.000 265.400 ;
        RECT 512.400 264.200 513.000 264.800 ;
        RECT 516.400 264.200 517.200 265.000 ;
        RECT 506.800 263.600 508.800 264.200 ;
        RECT 508.000 262.200 508.800 263.600 ;
        RECT 512.400 262.200 513.200 264.200 ;
        RECT 516.400 263.600 517.800 264.200 ;
        RECT 516.600 262.200 517.800 263.600 ;
        RECT 521.200 262.200 522.000 266.600 ;
        RECT 522.800 262.200 523.600 267.000 ;
        RECT 527.800 265.600 528.400 267.800 ;
        RECT 533.400 267.600 534.800 267.800 ;
        RECT 540.400 267.200 541.200 270.600 ;
        RECT 548.400 270.200 549.200 270.400 ;
        RECT 544.200 269.600 549.200 270.200 ;
        RECT 551.600 270.300 552.400 270.400 ;
        RECT 553.200 270.300 553.800 271.600 ;
        RECT 559.600 271.200 560.400 279.800 ;
        RECT 556.200 270.600 560.400 271.200 ;
        RECT 561.200 271.400 562.000 279.800 ;
        RECT 565.600 276.400 566.400 279.800 ;
        RECT 564.400 275.800 566.400 276.400 ;
        RECT 570.000 275.800 570.800 279.800 ;
        RECT 574.200 275.800 575.400 279.800 ;
        RECT 564.400 275.000 565.200 275.800 ;
        RECT 570.000 275.200 570.600 275.800 ;
        RECT 567.800 274.600 571.400 275.200 ;
        RECT 574.000 275.000 574.800 275.800 ;
        RECT 567.800 274.400 568.600 274.600 ;
        RECT 570.600 274.400 571.400 274.600 ;
        RECT 564.400 273.000 565.200 273.200 ;
        RECT 569.000 273.000 569.800 273.200 ;
        RECT 564.400 272.400 569.800 273.000 ;
        RECT 570.400 273.000 572.600 273.600 ;
        RECT 570.400 271.800 571.000 273.000 ;
        RECT 571.800 272.800 572.600 273.000 ;
        RECT 574.200 273.200 575.600 274.000 ;
        RECT 574.200 272.200 574.800 273.200 ;
        RECT 566.200 271.400 571.000 271.800 ;
        RECT 561.200 271.200 571.000 271.400 ;
        RECT 572.400 271.600 574.800 272.200 ;
        RECT 561.200 271.000 567.000 271.200 ;
        RECT 561.200 270.800 566.800 271.000 ;
        RECT 556.200 270.400 557.000 270.600 ;
        RECT 551.600 269.700 553.900 270.300 ;
        RECT 557.800 269.800 558.600 270.000 ;
        RECT 551.600 269.600 552.400 269.700 ;
        RECT 544.200 269.400 545.000 269.600 ;
        RECT 546.800 269.400 547.600 269.600 ;
        RECT 545.800 268.400 546.600 268.600 ;
        RECT 553.200 268.400 553.800 269.700 ;
        RECT 554.800 269.200 558.600 269.800 ;
        RECT 554.800 269.000 555.600 269.200 ;
        RECT 542.800 267.800 553.800 268.400 ;
        RECT 542.800 267.600 544.400 267.800 ;
        RECT 537.400 266.600 541.200 267.200 ;
        RECT 537.400 266.400 538.200 266.600 ;
        RECT 526.000 264.200 526.800 265.000 ;
        RECT 527.600 264.800 528.400 265.600 ;
        RECT 529.400 265.400 530.200 265.600 ;
        RECT 529.400 264.800 532.200 265.400 ;
        RECT 531.600 264.200 532.200 264.800 ;
        RECT 535.600 264.200 536.400 265.000 ;
        RECT 526.000 263.600 528.000 264.200 ;
        RECT 527.200 262.200 528.000 263.600 ;
        RECT 531.600 262.200 532.400 264.200 ;
        RECT 535.600 263.600 537.000 264.200 ;
        RECT 535.800 262.200 537.000 263.600 ;
        RECT 540.400 262.200 541.200 266.600 ;
        RECT 542.000 262.200 542.800 267.000 ;
        RECT 547.000 265.600 547.600 267.800 ;
        RECT 552.600 267.600 553.400 267.800 ;
        RECT 559.600 267.200 560.400 270.600 ;
        RECT 567.600 270.200 568.400 270.400 ;
        RECT 563.400 269.600 568.400 270.200 ;
        RECT 563.400 269.400 564.200 269.600 ;
        RECT 566.000 269.400 566.800 269.600 ;
        RECT 565.000 268.400 565.800 268.600 ;
        RECT 572.400 268.400 573.000 271.600 ;
        RECT 578.800 271.200 579.600 279.800 ;
        RECT 580.400 272.400 581.200 279.800 ;
        RECT 580.400 271.800 582.600 272.400 ;
        RECT 575.400 270.600 579.600 271.200 ;
        RECT 575.400 270.400 576.200 270.600 ;
        RECT 577.000 269.800 577.800 270.000 ;
        RECT 574.000 269.200 577.800 269.800 ;
        RECT 574.000 269.000 574.800 269.200 ;
        RECT 562.000 267.800 573.000 268.400 ;
        RECT 562.000 267.600 563.600 267.800 ;
        RECT 556.600 266.600 560.400 267.200 ;
        RECT 556.600 266.400 557.400 266.600 ;
        RECT 545.200 264.200 546.000 265.000 ;
        RECT 546.800 264.800 547.600 265.600 ;
        RECT 548.600 265.400 549.400 265.600 ;
        RECT 548.600 264.800 551.400 265.400 ;
        RECT 550.800 264.200 551.400 264.800 ;
        RECT 554.800 264.200 555.600 265.000 ;
        RECT 545.200 263.600 547.200 264.200 ;
        RECT 546.400 262.200 547.200 263.600 ;
        RECT 550.800 262.200 551.600 264.200 ;
        RECT 554.800 263.600 556.200 264.200 ;
        RECT 555.000 262.200 556.200 263.600 ;
        RECT 559.600 262.200 560.400 266.600 ;
        RECT 561.200 262.200 562.000 267.000 ;
        RECT 566.200 265.600 566.800 267.800 ;
        RECT 571.800 267.600 572.600 267.800 ;
        RECT 578.800 267.200 579.600 270.600 ;
        RECT 582.000 271.200 582.600 271.800 ;
        RECT 582.000 270.400 583.200 271.200 ;
        RECT 580.400 268.800 581.200 270.400 ;
        RECT 582.000 267.400 582.600 270.400 ;
        RECT 575.800 266.600 579.600 267.200 ;
        RECT 575.800 266.400 576.600 266.600 ;
        RECT 564.400 264.200 565.200 265.000 ;
        RECT 566.000 264.800 566.800 265.600 ;
        RECT 567.800 265.400 568.600 265.600 ;
        RECT 567.800 264.800 570.600 265.400 ;
        RECT 570.000 264.200 570.600 264.800 ;
        RECT 574.000 264.200 574.800 265.000 ;
        RECT 564.400 263.600 566.400 264.200 ;
        RECT 565.600 262.200 566.400 263.600 ;
        RECT 570.000 262.200 570.800 264.200 ;
        RECT 574.000 263.600 575.400 264.200 ;
        RECT 574.200 262.200 575.400 263.600 ;
        RECT 578.800 262.200 579.600 266.600 ;
        RECT 580.400 266.800 582.600 267.400 ;
        RECT 580.400 262.200 581.200 266.800 ;
        RECT 1.200 256.000 2.000 259.800 ;
        RECT 4.400 256.000 5.200 259.800 ;
        RECT 1.200 255.800 5.200 256.000 ;
        RECT 6.000 255.800 6.800 259.800 ;
        RECT 8.200 256.400 9.000 259.800 ;
        RECT 8.200 255.800 10.000 256.400 ;
        RECT 1.400 255.400 5.000 255.800 ;
        RECT 2.000 254.400 2.800 254.800 ;
        RECT 6.000 254.400 6.600 255.800 ;
        RECT 1.200 253.800 2.800 254.400 ;
        RECT 1.200 253.600 2.000 253.800 ;
        RECT 4.200 253.600 6.800 254.400 ;
        RECT 2.800 251.600 3.600 253.200 ;
        RECT 4.200 252.300 4.800 253.600 ;
        RECT 4.200 251.700 8.300 252.300 ;
        RECT 4.200 250.200 4.800 251.700 ;
        RECT 7.700 250.400 8.300 251.700 ;
        RECT 6.000 250.200 6.800 250.400 ;
        RECT 3.800 249.600 4.800 250.200 ;
        RECT 5.400 249.600 6.800 250.200 ;
        RECT 3.800 242.200 4.600 249.600 ;
        RECT 5.400 248.400 6.000 249.600 ;
        RECT 7.600 248.800 8.400 250.400 ;
        RECT 5.200 247.600 6.000 248.400 ;
        RECT 9.200 242.200 10.000 255.800 ;
        RECT 10.800 253.600 11.600 255.200 ;
        RECT 12.400 253.600 13.200 255.200 ;
        RECT 14.000 250.300 14.800 259.800 ;
        RECT 15.600 255.600 16.400 257.200 ;
        RECT 17.200 254.300 18.000 259.800 ;
        RECT 22.000 255.800 22.800 259.800 ;
        RECT 23.400 256.400 24.200 257.200 ;
        RECT 25.200 257.000 26.000 259.000 ;
        RECT 22.000 254.400 22.600 255.800 ;
        RECT 23.600 255.600 24.400 256.400 ;
        RECT 25.200 254.800 25.800 257.000 ;
        RECT 29.400 256.000 30.200 259.000 ;
        RECT 29.400 255.400 31.000 256.000 ;
        RECT 34.800 255.800 35.600 259.800 ;
        RECT 36.400 256.000 37.200 259.800 ;
        RECT 39.600 256.000 40.400 259.800 ;
        RECT 41.800 258.400 42.600 259.800 ;
        RECT 41.200 257.600 42.600 258.400 ;
        RECT 36.400 255.800 40.400 256.000 ;
        RECT 41.800 256.400 42.600 257.600 ;
        RECT 47.600 257.600 48.400 259.800 ;
        RECT 41.800 255.800 43.600 256.400 ;
        RECT 30.200 255.000 31.000 255.400 ;
        RECT 20.400 254.300 21.200 254.400 ;
        RECT 17.200 253.700 21.200 254.300 ;
        RECT 15.600 250.300 16.400 250.400 ;
        RECT 14.000 249.700 16.400 250.300 ;
        RECT 14.000 242.200 14.800 249.700 ;
        RECT 15.600 249.600 16.400 249.700 ;
        RECT 17.200 242.200 18.000 253.700 ;
        RECT 20.400 252.800 21.200 253.700 ;
        RECT 22.000 253.600 22.800 254.400 ;
        RECT 25.200 254.200 29.400 254.800 ;
        RECT 28.400 253.800 29.400 254.200 ;
        RECT 30.400 254.400 31.000 255.000 ;
        RECT 35.000 254.400 35.600 255.800 ;
        RECT 36.600 255.400 40.200 255.800 ;
        RECT 38.800 254.400 39.600 254.800 ;
        RECT 18.800 252.200 19.600 252.400 ;
        RECT 22.000 252.200 22.600 253.600 ;
        RECT 23.600 252.200 24.400 252.400 ;
        RECT 18.800 251.600 20.400 252.200 ;
        RECT 22.000 251.600 24.400 252.200 ;
        RECT 25.200 251.600 26.000 253.200 ;
        RECT 26.800 251.600 27.600 253.200 ;
        RECT 28.400 253.000 29.800 253.800 ;
        RECT 30.400 253.600 32.400 254.400 ;
        RECT 34.800 253.600 37.400 254.400 ;
        RECT 38.800 253.800 40.400 254.400 ;
        RECT 39.600 253.600 40.400 253.800 ;
        RECT 19.600 251.200 20.400 251.600 ;
        RECT 23.600 250.200 24.200 251.600 ;
        RECT 28.400 251.000 29.000 253.000 ;
        RECT 25.200 250.400 29.000 251.000 ;
        RECT 18.800 249.600 22.800 250.200 ;
        RECT 18.800 242.200 19.600 249.600 ;
        RECT 22.000 242.200 22.800 249.600 ;
        RECT 23.600 242.200 24.400 250.200 ;
        RECT 25.200 247.000 25.800 250.400 ;
        RECT 30.400 249.800 31.000 253.600 ;
        RECT 31.600 252.300 32.400 252.400 ;
        RECT 33.200 252.300 34.000 252.400 ;
        RECT 31.600 251.700 34.000 252.300 ;
        RECT 31.600 250.800 32.400 251.700 ;
        RECT 33.200 251.600 34.000 251.700 ;
        RECT 29.400 249.200 31.000 249.800 ;
        RECT 34.800 250.200 35.600 250.400 ;
        RECT 36.800 250.200 37.400 253.600 ;
        RECT 38.000 251.600 38.800 253.200 ;
        RECT 34.800 249.600 36.200 250.200 ;
        RECT 36.800 249.600 37.800 250.200 ;
        RECT 25.200 243.000 26.000 247.000 ;
        RECT 29.400 244.400 30.200 249.200 ;
        RECT 35.600 248.400 36.200 249.600 ;
        RECT 35.600 247.600 36.400 248.400 ;
        RECT 37.000 244.400 37.800 249.600 ;
        RECT 41.200 248.800 42.000 250.400 ;
        RECT 29.400 243.600 30.800 244.400 ;
        RECT 37.000 243.600 38.800 244.400 ;
        RECT 29.400 242.200 30.200 243.600 ;
        RECT 37.000 242.200 37.800 243.600 ;
        RECT 42.800 242.200 43.600 255.800 ;
        RECT 44.400 254.300 45.200 255.200 ;
        RECT 47.600 254.400 48.200 257.600 ;
        RECT 49.200 255.600 50.000 257.200 ;
        RECT 50.800 255.800 51.600 259.800 ;
        RECT 55.200 256.200 56.800 259.800 ;
        RECT 46.000 254.300 46.800 254.400 ;
        RECT 44.400 253.700 46.800 254.300 ;
        RECT 44.400 253.600 45.200 253.700 ;
        RECT 46.000 253.600 46.800 253.700 ;
        RECT 47.600 253.600 48.400 254.400 ;
        RECT 49.300 254.300 49.900 255.600 ;
        RECT 50.800 255.200 53.200 255.800 ;
        RECT 52.400 255.000 53.200 255.200 ;
        RECT 53.800 254.800 54.600 255.600 ;
        RECT 53.800 254.400 54.400 254.800 ;
        RECT 50.800 254.300 52.400 254.400 ;
        RECT 49.300 253.700 52.400 254.300 ;
        RECT 50.800 253.600 52.400 253.700 ;
        RECT 53.600 253.600 54.400 254.400 ;
        RECT 46.000 250.800 46.800 252.400 ;
        RECT 47.600 250.200 48.200 253.600 ;
        RECT 55.200 252.800 55.800 256.200 ;
        RECT 60.400 255.800 61.200 259.800 ;
        RECT 56.400 255.400 58.000 255.600 ;
        RECT 56.400 254.800 58.400 255.400 ;
        RECT 59.000 255.200 61.200 255.800 ;
        RECT 62.000 255.800 62.800 259.800 ;
        RECT 66.400 256.200 68.000 259.800 ;
        RECT 62.000 255.200 64.200 255.800 ;
        RECT 65.200 255.400 66.800 255.600 ;
        RECT 59.000 255.000 59.800 255.200 ;
        RECT 63.400 255.000 64.200 255.200 ;
        RECT 57.800 254.400 58.400 254.800 ;
        RECT 64.800 254.800 66.800 255.400 ;
        RECT 64.800 254.400 65.400 254.800 ;
        RECT 56.400 253.400 57.200 254.200 ;
        RECT 57.800 253.800 61.200 254.400 ;
        RECT 59.600 253.600 61.200 253.800 ;
        RECT 62.000 253.800 65.400 254.400 ;
        RECT 62.000 253.600 63.600 253.800 ;
        RECT 54.800 252.400 55.800 252.800 ;
        RECT 54.000 252.200 55.800 252.400 ;
        RECT 56.600 252.800 57.200 253.400 ;
        RECT 66.000 253.400 66.800 254.200 ;
        RECT 66.000 252.800 66.600 253.400 ;
        RECT 56.600 252.200 59.200 252.800 ;
        RECT 54.000 251.600 55.400 252.200 ;
        RECT 58.400 252.000 59.200 252.200 ;
        RECT 64.000 252.200 66.600 252.800 ;
        RECT 67.400 252.800 68.000 256.200 ;
        RECT 71.600 255.800 72.400 259.800 ;
        RECT 68.600 254.800 69.400 255.600 ;
        RECT 70.000 255.200 72.400 255.800 ;
        RECT 76.400 255.800 77.200 259.800 ;
        RECT 77.800 256.400 78.600 257.200 ;
        RECT 70.000 255.000 70.800 255.200 ;
        RECT 68.800 254.400 69.400 254.800 ;
        RECT 68.800 253.600 69.600 254.400 ;
        RECT 70.800 254.300 72.400 254.400 ;
        RECT 74.800 254.300 75.600 254.400 ;
        RECT 70.800 253.700 75.600 254.300 ;
        RECT 70.800 253.600 72.400 253.700 ;
        RECT 74.800 252.800 75.600 253.700 ;
        RECT 67.400 252.400 68.400 252.800 ;
        RECT 67.400 252.200 69.200 252.400 ;
        RECT 64.000 252.000 64.800 252.200 ;
        RECT 67.800 251.600 69.200 252.200 ;
        RECT 71.600 252.300 72.400 252.400 ;
        RECT 73.200 252.300 74.000 252.400 ;
        RECT 71.600 252.200 74.000 252.300 ;
        RECT 76.400 252.200 77.000 255.800 ;
        RECT 78.000 255.600 78.800 256.400 ;
        RECT 78.000 254.300 78.800 254.400 ;
        RECT 79.600 254.300 80.400 259.800 ;
        RECT 81.200 255.600 82.000 257.200 ;
        RECT 82.800 256.000 83.600 259.800 ;
        RECT 86.000 256.000 86.800 259.800 ;
        RECT 82.800 255.800 86.800 256.000 ;
        RECT 87.600 255.800 88.400 259.800 ;
        RECT 78.000 253.700 80.400 254.300 ;
        RECT 81.300 254.300 81.900 255.600 ;
        RECT 83.000 255.400 86.600 255.800 ;
        RECT 83.600 254.400 84.400 254.800 ;
        RECT 87.600 254.400 88.200 255.800 ;
        RECT 82.800 254.300 84.400 254.400 ;
        RECT 81.300 253.800 84.400 254.300 ;
        RECT 81.300 253.700 83.600 253.800 ;
        RECT 78.000 253.600 78.800 253.700 ;
        RECT 78.000 252.200 78.800 252.400 ;
        RECT 71.600 251.700 74.800 252.200 ;
        RECT 71.600 251.600 72.400 251.700 ;
        RECT 73.200 251.600 74.800 251.700 ;
        RECT 76.400 251.600 78.800 252.200 ;
        RECT 54.800 250.200 55.400 251.600 ;
        RECT 56.200 251.400 57.000 251.600 ;
        RECT 66.200 251.400 67.000 251.600 ;
        RECT 56.200 250.800 59.600 251.400 ;
        RECT 59.000 250.200 59.600 250.800 ;
        RECT 63.600 250.800 67.000 251.400 ;
        RECT 63.600 250.200 64.200 250.800 ;
        RECT 67.800 250.200 68.400 251.600 ;
        RECT 74.000 251.200 74.800 251.600 ;
        RECT 78.000 250.200 78.600 251.600 ;
        RECT 46.600 249.400 48.400 250.200 ;
        RECT 50.800 249.600 53.200 250.200 ;
        RECT 54.800 249.600 56.800 250.200 ;
        RECT 46.600 242.200 47.400 249.400 ;
        RECT 50.800 242.200 51.600 249.600 ;
        RECT 52.400 249.400 53.200 249.600 ;
        RECT 55.200 244.400 56.800 249.600 ;
        RECT 59.000 249.600 61.200 250.200 ;
        RECT 59.000 249.400 59.800 249.600 ;
        RECT 54.000 243.600 56.800 244.400 ;
        RECT 55.200 242.200 56.800 243.600 ;
        RECT 60.400 242.200 61.200 249.600 ;
        RECT 62.000 249.600 64.200 250.200 ;
        RECT 62.000 242.200 62.800 249.600 ;
        RECT 63.400 249.400 64.200 249.600 ;
        RECT 66.400 249.600 68.400 250.200 ;
        RECT 70.000 249.600 72.400 250.200 ;
        RECT 66.400 242.200 68.000 249.600 ;
        RECT 70.000 249.400 70.800 249.600 ;
        RECT 71.600 242.200 72.400 249.600 ;
        RECT 73.200 249.600 77.200 250.200 ;
        RECT 73.200 242.200 74.000 249.600 ;
        RECT 76.400 242.200 77.200 249.600 ;
        RECT 78.000 242.200 78.800 250.200 ;
        RECT 79.600 242.200 80.400 253.700 ;
        RECT 82.800 253.600 83.600 253.700 ;
        RECT 85.800 253.600 88.400 254.400 ;
        RECT 81.200 252.300 82.000 252.400 ;
        RECT 84.400 252.300 85.200 253.200 ;
        RECT 81.200 251.700 85.200 252.300 ;
        RECT 81.200 251.600 82.000 251.700 ;
        RECT 84.400 251.600 85.200 251.700 ;
        RECT 85.800 250.200 86.400 253.600 ;
        RECT 87.600 250.300 88.400 250.400 ;
        RECT 89.200 250.300 90.000 259.800 ;
        RECT 90.800 255.600 91.600 257.200 ;
        RECT 87.600 250.200 90.000 250.300 ;
        RECT 85.400 249.600 86.400 250.200 ;
        RECT 87.000 249.700 90.000 250.200 ;
        RECT 87.000 249.600 88.400 249.700 ;
        RECT 85.400 242.200 86.200 249.600 ;
        RECT 87.000 248.400 87.600 249.600 ;
        RECT 86.800 247.600 87.600 248.400 ;
        RECT 89.200 242.200 90.000 249.700 ;
        RECT 90.800 248.300 91.600 248.400 ;
        RECT 92.400 248.300 93.200 259.800 ;
        RECT 94.000 255.600 94.800 257.200 ;
        RECT 99.200 254.200 100.000 259.800 ;
        RECT 102.000 256.000 102.800 259.800 ;
        RECT 105.200 256.000 106.000 259.800 ;
        RECT 102.000 255.800 106.000 256.000 ;
        RECT 106.800 255.800 107.600 259.800 ;
        RECT 102.200 255.400 105.800 255.800 ;
        RECT 102.800 254.400 103.600 254.800 ;
        RECT 106.800 254.400 107.400 255.800 ;
        RECT 99.200 253.800 101.000 254.200 ;
        RECT 99.400 253.600 101.000 253.800 ;
        RECT 102.000 253.800 103.600 254.400 ;
        RECT 102.000 253.600 102.800 253.800 ;
        RECT 105.000 253.600 107.600 254.400 ;
        RECT 97.200 251.600 98.800 252.400 ;
        RECT 94.000 250.300 94.800 250.400 ;
        RECT 95.600 250.300 96.400 251.200 ;
        RECT 94.000 249.700 96.400 250.300 ;
        RECT 94.000 249.600 94.800 249.700 ;
        RECT 95.600 249.600 96.400 249.700 ;
        RECT 100.400 250.400 101.000 253.600 ;
        RECT 103.600 251.600 104.400 253.200 ;
        RECT 100.400 249.600 101.200 250.400 ;
        RECT 105.000 250.200 105.600 253.600 ;
        RECT 106.800 250.300 107.600 250.400 ;
        RECT 108.400 250.300 109.200 259.800 ;
        RECT 113.200 257.800 114.000 259.800 ;
        RECT 110.000 255.600 110.800 257.200 ;
        RECT 113.200 254.400 113.800 257.800 ;
        RECT 114.800 255.600 115.600 257.200 ;
        RECT 116.400 255.800 117.200 259.800 ;
        RECT 118.000 256.000 118.800 259.800 ;
        RECT 121.200 256.000 122.000 259.800 ;
        RECT 124.400 257.800 125.200 259.800 ;
        RECT 118.000 255.800 122.000 256.000 ;
        RECT 122.800 256.300 123.600 256.400 ;
        RECT 124.400 256.300 125.000 257.800 ;
        RECT 116.600 254.400 117.200 255.800 ;
        RECT 118.200 255.400 121.800 255.800 ;
        RECT 122.800 255.700 125.100 256.300 ;
        RECT 122.800 255.600 123.600 255.700 ;
        RECT 120.400 254.400 121.200 254.800 ;
        RECT 124.400 254.400 125.000 255.700 ;
        RECT 126.000 255.600 126.800 257.200 ;
        RECT 127.600 255.800 128.400 259.800 ;
        RECT 132.000 256.200 133.600 259.800 ;
        RECT 127.600 255.200 129.800 255.800 ;
        RECT 130.800 255.400 132.400 255.600 ;
        RECT 129.000 255.000 129.800 255.200 ;
        RECT 130.400 254.800 132.400 255.400 ;
        RECT 130.400 254.400 131.000 254.800 ;
        RECT 113.200 253.600 114.000 254.400 ;
        RECT 116.400 253.600 119.000 254.400 ;
        RECT 120.400 253.800 122.000 254.400 ;
        RECT 121.200 253.600 122.000 253.800 ;
        RECT 124.400 253.600 125.200 254.400 ;
        RECT 127.600 253.800 131.000 254.400 ;
        RECT 127.600 253.600 129.200 253.800 ;
        RECT 113.200 252.400 113.800 253.600 ;
        RECT 111.600 250.800 112.400 252.400 ;
        RECT 113.200 251.600 114.000 252.400 ;
        RECT 106.800 250.200 109.200 250.300 ;
        RECT 113.200 250.200 113.800 251.600 ;
        RECT 116.400 250.200 117.200 250.400 ;
        RECT 118.400 250.200 119.000 253.600 ;
        RECT 119.600 251.600 120.400 253.200 ;
        RECT 121.300 252.300 121.900 253.600 ;
        RECT 122.800 252.300 123.600 252.400 ;
        RECT 121.300 251.700 123.600 252.300 ;
        RECT 122.800 250.800 123.600 251.700 ;
        RECT 124.400 250.200 125.000 253.600 ;
        RECT 131.600 253.400 132.400 254.200 ;
        RECT 131.600 252.800 132.200 253.400 ;
        RECT 129.600 252.200 132.200 252.800 ;
        RECT 133.000 252.800 133.600 256.200 ;
        RECT 137.200 255.800 138.000 259.800 ;
        RECT 134.200 254.800 135.000 255.600 ;
        RECT 135.600 255.200 138.000 255.800 ;
        RECT 143.600 255.800 144.400 259.800 ;
        RECT 148.000 256.200 149.600 259.800 ;
        RECT 143.600 255.200 145.800 255.800 ;
        RECT 146.800 255.400 148.400 255.600 ;
        RECT 135.600 255.000 136.400 255.200 ;
        RECT 145.000 255.000 145.800 255.200 ;
        RECT 134.400 254.400 135.000 254.800 ;
        RECT 146.400 254.800 148.400 255.400 ;
        RECT 146.400 254.400 147.000 254.800 ;
        RECT 134.400 253.600 135.200 254.400 ;
        RECT 136.400 253.600 138.000 254.400 ;
        RECT 142.000 254.300 142.800 254.400 ;
        RECT 143.600 254.300 147.000 254.400 ;
        RECT 142.000 253.800 147.000 254.300 ;
        RECT 142.000 253.700 145.200 253.800 ;
        RECT 142.000 253.600 142.800 253.700 ;
        RECT 143.600 253.600 145.200 253.700 ;
        RECT 147.600 253.400 148.400 254.200 ;
        RECT 147.600 252.800 148.200 253.400 ;
        RECT 133.000 252.400 134.000 252.800 ;
        RECT 133.000 252.200 134.800 252.400 ;
        RECT 129.600 252.000 130.400 252.200 ;
        RECT 133.400 251.600 134.800 252.200 ;
        RECT 145.600 252.200 148.200 252.800 ;
        RECT 149.000 252.800 149.600 256.200 ;
        RECT 153.200 255.800 154.000 259.800 ;
        RECT 157.400 258.400 158.200 259.800 ;
        RECT 157.400 257.600 158.800 258.400 ;
        RECT 157.400 256.400 158.200 257.600 ;
        RECT 150.200 254.800 151.000 255.600 ;
        RECT 151.600 255.200 154.000 255.800 ;
        RECT 156.400 255.800 158.200 256.400 ;
        RECT 159.600 256.000 160.400 259.800 ;
        RECT 162.800 256.000 163.600 259.800 ;
        RECT 159.600 255.800 163.600 256.000 ;
        RECT 164.400 255.800 165.200 259.800 ;
        RECT 166.600 256.400 167.400 259.800 ;
        RECT 166.600 255.800 168.400 256.400 ;
        RECT 170.800 255.800 171.600 259.800 ;
        RECT 172.400 256.000 173.200 259.800 ;
        RECT 175.600 256.000 176.400 259.800 ;
        RECT 172.400 255.800 176.400 256.000 ;
        RECT 178.800 257.800 179.600 259.800 ;
        RECT 151.600 255.000 152.400 255.200 ;
        RECT 150.400 254.400 151.000 254.800 ;
        RECT 150.400 253.600 151.200 254.400 ;
        RECT 152.400 253.600 154.000 254.400 ;
        RECT 154.800 253.600 155.600 255.200 ;
        RECT 149.000 252.400 150.000 252.800 ;
        RECT 149.000 252.200 150.800 252.400 ;
        RECT 145.600 252.000 146.400 252.200 ;
        RECT 149.400 251.600 150.800 252.200 ;
        RECT 131.800 251.400 132.600 251.600 ;
        RECT 129.200 250.800 132.600 251.400 ;
        RECT 129.200 250.200 129.800 250.800 ;
        RECT 133.400 250.200 134.000 251.600 ;
        RECT 147.800 251.400 148.600 251.600 ;
        RECT 145.200 250.800 148.600 251.400 ;
        RECT 145.200 250.200 145.800 250.800 ;
        RECT 149.400 250.200 150.000 251.600 ;
        RECT 104.600 249.600 105.600 250.200 ;
        RECT 106.200 249.700 109.200 250.200 ;
        RECT 106.200 249.600 107.600 249.700 ;
        RECT 90.800 247.700 93.200 248.300 ;
        RECT 90.800 247.600 91.600 247.700 ;
        RECT 92.400 242.200 93.200 247.700 ;
        RECT 98.800 247.600 99.600 249.200 ;
        RECT 100.400 247.000 101.000 249.600 ;
        RECT 104.600 248.400 105.400 249.600 ;
        RECT 106.200 248.400 106.800 249.600 ;
        RECT 103.600 247.600 105.400 248.400 ;
        RECT 106.000 247.600 106.800 248.400 ;
        RECT 97.400 246.400 101.000 247.000 ;
        RECT 97.400 246.200 98.000 246.400 ;
        RECT 97.200 242.200 98.000 246.200 ;
        RECT 100.400 246.200 101.000 246.400 ;
        RECT 100.400 242.200 101.200 246.200 ;
        RECT 104.600 242.200 105.400 247.600 ;
        RECT 108.400 242.200 109.200 249.700 ;
        RECT 112.200 249.400 114.000 250.200 ;
        RECT 116.400 249.600 117.800 250.200 ;
        RECT 118.400 249.600 119.400 250.200 ;
        RECT 112.200 242.200 113.000 249.400 ;
        RECT 117.200 248.400 117.800 249.600 ;
        RECT 117.200 247.600 118.000 248.400 ;
        RECT 118.600 242.200 119.400 249.600 ;
        RECT 123.400 249.400 125.200 250.200 ;
        RECT 127.600 249.600 129.800 250.200 ;
        RECT 123.400 242.200 124.200 249.400 ;
        RECT 127.600 242.200 128.400 249.600 ;
        RECT 129.000 249.400 129.800 249.600 ;
        RECT 132.000 249.600 134.000 250.200 ;
        RECT 135.600 249.600 138.000 250.200 ;
        RECT 132.000 244.400 133.600 249.600 ;
        RECT 135.600 249.400 136.400 249.600 ;
        RECT 130.800 243.600 133.600 244.400 ;
        RECT 132.000 242.200 133.600 243.600 ;
        RECT 137.200 242.200 138.000 249.600 ;
        RECT 143.600 249.600 145.800 250.200 ;
        RECT 143.600 242.200 144.400 249.600 ;
        RECT 145.000 249.400 145.800 249.600 ;
        RECT 148.000 249.600 150.000 250.200 ;
        RECT 151.600 249.600 154.000 250.200 ;
        RECT 148.000 244.400 149.600 249.600 ;
        RECT 151.600 249.400 152.400 249.600 ;
        RECT 146.800 243.600 149.600 244.400 ;
        RECT 148.000 242.200 149.600 243.600 ;
        RECT 153.200 242.200 154.000 249.600 ;
        RECT 156.400 242.200 157.200 255.800 ;
        RECT 159.800 255.400 163.400 255.800 ;
        RECT 160.400 254.400 161.200 254.800 ;
        RECT 164.400 254.400 165.000 255.800 ;
        RECT 159.600 253.800 161.200 254.400 ;
        RECT 159.600 253.600 160.400 253.800 ;
        RECT 162.600 253.600 165.200 254.400 ;
        RECT 161.200 252.300 162.000 253.200 ;
        RECT 158.100 251.700 162.000 252.300 ;
        RECT 158.100 250.400 158.700 251.700 ;
        RECT 161.200 251.600 162.000 251.700 ;
        RECT 162.600 252.400 163.200 253.600 ;
        RECT 162.600 251.600 163.600 252.400 ;
        RECT 158.000 248.800 158.800 250.400 ;
        RECT 162.600 250.200 163.200 251.600 ;
        RECT 164.400 250.300 165.200 250.400 ;
        RECT 166.000 250.300 166.800 250.400 ;
        RECT 164.400 250.200 166.800 250.300 ;
        RECT 162.200 249.600 163.200 250.200 ;
        RECT 163.800 249.700 166.800 250.200 ;
        RECT 163.800 249.600 165.200 249.700 ;
        RECT 162.200 242.200 163.000 249.600 ;
        RECT 163.800 248.400 164.400 249.600 ;
        RECT 166.000 248.800 166.800 249.700 ;
        RECT 167.600 250.300 168.400 255.800 ;
        RECT 169.200 253.600 170.000 255.200 ;
        RECT 171.000 254.400 171.600 255.800 ;
        RECT 172.600 255.400 176.200 255.800 ;
        RECT 174.800 254.400 175.600 254.800 ;
        RECT 178.800 254.400 179.400 257.800 ;
        RECT 180.400 255.600 181.200 257.200 ;
        RECT 182.000 255.800 182.800 259.800 ;
        RECT 183.600 256.000 184.400 259.800 ;
        RECT 186.800 256.000 187.600 259.800 ;
        RECT 183.600 255.800 187.600 256.000 ;
        RECT 182.200 254.400 182.800 255.800 ;
        RECT 183.800 255.400 187.400 255.800 ;
        RECT 186.000 254.400 186.800 254.800 ;
        RECT 170.800 253.600 173.400 254.400 ;
        RECT 174.800 253.800 176.400 254.400 ;
        RECT 175.600 253.600 176.400 253.800 ;
        RECT 178.800 253.600 179.600 254.400 ;
        RECT 182.000 253.600 184.600 254.400 ;
        RECT 186.000 254.300 187.600 254.400 ;
        RECT 188.400 254.300 189.200 259.800 ;
        RECT 190.000 255.600 190.800 257.200 ;
        RECT 186.000 253.800 189.200 254.300 ;
        RECT 186.800 253.700 189.200 253.800 ;
        RECT 186.800 253.600 187.600 253.700 ;
        RECT 170.800 250.300 171.600 250.400 ;
        RECT 167.600 250.200 171.600 250.300 ;
        RECT 172.800 250.200 173.400 253.600 ;
        RECT 174.000 252.300 174.800 253.200 ;
        RECT 175.600 252.300 176.400 252.400 ;
        RECT 174.000 251.700 176.400 252.300 ;
        RECT 174.000 251.600 174.800 251.700 ;
        RECT 175.600 251.600 176.400 251.700 ;
        RECT 177.200 250.800 178.000 252.400 ;
        RECT 178.800 250.200 179.400 253.600 ;
        RECT 182.000 250.200 182.800 250.400 ;
        RECT 184.000 250.200 184.600 253.600 ;
        RECT 185.200 252.300 186.000 253.200 ;
        RECT 186.800 252.300 187.600 252.400 ;
        RECT 185.200 251.700 187.600 252.300 ;
        RECT 185.200 251.600 186.000 251.700 ;
        RECT 186.800 251.600 187.600 251.700 ;
        RECT 167.600 249.700 172.200 250.200 ;
        RECT 163.600 247.600 164.400 248.400 ;
        RECT 167.600 242.200 168.400 249.700 ;
        RECT 170.800 249.600 172.200 249.700 ;
        RECT 172.800 249.600 173.800 250.200 ;
        RECT 171.600 248.400 172.200 249.600 ;
        RECT 171.600 247.600 172.400 248.400 ;
        RECT 173.000 242.200 173.800 249.600 ;
        RECT 177.800 249.400 179.600 250.200 ;
        RECT 182.000 249.600 183.400 250.200 ;
        RECT 184.000 249.600 185.000 250.200 ;
        RECT 177.800 248.400 178.600 249.400 ;
        RECT 177.200 247.600 178.600 248.400 ;
        RECT 182.800 248.400 183.400 249.600 ;
        RECT 182.800 247.600 183.600 248.400 ;
        RECT 177.800 242.200 178.600 247.600 ;
        RECT 184.200 244.400 185.000 249.600 ;
        RECT 184.200 243.600 186.000 244.400 ;
        RECT 184.200 242.200 185.000 243.600 ;
        RECT 188.400 242.200 189.200 253.700 ;
        RECT 190.000 252.300 190.800 252.400 ;
        RECT 191.600 252.300 192.400 259.800 ;
        RECT 196.400 257.800 197.200 259.800 ;
        RECT 193.200 255.600 194.000 257.200 ;
        RECT 196.400 254.400 197.000 257.800 ;
        RECT 198.000 255.600 198.800 257.200 ;
        RECT 199.600 255.400 200.400 259.800 ;
        RECT 203.800 258.400 205.000 259.800 ;
        RECT 203.800 257.800 205.200 258.400 ;
        RECT 208.400 257.800 209.200 259.800 ;
        RECT 212.800 258.400 213.600 259.800 ;
        RECT 212.800 257.800 214.800 258.400 ;
        RECT 204.400 257.000 205.200 257.800 ;
        RECT 208.600 257.200 209.200 257.800 ;
        RECT 208.600 256.600 211.400 257.200 ;
        RECT 210.600 256.400 211.400 256.600 ;
        RECT 212.400 256.400 213.200 257.200 ;
        RECT 214.000 257.000 214.800 257.800 ;
        RECT 202.600 255.400 203.400 255.600 ;
        RECT 199.600 254.800 203.400 255.400 ;
        RECT 196.400 253.600 197.200 254.400 ;
        RECT 190.000 251.700 192.400 252.300 ;
        RECT 190.000 251.600 190.800 251.700 ;
        RECT 191.600 242.200 192.400 251.700 ;
        RECT 193.200 252.300 194.000 252.400 ;
        RECT 194.800 252.300 195.600 252.400 ;
        RECT 193.200 251.700 195.600 252.300 ;
        RECT 193.200 251.600 194.000 251.700 ;
        RECT 194.800 250.800 195.600 251.700 ;
        RECT 196.400 250.200 197.000 253.600 ;
        RECT 199.600 251.400 200.400 254.800 ;
        RECT 206.600 254.200 207.400 254.400 ;
        RECT 212.400 254.200 213.000 256.400 ;
        RECT 217.200 255.000 218.000 259.800 ;
        RECT 218.800 255.400 219.600 259.800 ;
        RECT 223.000 258.400 224.200 259.800 ;
        RECT 223.000 257.800 224.400 258.400 ;
        RECT 227.600 257.800 228.400 259.800 ;
        RECT 232.000 258.400 232.800 259.800 ;
        RECT 232.000 257.800 234.000 258.400 ;
        RECT 223.600 257.000 224.400 257.800 ;
        RECT 227.800 257.200 228.400 257.800 ;
        RECT 227.800 256.600 230.600 257.200 ;
        RECT 229.800 256.400 230.600 256.600 ;
        RECT 231.600 255.600 232.400 257.200 ;
        RECT 233.200 257.000 234.000 257.800 ;
        RECT 221.800 255.400 222.600 255.600 ;
        RECT 218.800 254.800 222.600 255.400 ;
        RECT 215.600 254.200 217.200 254.400 ;
        RECT 206.200 253.600 217.200 254.200 ;
        RECT 204.400 252.800 205.200 253.000 ;
        RECT 201.400 252.200 205.200 252.800 ;
        RECT 206.200 252.400 206.800 253.600 ;
        RECT 213.400 253.400 214.200 253.600 ;
        RECT 212.400 252.400 213.200 252.600 ;
        RECT 215.000 252.400 215.800 252.600 ;
        RECT 201.400 252.000 202.200 252.200 ;
        RECT 206.000 251.600 206.800 252.400 ;
        RECT 210.800 251.800 215.800 252.400 ;
        RECT 210.800 251.600 211.600 251.800 ;
        RECT 203.000 251.400 203.800 251.600 ;
        RECT 199.600 250.800 203.800 251.400 ;
        RECT 195.400 249.400 197.200 250.200 ;
        RECT 193.200 248.300 194.000 248.400 ;
        RECT 195.400 248.300 196.200 249.400 ;
        RECT 193.200 247.700 196.200 248.300 ;
        RECT 193.200 247.600 194.000 247.700 ;
        RECT 195.400 242.200 196.200 247.700 ;
        RECT 199.600 242.200 200.400 250.800 ;
        RECT 206.200 250.400 206.800 251.600 ;
        RECT 218.800 251.400 219.600 254.800 ;
        RECT 225.800 254.200 226.600 254.400 ;
        RECT 231.600 254.200 232.200 255.600 ;
        RECT 236.400 255.000 237.200 259.800 ;
        RECT 234.800 254.200 236.400 254.400 ;
        RECT 225.400 253.600 236.400 254.200 ;
        RECT 223.600 252.800 224.400 253.000 ;
        RECT 220.600 252.200 224.400 252.800 ;
        RECT 225.400 252.400 226.000 253.600 ;
        RECT 232.600 253.400 233.400 253.600 ;
        RECT 234.200 252.400 235.000 252.600 ;
        RECT 220.600 252.000 221.400 252.200 ;
        RECT 225.200 251.600 226.000 252.400 ;
        RECT 230.000 251.800 235.000 252.400 ;
        RECT 238.000 252.400 238.800 259.800 ;
        RECT 241.200 255.200 242.000 259.800 ;
        RECT 239.800 254.600 242.000 255.200 ;
        RECT 242.800 255.400 243.600 259.800 ;
        RECT 247.000 258.400 248.200 259.800 ;
        RECT 247.000 257.800 248.400 258.400 ;
        RECT 251.600 257.800 252.400 259.800 ;
        RECT 256.000 258.400 256.800 259.800 ;
        RECT 256.000 257.800 258.000 258.400 ;
        RECT 247.600 257.000 248.400 257.800 ;
        RECT 251.800 257.200 252.400 257.800 ;
        RECT 251.800 256.600 254.600 257.200 ;
        RECT 253.800 256.400 254.600 256.600 ;
        RECT 255.600 256.400 256.400 257.200 ;
        RECT 257.200 257.000 258.000 257.800 ;
        RECT 245.800 255.400 246.600 255.600 ;
        RECT 242.800 254.800 246.600 255.400 ;
        RECT 230.000 251.600 230.800 251.800 ;
        RECT 222.200 251.400 223.000 251.600 ;
        RECT 212.400 251.000 218.000 251.200 ;
        RECT 212.200 250.800 218.000 251.000 ;
        RECT 204.400 249.800 206.800 250.400 ;
        RECT 208.200 250.600 218.000 250.800 ;
        RECT 208.200 250.200 213.000 250.600 ;
        RECT 204.400 248.800 205.000 249.800 ;
        RECT 203.600 248.000 205.000 248.800 ;
        RECT 206.600 249.000 207.400 249.200 ;
        RECT 208.200 249.000 208.800 250.200 ;
        RECT 206.600 248.400 208.800 249.000 ;
        RECT 209.400 249.000 214.800 249.600 ;
        RECT 209.400 248.800 210.200 249.000 ;
        RECT 214.000 248.800 214.800 249.000 ;
        RECT 207.800 247.400 208.600 247.600 ;
        RECT 210.600 247.400 211.400 247.600 ;
        RECT 204.400 246.200 205.200 247.000 ;
        RECT 207.800 246.800 211.400 247.400 ;
        RECT 208.600 246.200 209.200 246.800 ;
        RECT 214.000 246.200 214.800 247.000 ;
        RECT 203.800 242.200 205.000 246.200 ;
        RECT 208.400 242.200 209.200 246.200 ;
        RECT 212.800 245.600 214.800 246.200 ;
        RECT 212.800 242.200 213.600 245.600 ;
        RECT 217.200 242.200 218.000 250.600 ;
        RECT 218.800 250.800 223.000 251.400 ;
        RECT 218.800 242.200 219.600 250.800 ;
        RECT 225.400 250.400 226.000 251.600 ;
        RECT 231.600 251.000 237.200 251.200 ;
        RECT 231.400 250.800 237.200 251.000 ;
        RECT 223.600 249.800 226.000 250.400 ;
        RECT 227.400 250.600 237.200 250.800 ;
        RECT 227.400 250.200 232.200 250.600 ;
        RECT 223.600 248.800 224.200 249.800 ;
        RECT 222.800 248.000 224.200 248.800 ;
        RECT 225.800 249.000 226.600 249.200 ;
        RECT 227.400 249.000 228.000 250.200 ;
        RECT 225.800 248.400 228.000 249.000 ;
        RECT 228.600 249.000 234.000 249.600 ;
        RECT 228.600 248.800 229.400 249.000 ;
        RECT 233.200 248.800 234.000 249.000 ;
        RECT 227.000 247.400 227.800 247.600 ;
        RECT 229.800 247.400 230.600 247.600 ;
        RECT 223.600 246.200 224.400 247.000 ;
        RECT 227.000 246.800 230.600 247.400 ;
        RECT 227.800 246.200 228.400 246.800 ;
        RECT 233.200 246.200 234.000 247.000 ;
        RECT 223.000 242.200 224.200 246.200 ;
        RECT 227.600 242.200 228.400 246.200 ;
        RECT 232.000 245.600 234.000 246.200 ;
        RECT 232.000 242.200 232.800 245.600 ;
        RECT 236.400 242.200 237.200 250.600 ;
        RECT 238.000 250.200 238.600 252.400 ;
        RECT 239.800 251.600 240.400 254.600 ;
        RECT 241.200 251.600 242.000 253.200 ;
        RECT 239.200 250.800 240.400 251.600 ;
        RECT 239.800 250.200 240.400 250.800 ;
        RECT 242.800 251.400 243.600 254.800 ;
        RECT 249.800 254.200 250.600 254.400 ;
        RECT 255.600 254.200 256.200 256.400 ;
        RECT 260.400 255.000 261.200 259.800 ;
        RECT 262.000 255.400 262.800 259.800 ;
        RECT 266.200 258.400 267.400 259.800 ;
        RECT 266.200 257.800 267.600 258.400 ;
        RECT 270.800 257.800 271.600 259.800 ;
        RECT 275.200 258.400 276.000 259.800 ;
        RECT 275.200 257.800 277.200 258.400 ;
        RECT 266.800 257.000 267.600 257.800 ;
        RECT 271.000 257.200 271.600 257.800 ;
        RECT 271.000 256.600 273.800 257.200 ;
        RECT 273.000 256.400 273.800 256.600 ;
        RECT 274.800 256.400 275.600 257.200 ;
        RECT 276.400 257.000 277.200 257.800 ;
        RECT 265.000 255.400 265.800 255.600 ;
        RECT 262.000 254.800 265.800 255.400 ;
        RECT 258.800 254.200 260.400 254.400 ;
        RECT 249.400 253.600 260.400 254.200 ;
        RECT 247.600 252.800 248.400 253.000 ;
        RECT 244.600 252.200 248.400 252.800 ;
        RECT 244.600 252.000 245.400 252.200 ;
        RECT 246.200 251.400 247.000 251.600 ;
        RECT 242.800 250.800 247.000 251.400 ;
        RECT 238.000 242.200 238.800 250.200 ;
        RECT 239.800 249.600 242.000 250.200 ;
        RECT 241.200 242.200 242.000 249.600 ;
        RECT 242.800 242.200 243.600 250.800 ;
        RECT 249.400 250.400 250.000 253.600 ;
        RECT 256.600 253.400 257.400 253.600 ;
        RECT 255.600 252.400 256.400 252.600 ;
        RECT 258.200 252.400 259.000 252.600 ;
        RECT 254.000 251.800 259.000 252.400 ;
        RECT 254.000 251.600 254.800 251.800 ;
        RECT 262.000 251.400 262.800 254.800 ;
        RECT 269.000 254.200 269.800 254.400 ;
        RECT 274.800 254.200 275.400 256.400 ;
        RECT 279.600 255.000 280.400 259.800 ;
        RECT 278.000 254.200 279.600 254.400 ;
        RECT 268.600 253.600 279.600 254.200 ;
        RECT 266.800 252.800 267.600 253.000 ;
        RECT 263.800 252.200 267.600 252.800 ;
        RECT 268.600 252.400 269.200 253.600 ;
        RECT 275.800 253.400 276.600 253.600 ;
        RECT 274.800 252.400 275.600 252.600 ;
        RECT 277.400 252.400 278.200 252.600 ;
        RECT 263.800 252.000 264.600 252.200 ;
        RECT 268.400 251.600 269.200 252.400 ;
        RECT 273.200 251.800 278.200 252.400 ;
        RECT 281.200 252.400 282.000 259.800 ;
        RECT 284.400 255.200 285.200 259.800 ;
        RECT 289.200 258.300 290.000 258.400 ;
        RECT 290.800 258.300 291.600 259.800 ;
        RECT 289.200 257.700 291.600 258.300 ;
        RECT 295.000 258.400 296.200 259.800 ;
        RECT 295.000 257.800 296.400 258.400 ;
        RECT 299.600 257.800 300.400 259.800 ;
        RECT 304.000 258.400 304.800 259.800 ;
        RECT 304.000 257.800 306.000 258.400 ;
        RECT 289.200 257.600 290.000 257.700 ;
        RECT 283.000 254.600 285.200 255.200 ;
        RECT 290.800 255.400 291.600 257.700 ;
        RECT 295.600 257.000 296.400 257.800 ;
        RECT 299.800 257.200 300.400 257.800 ;
        RECT 299.800 256.600 302.600 257.200 ;
        RECT 301.800 256.400 302.600 256.600 ;
        RECT 303.600 256.400 304.400 257.200 ;
        RECT 305.200 257.000 306.000 257.800 ;
        RECT 293.800 255.400 294.600 255.600 ;
        RECT 290.800 254.800 294.600 255.400 ;
        RECT 273.200 251.600 274.000 251.800 ;
        RECT 265.400 251.400 266.200 251.600 ;
        RECT 255.600 251.000 261.200 251.200 ;
        RECT 255.400 250.800 261.200 251.000 ;
        RECT 247.600 249.800 250.000 250.400 ;
        RECT 251.400 250.600 261.200 250.800 ;
        RECT 251.400 250.200 256.200 250.600 ;
        RECT 247.600 248.800 248.200 249.800 ;
        RECT 246.800 248.000 248.200 248.800 ;
        RECT 249.800 249.000 250.600 249.200 ;
        RECT 251.400 249.000 252.000 250.200 ;
        RECT 249.800 248.400 252.000 249.000 ;
        RECT 252.600 249.000 258.000 249.600 ;
        RECT 252.600 248.800 253.400 249.000 ;
        RECT 257.200 248.800 258.000 249.000 ;
        RECT 251.000 247.400 251.800 247.600 ;
        RECT 253.800 247.400 254.600 247.600 ;
        RECT 247.600 246.200 248.400 247.000 ;
        RECT 251.000 246.800 254.600 247.400 ;
        RECT 251.800 246.200 252.400 246.800 ;
        RECT 257.200 246.200 258.000 247.000 ;
        RECT 247.000 242.200 248.200 246.200 ;
        RECT 251.600 242.200 252.400 246.200 ;
        RECT 256.000 245.600 258.000 246.200 ;
        RECT 256.000 242.200 256.800 245.600 ;
        RECT 260.400 242.200 261.200 250.600 ;
        RECT 262.000 250.800 266.200 251.400 ;
        RECT 262.000 242.200 262.800 250.800 ;
        RECT 268.600 250.400 269.200 251.600 ;
        RECT 274.800 251.000 280.400 251.200 ;
        RECT 274.600 250.800 280.400 251.000 ;
        RECT 266.800 249.800 269.200 250.400 ;
        RECT 270.600 250.600 280.400 250.800 ;
        RECT 270.600 250.200 275.400 250.600 ;
        RECT 266.800 248.800 267.400 249.800 ;
        RECT 266.000 248.000 267.400 248.800 ;
        RECT 269.000 249.000 269.800 249.200 ;
        RECT 270.600 249.000 271.200 250.200 ;
        RECT 269.000 248.400 271.200 249.000 ;
        RECT 271.800 249.000 277.200 249.600 ;
        RECT 271.800 248.800 272.600 249.000 ;
        RECT 276.400 248.800 277.200 249.000 ;
        RECT 270.200 247.400 271.000 247.600 ;
        RECT 273.000 247.400 273.800 247.600 ;
        RECT 266.800 246.200 267.600 247.000 ;
        RECT 270.200 246.800 273.800 247.400 ;
        RECT 271.000 246.200 271.600 246.800 ;
        RECT 276.400 246.200 277.200 247.000 ;
        RECT 266.200 242.200 267.400 246.200 ;
        RECT 270.800 242.200 271.600 246.200 ;
        RECT 275.200 245.600 277.200 246.200 ;
        RECT 275.200 242.200 276.000 245.600 ;
        RECT 279.600 242.200 280.400 250.600 ;
        RECT 281.200 250.200 281.800 252.400 ;
        RECT 283.000 251.600 283.600 254.600 ;
        RECT 284.400 252.300 285.200 253.200 ;
        RECT 289.200 252.300 290.000 252.400 ;
        RECT 284.400 251.700 290.000 252.300 ;
        RECT 284.400 251.600 285.200 251.700 ;
        RECT 289.200 251.600 290.000 251.700 ;
        RECT 282.400 250.800 283.600 251.600 ;
        RECT 283.000 250.200 283.600 250.800 ;
        RECT 290.800 251.400 291.600 254.800 ;
        RECT 297.800 254.200 298.600 254.400 ;
        RECT 303.600 254.200 304.200 256.400 ;
        RECT 308.400 255.000 309.200 259.800 ;
        RECT 310.000 255.800 310.800 259.800 ;
        RECT 314.400 256.200 316.000 259.800 ;
        RECT 310.000 255.200 312.200 255.800 ;
        RECT 313.200 255.400 314.800 255.600 ;
        RECT 311.400 255.000 312.200 255.200 ;
        RECT 312.800 254.800 314.800 255.400 ;
        RECT 312.800 254.400 313.400 254.800 ;
        RECT 306.800 254.200 308.400 254.400 ;
        RECT 297.400 253.600 308.400 254.200 ;
        RECT 310.000 253.800 313.400 254.400 ;
        RECT 310.000 253.600 311.600 253.800 ;
        RECT 295.600 252.800 296.400 253.000 ;
        RECT 292.600 252.200 296.400 252.800 ;
        RECT 297.400 252.400 298.000 253.600 ;
        RECT 304.600 253.400 305.400 253.600 ;
        RECT 314.000 253.400 314.800 254.200 ;
        RECT 314.000 252.800 314.600 253.400 ;
        RECT 303.600 252.400 304.400 252.600 ;
        RECT 306.200 252.400 307.000 252.600 ;
        RECT 292.600 252.000 293.400 252.200 ;
        RECT 297.200 251.600 298.000 252.400 ;
        RECT 302.000 251.800 307.000 252.400 ;
        RECT 312.000 252.200 314.600 252.800 ;
        RECT 315.400 252.800 316.000 256.200 ;
        RECT 319.600 255.800 320.400 259.800 ;
        RECT 321.200 255.800 322.000 259.800 ;
        RECT 322.800 256.000 323.600 259.800 ;
        RECT 326.000 256.000 326.800 259.800 ;
        RECT 330.200 258.400 331.000 259.800 ;
        RECT 329.200 257.600 331.000 258.400 ;
        RECT 330.200 256.400 331.000 257.600 ;
        RECT 322.800 255.800 326.800 256.000 ;
        RECT 329.200 255.800 331.000 256.400 ;
        RECT 332.400 256.000 333.200 259.800 ;
        RECT 335.600 259.200 339.600 259.800 ;
        RECT 335.600 256.000 336.400 259.200 ;
        RECT 332.400 255.800 336.400 256.000 ;
        RECT 337.200 255.800 338.000 258.600 ;
        RECT 338.800 255.800 339.600 259.200 ;
        RECT 342.000 257.800 342.800 259.800 ;
        RECT 345.800 258.400 346.600 259.800 ;
        RECT 316.600 254.800 317.400 255.600 ;
        RECT 318.000 255.200 320.400 255.800 ;
        RECT 318.000 255.000 318.800 255.200 ;
        RECT 316.800 254.400 317.400 254.800 ;
        RECT 321.400 254.400 322.000 255.800 ;
        RECT 323.000 255.400 326.600 255.800 ;
        RECT 325.200 254.400 326.000 254.800 ;
        RECT 316.800 253.600 317.600 254.400 ;
        RECT 318.800 253.600 320.400 254.400 ;
        RECT 321.200 253.600 323.800 254.400 ;
        RECT 325.200 254.300 326.800 254.400 ;
        RECT 327.600 254.300 328.400 255.200 ;
        RECT 325.200 253.800 328.400 254.300 ;
        RECT 326.000 253.700 328.400 253.800 ;
        RECT 326.000 253.600 326.800 253.700 ;
        RECT 327.600 253.600 328.400 253.700 ;
        RECT 315.400 252.400 316.400 252.800 ;
        RECT 315.400 252.200 317.200 252.400 ;
        RECT 312.000 252.000 312.800 252.200 ;
        RECT 302.000 251.600 302.800 251.800 ;
        RECT 315.800 251.600 317.200 252.200 ;
        RECT 294.200 251.400 295.000 251.600 ;
        RECT 290.800 250.800 295.000 251.400 ;
        RECT 281.200 242.200 282.000 250.200 ;
        RECT 283.000 249.600 285.200 250.200 ;
        RECT 284.400 242.200 285.200 249.600 ;
        RECT 290.800 242.200 291.600 250.800 ;
        RECT 297.400 250.400 298.000 251.600 ;
        RECT 314.200 251.400 315.000 251.600 ;
        RECT 303.600 251.000 309.200 251.200 ;
        RECT 303.400 250.800 309.200 251.000 ;
        RECT 295.600 249.800 298.000 250.400 ;
        RECT 299.400 250.600 309.200 250.800 ;
        RECT 299.400 250.200 304.200 250.600 ;
        RECT 295.600 248.800 296.200 249.800 ;
        RECT 294.800 248.000 296.200 248.800 ;
        RECT 297.800 249.000 298.600 249.200 ;
        RECT 299.400 249.000 300.000 250.200 ;
        RECT 297.800 248.400 300.000 249.000 ;
        RECT 300.600 249.000 306.000 249.600 ;
        RECT 300.600 248.800 301.400 249.000 ;
        RECT 305.200 248.800 306.000 249.000 ;
        RECT 299.000 247.400 299.800 247.600 ;
        RECT 301.800 247.400 302.600 247.600 ;
        RECT 295.600 246.200 296.400 247.000 ;
        RECT 299.000 246.800 302.600 247.400 ;
        RECT 299.800 246.200 300.400 246.800 ;
        RECT 305.200 246.200 306.000 247.000 ;
        RECT 295.000 242.200 296.200 246.200 ;
        RECT 299.600 242.200 300.400 246.200 ;
        RECT 304.000 245.600 306.000 246.200 ;
        RECT 304.000 242.200 304.800 245.600 ;
        RECT 308.400 242.200 309.200 250.600 ;
        RECT 311.600 250.800 315.000 251.400 ;
        RECT 311.600 250.200 312.200 250.800 ;
        RECT 315.800 250.200 316.400 251.600 ;
        RECT 321.200 250.200 322.000 250.400 ;
        RECT 323.200 250.200 323.800 253.600 ;
        RECT 324.400 251.600 325.200 253.200 ;
        RECT 310.000 249.600 312.200 250.200 ;
        RECT 310.000 242.200 310.800 249.600 ;
        RECT 311.400 249.400 312.200 249.600 ;
        RECT 314.400 249.600 316.400 250.200 ;
        RECT 318.000 249.600 320.400 250.200 ;
        RECT 321.200 249.600 322.600 250.200 ;
        RECT 323.200 249.600 324.200 250.200 ;
        RECT 314.400 248.400 316.000 249.600 ;
        RECT 318.000 249.400 318.800 249.600 ;
        RECT 313.200 247.600 316.000 248.400 ;
        RECT 314.400 242.200 316.000 247.600 ;
        RECT 319.600 242.200 320.400 249.600 ;
        RECT 322.000 248.400 322.600 249.600 ;
        RECT 322.000 247.600 322.800 248.400 ;
        RECT 323.400 242.200 324.200 249.600 ;
        RECT 329.200 242.200 330.000 255.800 ;
        RECT 332.600 255.400 336.200 255.800 ;
        RECT 333.200 254.400 334.000 254.800 ;
        RECT 337.400 254.400 338.000 255.800 ;
        RECT 340.400 255.600 341.200 257.200 ;
        RECT 342.200 254.400 342.800 257.800 ;
        RECT 345.200 257.600 346.600 258.400 ;
        RECT 351.600 257.800 352.400 259.800 ;
        RECT 345.800 256.400 346.600 257.600 ;
        RECT 345.800 255.800 347.600 256.400 ;
        RECT 330.800 254.300 331.600 254.400 ;
        RECT 332.400 254.300 334.000 254.400 ;
        RECT 330.800 253.800 334.000 254.300 ;
        RECT 335.600 253.800 338.000 254.400 ;
        RECT 338.800 254.300 339.600 254.400 ;
        RECT 342.000 254.300 342.800 254.400 ;
        RECT 330.800 253.700 333.200 253.800 ;
        RECT 330.800 253.600 331.600 253.700 ;
        RECT 332.400 253.600 333.200 253.700 ;
        RECT 335.600 253.600 336.400 253.800 ;
        RECT 338.800 253.700 342.800 254.300 ;
        RECT 332.400 252.300 333.200 252.400 ;
        RECT 330.900 251.700 333.200 252.300 ;
        RECT 330.900 250.400 331.500 251.700 ;
        RECT 332.400 251.600 333.200 251.700 ;
        RECT 334.000 251.600 334.800 253.200 ;
        RECT 335.600 250.400 336.200 253.600 ;
        RECT 337.200 251.600 338.000 253.200 ;
        RECT 338.800 252.800 339.600 253.700 ;
        RECT 342.000 253.600 342.800 253.700 ;
        RECT 330.800 248.800 331.600 250.400 ;
        RECT 334.000 250.200 336.200 250.400 ;
        RECT 342.200 250.200 342.800 253.600 ;
        RECT 343.600 250.800 344.400 252.400 ;
        RECT 334.000 249.600 337.000 250.200 ;
        RECT 335.000 242.200 337.000 249.600 ;
        RECT 342.000 249.400 343.800 250.200 ;
        RECT 343.000 242.200 343.800 249.400 ;
        RECT 345.200 248.800 346.000 250.400 ;
        RECT 346.800 242.200 347.600 255.800 ;
        RECT 350.000 255.600 350.800 257.200 ;
        RECT 348.400 253.600 349.200 255.200 ;
        RECT 351.800 254.400 352.400 257.800 ;
        RECT 353.200 256.300 354.000 256.400 ;
        RECT 354.800 256.300 355.600 259.800 ;
        RECT 353.200 255.700 355.600 256.300 ;
        RECT 353.200 255.600 354.000 255.700 ;
        RECT 350.000 254.300 350.800 254.400 ;
        RECT 351.600 254.300 352.400 254.400 ;
        RECT 350.000 253.700 352.400 254.300 ;
        RECT 350.000 253.600 350.800 253.700 ;
        RECT 351.600 253.600 352.400 253.700 ;
        RECT 351.800 250.200 352.400 253.600 ;
        RECT 353.200 250.800 354.000 252.400 ;
        RECT 351.600 249.400 353.400 250.200 ;
        RECT 352.600 242.200 353.400 249.400 ;
        RECT 354.800 242.200 355.600 255.700 ;
        RECT 356.400 255.600 357.200 257.200 ;
        RECT 358.000 255.800 358.800 259.800 ;
        RECT 359.600 256.000 360.400 259.800 ;
        RECT 362.800 256.000 363.600 259.800 ;
        RECT 359.600 255.800 363.600 256.000 ;
        RECT 358.200 254.400 358.800 255.800 ;
        RECT 359.800 255.400 363.400 255.800 ;
        RECT 362.000 254.400 362.800 254.800 ;
        RECT 358.000 253.600 360.600 254.400 ;
        RECT 362.000 253.800 363.600 254.400 ;
        RECT 362.800 253.600 363.600 253.800 ;
        RECT 356.400 252.300 357.200 252.400 ;
        RECT 360.000 252.300 360.600 253.600 ;
        RECT 356.400 251.700 360.600 252.300 ;
        RECT 356.400 251.600 357.200 251.700 ;
        RECT 358.000 250.200 358.800 250.400 ;
        RECT 360.000 250.200 360.600 251.700 ;
        RECT 361.200 251.600 362.000 253.200 ;
        RECT 358.000 249.600 359.400 250.200 ;
        RECT 360.000 249.600 361.000 250.200 ;
        RECT 358.800 248.400 359.400 249.600 ;
        RECT 358.800 247.600 359.600 248.400 ;
        RECT 360.200 242.200 361.000 249.600 ;
        RECT 364.400 242.200 365.200 259.800 ;
        RECT 366.000 255.600 366.800 257.200 ;
        RECT 367.600 255.400 368.400 259.800 ;
        RECT 371.800 258.400 373.000 259.800 ;
        RECT 371.800 257.800 373.200 258.400 ;
        RECT 376.400 257.800 377.200 259.800 ;
        RECT 380.800 258.400 381.600 259.800 ;
        RECT 380.800 257.800 382.800 258.400 ;
        RECT 372.400 257.000 373.200 257.800 ;
        RECT 376.600 257.200 377.200 257.800 ;
        RECT 376.600 256.600 379.400 257.200 ;
        RECT 378.600 256.400 379.400 256.600 ;
        RECT 380.400 256.400 381.200 257.200 ;
        RECT 382.000 257.000 382.800 257.800 ;
        RECT 370.600 255.400 371.400 255.600 ;
        RECT 367.600 254.800 371.400 255.400 ;
        RECT 367.600 251.400 368.400 254.800 ;
        RECT 374.000 254.200 375.400 254.400 ;
        RECT 380.400 254.200 381.000 256.400 ;
        RECT 385.200 255.000 386.000 259.800 ;
        RECT 389.800 255.800 391.400 259.800 ;
        RECT 396.400 257.600 397.200 259.800 ;
        RECT 383.600 254.200 385.200 254.400 ;
        RECT 374.000 253.600 385.200 254.200 ;
        RECT 372.400 252.800 373.200 253.000 ;
        RECT 369.400 252.200 373.200 252.800 ;
        RECT 369.400 252.000 370.200 252.200 ;
        RECT 371.000 251.400 371.800 251.600 ;
        RECT 367.600 250.800 371.800 251.400 ;
        RECT 367.600 242.200 368.400 250.800 ;
        RECT 374.200 250.400 374.800 253.600 ;
        RECT 381.400 253.400 382.200 253.600 ;
        RECT 388.400 252.800 389.200 254.400 ;
        RECT 380.400 252.400 381.200 252.600 ;
        RECT 383.000 252.400 383.800 252.600 ;
        RECT 390.200 252.400 390.800 255.800 ;
        RECT 394.800 255.600 395.600 257.200 ;
        RECT 396.600 254.400 397.200 257.600 ;
        RECT 391.600 253.600 392.400 254.400 ;
        RECT 396.400 253.600 397.200 254.400 ;
        RECT 391.600 253.200 392.200 253.600 ;
        RECT 391.400 252.400 392.200 253.200 ;
        RECT 378.800 251.800 383.800 252.400 ;
        RECT 386.800 252.200 387.600 252.400 ;
        RECT 378.800 251.600 379.600 251.800 ;
        RECT 386.800 251.600 388.400 252.200 ;
        RECT 390.000 251.600 390.800 252.400 ;
        RECT 387.600 251.200 388.400 251.600 ;
        RECT 390.200 251.400 390.800 251.600 ;
        RECT 380.400 251.000 386.000 251.200 ;
        RECT 380.200 250.800 386.000 251.000 ;
        RECT 390.200 250.800 392.200 251.400 ;
        RECT 393.200 250.800 394.000 252.400 ;
        RECT 372.400 249.800 374.800 250.400 ;
        RECT 376.200 250.600 386.000 250.800 ;
        RECT 376.200 250.200 381.000 250.600 ;
        RECT 372.400 248.800 373.000 249.800 ;
        RECT 371.600 248.000 373.000 248.800 ;
        RECT 374.600 249.000 375.400 249.200 ;
        RECT 376.200 249.000 376.800 250.200 ;
        RECT 374.600 248.400 376.800 249.000 ;
        RECT 377.400 249.000 382.800 249.600 ;
        RECT 377.400 248.800 378.200 249.000 ;
        RECT 382.000 248.800 382.800 249.000 ;
        RECT 375.800 247.400 376.600 247.600 ;
        RECT 378.600 247.400 379.400 247.600 ;
        RECT 372.400 246.200 373.200 247.000 ;
        RECT 375.800 246.800 379.400 247.400 ;
        RECT 376.600 246.200 377.200 246.800 ;
        RECT 382.000 246.200 382.800 247.000 ;
        RECT 371.800 242.200 373.000 246.200 ;
        RECT 376.400 242.200 377.200 246.200 ;
        RECT 380.800 245.600 382.800 246.200 ;
        RECT 380.800 242.200 381.600 245.600 ;
        RECT 385.200 242.200 386.000 250.600 ;
        RECT 391.600 250.200 392.200 250.800 ;
        RECT 396.600 250.200 397.200 253.600 ;
        RECT 399.600 255.400 400.400 259.800 ;
        RECT 403.800 258.400 405.000 259.800 ;
        RECT 403.800 257.800 405.200 258.400 ;
        RECT 408.400 257.800 409.200 259.800 ;
        RECT 412.800 258.400 413.600 259.800 ;
        RECT 412.800 257.800 414.800 258.400 ;
        RECT 404.400 257.000 405.200 257.800 ;
        RECT 408.600 257.200 409.200 257.800 ;
        RECT 408.600 256.600 411.400 257.200 ;
        RECT 410.600 256.400 411.400 256.600 ;
        RECT 412.400 256.400 413.200 257.200 ;
        RECT 414.000 257.000 414.800 257.800 ;
        RECT 402.600 255.400 403.400 255.600 ;
        RECT 399.600 254.800 403.400 255.400 ;
        RECT 398.000 250.800 398.800 252.400 ;
        RECT 399.600 251.400 400.400 254.800 ;
        RECT 406.600 254.200 407.400 254.400 ;
        RECT 412.400 254.200 413.000 256.400 ;
        RECT 417.200 255.000 418.000 259.800 ;
        RECT 418.800 255.400 419.600 259.800 ;
        RECT 423.000 258.400 424.200 259.800 ;
        RECT 423.000 257.800 424.400 258.400 ;
        RECT 427.600 257.800 428.400 259.800 ;
        RECT 432.000 258.400 432.800 259.800 ;
        RECT 432.000 257.800 434.000 258.400 ;
        RECT 423.600 257.000 424.400 257.800 ;
        RECT 427.800 257.200 428.400 257.800 ;
        RECT 427.800 256.600 430.600 257.200 ;
        RECT 429.800 256.400 430.600 256.600 ;
        RECT 431.600 256.400 432.400 257.200 ;
        RECT 433.200 257.000 434.000 257.800 ;
        RECT 421.800 255.400 422.600 255.600 ;
        RECT 418.800 254.800 422.600 255.400 ;
        RECT 415.600 254.200 417.200 254.400 ;
        RECT 406.200 253.600 417.200 254.200 ;
        RECT 404.400 252.800 405.200 253.000 ;
        RECT 401.400 252.200 405.200 252.800 ;
        RECT 401.400 252.000 402.200 252.200 ;
        RECT 403.000 251.400 403.800 251.600 ;
        RECT 399.600 250.800 403.800 251.400 ;
        RECT 386.800 249.600 390.800 250.200 ;
        RECT 386.800 242.200 387.600 249.600 ;
        RECT 390.000 242.800 390.800 249.600 ;
        RECT 391.600 243.400 392.400 250.200 ;
        RECT 393.200 242.800 394.000 250.200 ;
        RECT 396.400 249.400 398.200 250.200 ;
        RECT 390.000 242.200 394.000 242.800 ;
        RECT 397.400 242.200 398.200 249.400 ;
        RECT 399.600 242.200 400.400 250.800 ;
        RECT 406.200 250.400 406.800 253.600 ;
        RECT 413.400 253.400 414.200 253.600 ;
        RECT 415.000 252.400 415.800 252.600 ;
        RECT 409.200 252.300 410.000 252.400 ;
        RECT 410.800 252.300 415.800 252.400 ;
        RECT 409.200 251.800 415.800 252.300 ;
        RECT 409.200 251.700 411.600 251.800 ;
        RECT 409.200 251.600 410.000 251.700 ;
        RECT 410.800 251.600 411.600 251.700 ;
        RECT 418.800 251.400 419.600 254.800 ;
        RECT 425.800 254.200 426.600 254.400 ;
        RECT 430.000 254.200 430.800 254.400 ;
        RECT 431.600 254.200 432.200 256.400 ;
        RECT 436.400 255.000 437.200 259.800 ;
        RECT 441.200 255.800 442.000 259.800 ;
        RECT 442.600 256.400 443.400 257.200 ;
        RECT 434.800 254.200 436.400 254.400 ;
        RECT 425.400 253.600 436.400 254.200 ;
        RECT 423.600 252.800 424.400 253.000 ;
        RECT 420.600 252.200 424.400 252.800 ;
        RECT 420.600 252.000 421.400 252.200 ;
        RECT 422.200 251.400 423.000 251.600 ;
        RECT 412.400 251.000 418.000 251.200 ;
        RECT 412.200 250.800 418.000 251.000 ;
        RECT 404.400 249.800 406.800 250.400 ;
        RECT 408.200 250.600 418.000 250.800 ;
        RECT 408.200 250.200 413.000 250.600 ;
        RECT 404.400 248.800 405.000 249.800 ;
        RECT 403.600 248.000 405.000 248.800 ;
        RECT 406.600 249.000 407.400 249.200 ;
        RECT 408.200 249.000 408.800 250.200 ;
        RECT 406.600 248.400 408.800 249.000 ;
        RECT 409.400 249.000 414.800 249.600 ;
        RECT 409.400 248.800 410.200 249.000 ;
        RECT 414.000 248.800 414.800 249.000 ;
        RECT 407.800 247.400 408.600 247.600 ;
        RECT 410.600 247.400 411.400 247.600 ;
        RECT 404.400 246.200 405.200 247.000 ;
        RECT 407.800 246.800 411.400 247.400 ;
        RECT 408.600 246.200 409.200 246.800 ;
        RECT 414.000 246.200 414.800 247.000 ;
        RECT 403.800 242.200 405.000 246.200 ;
        RECT 408.400 242.200 409.200 246.200 ;
        RECT 412.800 245.600 414.800 246.200 ;
        RECT 412.800 242.200 413.600 245.600 ;
        RECT 417.200 242.200 418.000 250.600 ;
        RECT 418.800 250.800 423.000 251.400 ;
        RECT 418.800 242.200 419.600 250.800 ;
        RECT 425.400 250.400 426.000 253.600 ;
        RECT 432.600 253.400 433.400 253.600 ;
        RECT 439.600 252.800 440.400 254.400 ;
        RECT 431.600 252.400 432.400 252.600 ;
        RECT 434.200 252.400 435.000 252.600 ;
        RECT 430.000 251.800 435.000 252.400 ;
        RECT 438.000 252.200 438.800 252.400 ;
        RECT 441.200 252.200 441.800 255.800 ;
        RECT 442.800 255.600 443.600 256.400 ;
        RECT 450.400 254.200 451.200 259.800 ;
        RECT 449.400 253.800 451.200 254.200 ;
        RECT 457.200 257.600 458.000 259.800 ;
        RECT 457.200 254.400 457.800 257.600 ;
        RECT 458.800 255.600 459.600 257.200 ;
        RECT 463.400 255.800 465.000 259.800 ;
        RECT 449.400 253.600 451.000 253.800 ;
        RECT 457.200 253.600 458.000 254.400 ;
        RECT 442.800 252.200 443.600 252.400 ;
        RECT 430.000 251.600 430.800 251.800 ;
        RECT 438.000 251.600 439.600 252.200 ;
        RECT 441.200 251.600 443.600 252.200 ;
        RECT 438.800 251.200 439.600 251.600 ;
        RECT 431.600 251.000 437.200 251.200 ;
        RECT 431.400 250.800 437.200 251.000 ;
        RECT 423.600 249.800 426.000 250.400 ;
        RECT 427.400 250.600 437.200 250.800 ;
        RECT 427.400 250.200 432.200 250.600 ;
        RECT 423.600 248.800 424.200 249.800 ;
        RECT 422.800 248.000 424.200 248.800 ;
        RECT 425.800 249.000 426.600 249.200 ;
        RECT 427.400 249.000 428.000 250.200 ;
        RECT 425.800 248.400 428.000 249.000 ;
        RECT 428.600 249.000 434.000 249.600 ;
        RECT 428.600 248.800 429.400 249.000 ;
        RECT 433.200 248.800 434.000 249.000 ;
        RECT 427.000 247.400 427.800 247.600 ;
        RECT 429.800 247.400 430.600 247.600 ;
        RECT 423.600 246.200 424.400 247.000 ;
        RECT 427.000 246.800 430.600 247.400 ;
        RECT 427.800 246.200 428.400 246.800 ;
        RECT 433.200 246.200 434.000 247.000 ;
        RECT 423.000 242.200 424.200 246.200 ;
        RECT 427.600 242.200 428.400 246.200 ;
        RECT 432.000 245.600 434.000 246.200 ;
        RECT 432.000 242.200 432.800 245.600 ;
        RECT 436.400 242.200 437.200 250.600 ;
        RECT 442.800 250.200 443.400 251.600 ;
        RECT 449.400 250.400 450.000 253.600 ;
        RECT 451.600 251.600 453.200 252.400 ;
        RECT 438.000 249.600 442.000 250.200 ;
        RECT 438.000 242.200 438.800 249.600 ;
        RECT 441.200 242.200 442.000 249.600 ;
        RECT 442.800 242.200 443.600 250.200 ;
        RECT 449.200 249.600 450.000 250.400 ;
        RECT 454.000 249.600 454.800 251.200 ;
        RECT 455.600 250.800 456.400 252.400 ;
        RECT 457.200 250.200 457.800 253.600 ;
        RECT 462.000 252.800 462.800 254.400 ;
        RECT 463.800 252.400 464.400 255.800 ;
        RECT 468.400 255.600 469.200 257.200 ;
        RECT 465.200 253.600 466.000 254.400 ;
        RECT 465.200 253.200 465.800 253.600 ;
        RECT 465.000 252.400 465.800 253.200 ;
        RECT 460.400 252.200 461.200 252.400 ;
        RECT 460.400 251.600 462.000 252.200 ;
        RECT 463.600 251.600 464.400 252.400 ;
        RECT 461.200 251.200 462.000 251.600 ;
        RECT 463.800 251.400 464.400 251.600 ;
        RECT 463.800 250.800 465.800 251.400 ;
        RECT 466.800 250.800 467.600 252.400 ;
        RECT 465.200 250.200 465.800 250.800 ;
        RECT 468.400 250.300 469.200 250.400 ;
        RECT 470.000 250.300 470.800 259.800 ;
        RECT 471.600 255.800 472.400 259.800 ;
        RECT 473.200 256.000 474.000 259.800 ;
        RECT 476.400 256.000 477.200 259.800 ;
        RECT 473.200 255.800 477.200 256.000 ;
        RECT 478.600 256.400 479.400 259.800 ;
        RECT 478.600 255.800 480.400 256.400 ;
        RECT 482.800 255.800 483.600 259.800 ;
        RECT 484.400 256.000 485.200 259.800 ;
        RECT 487.600 256.000 488.400 259.800 ;
        RECT 484.400 255.800 488.400 256.000 ;
        RECT 489.800 258.400 490.600 259.800 ;
        RECT 489.800 257.600 491.600 258.400 ;
        RECT 495.600 257.800 496.400 259.800 ;
        RECT 489.800 256.400 490.600 257.600 ;
        RECT 489.800 255.800 491.600 256.400 ;
        RECT 471.800 254.400 472.400 255.800 ;
        RECT 473.400 255.400 477.000 255.800 ;
        RECT 475.600 254.400 476.400 254.800 ;
        RECT 471.600 253.600 474.200 254.400 ;
        RECT 475.600 254.300 477.200 254.400 ;
        RECT 479.600 254.300 480.400 255.800 ;
        RECT 475.600 253.800 480.400 254.300 ;
        RECT 476.400 253.700 480.400 253.800 ;
        RECT 476.400 253.600 477.200 253.700 ;
        RECT 471.600 252.300 472.400 252.400 ;
        RECT 473.600 252.300 474.200 253.600 ;
        RECT 471.600 251.700 474.200 252.300 ;
        RECT 471.600 251.600 472.400 251.700 ;
        RECT 471.600 250.300 472.400 250.400 ;
        RECT 468.400 250.200 472.400 250.300 ;
        RECT 473.600 250.200 474.200 251.700 ;
        RECT 474.800 251.600 475.600 253.200 ;
        RECT 449.400 247.000 450.000 249.600 ;
        RECT 456.200 249.400 458.000 250.200 ;
        RECT 460.400 249.600 464.400 250.200 ;
        RECT 450.800 247.600 451.600 249.200 ;
        RECT 449.400 246.400 453.000 247.000 ;
        RECT 449.400 246.200 450.000 246.400 ;
        RECT 449.200 242.200 450.000 246.200 ;
        RECT 452.400 242.200 453.200 246.400 ;
        RECT 456.200 242.200 457.000 249.400 ;
        RECT 460.400 242.200 461.200 249.600 ;
        RECT 463.600 242.800 464.400 249.600 ;
        RECT 465.200 243.400 466.000 250.200 ;
        RECT 466.800 242.800 467.600 250.200 ;
        RECT 468.400 249.700 473.000 250.200 ;
        RECT 468.400 249.600 469.200 249.700 ;
        RECT 463.600 242.200 467.600 242.800 ;
        RECT 470.000 242.200 470.800 249.700 ;
        RECT 471.600 249.600 473.000 249.700 ;
        RECT 473.600 249.600 474.600 250.200 ;
        RECT 472.400 248.400 473.000 249.600 ;
        RECT 472.400 247.600 473.200 248.400 ;
        RECT 473.800 242.200 474.600 249.600 ;
        RECT 478.000 248.800 478.800 250.400 ;
        RECT 479.600 242.200 480.400 253.700 ;
        RECT 481.200 253.600 482.000 255.200 ;
        RECT 483.000 254.400 483.600 255.800 ;
        RECT 484.600 255.400 488.200 255.800 ;
        RECT 486.800 254.400 487.600 254.800 ;
        RECT 482.800 253.600 485.400 254.400 ;
        RECT 486.800 253.800 488.400 254.400 ;
        RECT 487.600 253.600 488.400 253.800 ;
        RECT 484.800 250.400 485.400 253.600 ;
        RECT 486.000 251.600 486.800 253.200 ;
        RECT 482.800 250.200 483.600 250.400 ;
        RECT 482.800 249.600 484.200 250.200 ;
        RECT 484.800 249.600 486.800 250.400 ;
        RECT 483.600 248.400 484.200 249.600 ;
        RECT 483.600 247.600 484.400 248.400 ;
        RECT 485.000 242.200 485.800 249.600 ;
        RECT 489.200 248.800 490.000 250.400 ;
        RECT 490.800 242.200 491.600 255.800 ;
        RECT 494.000 255.600 494.800 257.200 ;
        RECT 495.800 256.300 496.400 257.800 ;
        RECT 500.400 257.800 501.200 259.800 ;
        RECT 498.800 256.300 499.600 256.400 ;
        RECT 495.700 255.700 499.600 256.300 ;
        RECT 492.400 254.300 493.200 255.200 ;
        RECT 494.100 254.300 494.700 255.600 ;
        RECT 495.800 254.400 496.400 255.700 ;
        RECT 498.800 255.600 499.600 255.700 ;
        RECT 492.400 253.700 494.700 254.300 ;
        RECT 492.400 253.600 493.200 253.700 ;
        RECT 495.600 253.600 496.400 254.400 ;
        RECT 495.800 250.200 496.400 253.600 ;
        RECT 500.400 254.400 501.000 257.800 ;
        RECT 502.000 255.600 502.800 257.200 ;
        RECT 503.600 255.800 504.400 259.800 ;
        RECT 508.000 258.400 509.600 259.800 ;
        RECT 508.000 257.600 510.800 258.400 ;
        RECT 508.000 256.200 509.600 257.600 ;
        RECT 503.600 255.200 506.000 255.800 ;
        RECT 505.200 255.000 506.000 255.200 ;
        RECT 506.600 254.800 507.400 255.600 ;
        RECT 506.600 254.400 507.200 254.800 ;
        RECT 500.400 254.300 501.200 254.400 ;
        RECT 502.000 254.300 502.800 254.400 ;
        RECT 500.400 253.700 502.800 254.300 ;
        RECT 500.400 253.600 501.200 253.700 ;
        RECT 502.000 253.600 502.800 253.700 ;
        RECT 503.600 253.600 505.200 254.400 ;
        RECT 506.400 253.600 507.200 254.400 ;
        RECT 508.000 254.200 508.600 256.200 ;
        RECT 513.200 255.800 514.000 259.800 ;
        RECT 509.200 254.800 510.800 255.600 ;
        RECT 511.400 255.200 514.000 255.800 ;
        RECT 514.800 255.800 515.600 259.800 ;
        RECT 519.200 258.400 520.800 259.800 ;
        RECT 519.200 257.600 522.000 258.400 ;
        RECT 519.200 256.200 520.800 257.600 ;
        RECT 514.800 255.200 517.400 255.800 ;
        RECT 511.400 255.000 512.200 255.200 ;
        RECT 516.600 255.000 517.400 255.200 ;
        RECT 518.000 254.800 519.600 255.600 ;
        RECT 512.400 254.200 514.000 254.400 ;
        RECT 508.000 253.600 509.000 254.200 ;
        RECT 511.800 254.000 514.000 254.200 ;
        RECT 497.200 250.800 498.000 252.400 ;
        RECT 498.800 250.800 499.600 252.400 ;
        RECT 500.400 250.200 501.000 253.600 ;
        RECT 502.000 252.300 502.800 252.400 ;
        RECT 503.700 252.300 504.300 253.600 ;
        RECT 502.000 251.700 504.300 252.300 ;
        RECT 508.400 252.400 509.000 253.600 ;
        RECT 509.600 253.600 514.000 254.000 ;
        RECT 514.800 254.200 516.400 254.400 ;
        RECT 520.200 254.200 520.800 256.200 ;
        RECT 524.400 255.800 525.200 259.800 ;
        RECT 521.400 254.800 522.200 255.600 ;
        RECT 522.800 255.200 525.200 255.800 ;
        RECT 526.000 255.800 526.800 259.800 ;
        RECT 530.400 258.400 532.000 259.800 ;
        RECT 530.400 257.600 533.200 258.400 ;
        RECT 530.400 256.200 532.000 257.600 ;
        RECT 526.000 255.200 528.400 255.800 ;
        RECT 522.800 255.000 523.600 255.200 ;
        RECT 527.600 255.000 528.400 255.200 ;
        RECT 514.800 254.000 517.000 254.200 ;
        RECT 514.800 253.600 519.200 254.000 ;
        RECT 509.600 253.400 512.400 253.600 ;
        RECT 516.400 253.400 519.200 253.600 ;
        RECT 509.600 253.200 510.400 253.400 ;
        RECT 518.400 253.200 519.200 253.400 ;
        RECT 519.800 253.600 520.800 254.200 ;
        RECT 521.600 254.400 522.200 254.800 ;
        RECT 529.000 254.800 529.800 255.600 ;
        RECT 529.000 254.400 529.600 254.800 ;
        RECT 521.600 253.600 522.400 254.400 ;
        RECT 523.600 254.300 525.200 254.400 ;
        RECT 526.000 254.300 527.600 254.400 ;
        RECT 523.600 253.700 527.600 254.300 ;
        RECT 523.600 253.600 525.200 253.700 ;
        RECT 526.000 253.600 527.600 253.700 ;
        RECT 528.800 253.600 529.600 254.400 ;
        RECT 519.800 252.400 520.400 253.600 ;
        RECT 530.400 252.800 531.000 256.200 ;
        RECT 535.600 255.800 536.400 259.800 ;
        RECT 531.600 255.400 533.200 255.600 ;
        RECT 531.600 254.800 533.600 255.400 ;
        RECT 534.200 255.200 536.400 255.800 ;
        RECT 534.200 255.000 535.000 255.200 ;
        RECT 537.200 255.000 538.000 259.800 ;
        RECT 541.600 258.400 542.400 259.800 ;
        RECT 540.400 257.800 542.400 258.400 ;
        RECT 546.000 257.800 546.800 259.800 ;
        RECT 550.200 258.400 551.400 259.800 ;
        RECT 550.000 257.800 551.400 258.400 ;
        RECT 540.400 257.000 541.200 257.800 ;
        RECT 546.000 257.200 546.600 257.800 ;
        RECT 542.000 256.400 542.800 257.200 ;
        RECT 543.800 256.600 546.600 257.200 ;
        RECT 550.000 257.000 550.800 257.800 ;
        RECT 543.800 256.400 544.600 256.600 ;
        RECT 533.000 254.400 533.600 254.800 ;
        RECT 531.600 253.400 532.400 254.200 ;
        RECT 533.000 253.800 536.400 254.400 ;
        RECT 534.800 253.600 536.400 253.800 ;
        RECT 538.000 254.200 539.600 254.400 ;
        RECT 542.200 254.200 542.800 256.400 ;
        RECT 551.800 255.400 552.600 255.600 ;
        RECT 554.800 255.400 555.600 259.800 ;
        RECT 551.800 254.800 555.600 255.400 ;
        RECT 543.600 254.200 544.400 254.400 ;
        RECT 547.800 254.200 548.600 254.400 ;
        RECT 538.000 253.600 549.000 254.200 ;
        RECT 541.000 253.400 541.800 253.600 ;
        RECT 530.000 252.400 531.000 252.800 ;
        RECT 502.000 251.600 502.800 251.700 ;
        RECT 508.400 251.600 509.200 252.400 ;
        RECT 511.000 252.200 511.800 252.400 ;
        RECT 510.200 251.600 511.800 252.200 ;
        RECT 517.000 252.200 517.800 252.400 ;
        RECT 517.000 251.600 518.600 252.200 ;
        RECT 519.600 251.600 520.400 252.400 ;
        RECT 529.200 252.200 531.000 252.400 ;
        RECT 531.800 252.800 532.400 253.400 ;
        RECT 531.800 252.200 534.400 252.800 ;
        RECT 529.200 251.600 530.600 252.200 ;
        RECT 533.600 252.000 534.400 252.200 ;
        RECT 539.400 252.400 540.200 252.600 ;
        RECT 542.000 252.400 542.800 252.600 ;
        RECT 539.400 251.800 544.400 252.400 ;
        RECT 543.600 251.600 544.400 251.800 ;
        RECT 508.400 250.200 509.000 251.600 ;
        RECT 510.200 251.400 511.000 251.600 ;
        RECT 517.800 251.400 518.600 251.600 ;
        RECT 519.800 250.200 520.400 251.600 ;
        RECT 530.000 250.200 530.600 251.600 ;
        RECT 531.400 251.400 532.200 251.600 ;
        RECT 531.400 250.800 534.800 251.400 ;
        RECT 534.200 250.200 534.800 250.800 ;
        RECT 537.200 251.000 542.800 251.200 ;
        RECT 537.200 250.800 543.000 251.000 ;
        RECT 537.200 250.600 547.000 250.800 ;
        RECT 495.600 249.400 497.400 250.200 ;
        RECT 496.600 242.200 497.400 249.400 ;
        RECT 499.400 249.400 501.200 250.200 ;
        RECT 503.600 249.600 506.000 250.200 ;
        RECT 499.400 242.200 500.200 249.400 ;
        RECT 503.600 242.200 504.400 249.600 ;
        RECT 505.200 249.400 506.000 249.600 ;
        RECT 508.000 242.200 509.600 250.200 ;
        RECT 511.400 249.600 514.000 250.200 ;
        RECT 511.400 249.400 512.200 249.600 ;
        RECT 513.200 242.200 514.000 249.600 ;
        RECT 514.800 249.600 517.400 250.200 ;
        RECT 514.800 242.200 515.600 249.600 ;
        RECT 516.600 249.400 517.400 249.600 ;
        RECT 519.200 242.200 520.800 250.200 ;
        RECT 522.800 249.600 525.200 250.200 ;
        RECT 522.800 249.400 523.600 249.600 ;
        RECT 524.400 242.200 525.200 249.600 ;
        RECT 526.000 249.600 528.400 250.200 ;
        RECT 530.000 249.600 532.000 250.200 ;
        RECT 526.000 242.200 526.800 249.600 ;
        RECT 527.600 249.400 528.400 249.600 ;
        RECT 530.400 242.200 532.000 249.600 ;
        RECT 534.200 249.600 536.400 250.200 ;
        RECT 534.200 249.400 535.000 249.600 ;
        RECT 535.600 242.200 536.400 249.600 ;
        RECT 537.200 242.200 538.000 250.600 ;
        RECT 542.200 250.200 547.000 250.600 ;
        RECT 540.400 249.000 545.800 249.600 ;
        RECT 540.400 248.800 541.200 249.000 ;
        RECT 545.000 248.800 545.800 249.000 ;
        RECT 546.400 249.000 547.000 250.200 ;
        RECT 548.400 250.400 549.000 253.600 ;
        RECT 550.000 252.800 550.800 253.000 ;
        RECT 550.000 252.200 553.800 252.800 ;
        RECT 553.000 252.000 553.800 252.200 ;
        RECT 551.400 251.400 552.200 251.600 ;
        RECT 554.800 251.400 555.600 254.800 ;
        RECT 556.400 255.200 557.200 259.800 ;
        RECT 556.400 254.600 558.600 255.200 ;
        RECT 561.200 255.000 562.000 259.800 ;
        RECT 565.600 258.400 566.400 259.800 ;
        RECT 564.400 257.800 566.400 258.400 ;
        RECT 570.000 257.800 570.800 259.800 ;
        RECT 574.200 258.400 575.400 259.800 ;
        RECT 574.000 257.800 575.400 258.400 ;
        RECT 564.400 257.000 565.200 257.800 ;
        RECT 570.000 257.200 570.600 257.800 ;
        RECT 566.000 256.400 566.800 257.200 ;
        RECT 567.800 256.600 570.600 257.200 ;
        RECT 574.000 257.000 574.800 257.800 ;
        RECT 567.800 256.400 568.600 256.600 ;
        RECT 556.400 251.600 557.200 253.200 ;
        RECT 558.000 251.600 558.600 254.600 ;
        RECT 562.000 254.200 563.600 254.400 ;
        RECT 566.200 254.200 566.800 256.400 ;
        RECT 575.800 255.400 576.600 255.600 ;
        RECT 578.800 255.400 579.600 259.800 ;
        RECT 575.800 254.800 579.600 255.400 ;
        RECT 571.800 254.200 572.600 254.400 ;
        RECT 562.000 253.600 573.000 254.200 ;
        RECT 565.000 253.400 565.800 253.600 ;
        RECT 563.400 252.400 564.200 252.600 ;
        RECT 566.000 252.400 566.800 252.600 ;
        RECT 563.400 251.800 568.400 252.400 ;
        RECT 567.600 251.600 568.400 251.800 ;
        RECT 551.400 250.800 555.600 251.400 ;
        RECT 548.400 249.800 550.800 250.400 ;
        RECT 547.800 249.000 548.600 249.200 ;
        RECT 546.400 248.400 548.600 249.000 ;
        RECT 550.200 248.800 550.800 249.800 ;
        RECT 550.200 248.000 551.600 248.800 ;
        RECT 543.800 247.400 544.600 247.600 ;
        RECT 546.600 247.400 547.400 247.600 ;
        RECT 540.400 246.200 541.200 247.000 ;
        RECT 543.800 246.800 547.400 247.400 ;
        RECT 546.000 246.200 546.600 246.800 ;
        RECT 550.000 246.200 550.800 247.000 ;
        RECT 540.400 245.600 542.400 246.200 ;
        RECT 541.600 242.200 542.400 245.600 ;
        RECT 546.000 242.200 546.800 246.200 ;
        RECT 550.200 242.200 551.400 246.200 ;
        RECT 554.800 242.200 555.600 250.800 ;
        RECT 558.000 250.800 559.200 251.600 ;
        RECT 561.200 251.000 566.800 251.200 ;
        RECT 561.200 250.800 567.000 251.000 ;
        RECT 558.000 250.200 558.600 250.800 ;
        RECT 556.400 249.600 558.600 250.200 ;
        RECT 561.200 250.600 571.000 250.800 ;
        RECT 556.400 242.200 557.200 249.600 ;
        RECT 561.200 242.200 562.000 250.600 ;
        RECT 566.200 250.200 571.000 250.600 ;
        RECT 564.400 249.000 569.800 249.600 ;
        RECT 564.400 248.800 565.200 249.000 ;
        RECT 569.000 248.800 569.800 249.000 ;
        RECT 570.400 249.000 571.000 250.200 ;
        RECT 572.400 250.400 573.000 253.600 ;
        RECT 574.000 252.800 574.800 253.000 ;
        RECT 574.000 252.200 577.800 252.800 ;
        RECT 577.000 252.000 577.800 252.200 ;
        RECT 575.400 251.400 576.200 251.600 ;
        RECT 578.800 251.400 579.600 254.800 ;
        RECT 580.400 255.200 581.200 259.800 ;
        RECT 580.400 254.600 582.600 255.200 ;
        RECT 580.400 251.600 581.200 253.200 ;
        RECT 582.000 251.600 582.600 254.600 ;
        RECT 575.400 250.800 579.600 251.400 ;
        RECT 572.400 249.800 574.800 250.400 ;
        RECT 571.800 249.000 572.600 249.200 ;
        RECT 570.400 248.400 572.600 249.000 ;
        RECT 574.200 248.800 574.800 249.800 ;
        RECT 574.200 248.000 575.600 248.800 ;
        RECT 567.800 247.400 568.600 247.600 ;
        RECT 570.600 247.400 571.400 247.600 ;
        RECT 564.400 246.200 565.200 247.000 ;
        RECT 567.800 246.800 571.400 247.400 ;
        RECT 570.000 246.200 570.600 246.800 ;
        RECT 574.000 246.200 574.800 247.000 ;
        RECT 564.400 245.600 566.400 246.200 ;
        RECT 565.600 242.200 566.400 245.600 ;
        RECT 570.000 242.200 570.800 246.200 ;
        RECT 574.200 242.200 575.400 246.200 ;
        RECT 578.800 242.200 579.600 250.800 ;
        RECT 582.000 250.800 583.200 251.600 ;
        RECT 582.000 250.200 582.600 250.800 ;
        RECT 580.400 249.600 582.600 250.200 ;
        RECT 580.400 242.200 581.200 249.600 ;
        RECT 1.200 231.200 2.000 239.800 ;
        RECT 5.400 235.800 6.600 239.800 ;
        RECT 10.000 235.800 10.800 239.800 ;
        RECT 14.400 236.400 15.200 239.800 ;
        RECT 14.400 235.800 16.400 236.400 ;
        RECT 6.000 235.000 6.800 235.800 ;
        RECT 10.200 235.200 10.800 235.800 ;
        RECT 9.400 234.600 13.000 235.200 ;
        RECT 15.600 235.000 16.400 235.800 ;
        RECT 9.400 234.400 10.200 234.600 ;
        RECT 12.200 234.400 13.000 234.600 ;
        RECT 5.200 233.200 6.600 234.000 ;
        RECT 6.000 232.200 6.600 233.200 ;
        RECT 8.200 233.000 10.400 233.600 ;
        RECT 8.200 232.800 9.000 233.000 ;
        RECT 6.000 231.600 8.400 232.200 ;
        RECT 1.200 230.600 5.400 231.200 ;
        RECT 1.200 227.200 2.000 230.600 ;
        RECT 4.600 230.400 5.400 230.600 ;
        RECT 3.000 229.800 3.800 230.000 ;
        RECT 3.000 229.200 6.800 229.800 ;
        RECT 6.000 229.000 6.800 229.200 ;
        RECT 7.800 228.400 8.400 231.600 ;
        RECT 9.800 231.800 10.400 233.000 ;
        RECT 11.000 233.000 11.800 233.200 ;
        RECT 15.600 233.000 16.400 233.200 ;
        RECT 11.000 232.400 16.400 233.000 ;
        RECT 9.800 231.400 14.600 231.800 ;
        RECT 18.800 231.400 19.600 239.800 ;
        RECT 20.400 232.400 21.200 239.800 ;
        RECT 22.000 232.400 22.800 232.600 ;
        RECT 24.800 232.400 26.400 239.800 ;
        RECT 20.400 231.800 22.800 232.400 ;
        RECT 24.400 231.800 26.400 232.400 ;
        RECT 28.600 232.400 29.400 232.600 ;
        RECT 30.000 232.400 30.800 239.800 ;
        RECT 28.600 231.800 30.800 232.400 ;
        RECT 31.600 232.400 32.400 239.800 ;
        RECT 33.200 232.400 34.000 232.600 ;
        RECT 36.000 232.400 37.600 239.800 ;
        RECT 31.600 231.800 34.000 232.400 ;
        RECT 35.600 231.800 37.600 232.400 ;
        RECT 39.800 232.400 40.600 232.600 ;
        RECT 41.200 232.400 42.000 239.800 ;
        RECT 39.800 231.800 42.000 232.400 ;
        RECT 9.800 231.200 19.600 231.400 ;
        RECT 13.800 231.000 19.600 231.200 ;
        RECT 14.000 230.800 19.600 231.000 ;
        RECT 24.400 230.400 25.000 231.800 ;
        RECT 28.600 231.200 29.200 231.800 ;
        RECT 25.800 230.600 29.200 231.200 ;
        RECT 25.800 230.400 26.600 230.600 ;
        RECT 35.600 230.400 36.200 231.800 ;
        RECT 39.800 231.200 40.400 231.800 ;
        RECT 37.000 230.600 40.400 231.200 ;
        RECT 42.800 231.200 43.600 239.800 ;
        RECT 47.000 235.800 48.200 239.800 ;
        RECT 51.600 235.800 52.400 239.800 ;
        RECT 56.000 236.400 56.800 239.800 ;
        RECT 56.000 235.800 58.000 236.400 ;
        RECT 47.600 235.000 48.400 235.800 ;
        RECT 51.800 235.200 52.400 235.800 ;
        RECT 51.000 234.600 54.600 235.200 ;
        RECT 57.200 235.000 58.000 235.800 ;
        RECT 51.000 234.400 51.800 234.600 ;
        RECT 53.800 234.400 54.600 234.600 ;
        RECT 46.800 233.200 48.200 234.000 ;
        RECT 47.600 232.200 48.200 233.200 ;
        RECT 49.800 233.000 52.000 233.600 ;
        RECT 49.800 232.800 50.600 233.000 ;
        RECT 47.600 231.600 50.000 232.200 ;
        RECT 42.800 230.600 47.000 231.200 ;
        RECT 37.000 230.400 37.800 230.600 ;
        RECT 12.400 230.200 13.200 230.400 ;
        RECT 12.400 229.600 17.400 230.200 ;
        RECT 23.600 229.800 25.000 230.400 ;
        RECT 28.000 229.800 28.800 230.000 ;
        RECT 23.600 229.600 25.400 229.800 ;
        RECT 14.000 229.400 14.800 229.600 ;
        RECT 16.600 229.400 17.400 229.600 ;
        RECT 24.400 229.200 25.400 229.600 ;
        RECT 15.000 228.400 15.800 228.600 ;
        RECT 7.800 227.800 18.800 228.400 ;
        RECT 8.200 227.600 9.000 227.800 ;
        RECT 12.400 227.600 13.200 227.800 ;
        RECT 1.200 226.600 5.000 227.200 ;
        RECT 1.200 222.200 2.000 226.600 ;
        RECT 4.200 226.400 5.000 226.600 ;
        RECT 14.000 225.600 14.600 227.800 ;
        RECT 17.200 227.600 18.800 227.800 ;
        RECT 20.400 227.600 22.000 228.400 ;
        RECT 23.200 227.600 24.000 228.400 ;
        RECT 23.400 227.200 24.000 227.600 ;
        RECT 12.200 225.400 13.000 225.600 ;
        RECT 6.000 224.200 6.800 225.000 ;
        RECT 10.200 224.800 13.000 225.400 ;
        RECT 14.000 224.800 14.800 225.600 ;
        RECT 10.200 224.200 10.800 224.800 ;
        RECT 15.600 224.200 16.400 225.000 ;
        RECT 5.400 223.600 6.800 224.200 ;
        RECT 5.400 222.200 6.600 223.600 ;
        RECT 10.000 222.200 10.800 224.200 ;
        RECT 14.400 223.600 16.400 224.200 ;
        RECT 14.400 222.200 15.200 223.600 ;
        RECT 18.800 222.200 19.600 227.000 ;
        RECT 22.000 226.800 22.800 227.000 ;
        RECT 20.400 226.200 22.800 226.800 ;
        RECT 23.400 226.400 24.200 227.200 ;
        RECT 20.400 222.200 21.200 226.200 ;
        RECT 24.800 225.800 25.400 229.200 ;
        RECT 26.200 229.200 28.800 229.800 ;
        RECT 34.800 229.800 36.200 230.400 ;
        RECT 39.200 229.800 40.000 230.000 ;
        RECT 34.800 229.600 36.600 229.800 ;
        RECT 35.600 229.200 36.600 229.600 ;
        RECT 26.200 228.600 26.800 229.200 ;
        RECT 26.000 227.800 26.800 228.600 ;
        RECT 29.200 228.200 30.800 228.400 ;
        RECT 27.400 227.600 30.800 228.200 ;
        RECT 31.600 227.600 33.200 228.400 ;
        RECT 34.400 227.600 35.200 228.400 ;
        RECT 27.400 227.200 28.000 227.600 ;
        RECT 26.000 226.600 28.000 227.200 ;
        RECT 34.600 227.200 35.200 227.600 ;
        RECT 28.600 226.800 29.400 227.000 ;
        RECT 33.200 226.800 34.000 227.000 ;
        RECT 26.000 226.400 27.600 226.600 ;
        RECT 28.600 226.200 30.800 226.800 ;
        RECT 24.800 222.200 26.400 225.800 ;
        RECT 30.000 222.200 30.800 226.200 ;
        RECT 31.600 226.200 34.000 226.800 ;
        RECT 34.600 226.400 35.400 227.200 ;
        RECT 31.600 222.200 32.400 226.200 ;
        RECT 36.000 225.800 36.600 229.200 ;
        RECT 37.400 229.200 40.000 229.800 ;
        RECT 37.400 228.600 38.000 229.200 ;
        RECT 37.200 227.800 38.000 228.600 ;
        RECT 40.400 228.200 42.000 228.400 ;
        RECT 38.600 227.600 42.000 228.200 ;
        RECT 38.600 227.200 39.200 227.600 ;
        RECT 37.200 226.600 39.200 227.200 ;
        RECT 42.800 227.200 43.600 230.600 ;
        RECT 46.200 230.400 47.000 230.600 ;
        RECT 44.600 229.800 45.400 230.000 ;
        RECT 44.600 229.200 48.400 229.800 ;
        RECT 47.600 229.000 48.400 229.200 ;
        RECT 49.400 228.400 50.000 231.600 ;
        RECT 51.400 231.800 52.000 233.000 ;
        RECT 52.600 233.000 53.400 233.200 ;
        RECT 57.200 233.000 58.000 233.200 ;
        RECT 52.600 232.400 58.000 233.000 ;
        RECT 51.400 231.400 56.200 231.800 ;
        RECT 60.400 231.400 61.200 239.800 ;
        RECT 51.400 231.200 61.200 231.400 ;
        RECT 55.400 231.000 61.200 231.200 ;
        RECT 55.600 230.800 61.200 231.000 ;
        RECT 62.000 231.400 62.800 239.800 ;
        RECT 66.400 236.400 67.200 239.800 ;
        RECT 65.200 235.800 67.200 236.400 ;
        RECT 70.800 235.800 71.600 239.800 ;
        RECT 75.000 235.800 76.200 239.800 ;
        RECT 65.200 235.000 66.000 235.800 ;
        RECT 70.800 235.200 71.400 235.800 ;
        RECT 68.600 234.600 72.200 235.200 ;
        RECT 74.800 235.000 75.600 235.800 ;
        RECT 68.600 234.400 69.400 234.600 ;
        RECT 71.400 234.400 72.200 234.600 ;
        RECT 65.200 233.000 66.000 233.200 ;
        RECT 69.800 233.000 70.600 233.200 ;
        RECT 65.200 232.400 70.600 233.000 ;
        RECT 71.200 233.000 73.400 233.600 ;
        RECT 71.200 231.800 71.800 233.000 ;
        RECT 72.600 232.800 73.400 233.000 ;
        RECT 75.000 233.200 76.400 234.000 ;
        RECT 75.000 232.200 75.600 233.200 ;
        RECT 67.000 231.400 71.800 231.800 ;
        RECT 62.000 231.200 71.800 231.400 ;
        RECT 73.200 231.600 75.600 232.200 ;
        RECT 62.000 231.000 67.800 231.200 ;
        RECT 62.000 230.800 67.600 231.000 ;
        RECT 54.000 230.200 54.800 230.400 ;
        RECT 68.400 230.200 69.200 230.400 ;
        RECT 54.000 229.600 59.000 230.200 ;
        RECT 55.600 229.400 56.400 229.600 ;
        RECT 58.200 229.400 59.000 229.600 ;
        RECT 64.200 229.600 69.200 230.200 ;
        RECT 64.200 229.400 65.000 229.600 ;
        RECT 66.800 229.400 67.600 229.600 ;
        RECT 56.600 228.400 57.400 228.600 ;
        RECT 65.800 228.400 66.600 228.600 ;
        RECT 73.200 228.400 73.800 231.600 ;
        RECT 79.600 231.200 80.400 239.800 ;
        RECT 81.200 232.400 82.000 239.800 ;
        RECT 85.600 234.400 87.200 239.800 ;
        RECT 84.400 233.600 87.200 234.400 ;
        RECT 82.600 232.400 83.400 232.600 ;
        RECT 81.200 231.800 83.400 232.400 ;
        RECT 85.600 232.400 87.200 233.600 ;
        RECT 89.200 232.400 90.000 232.600 ;
        RECT 90.800 232.400 91.600 239.800 ;
        RECT 85.600 231.800 87.600 232.400 ;
        RECT 89.200 231.800 91.600 232.400 ;
        RECT 76.200 230.600 80.400 231.200 ;
        RECT 82.800 231.200 83.400 231.800 ;
        RECT 82.800 230.600 86.200 231.200 ;
        RECT 76.200 230.400 77.000 230.600 ;
        RECT 77.800 229.800 78.600 230.000 ;
        RECT 74.800 229.200 78.600 229.800 ;
        RECT 74.800 229.000 75.600 229.200 ;
        RECT 49.400 227.800 60.400 228.400 ;
        RECT 49.800 227.600 50.600 227.800 ;
        RECT 39.800 226.800 40.600 227.000 ;
        RECT 37.200 226.400 38.800 226.600 ;
        RECT 39.800 226.200 42.000 226.800 ;
        RECT 36.000 224.400 37.600 225.800 ;
        RECT 34.800 223.600 37.600 224.400 ;
        RECT 36.000 222.200 37.600 223.600 ;
        RECT 41.200 222.200 42.000 226.200 ;
        RECT 42.800 226.600 46.600 227.200 ;
        RECT 42.800 222.200 43.600 226.600 ;
        RECT 45.800 226.400 46.600 226.600 ;
        RECT 55.600 226.400 56.200 227.800 ;
        RECT 58.800 227.600 60.400 227.800 ;
        RECT 62.800 227.800 73.800 228.400 ;
        RECT 62.800 227.600 64.400 227.800 ;
        RECT 53.800 225.400 54.600 225.600 ;
        RECT 47.600 224.200 48.400 225.000 ;
        RECT 51.800 224.800 54.600 225.400 ;
        RECT 55.600 224.800 56.400 226.400 ;
        RECT 51.800 224.200 52.400 224.800 ;
        RECT 57.200 224.200 58.000 225.000 ;
        RECT 47.000 223.600 48.400 224.200 ;
        RECT 47.000 222.200 48.200 223.600 ;
        RECT 51.600 222.200 52.400 224.200 ;
        RECT 56.000 223.600 58.000 224.200 ;
        RECT 56.000 222.200 56.800 223.600 ;
        RECT 60.400 222.200 61.200 227.000 ;
        RECT 62.000 222.200 62.800 227.000 ;
        RECT 67.000 225.600 67.600 227.800 ;
        RECT 70.000 227.600 70.800 227.800 ;
        RECT 72.600 227.600 73.400 227.800 ;
        RECT 79.600 227.200 80.400 230.600 ;
        RECT 85.400 230.400 86.200 230.600 ;
        RECT 87.000 230.400 87.600 231.800 ;
        RECT 92.400 231.600 93.200 233.200 ;
        RECT 83.200 229.800 84.000 230.000 ;
        RECT 87.000 229.800 88.400 230.400 ;
        RECT 83.200 229.200 85.800 229.800 ;
        RECT 85.200 228.600 85.800 229.200 ;
        RECT 86.600 229.600 88.400 229.800 ;
        RECT 86.600 229.200 87.600 229.600 ;
        RECT 81.200 228.200 82.800 228.400 ;
        RECT 81.200 227.600 84.600 228.200 ;
        RECT 85.200 227.800 86.000 228.600 ;
        RECT 76.600 226.600 80.400 227.200 ;
        RECT 84.000 227.200 84.600 227.600 ;
        RECT 82.600 226.800 83.400 227.000 ;
        RECT 76.600 226.400 77.400 226.600 ;
        RECT 65.200 224.200 66.000 225.000 ;
        RECT 66.800 224.800 67.600 225.600 ;
        RECT 68.600 225.400 69.400 225.600 ;
        RECT 68.600 224.800 71.400 225.400 ;
        RECT 70.800 224.200 71.400 224.800 ;
        RECT 74.800 224.200 75.600 225.000 ;
        RECT 65.200 223.600 67.200 224.200 ;
        RECT 66.400 222.200 67.200 223.600 ;
        RECT 70.800 222.200 71.600 224.200 ;
        RECT 74.800 223.600 76.200 224.200 ;
        RECT 75.000 222.200 76.200 223.600 ;
        RECT 79.600 222.200 80.400 226.600 ;
        RECT 81.200 226.200 83.400 226.800 ;
        RECT 84.000 226.600 86.000 227.200 ;
        RECT 84.400 226.400 86.000 226.600 ;
        RECT 81.200 222.200 82.000 226.200 ;
        RECT 86.600 225.800 87.200 229.200 ;
        RECT 88.000 227.600 88.800 228.400 ;
        RECT 90.000 227.600 91.600 228.400 ;
        RECT 88.000 227.200 88.600 227.600 ;
        RECT 87.800 226.400 88.600 227.200 ;
        RECT 89.200 226.800 90.000 227.000 ;
        RECT 89.200 226.200 91.600 226.800 ;
        RECT 94.000 226.200 94.800 239.800 ;
        RECT 97.200 231.200 98.000 239.800 ;
        RECT 101.400 235.800 102.600 239.800 ;
        RECT 106.000 235.800 106.800 239.800 ;
        RECT 110.400 236.400 111.200 239.800 ;
        RECT 110.400 235.800 112.400 236.400 ;
        RECT 102.000 235.000 102.800 235.800 ;
        RECT 106.200 235.200 106.800 235.800 ;
        RECT 105.400 234.600 109.000 235.200 ;
        RECT 111.600 235.000 112.400 235.800 ;
        RECT 105.400 234.400 106.200 234.600 ;
        RECT 108.200 234.400 109.000 234.600 ;
        RECT 101.200 233.200 102.600 234.000 ;
        RECT 102.000 232.200 102.600 233.200 ;
        RECT 104.200 233.000 106.400 233.600 ;
        RECT 104.200 232.800 105.000 233.000 ;
        RECT 102.000 231.600 104.400 232.200 ;
        RECT 97.200 230.600 101.400 231.200 ;
        RECT 95.600 226.800 96.400 228.400 ;
        RECT 97.200 227.200 98.000 230.600 ;
        RECT 100.600 230.400 101.400 230.600 ;
        RECT 99.000 229.800 99.800 230.000 ;
        RECT 99.000 229.200 102.800 229.800 ;
        RECT 102.000 229.000 102.800 229.200 ;
        RECT 103.800 228.400 104.400 231.600 ;
        RECT 105.800 231.800 106.400 233.000 ;
        RECT 107.000 233.000 107.800 233.200 ;
        RECT 111.600 233.000 112.400 233.200 ;
        RECT 107.000 232.400 112.400 233.000 ;
        RECT 105.800 231.400 110.600 231.800 ;
        RECT 114.800 231.400 115.600 239.800 ;
        RECT 105.800 231.200 115.600 231.400 ;
        RECT 109.800 231.000 115.600 231.200 ;
        RECT 110.000 230.800 115.600 231.000 ;
        RECT 116.400 231.200 117.200 239.800 ;
        RECT 120.600 235.800 121.800 239.800 ;
        RECT 125.200 235.800 126.000 239.800 ;
        RECT 129.600 236.400 130.400 239.800 ;
        RECT 129.600 235.800 131.600 236.400 ;
        RECT 121.200 235.000 122.000 235.800 ;
        RECT 125.400 235.200 126.000 235.800 ;
        RECT 124.600 234.600 128.200 235.200 ;
        RECT 130.800 235.000 131.600 235.800 ;
        RECT 124.600 234.400 125.400 234.600 ;
        RECT 127.400 234.400 128.200 234.600 ;
        RECT 120.400 233.200 121.800 234.000 ;
        RECT 121.200 232.200 121.800 233.200 ;
        RECT 123.400 233.000 125.600 233.600 ;
        RECT 123.400 232.800 124.200 233.000 ;
        RECT 121.200 231.600 123.600 232.200 ;
        RECT 116.400 230.600 120.600 231.200 ;
        RECT 108.400 230.200 109.200 230.400 ;
        RECT 108.400 229.600 113.400 230.200 ;
        RECT 110.000 229.400 110.800 229.600 ;
        RECT 112.600 229.400 113.400 229.600 ;
        RECT 111.000 228.400 111.800 228.600 ;
        RECT 103.800 227.800 114.800 228.400 ;
        RECT 104.200 227.600 105.000 227.800 ;
        RECT 106.800 227.600 107.600 227.800 ;
        RECT 85.600 222.200 87.200 225.800 ;
        RECT 90.800 222.200 91.600 226.200 ;
        RECT 93.000 225.600 94.800 226.200 ;
        RECT 97.200 226.600 101.000 227.200 ;
        RECT 93.000 224.400 93.800 225.600 ;
        RECT 92.400 223.600 93.800 224.400 ;
        RECT 93.000 222.200 93.800 223.600 ;
        RECT 97.200 222.200 98.000 226.600 ;
        RECT 100.200 226.400 101.000 226.600 ;
        RECT 110.000 225.600 110.600 227.800 ;
        RECT 113.200 227.600 114.800 227.800 ;
        RECT 116.400 227.200 117.200 230.600 ;
        RECT 119.800 230.400 120.600 230.600 ;
        RECT 118.200 229.800 119.000 230.000 ;
        RECT 118.200 229.200 122.000 229.800 ;
        RECT 121.200 229.000 122.000 229.200 ;
        RECT 123.000 228.400 123.600 231.600 ;
        RECT 125.000 231.800 125.600 233.000 ;
        RECT 126.200 233.000 127.000 233.200 ;
        RECT 130.800 233.000 131.600 233.200 ;
        RECT 126.200 232.400 131.600 233.000 ;
        RECT 125.000 231.400 129.800 231.800 ;
        RECT 134.000 231.400 134.800 239.800 ;
        RECT 140.400 232.400 141.200 239.800 ;
        RECT 141.800 232.400 142.600 232.600 ;
        RECT 140.400 231.800 142.600 232.400 ;
        RECT 144.800 232.400 146.400 239.800 ;
        RECT 148.400 232.400 149.200 232.600 ;
        RECT 150.000 232.400 150.800 239.800 ;
        RECT 154.200 232.400 155.000 239.800 ;
        RECT 155.600 233.600 156.400 234.400 ;
        RECT 155.800 232.400 156.400 233.600 ;
        RECT 160.600 232.400 161.400 239.800 ;
        RECT 162.000 233.600 162.800 234.400 ;
        RECT 162.200 232.400 162.800 233.600 ;
        RECT 144.800 231.800 146.800 232.400 ;
        RECT 148.400 231.800 150.800 232.400 ;
        RECT 125.000 231.200 134.800 231.400 ;
        RECT 129.000 231.000 134.800 231.200 ;
        RECT 129.200 230.800 134.800 231.000 ;
        RECT 142.000 231.200 142.600 231.800 ;
        RECT 142.000 230.600 145.400 231.200 ;
        RECT 144.600 230.400 145.400 230.600 ;
        RECT 146.200 230.400 146.800 231.800 ;
        RECT 153.200 231.600 155.200 232.400 ;
        RECT 155.800 231.800 157.200 232.400 ;
        RECT 160.600 231.800 161.600 232.400 ;
        RECT 162.200 231.800 163.600 232.400 ;
        RECT 156.400 231.600 157.200 231.800 ;
        RECT 127.600 230.200 128.400 230.400 ;
        RECT 127.600 229.600 132.600 230.200 ;
        RECT 129.200 229.400 130.000 229.600 ;
        RECT 131.800 229.400 132.600 229.600 ;
        RECT 142.400 229.800 143.200 230.000 ;
        RECT 146.200 229.800 147.600 230.400 ;
        RECT 142.400 229.200 145.000 229.800 ;
        RECT 144.400 228.600 145.000 229.200 ;
        RECT 145.800 229.600 147.600 229.800 ;
        RECT 145.800 229.200 146.800 229.600 ;
        RECT 130.200 228.400 131.000 228.600 ;
        RECT 123.000 227.800 134.000 228.400 ;
        RECT 123.400 227.600 124.200 227.800 ;
        RECT 108.200 225.400 109.000 225.600 ;
        RECT 102.000 224.200 102.800 225.000 ;
        RECT 106.200 224.800 109.000 225.400 ;
        RECT 110.000 224.800 110.800 225.600 ;
        RECT 106.200 224.200 106.800 224.800 ;
        RECT 111.600 224.200 112.400 225.000 ;
        RECT 101.400 223.600 102.800 224.200 ;
        RECT 101.400 222.200 102.600 223.600 ;
        RECT 106.000 222.200 106.800 224.200 ;
        RECT 110.400 223.600 112.400 224.200 ;
        RECT 110.400 222.200 111.200 223.600 ;
        RECT 114.800 222.200 115.600 227.000 ;
        RECT 116.400 226.600 120.200 227.200 ;
        RECT 116.400 222.200 117.200 226.600 ;
        RECT 119.400 226.400 120.200 226.600 ;
        RECT 129.200 225.600 129.800 227.800 ;
        RECT 132.400 227.600 134.000 227.800 ;
        RECT 140.400 228.200 142.000 228.400 ;
        RECT 140.400 227.600 143.800 228.200 ;
        RECT 144.400 227.800 145.200 228.600 ;
        RECT 143.200 227.200 143.800 227.600 ;
        RECT 127.400 225.400 128.200 225.600 ;
        RECT 121.200 224.200 122.000 225.000 ;
        RECT 125.400 224.800 128.200 225.400 ;
        RECT 129.200 224.800 130.000 225.600 ;
        RECT 125.400 224.200 126.000 224.800 ;
        RECT 130.800 224.200 131.600 225.000 ;
        RECT 120.600 223.600 122.000 224.200 ;
        RECT 120.600 222.200 121.800 223.600 ;
        RECT 125.200 222.200 126.000 224.200 ;
        RECT 129.600 223.600 131.600 224.200 ;
        RECT 129.600 222.200 130.400 223.600 ;
        RECT 134.000 222.200 134.800 227.000 ;
        RECT 141.800 226.800 142.600 227.000 ;
        RECT 140.400 226.200 142.600 226.800 ;
        RECT 143.200 226.600 145.200 227.200 ;
        RECT 143.600 226.400 145.200 226.600 ;
        RECT 140.400 222.200 141.200 226.200 ;
        RECT 145.800 225.800 146.400 229.200 ;
        RECT 153.200 228.800 154.000 230.400 ;
        RECT 154.600 228.400 155.200 231.600 ;
        RECT 156.500 230.300 157.100 231.600 ;
        RECT 159.600 230.300 160.400 230.400 ;
        RECT 156.500 229.700 160.400 230.300 ;
        RECT 159.600 228.800 160.400 229.700 ;
        RECT 161.000 228.400 161.600 231.800 ;
        RECT 162.800 231.600 163.600 231.800 ;
        RECT 164.400 231.200 165.200 239.800 ;
        RECT 168.600 235.800 169.800 239.800 ;
        RECT 173.200 235.800 174.000 239.800 ;
        RECT 177.600 236.400 178.400 239.800 ;
        RECT 177.600 235.800 179.600 236.400 ;
        RECT 169.200 235.000 170.000 235.800 ;
        RECT 173.400 235.200 174.000 235.800 ;
        RECT 172.600 234.600 176.200 235.200 ;
        RECT 178.800 235.000 179.600 235.800 ;
        RECT 172.600 234.400 173.400 234.600 ;
        RECT 175.400 234.400 176.200 234.600 ;
        RECT 168.400 233.200 169.800 234.000 ;
        RECT 169.200 232.200 169.800 233.200 ;
        RECT 171.400 233.000 173.600 233.600 ;
        RECT 171.400 232.800 172.200 233.000 ;
        RECT 169.200 231.600 171.600 232.200 ;
        RECT 164.400 230.600 168.600 231.200 ;
        RECT 147.200 227.600 148.000 228.400 ;
        RECT 149.200 227.600 150.800 228.400 ;
        RECT 151.600 228.200 152.400 228.400 ;
        RECT 151.600 227.600 153.200 228.200 ;
        RECT 154.600 227.600 157.200 228.400 ;
        RECT 158.000 228.200 158.800 228.400 ;
        RECT 158.000 227.600 159.600 228.200 ;
        RECT 161.000 227.600 163.600 228.400 ;
        RECT 147.200 227.200 147.800 227.600 ;
        RECT 152.400 227.200 153.200 227.600 ;
        RECT 147.000 226.400 147.800 227.200 ;
        RECT 148.400 226.800 149.200 227.000 ;
        RECT 148.400 226.200 150.800 226.800 ;
        RECT 151.800 226.200 155.400 226.600 ;
        RECT 156.400 226.200 157.000 227.600 ;
        RECT 158.800 227.200 159.600 227.600 ;
        RECT 158.200 226.200 161.800 226.600 ;
        RECT 162.800 226.200 163.400 227.600 ;
        RECT 164.400 227.200 165.200 230.600 ;
        RECT 167.800 230.400 168.600 230.600 ;
        RECT 166.200 229.800 167.000 230.000 ;
        RECT 166.200 229.200 170.000 229.800 ;
        RECT 169.200 229.000 170.000 229.200 ;
        RECT 171.000 228.400 171.600 231.600 ;
        RECT 173.000 231.800 173.600 233.000 ;
        RECT 174.200 233.000 175.000 233.200 ;
        RECT 178.800 233.000 179.600 233.200 ;
        RECT 174.200 232.400 179.600 233.000 ;
        RECT 173.000 231.400 177.800 231.800 ;
        RECT 182.000 231.400 182.800 239.800 ;
        RECT 173.000 231.200 182.800 231.400 ;
        RECT 177.000 231.000 182.800 231.200 ;
        RECT 177.200 230.800 182.800 231.000 ;
        RECT 185.200 231.200 186.000 239.800 ;
        RECT 188.400 231.200 189.200 239.800 ;
        RECT 191.600 231.200 192.400 239.800 ;
        RECT 194.800 231.200 195.600 239.800 ;
        RECT 198.000 231.200 198.800 239.800 ;
        RECT 202.200 235.800 203.400 239.800 ;
        RECT 206.800 235.800 207.600 239.800 ;
        RECT 211.200 236.400 212.000 239.800 ;
        RECT 211.200 235.800 213.200 236.400 ;
        RECT 202.800 235.000 203.600 235.800 ;
        RECT 207.000 235.200 207.600 235.800 ;
        RECT 206.200 234.600 209.800 235.200 ;
        RECT 212.400 235.000 213.200 235.800 ;
        RECT 206.200 234.400 207.000 234.600 ;
        RECT 209.000 234.400 209.800 234.600 ;
        RECT 202.000 233.200 203.400 234.000 ;
        RECT 202.800 232.200 203.400 233.200 ;
        RECT 205.000 233.000 207.200 233.600 ;
        RECT 205.000 232.800 205.800 233.000 ;
        RECT 202.800 231.600 205.200 232.200 ;
        RECT 185.200 230.400 187.000 231.200 ;
        RECT 188.400 230.400 190.600 231.200 ;
        RECT 191.600 230.400 193.800 231.200 ;
        RECT 194.800 230.400 197.200 231.200 ;
        RECT 175.600 230.200 176.400 230.400 ;
        RECT 175.600 229.600 180.600 230.200 ;
        RECT 177.200 229.400 178.000 229.600 ;
        RECT 179.800 229.400 180.600 229.600 ;
        RECT 186.200 229.000 187.000 230.400 ;
        RECT 189.800 229.000 190.600 230.400 ;
        RECT 193.000 229.000 193.800 230.400 ;
        RECT 178.200 228.400 179.000 228.600 ;
        RECT 170.800 227.800 182.000 228.400 ;
        RECT 170.800 227.600 172.200 227.800 ;
        RECT 164.400 226.600 168.200 227.200 ;
        RECT 144.800 224.400 146.400 225.800 ;
        RECT 143.600 223.600 146.400 224.400 ;
        RECT 144.800 222.200 146.400 223.600 ;
        RECT 150.000 222.200 150.800 226.200 ;
        RECT 151.600 226.000 155.600 226.200 ;
        RECT 151.600 222.200 152.400 226.000 ;
        RECT 154.800 222.200 155.600 226.000 ;
        RECT 156.400 222.200 157.200 226.200 ;
        RECT 158.000 226.000 162.000 226.200 ;
        RECT 158.000 222.200 158.800 226.000 ;
        RECT 161.200 222.200 162.000 226.000 ;
        RECT 162.800 222.200 163.600 226.200 ;
        RECT 164.400 222.200 165.200 226.600 ;
        RECT 167.400 226.400 168.200 226.600 ;
        RECT 177.200 225.600 177.800 227.800 ;
        RECT 180.400 227.600 182.000 227.800 ;
        RECT 186.200 228.200 188.800 229.000 ;
        RECT 189.800 228.200 192.200 229.000 ;
        RECT 193.000 228.200 195.600 229.000 ;
        RECT 186.200 227.600 187.000 228.200 ;
        RECT 189.800 227.600 190.600 228.200 ;
        RECT 193.000 227.600 193.800 228.200 ;
        RECT 196.400 227.600 197.200 230.400 ;
        RECT 175.400 225.400 176.200 225.600 ;
        RECT 169.200 224.200 170.000 225.000 ;
        RECT 173.400 224.800 176.200 225.400 ;
        RECT 177.200 224.800 178.000 225.600 ;
        RECT 173.400 224.200 174.000 224.800 ;
        RECT 178.800 224.200 179.600 225.000 ;
        RECT 168.600 223.600 170.000 224.200 ;
        RECT 168.600 222.200 169.800 223.600 ;
        RECT 173.200 222.200 174.000 224.200 ;
        RECT 177.600 223.600 179.600 224.200 ;
        RECT 177.600 222.200 178.400 223.600 ;
        RECT 182.000 222.200 182.800 227.000 ;
        RECT 185.200 226.800 187.000 227.600 ;
        RECT 188.400 226.800 190.600 227.600 ;
        RECT 191.600 226.800 193.800 227.600 ;
        RECT 194.800 226.800 197.200 227.600 ;
        RECT 198.000 230.600 202.200 231.200 ;
        RECT 198.000 227.200 198.800 230.600 ;
        RECT 201.400 230.400 202.200 230.600 ;
        RECT 204.600 230.400 205.200 231.600 ;
        RECT 206.600 231.800 207.200 233.000 ;
        RECT 207.800 233.000 208.600 233.200 ;
        RECT 212.400 233.000 213.200 233.200 ;
        RECT 207.800 232.400 213.200 233.000 ;
        RECT 206.600 231.400 211.400 231.800 ;
        RECT 215.600 231.400 216.400 239.800 ;
        RECT 206.600 231.200 216.400 231.400 ;
        RECT 210.600 231.000 216.400 231.200 ;
        RECT 210.800 230.800 216.400 231.000 ;
        RECT 217.200 231.200 218.000 239.800 ;
        RECT 221.400 235.800 222.600 239.800 ;
        RECT 226.000 235.800 226.800 239.800 ;
        RECT 230.400 236.400 231.200 239.800 ;
        RECT 230.400 235.800 232.400 236.400 ;
        RECT 222.000 235.000 222.800 235.800 ;
        RECT 226.200 235.200 226.800 235.800 ;
        RECT 225.400 234.600 229.000 235.200 ;
        RECT 231.600 235.000 232.400 235.800 ;
        RECT 225.400 234.400 226.200 234.600 ;
        RECT 228.200 234.400 229.000 234.600 ;
        RECT 221.200 233.200 222.600 234.000 ;
        RECT 222.000 232.200 222.600 233.200 ;
        RECT 224.200 233.000 226.400 233.600 ;
        RECT 224.200 232.800 225.000 233.000 ;
        RECT 222.000 231.600 224.400 232.200 ;
        RECT 217.200 230.600 221.400 231.200 ;
        RECT 199.800 229.800 200.600 230.000 ;
        RECT 199.800 229.200 203.600 229.800 ;
        RECT 204.400 229.600 205.200 230.400 ;
        RECT 209.200 230.200 210.000 230.400 ;
        RECT 209.200 229.600 214.200 230.200 ;
        RECT 202.800 229.000 203.600 229.200 ;
        RECT 204.600 228.400 205.200 229.600 ;
        RECT 210.800 229.400 211.600 229.600 ;
        RECT 213.400 229.400 214.200 229.600 ;
        RECT 211.800 228.400 212.600 228.600 ;
        RECT 204.600 227.800 215.600 228.400 ;
        RECT 205.000 227.600 205.800 227.800 ;
        RECT 185.200 222.200 186.000 226.800 ;
        RECT 188.400 222.200 189.200 226.800 ;
        RECT 191.600 222.200 192.400 226.800 ;
        RECT 194.800 222.200 195.600 226.800 ;
        RECT 198.000 226.600 201.800 227.200 ;
        RECT 198.000 222.200 198.800 226.600 ;
        RECT 201.000 226.400 201.800 226.600 ;
        RECT 210.800 225.600 211.400 227.800 ;
        RECT 214.000 227.600 215.600 227.800 ;
        RECT 217.200 227.200 218.000 230.600 ;
        RECT 220.600 230.400 221.400 230.600 ;
        RECT 223.800 230.400 224.400 231.600 ;
        RECT 225.800 231.800 226.400 233.000 ;
        RECT 227.000 233.000 227.800 233.200 ;
        RECT 231.600 233.000 232.400 233.200 ;
        RECT 227.000 232.400 232.400 233.000 ;
        RECT 225.800 231.400 230.600 231.800 ;
        RECT 234.800 231.400 235.600 239.800 ;
        RECT 225.800 231.200 235.600 231.400 ;
        RECT 229.800 231.000 235.600 231.200 ;
        RECT 230.000 230.800 235.600 231.000 ;
        RECT 219.000 229.800 219.800 230.000 ;
        RECT 219.000 229.200 222.800 229.800 ;
        RECT 223.600 229.600 224.400 230.400 ;
        RECT 228.400 230.200 229.200 230.400 ;
        RECT 228.400 229.600 233.400 230.200 ;
        RECT 222.000 229.000 222.800 229.200 ;
        RECT 223.800 228.400 224.400 229.600 ;
        RECT 230.000 229.400 230.800 229.600 ;
        RECT 232.600 229.400 233.400 229.600 ;
        RECT 231.000 228.400 231.800 228.600 ;
        RECT 223.800 227.800 234.800 228.400 ;
        RECT 224.200 227.600 225.000 227.800 ;
        RECT 209.000 225.400 209.800 225.600 ;
        RECT 202.800 224.200 203.600 225.000 ;
        RECT 207.000 224.800 209.800 225.400 ;
        RECT 210.800 224.800 211.600 225.600 ;
        RECT 207.000 224.200 207.600 224.800 ;
        RECT 212.400 224.200 213.200 225.000 ;
        RECT 202.200 223.600 203.600 224.200 ;
        RECT 202.200 222.200 203.400 223.600 ;
        RECT 206.800 222.200 207.600 224.200 ;
        RECT 211.200 223.600 213.200 224.200 ;
        RECT 211.200 222.200 212.000 223.600 ;
        RECT 215.600 222.200 216.400 227.000 ;
        RECT 217.200 226.600 221.000 227.200 ;
        RECT 217.200 222.200 218.000 226.600 ;
        RECT 220.200 226.400 221.000 226.600 ;
        RECT 230.000 225.600 230.600 227.800 ;
        RECT 233.200 227.600 234.800 227.800 ;
        RECT 228.200 225.400 229.000 225.600 ;
        RECT 222.000 224.200 222.800 225.000 ;
        RECT 226.200 224.800 229.000 225.400 ;
        RECT 230.000 224.800 230.800 225.600 ;
        RECT 226.200 224.200 226.800 224.800 ;
        RECT 231.600 224.200 232.400 225.000 ;
        RECT 221.400 223.600 222.800 224.200 ;
        RECT 221.400 222.200 222.600 223.600 ;
        RECT 226.000 222.200 226.800 224.200 ;
        RECT 230.400 223.600 232.400 224.200 ;
        RECT 230.400 222.200 231.200 223.600 ;
        RECT 234.800 222.200 235.600 227.000 ;
        RECT 236.400 224.800 237.200 226.400 ;
        RECT 238.000 222.200 238.800 239.800 ;
        RECT 239.600 231.800 240.400 239.800 ;
        RECT 242.800 232.400 243.600 239.800 ;
        RECT 241.400 231.800 243.600 232.400 ;
        RECT 239.600 229.600 240.200 231.800 ;
        RECT 241.400 231.200 242.000 231.800 ;
        RECT 240.800 230.400 242.000 231.200 ;
        RECT 244.400 231.400 245.200 239.800 ;
        RECT 248.800 236.400 249.600 239.800 ;
        RECT 247.600 235.800 249.600 236.400 ;
        RECT 253.200 235.800 254.000 239.800 ;
        RECT 257.400 235.800 258.600 239.800 ;
        RECT 247.600 235.000 248.400 235.800 ;
        RECT 253.200 235.200 253.800 235.800 ;
        RECT 251.000 234.600 254.600 235.200 ;
        RECT 257.200 235.000 258.000 235.800 ;
        RECT 251.000 234.400 251.800 234.600 ;
        RECT 253.800 234.400 254.600 234.600 ;
        RECT 258.200 234.000 259.600 234.400 ;
        RECT 257.400 233.600 259.600 234.000 ;
        RECT 247.600 233.000 248.400 233.200 ;
        RECT 252.200 233.000 253.000 233.200 ;
        RECT 247.600 232.400 253.000 233.000 ;
        RECT 253.600 233.000 255.800 233.600 ;
        RECT 253.600 231.800 254.200 233.000 ;
        RECT 255.000 232.800 255.800 233.000 ;
        RECT 257.400 233.200 258.800 233.600 ;
        RECT 257.400 232.200 258.000 233.200 ;
        RECT 249.400 231.400 254.200 231.800 ;
        RECT 244.400 231.200 254.200 231.400 ;
        RECT 255.600 231.600 258.000 232.200 ;
        RECT 244.400 231.000 250.200 231.200 ;
        RECT 244.400 230.800 250.000 231.000 ;
        RECT 239.600 222.200 240.400 229.600 ;
        RECT 241.400 227.400 242.000 230.400 ;
        RECT 242.800 228.800 243.600 230.400 ;
        RECT 250.800 230.200 251.600 230.400 ;
        RECT 246.600 229.600 251.600 230.200 ;
        RECT 246.600 229.400 247.400 229.600 ;
        RECT 249.200 229.400 250.000 229.600 ;
        RECT 248.200 228.400 249.000 228.600 ;
        RECT 255.600 228.400 256.200 231.600 ;
        RECT 262.000 231.200 262.800 239.800 ;
        RECT 258.600 230.600 262.800 231.200 ;
        RECT 263.600 231.400 264.400 239.800 ;
        RECT 268.000 236.400 268.800 239.800 ;
        RECT 266.800 235.800 268.800 236.400 ;
        RECT 272.400 235.800 273.200 239.800 ;
        RECT 276.600 235.800 277.800 239.800 ;
        RECT 266.800 235.000 267.600 235.800 ;
        RECT 272.400 235.200 273.000 235.800 ;
        RECT 270.200 234.600 273.800 235.200 ;
        RECT 276.400 235.000 277.200 235.800 ;
        RECT 270.200 234.400 271.000 234.600 ;
        RECT 273.000 234.400 273.800 234.600 ;
        RECT 266.800 233.000 267.600 233.200 ;
        RECT 271.400 233.000 272.200 233.200 ;
        RECT 266.800 232.400 272.200 233.000 ;
        RECT 272.800 233.000 275.000 233.600 ;
        RECT 272.800 231.800 273.400 233.000 ;
        RECT 274.200 232.800 275.000 233.000 ;
        RECT 276.600 233.200 278.000 234.000 ;
        RECT 276.600 232.200 277.200 233.200 ;
        RECT 268.600 231.400 273.400 231.800 ;
        RECT 263.600 231.200 273.400 231.400 ;
        RECT 274.800 231.600 277.200 232.200 ;
        RECT 263.600 231.000 269.400 231.200 ;
        RECT 263.600 230.800 269.200 231.000 ;
        RECT 258.600 230.400 259.400 230.600 ;
        RECT 260.200 229.800 261.000 230.000 ;
        RECT 257.200 229.200 261.000 229.800 ;
        RECT 257.200 229.000 258.000 229.200 ;
        RECT 245.200 227.800 256.200 228.400 ;
        RECT 245.200 227.600 246.800 227.800 ;
        RECT 241.400 226.800 243.600 227.400 ;
        RECT 242.800 222.200 243.600 226.800 ;
        RECT 244.400 222.200 245.200 227.000 ;
        RECT 249.400 225.600 250.000 227.800 ;
        RECT 255.000 227.600 255.800 227.800 ;
        RECT 262.000 227.200 262.800 230.600 ;
        RECT 270.000 230.200 270.800 230.400 ;
        RECT 265.800 229.600 270.800 230.200 ;
        RECT 265.800 229.400 266.600 229.600 ;
        RECT 267.400 228.400 268.200 228.600 ;
        RECT 274.800 228.400 275.400 231.600 ;
        RECT 281.200 231.200 282.000 239.800 ;
        RECT 277.800 230.600 282.000 231.200 ;
        RECT 277.800 230.400 278.600 230.600 ;
        RECT 279.400 229.800 280.200 230.000 ;
        RECT 276.400 229.200 280.200 229.800 ;
        RECT 276.400 229.000 277.200 229.200 ;
        RECT 264.400 227.800 275.400 228.400 ;
        RECT 264.400 227.600 266.000 227.800 ;
        RECT 259.000 226.600 262.800 227.200 ;
        RECT 259.000 226.400 259.800 226.600 ;
        RECT 247.600 224.200 248.400 225.000 ;
        RECT 249.200 224.800 250.000 225.600 ;
        RECT 251.000 225.400 251.800 225.600 ;
        RECT 251.000 224.800 253.800 225.400 ;
        RECT 253.200 224.200 253.800 224.800 ;
        RECT 257.200 224.200 258.000 225.000 ;
        RECT 247.600 223.600 249.600 224.200 ;
        RECT 248.800 222.200 249.600 223.600 ;
        RECT 253.200 222.200 254.000 224.200 ;
        RECT 257.200 223.600 258.600 224.200 ;
        RECT 257.400 222.200 258.600 223.600 ;
        RECT 262.000 222.200 262.800 226.600 ;
        RECT 263.600 222.200 264.400 227.000 ;
        RECT 268.600 225.600 269.200 227.800 ;
        RECT 274.200 227.600 275.000 227.800 ;
        RECT 281.200 227.200 282.000 230.600 ;
        RECT 278.200 226.600 282.000 227.200 ;
        RECT 278.200 226.400 279.000 226.600 ;
        RECT 266.800 224.200 267.600 225.000 ;
        RECT 268.400 224.800 269.200 225.600 ;
        RECT 270.200 225.400 271.000 225.600 ;
        RECT 270.200 224.800 273.000 225.400 ;
        RECT 272.400 224.200 273.000 224.800 ;
        RECT 276.400 224.200 277.200 225.000 ;
        RECT 266.800 223.600 268.800 224.200 ;
        RECT 268.000 222.200 268.800 223.600 ;
        RECT 272.400 222.200 273.200 224.200 ;
        RECT 276.400 223.600 277.800 224.200 ;
        RECT 276.600 222.200 277.800 223.600 ;
        RECT 281.200 222.200 282.000 226.600 ;
        RECT 284.400 228.300 285.200 239.800 ;
        RECT 286.000 228.300 286.800 228.400 ;
        RECT 284.400 227.700 286.800 228.300 ;
        RECT 282.800 224.800 283.600 226.400 ;
        RECT 284.400 222.200 285.200 227.700 ;
        RECT 286.000 226.800 286.800 227.700 ;
        RECT 287.600 228.300 288.400 239.800 ;
        RECT 296.200 234.400 297.000 239.800 ;
        RECT 296.200 233.600 298.000 234.400 ;
        RECT 289.200 231.600 290.000 233.200 ;
        RECT 296.200 232.600 297.000 233.600 ;
        RECT 296.200 231.800 298.000 232.600 ;
        RECT 294.000 230.300 294.800 230.400 ;
        RECT 295.600 230.300 296.400 231.200 ;
        RECT 294.000 229.700 296.400 230.300 ;
        RECT 294.000 229.600 294.800 229.700 ;
        RECT 295.600 229.600 296.400 229.700 ;
        RECT 297.200 228.400 297.800 231.800 ;
        RECT 295.600 228.300 296.400 228.400 ;
        RECT 287.600 227.700 296.400 228.300 ;
        RECT 287.600 226.200 288.400 227.700 ;
        RECT 295.600 227.600 296.400 227.700 ;
        RECT 297.200 227.600 298.000 228.400 ;
        RECT 287.600 225.600 289.400 226.200 ;
        RECT 288.600 222.200 289.400 225.600 ;
        RECT 297.200 224.200 297.800 227.600 ;
        RECT 298.800 226.300 299.600 226.400 ;
        RECT 300.400 226.300 301.200 239.800 ;
        RECT 306.200 232.600 307.000 239.800 ;
        RECT 305.200 231.800 307.000 232.600 ;
        RECT 305.200 231.600 306.000 231.800 ;
        RECT 305.400 228.400 306.000 231.600 ;
        RECT 308.400 231.400 309.200 239.800 ;
        RECT 312.800 236.400 313.600 239.800 ;
        RECT 311.600 235.800 313.600 236.400 ;
        RECT 317.200 235.800 318.000 239.800 ;
        RECT 321.400 235.800 322.600 239.800 ;
        RECT 311.600 235.000 312.400 235.800 ;
        RECT 317.200 235.200 317.800 235.800 ;
        RECT 315.000 234.600 318.600 235.200 ;
        RECT 321.200 235.000 322.000 235.800 ;
        RECT 315.000 234.400 315.800 234.600 ;
        RECT 317.800 234.400 318.600 234.600 ;
        RECT 311.600 233.000 312.400 233.200 ;
        RECT 316.200 233.000 317.000 233.200 ;
        RECT 311.600 232.400 317.000 233.000 ;
        RECT 317.600 233.000 319.800 233.600 ;
        RECT 317.600 231.800 318.200 233.000 ;
        RECT 319.000 232.800 319.800 233.000 ;
        RECT 321.400 233.200 322.800 234.000 ;
        RECT 321.400 232.200 322.000 233.200 ;
        RECT 313.400 231.400 318.200 231.800 ;
        RECT 308.400 231.200 318.200 231.400 ;
        RECT 319.600 231.600 322.000 232.200 ;
        RECT 306.800 229.600 307.600 231.200 ;
        RECT 308.400 231.000 314.200 231.200 ;
        RECT 308.400 230.800 314.000 231.000 ;
        RECT 314.800 230.200 315.600 230.400 ;
        RECT 310.600 229.600 315.600 230.200 ;
        RECT 310.600 229.400 311.400 229.600 ;
        RECT 312.200 228.400 313.000 228.600 ;
        RECT 319.600 228.400 320.200 231.600 ;
        RECT 326.000 231.200 326.800 239.800 ;
        RECT 327.600 231.600 328.400 233.200 ;
        RECT 322.600 230.600 326.800 231.200 ;
        RECT 322.600 230.400 323.400 230.600 ;
        RECT 324.200 229.800 325.000 230.000 ;
        RECT 321.200 229.200 325.000 229.800 ;
        RECT 321.200 229.000 322.000 229.200 ;
        RECT 305.200 227.600 306.000 228.400 ;
        RECT 309.200 227.800 320.200 228.400 ;
        RECT 309.200 227.600 310.800 227.800 ;
        RECT 298.800 225.700 301.200 226.300 ;
        RECT 298.800 224.800 299.600 225.700 ;
        RECT 297.200 222.200 298.000 224.200 ;
        RECT 300.400 222.200 301.200 225.700 ;
        RECT 302.000 226.300 302.800 226.400 ;
        RECT 303.600 226.300 304.400 226.400 ;
        RECT 302.000 225.700 304.400 226.300 ;
        RECT 302.000 224.800 302.800 225.700 ;
        RECT 303.600 224.800 304.400 225.700 ;
        RECT 305.400 224.200 306.000 227.600 ;
        RECT 305.200 222.200 306.000 224.200 ;
        RECT 308.400 222.200 309.200 227.000 ;
        RECT 313.400 225.600 314.000 227.800 ;
        RECT 319.000 227.600 319.800 227.800 ;
        RECT 326.000 227.200 326.800 230.600 ;
        RECT 323.000 226.600 326.800 227.200 ;
        RECT 323.000 226.400 323.800 226.600 ;
        RECT 311.600 224.200 312.400 225.000 ;
        RECT 313.200 224.800 314.000 225.600 ;
        RECT 315.000 225.400 315.800 225.600 ;
        RECT 315.000 224.800 317.800 225.400 ;
        RECT 317.200 224.200 317.800 224.800 ;
        RECT 321.200 224.200 322.000 225.000 ;
        RECT 311.600 223.600 313.600 224.200 ;
        RECT 312.800 222.200 313.600 223.600 ;
        RECT 317.200 222.200 318.000 224.200 ;
        RECT 321.200 223.600 322.600 224.200 ;
        RECT 321.400 222.200 322.600 223.600 ;
        RECT 326.000 222.200 326.800 226.600 ;
        RECT 329.200 226.200 330.000 239.800 ;
        RECT 330.800 228.300 331.600 228.400 ;
        RECT 334.000 228.300 334.800 239.800 ;
        RECT 335.600 228.300 336.400 228.400 ;
        RECT 330.800 227.700 333.100 228.300 ;
        RECT 330.800 226.800 331.600 227.700 ;
        RECT 332.500 226.400 333.100 227.700 ;
        RECT 334.000 227.700 336.400 228.300 ;
        RECT 328.200 225.600 330.000 226.200 ;
        RECT 328.200 224.400 329.000 225.600 ;
        RECT 332.400 224.800 333.200 226.400 ;
        RECT 328.200 223.600 330.000 224.400 ;
        RECT 328.200 222.200 329.000 223.600 ;
        RECT 334.000 222.200 334.800 227.700 ;
        RECT 335.600 226.800 336.400 227.700 ;
        RECT 337.200 226.200 338.000 239.800 ;
        RECT 338.800 231.600 339.600 233.200 ;
        RECT 340.400 231.400 341.200 239.800 ;
        RECT 344.800 236.400 345.600 239.800 ;
        RECT 343.600 235.800 345.600 236.400 ;
        RECT 349.200 235.800 350.000 239.800 ;
        RECT 353.400 235.800 354.600 239.800 ;
        RECT 343.600 235.000 344.400 235.800 ;
        RECT 349.200 235.200 349.800 235.800 ;
        RECT 347.000 234.600 350.600 235.200 ;
        RECT 353.200 235.000 354.000 235.800 ;
        RECT 347.000 234.400 347.800 234.600 ;
        RECT 349.800 234.400 350.600 234.600 ;
        RECT 343.600 233.000 344.400 233.200 ;
        RECT 348.200 233.000 349.000 233.200 ;
        RECT 343.600 232.400 349.000 233.000 ;
        RECT 349.600 233.000 351.800 233.600 ;
        RECT 349.600 231.800 350.200 233.000 ;
        RECT 351.000 232.800 351.800 233.000 ;
        RECT 353.400 233.200 354.800 234.000 ;
        RECT 353.400 232.200 354.000 233.200 ;
        RECT 345.400 231.400 350.200 231.800 ;
        RECT 340.400 231.200 350.200 231.400 ;
        RECT 351.600 231.600 354.000 232.200 ;
        RECT 340.400 231.000 346.200 231.200 ;
        RECT 340.400 230.800 346.000 231.000 ;
        RECT 351.600 230.400 352.200 231.600 ;
        RECT 358.000 231.200 358.800 239.800 ;
        RECT 359.600 232.400 360.400 239.800 ;
        RECT 359.600 231.800 361.800 232.400 ;
        RECT 362.800 231.800 363.600 239.800 ;
        RECT 354.600 230.600 358.800 231.200 ;
        RECT 354.600 230.400 355.400 230.600 ;
        RECT 346.800 230.200 347.600 230.400 ;
        RECT 342.600 229.600 347.600 230.200 ;
        RECT 351.600 229.600 352.400 230.400 ;
        RECT 356.200 229.800 357.000 230.000 ;
        RECT 342.600 229.400 343.400 229.600 ;
        RECT 345.200 229.400 346.000 229.600 ;
        RECT 344.200 228.400 345.000 228.600 ;
        RECT 351.600 228.400 352.200 229.600 ;
        RECT 353.200 229.200 357.000 229.800 ;
        RECT 353.200 229.000 354.000 229.200 ;
        RECT 341.200 227.800 352.200 228.400 ;
        RECT 341.200 227.600 342.800 227.800 ;
        RECT 337.200 225.600 339.000 226.200 ;
        RECT 338.200 224.400 339.000 225.600 ;
        RECT 338.200 223.600 339.600 224.400 ;
        RECT 338.200 222.200 339.000 223.600 ;
        RECT 340.400 222.200 341.200 227.000 ;
        RECT 345.400 225.600 346.000 227.800 ;
        RECT 351.000 227.600 351.800 227.800 ;
        RECT 358.000 227.200 358.800 230.600 ;
        RECT 361.200 231.200 361.800 231.800 ;
        RECT 361.200 230.400 362.400 231.200 ;
        RECT 359.600 228.800 360.400 230.400 ;
        RECT 361.200 227.400 361.800 230.400 ;
        RECT 363.000 229.600 363.600 231.800 ;
        RECT 355.000 226.600 358.800 227.200 ;
        RECT 355.000 226.400 355.800 226.600 ;
        RECT 343.600 224.200 344.400 225.000 ;
        RECT 345.200 224.800 346.000 225.600 ;
        RECT 347.000 225.400 347.800 225.600 ;
        RECT 347.000 224.800 349.800 225.400 ;
        RECT 349.200 224.200 349.800 224.800 ;
        RECT 353.200 224.200 354.000 225.000 ;
        RECT 343.600 223.600 345.600 224.200 ;
        RECT 344.800 222.200 345.600 223.600 ;
        RECT 349.200 222.200 350.000 224.200 ;
        RECT 353.200 223.600 354.600 224.200 ;
        RECT 353.400 222.200 354.600 223.600 ;
        RECT 358.000 222.200 358.800 226.600 ;
        RECT 359.600 226.800 361.800 227.400 ;
        RECT 359.600 222.200 360.400 226.800 ;
        RECT 362.800 222.200 363.600 229.600 ;
        RECT 364.400 231.200 365.200 239.800 ;
        RECT 368.600 235.800 369.800 239.800 ;
        RECT 373.200 235.800 374.000 239.800 ;
        RECT 377.600 236.400 378.400 239.800 ;
        RECT 377.600 235.800 379.600 236.400 ;
        RECT 369.200 235.000 370.000 235.800 ;
        RECT 373.400 235.200 374.000 235.800 ;
        RECT 372.600 234.600 376.200 235.200 ;
        RECT 378.800 235.000 379.600 235.800 ;
        RECT 372.600 234.400 373.400 234.600 ;
        RECT 375.400 234.400 376.200 234.600 ;
        RECT 368.400 233.200 369.800 234.000 ;
        RECT 369.200 232.200 369.800 233.200 ;
        RECT 371.400 233.000 373.600 233.600 ;
        RECT 371.400 232.800 372.200 233.000 ;
        RECT 369.200 231.600 371.600 232.200 ;
        RECT 364.400 230.600 368.600 231.200 ;
        RECT 364.400 227.200 365.200 230.600 ;
        RECT 367.800 230.400 368.600 230.600 ;
        RECT 366.200 229.800 367.000 230.000 ;
        RECT 366.200 229.200 370.000 229.800 ;
        RECT 369.200 229.000 370.000 229.200 ;
        RECT 371.000 228.400 371.600 231.600 ;
        RECT 373.000 231.800 373.600 233.000 ;
        RECT 374.200 233.000 375.000 233.200 ;
        RECT 378.800 233.000 379.600 233.200 ;
        RECT 374.200 232.400 379.600 233.000 ;
        RECT 373.000 231.400 377.800 231.800 ;
        RECT 382.000 231.400 382.800 239.800 ;
        RECT 373.000 231.200 382.800 231.400 ;
        RECT 377.000 231.000 382.800 231.200 ;
        RECT 377.200 230.800 382.800 231.000 ;
        RECT 383.600 231.400 384.400 239.800 ;
        RECT 388.000 236.400 388.800 239.800 ;
        RECT 386.800 235.800 388.800 236.400 ;
        RECT 392.400 235.800 393.200 239.800 ;
        RECT 396.600 235.800 397.800 239.800 ;
        RECT 386.800 235.000 387.600 235.800 ;
        RECT 392.400 235.200 393.000 235.800 ;
        RECT 390.200 234.600 393.800 235.200 ;
        RECT 396.400 235.000 397.200 235.800 ;
        RECT 390.200 234.400 391.000 234.600 ;
        RECT 393.000 234.400 393.800 234.600 ;
        RECT 386.800 233.000 387.600 233.200 ;
        RECT 391.400 233.000 392.200 233.200 ;
        RECT 386.800 232.400 392.200 233.000 ;
        RECT 392.800 233.000 395.000 233.600 ;
        RECT 392.800 231.800 393.400 233.000 ;
        RECT 394.200 232.800 395.000 233.000 ;
        RECT 396.600 233.200 398.000 234.000 ;
        RECT 396.600 232.200 397.200 233.200 ;
        RECT 388.600 231.400 393.400 231.800 ;
        RECT 383.600 231.200 393.400 231.400 ;
        RECT 394.800 231.600 397.200 232.200 ;
        RECT 383.600 231.000 389.400 231.200 ;
        RECT 383.600 230.800 389.200 231.000 ;
        RECT 394.800 230.400 395.400 231.600 ;
        RECT 401.200 231.200 402.000 239.800 ;
        RECT 397.800 230.600 402.000 231.200 ;
        RECT 402.800 231.400 403.600 239.800 ;
        RECT 407.200 236.400 408.000 239.800 ;
        RECT 406.000 235.800 408.000 236.400 ;
        RECT 411.600 235.800 412.400 239.800 ;
        RECT 415.800 235.800 417.000 239.800 ;
        RECT 406.000 235.000 406.800 235.800 ;
        RECT 411.600 235.200 412.200 235.800 ;
        RECT 409.400 234.600 413.000 235.200 ;
        RECT 415.600 235.000 416.400 235.800 ;
        RECT 409.400 234.400 410.200 234.600 ;
        RECT 412.200 234.400 413.000 234.600 ;
        RECT 420.400 234.300 421.200 239.800 ;
        RECT 422.000 234.300 422.800 234.400 ;
        RECT 406.000 233.000 406.800 233.200 ;
        RECT 410.600 233.000 411.400 233.200 ;
        RECT 406.000 232.400 411.400 233.000 ;
        RECT 412.000 233.000 414.200 233.600 ;
        RECT 412.000 231.800 412.600 233.000 ;
        RECT 413.400 232.800 414.200 233.000 ;
        RECT 415.800 233.200 417.200 234.000 ;
        RECT 420.400 233.700 422.800 234.300 ;
        RECT 415.800 232.200 416.400 233.200 ;
        RECT 407.800 231.400 412.600 231.800 ;
        RECT 402.800 231.200 412.600 231.400 ;
        RECT 414.000 231.600 416.400 232.200 ;
        RECT 402.800 231.000 408.600 231.200 ;
        RECT 402.800 230.800 408.400 231.000 ;
        RECT 397.800 230.400 398.600 230.600 ;
        RECT 375.600 230.200 376.400 230.400 ;
        RECT 390.000 230.200 390.800 230.400 ;
        RECT 375.600 229.600 380.600 230.200 ;
        RECT 379.800 229.400 380.600 229.600 ;
        RECT 385.800 229.600 390.800 230.200 ;
        RECT 394.800 229.600 395.600 230.400 ;
        RECT 399.400 229.800 400.200 230.000 ;
        RECT 385.800 229.400 386.600 229.600 ;
        RECT 388.400 229.400 389.200 229.600 ;
        RECT 378.200 228.400 379.000 228.600 ;
        RECT 387.400 228.400 388.200 228.600 ;
        RECT 394.800 228.400 395.400 229.600 ;
        RECT 396.400 229.200 400.200 229.800 ;
        RECT 396.400 229.000 397.200 229.200 ;
        RECT 371.000 228.300 382.000 228.400 ;
        RECT 384.400 228.300 395.400 228.400 ;
        RECT 371.000 227.800 395.400 228.300 ;
        RECT 371.400 227.600 372.200 227.800 ;
        RECT 364.400 226.600 368.200 227.200 ;
        RECT 364.400 222.200 365.200 226.600 ;
        RECT 367.400 226.400 368.200 226.600 ;
        RECT 377.200 225.600 377.800 227.800 ;
        RECT 380.400 227.700 386.000 227.800 ;
        RECT 380.400 227.600 382.000 227.700 ;
        RECT 384.400 227.600 386.000 227.700 ;
        RECT 375.400 225.400 376.200 225.600 ;
        RECT 369.200 224.200 370.000 225.000 ;
        RECT 373.400 224.800 376.200 225.400 ;
        RECT 377.200 224.800 378.000 225.600 ;
        RECT 373.400 224.200 374.000 224.800 ;
        RECT 378.800 224.200 379.600 225.000 ;
        RECT 368.600 223.600 370.000 224.200 ;
        RECT 368.600 222.200 369.800 223.600 ;
        RECT 373.200 222.200 374.000 224.200 ;
        RECT 377.600 223.600 379.600 224.200 ;
        RECT 377.600 222.200 378.400 223.600 ;
        RECT 382.000 222.200 382.800 227.000 ;
        RECT 383.600 222.200 384.400 227.000 ;
        RECT 388.600 225.600 389.200 227.800 ;
        RECT 394.200 227.600 395.000 227.800 ;
        RECT 401.200 227.200 402.000 230.600 ;
        RECT 414.000 230.400 414.600 231.600 ;
        RECT 420.400 231.200 421.200 233.700 ;
        RECT 422.000 233.600 422.800 233.700 ;
        RECT 417.000 230.600 421.200 231.200 ;
        RECT 417.000 230.400 417.800 230.600 ;
        RECT 409.200 230.200 410.000 230.400 ;
        RECT 405.000 229.600 410.000 230.200 ;
        RECT 414.000 229.600 414.800 230.400 ;
        RECT 418.600 229.800 419.400 230.000 ;
        RECT 405.000 229.400 405.800 229.600 ;
        RECT 407.600 229.400 408.400 229.600 ;
        RECT 406.600 228.400 407.400 228.600 ;
        RECT 414.000 228.400 414.600 229.600 ;
        RECT 415.600 229.200 419.400 229.800 ;
        RECT 415.600 229.000 416.400 229.200 ;
        RECT 403.600 227.800 414.600 228.400 ;
        RECT 420.400 228.300 421.200 230.600 ;
        RECT 422.000 228.300 422.800 228.400 ;
        RECT 403.600 227.600 405.200 227.800 ;
        RECT 398.200 226.600 402.000 227.200 ;
        RECT 398.200 226.400 399.000 226.600 ;
        RECT 386.800 224.200 387.600 225.000 ;
        RECT 388.400 224.800 389.200 225.600 ;
        RECT 390.200 225.400 391.000 225.600 ;
        RECT 390.200 224.800 393.000 225.400 ;
        RECT 392.400 224.200 393.000 224.800 ;
        RECT 396.400 224.200 397.200 225.000 ;
        RECT 386.800 223.600 388.800 224.200 ;
        RECT 388.000 222.200 388.800 223.600 ;
        RECT 392.400 222.200 393.200 224.200 ;
        RECT 396.400 223.600 397.800 224.200 ;
        RECT 396.600 222.200 397.800 223.600 ;
        RECT 401.200 222.200 402.000 226.600 ;
        RECT 402.800 222.200 403.600 227.000 ;
        RECT 407.800 225.600 408.400 227.800 ;
        RECT 413.400 227.600 414.200 227.800 ;
        RECT 420.400 227.700 422.800 228.300 ;
        RECT 420.400 227.200 421.200 227.700 ;
        RECT 417.400 226.600 421.200 227.200 ;
        RECT 422.000 226.800 422.800 227.700 ;
        RECT 417.400 226.400 418.200 226.600 ;
        RECT 406.000 224.200 406.800 225.000 ;
        RECT 407.600 224.800 408.400 225.600 ;
        RECT 409.400 225.400 410.200 225.600 ;
        RECT 409.400 224.800 412.200 225.400 ;
        RECT 411.600 224.200 412.200 224.800 ;
        RECT 415.600 224.200 416.400 225.000 ;
        RECT 406.000 223.600 408.000 224.200 ;
        RECT 407.200 222.200 408.000 223.600 ;
        RECT 411.600 222.200 412.400 224.200 ;
        RECT 415.600 223.600 417.000 224.200 ;
        RECT 415.800 222.200 417.000 223.600 ;
        RECT 420.400 222.200 421.200 226.600 ;
        RECT 423.600 226.300 424.400 239.800 ;
        RECT 425.200 231.600 426.000 233.200 ;
        RECT 429.400 232.600 430.200 239.800 ;
        RECT 428.400 231.800 430.200 232.600 ;
        RECT 432.200 238.400 433.000 239.800 ;
        RECT 432.200 237.600 434.000 238.400 ;
        RECT 432.200 232.600 433.000 237.600 ;
        RECT 432.200 231.800 434.000 232.600 ;
        RECT 428.600 228.400 429.200 231.800 ;
        RECT 430.000 229.600 430.800 231.200 ;
        RECT 431.600 229.600 432.400 231.200 ;
        RECT 428.400 228.300 429.200 228.400 ;
        RECT 431.700 228.300 432.300 229.600 ;
        RECT 428.400 227.700 432.300 228.300 ;
        RECT 433.200 228.400 433.800 231.800 ;
        RECT 428.400 227.600 429.200 227.700 ;
        RECT 426.800 226.300 427.600 226.400 ;
        RECT 423.600 225.700 427.600 226.300 ;
        RECT 423.600 225.600 425.400 225.700 ;
        RECT 424.600 222.200 425.400 225.600 ;
        RECT 426.800 224.800 427.600 225.700 ;
        RECT 428.600 224.400 429.200 227.600 ;
        RECT 428.400 222.200 429.200 224.400 ;
        RECT 433.200 227.600 434.000 228.400 ;
        RECT 433.200 224.200 433.800 227.600 ;
        RECT 434.800 224.800 435.600 226.400 ;
        RECT 436.400 224.800 437.200 226.400 ;
        RECT 433.200 222.200 434.000 224.200 ;
        RECT 438.000 222.200 438.800 239.800 ;
        RECT 439.600 235.800 440.400 239.800 ;
        RECT 439.800 235.600 440.400 235.800 ;
        RECT 442.800 235.800 443.600 239.800 ;
        RECT 442.800 235.600 443.400 235.800 ;
        RECT 439.800 235.000 443.400 235.600 ;
        RECT 439.800 232.400 440.400 235.000 ;
        RECT 441.200 232.800 442.000 234.400 ;
        RECT 442.800 234.300 443.600 234.400 ;
        RECT 450.800 234.300 451.600 239.800 ;
        RECT 442.800 233.700 451.600 234.300 ;
        RECT 442.800 233.600 443.600 233.700 ;
        RECT 439.600 231.600 440.400 232.400 ;
        RECT 439.800 228.400 440.400 231.600 ;
        RECT 444.400 230.800 445.200 232.400 ;
        RECT 442.000 229.600 443.600 230.400 ;
        RECT 439.800 228.200 441.400 228.400 ;
        RECT 439.800 227.800 441.600 228.200 ;
        RECT 440.800 222.200 441.600 227.800 ;
        RECT 450.800 222.200 451.600 233.700 ;
        RECT 454.600 234.400 455.400 239.800 ;
        RECT 454.600 233.600 456.400 234.400 ;
        RECT 454.600 232.600 455.400 233.600 ;
        RECT 454.600 231.800 456.400 232.600 ;
        RECT 452.400 230.300 453.200 230.400 ;
        RECT 454.000 230.300 454.800 231.200 ;
        RECT 452.400 229.700 454.800 230.300 ;
        RECT 452.400 229.600 453.200 229.700 ;
        RECT 454.000 229.600 454.800 229.700 ;
        RECT 455.600 228.400 456.200 231.800 ;
        RECT 458.800 231.600 459.600 233.200 ;
        RECT 455.600 227.600 456.400 228.400 ;
        RECT 452.400 226.300 453.200 226.400 ;
        RECT 454.000 226.300 454.800 226.400 ;
        RECT 452.400 225.700 454.800 226.300 ;
        RECT 452.400 224.800 453.200 225.700 ;
        RECT 454.000 225.600 454.800 225.700 ;
        RECT 455.600 224.200 456.200 227.600 ;
        RECT 457.200 224.800 458.000 226.400 ;
        RECT 460.400 226.200 461.200 239.800 ;
        RECT 462.000 228.300 462.800 228.400 ;
        RECT 463.600 228.300 464.400 228.400 ;
        RECT 462.000 227.700 464.400 228.300 ;
        RECT 462.000 226.800 462.800 227.700 ;
        RECT 463.600 226.800 464.400 227.700 ;
        RECT 459.400 225.600 461.200 226.200 ;
        RECT 465.200 226.200 466.000 239.800 ;
        RECT 466.800 231.600 467.600 233.200 ;
        RECT 471.000 231.800 473.000 239.800 ;
        RECT 466.800 228.300 467.600 228.400 ;
        RECT 468.400 228.300 469.200 229.200 ;
        RECT 470.000 228.800 470.800 230.400 ;
        RECT 471.800 228.400 472.400 231.800 ;
        RECT 473.200 228.800 474.000 230.400 ;
        RECT 466.800 227.700 469.200 228.300 ;
        RECT 471.600 228.200 472.400 228.400 ;
        RECT 474.800 228.200 475.600 228.400 ;
        RECT 466.800 227.600 467.600 227.700 ;
        RECT 468.400 227.600 469.200 227.700 ;
        RECT 470.000 227.600 472.400 228.200 ;
        RECT 474.000 227.600 475.600 228.200 ;
        RECT 470.000 226.200 470.600 227.600 ;
        RECT 474.000 227.200 474.800 227.600 ;
        RECT 471.800 226.200 475.400 226.600 ;
        RECT 465.200 225.600 467.000 226.200 ;
        RECT 459.400 224.400 460.200 225.600 ;
        RECT 455.600 222.200 456.400 224.200 ;
        RECT 459.400 223.600 461.200 224.400 ;
        RECT 459.400 222.200 460.200 223.600 ;
        RECT 466.200 222.200 467.000 225.600 ;
        RECT 468.400 222.800 469.200 226.200 ;
        RECT 470.000 223.400 470.800 226.200 ;
        RECT 471.600 226.000 475.600 226.200 ;
        RECT 471.600 222.800 472.400 226.000 ;
        RECT 468.400 222.200 472.400 222.800 ;
        RECT 474.800 222.200 475.600 226.000 ;
        RECT 476.400 224.800 477.200 226.400 ;
        RECT 478.000 222.200 478.800 239.800 ;
        RECT 479.600 232.400 480.400 239.800 ;
        RECT 484.000 234.400 485.600 239.800 ;
        RECT 484.000 233.600 486.800 234.400 ;
        RECT 481.200 232.400 482.000 232.600 ;
        RECT 484.000 232.400 485.600 233.600 ;
        RECT 479.600 231.800 482.000 232.400 ;
        RECT 483.600 231.800 485.600 232.400 ;
        RECT 487.800 232.400 488.600 232.600 ;
        RECT 489.200 232.400 490.000 239.800 ;
        RECT 487.800 231.800 490.000 232.400 ;
        RECT 483.600 230.400 484.200 231.800 ;
        RECT 487.800 231.200 488.400 231.800 ;
        RECT 485.000 230.600 488.400 231.200 ;
        RECT 490.800 231.400 491.600 239.800 ;
        RECT 495.200 236.400 496.000 239.800 ;
        RECT 494.000 235.800 496.000 236.400 ;
        RECT 499.600 235.800 500.400 239.800 ;
        RECT 503.800 235.800 505.000 239.800 ;
        RECT 494.000 235.000 494.800 235.800 ;
        RECT 499.600 235.200 500.200 235.800 ;
        RECT 497.400 234.600 501.000 235.200 ;
        RECT 503.600 235.000 504.400 235.800 ;
        RECT 497.400 234.400 498.200 234.600 ;
        RECT 500.200 234.400 501.000 234.600 ;
        RECT 494.000 233.000 494.800 233.200 ;
        RECT 498.600 233.000 499.400 233.200 ;
        RECT 494.000 232.400 499.400 233.000 ;
        RECT 500.000 233.000 502.200 233.600 ;
        RECT 500.000 231.800 500.600 233.000 ;
        RECT 501.400 232.800 502.200 233.000 ;
        RECT 503.800 233.200 505.200 234.000 ;
        RECT 503.800 232.200 504.400 233.200 ;
        RECT 495.800 231.400 500.600 231.800 ;
        RECT 490.800 231.200 500.600 231.400 ;
        RECT 502.000 231.600 504.400 232.200 ;
        RECT 490.800 231.000 496.600 231.200 ;
        RECT 490.800 230.800 496.400 231.000 ;
        RECT 485.000 230.400 485.800 230.600 ;
        RECT 482.800 229.800 484.200 230.400 ;
        RECT 497.200 230.200 498.000 230.400 ;
        RECT 487.200 229.800 488.000 230.000 ;
        RECT 482.800 229.600 484.600 229.800 ;
        RECT 483.600 229.200 484.600 229.600 ;
        RECT 479.600 227.600 481.200 228.400 ;
        RECT 482.400 227.600 483.200 228.400 ;
        RECT 482.600 227.200 483.200 227.600 ;
        RECT 481.200 226.800 482.000 227.000 ;
        RECT 479.600 226.200 482.000 226.800 ;
        RECT 482.600 226.400 483.400 227.200 ;
        RECT 479.600 222.200 480.400 226.200 ;
        RECT 484.000 225.800 484.600 229.200 ;
        RECT 485.400 229.200 488.000 229.800 ;
        RECT 493.000 229.600 498.000 230.200 ;
        RECT 493.000 229.400 493.800 229.600 ;
        RECT 495.600 229.400 496.400 229.600 ;
        RECT 485.400 228.600 486.000 229.200 ;
        RECT 485.200 227.800 486.000 228.600 ;
        RECT 494.600 228.400 495.400 228.600 ;
        RECT 502.000 228.400 502.600 231.600 ;
        RECT 508.400 231.200 509.200 239.800 ;
        RECT 505.000 230.600 509.200 231.200 ;
        RECT 510.000 231.400 510.800 239.800 ;
        RECT 514.400 236.400 515.200 239.800 ;
        RECT 513.200 235.800 515.200 236.400 ;
        RECT 518.800 235.800 519.600 239.800 ;
        RECT 523.000 235.800 524.200 239.800 ;
        RECT 513.200 235.000 514.000 235.800 ;
        RECT 518.800 235.200 519.400 235.800 ;
        RECT 516.600 234.600 520.200 235.200 ;
        RECT 522.800 235.000 523.600 235.800 ;
        RECT 516.600 234.400 517.400 234.600 ;
        RECT 519.400 234.400 520.200 234.600 ;
        RECT 513.200 233.000 514.000 233.200 ;
        RECT 517.800 233.000 518.600 233.200 ;
        RECT 513.200 232.400 518.600 233.000 ;
        RECT 519.200 233.000 521.400 233.600 ;
        RECT 519.200 231.800 519.800 233.000 ;
        RECT 520.600 232.800 521.400 233.000 ;
        RECT 523.000 233.200 524.400 234.000 ;
        RECT 523.000 232.200 523.600 233.200 ;
        RECT 515.000 231.400 519.800 231.800 ;
        RECT 510.000 231.200 519.800 231.400 ;
        RECT 521.200 231.600 523.600 232.200 ;
        RECT 510.000 231.000 515.800 231.200 ;
        RECT 510.000 230.800 515.600 231.000 ;
        RECT 505.000 230.400 505.800 230.600 ;
        RECT 506.600 229.800 507.400 230.000 ;
        RECT 503.600 229.200 507.400 229.800 ;
        RECT 503.600 229.000 504.400 229.200 ;
        RECT 488.400 228.200 490.000 228.400 ;
        RECT 486.600 227.600 490.000 228.200 ;
        RECT 491.600 227.800 502.600 228.400 ;
        RECT 491.600 227.600 493.200 227.800 ;
        RECT 486.600 227.200 487.200 227.600 ;
        RECT 485.200 226.600 487.200 227.200 ;
        RECT 487.800 226.800 488.600 227.000 ;
        RECT 485.200 226.400 486.800 226.600 ;
        RECT 487.800 226.200 490.000 226.800 ;
        RECT 484.000 222.200 485.600 225.800 ;
        RECT 489.200 222.200 490.000 226.200 ;
        RECT 490.800 222.200 491.600 227.000 ;
        RECT 495.800 225.600 496.400 227.800 ;
        RECT 501.400 227.600 502.200 227.800 ;
        RECT 508.400 227.200 509.200 230.600 ;
        RECT 516.400 230.200 517.200 230.400 ;
        RECT 512.200 229.600 517.200 230.200 ;
        RECT 512.200 229.400 513.000 229.600 ;
        RECT 514.800 229.400 515.600 229.600 ;
        RECT 513.800 228.400 514.600 228.600 ;
        RECT 521.200 228.400 521.800 231.600 ;
        RECT 527.600 231.200 528.400 239.800 ;
        RECT 529.200 232.400 530.000 239.800 ;
        RECT 529.200 231.800 531.400 232.400 ;
        RECT 524.200 230.600 528.400 231.200 ;
        RECT 524.200 230.400 525.000 230.600 ;
        RECT 525.800 229.800 526.600 230.000 ;
        RECT 522.800 229.200 526.600 229.800 ;
        RECT 522.800 229.000 523.600 229.200 ;
        RECT 510.800 227.800 521.800 228.400 ;
        RECT 510.800 227.600 512.400 227.800 ;
        RECT 505.400 226.600 509.200 227.200 ;
        RECT 505.400 226.400 506.200 226.600 ;
        RECT 494.000 224.200 494.800 225.000 ;
        RECT 495.600 224.800 496.400 225.600 ;
        RECT 497.400 225.400 498.200 225.600 ;
        RECT 497.400 224.800 500.200 225.400 ;
        RECT 499.600 224.200 500.200 224.800 ;
        RECT 503.600 224.200 504.400 225.000 ;
        RECT 494.000 223.600 496.000 224.200 ;
        RECT 495.200 222.200 496.000 223.600 ;
        RECT 499.600 222.200 500.400 224.200 ;
        RECT 503.600 223.600 505.000 224.200 ;
        RECT 503.800 222.200 505.000 223.600 ;
        RECT 508.400 222.200 509.200 226.600 ;
        RECT 510.000 222.200 510.800 227.000 ;
        RECT 515.000 225.600 515.600 227.800 ;
        RECT 520.600 227.600 521.400 227.800 ;
        RECT 527.600 227.200 528.400 230.600 ;
        RECT 530.800 231.200 531.400 231.800 ;
        RECT 534.000 231.400 534.800 239.800 ;
        RECT 538.400 236.400 539.200 239.800 ;
        RECT 537.200 235.800 539.200 236.400 ;
        RECT 542.800 235.800 543.600 239.800 ;
        RECT 547.000 235.800 548.200 239.800 ;
        RECT 537.200 235.000 538.000 235.800 ;
        RECT 542.800 235.200 543.400 235.800 ;
        RECT 540.600 234.600 544.200 235.200 ;
        RECT 546.800 235.000 547.600 235.800 ;
        RECT 540.600 234.400 541.400 234.600 ;
        RECT 543.400 234.400 544.200 234.600 ;
        RECT 537.200 233.000 538.000 233.200 ;
        RECT 541.800 233.000 542.600 233.200 ;
        RECT 537.200 232.400 542.600 233.000 ;
        RECT 543.200 233.000 545.400 233.600 ;
        RECT 543.200 231.800 543.800 233.000 ;
        RECT 544.600 232.800 545.400 233.000 ;
        RECT 547.000 233.200 548.400 234.000 ;
        RECT 547.000 232.200 547.600 233.200 ;
        RECT 539.000 231.400 543.800 231.800 ;
        RECT 534.000 231.200 543.800 231.400 ;
        RECT 545.200 231.600 547.600 232.200 ;
        RECT 530.800 230.400 532.000 231.200 ;
        RECT 534.000 231.000 539.800 231.200 ;
        RECT 534.000 230.800 539.600 231.000 ;
        RECT 529.200 228.800 530.000 230.400 ;
        RECT 530.800 227.400 531.400 230.400 ;
        RECT 540.400 230.200 541.200 230.400 ;
        RECT 536.200 229.600 541.200 230.200 ;
        RECT 543.600 230.300 544.400 230.400 ;
        RECT 545.200 230.300 545.800 231.600 ;
        RECT 551.600 231.200 552.400 239.800 ;
        RECT 548.200 230.600 552.400 231.200 ;
        RECT 553.200 231.400 554.000 239.800 ;
        RECT 557.600 236.400 558.400 239.800 ;
        RECT 556.400 235.800 558.400 236.400 ;
        RECT 562.000 235.800 562.800 239.800 ;
        RECT 566.200 235.800 567.400 239.800 ;
        RECT 556.400 235.000 557.200 235.800 ;
        RECT 562.000 235.200 562.600 235.800 ;
        RECT 559.800 234.600 563.400 235.200 ;
        RECT 566.000 235.000 566.800 235.800 ;
        RECT 559.800 234.400 560.600 234.600 ;
        RECT 562.600 234.400 563.400 234.600 ;
        RECT 556.400 233.000 557.200 233.200 ;
        RECT 561.000 233.000 561.800 233.200 ;
        RECT 556.400 232.400 561.800 233.000 ;
        RECT 562.400 233.000 564.600 233.600 ;
        RECT 562.400 231.800 563.000 233.000 ;
        RECT 563.800 232.800 564.600 233.000 ;
        RECT 566.200 233.200 567.600 234.000 ;
        RECT 566.200 232.200 566.800 233.200 ;
        RECT 558.200 231.400 563.000 231.800 ;
        RECT 553.200 231.200 563.000 231.400 ;
        RECT 564.400 231.600 566.800 232.200 ;
        RECT 553.200 231.000 559.000 231.200 ;
        RECT 553.200 230.800 558.800 231.000 ;
        RECT 548.200 230.400 549.000 230.600 ;
        RECT 543.600 229.700 545.900 230.300 ;
        RECT 549.800 229.800 550.600 230.000 ;
        RECT 543.600 229.600 544.400 229.700 ;
        RECT 536.200 229.400 537.000 229.600 ;
        RECT 538.800 229.400 539.600 229.600 ;
        RECT 537.800 228.400 538.600 228.600 ;
        RECT 545.200 228.400 545.800 229.700 ;
        RECT 546.800 229.200 550.600 229.800 ;
        RECT 546.800 229.000 547.600 229.200 ;
        RECT 534.800 227.800 545.800 228.400 ;
        RECT 534.800 227.600 536.400 227.800 ;
        RECT 524.600 226.600 528.400 227.200 ;
        RECT 524.600 226.400 525.400 226.600 ;
        RECT 513.200 224.200 514.000 225.000 ;
        RECT 514.800 224.800 515.600 225.600 ;
        RECT 516.600 225.400 517.400 225.600 ;
        RECT 516.600 224.800 519.400 225.400 ;
        RECT 518.800 224.200 519.400 224.800 ;
        RECT 522.800 224.200 523.600 225.000 ;
        RECT 513.200 223.600 515.200 224.200 ;
        RECT 514.400 222.200 515.200 223.600 ;
        RECT 518.800 222.200 519.600 224.200 ;
        RECT 522.800 223.600 524.200 224.200 ;
        RECT 523.000 222.200 524.200 223.600 ;
        RECT 527.600 222.200 528.400 226.600 ;
        RECT 529.200 226.800 531.400 227.400 ;
        RECT 529.200 222.200 530.000 226.800 ;
        RECT 534.000 222.200 534.800 227.000 ;
        RECT 539.000 225.600 539.600 227.800 ;
        RECT 544.600 227.600 545.400 227.800 ;
        RECT 551.600 227.200 552.400 230.600 ;
        RECT 559.600 230.200 560.400 230.400 ;
        RECT 555.400 229.600 560.400 230.200 ;
        RECT 555.400 229.400 556.200 229.600 ;
        RECT 558.000 229.400 558.800 229.600 ;
        RECT 557.000 228.400 557.800 228.600 ;
        RECT 564.400 228.400 565.000 231.600 ;
        RECT 570.800 231.200 571.600 239.800 ;
        RECT 572.400 232.400 573.200 239.800 ;
        RECT 577.200 232.400 578.000 239.800 ;
        RECT 572.400 231.800 574.600 232.400 ;
        RECT 577.200 231.800 579.400 232.400 ;
        RECT 567.400 230.600 571.600 231.200 ;
        RECT 567.400 230.400 568.200 230.600 ;
        RECT 569.000 229.800 569.800 230.000 ;
        RECT 566.000 229.200 569.800 229.800 ;
        RECT 566.000 229.000 566.800 229.200 ;
        RECT 554.000 227.800 565.200 228.400 ;
        RECT 554.000 227.600 555.600 227.800 ;
        RECT 548.600 226.600 552.400 227.200 ;
        RECT 548.600 226.400 549.400 226.600 ;
        RECT 537.200 224.200 538.000 225.000 ;
        RECT 538.800 224.800 539.600 225.600 ;
        RECT 540.600 225.400 541.400 225.600 ;
        RECT 540.600 224.800 543.400 225.400 ;
        RECT 542.800 224.200 543.400 224.800 ;
        RECT 546.800 224.200 547.600 225.000 ;
        RECT 537.200 223.600 539.200 224.200 ;
        RECT 538.400 222.200 539.200 223.600 ;
        RECT 542.800 222.200 543.600 224.200 ;
        RECT 546.800 223.600 548.200 224.200 ;
        RECT 547.000 222.200 548.200 223.600 ;
        RECT 551.600 222.200 552.400 226.600 ;
        RECT 553.200 222.200 554.000 227.000 ;
        RECT 558.200 225.600 558.800 227.800 ;
        RECT 563.800 227.600 565.200 227.800 ;
        RECT 570.800 227.200 571.600 230.600 ;
        RECT 574.000 231.200 574.600 231.800 ;
        RECT 578.800 231.200 579.400 231.800 ;
        RECT 574.000 230.400 575.200 231.200 ;
        RECT 578.800 230.400 580.000 231.200 ;
        RECT 572.400 228.800 573.200 230.400 ;
        RECT 574.000 227.400 574.600 230.400 ;
        RECT 577.200 228.800 578.000 230.400 ;
        RECT 578.800 227.400 579.400 230.400 ;
        RECT 567.800 226.600 571.600 227.200 ;
        RECT 567.800 226.400 568.600 226.600 ;
        RECT 556.400 224.200 557.200 225.000 ;
        RECT 558.000 224.800 558.800 225.600 ;
        RECT 559.800 225.400 560.600 225.600 ;
        RECT 559.800 224.800 562.600 225.400 ;
        RECT 562.000 224.200 562.600 224.800 ;
        RECT 566.000 224.200 566.800 225.000 ;
        RECT 556.400 223.600 558.400 224.200 ;
        RECT 557.600 222.200 558.400 223.600 ;
        RECT 562.000 222.200 562.800 224.200 ;
        RECT 566.000 223.600 567.400 224.200 ;
        RECT 566.200 222.200 567.400 223.600 ;
        RECT 570.800 222.200 571.600 226.600 ;
        RECT 572.400 226.800 574.600 227.400 ;
        RECT 577.200 226.800 579.400 227.400 ;
        RECT 572.400 222.200 573.200 226.800 ;
        RECT 577.200 222.200 578.000 226.800 ;
        RECT 1.200 215.000 2.000 219.800 ;
        RECT 5.600 218.400 6.400 219.800 ;
        RECT 4.400 217.800 6.400 218.400 ;
        RECT 10.000 217.800 10.800 219.800 ;
        RECT 14.200 218.400 15.400 219.800 ;
        RECT 14.000 217.800 15.400 218.400 ;
        RECT 4.400 217.000 5.200 217.800 ;
        RECT 10.000 217.200 10.600 217.800 ;
        RECT 6.000 216.400 6.800 217.200 ;
        RECT 7.800 216.600 10.600 217.200 ;
        RECT 14.000 217.000 14.800 217.800 ;
        RECT 7.800 216.400 8.600 216.600 ;
        RECT 2.000 214.200 3.600 214.400 ;
        RECT 6.200 214.200 6.800 216.400 ;
        RECT 15.800 215.400 16.600 215.600 ;
        RECT 18.800 215.400 19.600 219.800 ;
        RECT 15.800 214.800 19.600 215.400 ;
        RECT 20.400 215.000 21.200 219.800 ;
        RECT 24.800 218.400 25.600 219.800 ;
        RECT 23.600 217.800 25.600 218.400 ;
        RECT 29.200 217.800 30.000 219.800 ;
        RECT 33.400 218.400 34.600 219.800 ;
        RECT 33.200 217.800 34.600 218.400 ;
        RECT 23.600 217.000 24.400 217.800 ;
        RECT 29.200 217.200 29.800 217.800 ;
        RECT 25.200 216.400 26.000 217.200 ;
        RECT 27.000 216.600 29.800 217.200 ;
        RECT 33.200 217.000 34.000 217.800 ;
        RECT 27.000 216.400 27.800 216.600 ;
        RECT 11.800 214.200 12.600 214.400 ;
        RECT 2.000 213.600 13.000 214.200 ;
        RECT 5.000 213.400 5.800 213.600 ;
        RECT 3.400 212.400 4.200 212.600 ;
        RECT 6.000 212.400 6.800 212.600 ;
        RECT 12.400 212.400 13.000 213.600 ;
        RECT 14.000 212.800 14.800 213.000 ;
        RECT 3.400 211.800 8.400 212.400 ;
        RECT 7.600 211.600 8.400 211.800 ;
        RECT 12.400 211.600 13.200 212.400 ;
        RECT 14.000 212.200 17.800 212.800 ;
        RECT 17.000 212.000 17.800 212.200 ;
        RECT 1.200 211.000 6.800 211.200 ;
        RECT 1.200 210.800 7.000 211.000 ;
        RECT 1.200 210.600 11.000 210.800 ;
        RECT 1.200 202.200 2.000 210.600 ;
        RECT 6.200 210.200 11.000 210.600 ;
        RECT 4.400 209.000 9.800 209.600 ;
        RECT 4.400 208.800 5.200 209.000 ;
        RECT 9.000 208.800 9.800 209.000 ;
        RECT 10.400 209.000 11.000 210.200 ;
        RECT 12.400 210.400 13.000 211.600 ;
        RECT 15.400 211.400 16.200 211.600 ;
        RECT 18.800 211.400 19.600 214.800 ;
        RECT 21.200 214.200 22.800 214.400 ;
        RECT 25.400 214.200 26.000 216.400 ;
        RECT 35.000 215.400 35.800 215.600 ;
        RECT 38.000 215.400 38.800 219.800 ;
        RECT 35.000 214.800 38.800 215.400 ;
        RECT 31.000 214.200 31.800 214.400 ;
        RECT 21.200 213.600 32.200 214.200 ;
        RECT 24.200 213.400 25.000 213.600 ;
        RECT 22.600 212.400 23.400 212.600 ;
        RECT 31.600 212.400 32.200 213.600 ;
        RECT 33.200 212.800 34.000 213.000 ;
        RECT 22.600 211.800 27.600 212.400 ;
        RECT 26.800 211.600 27.600 211.800 ;
        RECT 31.600 211.600 32.400 212.400 ;
        RECT 33.200 212.200 37.000 212.800 ;
        RECT 36.200 212.000 37.000 212.200 ;
        RECT 15.400 210.800 19.600 211.400 ;
        RECT 12.400 209.800 14.800 210.400 ;
        RECT 11.800 209.000 12.600 209.200 ;
        RECT 10.400 208.400 12.600 209.000 ;
        RECT 14.200 208.800 14.800 209.800 ;
        RECT 14.200 208.000 15.600 208.800 ;
        RECT 7.800 207.400 8.600 207.600 ;
        RECT 10.600 207.400 11.400 207.600 ;
        RECT 4.400 206.200 5.200 207.000 ;
        RECT 7.800 206.800 11.400 207.400 ;
        RECT 10.000 206.200 10.600 206.800 ;
        RECT 14.000 206.200 14.800 207.000 ;
        RECT 4.400 205.600 6.400 206.200 ;
        RECT 5.600 202.200 6.400 205.600 ;
        RECT 10.000 202.200 10.800 206.200 ;
        RECT 14.200 202.200 15.400 206.200 ;
        RECT 18.800 202.200 19.600 210.800 ;
        RECT 20.400 211.000 26.000 211.200 ;
        RECT 20.400 210.800 26.200 211.000 ;
        RECT 20.400 210.600 30.200 210.800 ;
        RECT 20.400 202.200 21.200 210.600 ;
        RECT 25.400 210.200 30.200 210.600 ;
        RECT 23.600 209.000 29.000 209.600 ;
        RECT 23.600 208.800 24.400 209.000 ;
        RECT 28.200 208.800 29.000 209.000 ;
        RECT 29.600 209.000 30.200 210.200 ;
        RECT 31.600 210.400 32.200 211.600 ;
        RECT 34.600 211.400 35.400 211.600 ;
        RECT 38.000 211.400 38.800 214.800 ;
        RECT 34.600 210.800 38.800 211.400 ;
        RECT 31.600 209.800 34.000 210.400 ;
        RECT 31.000 209.000 31.800 209.200 ;
        RECT 29.600 208.400 31.800 209.000 ;
        RECT 33.400 208.800 34.000 209.800 ;
        RECT 33.400 208.000 34.800 208.800 ;
        RECT 27.000 207.400 27.800 207.600 ;
        RECT 29.800 207.400 30.600 207.600 ;
        RECT 23.600 206.200 24.400 207.000 ;
        RECT 27.000 206.800 30.600 207.400 ;
        RECT 29.200 206.200 29.800 206.800 ;
        RECT 33.200 206.200 34.000 207.000 ;
        RECT 23.600 205.600 25.600 206.200 ;
        RECT 24.800 202.200 25.600 205.600 ;
        RECT 29.200 202.200 30.000 206.200 ;
        RECT 33.400 202.200 34.600 206.200 ;
        RECT 38.000 202.200 38.800 210.800 ;
        RECT 39.600 215.400 40.400 219.800 ;
        RECT 43.800 218.400 45.000 219.800 ;
        RECT 43.800 217.800 45.200 218.400 ;
        RECT 48.400 217.800 49.200 219.800 ;
        RECT 52.800 218.400 53.600 219.800 ;
        RECT 52.800 217.800 54.800 218.400 ;
        RECT 44.400 217.000 45.200 217.800 ;
        RECT 48.600 217.200 49.200 217.800 ;
        RECT 48.600 216.600 51.400 217.200 ;
        RECT 50.600 216.400 51.400 216.600 ;
        RECT 52.400 216.400 53.200 217.200 ;
        RECT 54.000 217.000 54.800 217.800 ;
        RECT 42.600 215.400 43.400 215.600 ;
        RECT 39.600 214.800 43.400 215.400 ;
        RECT 39.600 211.400 40.400 214.800 ;
        RECT 46.600 214.200 47.400 214.400 ;
        RECT 52.400 214.200 53.000 216.400 ;
        RECT 57.200 215.000 58.000 219.800 ;
        RECT 58.800 215.000 59.600 219.800 ;
        RECT 63.200 218.400 64.000 219.800 ;
        RECT 62.000 217.800 64.000 218.400 ;
        RECT 67.600 217.800 68.400 219.800 ;
        RECT 71.800 218.400 73.000 219.800 ;
        RECT 71.600 217.800 73.000 218.400 ;
        RECT 62.000 217.000 62.800 217.800 ;
        RECT 67.600 217.200 68.200 217.800 ;
        RECT 63.600 216.400 64.400 217.200 ;
        RECT 65.400 216.600 68.200 217.200 ;
        RECT 71.600 217.000 72.400 217.800 ;
        RECT 65.400 216.400 66.200 216.600 ;
        RECT 55.600 214.200 57.200 214.400 ;
        RECT 46.200 213.600 57.200 214.200 ;
        RECT 59.600 214.200 61.200 214.400 ;
        RECT 63.800 214.200 64.400 216.400 ;
        RECT 73.400 215.400 74.200 215.600 ;
        RECT 76.400 215.400 77.200 219.800 ;
        RECT 73.400 214.800 77.200 215.400 ;
        RECT 69.400 214.200 70.200 214.400 ;
        RECT 59.600 213.600 70.600 214.200 ;
        RECT 44.400 212.800 45.200 213.000 ;
        RECT 41.400 212.200 45.200 212.800 ;
        RECT 41.400 212.000 42.200 212.200 ;
        RECT 43.000 211.400 43.800 211.600 ;
        RECT 39.600 210.800 43.800 211.400 ;
        RECT 39.600 202.200 40.400 210.800 ;
        RECT 46.200 210.400 46.800 213.600 ;
        RECT 53.400 213.400 54.200 213.600 ;
        RECT 62.600 213.400 63.400 213.600 ;
        RECT 52.400 212.400 53.200 212.600 ;
        RECT 55.000 212.400 55.800 212.600 ;
        RECT 50.800 211.800 55.800 212.400 ;
        RECT 61.000 212.400 61.800 212.600 ;
        RECT 70.000 212.400 70.600 213.600 ;
        RECT 71.600 212.800 72.400 213.000 ;
        RECT 61.000 211.800 66.000 212.400 ;
        RECT 50.800 211.600 51.600 211.800 ;
        RECT 65.200 211.600 66.000 211.800 ;
        RECT 70.000 211.600 70.800 212.400 ;
        RECT 71.600 212.200 75.400 212.800 ;
        RECT 74.600 212.000 75.400 212.200 ;
        RECT 52.400 211.000 58.000 211.200 ;
        RECT 52.200 210.800 58.000 211.000 ;
        RECT 44.400 209.800 46.800 210.400 ;
        RECT 48.200 210.600 58.000 210.800 ;
        RECT 48.200 210.200 53.000 210.600 ;
        RECT 44.400 208.800 45.000 209.800 ;
        RECT 43.600 208.000 45.000 208.800 ;
        RECT 46.600 209.000 47.400 209.200 ;
        RECT 48.200 209.000 48.800 210.200 ;
        RECT 46.600 208.400 48.800 209.000 ;
        RECT 49.400 209.000 54.800 209.600 ;
        RECT 49.400 208.800 50.200 209.000 ;
        RECT 54.000 208.800 54.800 209.000 ;
        RECT 47.800 207.400 48.600 207.600 ;
        RECT 50.600 207.400 51.400 207.600 ;
        RECT 44.400 206.200 45.200 207.000 ;
        RECT 47.800 206.800 51.400 207.400 ;
        RECT 48.600 206.200 49.200 206.800 ;
        RECT 54.000 206.200 54.800 207.000 ;
        RECT 43.800 202.200 45.000 206.200 ;
        RECT 48.400 202.200 49.200 206.200 ;
        RECT 52.800 205.600 54.800 206.200 ;
        RECT 52.800 202.200 53.600 205.600 ;
        RECT 57.200 202.200 58.000 210.600 ;
        RECT 58.800 211.000 64.400 211.200 ;
        RECT 58.800 210.800 64.600 211.000 ;
        RECT 58.800 210.600 68.600 210.800 ;
        RECT 58.800 202.200 59.600 210.600 ;
        RECT 63.800 210.200 68.600 210.600 ;
        RECT 62.000 209.000 67.400 209.600 ;
        RECT 62.000 208.800 62.800 209.000 ;
        RECT 66.600 208.800 67.400 209.000 ;
        RECT 68.000 209.000 68.600 210.200 ;
        RECT 70.000 210.400 70.600 211.600 ;
        RECT 73.000 211.400 73.800 211.600 ;
        RECT 76.400 211.400 77.200 214.800 ;
        RECT 73.000 210.800 77.200 211.400 ;
        RECT 70.000 209.800 72.400 210.400 ;
        RECT 69.400 209.000 70.200 209.200 ;
        RECT 68.000 208.400 70.200 209.000 ;
        RECT 71.800 208.800 72.400 209.800 ;
        RECT 71.800 208.000 73.200 208.800 ;
        RECT 65.400 207.400 66.200 207.600 ;
        RECT 68.200 207.400 69.000 207.600 ;
        RECT 62.000 206.200 62.800 207.000 ;
        RECT 65.400 206.800 69.000 207.400 ;
        RECT 67.600 206.200 68.200 206.800 ;
        RECT 71.600 206.200 72.400 207.000 ;
        RECT 62.000 205.600 64.000 206.200 ;
        RECT 63.200 202.200 64.000 205.600 ;
        RECT 67.600 202.200 68.400 206.200 ;
        RECT 71.800 202.200 73.000 206.200 ;
        RECT 76.400 202.200 77.200 210.800 ;
        RECT 78.000 215.400 78.800 219.800 ;
        RECT 82.200 218.400 83.400 219.800 ;
        RECT 82.200 217.800 83.600 218.400 ;
        RECT 86.800 217.800 87.600 219.800 ;
        RECT 91.200 218.400 92.000 219.800 ;
        RECT 91.200 217.800 93.200 218.400 ;
        RECT 82.800 217.000 83.600 217.800 ;
        RECT 87.000 217.200 87.600 217.800 ;
        RECT 87.000 216.600 89.800 217.200 ;
        RECT 89.000 216.400 89.800 216.600 ;
        RECT 90.800 216.400 91.600 217.200 ;
        RECT 92.400 217.000 93.200 217.800 ;
        RECT 81.000 215.400 81.800 215.600 ;
        RECT 78.000 214.800 81.800 215.400 ;
        RECT 78.000 211.400 78.800 214.800 ;
        RECT 85.000 214.200 85.800 214.400 ;
        RECT 90.800 214.200 91.400 216.400 ;
        RECT 95.600 215.000 96.400 219.800 ;
        RECT 98.800 215.200 99.600 219.800 ;
        RECT 102.000 215.200 102.800 219.800 ;
        RECT 105.200 215.200 106.000 219.800 ;
        RECT 108.400 215.200 109.200 219.800 ;
        RECT 97.200 214.400 99.600 215.200 ;
        RECT 100.600 214.400 102.800 215.200 ;
        RECT 103.800 214.400 106.000 215.200 ;
        RECT 107.400 214.400 109.200 215.200 ;
        RECT 111.600 215.400 112.400 219.800 ;
        RECT 115.800 218.400 117.000 219.800 ;
        RECT 115.800 217.800 117.200 218.400 ;
        RECT 120.400 217.800 121.200 219.800 ;
        RECT 124.800 218.400 125.600 219.800 ;
        RECT 124.800 217.800 126.800 218.400 ;
        RECT 116.400 217.000 117.200 217.800 ;
        RECT 120.600 217.200 121.200 217.800 ;
        RECT 120.600 216.600 123.400 217.200 ;
        RECT 122.600 216.400 123.400 216.600 ;
        RECT 124.400 216.400 125.200 217.200 ;
        RECT 126.000 217.000 126.800 217.800 ;
        RECT 114.600 215.400 115.400 215.600 ;
        RECT 111.600 214.800 115.400 215.400 ;
        RECT 94.000 214.200 95.600 214.400 ;
        RECT 84.600 213.600 95.600 214.200 ;
        RECT 82.800 212.800 83.600 213.000 ;
        RECT 79.800 212.200 83.600 212.800 ;
        RECT 79.800 212.000 80.600 212.200 ;
        RECT 81.400 211.400 82.200 211.600 ;
        RECT 78.000 210.800 82.200 211.400 ;
        RECT 78.000 202.200 78.800 210.800 ;
        RECT 84.600 210.400 85.200 213.600 ;
        RECT 91.800 213.400 92.600 213.600 ;
        RECT 90.800 212.400 91.600 212.600 ;
        RECT 93.400 212.400 94.200 212.600 ;
        RECT 89.200 211.800 94.200 212.400 ;
        RECT 89.200 211.600 90.000 211.800 ;
        RECT 97.200 211.600 98.000 214.400 ;
        RECT 100.600 213.800 101.400 214.400 ;
        RECT 103.800 213.800 104.600 214.400 ;
        RECT 107.400 213.800 108.200 214.400 ;
        RECT 98.800 213.000 101.400 213.800 ;
        RECT 102.200 213.000 104.600 213.800 ;
        RECT 105.600 213.000 108.200 213.800 ;
        RECT 100.600 211.600 101.400 213.000 ;
        RECT 103.800 211.600 104.600 213.000 ;
        RECT 107.400 211.600 108.200 213.000 ;
        RECT 90.800 211.000 96.400 211.200 ;
        RECT 90.600 210.800 96.400 211.000 ;
        RECT 97.200 210.800 99.600 211.600 ;
        RECT 100.600 210.800 102.800 211.600 ;
        RECT 103.800 210.800 106.000 211.600 ;
        RECT 107.400 210.800 109.200 211.600 ;
        RECT 82.800 209.800 85.200 210.400 ;
        RECT 86.600 210.600 96.400 210.800 ;
        RECT 86.600 210.200 91.400 210.600 ;
        RECT 82.800 208.800 83.400 209.800 ;
        RECT 82.000 208.000 83.400 208.800 ;
        RECT 85.000 209.000 85.800 209.200 ;
        RECT 86.600 209.000 87.200 210.200 ;
        RECT 85.000 208.400 87.200 209.000 ;
        RECT 87.800 209.000 93.200 209.600 ;
        RECT 87.800 208.800 88.600 209.000 ;
        RECT 92.400 208.800 93.200 209.000 ;
        RECT 86.200 207.400 87.000 207.600 ;
        RECT 89.000 207.400 89.800 207.600 ;
        RECT 82.800 206.200 83.600 207.000 ;
        RECT 86.200 206.800 89.800 207.400 ;
        RECT 87.000 206.200 87.600 206.800 ;
        RECT 92.400 206.200 93.200 207.000 ;
        RECT 82.200 202.200 83.400 206.200 ;
        RECT 86.800 202.200 87.600 206.200 ;
        RECT 91.200 205.600 93.200 206.200 ;
        RECT 91.200 202.200 92.000 205.600 ;
        RECT 95.600 202.200 96.400 210.600 ;
        RECT 98.800 202.200 99.600 210.800 ;
        RECT 102.000 202.200 102.800 210.800 ;
        RECT 105.200 202.200 106.000 210.800 ;
        RECT 108.400 202.200 109.200 210.800 ;
        RECT 111.600 211.400 112.400 214.800 ;
        RECT 118.600 214.200 119.400 214.400 ;
        RECT 124.400 214.200 125.000 216.400 ;
        RECT 129.200 215.000 130.000 219.800 ;
        RECT 135.600 215.000 136.400 219.800 ;
        RECT 140.000 218.400 140.800 219.800 ;
        RECT 138.800 217.800 140.800 218.400 ;
        RECT 144.400 217.800 145.200 219.800 ;
        RECT 148.600 218.400 149.800 219.800 ;
        RECT 148.400 217.800 149.800 218.400 ;
        RECT 138.800 217.000 139.600 217.800 ;
        RECT 144.400 217.200 145.000 217.800 ;
        RECT 140.400 216.400 141.200 217.200 ;
        RECT 142.200 216.600 145.000 217.200 ;
        RECT 148.400 217.000 149.200 217.800 ;
        RECT 142.200 216.400 143.000 216.600 ;
        RECT 127.600 214.200 129.200 214.400 ;
        RECT 118.200 213.600 129.200 214.200 ;
        RECT 132.400 214.300 133.200 214.400 ;
        RECT 136.400 214.300 138.000 214.400 ;
        RECT 132.400 214.200 138.000 214.300 ;
        RECT 140.600 214.200 141.200 216.400 ;
        RECT 150.200 215.400 151.000 215.600 ;
        RECT 153.200 215.400 154.000 219.800 ;
        RECT 150.200 214.800 154.000 215.400 ;
        RECT 154.800 215.000 155.600 219.800 ;
        RECT 159.200 218.400 160.000 219.800 ;
        RECT 158.000 217.800 160.000 218.400 ;
        RECT 163.600 217.800 164.400 219.800 ;
        RECT 167.800 218.400 169.000 219.800 ;
        RECT 167.600 217.800 169.000 218.400 ;
        RECT 158.000 217.000 158.800 217.800 ;
        RECT 163.600 217.200 164.200 217.800 ;
        RECT 159.600 216.400 160.400 217.200 ;
        RECT 161.400 216.600 164.200 217.200 ;
        RECT 167.600 217.000 168.400 217.800 ;
        RECT 161.400 216.400 162.200 216.600 ;
        RECT 146.200 214.200 147.000 214.400 ;
        RECT 132.400 213.700 147.400 214.200 ;
        RECT 132.400 213.600 133.200 213.700 ;
        RECT 136.400 213.600 147.400 213.700 ;
        RECT 116.400 212.800 117.200 213.000 ;
        RECT 113.400 212.200 117.200 212.800 ;
        RECT 118.200 212.400 118.800 213.600 ;
        RECT 125.400 213.400 126.200 213.600 ;
        RECT 139.400 213.400 140.200 213.600 ;
        RECT 124.400 212.400 125.200 212.600 ;
        RECT 127.000 212.400 127.800 212.600 ;
        RECT 113.400 212.000 114.200 212.200 ;
        RECT 118.000 211.600 118.800 212.400 ;
        RECT 122.800 211.800 127.800 212.400 ;
        RECT 137.800 212.400 138.600 212.600 ;
        RECT 146.800 212.400 147.400 213.600 ;
        RECT 148.400 212.800 149.200 213.000 ;
        RECT 137.800 212.300 142.800 212.400 ;
        RECT 143.600 212.300 144.400 212.400 ;
        RECT 137.800 211.800 144.400 212.300 ;
        RECT 122.800 211.600 123.600 211.800 ;
        RECT 142.000 211.700 144.400 211.800 ;
        RECT 142.000 211.600 142.800 211.700 ;
        RECT 143.600 211.600 144.400 211.700 ;
        RECT 146.800 211.600 147.600 212.400 ;
        RECT 148.400 212.200 152.200 212.800 ;
        RECT 151.400 212.000 152.200 212.200 ;
        RECT 115.000 211.400 115.800 211.600 ;
        RECT 111.600 210.800 115.800 211.400 ;
        RECT 111.600 202.200 112.400 210.800 ;
        RECT 118.200 210.400 118.800 211.600 ;
        RECT 124.400 211.000 130.000 211.200 ;
        RECT 124.200 210.800 130.000 211.000 ;
        RECT 116.400 209.800 118.800 210.400 ;
        RECT 120.200 210.600 130.000 210.800 ;
        RECT 120.200 210.200 125.000 210.600 ;
        RECT 116.400 208.800 117.000 209.800 ;
        RECT 115.600 208.000 117.000 208.800 ;
        RECT 118.600 209.000 119.400 209.200 ;
        RECT 120.200 209.000 120.800 210.200 ;
        RECT 118.600 208.400 120.800 209.000 ;
        RECT 121.400 209.000 126.800 209.600 ;
        RECT 121.400 208.800 122.200 209.000 ;
        RECT 126.000 208.800 126.800 209.000 ;
        RECT 119.800 207.400 120.600 207.600 ;
        RECT 122.600 207.400 123.400 207.600 ;
        RECT 116.400 206.200 117.200 207.000 ;
        RECT 119.800 206.800 123.400 207.400 ;
        RECT 120.600 206.200 121.200 206.800 ;
        RECT 126.000 206.200 126.800 207.000 ;
        RECT 115.800 202.200 117.000 206.200 ;
        RECT 120.400 202.200 121.200 206.200 ;
        RECT 124.800 205.600 126.800 206.200 ;
        RECT 124.800 202.200 125.600 205.600 ;
        RECT 129.200 202.200 130.000 210.600 ;
        RECT 135.600 211.000 141.200 211.200 ;
        RECT 135.600 210.800 141.400 211.000 ;
        RECT 135.600 210.600 145.400 210.800 ;
        RECT 135.600 202.200 136.400 210.600 ;
        RECT 140.600 210.200 145.400 210.600 ;
        RECT 138.800 209.000 144.200 209.600 ;
        RECT 138.800 208.800 139.600 209.000 ;
        RECT 143.400 208.800 144.200 209.000 ;
        RECT 144.800 209.000 145.400 210.200 ;
        RECT 146.800 210.400 147.400 211.600 ;
        RECT 149.800 211.400 150.600 211.600 ;
        RECT 153.200 211.400 154.000 214.800 ;
        RECT 155.600 214.200 157.200 214.400 ;
        RECT 159.800 214.200 160.400 216.400 ;
        RECT 169.400 215.400 170.200 215.600 ;
        RECT 172.400 215.400 173.200 219.800 ;
        RECT 174.000 215.600 174.800 217.200 ;
        RECT 175.600 216.300 176.400 219.800 ;
        RECT 178.800 217.800 179.600 219.800 ;
        RECT 177.200 216.300 178.000 217.200 ;
        RECT 175.600 215.700 178.000 216.300 ;
        RECT 169.400 214.800 173.200 215.400 ;
        RECT 165.400 214.200 166.200 214.400 ;
        RECT 155.600 213.600 166.600 214.200 ;
        RECT 158.600 213.400 159.400 213.600 ;
        RECT 157.000 212.400 157.800 212.600 ;
        RECT 166.000 212.400 166.600 213.600 ;
        RECT 167.600 212.800 168.400 213.000 ;
        RECT 157.000 212.300 162.000 212.400 ;
        RECT 162.800 212.300 163.600 212.400 ;
        RECT 157.000 211.800 163.600 212.300 ;
        RECT 161.200 211.700 163.600 211.800 ;
        RECT 161.200 211.600 162.000 211.700 ;
        RECT 162.800 211.600 163.600 211.700 ;
        RECT 166.000 211.600 166.800 212.400 ;
        RECT 167.600 212.200 171.400 212.800 ;
        RECT 170.600 212.000 171.400 212.200 ;
        RECT 149.800 210.800 154.000 211.400 ;
        RECT 146.800 209.800 149.200 210.400 ;
        RECT 146.200 209.000 147.000 209.200 ;
        RECT 144.800 208.400 147.000 209.000 ;
        RECT 148.600 208.800 149.200 209.800 ;
        RECT 148.600 208.000 150.000 208.800 ;
        RECT 142.200 207.400 143.000 207.600 ;
        RECT 145.000 207.400 145.800 207.600 ;
        RECT 138.800 206.200 139.600 207.000 ;
        RECT 142.200 206.800 145.800 207.400 ;
        RECT 144.400 206.200 145.000 206.800 ;
        RECT 148.400 206.200 149.200 207.000 ;
        RECT 138.800 205.600 140.800 206.200 ;
        RECT 140.000 202.200 140.800 205.600 ;
        RECT 144.400 202.200 145.200 206.200 ;
        RECT 148.600 202.200 149.800 206.200 ;
        RECT 153.200 202.200 154.000 210.800 ;
        RECT 154.800 211.000 160.400 211.200 ;
        RECT 154.800 210.800 160.600 211.000 ;
        RECT 154.800 210.600 164.600 210.800 ;
        RECT 154.800 202.200 155.600 210.600 ;
        RECT 159.800 210.200 164.600 210.600 ;
        RECT 158.000 209.000 163.400 209.600 ;
        RECT 158.000 208.800 158.800 209.000 ;
        RECT 162.600 208.800 163.400 209.000 ;
        RECT 164.000 209.000 164.600 210.200 ;
        RECT 166.000 210.400 166.600 211.600 ;
        RECT 169.000 211.400 169.800 211.600 ;
        RECT 172.400 211.400 173.200 214.800 ;
        RECT 169.000 210.800 173.200 211.400 ;
        RECT 166.000 209.800 168.400 210.400 ;
        RECT 165.400 209.000 166.200 209.200 ;
        RECT 164.000 208.400 166.200 209.000 ;
        RECT 167.800 208.800 168.400 209.800 ;
        RECT 167.800 208.000 169.200 208.800 ;
        RECT 161.400 207.400 162.200 207.600 ;
        RECT 164.200 207.400 165.000 207.600 ;
        RECT 158.000 206.200 158.800 207.000 ;
        RECT 161.400 206.800 165.000 207.400 ;
        RECT 163.600 206.200 164.200 206.800 ;
        RECT 167.600 206.200 168.400 207.000 ;
        RECT 158.000 205.600 160.000 206.200 ;
        RECT 159.200 202.200 160.000 205.600 ;
        RECT 163.600 202.200 164.400 206.200 ;
        RECT 167.800 202.200 169.000 206.200 ;
        RECT 172.400 202.200 173.200 210.800 ;
        RECT 175.600 214.300 176.400 215.700 ;
        RECT 177.200 215.600 178.000 215.700 ;
        RECT 179.000 214.400 179.600 217.800 ;
        RECT 182.000 216.000 182.800 219.800 ;
        RECT 185.200 216.000 186.000 219.800 ;
        RECT 182.000 215.800 186.000 216.000 ;
        RECT 186.800 215.800 187.600 219.800 ;
        RECT 190.000 217.800 190.800 219.800 ;
        RECT 182.200 215.400 185.800 215.800 ;
        RECT 182.800 214.400 183.600 214.800 ;
        RECT 186.800 214.400 187.400 215.800 ;
        RECT 188.400 215.600 189.200 217.200 ;
        RECT 190.200 214.400 190.800 217.800 ;
        RECT 191.600 216.300 192.400 216.400 ;
        RECT 193.200 216.300 194.000 217.200 ;
        RECT 191.600 215.700 194.000 216.300 ;
        RECT 191.600 215.600 192.400 215.700 ;
        RECT 193.200 215.600 194.000 215.700 ;
        RECT 177.200 214.300 178.000 214.400 ;
        RECT 175.600 213.700 178.000 214.300 ;
        RECT 175.600 202.200 176.400 213.700 ;
        RECT 177.200 213.600 178.000 213.700 ;
        RECT 178.800 213.600 179.600 214.400 ;
        RECT 182.000 213.800 183.600 214.400 ;
        RECT 182.000 213.600 182.800 213.800 ;
        RECT 185.000 213.600 187.600 214.400 ;
        RECT 190.000 213.600 190.800 214.400 ;
        RECT 193.200 214.300 194.000 214.400 ;
        RECT 194.800 214.300 195.600 219.800 ;
        RECT 196.400 216.000 197.200 219.800 ;
        RECT 199.600 216.000 200.400 219.800 ;
        RECT 196.400 215.800 200.400 216.000 ;
        RECT 201.200 215.800 202.000 219.800 ;
        RECT 196.600 215.400 200.200 215.800 ;
        RECT 197.200 214.400 198.000 214.800 ;
        RECT 201.200 214.400 201.800 215.800 ;
        RECT 202.800 215.000 203.600 219.800 ;
        RECT 207.200 218.400 208.000 219.800 ;
        RECT 206.000 217.800 208.000 218.400 ;
        RECT 211.600 217.800 212.400 219.800 ;
        RECT 215.800 218.400 217.000 219.800 ;
        RECT 215.600 217.800 217.000 218.400 ;
        RECT 206.000 217.000 206.800 217.800 ;
        RECT 211.600 217.200 212.200 217.800 ;
        RECT 207.600 216.400 208.400 217.200 ;
        RECT 209.400 216.600 212.200 217.200 ;
        RECT 215.600 217.000 216.400 217.800 ;
        RECT 209.400 216.400 210.200 216.600 ;
        RECT 193.200 213.700 195.600 214.300 ;
        RECT 193.200 213.600 194.000 213.700 ;
        RECT 179.000 210.200 179.600 213.600 ;
        RECT 180.400 212.300 181.200 212.400 ;
        RECT 183.600 212.300 184.400 213.200 ;
        RECT 180.400 211.700 184.400 212.300 ;
        RECT 180.400 210.800 181.200 211.700 ;
        RECT 183.600 211.600 184.400 211.700 ;
        RECT 185.000 212.300 185.600 213.600 ;
        RECT 188.400 212.300 189.200 212.400 ;
        RECT 185.000 211.700 189.200 212.300 ;
        RECT 185.000 210.200 185.600 211.700 ;
        RECT 188.400 211.600 189.200 211.700 ;
        RECT 186.800 210.200 187.600 210.400 ;
        RECT 190.200 210.200 190.800 213.600 ;
        RECT 191.600 210.800 192.400 212.400 ;
        RECT 178.800 209.400 180.600 210.200 ;
        RECT 179.800 204.400 180.600 209.400 ;
        RECT 184.600 209.600 185.600 210.200 ;
        RECT 186.200 209.600 187.600 210.200 ;
        RECT 179.800 203.600 181.200 204.400 ;
        RECT 179.800 202.200 180.600 203.600 ;
        RECT 184.600 202.200 185.400 209.600 ;
        RECT 186.200 208.400 186.800 209.600 ;
        RECT 190.000 209.400 191.800 210.200 ;
        RECT 186.000 207.600 186.800 208.400 ;
        RECT 191.000 208.300 191.800 209.400 ;
        RECT 193.200 208.300 194.000 208.400 ;
        RECT 191.000 207.700 194.000 208.300 ;
        RECT 191.000 202.200 191.800 207.700 ;
        RECT 193.200 207.600 194.000 207.700 ;
        RECT 194.800 202.200 195.600 213.700 ;
        RECT 196.400 213.800 198.000 214.400 ;
        RECT 196.400 213.600 197.200 213.800 ;
        RECT 199.400 213.600 202.000 214.400 ;
        RECT 203.600 214.200 205.200 214.400 ;
        RECT 207.800 214.200 208.400 216.400 ;
        RECT 217.400 215.400 218.200 215.600 ;
        RECT 220.400 215.400 221.200 219.800 ;
        RECT 217.400 214.800 221.200 215.400 ;
        RECT 213.400 214.200 214.200 214.400 ;
        RECT 203.600 213.600 214.600 214.200 ;
        RECT 198.000 211.600 198.800 213.200 ;
        RECT 199.400 210.200 200.000 213.600 ;
        RECT 206.600 213.400 207.400 213.600 ;
        RECT 205.000 212.400 205.800 212.600 ;
        RECT 207.600 212.400 208.400 212.600 ;
        RECT 205.000 211.800 210.000 212.400 ;
        RECT 209.200 211.600 210.000 211.800 ;
        RECT 202.800 211.000 208.400 211.200 ;
        RECT 202.800 210.800 208.600 211.000 ;
        RECT 202.800 210.600 212.600 210.800 ;
        RECT 201.200 210.200 202.000 210.400 ;
        RECT 199.000 209.600 200.000 210.200 ;
        RECT 200.600 209.600 202.000 210.200 ;
        RECT 199.000 204.400 199.800 209.600 ;
        RECT 200.600 208.400 201.200 209.600 ;
        RECT 200.400 207.600 201.200 208.400 ;
        RECT 198.000 203.600 199.800 204.400 ;
        RECT 199.000 202.200 199.800 203.600 ;
        RECT 202.800 202.200 203.600 210.600 ;
        RECT 207.800 210.200 212.600 210.600 ;
        RECT 206.000 209.000 211.400 209.600 ;
        RECT 206.000 208.800 206.800 209.000 ;
        RECT 210.600 208.800 211.400 209.000 ;
        RECT 212.000 209.000 212.600 210.200 ;
        RECT 214.000 210.400 214.600 213.600 ;
        RECT 215.600 212.800 216.400 213.000 ;
        RECT 215.600 212.200 219.400 212.800 ;
        RECT 218.600 212.000 219.400 212.200 ;
        RECT 217.000 211.400 217.800 211.600 ;
        RECT 220.400 211.400 221.200 214.800 ;
        RECT 223.600 217.800 224.400 219.800 ;
        RECT 223.600 214.400 224.200 217.800 ;
        RECT 225.200 216.300 226.000 217.200 ;
        RECT 226.800 216.300 227.600 217.200 ;
        RECT 225.200 215.700 227.600 216.300 ;
        RECT 225.200 215.600 226.000 215.700 ;
        RECT 226.800 215.600 227.600 215.700 ;
        RECT 228.400 216.300 229.200 219.800 ;
        RECT 231.600 217.800 232.400 219.800 ;
        RECT 230.000 216.300 230.800 217.200 ;
        RECT 228.400 215.700 230.800 216.300 ;
        RECT 223.600 213.600 224.400 214.400 ;
        RECT 228.400 214.300 229.200 215.700 ;
        RECT 230.000 215.600 230.800 215.700 ;
        RECT 231.800 214.400 232.400 217.800 ;
        RECT 234.800 216.000 235.600 219.800 ;
        RECT 238.000 216.000 238.800 219.800 ;
        RECT 234.800 215.800 238.800 216.000 ;
        RECT 239.600 215.800 240.400 219.800 ;
        RECT 241.200 216.000 242.000 219.800 ;
        RECT 244.400 216.000 245.200 219.800 ;
        RECT 241.200 215.800 245.200 216.000 ;
        RECT 246.000 215.800 246.800 219.800 ;
        RECT 247.600 216.000 248.400 219.800 ;
        RECT 250.800 216.000 251.600 219.800 ;
        RECT 247.600 215.800 251.600 216.000 ;
        RECT 252.400 215.800 253.200 219.800 ;
        RECT 235.000 215.400 238.600 215.800 ;
        RECT 235.600 214.400 236.400 214.800 ;
        RECT 239.600 214.400 240.200 215.800 ;
        RECT 241.400 215.400 245.000 215.800 ;
        RECT 242.000 214.400 242.800 214.800 ;
        RECT 246.000 214.400 246.600 215.800 ;
        RECT 247.800 215.400 251.400 215.800 ;
        RECT 248.400 214.400 249.200 214.800 ;
        RECT 252.400 214.400 253.000 215.800 ;
        RECT 254.000 215.000 254.800 219.800 ;
        RECT 258.400 218.400 259.200 219.800 ;
        RECT 257.200 217.800 259.200 218.400 ;
        RECT 262.800 217.800 263.600 219.800 ;
        RECT 267.000 218.400 268.200 219.800 ;
        RECT 266.800 217.800 268.200 218.400 ;
        RECT 257.200 217.000 258.000 217.800 ;
        RECT 262.800 217.200 263.400 217.800 ;
        RECT 258.800 216.400 259.600 217.200 ;
        RECT 260.600 216.600 263.400 217.200 ;
        RECT 266.800 217.000 267.600 217.800 ;
        RECT 260.600 216.400 261.400 216.600 ;
        RECT 230.000 214.300 230.800 214.400 ;
        RECT 228.400 213.700 230.800 214.300 ;
        RECT 217.000 210.800 221.200 211.400 ;
        RECT 222.000 210.800 222.800 212.400 ;
        RECT 223.600 212.300 224.200 213.600 ;
        RECT 226.800 212.300 227.600 212.400 ;
        RECT 223.600 211.700 227.600 212.300 ;
        RECT 214.000 209.800 216.400 210.400 ;
        RECT 213.400 209.000 214.200 209.200 ;
        RECT 212.000 208.400 214.200 209.000 ;
        RECT 215.800 208.800 216.400 209.800 ;
        RECT 215.800 208.400 217.200 208.800 ;
        RECT 215.800 208.000 218.000 208.400 ;
        RECT 216.600 207.600 218.000 208.000 ;
        RECT 209.400 207.400 210.200 207.600 ;
        RECT 212.200 207.400 213.000 207.600 ;
        RECT 206.000 206.200 206.800 207.000 ;
        RECT 209.400 206.800 213.000 207.400 ;
        RECT 211.600 206.200 212.200 206.800 ;
        RECT 215.600 206.200 216.400 207.000 ;
        RECT 206.000 205.600 208.000 206.200 ;
        RECT 207.200 202.200 208.000 205.600 ;
        RECT 211.600 202.200 212.400 206.200 ;
        RECT 215.800 202.200 217.000 206.200 ;
        RECT 220.400 202.200 221.200 210.800 ;
        RECT 223.600 210.200 224.200 211.700 ;
        RECT 226.800 211.600 227.600 211.700 ;
        RECT 222.600 209.400 224.400 210.200 ;
        RECT 222.600 202.200 223.400 209.400 ;
        RECT 228.400 202.200 229.200 213.700 ;
        RECT 230.000 213.600 230.800 213.700 ;
        RECT 231.600 213.600 232.400 214.400 ;
        RECT 234.800 213.800 236.400 214.400 ;
        RECT 234.800 213.600 235.600 213.800 ;
        RECT 237.800 213.600 240.400 214.400 ;
        RECT 241.200 213.800 242.800 214.400 ;
        RECT 241.200 213.600 242.000 213.800 ;
        RECT 244.200 213.600 246.800 214.400 ;
        RECT 247.600 213.800 249.200 214.400 ;
        RECT 247.600 213.600 248.400 213.800 ;
        RECT 250.600 213.600 253.200 214.400 ;
        RECT 254.800 214.200 256.400 214.400 ;
        RECT 259.000 214.200 259.600 216.400 ;
        RECT 268.600 215.400 269.400 215.600 ;
        RECT 271.600 215.400 272.400 219.800 ;
        RECT 273.200 215.600 274.000 217.200 ;
        RECT 274.800 216.300 275.600 219.800 ;
        RECT 278.000 217.800 278.800 219.800 ;
        RECT 276.400 216.300 277.200 217.200 ;
        RECT 274.800 215.700 277.200 216.300 ;
        RECT 268.600 214.800 272.400 215.400 ;
        RECT 264.600 214.200 265.400 214.400 ;
        RECT 254.800 213.600 265.800 214.200 ;
        RECT 231.800 210.200 232.400 213.600 ;
        RECT 233.200 212.300 234.000 212.400 ;
        RECT 236.400 212.300 237.200 213.200 ;
        RECT 233.200 211.700 237.200 212.300 ;
        RECT 233.200 210.800 234.000 211.700 ;
        RECT 236.400 211.600 237.200 211.700 ;
        RECT 237.800 212.300 238.400 213.600 ;
        RECT 242.800 212.300 243.600 213.200 ;
        RECT 237.800 211.700 243.600 212.300 ;
        RECT 237.800 210.200 238.400 211.700 ;
        RECT 242.800 211.600 243.600 211.700 ;
        RECT 239.600 210.200 240.400 210.400 ;
        RECT 244.200 210.200 244.800 213.600 ;
        RECT 249.200 211.600 250.000 213.200 ;
        RECT 246.000 210.200 246.800 210.400 ;
        RECT 250.600 210.200 251.200 213.600 ;
        RECT 257.800 213.400 258.600 213.600 ;
        RECT 256.200 212.400 257.000 212.600 ;
        RECT 258.800 212.400 259.600 212.600 ;
        RECT 265.200 212.400 265.800 213.600 ;
        RECT 266.800 212.800 267.600 213.000 ;
        RECT 256.200 211.800 261.200 212.400 ;
        RECT 260.400 211.600 261.200 211.800 ;
        RECT 265.200 211.600 266.000 212.400 ;
        RECT 266.800 212.200 270.600 212.800 ;
        RECT 269.800 212.000 270.600 212.200 ;
        RECT 254.000 211.000 259.600 211.200 ;
        RECT 254.000 210.800 259.800 211.000 ;
        RECT 254.000 210.600 263.800 210.800 ;
        RECT 252.400 210.200 253.200 210.400 ;
        RECT 231.600 209.400 233.400 210.200 ;
        RECT 232.600 208.400 233.400 209.400 ;
        RECT 237.400 209.600 238.400 210.200 ;
        RECT 239.000 209.600 240.400 210.200 ;
        RECT 243.800 209.600 244.800 210.200 ;
        RECT 245.400 209.600 246.800 210.200 ;
        RECT 250.200 209.600 251.200 210.200 ;
        RECT 251.800 209.600 253.200 210.200 ;
        RECT 232.600 207.600 234.000 208.400 ;
        RECT 232.600 202.200 233.400 207.600 ;
        RECT 237.400 202.200 238.200 209.600 ;
        RECT 239.000 208.400 239.600 209.600 ;
        RECT 238.800 207.600 239.600 208.400 ;
        RECT 243.800 202.200 244.600 209.600 ;
        RECT 245.400 208.400 246.000 209.600 ;
        RECT 250.200 208.400 251.000 209.600 ;
        RECT 251.800 208.400 252.400 209.600 ;
        RECT 245.200 207.600 246.000 208.400 ;
        RECT 249.200 207.600 251.000 208.400 ;
        RECT 251.600 207.600 252.400 208.400 ;
        RECT 250.200 202.200 251.000 207.600 ;
        RECT 254.000 202.200 254.800 210.600 ;
        RECT 259.000 210.200 263.800 210.600 ;
        RECT 257.200 209.000 262.600 209.600 ;
        RECT 257.200 208.800 258.000 209.000 ;
        RECT 261.800 208.800 262.600 209.000 ;
        RECT 263.200 209.000 263.800 210.200 ;
        RECT 265.200 210.400 265.800 211.600 ;
        RECT 268.200 211.400 269.000 211.600 ;
        RECT 271.600 211.400 272.400 214.800 ;
        RECT 268.200 210.800 272.400 211.400 ;
        RECT 265.200 209.800 267.600 210.400 ;
        RECT 264.600 209.000 265.400 209.200 ;
        RECT 263.200 208.400 265.400 209.000 ;
        RECT 267.000 208.800 267.600 209.800 ;
        RECT 267.000 208.000 268.400 208.800 ;
        RECT 260.600 207.400 261.400 207.600 ;
        RECT 263.400 207.400 264.200 207.600 ;
        RECT 257.200 206.200 258.000 207.000 ;
        RECT 260.600 206.800 264.200 207.400 ;
        RECT 262.800 206.200 263.400 206.800 ;
        RECT 266.800 206.200 267.600 207.000 ;
        RECT 257.200 205.600 259.200 206.200 ;
        RECT 258.400 202.200 259.200 205.600 ;
        RECT 262.800 202.200 263.600 206.200 ;
        RECT 267.000 202.200 268.200 206.200 ;
        RECT 271.600 202.200 272.400 210.800 ;
        RECT 274.800 202.200 275.600 215.700 ;
        RECT 276.400 215.600 277.200 215.700 ;
        RECT 278.200 214.400 278.800 217.800 ;
        RECT 283.800 218.400 284.600 219.800 ;
        RECT 283.800 217.600 285.200 218.400 ;
        RECT 283.800 216.400 284.600 217.600 ;
        RECT 282.800 215.800 284.600 216.400 ;
        RECT 278.000 213.600 278.800 214.400 ;
        RECT 281.200 213.600 282.000 215.200 ;
        RECT 278.200 210.200 278.800 213.600 ;
        RECT 279.600 210.800 280.400 212.400 ;
        RECT 278.000 209.400 279.800 210.200 ;
        RECT 279.000 208.300 279.800 209.400 ;
        RECT 281.200 208.300 282.000 208.400 ;
        RECT 279.000 207.700 282.000 208.300 ;
        RECT 279.000 202.200 279.800 207.700 ;
        RECT 281.200 207.600 282.000 207.700 ;
        RECT 282.800 202.200 283.600 215.800 ;
        RECT 284.400 212.300 285.200 212.400 ;
        RECT 286.000 212.300 286.800 219.800 ;
        RECT 295.600 217.800 296.400 219.800 ;
        RECT 287.600 216.300 288.400 217.200 ;
        RECT 292.400 216.300 293.200 216.400 ;
        RECT 287.600 215.700 293.200 216.300 ;
        RECT 287.600 215.600 288.400 215.700 ;
        RECT 292.400 215.600 293.200 215.700 ;
        RECT 294.000 215.600 294.800 217.200 ;
        RECT 295.800 214.400 296.400 217.800 ;
        RECT 287.600 214.300 288.400 214.400 ;
        RECT 295.600 214.300 296.400 214.400 ;
        RECT 287.600 213.700 296.400 214.300 ;
        RECT 287.600 213.600 288.400 213.700 ;
        RECT 295.600 213.600 296.400 213.700 ;
        RECT 284.400 211.700 286.800 212.300 ;
        RECT 284.400 211.600 285.200 211.700 ;
        RECT 284.400 208.800 285.200 210.400 ;
        RECT 286.000 202.200 286.800 211.700 ;
        RECT 295.800 210.200 296.400 213.600 ;
        RECT 298.800 215.400 299.600 219.800 ;
        RECT 303.000 218.400 304.200 219.800 ;
        RECT 303.000 217.800 304.400 218.400 ;
        RECT 307.600 217.800 308.400 219.800 ;
        RECT 312.000 218.400 312.800 219.800 ;
        RECT 312.000 217.800 314.000 218.400 ;
        RECT 303.600 217.000 304.400 217.800 ;
        RECT 307.800 217.200 308.400 217.800 ;
        RECT 307.800 216.600 310.600 217.200 ;
        RECT 309.800 216.400 310.600 216.600 ;
        RECT 311.600 216.400 312.400 217.200 ;
        RECT 313.200 217.000 314.000 217.800 ;
        RECT 301.800 215.400 302.600 215.600 ;
        RECT 298.800 214.800 302.600 215.400 ;
        RECT 297.200 212.300 298.000 212.400 ;
        RECT 298.800 212.300 299.600 214.800 ;
        RECT 305.800 214.200 306.600 214.400 ;
        RECT 310.000 214.200 310.800 214.400 ;
        RECT 311.600 214.200 312.200 216.400 ;
        RECT 316.400 215.000 317.200 219.800 ;
        RECT 314.800 214.200 316.400 214.400 ;
        RECT 305.400 213.600 316.400 214.200 ;
        RECT 303.600 212.800 304.400 213.000 ;
        RECT 297.200 211.700 299.600 212.300 ;
        RECT 300.600 212.200 304.400 212.800 ;
        RECT 305.400 212.400 306.000 213.600 ;
        RECT 312.600 213.400 313.400 213.600 ;
        RECT 311.600 212.400 312.400 212.600 ;
        RECT 314.200 212.400 315.000 212.600 ;
        RECT 300.600 212.000 301.400 212.200 ;
        RECT 297.200 210.800 298.000 211.700 ;
        RECT 298.800 211.400 299.600 211.700 ;
        RECT 305.200 211.600 306.000 212.400 ;
        RECT 310.000 211.800 315.000 212.400 ;
        RECT 318.000 212.400 318.800 219.800 ;
        RECT 321.200 215.200 322.000 219.800 ;
        RECT 319.800 214.600 322.000 215.200 ;
        RECT 322.800 215.400 323.600 219.800 ;
        RECT 327.000 218.400 328.200 219.800 ;
        RECT 327.000 217.800 328.400 218.400 ;
        RECT 331.600 217.800 332.400 219.800 ;
        RECT 336.000 218.400 336.800 219.800 ;
        RECT 336.000 217.800 338.000 218.400 ;
        RECT 327.600 217.000 328.400 217.800 ;
        RECT 331.800 217.200 332.400 217.800 ;
        RECT 331.800 216.600 334.600 217.200 ;
        RECT 333.800 216.400 334.600 216.600 ;
        RECT 335.600 216.400 336.400 217.200 ;
        RECT 337.200 217.000 338.000 217.800 ;
        RECT 325.800 215.400 326.600 215.600 ;
        RECT 322.800 214.800 326.600 215.400 ;
        RECT 310.000 211.600 310.800 211.800 ;
        RECT 302.200 211.400 303.000 211.600 ;
        RECT 298.800 210.800 303.000 211.400 ;
        RECT 295.600 209.400 297.400 210.200 ;
        RECT 296.600 202.200 297.400 209.400 ;
        RECT 298.800 202.200 299.600 210.800 ;
        RECT 305.400 210.400 306.000 211.600 ;
        RECT 311.600 211.000 317.200 211.200 ;
        RECT 311.400 210.800 317.200 211.000 ;
        RECT 303.600 209.800 306.000 210.400 ;
        RECT 307.400 210.600 317.200 210.800 ;
        RECT 307.400 210.200 312.200 210.600 ;
        RECT 303.600 208.800 304.200 209.800 ;
        RECT 302.800 208.000 304.200 208.800 ;
        RECT 305.800 209.000 306.600 209.200 ;
        RECT 307.400 209.000 308.000 210.200 ;
        RECT 305.800 208.400 308.000 209.000 ;
        RECT 308.600 209.000 314.000 209.600 ;
        RECT 308.600 208.800 309.400 209.000 ;
        RECT 313.200 208.800 314.000 209.000 ;
        RECT 307.000 207.400 307.800 207.600 ;
        RECT 309.800 207.400 310.600 207.600 ;
        RECT 303.600 206.200 304.400 207.000 ;
        RECT 307.000 206.800 310.600 207.400 ;
        RECT 307.800 206.200 308.400 206.800 ;
        RECT 313.200 206.200 314.000 207.000 ;
        RECT 303.000 202.200 304.200 206.200 ;
        RECT 307.600 202.200 308.400 206.200 ;
        RECT 312.000 205.600 314.000 206.200 ;
        RECT 312.000 202.200 312.800 205.600 ;
        RECT 316.400 202.200 317.200 210.600 ;
        RECT 318.000 210.200 318.600 212.400 ;
        RECT 319.800 211.600 320.400 214.600 ;
        RECT 321.200 211.600 322.000 213.200 ;
        RECT 319.200 210.800 320.400 211.600 ;
        RECT 319.800 210.200 320.400 210.800 ;
        RECT 322.800 211.400 323.600 214.800 ;
        RECT 329.800 214.200 330.600 214.400 ;
        RECT 335.600 214.200 336.200 216.400 ;
        RECT 340.400 215.000 341.200 219.800 ;
        RECT 338.800 214.200 340.400 214.400 ;
        RECT 329.400 213.600 340.400 214.200 ;
        RECT 327.600 212.800 328.400 213.000 ;
        RECT 324.600 212.200 328.400 212.800 ;
        RECT 329.400 212.400 330.000 213.600 ;
        RECT 336.600 213.400 337.400 213.600 ;
        RECT 335.600 212.400 336.400 212.600 ;
        RECT 338.200 212.400 339.000 212.600 ;
        RECT 324.600 212.000 325.400 212.200 ;
        RECT 329.200 211.600 330.000 212.400 ;
        RECT 334.000 211.800 339.000 212.400 ;
        RECT 342.000 212.400 342.800 219.800 ;
        RECT 345.200 215.200 346.000 219.800 ;
        RECT 343.800 214.600 346.000 215.200 ;
        RECT 346.800 215.000 347.600 219.800 ;
        RECT 351.200 218.400 352.000 219.800 ;
        RECT 350.000 217.800 352.000 218.400 ;
        RECT 355.600 217.800 356.400 219.800 ;
        RECT 359.800 218.400 361.000 219.800 ;
        RECT 359.600 217.800 361.000 218.400 ;
        RECT 350.000 217.000 350.800 217.800 ;
        RECT 355.600 217.200 356.200 217.800 ;
        RECT 351.600 216.400 352.400 217.200 ;
        RECT 353.400 216.600 356.200 217.200 ;
        RECT 359.600 217.000 360.400 217.800 ;
        RECT 353.400 216.400 354.200 216.600 ;
        RECT 334.000 211.600 334.800 211.800 ;
        RECT 326.200 211.400 327.000 211.600 ;
        RECT 322.800 210.800 327.000 211.400 ;
        RECT 318.000 202.200 318.800 210.200 ;
        RECT 319.800 209.600 322.000 210.200 ;
        RECT 321.200 202.200 322.000 209.600 ;
        RECT 322.800 202.200 323.600 210.800 ;
        RECT 329.400 210.400 330.000 211.600 ;
        RECT 335.600 211.000 341.200 211.200 ;
        RECT 335.400 210.800 341.200 211.000 ;
        RECT 327.600 209.800 330.000 210.400 ;
        RECT 331.400 210.600 341.200 210.800 ;
        RECT 331.400 210.200 336.200 210.600 ;
        RECT 327.600 208.800 328.200 209.800 ;
        RECT 326.800 208.000 328.200 208.800 ;
        RECT 329.800 209.000 330.600 209.200 ;
        RECT 331.400 209.000 332.000 210.200 ;
        RECT 329.800 208.400 332.000 209.000 ;
        RECT 332.600 209.000 338.000 209.600 ;
        RECT 332.600 208.800 333.400 209.000 ;
        RECT 337.200 208.800 338.000 209.000 ;
        RECT 331.000 207.400 331.800 207.600 ;
        RECT 333.800 207.400 334.600 207.600 ;
        RECT 327.600 206.200 328.400 207.000 ;
        RECT 331.000 206.800 334.600 207.400 ;
        RECT 331.800 206.200 332.400 206.800 ;
        RECT 337.200 206.200 338.000 207.000 ;
        RECT 327.000 202.200 328.200 206.200 ;
        RECT 331.600 202.200 332.400 206.200 ;
        RECT 336.000 205.600 338.000 206.200 ;
        RECT 336.000 202.200 336.800 205.600 ;
        RECT 340.400 202.200 341.200 210.600 ;
        RECT 342.000 210.200 342.600 212.400 ;
        RECT 343.800 211.600 344.400 214.600 ;
        RECT 347.600 214.200 349.200 214.400 ;
        RECT 351.800 214.200 352.400 216.400 ;
        RECT 361.400 215.400 362.200 215.600 ;
        RECT 364.400 215.400 365.200 219.800 ;
        RECT 366.000 215.600 366.800 217.200 ;
        RECT 361.400 214.800 365.200 215.400 ;
        RECT 357.400 214.200 358.200 214.400 ;
        RECT 347.600 213.600 358.600 214.200 ;
        RECT 350.600 213.400 351.400 213.600 ;
        RECT 345.200 211.600 346.000 213.200 ;
        RECT 349.000 212.400 349.800 212.600 ;
        RECT 351.600 212.400 352.400 212.600 ;
        RECT 358.000 212.400 358.600 213.600 ;
        RECT 359.600 212.800 360.400 213.000 ;
        RECT 349.000 211.800 354.000 212.400 ;
        RECT 353.200 211.600 354.000 211.800 ;
        RECT 358.000 211.600 358.800 212.400 ;
        RECT 359.600 212.200 363.400 212.800 ;
        RECT 362.600 212.000 363.400 212.200 ;
        RECT 343.200 210.800 344.400 211.600 ;
        RECT 343.800 210.200 344.400 210.800 ;
        RECT 346.800 211.000 352.400 211.200 ;
        RECT 346.800 210.800 352.600 211.000 ;
        RECT 346.800 210.600 356.600 210.800 ;
        RECT 342.000 202.200 342.800 210.200 ;
        RECT 343.800 209.600 346.000 210.200 ;
        RECT 345.200 202.200 346.000 209.600 ;
        RECT 346.800 202.200 347.600 210.600 ;
        RECT 351.800 210.200 356.600 210.600 ;
        RECT 350.000 209.000 355.400 209.600 ;
        RECT 350.000 208.800 350.800 209.000 ;
        RECT 354.600 208.800 355.400 209.000 ;
        RECT 356.000 209.000 356.600 210.200 ;
        RECT 358.000 210.400 358.600 211.600 ;
        RECT 361.000 211.400 361.800 211.600 ;
        RECT 364.400 211.400 365.200 214.800 ;
        RECT 361.000 210.800 365.200 211.400 ;
        RECT 358.000 209.800 360.400 210.400 ;
        RECT 357.400 209.000 358.200 209.200 ;
        RECT 356.000 208.400 358.200 209.000 ;
        RECT 359.800 208.800 360.400 209.800 ;
        RECT 359.800 208.000 361.200 208.800 ;
        RECT 353.400 207.400 354.200 207.600 ;
        RECT 356.200 207.400 357.000 207.600 ;
        RECT 350.000 206.200 350.800 207.000 ;
        RECT 353.400 206.800 357.000 207.400 ;
        RECT 355.600 206.200 356.200 206.800 ;
        RECT 359.600 206.200 360.400 207.000 ;
        RECT 350.000 205.600 352.000 206.200 ;
        RECT 351.200 202.200 352.000 205.600 ;
        RECT 355.600 202.200 356.400 206.200 ;
        RECT 359.800 202.200 361.000 206.200 ;
        RECT 364.400 202.200 365.200 210.800 ;
        RECT 367.600 214.300 368.400 219.800 ;
        RECT 369.200 216.000 370.000 219.800 ;
        RECT 372.400 216.000 373.200 219.800 ;
        RECT 369.200 215.800 373.200 216.000 ;
        RECT 374.000 215.800 374.800 219.800 ;
        RECT 375.600 216.000 376.400 219.800 ;
        RECT 378.800 216.000 379.600 219.800 ;
        RECT 375.600 215.800 379.600 216.000 ;
        RECT 369.400 215.400 373.000 215.800 ;
        RECT 370.000 214.400 370.800 214.800 ;
        RECT 374.000 214.400 374.600 215.800 ;
        RECT 375.800 215.400 379.400 215.800 ;
        RECT 380.400 215.600 381.200 219.800 ;
        RECT 382.000 215.800 382.800 219.800 ;
        RECT 386.400 218.400 388.000 219.800 ;
        RECT 386.400 217.600 389.200 218.400 ;
        RECT 386.400 216.200 388.000 217.600 ;
        RECT 376.400 214.400 377.200 214.800 ;
        RECT 380.400 214.400 381.000 215.600 ;
        RECT 382.000 215.200 384.600 215.800 ;
        RECT 383.800 215.000 384.600 215.200 ;
        RECT 385.200 214.800 386.800 215.600 ;
        RECT 369.200 214.300 370.800 214.400 ;
        RECT 367.600 213.800 370.800 214.300 ;
        RECT 367.600 213.700 370.000 213.800 ;
        RECT 367.600 202.200 368.400 213.700 ;
        RECT 369.200 213.600 370.000 213.700 ;
        RECT 372.200 213.600 374.800 214.400 ;
        RECT 375.600 213.800 377.200 214.400 ;
        RECT 375.600 213.600 376.400 213.800 ;
        RECT 378.600 213.600 381.200 214.400 ;
        RECT 382.000 214.200 383.600 214.400 ;
        RECT 387.400 214.200 388.000 216.200 ;
        RECT 391.600 215.800 392.400 219.800 ;
        RECT 388.600 214.800 389.400 215.600 ;
        RECT 390.000 215.200 392.400 215.800 ;
        RECT 393.200 215.600 394.000 217.200 ;
        RECT 390.000 215.000 390.800 215.200 ;
        RECT 382.000 214.000 384.200 214.200 ;
        RECT 382.000 213.600 386.400 214.000 ;
        RECT 370.800 211.600 371.600 213.200 ;
        RECT 372.200 210.200 372.800 213.600 ;
        RECT 377.200 211.600 378.000 213.200 ;
        RECT 374.000 210.200 374.800 210.400 ;
        RECT 378.600 210.200 379.200 213.600 ;
        RECT 383.600 213.400 386.400 213.600 ;
        RECT 385.600 213.200 386.400 213.400 ;
        RECT 387.000 213.600 388.000 214.200 ;
        RECT 388.800 214.400 389.400 214.800 ;
        RECT 388.800 213.600 389.600 214.400 ;
        RECT 390.800 214.300 392.400 214.400 ;
        RECT 393.200 214.300 394.000 214.400 ;
        RECT 390.800 213.700 394.000 214.300 ;
        RECT 390.800 213.600 392.400 213.700 ;
        RECT 393.200 213.600 394.000 213.700 ;
        RECT 387.000 212.400 387.600 213.600 ;
        RECT 384.200 212.200 385.000 212.400 ;
        RECT 384.200 211.600 385.800 212.200 ;
        RECT 386.800 211.600 387.600 212.400 ;
        RECT 385.000 211.400 385.800 211.600 ;
        RECT 380.400 210.200 381.200 210.400 ;
        RECT 387.000 210.200 387.600 211.600 ;
        RECT 394.800 212.300 395.600 219.800 ;
        RECT 396.400 215.800 397.200 219.800 ;
        RECT 398.000 216.000 398.800 219.800 ;
        RECT 401.200 216.000 402.000 219.800 ;
        RECT 398.000 215.800 402.000 216.000 ;
        RECT 402.800 215.800 403.600 219.800 ;
        RECT 407.200 216.200 408.800 219.800 ;
        RECT 396.600 214.400 397.200 215.800 ;
        RECT 398.200 215.400 401.800 215.800 ;
        RECT 402.800 215.200 405.200 215.800 ;
        RECT 404.400 215.000 405.200 215.200 ;
        RECT 405.800 214.800 406.600 215.600 ;
        RECT 400.400 214.400 401.200 214.800 ;
        RECT 405.800 214.400 406.400 214.800 ;
        RECT 396.400 213.600 399.000 214.400 ;
        RECT 400.400 213.800 402.000 214.400 ;
        RECT 401.200 213.600 402.000 213.800 ;
        RECT 402.800 213.600 404.400 214.400 ;
        RECT 405.600 213.600 406.400 214.400 ;
        RECT 396.400 212.300 397.200 212.400 ;
        RECT 394.800 211.700 397.200 212.300 ;
        RECT 371.800 209.600 372.800 210.200 ;
        RECT 373.400 209.600 374.800 210.200 ;
        RECT 378.200 209.600 379.200 210.200 ;
        RECT 379.800 209.600 381.200 210.200 ;
        RECT 382.000 209.600 384.600 210.200 ;
        RECT 371.800 208.400 372.600 209.600 ;
        RECT 373.400 208.400 374.000 209.600 ;
        RECT 370.800 207.600 372.600 208.400 ;
        RECT 373.200 207.600 374.000 208.400 ;
        RECT 371.800 202.200 372.600 207.600 ;
        RECT 378.200 202.200 379.000 209.600 ;
        RECT 379.800 208.400 380.400 209.600 ;
        RECT 379.600 207.600 380.400 208.400 ;
        RECT 382.000 202.200 382.800 209.600 ;
        RECT 383.800 209.400 384.600 209.600 ;
        RECT 386.400 202.200 388.000 210.200 ;
        RECT 390.000 209.600 392.400 210.200 ;
        RECT 390.000 209.400 390.800 209.600 ;
        RECT 391.600 202.200 392.400 209.600 ;
        RECT 394.800 202.200 395.600 211.700 ;
        RECT 396.400 211.600 397.200 211.700 ;
        RECT 398.400 210.400 399.000 213.600 ;
        RECT 399.600 211.600 400.400 213.200 ;
        RECT 407.200 212.800 407.800 216.200 ;
        RECT 412.400 215.800 413.200 219.800 ;
        RECT 408.400 215.400 410.000 215.600 ;
        RECT 408.400 214.800 410.400 215.400 ;
        RECT 411.000 215.200 413.200 215.800 ;
        RECT 411.000 215.000 411.800 215.200 ;
        RECT 414.000 215.000 414.800 219.800 ;
        RECT 418.400 218.400 419.200 219.800 ;
        RECT 417.200 217.800 419.200 218.400 ;
        RECT 422.800 217.800 423.600 219.800 ;
        RECT 427.000 218.400 428.200 219.800 ;
        RECT 426.800 217.800 428.200 218.400 ;
        RECT 417.200 217.000 418.000 217.800 ;
        RECT 422.800 217.200 423.400 217.800 ;
        RECT 418.800 216.400 419.600 217.200 ;
        RECT 420.600 216.600 423.400 217.200 ;
        RECT 426.800 217.000 427.600 217.800 ;
        RECT 420.600 216.400 421.400 216.600 ;
        RECT 409.800 214.400 410.400 214.800 ;
        RECT 408.400 213.400 409.200 214.200 ;
        RECT 409.800 213.800 413.200 214.400 ;
        RECT 411.600 213.600 413.200 213.800 ;
        RECT 414.800 214.200 416.400 214.400 ;
        RECT 419.000 214.200 419.600 216.400 ;
        RECT 428.600 215.400 429.400 215.600 ;
        RECT 431.600 215.400 432.400 219.800 ;
        RECT 428.600 214.800 432.400 215.400 ;
        RECT 424.600 214.200 425.400 214.400 ;
        RECT 414.800 213.600 425.800 214.200 ;
        RECT 417.800 213.400 418.600 213.600 ;
        RECT 406.800 212.400 407.800 212.800 ;
        RECT 406.000 212.200 407.800 212.400 ;
        RECT 408.600 212.800 409.200 213.400 ;
        RECT 408.600 212.200 411.200 212.800 ;
        RECT 406.000 211.600 407.400 212.200 ;
        RECT 410.400 212.000 411.200 212.200 ;
        RECT 416.200 212.400 417.000 212.600 ;
        RECT 418.800 212.400 419.600 212.600 ;
        RECT 425.200 212.400 425.800 213.600 ;
        RECT 426.800 212.800 427.600 213.000 ;
        RECT 416.200 211.800 421.200 212.400 ;
        RECT 420.400 211.600 421.200 211.800 ;
        RECT 425.200 211.600 426.000 212.400 ;
        RECT 426.800 212.200 430.600 212.800 ;
        RECT 429.800 212.000 430.600 212.200 ;
        RECT 396.400 210.200 397.200 210.400 ;
        RECT 396.400 209.600 397.800 210.200 ;
        RECT 398.400 209.600 400.400 210.400 ;
        RECT 406.800 210.200 407.400 211.600 ;
        RECT 408.200 211.400 409.000 211.600 ;
        RECT 408.200 210.800 411.600 211.400 ;
        RECT 411.000 210.200 411.600 210.800 ;
        RECT 414.000 211.000 419.600 211.200 ;
        RECT 414.000 210.800 419.800 211.000 ;
        RECT 414.000 210.600 423.800 210.800 ;
        RECT 402.800 209.600 405.200 210.200 ;
        RECT 406.800 209.600 408.800 210.200 ;
        RECT 397.200 208.400 397.800 209.600 ;
        RECT 397.200 207.600 398.000 208.400 ;
        RECT 398.600 202.200 399.400 209.600 ;
        RECT 402.800 202.200 403.600 209.600 ;
        RECT 404.400 209.400 405.200 209.600 ;
        RECT 407.200 202.200 408.800 209.600 ;
        RECT 411.000 209.600 413.200 210.200 ;
        RECT 411.000 209.400 411.800 209.600 ;
        RECT 412.400 202.200 413.200 209.600 ;
        RECT 414.000 202.200 414.800 210.600 ;
        RECT 419.000 210.200 423.800 210.600 ;
        RECT 417.200 209.000 422.600 209.600 ;
        RECT 417.200 208.800 418.000 209.000 ;
        RECT 421.800 208.800 422.600 209.000 ;
        RECT 423.200 209.000 423.800 210.200 ;
        RECT 425.200 210.400 425.800 211.600 ;
        RECT 428.200 211.400 429.000 211.600 ;
        RECT 431.600 211.400 432.400 214.800 ;
        RECT 428.200 210.800 432.400 211.400 ;
        RECT 425.200 209.800 427.600 210.400 ;
        RECT 424.600 209.000 425.400 209.200 ;
        RECT 423.200 208.400 425.400 209.000 ;
        RECT 427.000 208.800 427.600 209.800 ;
        RECT 427.000 208.000 428.400 208.800 ;
        RECT 420.600 207.400 421.400 207.600 ;
        RECT 423.400 207.400 424.200 207.600 ;
        RECT 417.200 206.200 418.000 207.000 ;
        RECT 420.600 206.800 424.200 207.400 ;
        RECT 422.800 206.200 423.400 206.800 ;
        RECT 426.800 206.200 427.600 207.000 ;
        RECT 417.200 205.600 419.200 206.200 ;
        RECT 418.400 202.200 419.200 205.600 ;
        RECT 422.800 202.200 423.600 206.200 ;
        RECT 427.000 202.200 428.200 206.200 ;
        RECT 431.600 202.200 432.400 210.800 ;
        RECT 433.200 215.800 434.000 219.800 ;
        RECT 436.400 217.800 437.200 219.800 ;
        RECT 433.200 212.400 433.800 215.800 ;
        RECT 436.400 215.600 437.000 217.800 ;
        RECT 441.200 217.600 442.000 219.800 ;
        RECT 438.000 215.600 438.800 217.200 ;
        RECT 434.600 215.000 437.000 215.600 ;
        RECT 433.200 211.600 434.000 212.400 ;
        RECT 434.600 212.000 435.200 215.000 ;
        RECT 441.200 214.400 441.800 217.600 ;
        RECT 442.800 215.600 443.600 217.200 ;
        RECT 451.800 216.400 452.600 219.800 ;
        RECT 450.800 215.800 452.600 216.400 ;
        RECT 455.600 217.600 456.400 219.800 ;
        RECT 436.200 213.600 437.200 214.400 ;
        RECT 441.200 213.600 442.000 214.400 ;
        RECT 449.200 213.600 450.000 215.200 ;
        RECT 436.000 212.800 436.800 213.600 ;
        RECT 433.200 210.200 433.800 211.600 ;
        RECT 434.600 211.400 435.400 212.000 ;
        RECT 434.600 211.200 438.800 211.400 ;
        RECT 434.800 210.800 438.800 211.200 ;
        RECT 439.600 210.800 440.400 212.400 ;
        RECT 433.200 209.600 434.600 210.200 ;
        RECT 433.800 202.200 434.600 209.600 ;
        RECT 438.000 202.200 438.800 210.800 ;
        RECT 441.200 210.200 441.800 213.600 ;
        RECT 450.800 212.300 451.600 215.800 ;
        RECT 455.600 214.400 456.200 217.600 ;
        RECT 457.200 215.600 458.000 217.200 ;
        RECT 458.800 216.000 459.600 219.800 ;
        RECT 462.000 216.000 462.800 219.800 ;
        RECT 458.800 215.800 462.800 216.000 ;
        RECT 463.600 215.800 464.400 219.800 ;
        RECT 465.800 216.400 466.600 219.800 ;
        RECT 459.000 215.400 462.600 215.800 ;
        RECT 459.600 214.400 460.400 214.800 ;
        RECT 463.600 214.400 464.200 215.800 ;
        RECT 465.200 215.600 467.600 216.400 ;
        RECT 470.000 216.000 470.800 219.800 ;
        RECT 473.200 216.000 474.000 219.800 ;
        RECT 470.000 215.800 474.000 216.000 ;
        RECT 474.800 215.800 475.600 219.800 ;
        RECT 476.400 216.000 477.200 219.800 ;
        RECT 479.600 216.000 480.400 219.800 ;
        RECT 476.400 215.800 480.400 216.000 ;
        RECT 481.200 215.800 482.000 219.800 ;
        RECT 485.400 218.400 486.200 219.800 ;
        RECT 485.400 217.600 486.800 218.400 ;
        RECT 485.400 216.400 486.200 217.600 ;
        RECT 484.400 215.800 486.200 216.400 ;
        RECT 455.600 213.600 456.400 214.400 ;
        RECT 458.800 213.800 460.400 214.400 ;
        RECT 461.800 214.300 464.400 214.400 ;
        RECT 465.200 214.300 466.000 214.400 ;
        RECT 458.800 213.600 459.600 213.800 ;
        RECT 461.800 213.700 466.000 214.300 ;
        RECT 461.800 213.600 464.400 213.700 ;
        RECT 465.200 213.600 466.000 213.700 ;
        RECT 454.000 212.300 454.800 212.400 ;
        RECT 450.800 211.700 454.800 212.300 ;
        RECT 440.200 209.400 442.000 210.200 ;
        RECT 440.200 202.200 441.000 209.400 ;
        RECT 450.800 202.200 451.600 211.700 ;
        RECT 454.000 210.800 454.800 211.700 ;
        RECT 452.400 208.800 453.200 210.400 ;
        RECT 455.600 210.200 456.200 213.600 ;
        RECT 460.400 211.600 461.200 213.200 ;
        RECT 461.800 210.200 462.400 213.600 ;
        RECT 463.600 210.200 464.400 210.400 ;
        RECT 454.600 209.400 456.400 210.200 ;
        RECT 461.400 209.600 462.400 210.200 ;
        RECT 463.000 209.600 464.400 210.200 ;
        RECT 454.600 202.200 455.400 209.400 ;
        RECT 461.400 202.200 462.200 209.600 ;
        RECT 463.000 208.400 463.600 209.600 ;
        RECT 465.200 208.800 466.000 210.400 ;
        RECT 462.800 207.600 463.600 208.400 ;
        RECT 466.800 202.200 467.600 215.600 ;
        RECT 470.200 215.400 473.800 215.800 ;
        RECT 468.400 214.300 469.200 215.200 ;
        RECT 470.800 214.400 471.600 214.800 ;
        RECT 474.800 214.400 475.400 215.800 ;
        RECT 476.600 215.400 480.200 215.800 ;
        RECT 477.200 214.400 478.000 214.800 ;
        RECT 481.200 214.400 481.800 215.800 ;
        RECT 470.000 214.300 471.600 214.400 ;
        RECT 468.400 213.800 471.600 214.300 ;
        RECT 468.400 213.700 470.800 213.800 ;
        RECT 468.400 213.600 469.200 213.700 ;
        RECT 470.000 213.600 470.800 213.700 ;
        RECT 473.000 213.600 475.600 214.400 ;
        RECT 476.400 213.800 478.000 214.400 ;
        RECT 476.400 213.600 477.200 213.800 ;
        RECT 479.400 213.600 482.000 214.400 ;
        RECT 482.800 213.600 483.600 215.200 ;
        RECT 470.000 212.300 470.800 212.400 ;
        RECT 471.600 212.300 472.400 213.200 ;
        RECT 470.000 211.700 472.400 212.300 ;
        RECT 470.000 211.600 470.800 211.700 ;
        RECT 471.600 211.600 472.400 211.700 ;
        RECT 473.000 212.300 473.600 213.600 ;
        RECT 476.400 212.300 477.200 212.400 ;
        RECT 473.000 211.700 477.200 212.300 ;
        RECT 473.000 210.200 473.600 211.700 ;
        RECT 476.400 211.600 477.200 211.700 ;
        RECT 478.000 211.600 478.800 213.200 ;
        RECT 479.400 212.300 480.000 213.600 ;
        RECT 482.800 212.300 483.600 212.400 ;
        RECT 479.400 211.700 483.600 212.300 ;
        RECT 474.800 210.200 475.600 210.400 ;
        RECT 479.400 210.200 480.000 211.700 ;
        RECT 482.800 211.600 483.600 211.700 ;
        RECT 481.200 210.200 482.000 210.400 ;
        RECT 472.600 209.600 473.600 210.200 ;
        RECT 474.200 209.600 475.600 210.200 ;
        RECT 479.000 209.600 480.000 210.200 ;
        RECT 480.600 209.600 482.000 210.200 ;
        RECT 472.600 202.200 473.400 209.600 ;
        RECT 474.200 208.400 474.800 209.600 ;
        RECT 474.000 207.600 474.800 208.400 ;
        RECT 479.000 202.200 479.800 209.600 ;
        RECT 480.600 208.400 481.200 209.600 ;
        RECT 480.400 207.600 481.200 208.400 ;
        RECT 484.400 202.200 485.200 215.800 ;
        RECT 487.600 215.600 488.400 217.200 ;
        RECT 486.000 208.800 486.800 210.400 ;
        RECT 489.200 202.200 490.000 219.800 ;
        RECT 490.800 216.000 491.600 219.800 ;
        RECT 494.000 219.200 498.000 219.800 ;
        RECT 494.000 216.000 494.800 219.200 ;
        RECT 490.800 215.800 494.800 216.000 ;
        RECT 495.600 215.800 496.400 218.600 ;
        RECT 497.200 215.800 498.000 219.200 ;
        RECT 501.400 216.400 502.200 219.800 ;
        RECT 500.400 215.800 502.200 216.400 ;
        RECT 503.600 215.800 504.400 219.800 ;
        RECT 508.000 218.400 509.600 219.800 ;
        RECT 508.000 217.600 510.800 218.400 ;
        RECT 508.000 216.200 509.600 217.600 ;
        RECT 491.000 215.400 494.600 215.800 ;
        RECT 491.600 214.400 492.400 214.800 ;
        RECT 495.800 214.400 496.400 215.800 ;
        RECT 490.800 213.800 492.400 214.400 ;
        RECT 494.000 213.800 496.400 214.400 ;
        RECT 490.800 213.600 491.600 213.800 ;
        RECT 494.000 213.600 494.800 213.800 ;
        RECT 492.400 211.600 493.200 213.200 ;
        RECT 494.000 210.200 494.600 213.600 ;
        RECT 495.600 211.600 496.400 213.200 ;
        RECT 497.200 212.800 498.000 214.400 ;
        RECT 498.800 213.600 499.600 215.200 ;
        RECT 493.400 202.200 495.400 210.200 ;
        RECT 500.400 202.200 501.200 215.800 ;
        RECT 503.600 215.200 505.800 215.800 ;
        RECT 506.800 215.400 508.400 215.600 ;
        RECT 505.000 215.000 505.800 215.200 ;
        RECT 506.400 214.800 508.400 215.400 ;
        RECT 506.400 214.400 507.000 214.800 ;
        RECT 502.000 214.300 502.800 214.400 ;
        RECT 503.600 214.300 507.000 214.400 ;
        RECT 502.000 213.800 507.000 214.300 ;
        RECT 502.000 213.700 505.200 213.800 ;
        RECT 502.000 213.600 502.800 213.700 ;
        RECT 503.600 213.600 505.200 213.700 ;
        RECT 507.600 213.400 508.400 214.200 ;
        RECT 507.600 212.800 508.200 213.400 ;
        RECT 505.600 212.200 508.200 212.800 ;
        RECT 509.000 212.800 509.600 216.200 ;
        RECT 513.200 215.800 514.000 219.800 ;
        RECT 510.200 214.800 511.000 215.600 ;
        RECT 511.600 215.200 514.000 215.800 ;
        RECT 514.800 215.800 515.600 219.800 ;
        RECT 519.200 218.400 520.800 219.800 ;
        RECT 519.200 217.600 522.000 218.400 ;
        RECT 519.200 216.200 520.800 217.600 ;
        RECT 514.800 215.200 517.200 215.800 ;
        RECT 511.600 215.000 512.400 215.200 ;
        RECT 516.400 215.000 517.200 215.200 ;
        RECT 510.400 214.400 511.000 214.800 ;
        RECT 517.800 214.800 518.600 215.600 ;
        RECT 517.800 214.400 518.400 214.800 ;
        RECT 510.400 213.600 511.200 214.400 ;
        RECT 512.400 213.600 514.000 214.400 ;
        RECT 514.800 213.600 516.400 214.400 ;
        RECT 517.600 213.600 518.400 214.400 ;
        RECT 519.200 212.800 519.800 216.200 ;
        RECT 524.400 215.800 525.200 219.800 ;
        RECT 529.000 215.800 530.600 219.800 ;
        RECT 534.600 216.400 535.400 219.800 ;
        RECT 541.400 218.400 542.200 219.800 ;
        RECT 541.400 217.600 542.800 218.400 ;
        RECT 541.400 216.400 542.200 217.600 ;
        RECT 534.600 215.800 536.400 216.400 ;
        RECT 520.400 215.400 522.000 215.600 ;
        RECT 520.400 214.800 522.400 215.400 ;
        RECT 523.000 215.200 525.200 215.800 ;
        RECT 529.200 215.600 530.000 215.800 ;
        RECT 523.000 215.000 523.800 215.200 ;
        RECT 521.800 214.400 522.400 214.800 ;
        RECT 520.400 213.400 521.200 214.200 ;
        RECT 521.800 213.800 525.200 214.400 ;
        RECT 523.600 213.600 525.200 213.800 ;
        RECT 509.000 212.400 510.000 212.800 ;
        RECT 518.800 212.400 519.800 212.800 ;
        RECT 509.000 212.200 510.800 212.400 ;
        RECT 505.600 212.000 506.400 212.200 ;
        RECT 509.400 211.600 510.800 212.200 ;
        RECT 518.000 212.200 519.800 212.400 ;
        RECT 520.600 212.800 521.200 213.400 ;
        RECT 527.600 212.800 528.400 214.400 ;
        RECT 520.600 212.200 523.200 212.800 ;
        RECT 529.400 212.400 530.000 215.600 ;
        RECT 530.800 214.300 531.600 214.400 ;
        RECT 532.400 214.300 533.200 214.400 ;
        RECT 530.800 213.700 533.200 214.300 ;
        RECT 530.800 213.600 531.600 213.700 ;
        RECT 532.400 213.600 533.200 213.700 ;
        RECT 530.800 213.200 531.400 213.600 ;
        RECT 530.600 212.400 531.400 213.200 ;
        RECT 518.000 211.600 519.400 212.200 ;
        RECT 522.400 212.000 523.200 212.200 ;
        RECT 524.400 212.300 525.200 212.400 ;
        RECT 526.000 212.300 526.800 212.400 ;
        RECT 524.400 212.200 526.800 212.300 ;
        RECT 524.400 211.700 527.600 212.200 ;
        RECT 524.400 211.600 525.200 211.700 ;
        RECT 526.000 211.600 527.600 211.700 ;
        RECT 529.200 211.600 530.000 212.400 ;
        RECT 507.800 211.400 508.600 211.600 ;
        RECT 505.200 210.800 508.600 211.400 ;
        RECT 502.000 208.800 502.800 210.400 ;
        RECT 505.200 210.200 505.800 210.800 ;
        RECT 509.400 210.200 510.000 211.600 ;
        RECT 518.800 210.200 519.400 211.600 ;
        RECT 520.200 211.400 521.000 211.600 ;
        RECT 520.200 210.800 523.600 211.400 ;
        RECT 526.800 211.200 527.600 211.600 ;
        RECT 529.400 211.400 530.000 211.600 ;
        RECT 532.400 212.300 533.200 212.400 ;
        RECT 535.600 212.300 536.400 215.800 ;
        RECT 540.400 215.800 542.200 216.400 ;
        RECT 537.200 213.600 538.000 215.200 ;
        RECT 538.800 213.600 539.600 215.200 ;
        RECT 532.400 211.700 536.400 212.300 ;
        RECT 529.400 210.800 531.400 211.400 ;
        RECT 532.400 210.800 533.200 211.700 ;
        RECT 523.000 210.200 523.600 210.800 ;
        RECT 530.800 210.200 531.400 210.800 ;
        RECT 503.600 209.600 505.800 210.200 ;
        RECT 503.600 202.200 504.400 209.600 ;
        RECT 505.000 209.400 505.800 209.600 ;
        RECT 508.000 209.600 510.000 210.200 ;
        RECT 511.600 209.600 514.000 210.200 ;
        RECT 508.000 202.200 509.600 209.600 ;
        RECT 511.600 209.400 512.400 209.600 ;
        RECT 513.200 202.200 514.000 209.600 ;
        RECT 514.800 209.600 517.200 210.200 ;
        RECT 518.800 209.600 520.800 210.200 ;
        RECT 514.800 202.200 515.600 209.600 ;
        RECT 516.400 209.400 517.200 209.600 ;
        RECT 519.200 202.200 520.800 209.600 ;
        RECT 523.000 209.600 525.200 210.200 ;
        RECT 523.000 209.400 523.800 209.600 ;
        RECT 524.400 202.200 525.200 209.600 ;
        RECT 526.000 209.600 530.000 210.200 ;
        RECT 526.000 202.200 526.800 209.600 ;
        RECT 529.200 202.800 530.000 209.600 ;
        RECT 530.800 203.400 531.600 210.200 ;
        RECT 532.400 202.800 533.200 210.200 ;
        RECT 534.000 208.800 534.800 210.400 ;
        RECT 535.600 210.300 536.400 211.700 ;
        RECT 537.200 212.300 538.000 212.400 ;
        RECT 538.900 212.300 539.500 213.600 ;
        RECT 537.200 211.700 539.500 212.300 ;
        RECT 537.200 211.600 538.000 211.700 ;
        RECT 538.800 210.300 539.600 210.400 ;
        RECT 535.600 209.700 539.600 210.300 ;
        RECT 529.200 202.200 533.200 202.800 ;
        RECT 535.600 202.200 536.400 209.700 ;
        RECT 538.800 209.600 539.600 209.700 ;
        RECT 540.400 202.200 541.200 215.800 ;
        RECT 543.600 215.000 544.400 219.800 ;
        RECT 548.000 218.400 548.800 219.800 ;
        RECT 546.800 217.800 548.800 218.400 ;
        RECT 552.400 217.800 553.200 219.800 ;
        RECT 556.600 218.400 557.800 219.800 ;
        RECT 556.400 217.800 557.800 218.400 ;
        RECT 546.800 217.000 547.600 217.800 ;
        RECT 552.400 217.200 553.000 217.800 ;
        RECT 548.400 216.400 549.200 217.200 ;
        RECT 550.200 216.600 553.000 217.200 ;
        RECT 556.400 217.000 557.200 217.800 ;
        RECT 550.200 216.400 551.000 216.600 ;
        RECT 544.400 214.200 546.000 214.400 ;
        RECT 548.600 214.200 549.200 216.400 ;
        RECT 558.200 215.400 559.000 215.600 ;
        RECT 561.200 215.400 562.000 219.800 ;
        RECT 558.200 214.800 562.000 215.400 ;
        RECT 562.800 215.000 563.600 219.800 ;
        RECT 567.200 218.400 568.000 219.800 ;
        RECT 566.000 217.800 568.000 218.400 ;
        RECT 571.600 217.800 572.400 219.800 ;
        RECT 575.800 218.400 577.000 219.800 ;
        RECT 575.600 217.800 577.000 218.400 ;
        RECT 566.000 217.000 566.800 217.800 ;
        RECT 571.600 217.200 572.200 217.800 ;
        RECT 567.600 216.400 568.400 217.200 ;
        RECT 569.400 216.600 572.200 217.200 ;
        RECT 575.600 217.000 576.400 217.800 ;
        RECT 569.400 216.400 570.200 216.600 ;
        RECT 554.200 214.200 555.000 214.400 ;
        RECT 544.400 213.600 555.400 214.200 ;
        RECT 547.400 213.400 548.200 213.600 ;
        RECT 545.800 212.400 546.600 212.600 ;
        RECT 548.400 212.400 549.200 212.600 ;
        RECT 554.800 212.400 555.400 213.600 ;
        RECT 556.400 212.800 557.200 213.000 ;
        RECT 545.800 211.800 550.800 212.400 ;
        RECT 550.000 211.600 550.800 211.800 ;
        RECT 554.800 211.600 555.600 212.400 ;
        RECT 556.400 212.200 560.200 212.800 ;
        RECT 559.400 212.000 560.200 212.200 ;
        RECT 543.600 211.000 549.200 211.200 ;
        RECT 543.600 210.800 549.400 211.000 ;
        RECT 543.600 210.600 553.400 210.800 ;
        RECT 542.000 208.800 542.800 210.400 ;
        RECT 543.600 202.200 544.400 210.600 ;
        RECT 548.600 210.200 553.400 210.600 ;
        RECT 546.800 209.000 552.200 209.600 ;
        RECT 546.800 208.800 547.600 209.000 ;
        RECT 551.400 208.800 552.200 209.000 ;
        RECT 552.800 209.000 553.400 210.200 ;
        RECT 554.800 210.400 555.400 211.600 ;
        RECT 557.800 211.400 558.600 211.600 ;
        RECT 561.200 211.400 562.000 214.800 ;
        RECT 567.800 214.400 568.400 216.400 ;
        RECT 577.400 215.400 578.200 215.600 ;
        RECT 580.400 215.400 581.200 219.800 ;
        RECT 577.400 214.800 581.200 215.400 ;
        RECT 563.600 214.200 565.200 214.400 ;
        RECT 567.600 214.200 568.400 214.400 ;
        RECT 573.400 214.200 574.200 214.400 ;
        RECT 563.600 213.600 574.600 214.200 ;
        RECT 566.600 213.400 567.400 213.600 ;
        RECT 565.000 212.400 565.800 212.600 ;
        RECT 565.000 211.800 570.000 212.400 ;
        RECT 569.200 211.600 570.000 211.800 ;
        RECT 557.800 210.800 562.000 211.400 ;
        RECT 554.800 209.800 557.200 210.400 ;
        RECT 554.200 209.000 555.000 209.200 ;
        RECT 552.800 208.400 555.000 209.000 ;
        RECT 556.600 208.800 557.200 209.800 ;
        RECT 556.600 208.000 558.000 208.800 ;
        RECT 550.200 207.400 551.000 207.600 ;
        RECT 553.000 207.400 553.800 207.600 ;
        RECT 546.800 206.200 547.600 207.000 ;
        RECT 550.200 206.800 553.800 207.400 ;
        RECT 552.400 206.200 553.000 206.800 ;
        RECT 556.400 206.200 557.200 207.000 ;
        RECT 546.800 205.600 548.800 206.200 ;
        RECT 548.000 202.200 548.800 205.600 ;
        RECT 552.400 202.200 553.200 206.200 ;
        RECT 556.600 202.200 557.800 206.200 ;
        RECT 561.200 202.200 562.000 210.800 ;
        RECT 562.800 211.000 568.400 211.200 ;
        RECT 562.800 210.800 568.600 211.000 ;
        RECT 562.800 210.600 572.600 210.800 ;
        RECT 562.800 202.200 563.600 210.600 ;
        RECT 567.800 210.200 572.600 210.600 ;
        RECT 566.000 209.000 571.400 209.600 ;
        RECT 566.000 208.800 566.800 209.000 ;
        RECT 570.600 208.800 571.400 209.000 ;
        RECT 572.000 209.000 572.600 210.200 ;
        RECT 574.000 210.400 574.600 213.600 ;
        RECT 575.600 212.800 576.400 213.000 ;
        RECT 575.600 212.200 579.400 212.800 ;
        RECT 578.600 212.000 579.400 212.200 ;
        RECT 577.000 211.400 577.800 211.600 ;
        RECT 580.400 211.400 581.200 214.800 ;
        RECT 582.000 215.200 582.800 219.800 ;
        RECT 582.000 214.600 584.200 215.200 ;
        RECT 582.000 211.600 582.800 213.200 ;
        RECT 583.600 211.600 584.200 214.600 ;
        RECT 577.000 210.800 581.200 211.400 ;
        RECT 574.000 209.800 576.400 210.400 ;
        RECT 573.400 209.000 574.200 209.200 ;
        RECT 572.000 208.400 574.200 209.000 ;
        RECT 575.800 208.800 576.400 209.800 ;
        RECT 575.800 208.000 577.200 208.800 ;
        RECT 569.400 207.400 570.200 207.600 ;
        RECT 572.200 207.400 573.000 207.600 ;
        RECT 566.000 206.200 566.800 207.000 ;
        RECT 569.400 206.800 573.000 207.400 ;
        RECT 571.600 206.200 572.200 206.800 ;
        RECT 575.600 206.200 576.400 207.000 ;
        RECT 566.000 205.600 568.000 206.200 ;
        RECT 567.200 202.200 568.000 205.600 ;
        RECT 571.600 202.200 572.400 206.200 ;
        RECT 575.800 202.200 577.000 206.200 ;
        RECT 580.400 202.200 581.200 210.800 ;
        RECT 583.600 210.800 584.800 211.600 ;
        RECT 583.600 210.200 584.200 210.800 ;
        RECT 582.000 209.600 584.200 210.200 ;
        RECT 582.000 202.200 582.800 209.600 ;
        RECT 1.200 191.400 2.000 199.800 ;
        RECT 5.600 196.400 6.400 199.800 ;
        RECT 4.400 195.800 6.400 196.400 ;
        RECT 10.000 195.800 10.800 199.800 ;
        RECT 14.200 195.800 15.400 199.800 ;
        RECT 4.400 195.000 5.200 195.800 ;
        RECT 10.000 195.200 10.600 195.800 ;
        RECT 7.800 194.600 11.400 195.200 ;
        RECT 14.000 195.000 14.800 195.800 ;
        RECT 7.800 194.400 8.600 194.600 ;
        RECT 10.600 194.400 11.400 194.600 ;
        RECT 4.400 193.000 5.200 193.200 ;
        RECT 9.000 193.000 9.800 193.200 ;
        RECT 4.400 192.400 9.800 193.000 ;
        RECT 10.400 193.000 12.600 193.600 ;
        RECT 10.400 191.800 11.000 193.000 ;
        RECT 11.800 192.800 12.600 193.000 ;
        RECT 14.200 193.200 15.600 194.000 ;
        RECT 14.200 192.200 14.800 193.200 ;
        RECT 6.200 191.400 11.000 191.800 ;
        RECT 1.200 191.200 11.000 191.400 ;
        RECT 12.400 191.600 14.800 192.200 ;
        RECT 1.200 191.000 7.000 191.200 ;
        RECT 1.200 190.800 6.800 191.000 ;
        RECT 12.400 190.400 13.000 191.600 ;
        RECT 18.800 191.200 19.600 199.800 ;
        RECT 15.400 190.600 19.600 191.200 ;
        RECT 20.400 191.400 21.200 199.800 ;
        RECT 24.800 196.400 25.600 199.800 ;
        RECT 23.600 195.800 25.600 196.400 ;
        RECT 29.200 195.800 30.000 199.800 ;
        RECT 33.400 195.800 34.600 199.800 ;
        RECT 23.600 195.000 24.400 195.800 ;
        RECT 29.200 195.200 29.800 195.800 ;
        RECT 27.000 194.600 30.600 195.200 ;
        RECT 33.200 195.000 34.000 195.800 ;
        RECT 27.000 194.400 27.800 194.600 ;
        RECT 29.800 194.400 30.600 194.600 ;
        RECT 23.600 193.000 24.400 193.200 ;
        RECT 28.200 193.000 29.000 193.200 ;
        RECT 23.600 192.400 29.000 193.000 ;
        RECT 29.600 193.000 31.800 193.600 ;
        RECT 29.600 191.800 30.200 193.000 ;
        RECT 31.000 192.800 31.800 193.000 ;
        RECT 33.400 193.200 34.800 194.000 ;
        RECT 33.400 192.200 34.000 193.200 ;
        RECT 25.400 191.400 30.200 191.800 ;
        RECT 20.400 191.200 30.200 191.400 ;
        RECT 31.600 191.600 34.000 192.200 ;
        RECT 20.400 191.000 26.200 191.200 ;
        RECT 20.400 190.800 26.000 191.000 ;
        RECT 15.400 190.400 16.200 190.600 ;
        RECT 7.600 190.300 8.400 190.400 ;
        RECT 9.200 190.300 10.000 190.400 ;
        RECT 7.600 190.200 10.000 190.300 ;
        RECT 3.400 189.700 10.000 190.200 ;
        RECT 3.400 189.600 8.400 189.700 ;
        RECT 9.200 189.600 10.000 189.700 ;
        RECT 12.400 189.600 13.200 190.400 ;
        RECT 17.000 189.800 17.800 190.000 ;
        RECT 3.400 189.400 4.200 189.600 ;
        RECT 5.000 188.400 5.800 188.600 ;
        RECT 12.400 188.400 13.000 189.600 ;
        RECT 14.000 189.200 17.800 189.800 ;
        RECT 14.000 189.000 14.800 189.200 ;
        RECT 2.000 187.800 13.000 188.400 ;
        RECT 2.000 187.600 3.600 187.800 ;
        RECT 1.200 182.200 2.000 187.000 ;
        RECT 6.200 185.600 6.800 187.800 ;
        RECT 11.800 187.600 12.600 187.800 ;
        RECT 18.800 187.200 19.600 190.600 ;
        RECT 31.600 190.400 32.200 191.600 ;
        RECT 38.000 191.200 38.800 199.800 ;
        RECT 39.600 191.600 40.400 193.200 ;
        RECT 34.600 190.600 38.800 191.200 ;
        RECT 34.600 190.400 35.400 190.600 ;
        RECT 26.800 190.200 27.600 190.400 ;
        RECT 22.600 189.600 27.600 190.200 ;
        RECT 31.600 189.600 32.400 190.400 ;
        RECT 36.200 189.800 37.000 190.000 ;
        RECT 22.600 189.400 23.400 189.600 ;
        RECT 25.200 189.400 26.000 189.600 ;
        RECT 24.200 188.400 25.000 188.600 ;
        RECT 31.600 188.400 32.200 189.600 ;
        RECT 33.200 189.200 37.000 189.800 ;
        RECT 33.200 189.000 34.000 189.200 ;
        RECT 21.200 187.800 32.200 188.400 ;
        RECT 21.200 187.600 22.800 187.800 ;
        RECT 15.800 186.600 19.600 187.200 ;
        RECT 15.800 186.400 16.600 186.600 ;
        RECT 4.400 184.200 5.200 185.000 ;
        RECT 6.000 184.800 6.800 185.600 ;
        RECT 7.800 185.400 8.600 185.600 ;
        RECT 7.800 184.800 10.600 185.400 ;
        RECT 10.000 184.200 10.600 184.800 ;
        RECT 14.000 184.200 14.800 185.000 ;
        RECT 4.400 183.600 6.400 184.200 ;
        RECT 5.600 182.200 6.400 183.600 ;
        RECT 10.000 182.200 10.800 184.200 ;
        RECT 14.000 183.600 15.400 184.200 ;
        RECT 14.200 182.200 15.400 183.600 ;
        RECT 18.800 182.200 19.600 186.600 ;
        RECT 20.400 182.200 21.200 187.000 ;
        RECT 25.400 185.600 26.000 187.800 ;
        RECT 31.000 187.600 31.800 187.800 ;
        RECT 38.000 187.200 38.800 190.600 ;
        RECT 35.000 186.600 38.800 187.200 ;
        RECT 35.000 186.400 35.800 186.600 ;
        RECT 23.600 184.200 24.400 185.000 ;
        RECT 25.200 184.800 26.000 185.600 ;
        RECT 27.000 185.400 27.800 185.600 ;
        RECT 27.000 184.800 29.800 185.400 ;
        RECT 29.200 184.200 29.800 184.800 ;
        RECT 33.200 184.200 34.000 185.000 ;
        RECT 23.600 183.600 25.600 184.200 ;
        RECT 24.800 182.200 25.600 183.600 ;
        RECT 29.200 182.200 30.000 184.200 ;
        RECT 33.200 183.600 34.600 184.200 ;
        RECT 33.400 182.200 34.600 183.600 ;
        RECT 38.000 182.200 38.800 186.600 ;
        RECT 41.200 186.200 42.000 199.800 ;
        RECT 44.400 191.200 45.200 199.800 ;
        RECT 48.600 192.400 49.400 199.800 ;
        RECT 53.400 192.600 54.200 199.800 ;
        RECT 48.600 191.800 50.000 192.400 ;
        RECT 52.400 191.800 54.200 192.600 ;
        RECT 49.200 191.600 50.000 191.800 ;
        RECT 44.400 190.800 48.400 191.200 ;
        RECT 44.400 190.600 48.600 190.800 ;
        RECT 47.800 190.000 48.600 190.600 ;
        RECT 49.400 190.400 50.000 191.600 ;
        RECT 46.400 188.400 47.200 189.200 ;
        RECT 42.800 186.800 43.600 188.400 ;
        RECT 46.000 187.600 47.000 188.400 ;
        RECT 48.000 187.000 48.600 190.000 ;
        RECT 49.200 189.600 50.000 190.400 ;
        RECT 46.200 186.400 48.600 187.000 ;
        RECT 40.200 185.600 42.000 186.200 ;
        RECT 40.200 184.400 41.000 185.600 ;
        RECT 44.400 184.800 45.200 186.400 ;
        RECT 39.600 183.600 41.000 184.400 ;
        RECT 46.200 184.200 46.800 186.400 ;
        RECT 49.400 186.200 50.000 189.600 ;
        RECT 52.600 188.400 53.200 191.800 ;
        RECT 55.600 191.600 56.400 193.200 ;
        RECT 54.000 189.600 54.800 191.200 ;
        RECT 52.400 187.600 53.200 188.400 ;
        RECT 40.200 182.200 41.000 183.600 ;
        RECT 46.000 182.200 46.800 184.200 ;
        RECT 49.200 182.200 50.000 186.200 ;
        RECT 50.800 184.800 51.600 186.400 ;
        RECT 52.600 184.400 53.200 187.600 ;
        RECT 57.200 186.200 58.000 199.800 ;
        RECT 60.400 191.600 61.200 193.200 ;
        RECT 58.800 188.300 59.600 188.400 ;
        RECT 62.000 188.300 62.800 199.800 ;
        RECT 66.000 193.600 66.800 194.400 ;
        RECT 66.000 192.400 66.600 193.600 ;
        RECT 67.400 192.400 68.200 199.800 ;
        RECT 73.200 195.800 74.000 199.800 ;
        RECT 65.200 191.800 66.600 192.400 ;
        RECT 67.200 191.800 68.200 192.400 ;
        RECT 65.200 191.600 66.000 191.800 ;
        RECT 63.600 190.300 64.400 190.400 ;
        RECT 67.200 190.300 67.800 191.800 ;
        RECT 73.400 191.600 74.000 195.800 ;
        RECT 76.400 191.800 77.200 199.800 ;
        RECT 73.400 191.000 75.800 191.600 ;
        RECT 63.600 189.700 67.800 190.300 ;
        RECT 63.600 189.600 64.400 189.700 ;
        RECT 67.200 188.400 67.800 189.700 ;
        RECT 68.400 188.800 69.200 190.400 ;
        RECT 73.200 189.600 74.000 190.400 ;
        RECT 58.800 187.700 62.800 188.300 ;
        RECT 58.800 186.800 59.600 187.700 ;
        RECT 62.000 186.200 62.800 187.700 ;
        RECT 63.600 186.800 64.400 188.400 ;
        RECT 65.200 187.600 67.800 188.400 ;
        RECT 70.000 188.200 70.800 188.400 ;
        RECT 69.200 187.600 70.800 188.200 ;
        RECT 71.600 187.600 72.400 189.200 ;
        RECT 73.400 188.800 74.000 189.600 ;
        RECT 73.200 188.000 74.400 188.800 ;
        RECT 75.200 187.600 75.800 191.000 ;
        RECT 76.600 190.400 77.200 191.800 ;
        RECT 78.000 192.300 78.800 192.400 ;
        RECT 79.600 192.300 80.400 199.800 ;
        RECT 81.200 192.300 82.000 193.200 ;
        RECT 78.000 191.700 82.000 192.300 ;
        RECT 78.000 191.600 78.800 191.700 ;
        RECT 76.400 189.600 77.200 190.400 ;
        RECT 65.400 186.200 66.000 187.600 ;
        RECT 69.200 187.200 70.000 187.600 ;
        RECT 75.200 187.400 76.000 187.600 ;
        RECT 73.000 187.000 76.000 187.400 ;
        RECT 71.800 186.800 76.000 187.000 ;
        RECT 67.000 186.200 70.600 186.600 ;
        RECT 71.800 186.400 73.600 186.800 ;
        RECT 71.800 186.200 72.400 186.400 ;
        RECT 76.600 186.200 77.200 189.600 ;
        RECT 52.400 182.200 53.200 184.400 ;
        RECT 56.200 185.600 58.000 186.200 ;
        RECT 61.000 185.600 62.800 186.200 ;
        RECT 56.200 184.400 57.000 185.600 ;
        RECT 61.000 184.400 61.800 185.600 ;
        RECT 56.200 183.600 58.000 184.400 ;
        RECT 61.000 183.600 62.800 184.400 ;
        RECT 56.200 182.200 57.000 183.600 ;
        RECT 61.000 182.200 61.800 183.600 ;
        RECT 65.200 182.200 66.000 186.200 ;
        RECT 66.800 186.000 70.800 186.200 ;
        RECT 66.800 182.200 67.600 186.000 ;
        RECT 70.000 182.200 70.800 186.000 ;
        RECT 71.600 182.200 72.400 186.200 ;
        RECT 75.800 185.200 77.200 186.200 ;
        RECT 75.800 184.400 76.600 185.200 ;
        RECT 78.000 184.800 78.800 186.400 ;
        RECT 75.800 183.600 77.200 184.400 ;
        RECT 75.800 182.200 76.600 183.600 ;
        RECT 79.600 182.200 80.400 191.700 ;
        RECT 81.200 191.600 82.000 191.700 ;
        RECT 82.800 186.200 83.600 199.800 ;
        RECT 84.400 188.300 85.200 188.400 ;
        RECT 86.000 188.300 86.800 199.800 ;
        RECT 87.600 192.300 88.400 192.400 ;
        RECT 89.200 192.300 90.000 193.200 ;
        RECT 87.600 191.700 90.000 192.300 ;
        RECT 87.600 191.600 88.400 191.700 ;
        RECT 89.200 191.600 90.000 191.700 ;
        RECT 84.400 187.700 86.800 188.300 ;
        RECT 84.400 186.800 85.200 187.700 ;
        RECT 81.800 185.600 83.600 186.200 ;
        RECT 81.800 184.400 82.600 185.600 ;
        RECT 81.200 183.600 82.600 184.400 ;
        RECT 81.800 182.200 82.600 183.600 ;
        RECT 86.000 182.200 86.800 187.700 ;
        RECT 90.800 190.300 91.600 199.800 ;
        RECT 94.000 190.300 94.800 190.400 ;
        RECT 90.800 189.700 94.800 190.300 ;
        RECT 87.600 184.800 88.400 186.400 ;
        RECT 90.800 186.200 91.600 189.700 ;
        RECT 94.000 189.600 94.800 189.700 ;
        RECT 95.600 190.300 96.400 199.800 ;
        RECT 99.800 192.400 100.600 199.800 ;
        RECT 101.200 193.600 102.000 194.400 ;
        RECT 101.400 192.400 102.000 193.600 ;
        RECT 104.400 193.600 105.200 194.400 ;
        RECT 104.400 192.400 105.000 193.600 ;
        RECT 105.800 192.400 106.600 199.800 ;
        RECT 99.800 191.800 100.800 192.400 ;
        RECT 101.400 191.800 102.800 192.400 ;
        RECT 98.800 190.300 99.600 190.400 ;
        RECT 95.600 189.700 99.600 190.300 ;
        RECT 92.400 186.800 93.200 188.400 ;
        RECT 89.800 185.600 91.600 186.200 ;
        RECT 89.800 182.200 90.600 185.600 ;
        RECT 94.000 184.800 94.800 186.400 ;
        RECT 95.600 182.200 96.400 189.700 ;
        RECT 98.800 188.800 99.600 189.700 ;
        RECT 100.200 188.400 100.800 191.800 ;
        RECT 102.000 191.600 102.800 191.800 ;
        RECT 103.600 191.800 105.000 192.400 ;
        RECT 105.600 191.800 106.600 192.400 ;
        RECT 103.600 191.600 104.400 191.800 ;
        RECT 102.100 190.300 102.700 191.600 ;
        RECT 105.600 190.300 106.200 191.800 ;
        RECT 110.000 191.600 110.800 193.200 ;
        RECT 102.100 189.700 106.200 190.300 ;
        RECT 105.600 188.400 106.200 189.700 ;
        RECT 106.800 190.300 107.600 190.400 ;
        RECT 110.100 190.300 110.700 191.600 ;
        RECT 106.800 189.700 110.700 190.300 ;
        RECT 106.800 188.800 107.600 189.700 ;
        RECT 97.200 188.200 98.000 188.400 ;
        RECT 97.200 187.600 98.800 188.200 ;
        RECT 100.200 187.600 102.800 188.400 ;
        RECT 103.600 187.600 106.200 188.400 ;
        RECT 108.400 188.200 109.200 188.400 ;
        RECT 107.600 187.600 109.200 188.200 ;
        RECT 98.000 187.200 98.800 187.600 ;
        RECT 97.400 186.200 101.000 186.600 ;
        RECT 102.000 186.200 102.600 187.600 ;
        RECT 103.800 186.200 104.400 187.600 ;
        RECT 107.600 187.200 108.400 187.600 ;
        RECT 105.400 186.200 109.000 186.600 ;
        RECT 111.600 186.200 112.400 199.800 ;
        RECT 116.400 192.300 117.200 199.800 ;
        RECT 118.000 192.300 118.800 193.200 ;
        RECT 116.400 191.700 118.800 192.300 ;
        RECT 113.200 188.300 114.000 188.400 ;
        RECT 113.200 187.700 115.500 188.300 ;
        RECT 113.200 186.800 114.000 187.700 ;
        RECT 114.900 186.400 115.500 187.700 ;
        RECT 97.200 186.000 101.200 186.200 ;
        RECT 97.200 182.200 98.000 186.000 ;
        RECT 100.400 182.200 101.200 186.000 ;
        RECT 102.000 182.200 102.800 186.200 ;
        RECT 103.600 182.200 104.400 186.200 ;
        RECT 105.200 186.000 109.200 186.200 ;
        RECT 105.200 182.200 106.000 186.000 ;
        RECT 108.400 182.200 109.200 186.000 ;
        RECT 110.600 185.600 112.400 186.200 ;
        RECT 110.600 184.400 111.400 185.600 ;
        RECT 114.800 184.800 115.600 186.400 ;
        RECT 110.600 183.600 112.400 184.400 ;
        RECT 110.600 182.200 111.400 183.600 ;
        RECT 116.400 182.200 117.200 191.700 ;
        RECT 118.000 191.600 118.800 191.700 ;
        RECT 119.600 186.200 120.400 199.800 ;
        RECT 122.800 191.400 123.600 199.800 ;
        RECT 127.200 196.400 128.000 199.800 ;
        RECT 126.000 195.800 128.000 196.400 ;
        RECT 131.600 195.800 132.400 199.800 ;
        RECT 135.800 195.800 137.000 199.800 ;
        RECT 126.000 195.000 126.800 195.800 ;
        RECT 131.600 195.200 132.200 195.800 ;
        RECT 129.400 194.600 133.000 195.200 ;
        RECT 135.600 195.000 136.400 195.800 ;
        RECT 129.400 194.400 130.200 194.600 ;
        RECT 132.200 194.400 133.000 194.600 ;
        RECT 126.000 193.000 126.800 193.200 ;
        RECT 130.600 193.000 131.400 193.200 ;
        RECT 126.000 192.400 131.400 193.000 ;
        RECT 132.000 193.000 134.200 193.600 ;
        RECT 132.000 191.800 132.600 193.000 ;
        RECT 133.400 192.800 134.200 193.000 ;
        RECT 135.800 193.200 137.200 194.000 ;
        RECT 135.800 192.200 136.400 193.200 ;
        RECT 127.800 191.400 132.600 191.800 ;
        RECT 122.800 191.200 132.600 191.400 ;
        RECT 134.000 191.600 136.400 192.200 ;
        RECT 122.800 191.000 128.600 191.200 ;
        RECT 122.800 190.800 128.400 191.000 ;
        RECT 129.200 190.200 130.000 190.400 ;
        RECT 125.000 189.600 130.000 190.200 ;
        RECT 125.000 189.400 125.800 189.600 ;
        RECT 126.600 188.400 127.400 188.600 ;
        RECT 134.000 188.400 134.600 191.600 ;
        RECT 140.400 191.200 141.200 199.800 ;
        RECT 137.000 190.600 141.200 191.200 ;
        RECT 146.800 191.400 147.600 199.800 ;
        RECT 151.200 196.400 152.000 199.800 ;
        RECT 150.000 195.800 152.000 196.400 ;
        RECT 155.600 195.800 156.400 199.800 ;
        RECT 159.800 195.800 161.000 199.800 ;
        RECT 150.000 195.000 150.800 195.800 ;
        RECT 155.600 195.200 156.200 195.800 ;
        RECT 153.400 194.600 157.000 195.200 ;
        RECT 159.600 195.000 160.400 195.800 ;
        RECT 153.400 194.400 154.200 194.600 ;
        RECT 156.200 194.400 157.000 194.600 ;
        RECT 150.000 193.000 150.800 193.200 ;
        RECT 154.600 193.000 155.400 193.200 ;
        RECT 150.000 192.400 155.400 193.000 ;
        RECT 156.000 193.000 158.200 193.600 ;
        RECT 156.000 191.800 156.600 193.000 ;
        RECT 157.400 192.800 158.200 193.000 ;
        RECT 159.800 193.200 161.200 194.000 ;
        RECT 159.800 192.200 160.400 193.200 ;
        RECT 151.800 191.400 156.600 191.800 ;
        RECT 146.800 191.200 156.600 191.400 ;
        RECT 158.000 191.600 160.400 192.200 ;
        RECT 146.800 191.000 152.600 191.200 ;
        RECT 146.800 190.800 152.400 191.000 ;
        RECT 137.000 190.400 137.800 190.600 ;
        RECT 138.600 189.800 139.400 190.000 ;
        RECT 135.600 189.200 139.400 189.800 ;
        RECT 135.600 189.000 136.400 189.200 ;
        RECT 121.200 186.800 122.000 188.400 ;
        RECT 123.600 187.800 134.600 188.400 ;
        RECT 123.600 187.600 125.200 187.800 ;
        RECT 127.600 187.600 128.400 187.800 ;
        RECT 133.400 187.600 134.200 187.800 ;
        RECT 118.600 185.600 120.400 186.200 ;
        RECT 118.600 184.400 119.400 185.600 ;
        RECT 118.600 183.600 120.400 184.400 ;
        RECT 118.600 182.200 119.400 183.600 ;
        RECT 122.800 182.200 123.600 187.000 ;
        RECT 127.800 185.600 128.400 187.600 ;
        RECT 140.400 187.200 141.200 190.600 ;
        RECT 153.200 190.200 154.000 190.400 ;
        RECT 149.000 189.600 154.000 190.200 ;
        RECT 156.400 190.300 157.200 190.400 ;
        RECT 158.000 190.300 158.600 191.600 ;
        RECT 164.400 191.200 165.200 199.800 ;
        RECT 161.000 190.600 165.200 191.200 ;
        RECT 166.000 191.400 166.800 199.800 ;
        RECT 170.400 196.400 171.200 199.800 ;
        RECT 169.200 195.800 171.200 196.400 ;
        RECT 174.800 195.800 175.600 199.800 ;
        RECT 179.000 195.800 180.200 199.800 ;
        RECT 169.200 195.000 170.000 195.800 ;
        RECT 174.800 195.200 175.400 195.800 ;
        RECT 172.600 194.600 176.200 195.200 ;
        RECT 178.800 195.000 179.600 195.800 ;
        RECT 172.600 194.400 173.400 194.600 ;
        RECT 175.400 194.400 176.200 194.600 ;
        RECT 169.200 193.000 170.000 193.200 ;
        RECT 173.800 193.000 174.600 193.200 ;
        RECT 169.200 192.400 174.600 193.000 ;
        RECT 175.200 193.000 177.400 193.600 ;
        RECT 175.200 191.800 175.800 193.000 ;
        RECT 176.600 192.800 177.400 193.000 ;
        RECT 179.000 193.200 180.400 194.000 ;
        RECT 179.000 192.200 179.600 193.200 ;
        RECT 171.000 191.400 175.800 191.800 ;
        RECT 166.000 191.200 175.800 191.400 ;
        RECT 177.200 191.600 179.600 192.200 ;
        RECT 166.000 191.000 171.800 191.200 ;
        RECT 166.000 190.800 171.600 191.000 ;
        RECT 161.000 190.400 161.800 190.600 ;
        RECT 156.400 189.700 158.700 190.300 ;
        RECT 162.600 189.800 163.400 190.000 ;
        RECT 156.400 189.600 157.200 189.700 ;
        RECT 149.000 189.400 149.800 189.600 ;
        RECT 151.600 189.400 152.400 189.600 ;
        RECT 150.600 188.400 151.400 188.600 ;
        RECT 158.000 188.400 158.600 189.700 ;
        RECT 159.600 189.200 163.400 189.800 ;
        RECT 159.600 189.000 160.400 189.200 ;
        RECT 147.600 187.800 158.600 188.400 ;
        RECT 147.600 187.600 149.200 187.800 ;
        RECT 137.400 186.600 141.200 187.200 ;
        RECT 137.400 186.400 138.200 186.600 ;
        RECT 126.000 184.200 126.800 185.000 ;
        RECT 127.600 184.800 128.400 185.600 ;
        RECT 129.400 185.400 130.200 185.600 ;
        RECT 129.400 184.800 132.200 185.400 ;
        RECT 131.600 184.200 132.200 184.800 ;
        RECT 135.600 184.200 136.400 185.000 ;
        RECT 140.400 184.300 141.200 186.600 ;
        RECT 145.200 184.300 146.000 184.400 ;
        RECT 126.000 183.600 128.000 184.200 ;
        RECT 127.200 182.200 128.000 183.600 ;
        RECT 131.600 182.200 132.400 184.200 ;
        RECT 135.600 183.600 137.000 184.200 ;
        RECT 135.800 182.200 137.000 183.600 ;
        RECT 140.400 183.700 146.000 184.300 ;
        RECT 140.400 182.200 141.200 183.700 ;
        RECT 145.200 183.600 146.000 183.700 ;
        RECT 146.800 182.200 147.600 187.000 ;
        RECT 151.800 185.600 152.400 187.800 ;
        RECT 157.400 187.600 158.200 187.800 ;
        RECT 164.400 187.200 165.200 190.600 ;
        RECT 172.400 190.300 173.200 190.400 ;
        RECT 175.600 190.300 176.400 190.400 ;
        RECT 172.400 190.200 176.400 190.300 ;
        RECT 168.200 189.700 176.400 190.200 ;
        RECT 168.200 189.600 173.200 189.700 ;
        RECT 175.600 189.600 176.400 189.700 ;
        RECT 168.200 189.400 169.000 189.600 ;
        RECT 169.800 188.400 170.600 188.600 ;
        RECT 177.200 188.400 177.800 191.600 ;
        RECT 183.600 191.200 184.400 199.800 ;
        RECT 180.200 190.600 184.400 191.200 ;
        RECT 180.200 190.400 181.000 190.600 ;
        RECT 181.800 189.800 182.600 190.000 ;
        RECT 178.800 189.200 182.600 189.800 ;
        RECT 178.800 189.000 179.600 189.200 ;
        RECT 166.800 187.800 177.800 188.400 ;
        RECT 166.800 187.600 168.400 187.800 ;
        RECT 170.800 187.600 171.600 187.800 ;
        RECT 176.600 187.600 177.400 187.800 ;
        RECT 161.400 186.600 165.200 187.200 ;
        RECT 161.400 186.400 162.200 186.600 ;
        RECT 150.000 184.200 150.800 185.000 ;
        RECT 151.600 184.800 152.400 185.600 ;
        RECT 153.400 185.400 154.200 185.600 ;
        RECT 153.400 184.800 156.200 185.400 ;
        RECT 155.600 184.200 156.200 184.800 ;
        RECT 159.600 184.200 160.400 185.000 ;
        RECT 150.000 183.600 152.000 184.200 ;
        RECT 151.200 182.200 152.000 183.600 ;
        RECT 155.600 182.200 156.400 184.200 ;
        RECT 159.600 183.600 161.000 184.200 ;
        RECT 159.800 182.200 161.000 183.600 ;
        RECT 164.400 182.200 165.200 186.600 ;
        RECT 166.000 182.200 166.800 187.000 ;
        RECT 171.000 185.600 171.600 187.600 ;
        RECT 183.600 187.200 184.400 190.600 ;
        RECT 180.600 186.600 184.400 187.200 ;
        RECT 180.600 186.400 181.400 186.600 ;
        RECT 169.200 184.200 170.000 185.000 ;
        RECT 170.800 184.800 171.600 185.600 ;
        RECT 172.600 185.400 173.400 185.600 ;
        RECT 172.600 184.800 175.400 185.400 ;
        RECT 174.800 184.200 175.400 184.800 ;
        RECT 178.800 184.200 179.600 185.000 ;
        RECT 169.200 183.600 171.200 184.200 ;
        RECT 170.400 182.200 171.200 183.600 ;
        RECT 174.800 182.200 175.600 184.200 ;
        RECT 178.800 183.600 180.200 184.200 ;
        RECT 179.000 182.200 180.200 183.600 ;
        RECT 183.600 182.200 184.400 186.600 ;
        RECT 185.200 184.800 186.000 186.400 ;
        RECT 186.800 182.200 187.600 199.800 ;
        RECT 189.200 193.600 190.000 194.400 ;
        RECT 189.200 192.400 189.800 193.600 ;
        RECT 190.600 192.400 191.400 199.800 ;
        RECT 188.400 191.800 189.800 192.400 ;
        RECT 188.400 191.600 189.200 191.800 ;
        RECT 190.400 191.600 192.400 192.400 ;
        RECT 194.800 191.600 195.600 193.200 ;
        RECT 190.400 188.400 191.000 191.600 ;
        RECT 191.600 190.300 192.400 190.400 ;
        RECT 194.900 190.300 195.500 191.600 ;
        RECT 191.600 189.700 195.500 190.300 ;
        RECT 191.600 188.800 192.400 189.700 ;
        RECT 188.400 187.600 191.000 188.400 ;
        RECT 193.200 188.200 194.000 188.400 ;
        RECT 192.400 187.600 194.000 188.200 ;
        RECT 188.600 186.200 189.200 187.600 ;
        RECT 192.400 187.200 193.200 187.600 ;
        RECT 190.200 186.200 193.800 186.600 ;
        RECT 196.400 186.200 197.200 199.800 ;
        RECT 201.800 194.400 202.600 199.800 ;
        RECT 200.400 193.600 201.200 194.400 ;
        RECT 201.800 193.600 203.600 194.400 ;
        RECT 200.400 192.400 201.000 193.600 ;
        RECT 201.800 192.400 202.600 193.600 ;
        RECT 199.600 191.800 201.000 192.400 ;
        RECT 201.600 191.800 202.600 192.400 ;
        RECT 199.600 191.600 200.400 191.800 ;
        RECT 201.600 188.400 202.200 191.800 ;
        RECT 206.000 191.600 206.800 193.200 ;
        RECT 202.800 188.800 203.600 190.400 ;
        RECT 198.000 186.800 198.800 188.400 ;
        RECT 199.600 187.600 202.200 188.400 ;
        RECT 204.400 188.200 205.200 188.400 ;
        RECT 203.600 187.600 205.200 188.200 ;
        RECT 199.800 186.200 200.400 187.600 ;
        RECT 203.600 187.200 204.400 187.600 ;
        RECT 201.400 186.200 205.000 186.600 ;
        RECT 207.600 186.200 208.400 199.800 ;
        RECT 209.200 188.300 210.000 188.400 ;
        RECT 210.800 188.300 211.600 199.800 ;
        RECT 214.000 192.400 214.800 199.800 ;
        RECT 215.600 192.400 216.400 192.600 ;
        RECT 218.400 192.400 220.000 199.800 ;
        RECT 214.000 191.800 216.400 192.400 ;
        RECT 218.000 191.800 220.000 192.400 ;
        RECT 222.200 192.400 223.000 192.600 ;
        RECT 223.600 192.400 224.400 199.800 ;
        RECT 222.200 191.800 224.400 192.400 ;
        RECT 218.000 190.400 218.600 191.800 ;
        RECT 222.200 191.200 222.800 191.800 ;
        RECT 219.400 190.600 222.800 191.200 ;
        RECT 225.200 191.400 226.000 199.800 ;
        RECT 229.600 196.400 230.400 199.800 ;
        RECT 228.400 195.800 230.400 196.400 ;
        RECT 234.000 195.800 234.800 199.800 ;
        RECT 238.200 195.800 239.400 199.800 ;
        RECT 228.400 195.000 229.200 195.800 ;
        RECT 234.000 195.200 234.600 195.800 ;
        RECT 231.800 194.600 235.400 195.200 ;
        RECT 238.000 195.000 238.800 195.800 ;
        RECT 231.800 194.400 232.600 194.600 ;
        RECT 234.600 194.400 235.400 194.600 ;
        RECT 228.400 193.000 229.200 193.200 ;
        RECT 233.000 193.000 233.800 193.200 ;
        RECT 228.400 192.400 233.800 193.000 ;
        RECT 234.400 193.000 236.600 193.600 ;
        RECT 234.400 191.800 235.000 193.000 ;
        RECT 235.800 192.800 236.600 193.000 ;
        RECT 238.200 193.200 239.600 194.000 ;
        RECT 238.200 192.200 238.800 193.200 ;
        RECT 230.200 191.400 235.000 191.800 ;
        RECT 225.200 191.200 235.000 191.400 ;
        RECT 236.400 191.600 238.800 192.200 ;
        RECT 225.200 191.000 231.000 191.200 ;
        RECT 225.200 190.800 230.800 191.000 ;
        RECT 219.400 190.400 220.200 190.600 ;
        RECT 217.200 189.800 218.600 190.400 ;
        RECT 231.600 190.200 232.400 190.400 ;
        RECT 221.600 189.800 222.400 190.000 ;
        RECT 217.200 189.600 219.000 189.800 ;
        RECT 218.000 189.200 219.000 189.600 ;
        RECT 214.000 188.300 215.600 188.400 ;
        RECT 209.200 187.700 211.600 188.300 ;
        RECT 209.200 186.800 210.000 187.700 ;
        RECT 188.400 182.200 189.200 186.200 ;
        RECT 190.000 186.000 194.000 186.200 ;
        RECT 190.000 182.200 190.800 186.000 ;
        RECT 193.200 182.200 194.000 186.000 ;
        RECT 195.400 185.600 197.200 186.200 ;
        RECT 195.400 184.400 196.200 185.600 ;
        RECT 195.400 183.600 197.200 184.400 ;
        RECT 195.400 182.200 196.200 183.600 ;
        RECT 199.600 182.200 200.400 186.200 ;
        RECT 201.200 186.000 205.200 186.200 ;
        RECT 201.200 182.200 202.000 186.000 ;
        RECT 204.400 182.200 205.200 186.000 ;
        RECT 206.600 185.600 208.400 186.200 ;
        RECT 206.600 184.400 207.400 185.600 ;
        RECT 206.600 183.600 208.400 184.400 ;
        RECT 206.600 182.200 207.400 183.600 ;
        RECT 210.800 182.200 211.600 187.700 ;
        RECT 212.500 187.700 215.600 188.300 ;
        RECT 212.500 186.400 213.100 187.700 ;
        RECT 214.000 187.600 215.600 187.700 ;
        RECT 216.800 187.600 217.600 188.400 ;
        RECT 217.000 187.200 217.600 187.600 ;
        RECT 215.600 186.800 216.400 187.000 ;
        RECT 212.400 184.800 213.200 186.400 ;
        RECT 214.000 186.200 216.400 186.800 ;
        RECT 217.000 186.400 217.800 187.200 ;
        RECT 214.000 182.200 214.800 186.200 ;
        RECT 218.400 185.800 219.000 189.200 ;
        RECT 219.800 189.200 222.400 189.800 ;
        RECT 227.400 189.600 232.400 190.200 ;
        RECT 227.400 189.400 228.200 189.600 ;
        RECT 230.000 189.400 230.800 189.600 ;
        RECT 219.800 188.600 220.400 189.200 ;
        RECT 219.600 187.800 220.400 188.600 ;
        RECT 229.000 188.400 229.800 188.600 ;
        RECT 236.400 188.400 237.000 191.600 ;
        RECT 242.800 191.200 243.600 199.800 ;
        RECT 245.200 193.600 246.000 194.400 ;
        RECT 245.200 192.400 245.800 193.600 ;
        RECT 246.600 192.400 247.400 199.800 ;
        RECT 244.400 191.800 245.800 192.400 ;
        RECT 246.400 191.800 247.400 192.400 ;
        RECT 244.400 191.600 245.200 191.800 ;
        RECT 239.400 190.600 243.600 191.200 ;
        RECT 239.400 190.400 240.200 190.600 ;
        RECT 241.000 189.800 241.800 190.000 ;
        RECT 238.000 189.200 241.800 189.800 ;
        RECT 238.000 189.000 238.800 189.200 ;
        RECT 222.800 188.200 224.400 188.400 ;
        RECT 221.000 187.600 224.400 188.200 ;
        RECT 226.000 187.800 237.000 188.400 ;
        RECT 226.000 187.600 227.600 187.800 ;
        RECT 221.000 187.200 221.600 187.600 ;
        RECT 219.600 186.600 221.600 187.200 ;
        RECT 222.200 186.800 223.000 187.000 ;
        RECT 219.600 186.400 221.200 186.600 ;
        RECT 222.200 186.200 224.400 186.800 ;
        RECT 218.400 182.200 220.000 185.800 ;
        RECT 223.600 182.200 224.400 186.200 ;
        RECT 225.200 182.200 226.000 187.000 ;
        RECT 230.200 185.600 230.800 187.800 ;
        RECT 234.800 187.600 236.600 187.800 ;
        RECT 242.800 187.200 243.600 190.600 ;
        RECT 246.400 188.400 247.000 191.800 ;
        RECT 247.600 190.300 248.400 190.400 ;
        RECT 250.800 190.300 251.600 190.400 ;
        RECT 247.600 189.700 251.600 190.300 ;
        RECT 247.600 188.800 248.400 189.700 ;
        RECT 250.800 189.600 251.600 189.700 ;
        RECT 252.400 190.300 253.200 199.800 ;
        RECT 254.600 192.600 255.400 199.800 ;
        RECT 254.600 191.800 256.400 192.600 ;
        RECT 258.800 192.400 259.600 199.800 ;
        RECT 263.200 198.400 264.800 199.800 ;
        RECT 263.200 197.600 266.000 198.400 ;
        RECT 260.200 192.400 261.000 192.600 ;
        RECT 258.800 191.800 261.000 192.400 ;
        RECT 263.200 192.400 264.800 197.600 ;
        RECT 266.800 192.400 267.600 192.600 ;
        RECT 268.400 192.400 269.200 199.800 ;
        RECT 263.200 191.800 265.200 192.400 ;
        RECT 266.800 191.800 269.200 192.400 ;
        RECT 255.600 191.600 256.400 191.800 ;
        RECT 254.000 190.300 254.800 191.200 ;
        RECT 252.400 189.700 254.800 190.300 ;
        RECT 244.400 187.600 247.000 188.400 ;
        RECT 249.200 188.200 250.000 188.400 ;
        RECT 248.400 187.600 250.000 188.200 ;
        RECT 239.800 186.600 243.600 187.200 ;
        RECT 239.800 186.400 240.600 186.600 ;
        RECT 228.400 184.200 229.200 185.000 ;
        RECT 230.000 184.800 230.800 185.600 ;
        RECT 231.800 185.400 232.600 185.600 ;
        RECT 231.800 184.800 234.600 185.400 ;
        RECT 234.000 184.200 234.600 184.800 ;
        RECT 238.000 184.200 238.800 185.000 ;
        RECT 228.400 183.600 230.400 184.200 ;
        RECT 229.600 182.200 230.400 183.600 ;
        RECT 234.000 182.200 234.800 184.200 ;
        RECT 238.000 183.600 239.400 184.200 ;
        RECT 238.200 182.200 239.400 183.600 ;
        RECT 242.800 182.200 243.600 186.600 ;
        RECT 244.600 186.200 245.200 187.600 ;
        RECT 248.400 187.200 249.200 187.600 ;
        RECT 246.200 186.200 249.800 186.600 ;
        RECT 244.400 182.200 245.200 186.200 ;
        RECT 246.000 186.000 250.000 186.200 ;
        RECT 246.000 182.200 246.800 186.000 ;
        RECT 249.200 182.200 250.000 186.000 ;
        RECT 250.800 184.800 251.600 186.400 ;
        RECT 252.400 182.200 253.200 189.700 ;
        RECT 254.000 189.600 254.800 189.700 ;
        RECT 255.600 188.400 256.200 191.600 ;
        RECT 260.400 191.200 261.000 191.800 ;
        RECT 260.400 190.600 263.800 191.200 ;
        RECT 263.000 190.400 263.800 190.600 ;
        RECT 264.600 190.400 265.200 191.800 ;
        RECT 260.800 189.800 261.600 190.000 ;
        RECT 264.600 189.800 266.000 190.400 ;
        RECT 260.800 189.200 263.400 189.800 ;
        RECT 262.800 188.600 263.400 189.200 ;
        RECT 264.200 189.600 266.000 189.800 ;
        RECT 264.200 189.200 265.200 189.600 ;
        RECT 255.600 187.600 256.400 188.400 ;
        RECT 258.800 188.200 260.400 188.400 ;
        RECT 258.800 187.600 262.200 188.200 ;
        RECT 262.800 187.800 263.600 188.600 ;
        RECT 255.600 184.200 256.200 187.600 ;
        RECT 261.600 187.200 262.200 187.600 ;
        RECT 260.200 186.800 261.000 187.000 ;
        RECT 257.200 184.800 258.000 186.400 ;
        RECT 258.800 186.200 261.000 186.800 ;
        RECT 261.600 186.600 263.600 187.200 ;
        RECT 262.000 186.400 263.600 186.600 ;
        RECT 255.600 182.200 256.400 184.200 ;
        RECT 258.800 182.200 259.600 186.200 ;
        RECT 264.200 185.800 264.800 189.200 ;
        RECT 265.600 187.600 266.400 188.400 ;
        RECT 267.600 188.300 269.200 188.400 ;
        RECT 270.000 188.300 270.800 188.400 ;
        RECT 267.600 187.700 270.800 188.300 ;
        RECT 267.600 187.600 269.200 187.700 ;
        RECT 265.600 187.200 266.200 187.600 ;
        RECT 265.400 186.400 266.200 187.200 ;
        RECT 266.800 186.800 267.600 187.000 ;
        RECT 270.000 186.800 270.800 187.700 ;
        RECT 266.800 186.200 269.200 186.800 ;
        RECT 263.200 182.200 264.800 185.800 ;
        RECT 268.400 182.200 269.200 186.200 ;
        RECT 271.600 186.200 272.400 199.800 ;
        RECT 273.200 191.600 274.000 193.200 ;
        RECT 274.800 191.400 275.600 199.800 ;
        RECT 279.200 196.400 280.000 199.800 ;
        RECT 278.000 195.800 280.000 196.400 ;
        RECT 283.600 195.800 284.400 199.800 ;
        RECT 287.800 195.800 289.000 199.800 ;
        RECT 278.000 195.000 278.800 195.800 ;
        RECT 283.600 195.200 284.200 195.800 ;
        RECT 281.400 194.600 285.000 195.200 ;
        RECT 287.600 195.000 288.400 195.800 ;
        RECT 281.400 194.400 282.200 194.600 ;
        RECT 284.200 194.400 285.000 194.600 ;
        RECT 278.000 193.000 278.800 193.200 ;
        RECT 282.600 193.000 283.400 193.200 ;
        RECT 278.000 192.400 283.400 193.000 ;
        RECT 284.000 193.000 286.200 193.600 ;
        RECT 284.000 191.800 284.600 193.000 ;
        RECT 285.400 192.800 286.200 193.000 ;
        RECT 287.800 193.200 289.200 194.000 ;
        RECT 287.800 192.200 288.400 193.200 ;
        RECT 279.800 191.400 284.600 191.800 ;
        RECT 274.800 191.200 284.600 191.400 ;
        RECT 286.000 191.600 288.400 192.200 ;
        RECT 274.800 191.000 280.600 191.200 ;
        RECT 274.800 190.800 280.400 191.000 ;
        RECT 281.200 190.200 282.000 190.400 ;
        RECT 277.000 189.600 282.000 190.200 ;
        RECT 277.000 189.400 277.800 189.600 ;
        RECT 279.600 189.400 280.400 189.600 ;
        RECT 278.600 188.400 279.400 188.600 ;
        RECT 286.000 188.400 286.600 191.600 ;
        RECT 292.400 191.200 293.200 199.800 ;
        RECT 289.000 190.600 293.200 191.200 ;
        RECT 289.000 190.400 289.800 190.600 ;
        RECT 290.600 189.800 291.400 190.000 ;
        RECT 287.600 189.200 291.400 189.800 ;
        RECT 287.600 189.000 288.400 189.200 ;
        RECT 275.600 187.800 286.600 188.400 ;
        RECT 275.600 187.600 277.200 187.800 ;
        RECT 271.600 185.600 273.400 186.200 ;
        RECT 272.600 184.400 273.400 185.600 ;
        RECT 272.600 183.600 274.000 184.400 ;
        RECT 272.600 182.200 273.400 183.600 ;
        RECT 274.800 182.200 275.600 187.000 ;
        RECT 279.800 185.600 280.400 187.800 ;
        RECT 285.400 187.600 286.200 187.800 ;
        RECT 292.400 187.200 293.200 190.600 ;
        RECT 300.400 190.300 301.200 199.800 ;
        RECT 305.200 194.300 306.000 199.800 ;
        RECT 306.800 194.300 307.600 194.400 ;
        RECT 305.200 193.700 307.600 194.300 ;
        RECT 302.000 192.300 302.800 193.200 ;
        RECT 303.600 192.300 304.400 193.200 ;
        RECT 302.000 191.700 304.400 192.300 ;
        RECT 302.000 191.600 302.800 191.700 ;
        RECT 303.600 191.600 304.400 191.700 ;
        RECT 303.600 190.300 304.400 190.400 ;
        RECT 300.400 189.700 304.400 190.300 ;
        RECT 289.400 186.600 293.200 187.200 ;
        RECT 298.800 186.800 299.600 188.400 ;
        RECT 289.400 186.400 290.200 186.600 ;
        RECT 278.000 184.200 278.800 185.000 ;
        RECT 279.600 184.800 280.400 185.600 ;
        RECT 281.400 185.400 282.200 185.600 ;
        RECT 281.400 184.800 284.200 185.400 ;
        RECT 283.600 184.200 284.200 184.800 ;
        RECT 287.600 184.200 288.400 185.000 ;
        RECT 278.000 183.600 280.000 184.200 ;
        RECT 279.200 182.200 280.000 183.600 ;
        RECT 283.600 182.200 284.400 184.200 ;
        RECT 287.600 183.600 289.000 184.200 ;
        RECT 287.800 182.200 289.000 183.600 ;
        RECT 292.400 182.200 293.200 186.600 ;
        RECT 300.400 186.200 301.200 189.700 ;
        RECT 303.600 189.600 304.400 189.700 ;
        RECT 305.200 186.200 306.000 193.700 ;
        RECT 306.800 193.600 307.600 193.700 ;
        RECT 306.800 188.300 307.600 188.400 ;
        RECT 308.400 188.300 309.200 199.800 ;
        RECT 312.400 193.600 313.200 194.400 ;
        RECT 312.400 192.400 313.000 193.600 ;
        RECT 313.800 192.400 314.600 199.800 ;
        RECT 311.600 191.800 313.000 192.400 ;
        RECT 313.600 191.800 314.600 192.400 ;
        RECT 311.600 191.600 312.400 191.800 ;
        RECT 313.600 188.400 314.200 191.800 ;
        RECT 314.800 188.800 315.600 190.400 ;
        RECT 306.800 187.700 309.200 188.300 ;
        RECT 306.800 186.800 307.600 187.700 ;
        RECT 300.400 185.600 302.200 186.200 ;
        RECT 301.400 182.200 302.200 185.600 ;
        RECT 304.200 185.600 306.000 186.200 ;
        RECT 304.200 182.200 305.000 185.600 ;
        RECT 308.400 182.200 309.200 187.700 ;
        RECT 310.000 186.800 310.800 188.400 ;
        RECT 311.600 187.600 314.200 188.400 ;
        RECT 316.400 188.300 317.200 188.400 ;
        RECT 318.000 188.300 318.800 188.400 ;
        RECT 316.400 188.200 318.800 188.300 ;
        RECT 315.600 187.700 318.800 188.200 ;
        RECT 315.600 187.600 317.200 187.700 ;
        RECT 311.800 186.200 312.400 187.600 ;
        RECT 315.600 187.200 316.400 187.600 ;
        RECT 318.000 186.800 318.800 187.700 ;
        RECT 313.400 186.200 317.000 186.600 ;
        RECT 319.600 186.200 320.400 199.800 ;
        RECT 321.200 191.600 322.000 193.200 ;
        RECT 322.800 192.400 323.600 199.800 ;
        RECT 327.200 198.400 328.800 199.800 ;
        RECT 326.000 197.600 328.800 198.400 ;
        RECT 324.200 192.400 325.000 192.600 ;
        RECT 322.800 191.800 325.000 192.400 ;
        RECT 327.200 192.400 328.800 197.600 ;
        RECT 330.800 192.400 331.600 192.600 ;
        RECT 332.400 192.400 333.200 199.800 ;
        RECT 327.200 191.800 329.200 192.400 ;
        RECT 330.800 191.800 333.200 192.400 ;
        RECT 336.600 192.400 337.400 199.800 ;
        RECT 338.000 193.600 338.800 194.400 ;
        RECT 338.200 192.400 338.800 193.600 ;
        RECT 336.600 191.800 337.600 192.400 ;
        RECT 338.200 191.800 339.600 192.400 ;
        RECT 324.400 191.200 325.000 191.800 ;
        RECT 324.400 190.600 327.800 191.200 ;
        RECT 327.000 190.400 327.800 190.600 ;
        RECT 328.600 190.400 329.200 191.800 ;
        RECT 324.800 189.800 325.600 190.000 ;
        RECT 328.600 189.800 330.000 190.400 ;
        RECT 324.800 189.200 327.400 189.800 ;
        RECT 326.800 188.600 327.400 189.200 ;
        RECT 328.200 189.600 330.000 189.800 ;
        RECT 328.200 189.200 329.200 189.600 ;
        RECT 322.800 188.200 324.400 188.400 ;
        RECT 322.800 187.600 326.200 188.200 ;
        RECT 326.800 187.800 327.600 188.600 ;
        RECT 325.600 187.200 326.200 187.600 ;
        RECT 324.200 186.800 325.000 187.000 ;
        RECT 322.800 186.200 325.000 186.800 ;
        RECT 325.600 186.600 327.600 187.200 ;
        RECT 326.000 186.400 327.600 186.600 ;
        RECT 311.600 182.200 312.400 186.200 ;
        RECT 313.200 186.000 317.200 186.200 ;
        RECT 313.200 182.200 314.000 186.000 ;
        RECT 316.400 182.200 317.200 186.000 ;
        RECT 319.600 185.600 321.400 186.200 ;
        RECT 320.600 184.400 321.400 185.600 ;
        RECT 320.600 183.600 322.000 184.400 ;
        RECT 320.600 182.200 321.400 183.600 ;
        RECT 322.800 182.200 323.600 186.200 ;
        RECT 328.200 185.800 328.800 189.200 ;
        RECT 335.600 188.800 336.400 190.400 ;
        RECT 337.000 188.400 337.600 191.800 ;
        RECT 338.800 191.600 339.600 191.800 ;
        RECT 329.600 187.600 330.400 188.400 ;
        RECT 331.600 188.300 333.200 188.400 ;
        RECT 334.000 188.300 334.800 188.400 ;
        RECT 331.600 188.200 334.800 188.300 ;
        RECT 337.000 188.300 339.600 188.400 ;
        RECT 340.400 188.300 341.200 188.400 ;
        RECT 331.600 187.700 335.600 188.200 ;
        RECT 331.600 187.600 333.200 187.700 ;
        RECT 334.000 187.600 335.600 187.700 ;
        RECT 337.000 187.700 341.200 188.300 ;
        RECT 337.000 187.600 339.600 187.700 ;
        RECT 329.600 187.200 330.200 187.600 ;
        RECT 334.800 187.200 335.600 187.600 ;
        RECT 329.400 186.400 330.200 187.200 ;
        RECT 330.800 186.800 331.600 187.000 ;
        RECT 330.800 186.200 333.200 186.800 ;
        RECT 334.200 186.200 337.800 186.600 ;
        RECT 338.800 186.200 339.400 187.600 ;
        RECT 340.400 186.800 341.200 187.700 ;
        RECT 342.000 186.200 342.800 199.800 ;
        RECT 343.600 191.600 344.400 193.200 ;
        RECT 345.200 192.400 346.000 199.800 ;
        RECT 349.600 198.400 351.200 199.800 ;
        RECT 349.600 197.600 352.400 198.400 ;
        RECT 346.800 192.400 347.600 192.600 ;
        RECT 349.600 192.400 351.200 197.600 ;
        RECT 345.200 191.800 347.600 192.400 ;
        RECT 349.200 191.800 351.200 192.400 ;
        RECT 353.400 192.400 354.200 192.600 ;
        RECT 354.800 192.400 355.600 199.800 ;
        RECT 353.400 191.800 355.600 192.400 ;
        RECT 349.200 190.400 349.800 191.800 ;
        RECT 353.400 191.200 354.000 191.800 ;
        RECT 350.600 190.600 354.000 191.200 ;
        RECT 356.400 191.400 357.200 199.800 ;
        RECT 360.800 196.400 361.600 199.800 ;
        RECT 359.600 195.800 361.600 196.400 ;
        RECT 365.200 195.800 366.000 199.800 ;
        RECT 369.400 195.800 370.600 199.800 ;
        RECT 359.600 195.000 360.400 195.800 ;
        RECT 365.200 195.200 365.800 195.800 ;
        RECT 363.000 194.600 366.600 195.200 ;
        RECT 369.200 195.000 370.000 195.800 ;
        RECT 363.000 194.400 363.800 194.600 ;
        RECT 365.800 194.400 366.600 194.600 ;
        RECT 359.600 193.000 360.400 193.200 ;
        RECT 364.200 193.000 365.000 193.200 ;
        RECT 359.600 192.400 365.000 193.000 ;
        RECT 365.600 193.000 367.800 193.600 ;
        RECT 365.600 191.800 366.200 193.000 ;
        RECT 367.000 192.800 367.800 193.000 ;
        RECT 369.400 193.200 370.800 194.000 ;
        RECT 369.400 192.200 370.000 193.200 ;
        RECT 361.400 191.400 366.200 191.800 ;
        RECT 356.400 191.200 366.200 191.400 ;
        RECT 367.600 191.600 370.000 192.200 ;
        RECT 356.400 191.000 362.200 191.200 ;
        RECT 356.400 190.800 362.000 191.000 ;
        RECT 350.600 190.400 351.400 190.600 ;
        RECT 348.400 189.800 349.800 190.400 ;
        RECT 362.800 190.200 363.600 190.400 ;
        RECT 352.800 189.800 353.600 190.000 ;
        RECT 348.400 189.600 350.200 189.800 ;
        RECT 349.200 189.200 350.200 189.600 ;
        RECT 345.200 187.600 346.800 188.400 ;
        RECT 348.000 187.600 348.800 188.400 ;
        RECT 348.200 187.200 348.800 187.600 ;
        RECT 346.800 186.800 347.600 187.000 ;
        RECT 345.200 186.200 347.600 186.800 ;
        RECT 348.200 186.400 349.000 187.200 ;
        RECT 327.200 182.200 328.800 185.800 ;
        RECT 332.400 182.200 333.200 186.200 ;
        RECT 334.000 186.000 338.000 186.200 ;
        RECT 334.000 182.200 334.800 186.000 ;
        RECT 337.200 182.200 338.000 186.000 ;
        RECT 338.800 182.200 339.600 186.200 ;
        RECT 342.000 185.600 343.800 186.200 ;
        RECT 343.000 182.200 343.800 185.600 ;
        RECT 345.200 182.200 346.000 186.200 ;
        RECT 349.600 185.800 350.200 189.200 ;
        RECT 351.000 189.200 353.600 189.800 ;
        RECT 358.600 189.600 363.600 190.200 ;
        RECT 358.600 189.400 359.400 189.600 ;
        RECT 361.200 189.400 362.000 189.600 ;
        RECT 351.000 188.600 351.600 189.200 ;
        RECT 350.800 187.800 351.600 188.600 ;
        RECT 360.200 188.400 361.000 188.600 ;
        RECT 367.600 188.400 368.200 191.600 ;
        RECT 374.000 191.200 374.800 199.800 ;
        RECT 370.600 190.600 374.800 191.200 ;
        RECT 375.600 195.000 376.400 199.000 ;
        RECT 379.800 198.400 380.600 199.800 ;
        RECT 379.800 197.600 381.200 198.400 ;
        RECT 375.600 191.600 376.200 195.000 ;
        RECT 379.800 192.800 380.600 197.600 ;
        RECT 386.000 193.600 386.800 194.400 ;
        RECT 379.800 192.200 381.400 192.800 ;
        RECT 386.000 192.400 386.600 193.600 ;
        RECT 387.400 192.400 388.200 199.800 ;
        RECT 394.200 198.400 395.000 199.800 ;
        RECT 393.200 197.600 395.000 198.400 ;
        RECT 394.200 192.600 395.000 197.600 ;
        RECT 375.600 191.000 379.400 191.600 ;
        RECT 370.600 190.400 371.400 190.600 ;
        RECT 374.000 190.300 374.800 190.600 ;
        RECT 375.600 190.300 376.400 190.400 ;
        RECT 372.200 189.800 373.000 190.000 ;
        RECT 369.200 189.200 373.000 189.800 ;
        RECT 374.000 189.700 376.400 190.300 ;
        RECT 369.200 189.000 370.000 189.200 ;
        RECT 354.000 188.200 355.600 188.400 ;
        RECT 352.200 187.600 355.600 188.200 ;
        RECT 357.200 187.800 368.200 188.400 ;
        RECT 357.200 187.600 358.800 187.800 ;
        RECT 352.200 187.200 352.800 187.600 ;
        RECT 350.800 186.600 352.800 187.200 ;
        RECT 353.400 186.800 354.200 187.000 ;
        RECT 350.800 186.400 352.400 186.600 ;
        RECT 353.400 186.200 355.600 186.800 ;
        RECT 349.600 182.200 351.200 185.800 ;
        RECT 354.800 182.200 355.600 186.200 ;
        RECT 356.400 182.200 357.200 187.000 ;
        RECT 361.400 185.600 362.000 187.800 ;
        RECT 367.000 187.600 367.800 187.800 ;
        RECT 374.000 187.200 374.800 189.700 ;
        RECT 375.600 188.800 376.400 189.700 ;
        RECT 377.200 188.800 378.000 190.400 ;
        RECT 378.800 189.000 379.400 191.000 ;
        RECT 378.800 188.200 380.200 189.000 ;
        RECT 380.800 188.400 381.400 192.200 ;
        RECT 385.200 191.800 386.600 192.400 ;
        RECT 387.200 191.800 388.200 192.400 ;
        RECT 393.200 191.800 395.000 192.600 ;
        RECT 397.000 192.600 397.800 199.800 ;
        RECT 397.000 191.800 398.800 192.600 ;
        RECT 385.200 191.600 386.000 191.800 ;
        RECT 382.000 189.600 382.800 191.200 ;
        RECT 383.600 190.300 384.400 190.400 ;
        RECT 385.300 190.300 385.900 191.600 ;
        RECT 383.600 189.700 385.900 190.300 ;
        RECT 383.600 189.600 384.400 189.700 ;
        RECT 387.200 188.400 387.800 191.800 ;
        RECT 388.400 188.800 389.200 190.400 ;
        RECT 393.400 188.400 394.000 191.800 ;
        RECT 394.800 189.600 395.600 191.200 ;
        RECT 396.400 189.600 397.200 191.200 ;
        RECT 378.800 187.800 379.800 188.200 ;
        RECT 371.000 186.600 374.800 187.200 ;
        RECT 371.000 186.400 371.800 186.600 ;
        RECT 359.600 184.200 360.400 185.000 ;
        RECT 361.200 184.800 362.000 185.600 ;
        RECT 363.000 185.400 363.800 185.600 ;
        RECT 363.000 184.800 365.800 185.400 ;
        RECT 365.200 184.200 365.800 184.800 ;
        RECT 369.200 184.200 370.000 185.000 ;
        RECT 359.600 183.600 361.600 184.200 ;
        RECT 360.800 182.200 361.600 183.600 ;
        RECT 365.200 182.200 366.000 184.200 ;
        RECT 369.200 183.600 370.600 184.200 ;
        RECT 369.400 182.200 370.600 183.600 ;
        RECT 374.000 182.200 374.800 186.600 ;
        RECT 375.600 187.200 379.800 187.800 ;
        RECT 380.800 187.600 382.800 188.400 ;
        RECT 385.200 187.600 387.800 188.400 ;
        RECT 390.000 188.200 390.800 188.400 ;
        RECT 389.200 187.600 390.800 188.200 ;
        RECT 393.200 187.600 394.000 188.400 ;
        RECT 394.900 188.300 395.500 189.600 ;
        RECT 398.000 188.400 398.600 191.800 ;
        RECT 398.000 188.300 398.800 188.400 ;
        RECT 394.900 187.700 398.800 188.300 ;
        RECT 375.600 185.000 376.200 187.200 ;
        RECT 380.800 187.000 381.400 187.600 ;
        RECT 380.600 186.600 381.400 187.000 ;
        RECT 379.800 186.000 381.400 186.600 ;
        RECT 385.400 186.200 386.000 187.600 ;
        RECT 389.200 187.200 390.000 187.600 ;
        RECT 387.000 186.200 390.600 186.600 ;
        RECT 375.600 183.000 376.400 185.000 ;
        RECT 379.800 183.000 380.600 186.000 ;
        RECT 385.200 182.200 386.000 186.200 ;
        RECT 386.800 186.000 390.800 186.200 ;
        RECT 386.800 182.200 387.600 186.000 ;
        RECT 390.000 182.200 390.800 186.000 ;
        RECT 391.600 184.800 392.400 186.400 ;
        RECT 393.400 184.200 394.000 187.600 ;
        RECT 393.200 182.200 394.000 184.200 ;
        RECT 398.000 187.600 398.800 187.700 ;
        RECT 398.000 184.200 398.600 187.600 ;
        RECT 399.600 184.800 400.400 186.400 ;
        RECT 401.200 184.800 402.000 186.400 ;
        RECT 398.000 182.200 398.800 184.200 ;
        RECT 402.800 182.200 403.600 199.800 ;
        RECT 407.000 192.600 407.800 199.800 ;
        RECT 406.000 191.800 407.800 192.600 ;
        RECT 406.200 188.400 406.800 191.800 ;
        RECT 409.200 191.200 410.000 199.800 ;
        RECT 413.400 195.800 414.600 199.800 ;
        RECT 418.000 195.800 418.800 199.800 ;
        RECT 422.400 196.400 423.200 199.800 ;
        RECT 422.400 195.800 424.400 196.400 ;
        RECT 414.000 195.000 414.800 195.800 ;
        RECT 418.200 195.200 418.800 195.800 ;
        RECT 417.400 194.600 421.000 195.200 ;
        RECT 423.600 195.000 424.400 195.800 ;
        RECT 417.400 194.400 418.200 194.600 ;
        RECT 420.200 194.400 421.000 194.600 ;
        RECT 413.200 193.200 414.600 194.000 ;
        RECT 414.000 192.200 414.600 193.200 ;
        RECT 416.200 193.000 418.400 193.600 ;
        RECT 416.200 192.800 417.000 193.000 ;
        RECT 414.000 191.600 416.400 192.200 ;
        RECT 407.600 189.600 408.400 191.200 ;
        RECT 409.200 190.600 413.400 191.200 ;
        RECT 406.000 187.600 406.800 188.400 ;
        RECT 404.400 184.800 405.200 186.400 ;
        RECT 406.200 186.300 406.800 187.600 ;
        RECT 409.200 187.200 410.000 190.600 ;
        RECT 412.600 190.400 413.400 190.600 ;
        RECT 411.000 189.800 411.800 190.000 ;
        RECT 411.000 189.200 414.800 189.800 ;
        RECT 414.000 189.000 414.800 189.200 ;
        RECT 415.800 188.400 416.400 191.600 ;
        RECT 417.800 191.800 418.400 193.000 ;
        RECT 419.000 193.000 419.800 193.200 ;
        RECT 423.600 193.000 424.400 193.200 ;
        RECT 419.000 192.400 424.400 193.000 ;
        RECT 417.800 191.400 422.600 191.800 ;
        RECT 426.800 191.400 427.600 199.800 ;
        RECT 417.800 191.200 427.600 191.400 ;
        RECT 421.800 191.000 427.600 191.200 ;
        RECT 422.000 190.800 427.600 191.000 ;
        RECT 428.400 191.400 429.200 199.800 ;
        RECT 432.800 196.400 433.600 199.800 ;
        RECT 431.600 195.800 433.600 196.400 ;
        RECT 437.200 195.800 438.000 199.800 ;
        RECT 441.400 195.800 442.600 199.800 ;
        RECT 446.000 198.300 446.800 199.800 ;
        RECT 450.800 198.300 451.600 198.400 ;
        RECT 446.000 197.700 451.600 198.300 ;
        RECT 431.600 195.000 432.400 195.800 ;
        RECT 437.200 195.200 437.800 195.800 ;
        RECT 435.000 194.600 438.600 195.200 ;
        RECT 441.200 195.000 442.000 195.800 ;
        RECT 435.000 194.400 435.800 194.600 ;
        RECT 437.800 194.400 438.600 194.600 ;
        RECT 431.600 193.000 432.400 193.200 ;
        RECT 436.200 193.000 437.000 193.200 ;
        RECT 431.600 192.400 437.000 193.000 ;
        RECT 437.600 193.000 439.800 193.600 ;
        RECT 437.600 191.800 438.200 193.000 ;
        RECT 439.000 192.800 439.800 193.000 ;
        RECT 441.400 193.200 442.800 194.000 ;
        RECT 441.400 192.200 442.000 193.200 ;
        RECT 433.400 191.400 438.200 191.800 ;
        RECT 428.400 191.200 438.200 191.400 ;
        RECT 439.600 191.600 442.000 192.200 ;
        RECT 428.400 191.000 434.200 191.200 ;
        RECT 428.400 190.800 434.000 191.000 ;
        RECT 420.400 190.200 421.200 190.400 ;
        RECT 434.800 190.200 435.600 190.400 ;
        RECT 420.400 189.600 425.400 190.200 ;
        RECT 424.600 189.400 425.400 189.600 ;
        RECT 430.600 189.600 435.600 190.200 ;
        RECT 430.600 189.400 431.400 189.600 ;
        RECT 433.200 189.400 434.000 189.600 ;
        RECT 423.000 188.400 423.800 188.600 ;
        RECT 432.200 188.400 433.000 188.600 ;
        RECT 439.600 188.400 440.200 191.600 ;
        RECT 446.000 191.200 446.800 197.700 ;
        RECT 450.800 197.600 451.600 197.700 ;
        RECT 452.400 192.400 453.200 199.800 ;
        RECT 455.600 192.400 456.400 199.800 ;
        RECT 452.400 191.800 456.400 192.400 ;
        RECT 457.200 192.300 458.000 199.800 ;
        RECT 459.600 193.600 460.400 194.400 ;
        RECT 459.600 192.400 460.200 193.600 ;
        RECT 461.000 192.400 461.800 199.800 ;
        RECT 458.800 192.300 460.200 192.400 ;
        RECT 457.200 191.800 460.200 192.300 ;
        RECT 460.800 191.800 461.800 192.400 ;
        RECT 465.200 192.400 466.000 199.800 ;
        RECT 469.600 198.400 471.200 199.800 ;
        RECT 469.600 197.600 472.400 198.400 ;
        RECT 466.600 192.400 467.400 192.600 ;
        RECT 465.200 191.800 467.400 192.400 ;
        RECT 469.600 192.400 471.200 197.600 ;
        RECT 473.200 192.400 474.000 192.600 ;
        RECT 474.800 192.400 475.600 199.800 ;
        RECT 469.600 191.800 471.600 192.400 ;
        RECT 473.200 191.800 475.600 192.400 ;
        RECT 479.000 192.400 479.800 199.800 ;
        RECT 480.400 193.600 481.200 194.400 ;
        RECT 480.600 192.400 481.200 193.600 ;
        RECT 479.000 191.800 480.000 192.400 ;
        RECT 480.600 192.300 482.000 192.400 ;
        RECT 482.800 192.300 483.600 199.800 ;
        RECT 480.600 191.800 483.600 192.300 ;
        RECT 488.600 192.400 489.400 199.800 ;
        RECT 490.000 193.600 490.800 194.400 ;
        RECT 490.200 192.400 490.800 193.600 ;
        RECT 492.400 192.400 493.200 199.800 ;
        RECT 495.600 192.400 496.400 199.800 ;
        RECT 488.600 191.800 489.600 192.400 ;
        RECT 490.200 191.800 491.600 192.400 ;
        RECT 492.400 191.800 496.400 192.400 ;
        RECT 497.200 191.800 498.000 199.800 ;
        RECT 498.800 192.400 499.600 199.800 ;
        RECT 503.200 198.400 504.800 199.800 ;
        RECT 503.200 197.600 506.000 198.400 ;
        RECT 500.400 192.400 501.200 192.600 ;
        RECT 503.200 192.400 504.800 197.600 ;
        RECT 498.800 191.800 501.200 192.400 ;
        RECT 502.800 191.800 504.800 192.400 ;
        RECT 507.000 192.400 507.800 192.600 ;
        RECT 508.400 192.400 509.200 199.800 ;
        RECT 507.000 191.800 509.200 192.400 ;
        RECT 442.600 190.600 446.800 191.200 ;
        RECT 457.200 191.700 459.600 191.800 ;
        RECT 442.600 190.400 443.400 190.600 ;
        RECT 444.200 189.800 445.000 190.000 ;
        RECT 441.200 189.200 445.000 189.800 ;
        RECT 441.200 189.000 442.000 189.200 ;
        RECT 415.800 187.800 426.800 188.400 ;
        RECT 416.200 187.600 417.000 187.800 ;
        RECT 409.200 186.600 413.000 187.200 ;
        RECT 407.600 186.300 408.400 186.400 ;
        RECT 406.100 185.700 408.400 186.300 ;
        RECT 406.200 184.200 406.800 185.700 ;
        RECT 407.600 185.600 408.400 185.700 ;
        RECT 406.000 182.200 406.800 184.200 ;
        RECT 409.200 182.200 410.000 186.600 ;
        RECT 412.200 186.400 413.000 186.600 ;
        RECT 422.000 185.600 422.600 187.800 ;
        RECT 425.200 187.600 426.800 187.800 ;
        RECT 429.200 187.800 440.200 188.400 ;
        RECT 429.200 187.600 430.800 187.800 ;
        RECT 420.200 185.400 421.000 185.600 ;
        RECT 414.000 184.200 414.800 185.000 ;
        RECT 418.200 184.800 421.000 185.400 ;
        RECT 422.000 184.800 422.800 185.600 ;
        RECT 418.200 184.200 418.800 184.800 ;
        RECT 423.600 184.200 424.400 185.000 ;
        RECT 413.400 183.600 414.800 184.200 ;
        RECT 413.400 182.200 414.600 183.600 ;
        RECT 418.000 182.200 418.800 184.200 ;
        RECT 422.400 183.600 424.400 184.200 ;
        RECT 422.400 182.200 423.200 183.600 ;
        RECT 426.800 182.200 427.600 187.000 ;
        RECT 428.400 182.200 429.200 187.000 ;
        RECT 433.400 186.400 434.000 187.800 ;
        RECT 439.000 187.600 439.800 187.800 ;
        RECT 446.000 187.200 446.800 190.600 ;
        RECT 453.200 190.400 454.000 190.800 ;
        RECT 457.200 190.400 457.800 191.700 ;
        RECT 458.800 191.600 459.600 191.700 ;
        RECT 452.400 189.800 454.000 190.400 ;
        RECT 455.600 189.800 458.000 190.400 ;
        RECT 452.400 189.600 453.200 189.800 ;
        RECT 454.000 187.600 454.800 189.200 ;
        RECT 443.000 186.600 446.800 187.200 ;
        RECT 443.000 186.400 443.800 186.600 ;
        RECT 431.600 184.200 432.400 185.000 ;
        RECT 433.200 184.800 434.000 186.400 ;
        RECT 435.000 185.400 435.800 185.600 ;
        RECT 435.000 184.800 437.800 185.400 ;
        RECT 437.200 184.200 437.800 184.800 ;
        RECT 441.200 184.200 442.000 185.000 ;
        RECT 431.600 183.600 433.600 184.200 ;
        RECT 432.800 182.200 433.600 183.600 ;
        RECT 437.200 182.200 438.000 184.200 ;
        RECT 441.200 183.600 442.600 184.200 ;
        RECT 441.400 182.200 442.600 183.600 ;
        RECT 446.000 182.200 446.800 186.600 ;
        RECT 455.600 186.200 456.200 189.800 ;
        RECT 457.200 189.600 458.000 189.800 ;
        RECT 460.800 188.400 461.400 191.800 ;
        RECT 466.800 191.200 467.400 191.800 ;
        RECT 466.800 190.600 470.200 191.200 ;
        RECT 469.400 190.400 470.200 190.600 ;
        RECT 471.000 190.400 471.600 191.800 ;
        RECT 462.000 188.800 462.800 190.400 ;
        RECT 467.200 189.800 468.000 190.000 ;
        RECT 471.000 189.800 472.400 190.400 ;
        RECT 467.200 189.200 469.800 189.800 ;
        RECT 469.200 188.600 469.800 189.200 ;
        RECT 470.600 189.600 472.400 189.800 ;
        RECT 470.600 189.200 471.600 189.600 ;
        RECT 458.800 187.600 461.400 188.400 ;
        RECT 463.600 188.200 464.400 188.400 ;
        RECT 462.800 187.600 464.400 188.200 ;
        RECT 465.200 188.200 466.800 188.400 ;
        RECT 465.200 187.600 468.600 188.200 ;
        RECT 469.200 187.800 470.000 188.600 ;
        RECT 455.600 182.200 456.400 186.200 ;
        RECT 457.200 185.600 458.000 186.400 ;
        RECT 459.000 186.200 459.600 187.600 ;
        RECT 462.800 187.200 463.600 187.600 ;
        RECT 468.000 187.200 468.600 187.600 ;
        RECT 466.600 186.800 467.400 187.000 ;
        RECT 460.600 186.200 464.200 186.600 ;
        RECT 465.200 186.200 467.400 186.800 ;
        RECT 468.000 186.600 470.000 187.200 ;
        RECT 468.400 186.400 470.000 186.600 ;
        RECT 457.000 184.800 457.800 185.600 ;
        RECT 458.800 182.200 459.600 186.200 ;
        RECT 460.400 186.000 464.400 186.200 ;
        RECT 460.400 182.200 461.200 186.000 ;
        RECT 463.600 182.200 464.400 186.000 ;
        RECT 465.200 182.200 466.000 186.200 ;
        RECT 470.600 185.800 471.200 189.200 ;
        RECT 478.000 188.800 478.800 190.400 ;
        RECT 479.400 188.400 480.000 191.800 ;
        RECT 481.200 191.700 483.600 191.800 ;
        RECT 481.200 191.600 482.000 191.700 ;
        RECT 472.000 187.600 472.800 188.400 ;
        RECT 474.000 187.600 475.600 188.400 ;
        RECT 476.400 188.200 477.200 188.400 ;
        RECT 476.400 187.600 478.000 188.200 ;
        RECT 479.400 187.600 482.000 188.400 ;
        RECT 472.000 187.200 472.600 187.600 ;
        RECT 477.200 187.200 478.000 187.600 ;
        RECT 471.800 186.400 472.600 187.200 ;
        RECT 473.200 186.800 474.000 187.000 ;
        RECT 473.200 186.200 475.600 186.800 ;
        RECT 476.600 186.200 480.200 186.600 ;
        RECT 481.200 186.200 481.800 187.600 ;
        RECT 469.600 182.200 471.200 185.800 ;
        RECT 474.800 182.200 475.600 186.200 ;
        RECT 476.400 186.000 480.400 186.200 ;
        RECT 476.400 182.200 477.200 186.000 ;
        RECT 479.600 182.200 480.400 186.000 ;
        RECT 481.200 182.200 482.000 186.200 ;
        RECT 482.800 182.200 483.600 191.700 ;
        RECT 487.600 188.800 488.400 190.400 ;
        RECT 489.000 188.400 489.600 191.800 ;
        RECT 490.800 191.600 491.600 191.800 ;
        RECT 493.200 190.400 494.000 190.800 ;
        RECT 497.200 190.400 497.800 191.800 ;
        RECT 502.800 190.400 503.400 191.800 ;
        RECT 507.000 191.200 507.600 191.800 ;
        RECT 504.200 190.600 507.600 191.200 ;
        RECT 504.200 190.400 505.000 190.600 ;
        RECT 492.400 189.800 494.000 190.400 ;
        RECT 495.600 189.800 498.000 190.400 ;
        RECT 492.400 189.600 493.200 189.800 ;
        RECT 486.000 188.200 486.800 188.400 ;
        RECT 489.000 188.300 491.600 188.400 ;
        RECT 494.000 188.300 494.800 189.200 ;
        RECT 486.000 187.600 487.600 188.200 ;
        RECT 489.000 187.700 494.800 188.300 ;
        RECT 489.000 187.600 491.600 187.700 ;
        RECT 494.000 187.600 494.800 187.700 ;
        RECT 486.800 187.200 487.600 187.600 ;
        RECT 484.400 184.800 485.200 186.400 ;
        RECT 486.200 186.200 489.800 186.600 ;
        RECT 490.800 186.200 491.400 187.600 ;
        RECT 495.600 186.200 496.200 189.800 ;
        RECT 497.200 189.600 498.000 189.800 ;
        RECT 502.000 189.800 503.400 190.400 ;
        RECT 506.400 189.800 507.200 190.000 ;
        RECT 502.000 189.600 503.800 189.800 ;
        RECT 502.800 189.200 503.800 189.600 ;
        RECT 498.800 187.600 500.400 188.400 ;
        RECT 501.600 187.600 502.400 188.400 ;
        RECT 501.800 187.200 502.400 187.600 ;
        RECT 500.400 186.800 501.200 187.000 ;
        RECT 486.000 186.000 490.000 186.200 ;
        RECT 486.000 182.200 486.800 186.000 ;
        RECT 489.200 182.200 490.000 186.000 ;
        RECT 490.800 182.200 491.600 186.200 ;
        RECT 495.600 182.200 496.400 186.200 ;
        RECT 497.200 185.600 498.000 186.400 ;
        RECT 498.800 186.200 501.200 186.800 ;
        RECT 501.800 186.400 502.600 187.200 ;
        RECT 497.000 184.800 497.800 185.600 ;
        RECT 498.800 182.200 499.600 186.200 ;
        RECT 503.200 185.800 503.800 189.200 ;
        RECT 504.600 189.200 507.200 189.800 ;
        RECT 504.600 188.600 505.200 189.200 ;
        RECT 504.400 187.800 505.200 188.600 ;
        RECT 507.600 188.200 509.200 188.400 ;
        RECT 505.800 187.600 509.200 188.200 ;
        RECT 505.800 187.200 506.400 187.600 ;
        RECT 504.400 186.600 506.400 187.200 ;
        RECT 507.000 186.800 507.800 187.000 ;
        RECT 504.400 186.400 506.000 186.600 ;
        RECT 507.000 186.200 509.200 186.800 ;
        RECT 503.200 182.200 504.800 185.800 ;
        RECT 508.400 182.200 509.200 186.200 ;
        RECT 510.000 184.800 510.800 186.400 ;
        RECT 511.600 182.200 512.400 199.800 ;
        RECT 515.800 192.600 516.600 199.800 ;
        RECT 514.800 191.800 516.600 192.600 ;
        RECT 515.000 188.400 515.600 191.800 ;
        RECT 518.000 191.600 518.800 193.200 ;
        RECT 516.400 189.600 517.200 191.200 ;
        RECT 514.800 187.600 515.600 188.400 ;
        RECT 513.200 184.800 514.000 186.400 ;
        RECT 515.000 184.400 515.600 187.600 ;
        RECT 519.600 186.200 520.400 199.800 ;
        RECT 524.400 190.300 525.200 199.800 ;
        RECT 529.200 194.300 530.000 199.800 ;
        RECT 532.400 194.300 533.200 194.400 ;
        RECT 529.200 193.700 533.200 194.300 ;
        RECT 527.600 191.600 528.400 193.200 ;
        RECT 527.700 190.300 528.300 191.600 ;
        RECT 524.400 189.700 528.300 190.300 ;
        RECT 521.200 186.800 522.000 188.400 ;
        RECT 518.600 185.600 520.400 186.200 ;
        RECT 518.600 184.400 519.400 185.600 ;
        RECT 514.800 182.200 515.600 184.400 ;
        RECT 518.000 183.600 519.400 184.400 ;
        RECT 518.600 182.200 519.400 183.600 ;
        RECT 524.400 182.200 525.200 189.700 ;
        RECT 526.000 188.300 526.800 188.400 ;
        RECT 527.600 188.300 528.400 188.400 ;
        RECT 526.000 187.700 528.400 188.300 ;
        RECT 526.000 186.800 526.800 187.700 ;
        RECT 527.600 187.600 528.400 187.700 ;
        RECT 529.200 186.200 530.000 193.700 ;
        RECT 532.400 193.600 533.200 193.700 ;
        RECT 530.800 186.800 531.600 188.400 ;
        RECT 528.200 185.600 530.000 186.200 ;
        RECT 528.200 182.200 529.000 185.600 ;
        RECT 532.400 184.800 533.200 186.400 ;
        RECT 534.000 182.200 534.800 199.800 ;
        RECT 535.600 186.800 536.400 188.400 ;
        RECT 537.200 186.200 538.000 199.800 ;
        RECT 538.800 191.600 539.600 193.200 ;
        RECT 537.200 185.600 539.000 186.200 ;
        RECT 538.200 182.200 539.000 185.600 ;
        RECT 540.400 182.200 541.200 199.800 ;
        RECT 546.200 192.400 547.000 199.800 ;
        RECT 547.600 193.600 548.400 194.400 ;
        RECT 547.800 192.400 548.400 193.600 ;
        RECT 550.600 192.600 551.400 199.800 ;
        RECT 546.200 191.800 547.200 192.400 ;
        RECT 547.800 191.800 549.200 192.400 ;
        RECT 550.600 191.800 552.400 192.600 ;
        RECT 554.800 192.400 555.600 199.800 ;
        RECT 556.400 192.400 557.200 192.600 ;
        RECT 559.200 192.400 560.800 199.800 ;
        RECT 554.800 191.800 557.200 192.400 ;
        RECT 558.800 191.800 560.800 192.400 ;
        RECT 563.000 192.400 563.800 192.600 ;
        RECT 564.400 192.400 565.200 199.800 ;
        RECT 563.000 191.800 565.200 192.400 ;
        RECT 545.200 188.800 546.000 190.400 ;
        RECT 546.600 188.400 547.200 191.800 ;
        RECT 548.400 191.600 549.200 191.800 ;
        RECT 550.000 189.600 550.800 191.200 ;
        RECT 551.600 188.400 552.200 191.800 ;
        RECT 558.800 190.400 559.400 191.800 ;
        RECT 563.000 191.200 563.600 191.800 ;
        RECT 560.200 190.600 563.600 191.200 ;
        RECT 566.000 191.400 566.800 199.800 ;
        RECT 570.400 196.400 571.200 199.800 ;
        RECT 569.200 195.800 571.200 196.400 ;
        RECT 574.800 195.800 575.600 199.800 ;
        RECT 579.000 195.800 580.200 199.800 ;
        RECT 569.200 195.000 570.000 195.800 ;
        RECT 574.800 195.200 575.400 195.800 ;
        RECT 572.600 194.600 576.200 195.200 ;
        RECT 578.800 195.000 579.600 195.800 ;
        RECT 572.600 194.400 573.400 194.600 ;
        RECT 575.400 194.400 576.200 194.600 ;
        RECT 569.200 193.000 570.000 193.200 ;
        RECT 573.800 193.000 574.600 193.200 ;
        RECT 569.200 192.400 574.600 193.000 ;
        RECT 575.200 193.000 577.400 193.600 ;
        RECT 575.200 191.800 575.800 193.000 ;
        RECT 576.600 192.800 577.400 193.000 ;
        RECT 579.000 193.200 580.400 194.000 ;
        RECT 579.000 192.200 579.600 193.200 ;
        RECT 571.000 191.400 575.800 191.800 ;
        RECT 566.000 191.200 575.800 191.400 ;
        RECT 577.200 191.600 579.600 192.200 ;
        RECT 566.000 191.000 571.800 191.200 ;
        RECT 566.000 190.800 571.600 191.000 ;
        RECT 560.200 190.400 561.000 190.600 ;
        RECT 558.000 189.800 559.400 190.400 ;
        RECT 572.400 190.200 573.200 190.400 ;
        RECT 562.400 189.800 563.200 190.000 ;
        RECT 558.000 189.600 559.800 189.800 ;
        RECT 558.800 189.200 559.800 189.600 ;
        RECT 542.000 188.300 542.800 188.400 ;
        RECT 543.600 188.300 544.400 188.400 ;
        RECT 542.000 188.200 544.400 188.300 ;
        RECT 542.000 187.700 545.200 188.200 ;
        RECT 542.000 186.800 542.800 187.700 ;
        RECT 543.600 187.600 545.200 187.700 ;
        RECT 546.600 187.600 549.200 188.400 ;
        RECT 551.600 188.300 552.400 188.400 ;
        RECT 554.800 188.300 556.400 188.400 ;
        RECT 551.600 187.700 556.400 188.300 ;
        RECT 551.600 187.600 552.400 187.700 ;
        RECT 554.800 187.600 556.400 187.700 ;
        RECT 557.600 187.600 558.400 188.400 ;
        RECT 544.400 187.200 545.200 187.600 ;
        RECT 543.800 186.200 547.400 186.600 ;
        RECT 548.400 186.200 549.000 187.600 ;
        RECT 543.600 186.000 547.600 186.200 ;
        RECT 543.600 182.200 544.400 186.000 ;
        RECT 546.800 182.200 547.600 186.000 ;
        RECT 548.400 182.200 549.200 186.200 ;
        RECT 551.600 184.200 552.200 187.600 ;
        RECT 557.800 187.200 558.400 187.600 ;
        RECT 556.400 186.800 557.200 187.000 ;
        RECT 553.200 184.800 554.000 186.400 ;
        RECT 554.800 186.200 557.200 186.800 ;
        RECT 557.800 186.400 558.600 187.200 ;
        RECT 551.600 182.200 552.400 184.200 ;
        RECT 554.800 182.200 555.600 186.200 ;
        RECT 559.200 185.800 559.800 189.200 ;
        RECT 560.600 189.200 563.200 189.800 ;
        RECT 568.200 189.600 573.200 190.200 ;
        RECT 568.200 189.400 569.000 189.600 ;
        RECT 570.800 189.400 571.600 189.600 ;
        RECT 560.600 188.600 561.200 189.200 ;
        RECT 560.400 187.800 561.200 188.600 ;
        RECT 569.800 188.400 570.600 188.600 ;
        RECT 577.200 188.400 577.800 191.600 ;
        RECT 583.600 191.200 584.400 199.800 ;
        RECT 580.200 190.600 584.400 191.200 ;
        RECT 580.200 190.400 581.000 190.600 ;
        RECT 581.800 189.800 582.600 190.000 ;
        RECT 578.800 189.200 582.600 189.800 ;
        RECT 578.800 189.000 579.600 189.200 ;
        RECT 563.600 188.200 565.200 188.400 ;
        RECT 561.800 187.600 565.200 188.200 ;
        RECT 566.800 187.800 577.800 188.400 ;
        RECT 566.800 187.600 568.400 187.800 ;
        RECT 561.800 187.200 562.400 187.600 ;
        RECT 560.400 186.600 562.400 187.200 ;
        RECT 563.000 186.800 563.800 187.000 ;
        RECT 560.400 186.400 562.000 186.600 ;
        RECT 563.000 186.200 565.200 186.800 ;
        RECT 559.200 182.200 560.800 185.800 ;
        RECT 564.400 182.200 565.200 186.200 ;
        RECT 566.000 182.200 566.800 187.000 ;
        RECT 571.000 185.600 571.600 187.800 ;
        RECT 576.600 187.600 577.400 187.800 ;
        RECT 583.600 187.200 584.400 190.600 ;
        RECT 580.600 186.600 584.400 187.200 ;
        RECT 580.600 186.400 581.400 186.600 ;
        RECT 569.200 184.200 570.000 185.000 ;
        RECT 570.800 184.800 571.600 185.600 ;
        RECT 572.600 185.400 573.400 185.600 ;
        RECT 572.600 184.800 575.400 185.400 ;
        RECT 574.800 184.200 575.400 184.800 ;
        RECT 578.800 184.200 579.600 185.000 ;
        RECT 569.200 183.600 571.200 184.200 ;
        RECT 570.400 182.200 571.200 183.600 ;
        RECT 574.800 182.200 575.600 184.200 ;
        RECT 578.800 183.600 580.200 184.200 ;
        RECT 579.000 182.200 580.200 183.600 ;
        RECT 583.600 182.200 584.400 186.600 ;
        RECT 1.200 175.400 2.000 179.800 ;
        RECT 5.400 178.400 6.600 179.800 ;
        RECT 5.400 177.800 6.800 178.400 ;
        RECT 10.000 177.800 10.800 179.800 ;
        RECT 14.400 178.400 15.200 179.800 ;
        RECT 14.400 177.800 16.400 178.400 ;
        RECT 6.000 177.000 6.800 177.800 ;
        RECT 10.200 177.200 10.800 177.800 ;
        RECT 10.200 176.600 13.000 177.200 ;
        RECT 12.200 176.400 13.000 176.600 ;
        RECT 14.000 176.400 14.800 177.200 ;
        RECT 15.600 177.000 16.400 177.800 ;
        RECT 4.200 175.400 5.000 175.600 ;
        RECT 1.200 174.800 5.000 175.400 ;
        RECT 1.200 171.400 2.000 174.800 ;
        RECT 8.200 174.200 9.000 174.400 ;
        RECT 12.400 174.200 13.200 174.400 ;
        RECT 14.000 174.200 14.600 176.400 ;
        RECT 18.800 175.000 19.600 179.800 ;
        RECT 20.400 175.800 21.200 179.800 ;
        RECT 22.000 176.000 22.800 179.800 ;
        RECT 25.200 176.000 26.000 179.800 ;
        RECT 22.000 175.800 26.000 176.000 ;
        RECT 26.800 175.800 27.600 179.800 ;
        RECT 31.200 176.200 32.800 179.800 ;
        RECT 20.600 174.400 21.200 175.800 ;
        RECT 22.200 175.400 25.800 175.800 ;
        RECT 26.800 175.200 29.200 175.800 ;
        RECT 28.400 175.000 29.200 175.200 ;
        RECT 29.800 174.800 30.600 175.600 ;
        RECT 24.400 174.400 25.200 174.800 ;
        RECT 29.800 174.400 30.400 174.800 ;
        RECT 17.200 174.200 18.800 174.400 ;
        RECT 7.800 173.600 18.800 174.200 ;
        RECT 20.400 173.600 23.000 174.400 ;
        RECT 24.400 173.800 26.000 174.400 ;
        RECT 25.200 173.600 26.000 173.800 ;
        RECT 26.800 173.600 28.400 174.400 ;
        RECT 29.600 173.600 30.400 174.400 ;
        RECT 6.000 172.800 6.800 173.000 ;
        RECT 3.000 172.200 6.800 172.800 ;
        RECT 3.000 172.000 3.800 172.200 ;
        RECT 4.600 171.400 5.400 171.600 ;
        RECT 1.200 170.800 5.400 171.400 ;
        RECT 1.200 162.200 2.000 170.800 ;
        RECT 7.800 170.400 8.400 173.600 ;
        RECT 15.000 173.400 15.800 173.600 ;
        RECT 14.000 172.400 14.800 172.600 ;
        RECT 16.600 172.400 17.400 172.600 ;
        RECT 22.400 172.400 23.000 173.600 ;
        RECT 12.400 171.800 17.400 172.400 ;
        RECT 12.400 171.600 13.200 171.800 ;
        RECT 22.000 171.600 23.000 172.400 ;
        RECT 23.600 171.600 24.400 173.200 ;
        RECT 25.300 172.300 25.900 173.600 ;
        RECT 31.200 172.800 31.800 176.200 ;
        RECT 36.400 175.800 37.200 179.800 ;
        RECT 32.400 175.400 34.000 175.600 ;
        RECT 32.400 174.800 34.400 175.400 ;
        RECT 35.000 175.200 37.200 175.800 ;
        RECT 38.000 175.800 38.800 179.800 ;
        RECT 42.400 176.200 44.000 179.800 ;
        RECT 38.000 175.200 40.400 175.800 ;
        RECT 35.000 175.000 35.800 175.200 ;
        RECT 39.600 175.000 40.400 175.200 ;
        RECT 33.800 174.400 34.400 174.800 ;
        RECT 41.000 174.800 41.800 175.600 ;
        RECT 41.000 174.400 41.600 174.800 ;
        RECT 32.400 173.400 33.200 174.200 ;
        RECT 33.800 173.800 37.200 174.400 ;
        RECT 35.600 173.600 37.200 173.800 ;
        RECT 38.000 173.600 39.600 174.400 ;
        RECT 40.800 173.600 41.600 174.400 ;
        RECT 30.800 172.400 31.800 172.800 ;
        RECT 30.000 172.300 31.800 172.400 ;
        RECT 25.300 172.200 31.800 172.300 ;
        RECT 32.600 172.800 33.200 173.400 ;
        RECT 42.400 172.800 43.000 176.200 ;
        RECT 47.600 175.800 48.400 179.800 ;
        RECT 49.200 175.800 50.000 179.800 ;
        RECT 50.800 176.000 51.600 179.800 ;
        RECT 54.000 176.000 54.800 179.800 ;
        RECT 55.800 176.400 56.600 177.200 ;
        RECT 50.800 175.800 54.800 176.000 ;
        RECT 43.600 175.400 45.200 175.600 ;
        RECT 43.600 174.800 45.600 175.400 ;
        RECT 46.200 175.200 48.400 175.800 ;
        RECT 46.200 175.000 47.000 175.200 ;
        RECT 45.000 174.400 45.600 174.800 ;
        RECT 49.400 174.400 50.000 175.800 ;
        RECT 51.000 175.400 54.600 175.800 ;
        RECT 55.600 175.600 56.400 176.400 ;
        RECT 57.200 175.800 58.000 179.800 ;
        RECT 62.000 175.800 62.800 179.800 ;
        RECT 63.600 176.000 64.400 179.800 ;
        RECT 66.800 176.000 67.600 179.800 ;
        RECT 63.600 175.800 67.600 176.000 ;
        RECT 53.200 174.400 54.000 174.800 ;
        RECT 43.600 173.400 44.400 174.200 ;
        RECT 45.000 173.800 48.400 174.400 ;
        RECT 46.800 173.600 48.400 173.800 ;
        RECT 49.200 173.600 51.800 174.400 ;
        RECT 53.200 173.800 54.800 174.400 ;
        RECT 54.000 173.600 54.800 173.800 ;
        RECT 32.600 172.200 35.200 172.800 ;
        RECT 42.000 172.400 43.000 172.800 ;
        RECT 25.300 171.700 31.400 172.200 ;
        RECT 34.400 172.000 35.200 172.200 ;
        RECT 41.200 172.200 43.000 172.400 ;
        RECT 43.800 172.800 44.400 173.400 ;
        RECT 43.800 172.200 46.400 172.800 ;
        RECT 30.000 171.600 31.400 171.700 ;
        RECT 41.200 171.600 42.600 172.200 ;
        RECT 45.600 172.000 46.400 172.200 ;
        RECT 47.600 172.300 48.400 172.400 ;
        RECT 51.200 172.300 51.800 173.600 ;
        RECT 47.600 171.700 51.800 172.300 ;
        RECT 47.600 171.600 48.400 171.700 ;
        RECT 14.000 171.000 19.600 171.200 ;
        RECT 13.800 170.800 19.600 171.000 ;
        RECT 6.000 169.800 8.400 170.400 ;
        RECT 9.800 170.600 19.600 170.800 ;
        RECT 9.800 170.200 14.600 170.600 ;
        RECT 6.000 168.800 6.600 169.800 ;
        RECT 5.200 168.000 6.600 168.800 ;
        RECT 8.200 169.000 9.000 169.200 ;
        RECT 9.800 169.000 10.400 170.200 ;
        RECT 8.200 168.400 10.400 169.000 ;
        RECT 11.000 169.000 16.400 169.600 ;
        RECT 11.000 168.800 11.800 169.000 ;
        RECT 15.600 168.800 16.400 169.000 ;
        RECT 9.400 167.400 10.200 167.600 ;
        RECT 12.200 167.400 13.000 167.600 ;
        RECT 6.000 166.200 6.800 167.000 ;
        RECT 9.400 166.800 13.000 167.400 ;
        RECT 10.200 166.200 10.800 166.800 ;
        RECT 15.600 166.200 16.400 167.000 ;
        RECT 5.400 162.200 6.600 166.200 ;
        RECT 10.000 162.200 10.800 166.200 ;
        RECT 14.400 165.600 16.400 166.200 ;
        RECT 14.400 162.200 15.200 165.600 ;
        RECT 18.800 162.200 19.600 170.600 ;
        RECT 20.400 170.200 21.200 170.400 ;
        RECT 22.400 170.200 23.000 171.600 ;
        RECT 30.800 170.200 31.400 171.600 ;
        RECT 32.200 171.400 33.000 171.600 ;
        RECT 32.200 170.800 35.600 171.400 ;
        RECT 35.000 170.200 35.600 170.800 ;
        RECT 42.000 170.200 42.600 171.600 ;
        RECT 43.400 171.400 44.200 171.600 ;
        RECT 43.400 170.800 46.800 171.400 ;
        RECT 46.200 170.200 46.800 170.800 ;
        RECT 49.200 170.200 50.000 170.400 ;
        RECT 51.200 170.200 51.800 171.700 ;
        RECT 52.400 171.600 53.200 173.200 ;
        RECT 55.600 172.200 56.400 172.400 ;
        RECT 57.400 172.200 58.000 175.800 ;
        RECT 62.200 174.400 62.800 175.800 ;
        RECT 63.800 175.400 67.400 175.800 ;
        RECT 66.000 174.400 66.800 174.800 ;
        RECT 58.800 172.800 59.600 174.400 ;
        RECT 62.000 173.600 64.600 174.400 ;
        RECT 66.000 173.800 67.600 174.400 ;
        RECT 66.800 173.600 67.600 173.800 ;
        RECT 68.400 174.300 69.200 179.800 ;
        RECT 73.200 177.800 74.000 179.800 ;
        RECT 70.000 176.300 70.800 177.200 ;
        RECT 71.600 176.300 72.400 177.200 ;
        RECT 70.000 175.700 72.400 176.300 ;
        RECT 70.000 175.600 70.800 175.700 ;
        RECT 71.600 175.600 72.400 175.700 ;
        RECT 73.400 174.400 74.000 177.800 ;
        RECT 76.400 176.000 77.200 179.800 ;
        RECT 79.600 176.000 80.400 179.800 ;
        RECT 76.400 175.800 80.400 176.000 ;
        RECT 81.200 175.800 82.000 179.800 ;
        RECT 82.800 175.800 83.600 179.800 ;
        RECT 87.200 176.200 88.800 179.800 ;
        RECT 76.600 175.400 80.200 175.800 ;
        RECT 77.200 174.400 78.000 174.800 ;
        RECT 81.200 174.400 81.800 175.800 ;
        RECT 82.800 175.200 85.200 175.800 ;
        RECT 84.400 175.000 85.200 175.200 ;
        RECT 85.800 174.800 86.600 175.600 ;
        RECT 85.800 174.400 86.400 174.800 ;
        RECT 70.000 174.300 70.800 174.400 ;
        RECT 68.400 173.700 70.800 174.300 ;
        RECT 64.000 172.400 64.600 173.600 ;
        RECT 60.400 172.200 61.200 172.400 ;
        RECT 55.600 171.600 58.000 172.200 ;
        RECT 59.600 171.600 61.200 172.200 ;
        RECT 63.600 171.600 64.600 172.400 ;
        RECT 65.200 171.600 66.000 173.200 ;
        RECT 55.800 170.200 56.400 171.600 ;
        RECT 59.600 171.200 60.400 171.600 ;
        RECT 62.000 170.200 62.800 170.400 ;
        RECT 64.000 170.200 64.600 171.600 ;
        RECT 20.400 169.600 21.800 170.200 ;
        RECT 22.400 169.600 23.400 170.200 ;
        RECT 21.200 168.400 21.800 169.600 ;
        RECT 21.200 167.600 22.000 168.400 ;
        RECT 22.600 162.200 23.400 169.600 ;
        RECT 26.800 169.600 29.200 170.200 ;
        RECT 30.800 169.600 32.800 170.200 ;
        RECT 26.800 162.200 27.600 169.600 ;
        RECT 28.400 169.400 29.200 169.600 ;
        RECT 31.200 168.400 32.800 169.600 ;
        RECT 35.000 169.600 37.200 170.200 ;
        RECT 35.000 169.400 35.800 169.600 ;
        RECT 31.200 167.600 34.000 168.400 ;
        RECT 31.200 162.200 32.800 167.600 ;
        RECT 36.400 162.200 37.200 169.600 ;
        RECT 38.000 169.600 40.400 170.200 ;
        RECT 42.000 169.600 44.000 170.200 ;
        RECT 38.000 162.200 38.800 169.600 ;
        RECT 39.600 169.400 40.400 169.600 ;
        RECT 42.400 166.400 44.000 169.600 ;
        RECT 46.200 169.600 48.400 170.200 ;
        RECT 49.200 169.600 50.600 170.200 ;
        RECT 51.200 169.600 52.200 170.200 ;
        RECT 46.200 169.400 47.000 169.600 ;
        RECT 42.400 165.600 45.200 166.400 ;
        RECT 42.400 162.200 44.000 165.600 ;
        RECT 47.600 162.200 48.400 169.600 ;
        RECT 50.000 168.400 50.600 169.600 ;
        RECT 50.000 167.600 50.800 168.400 ;
        RECT 51.400 162.200 52.200 169.600 ;
        RECT 55.600 162.200 56.400 170.200 ;
        RECT 57.200 169.600 61.200 170.200 ;
        RECT 62.000 169.600 63.400 170.200 ;
        RECT 64.000 169.600 65.000 170.200 ;
        RECT 57.200 162.200 58.000 169.600 ;
        RECT 60.400 162.200 61.200 169.600 ;
        RECT 62.800 168.400 63.400 169.600 ;
        RECT 62.800 167.600 63.600 168.400 ;
        RECT 64.200 162.200 65.000 169.600 ;
        RECT 68.400 162.200 69.200 173.700 ;
        RECT 70.000 173.600 70.800 173.700 ;
        RECT 73.200 174.300 74.000 174.400 ;
        RECT 76.400 174.300 78.000 174.400 ;
        RECT 73.200 173.800 78.000 174.300 ;
        RECT 73.200 173.700 77.200 173.800 ;
        RECT 73.200 173.600 74.000 173.700 ;
        RECT 76.400 173.600 77.200 173.700 ;
        RECT 79.400 173.600 82.000 174.400 ;
        RECT 82.800 173.600 84.400 174.400 ;
        RECT 85.600 173.600 86.400 174.400 ;
        RECT 87.200 174.200 87.800 176.200 ;
        RECT 92.400 175.800 93.200 179.800 ;
        RECT 88.400 174.800 90.000 175.600 ;
        RECT 90.600 175.200 93.200 175.800 ;
        RECT 94.000 175.800 94.800 179.800 ;
        RECT 98.400 176.200 100.000 179.800 ;
        RECT 94.000 175.200 96.600 175.800 ;
        RECT 90.600 175.000 91.400 175.200 ;
        RECT 95.800 175.000 96.600 175.200 ;
        RECT 97.200 174.800 98.800 175.600 ;
        RECT 91.600 174.200 93.200 174.400 ;
        RECT 87.200 173.600 88.200 174.200 ;
        RECT 91.000 174.000 93.200 174.200 ;
        RECT 70.000 172.300 70.800 172.400 ;
        RECT 73.400 172.300 74.000 173.600 ;
        RECT 70.000 171.700 74.000 172.300 ;
        RECT 70.000 171.600 70.800 171.700 ;
        RECT 73.400 170.200 74.000 171.700 ;
        RECT 74.800 170.800 75.600 172.400 ;
        RECT 76.400 172.300 77.200 172.400 ;
        RECT 78.000 172.300 78.800 173.200 ;
        RECT 76.400 171.700 78.800 172.300 ;
        RECT 76.400 171.600 77.200 171.700 ;
        RECT 78.000 171.600 78.800 171.700 ;
        RECT 79.400 170.200 80.000 173.600 ;
        RECT 87.600 172.400 88.200 173.600 ;
        RECT 88.800 173.600 93.200 174.000 ;
        RECT 94.000 174.200 95.600 174.400 ;
        RECT 99.400 174.200 100.000 176.200 ;
        RECT 103.600 175.800 104.400 179.800 ;
        RECT 100.600 174.800 101.400 175.600 ;
        RECT 102.000 175.200 104.400 175.800 ;
        RECT 102.000 175.000 102.800 175.200 ;
        RECT 105.200 175.000 106.000 179.800 ;
        RECT 109.600 178.400 110.400 179.800 ;
        RECT 108.400 177.800 110.400 178.400 ;
        RECT 114.000 177.800 114.800 179.800 ;
        RECT 118.200 178.400 119.400 179.800 ;
        RECT 118.000 177.800 119.400 178.400 ;
        RECT 108.400 177.000 109.200 177.800 ;
        RECT 114.000 177.200 114.600 177.800 ;
        RECT 110.000 176.400 110.800 177.200 ;
        RECT 111.800 176.600 114.600 177.200 ;
        RECT 118.000 177.000 118.800 177.800 ;
        RECT 111.800 176.400 112.600 176.600 ;
        RECT 94.000 174.000 96.200 174.200 ;
        RECT 94.000 173.600 98.400 174.000 ;
        RECT 88.800 173.400 91.600 173.600 ;
        RECT 95.600 173.400 98.400 173.600 ;
        RECT 88.800 173.200 89.600 173.400 ;
        RECT 97.600 173.200 98.400 173.400 ;
        RECT 99.000 173.600 100.000 174.200 ;
        RECT 100.800 174.400 101.400 174.800 ;
        RECT 100.800 173.600 101.600 174.400 ;
        RECT 102.800 173.600 104.400 174.400 ;
        RECT 106.000 174.200 107.600 174.400 ;
        RECT 110.200 174.200 110.800 176.400 ;
        RECT 119.800 175.400 120.600 175.600 ;
        RECT 122.800 175.400 123.600 179.800 ;
        RECT 127.000 176.400 127.800 179.800 ;
        RECT 119.800 174.800 123.600 175.400 ;
        RECT 126.000 175.800 127.800 176.400 ;
        RECT 115.800 174.200 116.600 174.400 ;
        RECT 106.000 173.600 117.000 174.200 ;
        RECT 99.000 172.400 99.600 173.600 ;
        RECT 109.000 173.400 109.800 173.600 ;
        RECT 87.600 171.600 88.400 172.400 ;
        RECT 90.200 172.200 91.000 172.400 ;
        RECT 89.400 171.600 91.000 172.200 ;
        RECT 96.200 172.200 97.000 172.400 ;
        RECT 96.200 171.600 97.800 172.200 ;
        RECT 98.800 171.600 99.600 172.400 ;
        RECT 107.400 172.400 108.200 172.600 ;
        RECT 110.000 172.400 110.800 172.600 ;
        RECT 107.400 171.800 112.400 172.400 ;
        RECT 111.600 171.600 112.400 171.800 ;
        RECT 81.200 170.200 82.000 170.400 ;
        RECT 87.600 170.200 88.200 171.600 ;
        RECT 89.400 171.400 90.200 171.600 ;
        RECT 97.000 171.400 97.800 171.600 ;
        RECT 99.000 170.200 99.600 171.600 ;
        RECT 105.200 171.000 110.800 171.200 ;
        RECT 105.200 170.800 111.000 171.000 ;
        RECT 105.200 170.600 115.000 170.800 ;
        RECT 73.200 169.400 75.000 170.200 ;
        RECT 74.200 162.200 75.000 169.400 ;
        RECT 79.000 169.600 80.000 170.200 ;
        RECT 80.600 169.600 82.000 170.200 ;
        RECT 82.800 169.600 85.200 170.200 ;
        RECT 79.000 168.400 79.800 169.600 ;
        RECT 80.600 168.400 81.200 169.600 ;
        RECT 78.000 167.600 79.800 168.400 ;
        RECT 80.400 167.600 81.200 168.400 ;
        RECT 79.000 162.200 79.800 167.600 ;
        RECT 82.800 162.200 83.600 169.600 ;
        RECT 84.400 169.400 85.200 169.600 ;
        RECT 87.200 162.200 88.800 170.200 ;
        RECT 90.600 169.600 93.200 170.200 ;
        RECT 90.600 169.400 91.400 169.600 ;
        RECT 92.400 162.200 93.200 169.600 ;
        RECT 94.000 169.600 96.600 170.200 ;
        RECT 94.000 162.200 94.800 169.600 ;
        RECT 95.800 169.400 96.600 169.600 ;
        RECT 98.400 164.400 100.000 170.200 ;
        RECT 102.000 169.600 104.400 170.200 ;
        RECT 102.000 169.400 102.800 169.600 ;
        RECT 98.400 163.600 101.200 164.400 ;
        RECT 98.400 162.200 100.000 163.600 ;
        RECT 103.600 162.200 104.400 169.600 ;
        RECT 105.200 162.200 106.000 170.600 ;
        RECT 110.200 170.200 115.000 170.600 ;
        RECT 108.400 169.000 113.800 169.600 ;
        RECT 108.400 168.800 109.200 169.000 ;
        RECT 113.000 168.800 113.800 169.000 ;
        RECT 114.400 169.000 115.000 170.200 ;
        RECT 116.400 170.400 117.000 173.600 ;
        RECT 118.000 172.800 118.800 173.000 ;
        RECT 118.000 172.200 121.800 172.800 ;
        RECT 121.000 172.000 121.800 172.200 ;
        RECT 119.400 171.400 120.200 171.600 ;
        RECT 122.800 171.400 123.600 174.800 ;
        RECT 124.400 173.600 125.200 175.200 ;
        RECT 119.400 170.800 123.600 171.400 ;
        RECT 116.400 169.800 118.800 170.400 ;
        RECT 115.800 169.000 116.600 169.200 ;
        RECT 114.400 168.400 116.600 169.000 ;
        RECT 118.200 168.800 118.800 169.800 ;
        RECT 118.200 168.000 119.600 168.800 ;
        RECT 111.800 167.400 112.600 167.600 ;
        RECT 114.600 167.400 115.400 167.600 ;
        RECT 108.400 166.200 109.200 167.000 ;
        RECT 111.800 166.800 115.400 167.400 ;
        RECT 114.000 166.200 114.600 166.800 ;
        RECT 118.000 166.200 118.800 167.000 ;
        RECT 108.400 165.600 110.400 166.200 ;
        RECT 109.600 162.200 110.400 165.600 ;
        RECT 114.000 162.200 114.800 166.200 ;
        RECT 118.200 162.200 119.400 166.200 ;
        RECT 122.800 162.200 123.600 170.800 ;
        RECT 126.000 172.300 126.800 175.800 ;
        RECT 134.000 175.000 134.800 179.800 ;
        RECT 138.400 178.400 139.200 179.800 ;
        RECT 137.200 177.800 139.200 178.400 ;
        RECT 142.800 177.800 143.600 179.800 ;
        RECT 147.000 178.400 148.200 179.800 ;
        RECT 146.800 177.800 148.200 178.400 ;
        RECT 137.200 177.000 138.000 177.800 ;
        RECT 142.800 177.200 143.400 177.800 ;
        RECT 138.800 176.400 139.600 177.200 ;
        RECT 140.600 176.600 143.400 177.200 ;
        RECT 146.800 177.000 147.600 177.800 ;
        RECT 140.600 176.400 141.400 176.600 ;
        RECT 134.800 174.200 136.400 174.400 ;
        RECT 139.000 174.200 139.600 176.400 ;
        RECT 148.600 175.400 149.400 175.600 ;
        RECT 151.600 175.400 152.400 179.800 ;
        RECT 148.600 174.800 152.400 175.400 ;
        RECT 153.200 175.000 154.000 179.800 ;
        RECT 157.600 178.400 158.400 179.800 ;
        RECT 156.400 177.800 158.400 178.400 ;
        RECT 162.000 177.800 162.800 179.800 ;
        RECT 166.200 178.400 167.400 179.800 ;
        RECT 166.000 177.800 167.400 178.400 ;
        RECT 156.400 177.000 157.200 177.800 ;
        RECT 162.000 177.200 162.600 177.800 ;
        RECT 158.000 176.400 158.800 177.200 ;
        RECT 159.800 176.600 162.600 177.200 ;
        RECT 166.000 177.000 166.800 177.800 ;
        RECT 159.800 176.400 160.600 176.600 ;
        RECT 144.600 174.200 145.400 174.400 ;
        RECT 134.800 173.600 145.800 174.200 ;
        RECT 137.800 173.400 138.600 173.600 ;
        RECT 136.200 172.400 137.000 172.600 ;
        RECT 138.800 172.400 139.600 172.600 ;
        RECT 145.200 172.400 145.800 173.600 ;
        RECT 146.800 172.800 147.600 173.000 ;
        RECT 132.400 172.300 133.200 172.400 ;
        RECT 126.000 171.700 133.200 172.300 ;
        RECT 136.200 171.800 141.200 172.400 ;
        RECT 126.000 162.200 126.800 171.700 ;
        RECT 132.400 171.600 133.200 171.700 ;
        RECT 140.400 171.600 141.200 171.800 ;
        RECT 145.200 171.600 146.000 172.400 ;
        RECT 146.800 172.200 150.600 172.800 ;
        RECT 149.800 172.000 150.600 172.200 ;
        RECT 134.000 171.000 139.600 171.200 ;
        RECT 134.000 170.800 139.800 171.000 ;
        RECT 134.000 170.600 143.800 170.800 ;
        RECT 127.600 168.800 128.400 170.400 ;
        RECT 134.000 162.200 134.800 170.600 ;
        RECT 139.000 170.200 143.800 170.600 ;
        RECT 137.200 169.000 142.600 169.600 ;
        RECT 137.200 168.800 138.000 169.000 ;
        RECT 141.800 168.800 142.600 169.000 ;
        RECT 143.200 169.000 143.800 170.200 ;
        RECT 145.200 170.400 145.800 171.600 ;
        RECT 148.200 171.400 149.000 171.600 ;
        RECT 151.600 171.400 152.400 174.800 ;
        RECT 154.000 174.200 155.600 174.400 ;
        RECT 158.200 174.200 158.800 176.400 ;
        RECT 167.800 175.400 168.600 175.600 ;
        RECT 170.800 175.400 171.600 179.800 ;
        RECT 167.800 174.800 171.600 175.400 ;
        RECT 172.400 175.800 173.200 179.800 ;
        RECT 176.800 176.200 178.400 179.800 ;
        RECT 172.400 175.200 174.800 175.800 ;
        RECT 174.000 175.000 174.800 175.200 ;
        RECT 163.800 174.200 164.600 174.400 ;
        RECT 154.000 173.600 165.000 174.200 ;
        RECT 157.000 173.400 157.800 173.600 ;
        RECT 155.400 172.400 156.200 172.600 ;
        RECT 158.000 172.400 158.800 172.600 ;
        RECT 164.400 172.400 165.000 173.600 ;
        RECT 166.000 172.800 166.800 173.000 ;
        RECT 155.400 171.800 160.400 172.400 ;
        RECT 159.600 171.600 160.400 171.800 ;
        RECT 164.400 171.600 165.200 172.400 ;
        RECT 166.000 172.200 169.800 172.800 ;
        RECT 169.000 172.000 169.800 172.200 ;
        RECT 148.200 170.800 152.400 171.400 ;
        RECT 145.200 169.800 147.600 170.400 ;
        RECT 144.600 169.000 145.400 169.200 ;
        RECT 143.200 168.400 145.400 169.000 ;
        RECT 147.000 168.800 147.600 169.800 ;
        RECT 147.000 168.000 148.400 168.800 ;
        RECT 140.600 167.400 141.400 167.600 ;
        RECT 143.400 167.400 144.200 167.600 ;
        RECT 137.200 166.200 138.000 167.000 ;
        RECT 140.600 166.800 144.200 167.400 ;
        RECT 142.800 166.200 143.400 166.800 ;
        RECT 146.800 166.200 147.600 167.000 ;
        RECT 137.200 165.600 139.200 166.200 ;
        RECT 138.400 162.200 139.200 165.600 ;
        RECT 142.800 162.200 143.600 166.200 ;
        RECT 147.000 162.200 148.200 166.200 ;
        RECT 151.600 162.200 152.400 170.800 ;
        RECT 153.200 171.000 158.800 171.200 ;
        RECT 153.200 170.800 159.000 171.000 ;
        RECT 153.200 170.600 163.000 170.800 ;
        RECT 153.200 162.200 154.000 170.600 ;
        RECT 158.200 170.200 163.000 170.600 ;
        RECT 156.400 169.000 161.800 169.600 ;
        RECT 156.400 168.800 157.200 169.000 ;
        RECT 161.000 168.800 161.800 169.000 ;
        RECT 162.400 169.000 163.000 170.200 ;
        RECT 164.400 170.400 165.000 171.600 ;
        RECT 167.400 171.400 168.200 171.600 ;
        RECT 170.800 171.400 171.600 174.800 ;
        RECT 175.400 174.800 176.200 175.600 ;
        RECT 175.400 174.400 176.000 174.800 ;
        RECT 172.400 173.600 174.000 174.400 ;
        RECT 175.200 173.600 176.000 174.400 ;
        RECT 176.800 172.800 177.400 176.200 ;
        RECT 182.000 175.800 182.800 179.800 ;
        RECT 183.600 176.000 184.400 179.800 ;
        RECT 186.800 176.000 187.600 179.800 ;
        RECT 183.600 175.800 187.600 176.000 ;
        RECT 188.400 175.800 189.200 179.800 ;
        RECT 192.600 176.400 193.400 179.800 ;
        RECT 191.600 175.800 193.400 176.400 ;
        RECT 194.800 176.000 195.600 179.800 ;
        RECT 198.000 176.000 198.800 179.800 ;
        RECT 194.800 175.800 198.800 176.000 ;
        RECT 199.600 175.800 200.400 179.800 ;
        RECT 201.400 176.400 202.200 177.200 ;
        RECT 178.000 175.400 179.600 175.600 ;
        RECT 178.000 174.800 180.000 175.400 ;
        RECT 180.600 175.200 182.800 175.800 ;
        RECT 183.800 175.400 187.400 175.800 ;
        RECT 180.600 175.000 181.400 175.200 ;
        RECT 179.400 174.400 180.000 174.800 ;
        RECT 184.400 174.400 185.200 174.800 ;
        RECT 188.400 174.400 189.000 175.800 ;
        RECT 178.000 173.400 178.800 174.200 ;
        RECT 179.400 173.800 182.800 174.400 ;
        RECT 181.200 173.600 182.800 173.800 ;
        RECT 183.600 173.800 185.200 174.400 ;
        RECT 183.600 173.600 184.400 173.800 ;
        RECT 186.600 173.600 189.200 174.400 ;
        RECT 190.000 173.600 190.800 175.200 ;
        RECT 176.400 172.400 177.400 172.800 ;
        RECT 175.600 172.200 177.400 172.400 ;
        RECT 178.200 172.800 178.800 173.400 ;
        RECT 178.200 172.200 180.800 172.800 ;
        RECT 175.600 171.600 177.000 172.200 ;
        RECT 180.000 172.000 180.800 172.200 ;
        RECT 185.200 171.600 186.000 173.200 ;
        RECT 186.600 172.400 187.200 173.600 ;
        RECT 186.600 171.600 187.600 172.400 ;
        RECT 167.400 170.800 171.600 171.400 ;
        RECT 164.400 169.800 166.800 170.400 ;
        RECT 163.800 169.000 164.600 169.200 ;
        RECT 162.400 168.400 164.600 169.000 ;
        RECT 166.200 168.800 166.800 169.800 ;
        RECT 166.200 168.000 167.600 168.800 ;
        RECT 159.800 167.400 160.600 167.600 ;
        RECT 162.600 167.400 163.400 167.600 ;
        RECT 156.400 166.200 157.200 167.000 ;
        RECT 159.800 166.800 163.400 167.400 ;
        RECT 162.000 166.200 162.600 166.800 ;
        RECT 166.000 166.200 166.800 167.000 ;
        RECT 156.400 165.600 158.400 166.200 ;
        RECT 157.600 162.200 158.400 165.600 ;
        RECT 162.000 162.200 162.800 166.200 ;
        RECT 166.200 162.200 167.400 166.200 ;
        RECT 170.800 162.200 171.600 170.800 ;
        RECT 176.400 170.200 177.000 171.600 ;
        RECT 177.800 171.400 178.600 171.600 ;
        RECT 177.800 170.800 181.200 171.400 ;
        RECT 180.600 170.200 181.200 170.800 ;
        RECT 186.600 170.200 187.200 171.600 ;
        RECT 188.400 170.300 189.200 170.400 ;
        RECT 191.600 170.300 192.400 175.800 ;
        RECT 195.000 175.400 198.600 175.800 ;
        RECT 195.600 174.400 196.400 174.800 ;
        RECT 199.600 174.400 200.200 175.800 ;
        RECT 201.200 175.600 202.000 176.400 ;
        RECT 202.800 175.800 203.600 179.800 ;
        RECT 193.200 174.300 194.000 174.400 ;
        RECT 194.800 174.300 196.400 174.400 ;
        RECT 193.200 173.800 196.400 174.300 ;
        RECT 193.200 173.700 195.600 173.800 ;
        RECT 193.200 173.600 194.000 173.700 ;
        RECT 194.800 173.600 195.600 173.700 ;
        RECT 197.800 173.600 200.400 174.400 ;
        RECT 196.400 172.300 197.200 173.200 ;
        RECT 193.300 171.700 197.200 172.300 ;
        RECT 193.300 170.400 193.900 171.700 ;
        RECT 196.400 171.600 197.200 171.700 ;
        RECT 197.800 172.400 198.400 173.600 ;
        RECT 203.000 172.400 203.600 175.800 ;
        RECT 204.400 172.800 205.200 174.400 ;
        RECT 197.800 171.600 198.800 172.400 ;
        RECT 201.200 172.200 202.000 172.400 ;
        RECT 202.800 172.200 203.600 172.400 ;
        RECT 206.000 172.300 206.800 172.400 ;
        RECT 207.600 172.300 208.400 179.800 ;
        RECT 209.200 175.600 210.000 177.200 ;
        RECT 210.800 176.000 211.600 179.800 ;
        RECT 214.000 176.000 214.800 179.800 ;
        RECT 210.800 175.800 214.800 176.000 ;
        RECT 215.600 175.800 216.400 179.800 ;
        RECT 217.200 175.800 218.000 179.800 ;
        RECT 218.800 176.000 219.600 179.800 ;
        RECT 222.000 176.000 222.800 179.800 ;
        RECT 226.200 176.400 227.000 179.800 ;
        RECT 231.000 176.400 231.800 179.800 ;
        RECT 218.800 175.800 222.800 176.000 ;
        RECT 225.200 175.800 227.000 176.400 ;
        RECT 230.000 175.800 231.800 176.400 ;
        RECT 211.000 175.400 214.600 175.800 ;
        RECT 211.600 174.400 212.400 174.800 ;
        RECT 215.600 174.400 216.200 175.800 ;
        RECT 217.400 174.400 218.000 175.800 ;
        RECT 219.000 175.400 222.600 175.800 ;
        RECT 221.200 174.400 222.000 174.800 ;
        RECT 210.800 173.800 212.400 174.400 ;
        RECT 210.800 173.600 211.600 173.800 ;
        RECT 213.800 173.600 216.400 174.400 ;
        RECT 217.200 173.600 219.800 174.400 ;
        RECT 221.200 173.800 222.800 174.400 ;
        RECT 222.000 173.600 222.800 173.800 ;
        RECT 223.600 173.600 224.400 175.200 ;
        RECT 225.200 174.300 226.000 175.800 ;
        RECT 228.400 174.300 229.200 175.200 ;
        RECT 225.200 173.700 229.200 174.300 ;
        RECT 206.000 172.200 208.400 172.300 ;
        RECT 201.200 171.600 203.600 172.200 ;
        RECT 205.200 171.700 208.400 172.200 ;
        RECT 205.200 171.600 206.800 171.700 ;
        RECT 188.400 170.200 192.400 170.300 ;
        RECT 172.400 169.600 174.800 170.200 ;
        RECT 176.400 169.600 178.400 170.200 ;
        RECT 172.400 162.200 173.200 169.600 ;
        RECT 174.000 169.400 174.800 169.600 ;
        RECT 176.800 166.400 178.400 169.600 ;
        RECT 180.600 169.600 182.800 170.200 ;
        RECT 180.600 169.400 181.400 169.600 ;
        RECT 176.800 165.600 179.600 166.400 ;
        RECT 176.800 162.200 178.400 165.600 ;
        RECT 182.000 162.200 182.800 169.600 ;
        RECT 186.200 169.600 187.200 170.200 ;
        RECT 187.800 169.700 192.400 170.200 ;
        RECT 187.800 169.600 189.200 169.700 ;
        RECT 186.200 162.200 187.000 169.600 ;
        RECT 187.800 168.400 188.400 169.600 ;
        RECT 187.600 167.600 188.400 168.400 ;
        RECT 191.600 162.200 192.400 169.700 ;
        RECT 193.200 168.800 194.000 170.400 ;
        RECT 197.800 170.200 198.400 171.600 ;
        RECT 199.600 170.200 200.400 170.400 ;
        RECT 201.400 170.200 202.000 171.600 ;
        RECT 205.200 171.200 206.000 171.600 ;
        RECT 197.400 169.600 198.400 170.200 ;
        RECT 199.000 169.600 200.400 170.200 ;
        RECT 197.400 162.200 198.200 169.600 ;
        RECT 199.000 168.400 199.600 169.600 ;
        RECT 198.800 167.600 199.600 168.400 ;
        RECT 201.200 162.200 202.000 170.200 ;
        RECT 202.800 169.600 206.800 170.200 ;
        RECT 202.800 162.200 203.600 169.600 ;
        RECT 206.000 162.200 206.800 169.600 ;
        RECT 207.600 162.200 208.400 171.700 ;
        RECT 212.400 171.600 213.200 173.200 ;
        RECT 213.800 172.300 214.400 173.600 ;
        RECT 215.600 172.300 216.400 172.400 ;
        RECT 213.800 171.700 216.400 172.300 ;
        RECT 213.800 170.200 214.400 171.700 ;
        RECT 215.600 171.600 216.400 171.700 ;
        RECT 215.600 170.200 216.400 170.400 ;
        RECT 213.400 169.600 214.400 170.200 ;
        RECT 215.000 169.600 216.400 170.200 ;
        RECT 217.200 170.200 218.000 170.400 ;
        RECT 219.200 170.200 219.800 173.600 ;
        RECT 220.400 171.600 221.200 173.200 ;
        RECT 217.200 169.600 218.600 170.200 ;
        RECT 219.200 169.600 220.200 170.200 ;
        RECT 213.400 162.200 214.200 169.600 ;
        RECT 215.000 168.400 215.600 169.600 ;
        RECT 214.800 167.600 215.600 168.400 ;
        RECT 218.000 168.400 218.600 169.600 ;
        RECT 219.400 168.400 220.200 169.600 ;
        RECT 218.000 167.600 218.800 168.400 ;
        RECT 219.400 167.600 221.200 168.400 ;
        RECT 219.400 162.200 220.200 167.600 ;
        RECT 225.200 162.200 226.000 173.700 ;
        RECT 228.400 173.600 229.200 173.700 ;
        RECT 226.800 168.800 227.600 170.400 ;
        RECT 230.000 162.200 230.800 175.800 ;
        RECT 233.200 175.000 234.000 179.800 ;
        RECT 237.600 178.400 238.400 179.800 ;
        RECT 236.400 177.800 238.400 178.400 ;
        RECT 242.000 177.800 242.800 179.800 ;
        RECT 246.200 178.400 247.400 179.800 ;
        RECT 246.000 177.800 247.400 178.400 ;
        RECT 236.400 177.000 237.200 177.800 ;
        RECT 242.000 177.200 242.600 177.800 ;
        RECT 238.000 176.400 238.800 177.200 ;
        RECT 239.800 176.600 242.600 177.200 ;
        RECT 246.000 177.000 246.800 177.800 ;
        RECT 239.800 176.400 240.600 176.600 ;
        RECT 234.000 174.200 235.600 174.400 ;
        RECT 238.200 174.200 238.800 176.400 ;
        RECT 247.800 175.400 248.600 175.600 ;
        RECT 250.800 175.400 251.600 179.800 ;
        RECT 247.800 174.800 251.600 175.400 ;
        RECT 243.800 174.200 244.600 174.400 ;
        RECT 234.000 173.600 245.000 174.200 ;
        RECT 249.200 173.600 250.000 174.800 ;
        RECT 237.000 173.400 237.800 173.600 ;
        RECT 235.400 172.400 236.200 172.600 ;
        RECT 238.000 172.400 238.800 172.600 ;
        RECT 235.400 171.800 240.400 172.400 ;
        RECT 239.600 171.600 240.400 171.800 ;
        RECT 233.200 171.000 238.800 171.200 ;
        RECT 233.200 170.800 239.000 171.000 ;
        RECT 233.200 170.600 243.000 170.800 ;
        RECT 231.600 168.800 232.400 170.400 ;
        RECT 233.200 162.200 234.000 170.600 ;
        RECT 238.200 170.200 243.000 170.600 ;
        RECT 236.400 169.000 241.800 169.600 ;
        RECT 236.400 168.800 237.200 169.000 ;
        RECT 241.000 168.800 241.800 169.000 ;
        RECT 242.400 169.000 243.000 170.200 ;
        RECT 244.400 170.400 245.000 173.600 ;
        RECT 246.000 172.800 246.800 173.000 ;
        RECT 246.000 172.200 249.800 172.800 ;
        RECT 249.000 172.000 249.800 172.200 ;
        RECT 247.400 171.400 248.200 171.600 ;
        RECT 250.800 171.400 251.600 174.800 ;
        RECT 254.000 175.200 254.800 179.800 ;
        RECT 257.200 175.200 258.000 179.800 ;
        RECT 260.400 175.200 261.200 179.800 ;
        RECT 263.600 175.200 264.400 179.800 ;
        RECT 254.000 174.400 255.800 175.200 ;
        RECT 257.200 174.400 259.400 175.200 ;
        RECT 260.400 174.400 262.600 175.200 ;
        RECT 263.600 174.400 266.000 175.200 ;
        RECT 266.800 175.000 267.600 179.800 ;
        RECT 271.200 178.400 272.000 179.800 ;
        RECT 270.000 177.800 272.000 178.400 ;
        RECT 275.600 177.800 276.400 179.800 ;
        RECT 279.800 178.400 281.000 179.800 ;
        RECT 279.600 177.800 281.000 178.400 ;
        RECT 270.000 177.000 270.800 177.800 ;
        RECT 275.600 177.200 276.200 177.800 ;
        RECT 271.600 176.400 272.400 177.200 ;
        RECT 273.400 176.600 276.200 177.200 ;
        RECT 279.600 177.000 280.400 177.800 ;
        RECT 273.400 176.400 274.200 176.600 ;
        RECT 255.000 173.800 255.800 174.400 ;
        RECT 258.600 173.800 259.400 174.400 ;
        RECT 261.800 173.800 262.600 174.400 ;
        RECT 255.000 173.000 257.600 173.800 ;
        RECT 258.600 173.000 261.000 173.800 ;
        RECT 261.800 173.000 264.400 173.800 ;
        RECT 255.000 171.600 255.800 173.000 ;
        RECT 258.600 171.600 259.400 173.000 ;
        RECT 261.800 171.600 262.600 173.000 ;
        RECT 265.200 171.600 266.000 174.400 ;
        RECT 267.600 174.200 269.200 174.400 ;
        RECT 271.800 174.200 272.400 176.400 ;
        RECT 281.400 175.400 282.200 175.600 ;
        RECT 284.400 175.400 285.200 179.800 ;
        RECT 281.400 174.800 285.200 175.400 ;
        RECT 290.800 175.000 291.600 179.800 ;
        RECT 295.200 178.400 296.000 179.800 ;
        RECT 294.000 177.800 296.000 178.400 ;
        RECT 299.600 177.800 300.400 179.800 ;
        RECT 303.800 178.400 305.000 179.800 ;
        RECT 303.600 177.800 305.000 178.400 ;
        RECT 294.000 177.000 294.800 177.800 ;
        RECT 299.600 177.200 300.200 177.800 ;
        RECT 295.600 176.400 296.400 177.200 ;
        RECT 297.400 176.600 300.200 177.200 ;
        RECT 303.600 177.000 304.400 177.800 ;
        RECT 297.400 176.400 298.200 176.600 ;
        RECT 276.400 174.200 278.200 174.400 ;
        RECT 267.600 173.600 278.600 174.200 ;
        RECT 270.600 173.400 271.400 173.600 ;
        RECT 269.000 172.400 269.800 172.600 ;
        RECT 271.600 172.400 272.400 172.600 ;
        RECT 269.000 171.800 274.000 172.400 ;
        RECT 273.200 171.600 274.000 171.800 ;
        RECT 247.400 170.800 251.600 171.400 ;
        RECT 244.400 169.800 246.800 170.400 ;
        RECT 243.800 169.000 244.600 169.200 ;
        RECT 242.400 168.400 244.600 169.000 ;
        RECT 246.200 168.800 246.800 169.800 ;
        RECT 246.200 168.000 247.600 168.800 ;
        RECT 239.800 167.400 240.600 167.600 ;
        RECT 242.600 167.400 243.400 167.600 ;
        RECT 236.400 166.200 237.200 167.000 ;
        RECT 239.800 166.800 243.400 167.400 ;
        RECT 242.000 166.200 242.600 166.800 ;
        RECT 246.000 166.200 246.800 167.000 ;
        RECT 236.400 165.600 238.400 166.200 ;
        RECT 237.600 162.200 238.400 165.600 ;
        RECT 242.000 162.200 242.800 166.200 ;
        RECT 246.200 162.200 247.400 166.200 ;
        RECT 250.800 162.200 251.600 170.800 ;
        RECT 254.000 170.800 255.800 171.600 ;
        RECT 257.200 170.800 259.400 171.600 ;
        RECT 260.400 170.800 262.600 171.600 ;
        RECT 263.600 170.800 266.000 171.600 ;
        RECT 266.800 171.000 272.400 171.200 ;
        RECT 266.800 170.800 272.600 171.000 ;
        RECT 254.000 162.200 254.800 170.800 ;
        RECT 257.200 162.200 258.000 170.800 ;
        RECT 260.400 162.200 261.200 170.800 ;
        RECT 263.600 162.200 264.400 170.800 ;
        RECT 266.800 170.600 276.600 170.800 ;
        RECT 266.800 162.200 267.600 170.600 ;
        RECT 271.800 170.200 276.600 170.600 ;
        RECT 270.000 169.000 275.400 169.600 ;
        RECT 270.000 168.800 270.800 169.000 ;
        RECT 274.600 168.800 275.400 169.000 ;
        RECT 276.000 169.000 276.600 170.200 ;
        RECT 278.000 170.400 278.600 173.600 ;
        RECT 279.600 172.800 280.400 173.000 ;
        RECT 279.600 172.200 283.400 172.800 ;
        RECT 282.600 172.000 283.400 172.200 ;
        RECT 281.000 171.400 281.800 171.600 ;
        RECT 284.400 171.400 285.200 174.800 ;
        RECT 291.600 174.200 293.200 174.400 ;
        RECT 295.800 174.200 296.400 176.400 ;
        RECT 305.400 175.400 306.200 175.600 ;
        RECT 308.400 175.400 309.200 179.800 ;
        RECT 310.600 176.400 311.400 179.800 ;
        RECT 310.600 175.800 312.400 176.400 ;
        RECT 314.800 176.000 315.600 179.800 ;
        RECT 318.000 176.000 318.800 179.800 ;
        RECT 314.800 175.800 318.800 176.000 ;
        RECT 319.600 175.800 320.400 179.800 ;
        RECT 323.800 176.400 324.600 179.800 ;
        RECT 322.800 175.800 324.600 176.400 ;
        RECT 326.000 175.800 326.800 179.800 ;
        RECT 327.600 176.000 328.400 179.800 ;
        RECT 330.800 176.000 331.600 179.800 ;
        RECT 327.600 175.800 331.600 176.000 ;
        RECT 332.400 175.800 333.200 179.800 ;
        RECT 334.000 176.000 334.800 179.800 ;
        RECT 337.200 176.000 338.000 179.800 ;
        RECT 334.000 175.800 338.000 176.000 ;
        RECT 305.400 174.800 309.200 175.400 ;
        RECT 301.400 174.200 302.200 174.400 ;
        RECT 291.600 173.600 302.600 174.200 ;
        RECT 294.600 173.400 295.400 173.600 ;
        RECT 293.000 172.400 293.800 172.600 ;
        RECT 295.600 172.400 296.400 172.600 ;
        RECT 293.000 171.800 298.000 172.400 ;
        RECT 297.200 171.600 298.000 171.800 ;
        RECT 281.000 170.800 285.200 171.400 ;
        RECT 278.000 169.800 280.400 170.400 ;
        RECT 277.400 169.000 278.200 169.200 ;
        RECT 276.000 168.400 278.200 169.000 ;
        RECT 279.800 168.800 280.400 169.800 ;
        RECT 279.800 168.000 281.200 168.800 ;
        RECT 273.400 167.400 274.200 167.600 ;
        RECT 276.200 167.400 277.000 167.600 ;
        RECT 270.000 166.200 270.800 167.000 ;
        RECT 273.400 166.800 277.000 167.400 ;
        RECT 275.600 166.200 276.200 166.800 ;
        RECT 279.600 166.200 280.400 167.000 ;
        RECT 270.000 165.600 272.000 166.200 ;
        RECT 271.200 162.200 272.000 165.600 ;
        RECT 275.600 162.200 276.400 166.200 ;
        RECT 279.800 162.200 281.000 166.200 ;
        RECT 284.400 162.200 285.200 170.800 ;
        RECT 290.800 171.000 296.400 171.200 ;
        RECT 290.800 170.800 296.600 171.000 ;
        RECT 290.800 170.600 300.600 170.800 ;
        RECT 290.800 162.200 291.600 170.600 ;
        RECT 295.800 170.200 300.600 170.600 ;
        RECT 294.000 169.000 299.400 169.600 ;
        RECT 294.000 168.800 294.800 169.000 ;
        RECT 298.600 168.800 299.400 169.000 ;
        RECT 300.000 169.000 300.600 170.200 ;
        RECT 302.000 170.400 302.600 173.600 ;
        RECT 303.600 172.800 304.400 173.000 ;
        RECT 303.600 172.200 307.400 172.800 ;
        RECT 306.600 172.000 307.400 172.200 ;
        RECT 305.000 171.400 305.800 171.600 ;
        RECT 308.400 171.400 309.200 174.800 ;
        RECT 305.000 170.800 309.200 171.400 ;
        RECT 302.000 169.800 304.400 170.400 ;
        RECT 301.400 169.000 302.200 169.200 ;
        RECT 300.000 168.400 302.200 169.000 ;
        RECT 303.800 168.800 304.400 169.800 ;
        RECT 303.800 168.400 305.200 168.800 ;
        RECT 303.800 168.000 306.000 168.400 ;
        RECT 304.600 167.600 306.000 168.000 ;
        RECT 297.400 167.400 298.200 167.600 ;
        RECT 300.200 167.400 301.000 167.600 ;
        RECT 294.000 166.200 294.800 167.000 ;
        RECT 297.400 166.800 301.000 167.400 ;
        RECT 299.600 166.200 300.200 166.800 ;
        RECT 303.600 166.200 304.400 167.000 ;
        RECT 294.000 165.600 296.000 166.200 ;
        RECT 295.200 162.200 296.000 165.600 ;
        RECT 299.600 162.200 300.400 166.200 ;
        RECT 303.800 162.200 305.000 166.200 ;
        RECT 308.400 162.200 309.200 170.800 ;
        RECT 311.600 172.300 312.400 175.800 ;
        RECT 315.000 175.400 318.600 175.800 ;
        RECT 313.200 173.600 314.000 175.200 ;
        RECT 315.600 174.400 316.400 174.800 ;
        RECT 319.600 174.400 320.200 175.800 ;
        RECT 314.800 173.800 316.400 174.400 ;
        RECT 317.800 174.300 320.400 174.400 ;
        RECT 321.200 174.300 322.000 175.200 ;
        RECT 314.800 173.600 315.600 173.800 ;
        RECT 317.800 173.700 322.000 174.300 ;
        RECT 317.800 173.600 320.400 173.700 ;
        RECT 321.200 173.600 322.000 173.700 ;
        RECT 322.800 174.300 323.600 175.800 ;
        RECT 326.200 174.400 326.800 175.800 ;
        RECT 327.800 175.400 331.400 175.800 ;
        RECT 330.000 174.400 330.800 174.800 ;
        RECT 332.600 174.400 333.200 175.800 ;
        RECT 334.200 175.400 337.800 175.800 ;
        RECT 336.400 174.400 337.200 174.800 ;
        RECT 324.400 174.300 325.200 174.400 ;
        RECT 322.800 173.700 325.200 174.300 ;
        RECT 314.900 172.300 315.500 173.600 ;
        RECT 311.600 171.700 315.500 172.300 ;
        RECT 310.000 168.800 310.800 170.400 ;
        RECT 311.600 162.200 312.400 171.700 ;
        RECT 316.400 171.600 317.200 173.200 ;
        RECT 317.800 170.200 318.400 173.600 ;
        RECT 319.600 170.200 320.400 170.400 ;
        RECT 317.400 169.600 318.400 170.200 ;
        RECT 319.000 169.600 320.400 170.200 ;
        RECT 317.400 162.200 318.200 169.600 ;
        RECT 319.000 168.400 319.600 169.600 ;
        RECT 318.800 167.600 319.600 168.400 ;
        RECT 322.800 162.200 323.600 173.700 ;
        RECT 324.400 173.600 325.200 173.700 ;
        RECT 326.000 173.600 328.600 174.400 ;
        RECT 330.000 173.800 331.600 174.400 ;
        RECT 330.800 173.600 331.600 173.800 ;
        RECT 332.400 173.600 335.000 174.400 ;
        RECT 336.400 173.800 338.000 174.400 ;
        RECT 337.200 173.600 338.000 173.800 ;
        RECT 328.000 172.300 328.600 173.600 ;
        RECT 324.500 171.700 328.600 172.300 ;
        RECT 324.500 170.400 325.100 171.700 ;
        RECT 324.400 168.800 325.200 170.400 ;
        RECT 326.000 170.200 326.800 170.400 ;
        RECT 328.000 170.200 328.600 171.700 ;
        RECT 329.200 172.300 330.000 173.200 ;
        RECT 334.400 172.300 335.000 173.600 ;
        RECT 329.200 171.700 335.000 172.300 ;
        RECT 329.200 171.600 330.000 171.700 ;
        RECT 334.400 170.400 335.000 171.700 ;
        RECT 335.600 172.300 336.400 173.200 ;
        RECT 338.800 172.300 339.600 179.800 ;
        RECT 340.400 175.600 341.200 177.200 ;
        RECT 342.000 176.000 342.800 179.800 ;
        RECT 345.200 176.000 346.000 179.800 ;
        RECT 342.000 175.800 346.000 176.000 ;
        RECT 346.800 175.800 347.600 179.800 ;
        RECT 351.000 178.400 351.800 179.800 ;
        RECT 351.000 177.600 352.400 178.400 ;
        RECT 354.800 177.800 355.600 179.800 ;
        RECT 359.600 177.800 360.400 179.800 ;
        RECT 351.000 176.400 351.800 177.600 ;
        RECT 350.000 175.800 351.800 176.400 ;
        RECT 342.200 175.400 345.800 175.800 ;
        RECT 342.800 174.400 343.600 174.800 ;
        RECT 346.800 174.400 347.400 175.800 ;
        RECT 342.000 173.800 343.600 174.400 ;
        RECT 342.000 173.600 342.800 173.800 ;
        RECT 345.000 173.600 347.600 174.400 ;
        RECT 348.400 173.600 349.200 175.200 ;
        RECT 335.600 171.700 339.600 172.300 ;
        RECT 335.600 171.600 336.400 171.700 ;
        RECT 332.400 170.200 333.200 170.400 ;
        RECT 326.000 169.600 327.400 170.200 ;
        RECT 328.000 169.600 329.000 170.200 ;
        RECT 332.400 169.600 333.800 170.200 ;
        RECT 334.400 169.600 336.400 170.400 ;
        RECT 326.800 168.400 327.400 169.600 ;
        RECT 326.800 167.600 327.600 168.400 ;
        RECT 328.200 162.200 329.000 169.600 ;
        RECT 333.200 168.400 333.800 169.600 ;
        RECT 333.200 167.600 334.000 168.400 ;
        RECT 334.600 162.200 335.400 169.600 ;
        RECT 338.800 162.200 339.600 171.700 ;
        RECT 343.600 171.600 344.400 173.200 ;
        RECT 345.000 172.300 345.600 173.600 ;
        RECT 348.400 172.300 349.200 172.400 ;
        RECT 345.000 171.700 349.200 172.300 ;
        RECT 345.000 170.200 345.600 171.700 ;
        RECT 348.400 171.600 349.200 171.700 ;
        RECT 346.800 170.200 347.600 170.400 ;
        RECT 344.600 169.600 345.600 170.200 ;
        RECT 346.200 169.600 347.600 170.200 ;
        RECT 344.600 162.200 345.400 169.600 ;
        RECT 346.200 168.400 346.800 169.600 ;
        RECT 346.000 167.600 346.800 168.400 ;
        RECT 350.000 162.200 350.800 175.800 ;
        RECT 354.800 174.400 355.400 177.800 ;
        RECT 356.400 175.600 357.200 177.200 ;
        RECT 358.000 175.600 358.800 177.200 ;
        RECT 354.800 174.300 355.600 174.400 ;
        RECT 358.100 174.300 358.700 175.600 ;
        RECT 359.800 174.400 360.400 177.800 ;
        RECT 354.800 173.700 358.700 174.300 ;
        RECT 354.800 173.600 355.600 173.700 ;
        RECT 359.600 173.600 360.400 174.400 ;
        RECT 353.200 170.800 354.000 172.400 ;
        RECT 351.600 168.800 352.400 170.400 ;
        RECT 354.800 170.200 355.400 173.600 ;
        RECT 359.800 170.200 360.400 173.600 ;
        RECT 361.200 170.800 362.000 172.400 ;
        RECT 362.800 172.300 363.600 179.800 ;
        RECT 367.600 177.800 368.400 179.800 ;
        RECT 364.400 175.600 365.200 177.200 ;
        RECT 367.600 174.400 368.200 177.800 ;
        RECT 369.200 175.600 370.000 177.200 ;
        RECT 371.000 176.400 371.800 177.200 ;
        RECT 370.800 175.600 371.600 176.400 ;
        RECT 372.400 175.800 373.200 179.800 ;
        RECT 378.800 177.600 379.600 179.800 ;
        RECT 384.600 178.400 385.400 179.800 ;
        RECT 383.600 177.600 385.400 178.400 ;
        RECT 366.000 174.300 366.800 174.400 ;
        RECT 367.600 174.300 368.400 174.400 ;
        RECT 370.900 174.300 371.500 175.600 ;
        RECT 366.000 173.700 371.500 174.300 ;
        RECT 366.000 173.600 366.800 173.700 ;
        RECT 367.600 173.600 368.400 173.700 ;
        RECT 366.000 172.300 366.800 172.400 ;
        RECT 362.800 171.700 366.800 172.300 ;
        RECT 353.800 169.400 355.600 170.200 ;
        RECT 359.600 169.400 361.400 170.200 ;
        RECT 353.800 162.200 354.600 169.400 ;
        RECT 360.600 168.400 361.400 169.400 ;
        RECT 360.600 167.600 362.000 168.400 ;
        RECT 360.600 162.200 361.400 167.600 ;
        RECT 362.800 162.200 363.600 171.700 ;
        RECT 366.000 170.800 366.800 171.700 ;
        RECT 367.600 170.200 368.200 173.600 ;
        RECT 370.800 172.200 371.600 172.400 ;
        RECT 372.600 172.200 373.200 175.800 ;
        RECT 377.200 175.600 378.000 177.200 ;
        RECT 379.000 174.400 379.600 177.600 ;
        RECT 384.600 176.400 385.400 177.600 ;
        RECT 383.600 175.800 385.400 176.400 ;
        RECT 386.800 176.000 387.600 179.800 ;
        RECT 390.000 176.000 390.800 179.800 ;
        RECT 386.800 175.800 390.800 176.000 ;
        RECT 391.600 175.800 392.400 179.800 ;
        RECT 374.000 172.800 374.800 174.400 ;
        RECT 378.800 173.600 379.600 174.400 ;
        RECT 382.000 173.600 382.800 175.200 ;
        RECT 375.600 172.200 376.400 172.400 ;
        RECT 370.800 171.600 373.200 172.200 ;
        RECT 374.800 171.600 376.400 172.200 ;
        RECT 371.000 170.200 371.600 171.600 ;
        RECT 374.800 171.200 375.600 171.600 ;
        RECT 379.000 170.200 379.600 173.600 ;
        RECT 380.400 170.800 381.200 172.400 ;
        RECT 366.600 169.400 368.400 170.200 ;
        RECT 366.600 162.200 367.400 169.400 ;
        RECT 370.800 162.200 371.600 170.200 ;
        RECT 372.400 169.600 376.400 170.200 ;
        RECT 372.400 162.200 373.200 169.600 ;
        RECT 375.600 162.200 376.400 169.600 ;
        RECT 378.800 169.400 380.600 170.200 ;
        RECT 379.800 162.200 380.600 169.400 ;
        RECT 383.600 162.200 384.400 175.800 ;
        RECT 387.000 175.400 390.600 175.800 ;
        RECT 387.600 174.400 388.400 174.800 ;
        RECT 391.600 174.400 392.200 175.800 ;
        RECT 393.200 175.600 394.000 177.200 ;
        RECT 386.800 173.800 388.400 174.400 ;
        RECT 386.800 173.600 387.600 173.800 ;
        RECT 389.800 173.600 392.400 174.400 ;
        RECT 388.400 171.600 389.200 173.200 ;
        RECT 389.800 172.400 390.400 173.600 ;
        RECT 389.800 171.600 390.800 172.400 ;
        RECT 385.200 168.800 386.000 170.400 ;
        RECT 389.800 170.200 390.400 171.600 ;
        RECT 391.600 170.200 392.400 170.400 ;
        RECT 389.400 169.600 390.400 170.200 ;
        RECT 391.000 169.600 392.400 170.200 ;
        RECT 394.800 170.300 395.600 179.800 ;
        RECT 399.000 176.400 399.800 179.800 ;
        RECT 398.000 175.800 399.800 176.400 ;
        RECT 401.200 175.800 402.000 179.800 ;
        RECT 402.800 176.000 403.600 179.800 ;
        RECT 406.000 176.000 406.800 179.800 ;
        RECT 402.800 175.800 406.800 176.000 ;
        RECT 396.400 173.600 397.200 175.200 ;
        RECT 396.400 170.300 397.200 170.400 ;
        RECT 394.800 169.700 397.200 170.300 ;
        RECT 389.400 162.200 390.200 169.600 ;
        RECT 391.000 168.400 391.600 169.600 ;
        RECT 390.800 167.600 391.600 168.400 ;
        RECT 394.800 162.200 395.600 169.700 ;
        RECT 396.400 169.600 397.200 169.700 ;
        RECT 398.000 162.200 398.800 175.800 ;
        RECT 401.400 174.400 402.000 175.800 ;
        RECT 403.000 175.400 406.600 175.800 ;
        RECT 405.200 174.400 406.000 174.800 ;
        RECT 401.200 173.600 403.800 174.400 ;
        RECT 405.200 173.800 406.800 174.400 ;
        RECT 406.000 173.600 406.800 173.800 ;
        RECT 399.600 168.800 400.400 170.400 ;
        RECT 401.200 170.200 402.000 170.400 ;
        RECT 403.200 170.200 403.800 173.600 ;
        RECT 404.400 172.300 405.200 173.200 ;
        RECT 407.600 172.300 408.400 179.800 ;
        RECT 409.200 175.600 410.000 177.200 ;
        RECT 410.800 176.000 411.600 179.800 ;
        RECT 414.000 176.000 414.800 179.800 ;
        RECT 410.800 175.800 414.800 176.000 ;
        RECT 415.600 175.800 416.400 179.800 ;
        RECT 417.800 176.400 418.600 179.800 ;
        RECT 417.800 175.800 419.600 176.400 ;
        RECT 411.000 175.400 414.600 175.800 ;
        RECT 411.600 174.400 412.400 174.800 ;
        RECT 415.600 174.400 416.200 175.800 ;
        RECT 410.800 173.800 412.400 174.400 ;
        RECT 410.800 173.600 411.600 173.800 ;
        RECT 413.800 173.600 416.400 174.400 ;
        RECT 404.400 171.700 408.400 172.300 ;
        RECT 404.400 171.600 405.200 171.700 ;
        RECT 401.200 169.600 402.600 170.200 ;
        RECT 403.200 169.600 404.200 170.200 ;
        RECT 402.000 168.400 402.600 169.600 ;
        RECT 402.000 167.600 402.800 168.400 ;
        RECT 403.400 164.400 404.200 169.600 ;
        RECT 403.400 163.600 405.200 164.400 ;
        RECT 403.400 162.200 404.200 163.600 ;
        RECT 407.600 162.200 408.400 171.700 ;
        RECT 412.400 171.600 413.200 173.200 ;
        RECT 413.800 170.200 414.400 173.600 ;
        RECT 418.800 172.300 419.600 175.800 ;
        RECT 420.400 173.600 421.200 175.200 ;
        RECT 422.000 175.000 422.800 179.800 ;
        RECT 426.400 178.400 427.200 179.800 ;
        RECT 425.200 177.800 427.200 178.400 ;
        RECT 430.800 177.800 431.600 179.800 ;
        RECT 435.000 178.400 436.200 179.800 ;
        RECT 434.800 177.800 436.200 178.400 ;
        RECT 425.200 177.000 426.000 177.800 ;
        RECT 430.800 177.200 431.400 177.800 ;
        RECT 426.800 176.400 427.600 177.200 ;
        RECT 428.600 176.600 431.400 177.200 ;
        RECT 434.800 177.000 435.600 177.800 ;
        RECT 428.600 176.400 429.400 176.600 ;
        RECT 422.800 174.200 424.400 174.400 ;
        RECT 427.000 174.200 427.600 176.400 ;
        RECT 436.600 175.400 437.400 175.600 ;
        RECT 439.600 175.400 440.400 179.800 ;
        RECT 436.600 174.800 440.400 175.400 ;
        RECT 446.000 175.800 446.800 179.800 ;
        RECT 450.400 176.200 452.000 179.800 ;
        RECT 446.000 175.200 448.200 175.800 ;
        RECT 449.200 175.400 450.800 175.600 ;
        RECT 447.400 175.000 448.200 175.200 ;
        RECT 432.600 174.200 434.000 174.400 ;
        RECT 422.800 173.600 434.000 174.200 ;
        RECT 425.800 173.400 426.600 173.600 ;
        RECT 415.700 171.700 419.600 172.300 ;
        RECT 424.200 172.400 425.000 172.600 ;
        RECT 426.800 172.400 427.600 172.600 ;
        RECT 424.200 171.800 429.200 172.400 ;
        RECT 415.700 170.400 416.300 171.700 ;
        RECT 415.600 170.200 416.400 170.400 ;
        RECT 413.400 169.600 414.400 170.200 ;
        RECT 415.000 169.600 416.400 170.200 ;
        RECT 413.400 162.200 414.200 169.600 ;
        RECT 415.000 168.400 415.600 169.600 ;
        RECT 417.200 168.800 418.000 170.400 ;
        RECT 414.800 167.600 415.600 168.400 ;
        RECT 418.800 162.200 419.600 171.700 ;
        RECT 428.400 171.600 429.200 171.800 ;
        RECT 431.600 172.300 432.400 172.400 ;
        RECT 433.200 172.300 433.800 173.600 ;
        RECT 434.800 172.800 435.600 173.000 ;
        RECT 431.600 171.700 433.900 172.300 ;
        RECT 434.800 172.200 438.600 172.800 ;
        RECT 437.800 172.000 438.600 172.200 ;
        RECT 431.600 171.600 432.400 171.700 ;
        RECT 422.000 171.000 427.600 171.200 ;
        RECT 422.000 170.800 427.800 171.000 ;
        RECT 422.000 170.600 431.800 170.800 ;
        RECT 422.000 162.200 422.800 170.600 ;
        RECT 427.000 170.200 431.800 170.600 ;
        RECT 425.200 169.000 430.600 169.600 ;
        RECT 425.200 168.800 426.000 169.000 ;
        RECT 429.800 168.800 430.600 169.000 ;
        RECT 431.200 169.000 431.800 170.200 ;
        RECT 433.200 170.400 433.800 171.700 ;
        RECT 436.200 171.400 437.000 171.600 ;
        RECT 439.600 171.400 440.400 174.800 ;
        RECT 448.800 174.800 450.800 175.400 ;
        RECT 448.800 174.400 449.400 174.800 ;
        RECT 446.000 173.800 449.400 174.400 ;
        RECT 446.000 173.600 447.600 173.800 ;
        RECT 450.000 173.400 450.800 174.200 ;
        RECT 450.000 172.800 450.600 173.400 ;
        RECT 448.000 172.200 450.600 172.800 ;
        RECT 451.400 172.800 452.000 176.200 ;
        RECT 455.600 175.800 456.400 179.800 ;
        RECT 452.600 174.800 453.400 175.600 ;
        RECT 454.000 175.200 456.400 175.800 ;
        RECT 454.000 175.000 454.800 175.200 ;
        RECT 457.200 175.000 458.000 179.800 ;
        RECT 461.600 178.400 462.400 179.800 ;
        RECT 460.400 177.800 462.400 178.400 ;
        RECT 466.000 177.800 466.800 179.800 ;
        RECT 470.200 178.400 471.400 179.800 ;
        RECT 470.000 177.800 471.400 178.400 ;
        RECT 460.400 177.000 461.200 177.800 ;
        RECT 466.000 177.200 466.600 177.800 ;
        RECT 462.000 176.400 462.800 177.200 ;
        RECT 463.800 176.600 466.600 177.200 ;
        RECT 470.000 177.000 470.800 177.800 ;
        RECT 463.800 176.400 464.600 176.600 ;
        RECT 452.800 174.400 453.400 174.800 ;
        RECT 452.800 173.600 453.600 174.400 ;
        RECT 454.800 173.600 456.400 174.400 ;
        RECT 458.000 174.200 459.600 174.400 ;
        RECT 462.200 174.200 462.800 176.400 ;
        RECT 471.800 175.400 472.600 175.600 ;
        RECT 474.800 175.400 475.600 179.800 ;
        RECT 471.800 174.800 475.600 175.400 ;
        RECT 467.800 174.200 468.600 174.400 ;
        RECT 458.000 173.600 469.000 174.200 ;
        RECT 461.000 173.400 461.800 173.600 ;
        RECT 451.400 172.400 452.400 172.800 ;
        RECT 459.400 172.400 460.200 172.600 ;
        RECT 462.000 172.400 462.800 172.600 ;
        RECT 468.400 172.400 469.000 173.600 ;
        RECT 470.000 172.800 470.800 173.000 ;
        RECT 451.400 172.200 453.200 172.400 ;
        RECT 448.000 172.000 448.800 172.200 ;
        RECT 451.800 171.600 453.200 172.200 ;
        RECT 459.400 171.800 464.400 172.400 ;
        RECT 463.600 171.600 464.400 171.800 ;
        RECT 468.400 171.600 469.200 172.400 ;
        RECT 470.000 172.200 473.800 172.800 ;
        RECT 473.000 172.000 473.800 172.200 ;
        RECT 450.200 171.400 451.000 171.600 ;
        RECT 436.200 170.800 440.400 171.400 ;
        RECT 433.200 169.800 435.600 170.400 ;
        RECT 432.600 169.000 433.400 169.200 ;
        RECT 431.200 168.400 433.400 169.000 ;
        RECT 435.000 168.800 435.600 169.800 ;
        RECT 435.000 168.000 436.400 168.800 ;
        RECT 428.600 167.400 429.400 167.600 ;
        RECT 431.400 167.400 432.200 167.600 ;
        RECT 425.200 166.200 426.000 167.000 ;
        RECT 428.600 166.800 432.200 167.400 ;
        RECT 430.800 166.200 431.400 166.800 ;
        RECT 434.800 166.200 435.600 167.000 ;
        RECT 425.200 165.600 427.200 166.200 ;
        RECT 426.400 162.200 427.200 165.600 ;
        RECT 430.800 162.200 431.600 166.200 ;
        RECT 435.000 162.200 436.200 166.200 ;
        RECT 439.600 162.200 440.400 170.800 ;
        RECT 447.600 170.800 451.000 171.400 ;
        RECT 447.600 170.200 448.200 170.800 ;
        RECT 451.800 170.200 452.400 171.600 ;
        RECT 457.200 171.000 462.800 171.200 ;
        RECT 457.200 170.800 463.000 171.000 ;
        RECT 457.200 170.600 467.000 170.800 ;
        RECT 446.000 169.600 448.200 170.200 ;
        RECT 446.000 162.200 446.800 169.600 ;
        RECT 447.400 169.400 448.200 169.600 ;
        RECT 450.400 169.600 452.400 170.200 ;
        RECT 454.000 169.600 456.400 170.200 ;
        RECT 450.400 162.200 452.000 169.600 ;
        RECT 454.000 169.400 454.800 169.600 ;
        RECT 455.600 162.200 456.400 169.600 ;
        RECT 457.200 162.200 458.000 170.600 ;
        RECT 462.200 170.200 467.000 170.600 ;
        RECT 460.400 169.000 465.800 169.600 ;
        RECT 460.400 168.800 461.200 169.000 ;
        RECT 465.000 168.800 465.800 169.000 ;
        RECT 466.400 169.000 467.000 170.200 ;
        RECT 468.400 170.400 469.000 171.600 ;
        RECT 471.400 171.400 472.200 171.600 ;
        RECT 474.800 171.400 475.600 174.800 ;
        RECT 471.400 170.800 475.600 171.400 ;
        RECT 468.400 169.800 470.800 170.400 ;
        RECT 467.800 169.000 468.600 169.200 ;
        RECT 466.400 168.400 468.600 169.000 ;
        RECT 470.200 168.800 470.800 169.800 ;
        RECT 470.200 168.000 471.600 168.800 ;
        RECT 463.800 167.400 464.600 167.600 ;
        RECT 466.600 167.400 467.400 167.600 ;
        RECT 460.400 166.200 461.200 167.000 ;
        RECT 463.800 166.800 467.400 167.400 ;
        RECT 466.000 166.200 466.600 166.800 ;
        RECT 470.000 166.200 470.800 167.000 ;
        RECT 460.400 165.600 462.400 166.200 ;
        RECT 461.600 162.200 462.400 165.600 ;
        RECT 466.000 162.200 466.800 166.200 ;
        RECT 470.200 162.200 471.400 166.200 ;
        RECT 474.800 162.200 475.600 170.800 ;
        RECT 476.400 162.200 477.200 179.800 ;
        RECT 479.600 175.800 480.400 179.800 ;
        RECT 484.000 178.400 485.600 179.800 ;
        RECT 484.000 177.600 486.800 178.400 ;
        RECT 484.000 176.200 485.600 177.600 ;
        RECT 479.600 175.200 481.800 175.800 ;
        RECT 482.800 175.400 484.400 175.600 ;
        RECT 478.000 174.300 478.800 175.200 ;
        RECT 481.000 175.000 481.800 175.200 ;
        RECT 482.400 174.800 484.400 175.400 ;
        RECT 482.400 174.400 483.000 174.800 ;
        RECT 479.600 174.300 483.000 174.400 ;
        RECT 478.000 173.800 483.000 174.300 ;
        RECT 478.000 173.700 481.200 173.800 ;
        RECT 478.000 173.600 478.800 173.700 ;
        RECT 479.600 173.600 481.200 173.700 ;
        RECT 483.600 173.400 484.400 174.200 ;
        RECT 483.600 172.800 484.200 173.400 ;
        RECT 481.600 172.200 484.200 172.800 ;
        RECT 485.000 172.800 485.600 176.200 ;
        RECT 489.200 175.800 490.000 179.800 ;
        RECT 486.200 174.800 487.000 175.600 ;
        RECT 487.600 175.200 490.000 175.800 ;
        RECT 487.600 175.000 488.400 175.200 ;
        RECT 486.400 174.400 487.000 174.800 ;
        RECT 486.400 173.600 487.200 174.400 ;
        RECT 488.400 173.600 490.000 174.400 ;
        RECT 490.800 173.600 491.600 175.200 ;
        RECT 485.000 172.400 486.000 172.800 ;
        RECT 485.000 172.200 486.800 172.400 ;
        RECT 481.600 172.000 482.400 172.200 ;
        RECT 485.400 171.600 486.800 172.200 ;
        RECT 492.400 172.300 493.200 179.800 ;
        RECT 494.000 176.000 494.800 179.800 ;
        RECT 497.200 176.000 498.000 179.800 ;
        RECT 494.000 175.800 498.000 176.000 ;
        RECT 498.800 175.800 499.600 179.800 ;
        RECT 500.400 175.800 501.200 179.800 ;
        RECT 502.000 176.000 502.800 179.800 ;
        RECT 505.200 176.000 506.000 179.800 ;
        RECT 509.400 178.400 510.200 179.800 ;
        RECT 508.400 177.600 510.200 178.400 ;
        RECT 509.400 176.400 510.200 177.600 ;
        RECT 502.000 175.800 506.000 176.000 ;
        RECT 508.400 175.800 510.200 176.400 ;
        RECT 514.200 175.800 515.800 179.800 ;
        RECT 519.600 175.800 520.400 179.800 ;
        RECT 521.200 176.000 522.000 179.800 ;
        RECT 524.400 176.000 525.200 179.800 ;
        RECT 521.200 175.800 525.200 176.000 ;
        RECT 527.600 177.800 528.400 179.800 ;
        RECT 494.200 175.400 497.800 175.800 ;
        RECT 494.800 174.400 495.600 174.800 ;
        RECT 498.800 174.400 499.400 175.800 ;
        RECT 500.600 174.400 501.200 175.800 ;
        RECT 502.200 175.400 505.800 175.800 ;
        RECT 504.400 174.400 505.200 174.800 ;
        RECT 494.000 173.800 495.600 174.400 ;
        RECT 494.000 173.600 494.800 173.800 ;
        RECT 497.000 173.600 499.600 174.400 ;
        RECT 500.400 173.600 503.000 174.400 ;
        RECT 504.400 173.800 506.000 174.400 ;
        RECT 505.200 173.600 506.000 173.800 ;
        RECT 506.800 173.600 507.600 175.200 ;
        RECT 495.600 172.300 496.400 173.200 ;
        RECT 492.400 171.700 496.400 172.300 ;
        RECT 483.800 171.400 484.600 171.600 ;
        RECT 481.200 170.800 484.600 171.400 ;
        RECT 481.200 170.200 481.800 170.800 ;
        RECT 485.400 170.200 486.000 171.600 ;
        RECT 479.600 169.600 481.800 170.200 ;
        RECT 479.600 162.200 480.400 169.600 ;
        RECT 481.000 169.400 481.800 169.600 ;
        RECT 484.000 169.600 486.000 170.200 ;
        RECT 487.600 169.600 490.000 170.200 ;
        RECT 484.000 162.200 485.600 169.600 ;
        RECT 487.600 169.400 488.400 169.600 ;
        RECT 489.200 162.200 490.000 169.600 ;
        RECT 492.400 162.200 493.200 171.700 ;
        RECT 495.600 171.600 496.400 171.700 ;
        RECT 497.000 172.300 497.600 173.600 ;
        RECT 497.000 171.700 501.100 172.300 ;
        RECT 497.000 170.200 497.600 171.700 ;
        RECT 500.500 170.400 501.100 171.700 ;
        RECT 498.800 170.200 499.600 170.400 ;
        RECT 496.600 169.600 497.600 170.200 ;
        RECT 498.200 169.600 499.600 170.200 ;
        RECT 500.400 170.200 501.200 170.400 ;
        RECT 502.400 170.200 503.000 173.600 ;
        RECT 503.600 171.600 504.400 173.200 ;
        RECT 500.400 169.600 501.800 170.200 ;
        RECT 502.400 169.600 503.400 170.200 ;
        RECT 496.600 162.200 497.400 169.600 ;
        RECT 498.200 168.400 498.800 169.600 ;
        RECT 498.000 167.600 498.800 168.400 ;
        RECT 501.200 168.400 501.800 169.600 ;
        RECT 501.200 167.600 502.000 168.400 ;
        RECT 502.600 162.200 503.400 169.600 ;
        RECT 508.400 162.200 509.200 175.800 ;
        RECT 513.200 173.600 514.000 174.400 ;
        RECT 513.400 173.200 514.000 173.600 ;
        RECT 513.400 172.400 514.200 173.200 ;
        RECT 514.800 172.400 515.400 175.800 ;
        RECT 519.800 174.400 520.400 175.800 ;
        RECT 521.400 175.400 525.000 175.800 ;
        RECT 523.600 174.400 524.400 174.800 ;
        RECT 527.600 174.400 528.200 177.800 ;
        RECT 529.200 175.600 530.000 177.200 ;
        RECT 531.400 176.400 532.200 179.800 ;
        RECT 531.400 175.800 533.200 176.400 ;
        RECT 516.400 172.800 517.200 174.400 ;
        RECT 519.600 173.600 522.200 174.400 ;
        RECT 523.600 173.800 525.200 174.400 ;
        RECT 524.400 173.600 525.200 173.800 ;
        RECT 527.600 173.600 528.400 174.400 ;
        RECT 511.600 170.800 512.400 172.400 ;
        RECT 514.800 171.600 515.600 172.400 ;
        RECT 518.000 172.200 518.800 172.400 ;
        RECT 517.200 171.600 518.800 172.200 ;
        RECT 514.800 171.400 515.400 171.600 ;
        RECT 513.400 170.800 515.400 171.400 ;
        RECT 517.200 171.200 518.000 171.600 ;
        RECT 510.000 168.800 510.800 170.400 ;
        RECT 513.400 170.200 514.000 170.800 ;
        RECT 519.600 170.200 520.400 170.400 ;
        RECT 521.600 170.200 522.200 173.600 ;
        RECT 522.800 172.300 523.600 173.200 ;
        RECT 526.000 172.300 526.800 172.400 ;
        RECT 522.800 171.700 526.800 172.300 ;
        RECT 522.800 171.600 523.600 171.700 ;
        RECT 526.000 170.800 526.800 171.700 ;
        RECT 527.600 170.200 528.200 173.600 ;
        RECT 529.200 172.300 530.000 172.400 ;
        RECT 532.400 172.300 533.200 175.800 ;
        RECT 534.000 173.600 534.800 175.200 ;
        RECT 536.800 174.200 537.600 179.800 ;
        RECT 543.600 177.800 544.400 179.800 ;
        RECT 542.000 175.600 542.800 177.200 ;
        RECT 543.800 176.400 544.400 177.800 ;
        RECT 543.600 175.600 544.400 176.400 ;
        RECT 543.800 174.400 544.400 175.600 ;
        RECT 535.800 173.800 537.600 174.200 ;
        RECT 535.800 173.600 537.400 173.800 ;
        RECT 543.600 173.600 544.400 174.400 ;
        RECT 550.400 174.200 551.200 179.800 ;
        RECT 554.800 177.800 555.600 179.800 ;
        RECT 553.200 176.300 554.000 176.400 ;
        RECT 554.800 176.300 555.400 177.800 ;
        RECT 553.200 175.700 555.500 176.300 ;
        RECT 553.200 175.600 554.000 175.700 ;
        RECT 554.800 174.400 555.400 175.700 ;
        RECT 556.400 175.600 557.200 177.200 ;
        RECT 558.000 175.000 558.800 179.800 ;
        RECT 562.400 178.400 563.200 179.800 ;
        RECT 561.200 177.800 563.200 178.400 ;
        RECT 566.800 177.800 567.600 179.800 ;
        RECT 571.000 178.400 572.200 179.800 ;
        RECT 570.800 177.800 572.200 178.400 ;
        RECT 561.200 177.000 562.000 177.800 ;
        RECT 566.800 177.200 567.400 177.800 ;
        RECT 562.800 176.400 563.600 177.200 ;
        RECT 564.600 176.600 567.400 177.200 ;
        RECT 570.800 177.000 571.600 177.800 ;
        RECT 564.600 176.400 565.400 176.600 ;
        RECT 550.400 173.800 552.200 174.200 ;
        RECT 550.600 173.600 552.200 173.800 ;
        RECT 529.200 171.700 533.200 172.300 ;
        RECT 529.200 171.600 530.000 171.700 ;
        RECT 511.600 162.800 512.400 170.200 ;
        RECT 513.200 163.400 514.000 170.200 ;
        RECT 514.800 169.600 518.800 170.200 ;
        RECT 519.600 169.600 521.000 170.200 ;
        RECT 521.600 169.600 522.600 170.200 ;
        RECT 514.800 162.800 515.600 169.600 ;
        RECT 511.600 162.200 515.600 162.800 ;
        RECT 518.000 162.200 518.800 169.600 ;
        RECT 520.400 168.400 521.000 169.600 ;
        RECT 520.400 167.600 521.200 168.400 ;
        RECT 521.800 162.200 522.600 169.600 ;
        RECT 526.600 169.400 528.400 170.200 ;
        RECT 526.600 166.400 527.400 169.400 ;
        RECT 530.800 168.800 531.600 170.400 ;
        RECT 526.600 165.600 528.400 166.400 ;
        RECT 526.600 162.200 527.400 165.600 ;
        RECT 532.400 162.200 533.200 171.700 ;
        RECT 535.800 170.400 536.400 173.600 ;
        RECT 538.000 171.600 539.600 172.400 ;
        RECT 542.000 172.300 542.800 172.400 ;
        RECT 540.400 171.700 542.800 172.300 ;
        RECT 535.600 169.600 536.400 170.400 ;
        RECT 540.400 169.600 541.200 171.700 ;
        RECT 542.000 171.600 542.800 171.700 ;
        RECT 543.800 170.200 544.400 173.600 ;
        RECT 545.200 170.800 546.000 172.400 ;
        RECT 548.400 171.600 550.800 172.400 ;
        RECT 535.800 167.000 536.400 169.600 ;
        RECT 543.600 169.400 545.400 170.200 ;
        RECT 546.800 169.600 547.600 171.200 ;
        RECT 551.600 170.400 552.200 173.600 ;
        RECT 554.800 173.600 555.600 174.400 ;
        RECT 558.800 174.200 560.400 174.400 ;
        RECT 563.000 174.200 563.600 176.400 ;
        RECT 572.600 175.400 573.400 175.600 ;
        RECT 575.600 175.400 576.400 179.800 ;
        RECT 572.600 174.800 576.400 175.400 ;
        RECT 568.600 174.200 569.400 174.400 ;
        RECT 558.800 173.600 569.800 174.200 ;
        RECT 553.200 170.800 554.000 172.400 ;
        RECT 551.600 169.600 552.400 170.400 ;
        RECT 554.800 170.200 555.400 173.600 ;
        RECT 561.800 173.400 562.600 173.600 ;
        RECT 560.200 172.400 561.000 172.600 ;
        RECT 569.200 172.400 569.800 173.600 ;
        RECT 570.800 172.800 571.600 173.000 ;
        RECT 560.200 172.300 565.200 172.400 ;
        RECT 566.000 172.300 566.800 172.400 ;
        RECT 560.200 171.800 566.800 172.300 ;
        RECT 564.400 171.700 566.800 171.800 ;
        RECT 564.400 171.600 565.200 171.700 ;
        RECT 566.000 171.600 566.800 171.700 ;
        RECT 569.200 171.600 570.000 172.400 ;
        RECT 570.800 172.200 574.600 172.800 ;
        RECT 573.800 172.000 574.600 172.200 ;
        RECT 558.000 171.000 563.600 171.200 ;
        RECT 558.000 170.800 563.800 171.000 ;
        RECT 558.000 170.600 567.800 170.800 ;
        RECT 537.200 167.600 538.000 169.200 ;
        RECT 535.800 166.400 539.400 167.000 ;
        RECT 535.800 166.200 536.400 166.400 ;
        RECT 535.600 162.200 536.400 166.200 ;
        RECT 538.800 166.200 539.400 166.400 ;
        RECT 538.800 162.200 539.600 166.200 ;
        RECT 544.600 162.200 545.400 169.400 ;
        RECT 550.000 167.600 550.800 169.200 ;
        RECT 551.600 167.000 552.200 169.600 ;
        RECT 548.600 166.400 552.200 167.000 ;
        RECT 548.600 166.200 549.200 166.400 ;
        RECT 548.400 162.200 549.200 166.200 ;
        RECT 551.600 166.200 552.200 166.400 ;
        RECT 553.800 169.400 555.600 170.200 ;
        RECT 551.600 162.200 552.400 166.200 ;
        RECT 553.800 162.200 554.600 169.400 ;
        RECT 558.000 162.200 558.800 170.600 ;
        RECT 563.000 170.200 567.800 170.600 ;
        RECT 561.200 169.000 566.600 169.600 ;
        RECT 561.200 168.800 562.000 169.000 ;
        RECT 565.800 168.800 566.600 169.000 ;
        RECT 567.200 169.000 567.800 170.200 ;
        RECT 569.200 170.400 569.800 171.600 ;
        RECT 572.200 171.400 573.000 171.600 ;
        RECT 575.600 171.400 576.400 174.800 ;
        RECT 577.200 175.200 578.000 179.800 ;
        RECT 577.200 174.600 579.400 175.200 ;
        RECT 577.200 171.600 578.000 173.200 ;
        RECT 578.800 171.600 579.400 174.600 ;
        RECT 572.200 170.800 576.400 171.400 ;
        RECT 569.200 169.800 571.600 170.400 ;
        RECT 568.600 169.000 569.400 169.200 ;
        RECT 567.200 168.400 569.400 169.000 ;
        RECT 571.000 168.800 571.600 169.800 ;
        RECT 571.000 168.000 572.400 168.800 ;
        RECT 564.600 167.400 565.400 167.600 ;
        RECT 567.400 167.400 568.200 167.600 ;
        RECT 561.200 166.200 562.000 167.000 ;
        RECT 564.600 166.800 568.200 167.400 ;
        RECT 566.800 166.200 567.400 166.800 ;
        RECT 570.800 166.200 571.600 167.000 ;
        RECT 561.200 165.600 563.200 166.200 ;
        RECT 562.400 162.200 563.200 165.600 ;
        RECT 566.800 162.200 567.600 166.200 ;
        RECT 571.000 162.200 572.200 166.200 ;
        RECT 575.600 162.200 576.400 170.800 ;
        RECT 578.800 170.800 580.000 171.600 ;
        RECT 578.800 170.200 579.400 170.800 ;
        RECT 577.200 169.600 579.400 170.200 ;
        RECT 577.200 162.200 578.000 169.600 ;
        RECT 2.800 155.800 3.600 159.800 ;
        RECT 3.000 151.600 3.600 155.800 ;
        RECT 6.000 151.800 6.800 159.800 ;
        RECT 3.000 151.000 5.400 151.600 ;
        RECT 2.800 149.600 3.600 150.400 ;
        RECT 1.200 147.600 2.000 149.200 ;
        RECT 3.000 148.800 3.600 149.600 ;
        RECT 3.000 148.200 4.000 148.800 ;
        RECT 3.200 148.000 4.000 148.200 ;
        RECT 4.800 147.600 5.400 151.000 ;
        RECT 6.200 150.400 6.800 151.800 ;
        RECT 7.600 151.200 8.400 159.800 ;
        RECT 11.800 152.400 12.600 159.800 ;
        RECT 16.600 152.400 17.400 159.800 ;
        RECT 18.000 153.600 18.800 154.400 ;
        RECT 18.200 152.400 18.800 153.600 ;
        RECT 11.800 151.800 13.200 152.400 ;
        RECT 16.600 151.800 17.600 152.400 ;
        RECT 18.200 151.800 19.600 152.400 ;
        RECT 20.400 151.800 21.200 159.800 ;
        RECT 22.000 152.400 22.800 159.800 ;
        RECT 25.200 152.400 26.000 159.800 ;
        RECT 22.000 151.800 26.000 152.400 ;
        RECT 26.800 151.800 27.600 159.800 ;
        RECT 28.400 152.400 29.200 159.800 ;
        RECT 31.600 152.400 32.400 159.800 ;
        RECT 34.000 153.600 34.800 154.400 ;
        RECT 34.000 152.400 34.600 153.600 ;
        RECT 35.400 152.400 36.200 159.800 ;
        RECT 42.200 158.400 43.000 159.800 ;
        RECT 41.200 157.600 43.000 158.400 ;
        RECT 28.400 151.800 32.400 152.400 ;
        RECT 33.200 151.800 34.600 152.400 ;
        RECT 35.200 151.800 36.200 152.400 ;
        RECT 42.200 152.400 43.000 157.600 ;
        RECT 43.600 153.600 44.400 154.400 ;
        RECT 43.800 152.400 44.400 153.600 ;
        RECT 42.200 151.800 43.200 152.400 ;
        RECT 43.800 152.300 45.200 152.400 ;
        RECT 47.600 152.300 48.400 159.800 ;
        RECT 43.800 151.800 48.400 152.300 ;
        RECT 12.400 151.600 13.200 151.800 ;
        RECT 7.600 150.800 11.600 151.200 ;
        RECT 7.600 150.600 11.800 150.800 ;
        RECT 6.000 149.600 6.800 150.400 ;
        RECT 11.000 150.000 11.800 150.600 ;
        RECT 12.600 150.400 13.200 151.600 ;
        RECT 4.800 147.400 5.600 147.600 ;
        RECT 2.600 147.000 5.600 147.400 ;
        RECT 1.400 146.800 5.600 147.000 ;
        RECT 1.400 146.400 3.200 146.800 ;
        RECT 1.400 146.200 2.000 146.400 ;
        RECT 6.200 146.200 6.800 149.600 ;
        RECT 9.600 148.400 10.400 149.200 ;
        RECT 9.200 147.600 10.200 148.400 ;
        RECT 11.200 147.000 11.800 150.000 ;
        RECT 12.400 149.600 13.200 150.400 ;
        RECT 9.400 146.400 11.800 147.000 ;
        RECT 1.200 142.200 2.000 146.200 ;
        RECT 5.400 145.200 6.800 146.200 ;
        RECT 5.400 144.400 6.200 145.200 ;
        RECT 7.600 144.800 8.400 146.400 ;
        RECT 5.400 143.600 6.800 144.400 ;
        RECT 9.400 144.200 10.000 146.400 ;
        RECT 12.600 146.200 13.200 149.600 ;
        RECT 15.600 148.800 16.400 150.400 ;
        RECT 17.000 148.400 17.600 151.800 ;
        RECT 18.800 151.600 19.600 151.800 ;
        RECT 20.600 150.400 21.200 151.800 ;
        RECT 24.400 150.400 25.200 150.800 ;
        RECT 27.000 150.400 27.600 151.800 ;
        RECT 33.200 151.600 34.000 151.800 ;
        RECT 30.800 150.400 31.600 150.800 ;
        RECT 20.400 149.800 22.800 150.400 ;
        RECT 24.400 149.800 26.000 150.400 ;
        RECT 20.400 149.600 21.200 149.800 ;
        RECT 14.000 148.200 14.800 148.400 ;
        RECT 14.000 147.600 15.600 148.200 ;
        RECT 17.000 147.600 19.600 148.400 ;
        RECT 14.800 147.200 15.600 147.600 ;
        RECT 14.200 146.200 17.800 146.600 ;
        RECT 18.800 146.400 19.400 147.600 ;
        RECT 5.400 142.200 6.200 143.600 ;
        RECT 9.200 142.200 10.000 144.200 ;
        RECT 12.400 142.200 13.200 146.200 ;
        RECT 14.000 146.000 18.000 146.200 ;
        RECT 14.000 142.200 14.800 146.000 ;
        RECT 17.200 142.200 18.000 146.000 ;
        RECT 18.800 142.200 19.600 146.400 ;
        RECT 20.400 145.600 21.200 146.400 ;
        RECT 22.200 146.200 22.800 149.800 ;
        RECT 25.200 149.600 26.000 149.800 ;
        RECT 26.800 149.800 29.200 150.400 ;
        RECT 30.800 149.800 32.400 150.400 ;
        RECT 26.800 149.600 27.600 149.800 ;
        RECT 28.400 149.600 29.200 149.800 ;
        RECT 31.600 149.600 32.400 149.800 ;
        RECT 23.600 147.600 24.400 149.200 ;
        RECT 20.600 144.800 21.400 145.600 ;
        RECT 22.000 142.200 22.800 146.200 ;
        RECT 26.800 145.600 27.600 146.400 ;
        RECT 28.600 146.200 29.200 149.600 ;
        RECT 30.000 147.600 30.800 149.200 ;
        RECT 35.200 148.400 35.800 151.800 ;
        RECT 36.400 148.800 37.200 150.400 ;
        RECT 41.200 148.800 42.000 150.400 ;
        RECT 42.600 148.400 43.200 151.800 ;
        RECT 44.400 151.700 48.400 151.800 ;
        RECT 44.400 151.600 45.200 151.700 ;
        RECT 33.200 147.600 35.800 148.400 ;
        RECT 38.000 148.200 38.800 148.400 ;
        RECT 37.200 147.600 38.800 148.200 ;
        RECT 39.600 148.200 40.400 148.400 ;
        RECT 39.600 147.600 41.200 148.200 ;
        RECT 42.600 147.600 45.200 148.400 ;
        RECT 33.400 146.200 34.000 147.600 ;
        RECT 37.200 147.200 38.000 147.600 ;
        RECT 40.400 147.200 41.200 147.600 ;
        RECT 35.000 146.200 38.600 146.600 ;
        RECT 39.800 146.200 43.400 146.600 ;
        RECT 44.400 146.200 45.000 147.600 ;
        RECT 46.000 146.800 46.800 148.400 ;
        RECT 47.600 146.200 48.400 151.700 ;
        RECT 49.200 151.600 50.000 153.200 ;
        RECT 50.800 146.800 51.600 148.400 ;
        RECT 52.400 146.200 53.200 159.800 ;
        RECT 54.000 151.600 54.800 153.200 ;
        RECT 58.200 152.400 59.000 159.800 ;
        RECT 59.600 153.600 60.400 154.400 ;
        RECT 59.800 152.400 60.400 153.600 ;
        RECT 64.600 152.400 65.400 159.800 ;
        RECT 66.000 153.600 66.800 154.400 ;
        RECT 66.200 152.400 66.800 153.600 ;
        RECT 68.400 152.400 69.200 159.800 ;
        RECT 72.800 154.400 74.400 159.800 ;
        RECT 72.800 153.600 75.600 154.400 ;
        RECT 70.000 152.400 70.800 152.600 ;
        RECT 72.800 152.400 74.400 153.600 ;
        RECT 58.200 151.800 59.200 152.400 ;
        RECT 59.800 151.800 61.200 152.400 ;
        RECT 64.600 151.800 65.600 152.400 ;
        RECT 66.200 151.800 67.600 152.400 ;
        RECT 68.400 151.800 70.800 152.400 ;
        RECT 72.400 151.800 74.400 152.400 ;
        RECT 76.600 152.400 77.400 152.600 ;
        RECT 78.000 152.400 78.800 159.800 ;
        RECT 76.600 151.800 78.800 152.400 ;
        RECT 79.600 152.400 80.400 159.800 ;
        RECT 82.800 159.200 86.800 159.800 ;
        RECT 82.800 152.400 83.600 159.200 ;
        RECT 79.600 151.800 83.600 152.400 ;
        RECT 84.400 151.800 85.200 158.600 ;
        RECT 86.000 151.800 86.800 159.200 ;
        RECT 87.600 152.400 88.400 159.800 ;
        RECT 90.800 159.200 94.800 159.800 ;
        RECT 90.800 152.400 91.600 159.200 ;
        RECT 87.600 151.800 91.600 152.400 ;
        RECT 92.400 151.800 93.200 158.600 ;
        RECT 94.000 151.800 94.800 159.200 ;
        RECT 55.600 150.300 56.400 150.400 ;
        RECT 57.200 150.300 58.000 150.400 ;
        RECT 55.600 149.700 58.000 150.300 ;
        RECT 55.600 149.600 56.400 149.700 ;
        RECT 57.200 148.800 58.000 149.700 ;
        RECT 58.600 150.300 59.200 151.800 ;
        RECT 60.400 151.600 61.200 151.800 ;
        RECT 63.600 150.300 64.400 150.400 ;
        RECT 58.600 149.700 64.400 150.300 ;
        RECT 58.600 148.400 59.200 149.700 ;
        RECT 63.600 148.800 64.400 149.700 ;
        RECT 65.000 148.400 65.600 151.800 ;
        RECT 66.800 151.600 67.600 151.800 ;
        RECT 72.400 150.400 73.000 151.800 ;
        RECT 76.600 151.200 77.200 151.800 ;
        RECT 84.400 151.200 85.000 151.800 ;
        RECT 92.400 151.200 93.000 151.800 ;
        RECT 73.800 150.600 77.200 151.200 ;
        RECT 73.800 150.400 74.600 150.600 ;
        RECT 80.400 150.400 81.200 150.800 ;
        RECT 83.000 150.600 85.000 151.200 ;
        RECT 83.000 150.400 83.600 150.600 ;
        RECT 71.600 149.800 73.000 150.400 ;
        RECT 76.000 149.800 76.800 150.000 ;
        RECT 71.600 149.600 73.400 149.800 ;
        RECT 72.400 149.200 73.400 149.600 ;
        RECT 55.600 148.200 56.400 148.400 ;
        RECT 55.600 147.600 57.200 148.200 ;
        RECT 58.600 147.600 61.200 148.400 ;
        RECT 62.000 148.200 62.800 148.400 ;
        RECT 62.000 147.600 63.600 148.200 ;
        RECT 65.000 147.600 67.600 148.400 ;
        RECT 68.400 147.600 70.000 148.400 ;
        RECT 71.200 147.600 72.000 148.400 ;
        RECT 56.400 147.200 57.200 147.600 ;
        RECT 55.800 146.200 59.400 146.600 ;
        RECT 60.400 146.200 61.000 147.600 ;
        RECT 62.800 147.200 63.600 147.600 ;
        RECT 62.200 146.200 65.800 146.600 ;
        RECT 66.800 146.400 67.400 147.600 ;
        RECT 71.400 147.200 72.000 147.600 ;
        RECT 70.000 146.800 70.800 147.000 ;
        RECT 27.000 144.800 27.800 145.600 ;
        RECT 28.400 142.200 29.200 146.200 ;
        RECT 33.200 142.200 34.000 146.200 ;
        RECT 34.800 146.000 38.800 146.200 ;
        RECT 34.800 142.200 35.600 146.000 ;
        RECT 38.000 142.200 38.800 146.000 ;
        RECT 39.600 146.000 43.600 146.200 ;
        RECT 39.600 142.200 40.400 146.000 ;
        RECT 42.800 142.200 43.600 146.000 ;
        RECT 44.400 142.200 45.200 146.200 ;
        RECT 47.600 145.600 49.400 146.200 ;
        RECT 52.400 145.600 54.200 146.200 ;
        RECT 48.600 142.200 49.400 145.600 ;
        RECT 53.400 144.400 54.200 145.600 ;
        RECT 55.600 146.000 59.600 146.200 ;
        RECT 53.400 143.600 54.800 144.400 ;
        RECT 53.400 142.200 54.200 143.600 ;
        RECT 55.600 142.200 56.400 146.000 ;
        RECT 58.800 142.200 59.600 146.000 ;
        RECT 60.400 142.200 61.200 146.200 ;
        RECT 62.000 146.000 66.000 146.200 ;
        RECT 62.000 142.200 62.800 146.000 ;
        RECT 65.200 142.200 66.000 146.000 ;
        RECT 66.800 142.200 67.600 146.400 ;
        RECT 68.400 146.200 70.800 146.800 ;
        RECT 71.400 146.400 72.200 147.200 ;
        RECT 68.400 142.200 69.200 146.200 ;
        RECT 72.800 145.800 73.400 149.200 ;
        RECT 74.200 149.200 76.800 149.800 ;
        RECT 79.600 149.800 81.200 150.400 ;
        RECT 79.600 149.600 80.400 149.800 ;
        RECT 82.800 149.600 83.600 150.400 ;
        RECT 86.000 149.600 86.800 151.200 ;
        RECT 88.400 150.400 89.200 150.800 ;
        RECT 91.000 150.600 93.000 151.200 ;
        RECT 91.000 150.400 91.600 150.600 ;
        RECT 87.600 149.800 89.200 150.400 ;
        RECT 87.600 149.600 88.400 149.800 ;
        RECT 90.800 149.600 91.600 150.400 ;
        RECT 94.000 150.300 94.800 151.200 ;
        RECT 95.600 150.300 96.400 159.800 ;
        RECT 101.400 152.600 102.200 159.800 ;
        RECT 100.400 151.800 102.200 152.600 ;
        RECT 94.000 149.700 96.400 150.300 ;
        RECT 94.000 149.600 94.800 149.700 ;
        RECT 74.200 148.600 74.800 149.200 ;
        RECT 74.000 147.800 74.800 148.600 ;
        RECT 77.200 148.200 78.800 148.400 ;
        RECT 75.400 147.600 78.800 148.200 ;
        RECT 81.200 147.600 82.000 149.200 ;
        RECT 75.400 147.200 76.000 147.600 ;
        RECT 74.000 146.600 76.000 147.200 ;
        RECT 76.600 146.800 77.400 147.000 ;
        RECT 74.000 146.400 75.600 146.600 ;
        RECT 76.600 146.200 78.800 146.800 ;
        RECT 83.000 146.200 83.600 149.600 ;
        RECT 84.200 148.800 85.000 149.600 ;
        RECT 84.400 148.400 85.000 148.800 ;
        RECT 84.400 147.600 85.200 148.400 ;
        RECT 89.200 147.600 90.000 149.200 ;
        RECT 91.000 146.200 91.600 149.600 ;
        RECT 92.200 148.800 93.000 149.600 ;
        RECT 92.400 148.400 93.000 148.800 ;
        RECT 92.400 147.600 93.200 148.400 ;
        RECT 72.800 142.200 74.400 145.800 ;
        RECT 78.000 142.200 78.800 146.200 ;
        RECT 82.600 142.200 84.200 146.200 ;
        RECT 90.600 142.200 92.200 146.200 ;
        RECT 95.600 142.200 96.400 149.700 ;
        RECT 97.200 150.300 98.000 150.400 ;
        RECT 100.600 150.300 101.200 151.800 ;
        RECT 103.600 151.600 104.400 153.200 ;
        RECT 97.200 149.700 101.200 150.300 ;
        RECT 97.200 149.600 98.000 149.700 ;
        RECT 100.600 148.400 101.200 149.700 ;
        RECT 102.000 150.300 102.800 151.200 ;
        RECT 103.700 150.300 104.300 151.600 ;
        RECT 102.000 149.700 104.300 150.300 ;
        RECT 102.000 149.600 102.800 149.700 ;
        RECT 100.400 147.600 101.200 148.400 ;
        RECT 97.200 144.800 98.000 146.400 ;
        RECT 98.800 144.800 99.600 146.400 ;
        RECT 100.600 144.200 101.200 147.600 ;
        RECT 105.200 146.200 106.000 159.800 ;
        RECT 106.800 154.300 107.600 154.400 ;
        RECT 108.400 154.300 109.200 159.800 ;
        RECT 106.800 153.700 109.200 154.300 ;
        RECT 106.800 153.600 107.600 153.700 ;
        RECT 106.800 146.800 107.600 148.400 ;
        RECT 104.200 145.600 106.000 146.200 ;
        RECT 104.200 144.400 105.000 145.600 ;
        RECT 100.400 142.200 101.200 144.200 ;
        RECT 103.600 143.600 105.000 144.400 ;
        RECT 104.200 142.200 105.000 143.600 ;
        RECT 108.400 142.200 109.200 153.700 ;
        RECT 111.600 152.400 112.400 159.800 ;
        RECT 113.200 152.400 114.000 152.600 ;
        RECT 116.000 152.400 117.600 159.800 ;
        RECT 111.600 151.800 114.000 152.400 ;
        RECT 115.600 151.800 117.600 152.400 ;
        RECT 119.800 152.400 120.600 152.600 ;
        RECT 121.200 152.400 122.000 159.800 ;
        RECT 119.800 151.800 122.000 152.400 ;
        RECT 122.800 152.400 123.600 159.800 ;
        RECT 126.000 152.400 126.800 159.800 ;
        RECT 122.800 151.800 126.800 152.400 ;
        RECT 127.600 151.800 128.400 159.800 ;
        RECT 129.200 152.400 130.000 159.800 ;
        RECT 132.400 159.200 136.400 159.800 ;
        RECT 132.400 152.400 133.200 159.200 ;
        RECT 129.200 151.800 133.200 152.400 ;
        RECT 134.000 151.800 134.800 158.600 ;
        RECT 135.600 151.800 136.400 159.200 ;
        RECT 142.000 152.400 142.800 159.800 ;
        RECT 143.600 152.400 144.400 152.600 ;
        RECT 146.400 152.400 148.000 159.800 ;
        RECT 142.000 151.800 144.400 152.400 ;
        RECT 146.000 151.800 148.000 152.400 ;
        RECT 150.200 152.400 151.000 152.600 ;
        RECT 151.600 152.400 152.400 159.800 ;
        RECT 150.200 151.800 152.400 152.400 ;
        RECT 115.600 150.400 116.200 151.800 ;
        RECT 119.800 151.200 120.400 151.800 ;
        RECT 117.000 150.600 120.400 151.200 ;
        RECT 117.000 150.400 117.800 150.600 ;
        RECT 123.600 150.400 124.400 150.800 ;
        RECT 127.600 150.400 128.200 151.800 ;
        RECT 134.000 151.200 134.600 151.800 ;
        RECT 130.000 150.400 130.800 150.800 ;
        RECT 132.600 150.600 134.600 151.200 ;
        RECT 132.600 150.400 133.200 150.600 ;
        RECT 114.800 149.800 116.200 150.400 ;
        RECT 119.200 149.800 120.000 150.000 ;
        RECT 114.800 149.600 116.600 149.800 ;
        RECT 115.600 149.200 116.600 149.600 ;
        RECT 111.600 147.600 113.200 148.400 ;
        RECT 114.400 147.600 115.200 148.400 ;
        RECT 114.600 147.200 115.200 147.600 ;
        RECT 113.200 146.800 114.000 147.000 ;
        RECT 110.000 144.800 110.800 146.400 ;
        RECT 111.600 146.200 114.000 146.800 ;
        RECT 114.600 146.400 115.400 147.200 ;
        RECT 111.600 142.200 112.400 146.200 ;
        RECT 116.000 145.800 116.600 149.200 ;
        RECT 117.400 149.200 120.000 149.800 ;
        RECT 122.800 149.800 124.400 150.400 ;
        RECT 126.000 149.800 128.400 150.400 ;
        RECT 122.800 149.600 123.600 149.800 ;
        RECT 117.400 148.600 118.000 149.200 ;
        RECT 117.200 147.800 118.000 148.600 ;
        RECT 120.400 148.300 122.000 148.400 ;
        RECT 124.400 148.300 125.200 149.200 ;
        RECT 120.400 148.200 125.200 148.300 ;
        RECT 118.600 147.700 125.200 148.200 ;
        RECT 118.600 147.600 122.000 147.700 ;
        RECT 124.400 147.600 125.200 147.700 ;
        RECT 126.000 148.300 126.600 149.800 ;
        RECT 127.600 149.600 128.400 149.800 ;
        RECT 129.200 149.800 130.800 150.400 ;
        RECT 129.200 149.600 130.000 149.800 ;
        RECT 132.400 149.600 133.200 150.400 ;
        RECT 135.600 149.600 136.400 151.200 ;
        RECT 146.000 150.400 146.600 151.800 ;
        RECT 150.200 151.200 150.800 151.800 ;
        RECT 147.400 150.600 150.800 151.200 ;
        RECT 153.200 151.400 154.000 159.800 ;
        RECT 157.600 156.400 158.400 159.800 ;
        RECT 156.400 155.800 158.400 156.400 ;
        RECT 162.000 155.800 162.800 159.800 ;
        RECT 166.200 155.800 167.400 159.800 ;
        RECT 156.400 155.000 157.200 155.800 ;
        RECT 162.000 155.200 162.600 155.800 ;
        RECT 159.800 154.600 163.400 155.200 ;
        RECT 166.000 155.000 166.800 155.800 ;
        RECT 159.800 154.400 160.600 154.600 ;
        RECT 162.600 154.400 163.400 154.600 ;
        RECT 156.400 153.000 157.200 153.200 ;
        RECT 161.000 153.000 161.800 153.200 ;
        RECT 156.400 152.400 161.800 153.000 ;
        RECT 162.400 153.000 164.600 153.600 ;
        RECT 162.400 151.800 163.000 153.000 ;
        RECT 163.800 152.800 164.600 153.000 ;
        RECT 166.200 153.200 167.600 154.000 ;
        RECT 166.200 152.200 166.800 153.200 ;
        RECT 158.200 151.400 163.000 151.800 ;
        RECT 153.200 151.200 163.000 151.400 ;
        RECT 164.400 151.600 166.800 152.200 ;
        RECT 153.200 151.000 159.000 151.200 ;
        RECT 153.200 150.800 158.800 151.000 ;
        RECT 147.400 150.400 148.200 150.600 ;
        RECT 164.400 150.400 165.000 151.600 ;
        RECT 170.800 151.200 171.600 159.800 ;
        RECT 174.000 151.200 174.800 159.800 ;
        RECT 177.200 151.200 178.000 159.800 ;
        RECT 180.400 151.200 181.200 159.800 ;
        RECT 183.600 151.200 184.400 159.800 ;
        RECT 186.800 152.400 187.600 159.800 ;
        RECT 188.200 152.400 189.000 152.600 ;
        RECT 186.800 151.800 189.000 152.400 ;
        RECT 191.200 152.400 192.800 159.800 ;
        RECT 194.800 152.400 195.600 152.600 ;
        RECT 196.400 152.400 197.200 159.800 ;
        RECT 191.200 151.800 193.200 152.400 ;
        RECT 194.800 151.800 197.200 152.400 ;
        RECT 198.000 152.400 198.800 159.800 ;
        RECT 199.800 152.400 200.600 152.600 ;
        RECT 198.000 151.800 200.600 152.400 ;
        RECT 202.400 151.800 204.000 159.800 ;
        RECT 206.000 152.400 206.800 152.600 ;
        RECT 207.600 152.400 208.400 159.800 ;
        RECT 206.000 151.800 208.400 152.400 ;
        RECT 167.400 150.600 171.600 151.200 ;
        RECT 167.400 150.400 168.200 150.600 ;
        RECT 145.200 149.800 146.600 150.400 ;
        RECT 159.600 150.200 160.400 150.400 ;
        RECT 149.600 149.800 150.400 150.000 ;
        RECT 145.200 149.600 147.000 149.800 ;
        RECT 130.800 148.300 131.600 149.200 ;
        RECT 126.000 147.700 131.600 148.300 ;
        RECT 118.600 147.200 119.200 147.600 ;
        RECT 117.200 146.600 119.200 147.200 ;
        RECT 119.800 146.800 120.600 147.000 ;
        RECT 117.200 146.400 118.800 146.600 ;
        RECT 119.800 146.200 122.000 146.800 ;
        RECT 116.000 142.200 117.600 145.800 ;
        RECT 121.200 142.200 122.000 146.200 ;
        RECT 126.000 146.200 126.600 147.700 ;
        RECT 130.800 147.600 131.600 147.700 ;
        RECT 132.600 146.400 133.200 149.600 ;
        RECT 133.800 148.800 134.600 149.600 ;
        RECT 146.000 149.200 147.000 149.600 ;
        RECT 134.000 148.400 134.600 148.800 ;
        RECT 134.000 147.600 134.800 148.400 ;
        RECT 142.000 147.600 143.600 148.400 ;
        RECT 144.800 147.600 145.600 148.400 ;
        RECT 145.000 147.200 145.600 147.600 ;
        RECT 143.600 146.800 144.400 147.000 ;
        RECT 126.000 142.200 126.800 146.200 ;
        RECT 127.600 145.600 128.400 146.400 ;
        RECT 132.600 146.200 134.800 146.400 ;
        RECT 132.200 145.600 134.800 146.200 ;
        RECT 142.000 146.200 144.400 146.800 ;
        RECT 145.000 146.400 145.800 147.200 ;
        RECT 127.400 144.800 128.200 145.600 ;
        RECT 132.200 142.200 133.800 145.600 ;
        RECT 142.000 142.200 142.800 146.200 ;
        RECT 146.400 145.800 147.000 149.200 ;
        RECT 147.800 149.200 150.400 149.800 ;
        RECT 155.400 149.600 160.400 150.200 ;
        RECT 164.400 149.600 165.200 150.400 ;
        RECT 169.000 149.800 169.800 150.000 ;
        RECT 155.400 149.400 156.200 149.600 ;
        RECT 158.000 149.400 158.800 149.600 ;
        RECT 147.800 148.600 148.400 149.200 ;
        RECT 147.600 147.800 148.400 148.600 ;
        RECT 157.000 148.400 157.800 148.600 ;
        RECT 164.400 148.400 165.000 149.600 ;
        RECT 166.000 149.200 169.800 149.800 ;
        RECT 166.000 149.000 166.800 149.200 ;
        RECT 150.800 148.200 152.400 148.400 ;
        RECT 149.000 147.600 152.400 148.200 ;
        RECT 154.000 147.800 165.000 148.400 ;
        RECT 154.000 147.600 155.600 147.800 ;
        RECT 149.000 147.200 149.600 147.600 ;
        RECT 147.600 146.600 149.600 147.200 ;
        RECT 150.200 146.800 151.000 147.000 ;
        RECT 147.600 146.400 149.200 146.600 ;
        RECT 150.200 146.200 152.400 146.800 ;
        RECT 146.400 144.400 148.000 145.800 ;
        RECT 146.400 143.600 149.200 144.400 ;
        RECT 146.400 142.200 148.000 143.600 ;
        RECT 151.600 142.200 152.400 146.200 ;
        RECT 153.200 142.200 154.000 147.000 ;
        RECT 158.200 145.600 158.800 147.800 ;
        RECT 163.800 147.600 164.600 147.800 ;
        RECT 170.800 147.200 171.600 150.600 ;
        RECT 167.800 146.600 171.600 147.200 ;
        RECT 172.400 150.400 174.800 151.200 ;
        RECT 175.800 150.400 178.000 151.200 ;
        RECT 179.000 150.400 181.200 151.200 ;
        RECT 182.600 150.400 184.400 151.200 ;
        RECT 188.400 151.200 189.000 151.800 ;
        RECT 188.400 150.600 191.800 151.200 ;
        RECT 191.000 150.400 191.800 150.600 ;
        RECT 192.600 150.400 193.200 151.800 ;
        RECT 201.000 150.400 201.800 150.600 ;
        RECT 203.000 150.400 203.600 151.800 ;
        RECT 209.200 151.600 210.000 153.200 ;
        RECT 172.400 147.600 173.200 150.400 ;
        RECT 175.800 149.000 176.600 150.400 ;
        RECT 179.000 149.000 179.800 150.400 ;
        RECT 182.600 149.000 183.400 150.400 ;
        RECT 188.800 149.800 189.600 150.000 ;
        RECT 192.600 149.800 194.000 150.400 ;
        RECT 188.800 149.200 191.400 149.800 ;
        RECT 174.000 148.200 176.600 149.000 ;
        RECT 177.400 148.200 179.800 149.000 ;
        RECT 180.800 148.200 183.400 149.000 ;
        RECT 190.800 148.600 191.400 149.200 ;
        RECT 192.200 149.600 194.000 149.800 ;
        RECT 200.200 149.800 201.800 150.400 ;
        RECT 202.800 150.300 203.600 150.400 ;
        RECT 209.300 150.300 209.900 151.600 ;
        RECT 200.200 149.600 201.000 149.800 ;
        RECT 202.800 149.700 209.900 150.300 ;
        RECT 202.800 149.600 203.600 149.700 ;
        RECT 192.200 149.200 193.200 149.600 ;
        RECT 175.800 147.600 176.600 148.200 ;
        RECT 179.000 147.600 179.800 148.200 ;
        RECT 182.600 147.600 183.400 148.200 ;
        RECT 186.800 148.200 188.400 148.400 ;
        RECT 186.800 147.600 190.200 148.200 ;
        RECT 190.800 147.800 191.600 148.600 ;
        RECT 172.400 146.800 174.800 147.600 ;
        RECT 175.800 146.800 178.000 147.600 ;
        RECT 179.000 146.800 181.200 147.600 ;
        RECT 182.600 146.800 184.400 147.600 ;
        RECT 189.600 147.200 190.200 147.600 ;
        RECT 188.200 146.800 189.000 147.000 ;
        RECT 167.800 146.400 168.600 146.600 ;
        RECT 156.400 144.200 157.200 145.000 ;
        RECT 158.000 144.800 158.800 145.600 ;
        RECT 159.800 145.400 160.600 145.600 ;
        RECT 159.800 144.800 162.600 145.400 ;
        RECT 162.000 144.200 162.600 144.800 ;
        RECT 166.000 144.200 166.800 145.000 ;
        RECT 156.400 143.600 158.400 144.200 ;
        RECT 157.600 142.200 158.400 143.600 ;
        RECT 162.000 142.200 162.800 144.200 ;
        RECT 166.000 143.600 167.400 144.200 ;
        RECT 166.200 142.200 167.400 143.600 ;
        RECT 170.800 142.200 171.600 146.600 ;
        RECT 174.000 142.200 174.800 146.800 ;
        RECT 177.200 142.200 178.000 146.800 ;
        RECT 180.400 142.200 181.200 146.800 ;
        RECT 183.600 142.200 184.400 146.800 ;
        RECT 186.800 146.200 189.000 146.800 ;
        RECT 189.600 146.600 191.600 147.200 ;
        RECT 190.000 146.400 191.600 146.600 ;
        RECT 186.800 142.200 187.600 146.200 ;
        RECT 192.200 145.800 192.800 149.200 ;
        RECT 201.600 148.600 202.400 148.800 ;
        RECT 199.600 148.400 202.400 148.600 ;
        RECT 193.600 147.600 194.400 148.400 ;
        RECT 195.600 147.600 197.200 148.400 ;
        RECT 198.000 148.000 202.400 148.400 ;
        RECT 203.000 148.400 203.600 149.600 ;
        RECT 198.000 147.800 200.200 148.000 ;
        RECT 203.000 147.800 204.000 148.400 ;
        RECT 198.000 147.600 199.600 147.800 ;
        RECT 193.600 147.200 194.200 147.600 ;
        RECT 193.400 146.400 194.200 147.200 ;
        RECT 194.800 146.800 195.600 147.000 ;
        RECT 199.800 146.800 200.600 147.000 ;
        RECT 194.800 146.200 197.200 146.800 ;
        RECT 191.200 144.400 192.800 145.800 ;
        RECT 191.200 143.600 194.000 144.400 ;
        RECT 191.200 142.200 192.800 143.600 ;
        RECT 196.400 142.200 197.200 146.200 ;
        RECT 198.000 146.200 200.600 146.800 ;
        RECT 201.200 146.400 202.800 147.200 ;
        RECT 198.000 142.200 198.800 146.200 ;
        RECT 203.400 145.800 204.000 147.800 ;
        RECT 204.800 147.600 205.600 148.400 ;
        RECT 206.800 147.600 208.400 148.400 ;
        RECT 204.800 147.200 205.400 147.600 ;
        RECT 204.600 146.400 205.400 147.200 ;
        RECT 206.000 146.800 206.800 147.000 ;
        RECT 206.000 146.200 208.400 146.800 ;
        RECT 210.800 146.200 211.600 159.800 ;
        RECT 214.000 152.400 214.800 159.800 ;
        RECT 215.600 152.400 216.400 152.600 ;
        RECT 214.000 151.800 216.400 152.400 ;
        RECT 218.400 151.800 220.000 159.800 ;
        RECT 221.800 152.400 222.600 152.600 ;
        RECT 223.600 152.400 224.400 159.800 ;
        RECT 221.800 151.800 224.400 152.400 ;
        RECT 225.800 152.600 226.600 159.800 ;
        RECT 225.800 151.800 227.600 152.600 ;
        RECT 218.800 150.400 219.400 151.800 ;
        RECT 220.600 150.400 221.400 150.600 ;
        RECT 218.800 149.600 219.600 150.400 ;
        RECT 220.600 149.800 222.200 150.400 ;
        RECT 221.400 149.600 222.200 149.800 ;
        RECT 225.200 149.600 226.000 151.200 ;
        RECT 218.800 148.400 219.400 149.600 ;
        RECT 212.400 146.800 213.200 148.400 ;
        RECT 214.000 147.600 215.600 148.400 ;
        RECT 216.800 147.600 217.600 148.400 ;
        RECT 217.000 147.200 217.600 147.600 ;
        RECT 218.400 147.800 219.400 148.400 ;
        RECT 220.000 148.600 220.800 148.800 ;
        RECT 220.000 148.400 222.800 148.600 ;
        RECT 226.800 148.400 227.400 151.800 ;
        RECT 220.000 148.000 224.400 148.400 ;
        RECT 222.200 147.800 224.400 148.000 ;
        RECT 215.600 146.800 216.400 147.000 ;
        RECT 202.400 142.200 204.000 145.800 ;
        RECT 207.600 142.200 208.400 146.200 ;
        RECT 209.800 145.600 211.600 146.200 ;
        RECT 214.000 146.200 216.400 146.800 ;
        RECT 217.000 146.400 217.800 147.200 ;
        RECT 209.800 144.400 210.600 145.600 ;
        RECT 209.200 143.600 210.600 144.400 ;
        RECT 209.800 142.200 210.600 143.600 ;
        RECT 214.000 142.200 214.800 146.200 ;
        RECT 218.400 145.800 219.000 147.800 ;
        RECT 222.800 147.600 224.400 147.800 ;
        RECT 226.800 147.600 227.600 148.400 ;
        RECT 219.600 146.400 221.200 147.200 ;
        RECT 221.800 146.800 222.600 147.000 ;
        RECT 221.800 146.200 224.400 146.800 ;
        RECT 218.400 144.400 220.000 145.800 ;
        RECT 218.400 143.600 221.200 144.400 ;
        RECT 218.400 142.200 220.000 143.600 ;
        RECT 223.600 142.200 224.400 146.200 ;
        RECT 226.800 144.400 227.400 147.600 ;
        RECT 228.400 144.800 229.200 146.400 ;
        RECT 226.800 142.200 227.600 144.400 ;
        RECT 230.000 142.200 230.800 159.800 ;
        RECT 233.200 152.400 234.000 159.800 ;
        RECT 237.600 154.400 239.200 159.800 ;
        RECT 237.600 153.600 240.400 154.400 ;
        RECT 234.800 152.400 235.600 152.600 ;
        RECT 237.600 152.400 239.200 153.600 ;
        RECT 233.200 151.800 235.600 152.400 ;
        RECT 237.200 151.800 239.200 152.400 ;
        RECT 241.400 152.400 242.200 152.600 ;
        RECT 242.800 152.400 243.600 159.800 ;
        RECT 241.400 151.800 243.600 152.400 ;
        RECT 237.200 150.400 237.800 151.800 ;
        RECT 241.400 151.200 242.000 151.800 ;
        RECT 238.600 150.600 242.000 151.200 ;
        RECT 244.400 151.200 245.200 159.800 ;
        RECT 248.600 152.400 249.400 159.800 ;
        RECT 248.600 152.300 250.000 152.400 ;
        RECT 250.800 152.300 251.600 153.200 ;
        RECT 248.600 151.800 251.600 152.300 ;
        RECT 249.300 151.700 251.600 151.800 ;
        RECT 244.400 150.800 248.400 151.200 ;
        RECT 244.400 150.600 248.600 150.800 ;
        RECT 238.600 150.400 239.400 150.600 ;
        RECT 236.400 149.800 237.800 150.400 ;
        RECT 247.800 150.000 248.600 150.600 ;
        RECT 249.400 150.400 250.000 151.700 ;
        RECT 250.800 151.600 251.600 151.700 ;
        RECT 240.800 149.800 241.600 150.000 ;
        RECT 236.400 149.600 238.200 149.800 ;
        RECT 237.200 149.200 238.200 149.600 ;
        RECT 231.600 148.300 232.400 148.400 ;
        RECT 233.200 148.300 234.800 148.400 ;
        RECT 231.600 147.700 234.800 148.300 ;
        RECT 231.600 147.600 232.400 147.700 ;
        RECT 233.200 147.600 234.800 147.700 ;
        RECT 236.000 147.600 236.800 148.400 ;
        RECT 236.200 147.200 236.800 147.600 ;
        RECT 234.800 146.800 235.600 147.000 ;
        RECT 231.600 144.800 232.400 146.400 ;
        RECT 233.200 146.200 235.600 146.800 ;
        RECT 236.200 146.400 237.000 147.200 ;
        RECT 233.200 142.200 234.000 146.200 ;
        RECT 237.600 145.800 238.200 149.200 ;
        RECT 239.000 149.200 241.600 149.800 ;
        RECT 239.000 148.600 239.600 149.200 ;
        RECT 238.800 147.800 239.600 148.600 ;
        RECT 246.400 148.400 247.200 149.200 ;
        RECT 242.000 148.200 243.600 148.400 ;
        RECT 240.200 147.600 243.600 148.200 ;
        RECT 246.000 147.600 247.000 148.400 ;
        RECT 240.200 147.200 240.800 147.600 ;
        RECT 238.800 146.600 240.800 147.200 ;
        RECT 248.000 147.000 248.600 150.000 ;
        RECT 249.200 149.600 250.000 150.400 ;
        RECT 241.400 146.800 242.200 147.000 ;
        RECT 238.800 146.400 240.400 146.600 ;
        RECT 241.400 146.200 243.600 146.800 ;
        RECT 246.200 146.400 248.600 147.000 ;
        RECT 237.600 142.200 239.200 145.800 ;
        RECT 242.800 142.200 243.600 146.200 ;
        RECT 244.400 144.800 245.200 146.400 ;
        RECT 246.200 144.200 246.800 146.400 ;
        RECT 249.400 146.200 250.000 149.600 ;
        RECT 252.400 146.200 253.200 159.800 ;
        RECT 255.600 151.600 256.400 153.200 ;
        RECT 254.000 148.300 254.800 148.400 ;
        RECT 257.200 148.300 258.000 159.800 ;
        RECT 263.000 152.600 263.800 159.800 ;
        RECT 266.800 155.800 267.600 159.800 ;
        RECT 262.000 151.800 263.800 152.600 ;
        RECT 262.200 148.400 262.800 151.800 ;
        RECT 267.000 151.600 267.600 155.800 ;
        RECT 270.000 151.800 270.800 159.800 ;
        RECT 272.400 153.600 273.200 154.400 ;
        RECT 272.400 152.400 273.000 153.600 ;
        RECT 273.800 152.400 274.600 159.800 ;
        RECT 263.600 149.600 264.400 151.200 ;
        RECT 267.000 151.000 269.400 151.600 ;
        RECT 266.800 149.600 267.600 150.400 ;
        RECT 254.000 147.700 258.000 148.300 ;
        RECT 254.000 146.800 254.800 147.700 ;
        RECT 257.200 146.200 258.000 147.700 ;
        RECT 258.800 148.300 259.600 148.400 ;
        RECT 258.800 147.700 261.100 148.300 ;
        RECT 258.800 146.800 259.600 147.700 ;
        RECT 260.500 146.400 261.100 147.700 ;
        RECT 262.000 147.600 262.800 148.400 ;
        RECT 265.200 147.600 266.000 149.200 ;
        RECT 267.000 148.800 267.600 149.600 ;
        RECT 267.000 148.200 268.000 148.800 ;
        RECT 267.200 148.000 268.000 148.200 ;
        RECT 268.800 147.600 269.400 151.000 ;
        RECT 270.200 150.400 270.800 151.800 ;
        RECT 271.600 151.800 273.000 152.400 ;
        RECT 273.600 151.800 274.600 152.400 ;
        RECT 278.000 152.400 278.800 159.800 ;
        RECT 279.600 152.400 280.400 152.600 ;
        RECT 282.400 152.400 284.000 159.800 ;
        RECT 278.000 151.800 280.400 152.400 ;
        RECT 282.000 151.800 284.000 152.400 ;
        RECT 286.200 152.400 287.000 152.600 ;
        RECT 287.600 152.400 288.400 159.800 ;
        RECT 286.200 151.800 288.400 152.400 ;
        RECT 271.600 151.600 272.400 151.800 ;
        RECT 270.000 149.600 270.800 150.400 ;
        RECT 246.000 142.200 246.800 144.200 ;
        RECT 249.200 142.200 250.000 146.200 ;
        RECT 251.400 145.600 253.200 146.200 ;
        RECT 256.200 145.600 258.000 146.200 ;
        RECT 251.400 144.400 252.200 145.600 ;
        RECT 250.800 143.600 252.200 144.400 ;
        RECT 251.400 142.200 252.200 143.600 ;
        RECT 256.200 142.200 257.000 145.600 ;
        RECT 260.400 144.800 261.200 146.400 ;
        RECT 262.200 146.300 262.800 147.600 ;
        RECT 268.800 147.400 269.600 147.600 ;
        RECT 266.600 147.000 269.600 147.400 ;
        RECT 265.400 146.800 269.600 147.000 ;
        RECT 265.400 146.400 267.200 146.800 ;
        RECT 263.600 146.300 264.400 146.400 ;
        RECT 262.100 145.700 264.400 146.300 ;
        RECT 265.400 146.200 266.000 146.400 ;
        RECT 270.200 146.200 270.800 149.600 ;
        RECT 273.600 148.400 274.200 151.800 ;
        RECT 282.000 150.400 282.600 151.800 ;
        RECT 286.200 151.200 286.800 151.800 ;
        RECT 283.400 150.600 286.800 151.200 ;
        RECT 294.000 151.400 294.800 159.800 ;
        RECT 298.400 156.400 299.200 159.800 ;
        RECT 297.200 155.800 299.200 156.400 ;
        RECT 302.800 155.800 303.600 159.800 ;
        RECT 307.000 155.800 308.200 159.800 ;
        RECT 297.200 155.000 298.000 155.800 ;
        RECT 302.800 155.200 303.400 155.800 ;
        RECT 300.600 154.600 304.200 155.200 ;
        RECT 306.800 155.000 307.600 155.800 ;
        RECT 300.600 154.400 301.400 154.600 ;
        RECT 303.400 154.400 304.200 154.600 ;
        RECT 307.800 154.000 309.200 154.400 ;
        RECT 307.000 153.600 309.200 154.000 ;
        RECT 297.200 153.000 298.000 153.200 ;
        RECT 301.800 153.000 302.600 153.200 ;
        RECT 297.200 152.400 302.600 153.000 ;
        RECT 303.200 153.000 305.400 153.600 ;
        RECT 303.200 151.800 303.800 153.000 ;
        RECT 304.600 152.800 305.400 153.000 ;
        RECT 307.000 153.200 308.400 153.600 ;
        RECT 307.000 152.200 307.600 153.200 ;
        RECT 299.000 151.400 303.800 151.800 ;
        RECT 294.000 151.200 303.800 151.400 ;
        RECT 305.200 151.600 307.600 152.200 ;
        RECT 294.000 151.000 299.800 151.200 ;
        RECT 294.000 150.800 299.600 151.000 ;
        RECT 283.400 150.400 284.200 150.600 ;
        RECT 305.200 150.400 305.800 151.600 ;
        RECT 311.600 151.200 312.400 159.800 ;
        RECT 308.200 150.600 312.400 151.200 ;
        RECT 313.200 151.400 314.000 159.800 ;
        RECT 317.600 156.400 318.400 159.800 ;
        RECT 316.400 155.800 318.400 156.400 ;
        RECT 322.000 155.800 322.800 159.800 ;
        RECT 326.200 155.800 327.400 159.800 ;
        RECT 316.400 155.000 317.200 155.800 ;
        RECT 322.000 155.200 322.600 155.800 ;
        RECT 319.800 154.600 323.400 155.200 ;
        RECT 326.000 155.000 326.800 155.800 ;
        RECT 319.800 154.400 320.600 154.600 ;
        RECT 322.600 154.400 323.400 154.600 ;
        RECT 316.400 153.000 317.200 153.200 ;
        RECT 321.000 153.000 321.800 153.200 ;
        RECT 316.400 152.400 321.800 153.000 ;
        RECT 322.400 153.000 324.600 153.600 ;
        RECT 322.400 151.800 323.000 153.000 ;
        RECT 323.800 152.800 324.600 153.000 ;
        RECT 326.200 153.200 327.600 154.000 ;
        RECT 326.200 152.200 326.800 153.200 ;
        RECT 318.200 151.400 323.000 151.800 ;
        RECT 313.200 151.200 323.000 151.400 ;
        RECT 324.400 151.600 326.800 152.200 ;
        RECT 313.200 151.000 319.000 151.200 ;
        RECT 313.200 150.800 318.800 151.000 ;
        RECT 308.200 150.400 309.000 150.600 ;
        RECT 274.800 148.800 275.600 150.400 ;
        RECT 281.200 149.800 282.600 150.400 ;
        RECT 300.400 150.200 301.200 150.400 ;
        RECT 285.600 149.800 286.400 150.000 ;
        RECT 281.200 149.600 283.000 149.800 ;
        RECT 282.000 149.200 283.000 149.600 ;
        RECT 271.600 147.600 274.200 148.400 ;
        RECT 276.400 148.200 277.200 148.400 ;
        RECT 275.600 147.600 277.200 148.200 ;
        RECT 278.000 147.600 279.600 148.400 ;
        RECT 280.800 147.600 281.600 148.400 ;
        RECT 271.800 146.200 272.400 147.600 ;
        RECT 275.600 147.200 276.400 147.600 ;
        RECT 281.000 147.200 281.600 147.600 ;
        RECT 279.600 146.800 280.400 147.000 ;
        RECT 273.400 146.200 277.000 146.600 ;
        RECT 278.000 146.200 280.400 146.800 ;
        RECT 281.000 146.400 281.800 147.200 ;
        RECT 262.200 144.200 262.800 145.700 ;
        RECT 263.600 145.600 264.400 145.700 ;
        RECT 262.000 142.200 262.800 144.200 ;
        RECT 265.200 142.200 266.000 146.200 ;
        RECT 269.400 145.200 270.800 146.200 ;
        RECT 269.400 142.200 270.200 145.200 ;
        RECT 271.600 142.200 272.400 146.200 ;
        RECT 273.200 146.000 277.200 146.200 ;
        RECT 273.200 142.200 274.000 146.000 ;
        RECT 276.400 142.200 277.200 146.000 ;
        RECT 278.000 142.200 278.800 146.200 ;
        RECT 282.400 145.800 283.000 149.200 ;
        RECT 283.800 149.200 286.400 149.800 ;
        RECT 296.200 149.600 301.200 150.200 ;
        RECT 305.200 149.600 306.000 150.400 ;
        RECT 309.800 149.800 310.600 150.000 ;
        RECT 296.200 149.400 297.000 149.600 ;
        RECT 298.800 149.400 299.600 149.600 ;
        RECT 283.800 148.600 284.400 149.200 ;
        RECT 283.600 147.800 284.400 148.600 ;
        RECT 297.800 148.400 298.600 148.600 ;
        RECT 305.200 148.400 305.800 149.600 ;
        RECT 306.800 149.200 310.600 149.800 ;
        RECT 306.800 149.000 307.600 149.200 ;
        RECT 286.800 148.200 288.400 148.400 ;
        RECT 285.000 147.600 288.400 148.200 ;
        RECT 294.800 147.800 305.800 148.400 ;
        RECT 294.800 147.600 296.400 147.800 ;
        RECT 285.000 147.200 285.600 147.600 ;
        RECT 283.600 146.600 285.600 147.200 ;
        RECT 286.200 146.800 287.000 147.000 ;
        RECT 283.600 146.400 285.200 146.600 ;
        RECT 286.200 146.200 288.400 146.800 ;
        RECT 282.400 142.200 284.000 145.800 ;
        RECT 287.600 142.200 288.400 146.200 ;
        RECT 294.000 142.200 294.800 147.000 ;
        RECT 299.000 145.600 299.600 147.800 ;
        RECT 304.600 147.600 305.400 147.800 ;
        RECT 311.600 147.200 312.400 150.600 ;
        RECT 319.600 150.200 320.400 150.400 ;
        RECT 315.400 149.600 320.400 150.200 ;
        RECT 315.400 149.400 316.200 149.600 ;
        RECT 318.000 149.400 318.800 149.600 ;
        RECT 317.000 148.400 317.800 148.600 ;
        RECT 324.400 148.400 325.000 151.600 ;
        RECT 330.800 151.200 331.600 159.800 ;
        RECT 327.400 150.600 331.600 151.200 ;
        RECT 327.400 150.400 328.200 150.600 ;
        RECT 329.000 149.800 329.800 150.000 ;
        RECT 326.000 149.200 329.800 149.800 ;
        RECT 326.000 149.000 326.800 149.200 ;
        RECT 314.000 147.800 325.000 148.400 ;
        RECT 314.000 147.600 315.600 147.800 ;
        RECT 308.600 146.600 312.400 147.200 ;
        RECT 308.600 146.400 309.400 146.600 ;
        RECT 297.200 144.200 298.000 145.000 ;
        RECT 298.800 144.800 299.600 145.600 ;
        RECT 300.600 145.400 301.400 145.600 ;
        RECT 300.600 144.800 303.400 145.400 ;
        RECT 302.800 144.200 303.400 144.800 ;
        RECT 306.800 144.200 307.600 145.000 ;
        RECT 297.200 143.600 299.200 144.200 ;
        RECT 298.400 142.200 299.200 143.600 ;
        RECT 302.800 142.200 303.600 144.200 ;
        RECT 306.800 143.600 308.200 144.200 ;
        RECT 307.000 142.200 308.200 143.600 ;
        RECT 311.600 142.200 312.400 146.600 ;
        RECT 313.200 142.200 314.000 147.000 ;
        RECT 318.200 145.600 318.800 147.800 ;
        RECT 323.800 147.600 324.600 147.800 ;
        RECT 330.800 147.200 331.600 150.600 ;
        RECT 334.000 151.200 334.800 159.800 ;
        RECT 337.200 151.200 338.000 159.800 ;
        RECT 340.400 151.200 341.200 159.800 ;
        RECT 343.600 151.200 344.400 159.800 ;
        RECT 349.400 152.400 350.200 159.800 ;
        RECT 355.400 158.400 356.200 159.800 ;
        RECT 355.400 157.600 357.200 158.400 ;
        RECT 350.800 153.600 351.600 154.400 ;
        RECT 351.000 152.400 351.600 153.600 ;
        RECT 354.000 153.600 354.800 154.400 ;
        RECT 354.000 152.400 354.600 153.600 ;
        RECT 355.400 152.400 356.200 157.600 ;
        RECT 349.400 151.800 350.400 152.400 ;
        RECT 351.000 151.800 352.400 152.400 ;
        RECT 334.000 150.400 335.800 151.200 ;
        RECT 337.200 150.400 339.400 151.200 ;
        RECT 340.400 150.400 342.600 151.200 ;
        RECT 343.600 150.400 346.000 151.200 ;
        RECT 335.000 149.000 335.800 150.400 ;
        RECT 338.600 149.000 339.400 150.400 ;
        RECT 341.800 149.000 342.600 150.400 ;
        RECT 335.000 148.200 337.600 149.000 ;
        RECT 338.600 148.200 341.000 149.000 ;
        RECT 341.800 148.200 344.400 149.000 ;
        RECT 335.000 147.600 335.800 148.200 ;
        RECT 338.600 147.600 339.400 148.200 ;
        RECT 341.800 147.600 342.600 148.200 ;
        RECT 345.200 147.600 346.000 150.400 ;
        RECT 348.400 148.800 349.200 150.400 ;
        RECT 349.800 150.300 350.400 151.800 ;
        RECT 351.600 151.600 352.400 151.800 ;
        RECT 353.200 151.800 354.600 152.400 ;
        RECT 355.200 151.800 356.200 152.400 ;
        RECT 353.200 151.600 354.000 151.800 ;
        RECT 353.300 150.300 353.900 151.600 ;
        RECT 349.800 149.700 353.900 150.300 ;
        RECT 349.800 148.400 350.400 149.700 ;
        RECT 355.200 148.400 355.800 151.800 ;
        RECT 356.400 148.800 357.200 150.400 ;
        RECT 346.800 148.200 347.600 148.400 ;
        RECT 346.800 147.600 348.400 148.200 ;
        RECT 349.800 147.600 352.400 148.400 ;
        RECT 353.200 147.600 355.800 148.400 ;
        RECT 358.000 148.300 358.800 148.400 ;
        RECT 359.600 148.300 360.400 159.800 ;
        RECT 365.400 152.400 366.200 159.800 ;
        RECT 366.800 153.600 367.600 154.400 ;
        RECT 367.000 152.400 367.600 153.600 ;
        RECT 371.800 152.400 372.600 159.800 ;
        RECT 373.200 153.600 374.000 154.400 ;
        RECT 373.400 152.400 374.000 153.600 ;
        RECT 378.200 152.400 379.000 159.800 ;
        RECT 379.600 153.600 380.400 154.400 ;
        RECT 379.800 152.400 380.400 153.600 ;
        RECT 382.800 153.600 383.600 154.400 ;
        RECT 382.800 152.400 383.400 153.600 ;
        RECT 384.200 152.400 385.000 159.800 ;
        RECT 389.200 153.600 390.000 154.400 ;
        RECT 389.200 152.400 389.800 153.600 ;
        RECT 390.600 152.400 391.400 159.800 ;
        RECT 365.400 151.800 366.400 152.400 ;
        RECT 367.000 151.800 368.400 152.400 ;
        RECT 371.800 151.800 372.800 152.400 ;
        RECT 373.400 151.800 374.800 152.400 ;
        RECT 378.200 151.800 379.200 152.400 ;
        RECT 379.800 151.800 381.200 152.400 ;
        RECT 364.400 148.800 365.200 150.400 ;
        RECT 365.800 150.300 366.400 151.800 ;
        RECT 367.600 151.600 368.400 151.800 ;
        RECT 367.600 150.300 368.400 150.400 ;
        RECT 365.800 149.700 368.400 150.300 ;
        RECT 365.800 148.400 366.400 149.700 ;
        RECT 367.600 149.600 368.400 149.700 ;
        RECT 370.800 148.800 371.600 150.400 ;
        RECT 372.200 148.400 372.800 151.800 ;
        RECT 374.000 151.600 374.800 151.800 ;
        RECT 375.600 150.300 376.400 150.400 ;
        RECT 377.200 150.300 378.000 150.400 ;
        RECT 375.600 149.700 378.000 150.300 ;
        RECT 375.600 149.600 376.400 149.700 ;
        RECT 377.200 148.800 378.000 149.700 ;
        RECT 378.600 148.400 379.200 151.800 ;
        RECT 380.400 151.600 381.200 151.800 ;
        RECT 382.000 151.800 383.400 152.400 ;
        RECT 382.000 151.600 382.800 151.800 ;
        RECT 384.000 151.600 386.000 152.400 ;
        RECT 388.400 151.800 389.800 152.400 ;
        RECT 390.400 151.800 391.400 152.400 ;
        RECT 388.400 151.600 389.200 151.800 ;
        RECT 384.000 148.400 384.600 151.600 ;
        RECT 385.200 148.800 386.000 150.400 ;
        RECT 390.400 148.400 391.000 151.800 ;
        RECT 391.600 148.800 392.400 150.400 ;
        RECT 358.000 148.200 360.400 148.300 ;
        RECT 357.200 147.700 360.400 148.200 ;
        RECT 357.200 147.600 358.800 147.700 ;
        RECT 327.800 146.600 331.600 147.200 ;
        RECT 327.800 146.400 328.600 146.600 ;
        RECT 316.400 144.200 317.200 145.000 ;
        RECT 318.000 144.800 318.800 145.600 ;
        RECT 319.800 145.400 320.600 145.600 ;
        RECT 319.800 144.800 322.600 145.400 ;
        RECT 322.000 144.200 322.600 144.800 ;
        RECT 326.000 144.200 326.800 145.000 ;
        RECT 316.400 143.600 318.400 144.200 ;
        RECT 317.600 142.200 318.400 143.600 ;
        RECT 322.000 142.200 322.800 144.200 ;
        RECT 326.000 143.600 327.400 144.200 ;
        RECT 326.200 142.200 327.400 143.600 ;
        RECT 330.800 142.200 331.600 146.600 ;
        RECT 334.000 146.800 335.800 147.600 ;
        RECT 337.200 146.800 339.400 147.600 ;
        RECT 340.400 146.800 342.600 147.600 ;
        RECT 343.600 146.800 346.000 147.600 ;
        RECT 347.600 147.200 348.400 147.600 ;
        RECT 334.000 142.200 334.800 146.800 ;
        RECT 337.200 142.200 338.000 146.800 ;
        RECT 340.400 142.200 341.200 146.800 ;
        RECT 343.600 142.200 344.400 146.800 ;
        RECT 347.000 146.200 350.600 146.600 ;
        RECT 351.600 146.200 352.200 147.600 ;
        RECT 353.400 146.200 354.000 147.600 ;
        RECT 357.200 147.200 358.000 147.600 ;
        RECT 355.000 146.200 358.600 146.600 ;
        RECT 346.800 146.000 350.800 146.200 ;
        RECT 346.800 142.200 347.600 146.000 ;
        RECT 350.000 142.200 350.800 146.000 ;
        RECT 351.600 142.200 352.400 146.200 ;
        RECT 353.200 142.200 354.000 146.200 ;
        RECT 354.800 146.000 358.800 146.200 ;
        RECT 354.800 142.200 355.600 146.000 ;
        RECT 358.000 142.200 358.800 146.000 ;
        RECT 359.600 142.200 360.400 147.700 ;
        RECT 362.800 148.200 363.600 148.400 ;
        RECT 362.800 147.600 364.400 148.200 ;
        RECT 365.800 147.600 368.400 148.400 ;
        RECT 369.200 148.200 370.000 148.400 ;
        RECT 369.200 147.600 370.800 148.200 ;
        RECT 372.200 147.600 374.800 148.400 ;
        RECT 375.600 148.200 376.400 148.400 ;
        RECT 375.600 147.600 377.200 148.200 ;
        RECT 378.600 147.600 381.200 148.400 ;
        RECT 382.000 147.600 384.600 148.400 ;
        RECT 386.800 148.200 387.600 148.400 ;
        RECT 386.000 147.600 387.600 148.200 ;
        RECT 388.400 147.600 391.000 148.400 ;
        RECT 393.200 148.200 394.000 148.400 ;
        RECT 392.400 147.600 394.000 148.200 ;
        RECT 396.400 148.300 397.200 159.800 ;
        RECT 398.000 159.200 402.000 159.800 ;
        RECT 398.000 151.800 398.800 159.200 ;
        RECT 399.600 151.800 400.400 158.600 ;
        RECT 401.200 152.400 402.000 159.200 ;
        RECT 404.400 152.400 405.200 159.800 ;
        RECT 401.200 151.800 405.200 152.400 ;
        RECT 406.000 152.400 406.800 159.800 ;
        RECT 409.200 159.200 413.200 159.800 ;
        RECT 409.200 152.400 410.000 159.200 ;
        RECT 406.000 151.800 410.000 152.400 ;
        RECT 410.800 151.800 411.600 158.600 ;
        RECT 412.400 151.800 413.200 159.200 ;
        RECT 414.000 155.000 414.800 159.000 ;
        RECT 418.200 158.400 419.000 159.800 ;
        RECT 418.200 157.600 419.600 158.400 ;
        RECT 399.800 151.200 400.400 151.800 ;
        RECT 410.800 151.200 411.400 151.800 ;
        RECT 414.000 151.600 414.600 155.000 ;
        RECT 418.200 152.800 419.000 157.600 ;
        RECT 418.200 152.200 419.800 152.800 ;
        RECT 398.000 149.600 398.800 151.200 ;
        RECT 399.800 150.600 401.800 151.200 ;
        RECT 401.200 150.400 401.800 150.600 ;
        RECT 403.600 150.400 404.400 150.800 ;
        RECT 406.800 150.400 407.600 150.800 ;
        RECT 409.400 150.600 411.400 151.200 ;
        RECT 409.400 150.400 410.000 150.600 ;
        RECT 401.200 149.600 402.000 150.400 ;
        RECT 403.600 149.800 405.200 150.400 ;
        RECT 404.400 149.600 405.200 149.800 ;
        RECT 406.000 149.800 407.600 150.400 ;
        RECT 406.000 149.600 406.800 149.800 ;
        RECT 409.200 149.600 410.000 150.400 ;
        RECT 412.400 149.600 413.200 151.200 ;
        RECT 414.000 151.000 417.800 151.600 ;
        RECT 399.800 148.800 400.600 149.600 ;
        RECT 399.800 148.400 400.400 148.800 ;
        RECT 399.600 148.300 400.400 148.400 ;
        RECT 396.400 147.700 400.400 148.300 ;
        RECT 363.600 147.200 364.400 147.600 ;
        RECT 361.200 144.800 362.000 146.400 ;
        RECT 363.000 146.200 366.600 146.600 ;
        RECT 367.600 146.200 368.200 147.600 ;
        RECT 370.000 147.200 370.800 147.600 ;
        RECT 369.400 146.200 373.000 146.600 ;
        RECT 374.000 146.400 374.600 147.600 ;
        RECT 376.400 147.200 377.200 147.600 ;
        RECT 362.800 146.000 366.800 146.200 ;
        RECT 362.800 142.200 363.600 146.000 ;
        RECT 366.000 142.200 366.800 146.000 ;
        RECT 367.600 142.200 368.400 146.200 ;
        RECT 369.200 146.000 373.200 146.200 ;
        RECT 369.200 142.200 370.000 146.000 ;
        RECT 372.400 142.200 373.200 146.000 ;
        RECT 374.000 142.200 374.800 146.400 ;
        RECT 375.800 146.200 379.400 146.600 ;
        RECT 380.400 146.200 381.000 147.600 ;
        RECT 382.200 146.200 382.800 147.600 ;
        RECT 386.000 147.200 386.800 147.600 ;
        RECT 383.800 146.200 387.400 146.600 ;
        RECT 388.600 146.200 389.200 147.600 ;
        RECT 392.400 147.200 393.200 147.600 ;
        RECT 390.200 146.200 393.800 146.600 ;
        RECT 375.600 146.000 379.600 146.200 ;
        RECT 375.600 142.200 376.400 146.000 ;
        RECT 378.800 142.200 379.600 146.000 ;
        RECT 380.400 142.200 381.200 146.200 ;
        RECT 382.000 142.200 382.800 146.200 ;
        RECT 383.600 146.000 387.600 146.200 ;
        RECT 383.600 142.200 384.400 146.000 ;
        RECT 386.800 142.200 387.600 146.000 ;
        RECT 388.400 142.200 389.200 146.200 ;
        RECT 390.000 146.000 394.000 146.200 ;
        RECT 390.000 142.200 390.800 146.000 ;
        RECT 393.200 142.200 394.000 146.000 ;
        RECT 394.800 144.800 395.600 146.400 ;
        RECT 396.400 142.200 397.200 147.700 ;
        RECT 399.600 147.600 400.400 147.700 ;
        RECT 401.200 146.200 401.800 149.600 ;
        RECT 402.800 148.300 403.600 149.200 ;
        RECT 407.600 148.300 408.400 149.200 ;
        RECT 402.800 147.700 408.400 148.300 ;
        RECT 402.800 147.600 403.600 147.700 ;
        RECT 407.600 147.600 408.400 147.700 ;
        RECT 409.400 146.400 410.000 149.600 ;
        RECT 410.600 148.800 411.400 149.600 ;
        RECT 414.000 148.800 414.800 150.400 ;
        RECT 415.600 148.800 416.400 150.400 ;
        RECT 417.200 149.000 417.800 151.000 ;
        RECT 410.800 148.400 411.400 148.800 ;
        RECT 410.800 147.600 411.600 148.400 ;
        RECT 417.200 148.200 418.600 149.000 ;
        RECT 419.200 148.400 419.800 152.200 ;
        RECT 423.600 152.400 424.400 159.800 ;
        RECT 426.800 152.400 427.600 159.800 ;
        RECT 423.600 151.800 427.600 152.400 ;
        RECT 428.400 151.800 429.200 159.800 ;
        RECT 420.400 150.300 421.200 151.200 ;
        RECT 424.400 150.400 425.200 150.800 ;
        RECT 428.400 150.400 429.000 151.800 ;
        RECT 423.600 150.300 425.200 150.400 ;
        RECT 420.400 149.800 425.200 150.300 ;
        RECT 426.800 149.800 429.200 150.400 ;
        RECT 420.400 149.700 424.400 149.800 ;
        RECT 420.400 149.600 421.200 149.700 ;
        RECT 423.600 149.600 424.400 149.700 ;
        RECT 417.200 147.800 418.200 148.200 ;
        RECT 414.000 147.200 418.200 147.800 ;
        RECT 419.200 147.600 421.200 148.400 ;
        RECT 425.200 147.600 426.000 149.200 ;
        RECT 409.400 146.200 411.600 146.400 ;
        RECT 400.600 144.400 402.200 146.200 ;
        RECT 399.600 143.600 402.200 144.400 ;
        RECT 400.600 142.200 402.200 143.600 ;
        RECT 409.000 145.600 411.600 146.200 ;
        RECT 409.000 142.200 410.600 145.600 ;
        RECT 414.000 145.000 414.600 147.200 ;
        RECT 419.200 147.000 419.800 147.600 ;
        RECT 419.000 146.600 419.800 147.000 ;
        RECT 418.200 146.000 419.800 146.600 ;
        RECT 426.800 146.200 427.400 149.800 ;
        RECT 428.400 149.600 429.200 149.800 ;
        RECT 428.400 148.300 429.200 148.400 ;
        RECT 430.000 148.300 430.800 159.800 ;
        RECT 428.400 147.700 430.800 148.300 ;
        RECT 428.400 147.600 429.200 147.700 ;
        RECT 414.000 143.000 414.800 145.000 ;
        RECT 418.200 143.000 419.000 146.000 ;
        RECT 426.800 142.200 427.600 146.200 ;
        RECT 428.400 145.600 429.200 146.400 ;
        RECT 428.200 144.800 429.000 145.600 ;
        RECT 430.000 142.200 430.800 147.700 ;
        RECT 434.800 152.300 435.600 159.800 ;
        RECT 437.200 153.600 438.000 154.400 ;
        RECT 437.200 152.400 437.800 153.600 ;
        RECT 438.600 152.400 439.400 159.800 ;
        RECT 436.400 152.300 437.800 152.400 ;
        RECT 434.800 151.800 437.800 152.300 ;
        RECT 438.400 151.800 439.400 152.400 ;
        RECT 434.800 151.700 437.200 151.800 ;
        RECT 431.600 144.800 432.400 146.400 ;
        RECT 433.200 144.800 434.000 146.400 ;
        RECT 434.800 142.200 435.600 151.700 ;
        RECT 436.400 151.600 437.200 151.700 ;
        RECT 438.400 148.400 439.000 151.800 ;
        RECT 439.600 148.800 440.400 150.400 ;
        RECT 436.400 147.600 439.000 148.400 ;
        RECT 441.200 148.300 442.000 148.400 ;
        RECT 444.400 148.300 445.200 148.400 ;
        RECT 441.200 148.200 445.200 148.300 ;
        RECT 440.400 147.700 445.200 148.200 ;
        RECT 440.400 147.600 442.000 147.700 ;
        RECT 444.400 147.600 445.200 147.700 ;
        RECT 447.600 148.300 448.400 159.800 ;
        RECT 450.800 152.400 451.600 159.800 ;
        RECT 454.000 152.400 454.800 159.800 ;
        RECT 450.800 151.800 454.800 152.400 ;
        RECT 455.600 151.800 456.400 159.800 ;
        RECT 459.800 152.400 460.600 159.800 ;
        RECT 461.200 153.600 462.000 154.400 ;
        RECT 461.400 152.400 462.000 153.600 ;
        RECT 459.800 151.800 460.800 152.400 ;
        RECT 461.400 151.800 462.800 152.400 ;
        RECT 451.600 150.400 452.400 150.800 ;
        RECT 455.600 150.400 456.200 151.800 ;
        RECT 450.800 149.800 452.400 150.400 ;
        RECT 454.000 149.800 456.400 150.400 ;
        RECT 450.800 149.600 451.600 149.800 ;
        RECT 452.400 148.300 453.200 149.200 ;
        RECT 447.600 147.700 453.200 148.300 ;
        RECT 436.600 146.200 437.200 147.600 ;
        RECT 440.400 147.200 441.200 147.600 ;
        RECT 438.200 146.200 441.800 146.600 ;
        RECT 436.400 142.200 437.200 146.200 ;
        RECT 438.000 146.000 442.000 146.200 ;
        RECT 438.000 142.200 438.800 146.000 ;
        RECT 441.200 142.200 442.000 146.000 ;
        RECT 447.600 142.200 448.400 147.700 ;
        RECT 452.400 147.600 453.200 147.700 ;
        RECT 454.000 148.300 454.600 149.800 ;
        RECT 455.600 149.600 456.400 149.800 ;
        RECT 458.800 148.800 459.600 150.400 ;
        RECT 460.200 150.300 460.800 151.800 ;
        RECT 462.000 151.600 462.800 151.800 ;
        RECT 463.600 151.600 464.400 153.200 ;
        RECT 463.700 150.300 464.300 151.600 ;
        RECT 460.200 149.700 464.300 150.300 ;
        RECT 465.200 150.300 466.000 159.800 ;
        RECT 468.400 151.400 469.200 159.800 ;
        RECT 472.800 156.400 473.600 159.800 ;
        RECT 471.600 155.800 473.600 156.400 ;
        RECT 477.200 155.800 478.000 159.800 ;
        RECT 481.400 155.800 482.600 159.800 ;
        RECT 471.600 155.000 472.400 155.800 ;
        RECT 477.200 155.200 477.800 155.800 ;
        RECT 475.000 154.600 478.600 155.200 ;
        RECT 481.200 155.000 482.000 155.800 ;
        RECT 475.000 154.400 475.800 154.600 ;
        RECT 477.800 154.400 478.600 154.600 ;
        RECT 471.600 153.000 472.400 153.200 ;
        RECT 476.200 153.000 477.000 153.200 ;
        RECT 471.600 152.400 477.000 153.000 ;
        RECT 477.600 153.000 479.800 153.600 ;
        RECT 477.600 151.800 478.200 153.000 ;
        RECT 479.000 152.800 479.800 153.000 ;
        RECT 481.400 153.200 482.800 154.000 ;
        RECT 481.400 152.200 482.000 153.200 ;
        RECT 473.400 151.400 478.200 151.800 ;
        RECT 468.400 151.200 478.200 151.400 ;
        RECT 479.600 151.600 482.000 152.200 ;
        RECT 468.400 151.000 474.200 151.200 ;
        RECT 468.400 150.800 474.000 151.000 ;
        RECT 466.800 150.300 467.600 150.400 ;
        RECT 465.200 149.700 467.600 150.300 ;
        RECT 474.800 150.200 475.600 150.400 ;
        RECT 460.200 148.400 460.800 149.700 ;
        RECT 457.200 148.300 458.000 148.400 ;
        RECT 454.000 148.200 458.000 148.300 ;
        RECT 454.000 147.700 458.800 148.200 ;
        RECT 449.200 144.800 450.000 146.400 ;
        RECT 454.000 146.200 454.600 147.700 ;
        RECT 457.200 147.600 458.800 147.700 ;
        RECT 460.200 147.600 462.800 148.400 ;
        RECT 458.000 147.200 458.800 147.600 ;
        RECT 454.000 142.200 454.800 146.200 ;
        RECT 455.600 145.600 456.400 146.400 ;
        RECT 457.400 146.200 461.000 146.600 ;
        RECT 462.000 146.200 462.600 147.600 ;
        RECT 465.200 146.200 466.000 149.700 ;
        RECT 466.800 149.600 467.600 149.700 ;
        RECT 470.600 149.600 475.600 150.200 ;
        RECT 478.000 150.300 478.800 150.400 ;
        RECT 479.600 150.300 480.200 151.600 ;
        RECT 486.000 151.200 486.800 159.800 ;
        RECT 489.200 151.200 490.000 159.800 ;
        RECT 492.400 151.200 493.200 159.800 ;
        RECT 495.600 151.200 496.400 159.800 ;
        RECT 498.800 151.200 499.600 159.800 ;
        RECT 502.000 151.600 502.800 153.200 ;
        RECT 482.600 150.600 486.800 151.200 ;
        RECT 482.600 150.400 483.400 150.600 ;
        RECT 478.000 149.700 480.300 150.300 ;
        RECT 484.200 149.800 485.000 150.000 ;
        RECT 478.000 149.600 478.800 149.700 ;
        RECT 470.600 149.400 471.400 149.600 ;
        RECT 473.200 149.400 474.000 149.600 ;
        RECT 472.200 148.400 473.000 148.600 ;
        RECT 479.600 148.400 480.200 149.700 ;
        RECT 481.200 149.200 485.000 149.800 ;
        RECT 481.200 149.000 482.000 149.200 ;
        RECT 466.800 146.800 467.600 148.400 ;
        RECT 469.200 147.800 480.200 148.400 ;
        RECT 469.200 147.600 470.800 147.800 ;
        RECT 457.200 146.000 461.200 146.200 ;
        RECT 455.400 144.800 456.200 145.600 ;
        RECT 457.200 142.200 458.000 146.000 ;
        RECT 460.400 142.200 461.200 146.000 ;
        RECT 462.000 142.200 462.800 146.200 ;
        RECT 464.200 145.600 466.000 146.200 ;
        RECT 464.200 142.200 465.000 145.600 ;
        RECT 468.400 142.200 469.200 147.000 ;
        RECT 473.400 145.600 474.000 147.800 ;
        RECT 479.000 147.600 479.800 147.800 ;
        RECT 486.000 147.200 486.800 150.600 ;
        RECT 483.000 146.600 486.800 147.200 ;
        RECT 487.600 150.400 490.000 151.200 ;
        RECT 491.000 150.400 493.200 151.200 ;
        RECT 494.200 150.400 496.400 151.200 ;
        RECT 497.800 150.400 499.600 151.200 ;
        RECT 487.600 147.600 488.400 150.400 ;
        RECT 491.000 149.000 491.800 150.400 ;
        RECT 494.200 149.000 495.000 150.400 ;
        RECT 497.800 149.000 498.600 150.400 ;
        RECT 489.200 148.200 491.800 149.000 ;
        RECT 492.600 148.200 495.000 149.000 ;
        RECT 496.000 148.200 498.600 149.000 ;
        RECT 491.000 147.600 491.800 148.200 ;
        RECT 494.200 147.600 495.000 148.200 ;
        RECT 497.800 147.600 498.600 148.200 ;
        RECT 503.600 150.300 504.400 159.800 ;
        RECT 506.800 159.200 510.800 159.800 ;
        RECT 506.800 151.800 507.600 159.200 ;
        RECT 508.400 151.800 509.200 158.600 ;
        RECT 510.000 152.400 510.800 159.200 ;
        RECT 513.200 152.400 514.000 159.800 ;
        RECT 510.000 151.800 514.000 152.400 ;
        RECT 517.400 152.400 518.200 159.800 ;
        RECT 518.800 153.600 519.600 154.400 ;
        RECT 519.000 152.400 519.600 153.600 ;
        RECT 517.400 151.800 518.400 152.400 ;
        RECT 519.000 152.300 520.400 152.400 ;
        RECT 521.200 152.300 522.000 152.400 ;
        RECT 519.000 151.800 522.000 152.300 ;
        RECT 508.600 151.200 509.200 151.800 ;
        RECT 506.800 150.300 507.600 151.200 ;
        RECT 508.600 150.600 510.600 151.200 ;
        RECT 503.600 149.700 507.600 150.300 ;
        RECT 487.600 146.800 490.000 147.600 ;
        RECT 491.000 146.800 493.200 147.600 ;
        RECT 494.200 146.800 496.400 147.600 ;
        RECT 497.800 146.800 499.600 147.600 ;
        RECT 483.000 146.400 483.800 146.600 ;
        RECT 471.600 144.200 472.400 145.000 ;
        RECT 473.200 144.800 474.000 145.600 ;
        RECT 475.000 145.400 475.800 145.600 ;
        RECT 475.000 144.800 477.800 145.400 ;
        RECT 477.200 144.200 477.800 144.800 ;
        RECT 481.200 144.200 482.000 145.000 ;
        RECT 471.600 143.600 473.600 144.200 ;
        RECT 472.800 142.200 473.600 143.600 ;
        RECT 477.200 142.200 478.000 144.200 ;
        RECT 481.200 143.600 482.600 144.200 ;
        RECT 481.400 142.200 482.600 143.600 ;
        RECT 486.000 142.200 486.800 146.600 ;
        RECT 489.200 142.200 490.000 146.800 ;
        RECT 492.400 142.200 493.200 146.800 ;
        RECT 495.600 142.200 496.400 146.800 ;
        RECT 498.800 142.200 499.600 146.800 ;
        RECT 503.600 146.200 504.400 149.700 ;
        RECT 506.800 149.600 507.600 149.700 ;
        RECT 510.000 150.400 510.600 150.600 ;
        RECT 512.400 150.400 513.200 150.800 ;
        RECT 510.000 149.600 510.800 150.400 ;
        RECT 512.400 149.800 514.000 150.400 ;
        RECT 513.200 149.600 514.000 149.800 ;
        RECT 508.600 148.800 509.400 149.600 ;
        RECT 508.600 148.400 509.200 148.800 ;
        RECT 505.200 146.800 506.000 148.400 ;
        RECT 508.400 147.600 509.200 148.400 ;
        RECT 510.000 146.200 510.600 149.600 ;
        RECT 511.600 147.600 512.400 149.200 ;
        RECT 516.400 148.800 517.200 150.400 ;
        RECT 517.800 148.400 518.400 151.800 ;
        RECT 519.600 151.700 522.000 151.800 ;
        RECT 519.600 151.600 520.400 151.700 ;
        RECT 521.200 151.600 522.000 151.700 ;
        RECT 514.800 148.200 515.600 148.400 ;
        RECT 517.800 148.300 520.400 148.400 ;
        RECT 521.200 148.300 522.000 148.400 ;
        RECT 514.800 147.600 516.400 148.200 ;
        RECT 517.800 147.700 522.000 148.300 ;
        RECT 517.800 147.600 520.400 147.700 ;
        RECT 515.600 147.200 516.400 147.600 ;
        RECT 515.000 146.200 518.600 146.600 ;
        RECT 519.600 146.200 520.200 147.600 ;
        RECT 521.200 146.800 522.000 147.700 ;
        RECT 522.800 146.200 523.600 159.800 ;
        RECT 524.400 151.600 525.200 153.200 ;
        RECT 528.600 152.400 529.400 159.800 ;
        RECT 530.000 153.600 530.800 154.400 ;
        RECT 530.200 152.400 530.800 153.600 ;
        RECT 535.000 152.600 535.800 159.800 ;
        RECT 537.200 155.800 538.000 159.800 ;
        RECT 528.600 151.800 529.600 152.400 ;
        RECT 530.200 151.800 531.600 152.400 ;
        RECT 534.000 151.800 535.800 152.600 ;
        RECT 537.400 155.600 538.000 155.800 ;
        RECT 540.400 155.800 541.200 159.800 ;
        RECT 540.400 155.600 541.000 155.800 ;
        RECT 537.400 155.000 541.000 155.600 ;
        RECT 537.400 152.400 538.000 155.000 ;
        RECT 538.800 152.800 539.600 154.400 ;
        RECT 529.000 150.400 529.600 151.800 ;
        RECT 530.800 151.600 531.600 151.800 ;
        RECT 534.200 150.400 534.800 151.800 ;
        RECT 537.200 151.600 538.000 152.400 ;
        RECT 527.600 148.800 528.400 150.400 ;
        RECT 529.000 149.600 530.000 150.400 ;
        RECT 534.000 149.600 534.800 150.400 ;
        RECT 535.600 149.600 536.400 151.200 ;
        RECT 529.000 148.400 529.600 149.600 ;
        RECT 534.200 148.400 534.800 149.600 ;
        RECT 526.000 148.200 526.800 148.400 ;
        RECT 526.000 147.600 527.600 148.200 ;
        RECT 529.000 147.600 531.600 148.400 ;
        RECT 534.000 147.600 534.800 148.400 ;
        RECT 537.400 148.400 538.000 151.600 ;
        RECT 542.000 150.800 542.800 152.400 ;
        RECT 539.600 149.600 541.200 150.400 ;
        RECT 537.400 148.300 539.000 148.400 ;
        RECT 540.400 148.300 541.200 148.400 ;
        RECT 537.400 147.800 541.200 148.300 ;
        RECT 526.800 147.200 527.600 147.600 ;
        RECT 526.200 146.200 529.800 146.600 ;
        RECT 530.800 146.200 531.400 147.600 ;
        RECT 502.600 145.600 504.400 146.200 ;
        RECT 502.600 142.200 503.400 145.600 ;
        RECT 509.400 142.200 511.000 146.200 ;
        RECT 514.800 146.000 518.800 146.200 ;
        RECT 514.800 142.200 515.600 146.000 ;
        RECT 518.000 142.200 518.800 146.000 ;
        RECT 519.600 142.200 520.400 146.200 ;
        RECT 522.800 145.600 524.600 146.200 ;
        RECT 523.800 144.400 524.600 145.600 ;
        RECT 526.000 146.000 530.000 146.200 ;
        RECT 523.800 143.600 525.200 144.400 ;
        RECT 523.800 142.200 524.600 143.600 ;
        RECT 526.000 142.200 526.800 146.000 ;
        RECT 529.200 142.200 530.000 146.000 ;
        RECT 530.800 142.200 531.600 146.200 ;
        RECT 532.400 144.800 533.200 146.400 ;
        RECT 534.200 144.200 534.800 147.600 ;
        RECT 534.000 142.200 534.800 144.200 ;
        RECT 538.400 147.700 541.200 147.800 ;
        RECT 538.400 142.200 539.200 147.700 ;
        RECT 540.400 147.600 541.200 147.700 ;
        RECT 543.600 146.800 544.400 148.400 ;
        RECT 545.200 146.200 546.000 159.800 ;
        RECT 549.000 158.400 549.800 159.800 ;
        RECT 548.400 157.600 549.800 158.400 ;
        RECT 546.800 151.600 547.600 153.200 ;
        RECT 549.000 152.600 549.800 157.600 ;
        RECT 549.000 151.800 550.800 152.600 ;
        RECT 553.200 152.400 554.000 159.800 ;
        RECT 557.600 158.400 559.200 159.800 ;
        RECT 557.600 157.600 560.400 158.400 ;
        RECT 554.600 152.400 555.400 152.600 ;
        RECT 553.200 151.800 555.400 152.400 ;
        RECT 557.600 152.400 559.200 157.600 ;
        RECT 561.200 152.400 562.000 152.600 ;
        RECT 562.800 152.400 563.600 159.800 ;
        RECT 557.600 151.800 559.600 152.400 ;
        RECT 561.200 151.800 563.600 152.400 ;
        RECT 548.400 149.600 549.200 151.200 ;
        RECT 550.000 148.400 550.600 151.800 ;
        RECT 554.800 151.200 555.400 151.800 ;
        RECT 554.800 150.600 558.200 151.200 ;
        RECT 557.400 150.400 558.200 150.600 ;
        RECT 559.000 150.400 559.600 151.800 ;
        RECT 564.400 151.400 565.200 159.800 ;
        RECT 568.800 156.400 569.600 159.800 ;
        RECT 567.600 155.800 569.600 156.400 ;
        RECT 573.200 155.800 574.000 159.800 ;
        RECT 577.400 155.800 578.600 159.800 ;
        RECT 567.600 155.000 568.400 155.800 ;
        RECT 573.200 155.200 573.800 155.800 ;
        RECT 571.000 154.600 574.600 155.200 ;
        RECT 577.200 155.000 578.000 155.800 ;
        RECT 571.000 154.400 571.800 154.600 ;
        RECT 573.800 154.400 574.600 154.600 ;
        RECT 567.600 153.000 568.400 153.200 ;
        RECT 572.200 153.000 573.000 153.200 ;
        RECT 567.600 152.400 573.000 153.000 ;
        RECT 573.600 153.000 575.800 153.600 ;
        RECT 573.600 151.800 574.200 153.000 ;
        RECT 575.000 152.800 575.800 153.000 ;
        RECT 577.400 153.200 578.800 154.000 ;
        RECT 577.400 152.200 578.000 153.200 ;
        RECT 569.400 151.400 574.200 151.800 ;
        RECT 564.400 151.200 574.200 151.400 ;
        RECT 575.600 151.600 578.000 152.200 ;
        RECT 564.400 151.000 570.200 151.200 ;
        RECT 564.400 150.800 570.000 151.000 ;
        RECT 555.200 149.800 556.000 150.000 ;
        RECT 559.000 149.800 560.400 150.400 ;
        RECT 570.800 150.200 571.600 150.400 ;
        RECT 555.200 149.200 557.800 149.800 ;
        RECT 557.200 148.600 557.800 149.200 ;
        RECT 558.600 149.600 560.400 149.800 ;
        RECT 566.600 149.600 571.600 150.200 ;
        RECT 558.600 149.200 559.600 149.600 ;
        RECT 566.600 149.400 567.400 149.600 ;
        RECT 550.000 147.600 550.800 148.400 ;
        RECT 551.600 148.300 552.400 148.400 ;
        RECT 553.200 148.300 554.800 148.400 ;
        RECT 551.600 148.200 554.800 148.300 ;
        RECT 551.600 147.700 556.600 148.200 ;
        RECT 557.200 147.800 558.000 148.600 ;
        RECT 551.600 147.600 552.400 147.700 ;
        RECT 553.200 147.600 556.600 147.700 ;
        RECT 545.200 145.600 547.000 146.200 ;
        RECT 546.200 144.400 547.000 145.600 ;
        RECT 545.200 143.600 547.000 144.400 ;
        RECT 546.200 142.200 547.000 143.600 ;
        RECT 550.000 144.200 550.600 147.600 ;
        RECT 556.000 147.200 556.600 147.600 ;
        RECT 554.600 146.800 555.400 147.000 ;
        RECT 551.600 144.800 552.400 146.400 ;
        RECT 553.200 146.200 555.400 146.800 ;
        RECT 556.000 146.600 558.000 147.200 ;
        RECT 556.400 146.400 558.000 146.600 ;
        RECT 550.000 142.200 550.800 144.200 ;
        RECT 553.200 142.200 554.000 146.200 ;
        RECT 558.600 145.800 559.200 149.200 ;
        RECT 568.200 148.400 569.000 148.600 ;
        RECT 575.600 148.400 576.200 151.600 ;
        RECT 582.000 151.200 582.800 159.800 ;
        RECT 578.600 150.600 582.800 151.200 ;
        RECT 578.600 150.400 579.400 150.600 ;
        RECT 580.200 149.800 581.000 150.000 ;
        RECT 577.200 149.200 581.000 149.800 ;
        RECT 577.200 149.000 578.000 149.200 ;
        RECT 560.000 147.600 560.800 148.400 ;
        RECT 562.000 147.600 563.600 148.400 ;
        RECT 565.200 147.800 576.200 148.400 ;
        RECT 565.200 147.600 566.800 147.800 ;
        RECT 569.200 147.600 570.000 147.800 ;
        RECT 575.000 147.600 575.800 147.800 ;
        RECT 560.000 147.200 560.600 147.600 ;
        RECT 559.800 146.400 560.600 147.200 ;
        RECT 561.200 146.800 562.000 147.000 ;
        RECT 561.200 146.200 563.600 146.800 ;
        RECT 557.600 142.200 559.200 145.800 ;
        RECT 562.800 142.200 563.600 146.200 ;
        RECT 564.400 142.200 565.200 147.000 ;
        RECT 569.400 145.600 570.000 147.600 ;
        RECT 582.000 147.200 582.800 150.600 ;
        RECT 579.000 146.600 582.800 147.200 ;
        RECT 579.000 146.400 579.800 146.600 ;
        RECT 567.600 144.200 568.400 145.000 ;
        RECT 569.200 144.800 570.000 145.600 ;
        RECT 571.000 145.400 571.800 145.600 ;
        RECT 571.000 144.800 573.800 145.400 ;
        RECT 573.200 144.200 573.800 144.800 ;
        RECT 577.200 144.200 578.000 145.000 ;
        RECT 582.000 144.300 582.800 146.600 ;
        RECT 583.600 144.300 584.400 144.400 ;
        RECT 567.600 143.600 569.600 144.200 ;
        RECT 568.800 142.200 569.600 143.600 ;
        RECT 573.200 142.200 574.000 144.200 ;
        RECT 577.200 143.600 578.600 144.200 ;
        RECT 577.400 142.200 578.600 143.600 ;
        RECT 582.000 143.700 584.400 144.300 ;
        RECT 582.000 142.200 582.800 143.700 ;
        RECT 583.600 143.600 584.400 143.700 ;
        RECT 1.200 135.600 2.000 137.200 ;
        RECT 1.200 128.300 2.000 128.400 ;
        RECT 2.800 128.300 3.600 139.800 ;
        RECT 6.000 137.800 6.800 139.800 ;
        RECT 6.000 134.400 6.600 137.800 ;
        RECT 7.600 135.600 8.400 137.200 ;
        RECT 9.200 136.000 10.000 139.800 ;
        RECT 12.400 136.000 13.200 139.800 ;
        RECT 9.200 135.800 13.200 136.000 ;
        RECT 14.000 135.800 14.800 139.800 ;
        RECT 17.200 137.800 18.000 139.800 ;
        RECT 22.000 137.800 22.800 139.800 ;
        RECT 9.400 135.400 13.000 135.800 ;
        RECT 10.000 134.400 10.800 134.800 ;
        RECT 14.000 134.400 14.600 135.800 ;
        RECT 15.600 135.600 16.400 137.200 ;
        RECT 17.400 136.300 18.000 137.800 ;
        RECT 20.400 136.300 21.200 137.200 ;
        RECT 17.300 135.700 21.200 136.300 ;
        RECT 17.400 134.400 18.000 135.700 ;
        RECT 20.400 135.600 21.200 135.700 ;
        RECT 22.200 134.400 22.800 137.800 ;
        RECT 6.000 134.300 6.800 134.400 ;
        RECT 9.200 134.300 10.800 134.400 ;
        RECT 6.000 133.800 10.800 134.300 ;
        RECT 6.000 133.700 10.000 133.800 ;
        RECT 6.000 133.600 6.800 133.700 ;
        RECT 9.200 133.600 10.000 133.700 ;
        RECT 12.200 133.600 14.800 134.400 ;
        RECT 17.200 133.600 18.000 134.400 ;
        RECT 22.000 133.600 22.800 134.400 ;
        RECT 4.400 130.800 5.200 132.400 ;
        RECT 6.000 130.200 6.600 133.600 ;
        RECT 10.800 131.600 11.600 133.200 ;
        RECT 12.200 130.200 12.800 133.600 ;
        RECT 14.000 130.200 14.800 130.400 ;
        RECT 17.400 130.200 18.000 133.600 ;
        RECT 18.800 132.300 19.600 132.400 ;
        RECT 20.400 132.300 21.200 132.400 ;
        RECT 18.800 131.700 21.200 132.300 ;
        RECT 18.800 130.800 19.600 131.700 ;
        RECT 20.400 131.600 21.200 131.700 ;
        RECT 22.200 130.200 22.800 133.600 ;
        RECT 26.800 137.600 27.600 139.800 ;
        RECT 31.600 137.800 32.400 139.800 ;
        RECT 26.800 134.400 27.400 137.600 ;
        RECT 28.400 135.600 29.200 137.200 ;
        RECT 30.000 136.300 30.800 136.400 ;
        RECT 31.600 136.300 32.200 137.800 ;
        RECT 30.000 135.700 32.300 136.300 ;
        RECT 30.000 135.600 30.800 135.700 ;
        RECT 31.600 134.400 32.200 135.700 ;
        RECT 33.200 135.600 34.000 137.200 ;
        RECT 34.800 135.600 35.600 137.200 ;
        RECT 26.800 133.600 27.600 134.400 ;
        RECT 31.600 133.600 32.400 134.400 ;
        RECT 23.600 130.800 24.400 132.400 ;
        RECT 25.200 130.800 26.000 132.400 ;
        RECT 26.800 130.200 27.400 133.600 ;
        RECT 30.000 130.800 30.800 132.400 ;
        RECT 31.600 130.200 32.200 133.600 ;
        RECT 36.400 130.300 37.200 139.800 ;
        RECT 40.600 136.400 41.400 139.800 ;
        RECT 39.600 135.800 41.400 136.400 ;
        RECT 43.400 138.400 44.200 139.800 ;
        RECT 50.200 138.400 51.000 139.800 ;
        RECT 43.400 137.600 45.200 138.400 ;
        RECT 49.200 137.600 51.000 138.400 ;
        RECT 43.400 136.400 44.200 137.600 ;
        RECT 50.200 136.400 51.000 137.600 ;
        RECT 43.400 135.800 45.200 136.400 ;
        RECT 38.000 133.600 38.800 135.200 ;
        RECT 39.600 132.300 40.400 135.800 ;
        RECT 39.600 131.700 43.500 132.300 ;
        RECT 38.000 130.300 38.800 130.400 ;
        RECT 1.200 127.700 3.600 128.300 ;
        RECT 1.200 127.600 2.000 127.700 ;
        RECT 2.800 122.200 3.600 127.700 ;
        RECT 5.000 129.400 6.800 130.200 ;
        RECT 11.800 129.600 12.800 130.200 ;
        RECT 13.400 129.600 14.800 130.200 ;
        RECT 5.000 124.400 5.800 129.400 ;
        RECT 11.800 124.400 12.600 129.600 ;
        RECT 13.400 128.400 14.000 129.600 ;
        RECT 17.200 129.400 19.000 130.200 ;
        RECT 22.000 129.400 23.800 130.200 ;
        RECT 13.200 127.600 14.000 128.400 ;
        RECT 4.400 123.600 5.800 124.400 ;
        RECT 10.800 123.600 12.600 124.400 ;
        RECT 5.000 122.200 5.800 123.600 ;
        RECT 11.800 122.200 12.600 123.600 ;
        RECT 18.200 122.200 19.000 129.400 ;
        RECT 23.000 124.400 23.800 129.400 ;
        RECT 22.000 123.600 23.800 124.400 ;
        RECT 23.000 122.200 23.800 123.600 ;
        RECT 25.800 129.400 27.600 130.200 ;
        RECT 30.600 129.400 32.400 130.200 ;
        RECT 36.400 129.700 38.800 130.300 ;
        RECT 25.800 122.200 26.600 129.400 ;
        RECT 30.600 122.200 31.400 129.400 ;
        RECT 36.400 122.200 37.200 129.700 ;
        RECT 38.000 129.600 38.800 129.700 ;
        RECT 39.600 122.200 40.400 131.700 ;
        RECT 42.900 130.400 43.500 131.700 ;
        RECT 41.200 128.800 42.000 130.400 ;
        RECT 42.800 128.800 43.600 130.400 ;
        RECT 44.400 122.200 45.200 135.800 ;
        RECT 49.200 135.800 51.000 136.400 ;
        RECT 52.400 136.000 53.200 139.800 ;
        RECT 55.600 136.000 56.400 139.800 ;
        RECT 52.400 135.800 56.400 136.000 ;
        RECT 57.200 135.800 58.000 139.800 ;
        RECT 61.400 138.400 62.200 139.800 ;
        RECT 60.400 137.600 62.200 138.400 ;
        RECT 61.400 136.400 62.200 137.600 ;
        RECT 60.400 135.800 62.200 136.400 ;
        RECT 46.000 133.600 46.800 135.200 ;
        RECT 47.600 133.600 48.400 135.200 ;
        RECT 46.100 132.300 46.700 133.600 ;
        RECT 49.200 132.300 50.000 135.800 ;
        RECT 52.600 135.400 56.200 135.800 ;
        RECT 53.200 134.400 54.000 134.800 ;
        RECT 57.200 134.400 57.800 135.800 ;
        RECT 52.400 133.800 54.000 134.400 ;
        RECT 52.400 133.600 53.200 133.800 ;
        RECT 55.400 133.600 58.000 134.400 ;
        RECT 58.800 133.600 59.600 135.200 ;
        RECT 54.000 132.300 54.800 133.200 ;
        RECT 46.100 131.700 50.000 132.300 ;
        RECT 49.200 122.200 50.000 131.700 ;
        RECT 50.900 131.700 54.800 132.300 ;
        RECT 50.900 130.400 51.500 131.700 ;
        RECT 54.000 131.600 54.800 131.700 ;
        RECT 50.800 128.800 51.600 130.400 ;
        RECT 55.400 130.200 56.000 133.600 ;
        RECT 57.200 130.200 58.000 130.400 ;
        RECT 55.000 129.600 56.000 130.200 ;
        RECT 56.600 129.600 58.000 130.200 ;
        RECT 55.000 122.200 55.800 129.600 ;
        RECT 56.600 128.400 57.200 129.600 ;
        RECT 56.400 127.600 57.200 128.400 ;
        RECT 60.400 122.200 61.200 135.800 ;
        RECT 62.000 128.800 62.800 130.400 ;
        RECT 63.600 122.200 64.400 139.800 ;
        RECT 70.600 136.000 71.400 139.000 ;
        RECT 74.800 137.000 75.600 139.000 ;
        RECT 69.800 135.400 71.400 136.000 ;
        RECT 65.200 133.600 66.000 135.200 ;
        RECT 69.800 135.000 70.600 135.400 ;
        RECT 69.800 134.400 70.400 135.000 ;
        RECT 75.000 134.800 75.600 137.000 ;
        RECT 76.400 136.000 77.200 139.800 ;
        RECT 79.600 136.000 80.400 139.800 ;
        RECT 76.400 135.800 80.400 136.000 ;
        RECT 81.200 135.800 82.000 139.800 ;
        RECT 82.800 135.800 83.600 139.800 ;
        RECT 84.400 136.000 85.200 139.800 ;
        RECT 87.600 136.000 88.400 139.800 ;
        RECT 84.400 135.800 88.400 136.000 ;
        RECT 76.600 135.400 80.200 135.800 ;
        RECT 68.400 133.600 70.400 134.400 ;
        RECT 71.400 134.200 75.600 134.800 ;
        RECT 77.200 134.400 78.000 134.800 ;
        RECT 81.200 134.400 81.800 135.800 ;
        RECT 83.000 134.400 83.600 135.800 ;
        RECT 84.600 135.400 88.200 135.800 ;
        RECT 86.800 134.400 87.600 134.800 ;
        RECT 71.400 133.800 72.400 134.200 ;
        RECT 68.400 130.800 69.200 132.400 ;
        RECT 69.800 129.800 70.400 133.600 ;
        RECT 71.000 133.000 72.400 133.800 ;
        RECT 76.400 133.800 78.000 134.400 ;
        RECT 76.400 133.600 77.200 133.800 ;
        RECT 79.400 133.600 82.000 134.400 ;
        RECT 82.800 133.600 85.400 134.400 ;
        RECT 86.800 133.800 88.400 134.400 ;
        RECT 87.600 133.600 88.400 133.800 ;
        RECT 71.800 131.000 72.400 133.000 ;
        RECT 73.200 131.600 74.000 133.200 ;
        RECT 74.800 131.600 75.600 133.200 ;
        RECT 78.000 131.600 78.800 133.200 ;
        RECT 79.400 132.300 80.000 133.600 ;
        RECT 79.400 131.700 83.500 132.300 ;
        RECT 71.800 130.400 75.600 131.000 ;
        RECT 69.800 129.200 71.400 129.800 ;
        RECT 70.600 124.400 71.400 129.200 ;
        RECT 75.000 127.000 75.600 130.400 ;
        RECT 79.400 130.200 80.000 131.700 ;
        RECT 82.900 130.400 83.500 131.700 ;
        RECT 81.200 130.200 82.000 130.400 ;
        RECT 70.600 123.600 72.400 124.400 ;
        RECT 70.600 122.200 71.400 123.600 ;
        RECT 74.800 123.000 75.600 127.000 ;
        RECT 79.000 129.600 80.000 130.200 ;
        RECT 80.600 129.600 82.000 130.200 ;
        RECT 82.800 130.200 83.600 130.400 ;
        RECT 84.800 130.200 85.400 133.600 ;
        RECT 86.000 132.300 86.800 133.200 ;
        RECT 89.200 132.300 90.000 139.800 ;
        RECT 90.800 135.600 91.600 137.200 ;
        RECT 92.400 136.000 93.200 139.800 ;
        RECT 95.600 136.000 96.400 139.800 ;
        RECT 92.400 135.800 96.400 136.000 ;
        RECT 97.200 135.800 98.000 139.800 ;
        RECT 98.800 135.800 99.600 139.800 ;
        RECT 100.400 136.000 101.200 139.800 ;
        RECT 103.600 136.000 104.400 139.800 ;
        RECT 100.400 135.800 104.400 136.000 ;
        RECT 105.800 136.400 106.600 139.800 ;
        RECT 105.800 135.800 107.600 136.400 ;
        RECT 92.600 135.400 96.200 135.800 ;
        RECT 93.200 134.400 94.000 134.800 ;
        RECT 97.200 134.400 97.800 135.800 ;
        RECT 99.000 134.400 99.600 135.800 ;
        RECT 100.600 135.400 104.200 135.800 ;
        RECT 102.800 134.400 103.600 134.800 ;
        RECT 92.400 133.800 94.000 134.400 ;
        RECT 92.400 133.600 93.200 133.800 ;
        RECT 95.400 133.600 98.000 134.400 ;
        RECT 98.800 133.600 101.400 134.400 ;
        RECT 102.800 133.800 104.400 134.400 ;
        RECT 103.600 133.600 104.400 133.800 ;
        RECT 86.000 131.700 90.000 132.300 ;
        RECT 86.000 131.600 86.800 131.700 ;
        RECT 82.800 129.600 84.200 130.200 ;
        RECT 84.800 129.600 85.800 130.200 ;
        RECT 79.000 122.200 79.800 129.600 ;
        RECT 80.600 128.400 81.200 129.600 ;
        RECT 80.400 127.600 81.200 128.400 ;
        RECT 83.600 128.400 84.200 129.600 ;
        RECT 83.600 127.600 84.400 128.400 ;
        RECT 85.000 122.200 85.800 129.600 ;
        RECT 89.200 122.200 90.000 131.700 ;
        RECT 94.000 131.600 94.800 133.200 ;
        RECT 95.400 132.300 96.000 133.600 ;
        RECT 95.400 131.700 99.500 132.300 ;
        RECT 95.400 130.200 96.000 131.700 ;
        RECT 98.900 130.400 99.500 131.700 ;
        RECT 97.200 130.200 98.000 130.400 ;
        RECT 95.000 129.600 96.000 130.200 ;
        RECT 96.600 129.600 98.000 130.200 ;
        RECT 98.800 130.200 99.600 130.400 ;
        RECT 100.800 130.200 101.400 133.600 ;
        RECT 102.000 132.300 102.800 133.200 ;
        RECT 102.000 131.700 105.900 132.300 ;
        RECT 102.000 131.600 102.800 131.700 ;
        RECT 105.300 130.400 105.900 131.700 ;
        RECT 98.800 129.600 100.200 130.200 ;
        RECT 100.800 129.600 101.800 130.200 ;
        RECT 95.000 122.200 95.800 129.600 ;
        RECT 96.600 128.400 97.200 129.600 ;
        RECT 96.400 127.600 97.200 128.400 ;
        RECT 99.600 128.400 100.200 129.600 ;
        RECT 99.600 127.600 100.400 128.400 ;
        RECT 101.000 124.400 101.800 129.600 ;
        RECT 105.200 128.800 106.000 130.400 ;
        RECT 106.800 130.300 107.600 135.800 ;
        RECT 110.000 135.600 110.800 139.800 ;
        RECT 111.600 136.000 112.400 139.800 ;
        RECT 114.800 136.000 115.600 139.800 ;
        RECT 119.000 136.400 119.800 139.800 ;
        RECT 111.600 135.800 115.600 136.000 ;
        RECT 118.000 135.800 119.800 136.400 ;
        RECT 121.200 135.800 122.000 139.800 ;
        RECT 122.800 136.000 123.600 139.800 ;
        RECT 126.000 136.000 126.800 139.800 ;
        RECT 122.800 135.800 126.800 136.000 ;
        RECT 128.200 138.400 129.000 139.800 ;
        RECT 128.200 137.600 130.000 138.400 ;
        RECT 128.200 136.400 129.000 137.600 ;
        RECT 128.200 135.800 130.000 136.400 ;
        RECT 108.400 133.600 109.200 135.200 ;
        RECT 110.200 134.400 110.800 135.600 ;
        RECT 111.800 135.400 115.400 135.800 ;
        RECT 114.000 134.400 114.800 134.800 ;
        RECT 110.000 133.600 112.600 134.400 ;
        RECT 114.000 133.800 115.600 134.400 ;
        RECT 114.800 133.600 115.600 133.800 ;
        RECT 116.400 133.600 117.200 135.200 ;
        RECT 110.000 130.300 110.800 130.400 ;
        RECT 106.800 130.200 110.800 130.300 ;
        RECT 112.000 130.200 112.600 133.600 ;
        RECT 113.200 132.300 114.000 133.200 ;
        RECT 114.800 132.300 115.600 132.400 ;
        RECT 113.200 131.700 115.600 132.300 ;
        RECT 113.200 131.600 114.000 131.700 ;
        RECT 114.800 131.600 115.600 131.700 ;
        RECT 118.000 132.300 118.800 135.800 ;
        RECT 121.400 134.400 122.000 135.800 ;
        RECT 123.000 135.400 126.600 135.800 ;
        RECT 125.200 134.400 126.000 134.800 ;
        RECT 121.200 133.600 123.800 134.400 ;
        RECT 125.200 133.800 126.800 134.400 ;
        RECT 126.000 133.600 126.800 133.800 ;
        RECT 118.000 131.700 121.900 132.300 ;
        RECT 106.800 129.700 111.400 130.200 ;
        RECT 101.000 123.600 102.800 124.400 ;
        RECT 101.000 122.200 101.800 123.600 ;
        RECT 106.800 122.200 107.600 129.700 ;
        RECT 110.000 129.600 111.400 129.700 ;
        RECT 112.000 129.600 113.000 130.200 ;
        RECT 110.800 128.400 111.400 129.600 ;
        RECT 110.800 127.600 111.600 128.400 ;
        RECT 112.200 122.200 113.000 129.600 ;
        RECT 118.000 122.200 118.800 131.700 ;
        RECT 121.300 130.400 121.900 131.700 ;
        RECT 119.600 128.800 120.400 130.400 ;
        RECT 121.200 130.200 122.000 130.400 ;
        RECT 123.200 130.200 123.800 133.600 ;
        RECT 124.400 132.300 125.200 133.200 ;
        RECT 126.000 132.300 126.800 132.400 ;
        RECT 124.400 131.700 126.800 132.300 ;
        RECT 124.400 131.600 125.200 131.700 ;
        RECT 126.000 131.600 126.800 131.700 ;
        RECT 121.200 129.600 122.600 130.200 ;
        RECT 123.200 129.600 124.200 130.200 ;
        RECT 122.000 128.400 122.600 129.600 ;
        RECT 122.000 127.600 122.800 128.400 ;
        RECT 123.400 122.200 124.200 129.600 ;
        RECT 127.600 128.800 128.400 130.400 ;
        RECT 129.200 122.200 130.000 135.800 ;
        RECT 137.200 135.800 138.000 139.800 ;
        RECT 141.600 136.200 143.200 139.800 ;
        RECT 137.200 135.200 139.600 135.800 ;
        RECT 130.800 134.300 131.600 135.200 ;
        RECT 138.800 135.000 139.600 135.200 ;
        RECT 140.200 134.800 141.000 135.600 ;
        RECT 140.200 134.400 140.800 134.800 ;
        RECT 137.200 134.300 138.800 134.400 ;
        RECT 130.800 133.700 138.800 134.300 ;
        RECT 130.800 133.600 131.600 133.700 ;
        RECT 137.200 133.600 138.800 133.700 ;
        RECT 140.000 133.600 140.800 134.400 ;
        RECT 141.600 132.800 142.200 136.200 ;
        RECT 146.800 135.800 147.600 139.800 ;
        RECT 142.800 135.400 144.400 135.600 ;
        RECT 142.800 134.800 144.800 135.400 ;
        RECT 145.400 135.200 147.600 135.800 ;
        RECT 148.400 135.800 149.200 139.800 ;
        RECT 152.800 136.200 154.400 139.800 ;
        RECT 148.400 135.200 150.600 135.800 ;
        RECT 151.600 135.400 153.200 135.600 ;
        RECT 145.400 135.000 146.200 135.200 ;
        RECT 149.800 135.000 150.600 135.200 ;
        RECT 144.200 134.400 144.800 134.800 ;
        RECT 151.200 134.800 153.200 135.400 ;
        RECT 151.200 134.400 151.800 134.800 ;
        RECT 142.800 133.400 143.600 134.200 ;
        RECT 144.200 133.800 147.600 134.400 ;
        RECT 146.000 133.600 147.600 133.800 ;
        RECT 148.400 133.800 151.800 134.400 ;
        RECT 148.400 133.600 150.000 133.800 ;
        RECT 141.200 132.400 142.200 132.800 ;
        RECT 140.400 132.200 142.200 132.400 ;
        RECT 143.000 132.800 143.600 133.400 ;
        RECT 152.400 133.400 153.200 134.200 ;
        RECT 152.400 132.800 153.000 133.400 ;
        RECT 143.000 132.200 145.600 132.800 ;
        RECT 140.400 131.600 141.800 132.200 ;
        RECT 144.800 132.000 145.600 132.200 ;
        RECT 150.400 132.200 153.000 132.800 ;
        RECT 153.800 132.800 154.400 136.200 ;
        RECT 158.000 135.800 158.800 139.800 ;
        RECT 155.000 134.800 155.800 135.600 ;
        RECT 156.400 135.200 158.800 135.800 ;
        RECT 156.400 135.000 157.200 135.200 ;
        RECT 159.600 135.000 160.400 139.800 ;
        RECT 164.000 138.400 164.800 139.800 ;
        RECT 162.800 137.800 164.800 138.400 ;
        RECT 168.400 137.800 169.200 139.800 ;
        RECT 172.600 138.400 173.800 139.800 ;
        RECT 172.400 137.800 173.800 138.400 ;
        RECT 162.800 137.000 163.600 137.800 ;
        RECT 168.400 137.200 169.000 137.800 ;
        RECT 164.400 135.600 165.200 137.200 ;
        RECT 166.200 136.600 169.000 137.200 ;
        RECT 172.400 137.000 173.200 137.800 ;
        RECT 166.200 136.400 167.000 136.600 ;
        RECT 155.200 134.400 155.800 134.800 ;
        RECT 155.200 133.600 156.000 134.400 ;
        RECT 157.200 133.600 158.800 134.400 ;
        RECT 160.400 134.200 162.000 134.400 ;
        RECT 164.600 134.200 165.200 135.600 ;
        RECT 174.200 135.400 175.000 135.600 ;
        RECT 177.200 135.400 178.000 139.800 ;
        RECT 181.400 136.400 182.200 139.800 ;
        RECT 186.200 136.400 187.000 139.800 ;
        RECT 174.200 134.800 178.000 135.400 ;
        RECT 180.400 135.800 182.200 136.400 ;
        RECT 185.200 135.800 187.000 136.400 ;
        RECT 170.200 134.200 171.000 134.400 ;
        RECT 160.400 133.600 171.400 134.200 ;
        RECT 163.400 133.400 164.200 133.600 ;
        RECT 153.800 132.400 154.800 132.800 ;
        RECT 161.800 132.400 162.600 132.600 ;
        RECT 164.400 132.400 165.200 132.600 ;
        RECT 153.800 132.200 155.600 132.400 ;
        RECT 150.400 132.000 151.200 132.200 ;
        RECT 154.200 131.600 155.600 132.200 ;
        RECT 161.800 131.800 166.800 132.400 ;
        RECT 166.000 131.600 166.800 131.800 ;
        RECT 141.200 130.200 141.800 131.600 ;
        RECT 142.600 131.400 143.400 131.600 ;
        RECT 152.600 131.400 153.400 131.600 ;
        RECT 142.600 130.800 146.000 131.400 ;
        RECT 145.400 130.200 146.000 130.800 ;
        RECT 150.000 130.800 153.400 131.400 ;
        RECT 150.000 130.200 150.600 130.800 ;
        RECT 154.200 130.200 154.800 131.600 ;
        RECT 159.600 131.000 165.200 131.200 ;
        RECT 159.600 130.800 165.400 131.000 ;
        RECT 159.600 130.600 169.400 130.800 ;
        RECT 137.200 129.600 139.600 130.200 ;
        RECT 141.200 129.600 143.200 130.200 ;
        RECT 137.200 122.200 138.000 129.600 ;
        RECT 138.800 129.400 139.600 129.600 ;
        RECT 141.600 122.200 143.200 129.600 ;
        RECT 145.400 129.600 147.600 130.200 ;
        RECT 145.400 129.400 146.200 129.600 ;
        RECT 146.800 122.200 147.600 129.600 ;
        RECT 148.400 129.600 150.600 130.200 ;
        RECT 148.400 122.200 149.200 129.600 ;
        RECT 149.800 129.400 150.600 129.600 ;
        RECT 152.800 129.600 154.800 130.200 ;
        RECT 156.400 129.600 158.800 130.200 ;
        RECT 152.800 124.400 154.400 129.600 ;
        RECT 156.400 129.400 157.200 129.600 ;
        RECT 151.600 123.600 154.400 124.400 ;
        RECT 152.800 122.200 154.400 123.600 ;
        RECT 158.000 122.200 158.800 129.600 ;
        RECT 159.600 122.200 160.400 130.600 ;
        RECT 164.600 130.200 169.400 130.600 ;
        RECT 162.800 129.000 168.200 129.600 ;
        RECT 162.800 128.800 163.600 129.000 ;
        RECT 167.400 128.800 168.200 129.000 ;
        RECT 168.800 129.000 169.400 130.200 ;
        RECT 170.800 130.400 171.400 133.600 ;
        RECT 172.400 132.800 173.200 133.000 ;
        RECT 172.400 132.200 176.200 132.800 ;
        RECT 175.400 132.000 176.200 132.200 ;
        RECT 173.800 131.400 174.600 131.600 ;
        RECT 177.200 131.400 178.000 134.800 ;
        RECT 178.800 133.600 179.600 135.200 ;
        RECT 180.400 134.300 181.200 135.800 ;
        RECT 183.600 134.300 184.400 135.200 ;
        RECT 180.400 133.700 184.400 134.300 ;
        RECT 173.800 130.800 178.000 131.400 ;
        RECT 170.800 129.800 173.200 130.400 ;
        RECT 170.200 129.000 171.000 129.200 ;
        RECT 168.800 128.400 171.000 129.000 ;
        RECT 172.600 128.800 173.200 129.800 ;
        RECT 172.600 128.400 174.000 128.800 ;
        RECT 172.600 128.000 174.800 128.400 ;
        RECT 173.400 127.600 174.800 128.000 ;
        RECT 166.200 127.400 167.000 127.600 ;
        RECT 169.000 127.400 169.800 127.600 ;
        RECT 162.800 126.200 163.600 127.000 ;
        RECT 166.200 126.800 169.800 127.400 ;
        RECT 168.400 126.200 169.000 126.800 ;
        RECT 172.400 126.200 173.200 127.000 ;
        RECT 162.800 125.600 164.800 126.200 ;
        RECT 164.000 122.200 164.800 125.600 ;
        RECT 168.400 122.200 169.200 126.200 ;
        RECT 172.600 122.200 173.800 126.200 ;
        RECT 177.200 122.200 178.000 130.800 ;
        RECT 180.400 122.200 181.200 133.700 ;
        RECT 183.600 133.600 184.400 133.700 ;
        RECT 182.000 128.800 182.800 130.400 ;
        RECT 185.200 122.200 186.000 135.800 ;
        RECT 188.400 135.600 189.200 137.200 ;
        RECT 190.000 132.300 190.800 139.800 ;
        RECT 191.600 136.000 192.400 139.800 ;
        RECT 194.800 136.000 195.600 139.800 ;
        RECT 191.600 135.800 195.600 136.000 ;
        RECT 196.400 135.800 197.200 139.800 ;
        RECT 200.600 138.400 201.400 139.800 ;
        RECT 200.600 137.600 202.000 138.400 ;
        RECT 204.400 137.800 205.200 139.800 ;
        RECT 200.600 136.400 201.400 137.600 ;
        RECT 199.600 135.800 201.400 136.400 ;
        RECT 191.800 135.400 195.400 135.800 ;
        RECT 192.400 134.400 193.200 134.800 ;
        RECT 196.400 134.400 197.000 135.800 ;
        RECT 191.600 133.800 193.200 134.400 ;
        RECT 191.600 133.600 192.400 133.800 ;
        RECT 194.600 133.600 197.200 134.400 ;
        RECT 198.000 133.600 198.800 135.200 ;
        RECT 191.600 132.300 192.400 132.400 ;
        RECT 190.000 131.700 192.400 132.300 ;
        RECT 186.800 130.300 187.600 130.400 ;
        RECT 188.400 130.300 189.200 130.400 ;
        RECT 186.800 129.700 189.200 130.300 ;
        RECT 186.800 128.800 187.600 129.700 ;
        RECT 188.400 129.600 189.200 129.700 ;
        RECT 190.000 122.200 190.800 131.700 ;
        RECT 191.600 131.600 192.400 131.700 ;
        RECT 193.200 131.600 194.000 133.200 ;
        RECT 194.600 130.200 195.200 133.600 ;
        RECT 196.400 130.200 197.200 130.400 ;
        RECT 194.200 129.600 195.200 130.200 ;
        RECT 195.800 129.600 197.200 130.200 ;
        RECT 194.200 124.400 195.000 129.600 ;
        RECT 195.800 128.400 196.400 129.600 ;
        RECT 195.600 127.600 196.400 128.400 ;
        RECT 193.200 123.600 195.000 124.400 ;
        RECT 194.200 122.200 195.000 123.600 ;
        RECT 199.600 122.200 200.400 135.800 ;
        RECT 204.400 134.400 205.000 137.800 ;
        RECT 206.000 135.600 206.800 137.200 ;
        RECT 207.600 135.800 208.400 139.800 ;
        RECT 209.200 136.000 210.000 139.800 ;
        RECT 212.400 136.000 213.200 139.800 ;
        RECT 209.200 135.800 213.200 136.000 ;
        RECT 214.000 136.000 214.800 139.800 ;
        RECT 217.200 136.000 218.000 139.800 ;
        RECT 214.000 135.800 218.000 136.000 ;
        RECT 218.800 135.800 219.600 139.800 ;
        RECT 220.400 135.800 221.200 139.800 ;
        RECT 222.000 136.000 222.800 139.800 ;
        RECT 225.200 136.000 226.000 139.800 ;
        RECT 222.000 135.800 226.000 136.000 ;
        RECT 226.800 136.000 227.600 139.800 ;
        RECT 230.000 136.000 230.800 139.800 ;
        RECT 226.800 135.800 230.800 136.000 ;
        RECT 231.600 135.800 232.400 139.800 ;
        RECT 233.200 136.000 234.000 139.800 ;
        RECT 236.400 136.000 237.200 139.800 ;
        RECT 233.200 135.800 237.200 136.000 ;
        RECT 238.000 135.800 238.800 139.800 ;
        RECT 243.400 138.400 244.200 139.000 ;
        RECT 242.800 137.600 244.200 138.400 ;
        RECT 243.400 136.000 244.200 137.600 ;
        RECT 247.600 137.000 248.400 139.000 ;
        RECT 207.800 134.400 208.400 135.800 ;
        RECT 209.400 135.400 213.000 135.800 ;
        RECT 214.200 135.400 217.800 135.800 ;
        RECT 211.600 134.400 212.400 134.800 ;
        RECT 214.800 134.400 215.600 134.800 ;
        RECT 218.800 134.400 219.400 135.800 ;
        RECT 220.600 134.400 221.200 135.800 ;
        RECT 222.200 135.400 225.800 135.800 ;
        RECT 227.000 135.400 230.600 135.800 ;
        RECT 224.400 134.400 225.200 134.800 ;
        RECT 227.600 134.400 228.400 134.800 ;
        RECT 231.600 134.400 232.200 135.800 ;
        RECT 233.400 135.400 237.000 135.800 ;
        RECT 234.000 134.400 234.800 134.800 ;
        RECT 238.000 134.400 238.600 135.800 ;
        RECT 242.600 135.400 244.200 136.000 ;
        RECT 242.600 135.000 243.400 135.400 ;
        RECT 242.600 134.400 243.200 135.000 ;
        RECT 247.800 134.800 248.400 137.000 ;
        RECT 204.400 133.600 205.200 134.400 ;
        RECT 207.600 133.600 210.200 134.400 ;
        RECT 211.600 133.800 213.200 134.400 ;
        RECT 212.400 133.600 213.200 133.800 ;
        RECT 214.000 133.800 215.600 134.400 ;
        RECT 214.000 133.600 214.800 133.800 ;
        RECT 217.000 133.600 219.600 134.400 ;
        RECT 220.400 133.600 223.000 134.400 ;
        RECT 224.400 133.800 226.000 134.400 ;
        RECT 225.200 133.600 226.000 133.800 ;
        RECT 226.800 133.800 228.400 134.400 ;
        RECT 226.800 133.600 227.600 133.800 ;
        RECT 229.800 133.600 232.400 134.400 ;
        RECT 233.200 133.800 234.800 134.400 ;
        RECT 233.200 133.600 234.000 133.800 ;
        RECT 236.200 133.600 238.800 134.400 ;
        RECT 241.200 133.600 243.200 134.400 ;
        RECT 244.200 134.200 248.400 134.800 ;
        RECT 252.400 135.800 253.200 139.800 ;
        RECT 257.200 137.800 258.000 139.800 ;
        RECT 253.800 136.400 254.600 137.200 ;
        RECT 244.200 133.800 245.200 134.200 ;
        RECT 202.800 132.300 203.600 132.400 ;
        RECT 201.300 131.700 203.600 132.300 ;
        RECT 201.300 130.400 201.900 131.700 ;
        RECT 202.800 130.800 203.600 131.700 ;
        RECT 201.200 128.800 202.000 130.400 ;
        RECT 204.400 130.200 205.000 133.600 ;
        RECT 207.600 130.200 208.400 130.400 ;
        RECT 209.600 130.200 210.200 133.600 ;
        RECT 210.800 131.600 211.600 133.200 ;
        RECT 212.500 132.300 213.100 133.600 ;
        RECT 214.000 132.300 214.800 132.400 ;
        RECT 212.500 131.700 214.800 132.300 ;
        RECT 214.000 131.600 214.800 131.700 ;
        RECT 215.600 131.600 216.400 133.200 ;
        RECT 217.000 132.300 217.600 133.600 ;
        RECT 217.000 131.700 221.100 132.300 ;
        RECT 217.000 130.200 217.600 131.700 ;
        RECT 220.500 130.400 221.100 131.700 ;
        RECT 218.800 130.200 219.600 130.400 ;
        RECT 203.400 129.400 205.200 130.200 ;
        RECT 207.600 129.600 209.000 130.200 ;
        RECT 209.600 129.600 210.600 130.200 ;
        RECT 203.400 124.400 204.200 129.400 ;
        RECT 208.400 128.400 209.000 129.600 ;
        RECT 209.800 128.400 210.600 129.600 ;
        RECT 216.600 129.600 217.600 130.200 ;
        RECT 218.200 129.600 219.600 130.200 ;
        RECT 220.400 130.200 221.200 130.400 ;
        RECT 222.400 130.200 223.000 133.600 ;
        RECT 223.600 131.600 224.400 133.200 ;
        RECT 228.400 131.600 229.200 133.200 ;
        RECT 229.800 130.200 230.400 133.600 ;
        RECT 234.800 131.600 235.600 133.200 ;
        RECT 236.200 132.300 236.800 133.600 ;
        RECT 241.200 132.300 242.000 132.400 ;
        RECT 236.200 131.700 242.000 132.300 ;
        RECT 231.600 130.200 232.400 130.400 ;
        RECT 236.200 130.200 236.800 131.700 ;
        RECT 241.200 130.800 242.000 131.700 ;
        RECT 238.000 130.200 238.800 130.400 ;
        RECT 220.400 129.600 221.800 130.200 ;
        RECT 222.400 129.600 223.400 130.200 ;
        RECT 208.400 127.600 209.200 128.400 ;
        RECT 209.800 127.600 211.600 128.400 ;
        RECT 203.400 123.600 205.200 124.400 ;
        RECT 203.400 122.200 204.200 123.600 ;
        RECT 209.800 122.200 210.600 127.600 ;
        RECT 216.600 122.200 217.400 129.600 ;
        RECT 218.200 128.400 218.800 129.600 ;
        RECT 218.000 127.600 218.800 128.400 ;
        RECT 221.200 128.400 221.800 129.600 ;
        RECT 221.200 127.600 222.000 128.400 ;
        RECT 222.600 124.400 223.400 129.600 ;
        RECT 229.400 129.600 230.400 130.200 ;
        RECT 231.000 129.600 232.400 130.200 ;
        RECT 235.800 129.600 236.800 130.200 ;
        RECT 237.400 129.600 238.800 130.200 ;
        RECT 242.600 129.800 243.200 133.600 ;
        RECT 243.800 133.000 245.200 133.800 ;
        RECT 244.600 131.000 245.200 133.000 ;
        RECT 246.000 131.600 246.800 133.200 ;
        RECT 247.600 131.600 248.400 133.200 ;
        RECT 250.800 132.800 251.600 134.400 ;
        RECT 252.400 132.400 253.000 135.800 ;
        RECT 254.000 135.600 254.800 136.400 ;
        RECT 255.600 135.600 256.400 137.200 ;
        RECT 254.100 134.300 254.700 135.600 ;
        RECT 257.400 134.400 258.000 137.800 ;
        RECT 258.800 136.300 259.600 136.400 ;
        RECT 260.400 136.300 261.200 137.200 ;
        RECT 258.800 135.700 261.200 136.300 ;
        RECT 258.800 135.600 259.600 135.700 ;
        RECT 260.400 135.600 261.200 135.700 ;
        RECT 257.200 134.300 258.000 134.400 ;
        RECT 254.100 133.700 258.000 134.300 ;
        RECT 257.200 133.600 258.000 133.700 ;
        RECT 249.200 132.200 250.000 132.400 ;
        RECT 252.400 132.200 253.200 132.400 ;
        RECT 254.000 132.200 254.800 132.400 ;
        RECT 249.200 131.600 250.800 132.200 ;
        RECT 252.400 131.600 254.800 132.200 ;
        RECT 250.000 131.200 250.800 131.600 ;
        RECT 244.600 130.400 248.400 131.000 ;
        RECT 222.600 123.600 224.400 124.400 ;
        RECT 222.600 122.200 223.400 123.600 ;
        RECT 229.400 122.200 230.200 129.600 ;
        RECT 231.000 128.400 231.600 129.600 ;
        RECT 230.800 127.600 231.600 128.400 ;
        RECT 235.800 122.200 236.600 129.600 ;
        RECT 237.400 128.400 238.000 129.600 ;
        RECT 242.600 129.200 244.200 129.800 ;
        RECT 237.200 127.600 238.000 128.400 ;
        RECT 243.400 122.200 244.200 129.200 ;
        RECT 247.800 127.000 248.400 130.400 ;
        RECT 254.000 130.200 254.600 131.600 ;
        RECT 257.400 130.200 258.000 133.600 ;
        RECT 262.000 134.300 262.800 139.800 ;
        RECT 263.600 136.000 264.400 139.800 ;
        RECT 266.800 136.000 267.600 139.800 ;
        RECT 263.600 135.800 267.600 136.000 ;
        RECT 268.400 135.800 269.200 139.800 ;
        RECT 270.000 136.000 270.800 139.800 ;
        RECT 273.200 136.000 274.000 139.800 ;
        RECT 270.000 135.800 274.000 136.000 ;
        RECT 274.800 135.800 275.600 139.800 ;
        RECT 277.000 138.400 277.800 139.800 ;
        RECT 276.400 137.600 277.800 138.400 ;
        RECT 277.000 136.400 277.800 137.600 ;
        RECT 277.000 135.800 278.800 136.400 ;
        RECT 263.800 135.400 267.400 135.800 ;
        RECT 264.400 134.400 265.200 134.800 ;
        RECT 268.400 134.400 269.000 135.800 ;
        RECT 270.200 135.400 273.800 135.800 ;
        RECT 270.800 134.400 271.600 134.800 ;
        RECT 274.800 134.400 275.400 135.800 ;
        RECT 263.600 134.300 265.200 134.400 ;
        RECT 262.000 133.800 265.200 134.300 ;
        RECT 262.000 133.700 264.400 133.800 ;
        RECT 258.800 132.300 259.600 132.400 ;
        RECT 262.000 132.300 262.800 133.700 ;
        RECT 263.600 133.600 264.400 133.700 ;
        RECT 266.600 133.600 269.200 134.400 ;
        RECT 270.000 133.800 271.600 134.400 ;
        RECT 270.000 133.600 270.800 133.800 ;
        RECT 273.000 133.600 275.600 134.400 ;
        RECT 258.800 131.700 262.800 132.300 ;
        RECT 258.800 130.800 259.600 131.700 ;
        RECT 247.600 123.000 248.400 127.000 ;
        RECT 249.200 129.600 253.200 130.200 ;
        RECT 249.200 122.200 250.000 129.600 ;
        RECT 252.400 122.200 253.200 129.600 ;
        RECT 254.000 122.200 254.800 130.200 ;
        RECT 257.200 129.400 259.000 130.200 ;
        RECT 258.200 122.200 259.000 129.400 ;
        RECT 262.000 122.200 262.800 131.700 ;
        RECT 265.200 131.600 266.000 133.200 ;
        RECT 266.600 130.200 267.200 133.600 ;
        RECT 268.400 132.300 269.200 132.400 ;
        RECT 271.600 132.300 272.400 133.200 ;
        RECT 268.400 131.700 272.400 132.300 ;
        RECT 268.400 131.600 269.200 131.700 ;
        RECT 271.600 131.600 272.400 131.700 ;
        RECT 273.000 130.400 273.600 133.600 ;
        RECT 268.400 130.200 269.200 130.400 ;
        RECT 266.200 129.600 267.200 130.200 ;
        RECT 267.800 129.600 269.200 130.200 ;
        RECT 271.600 129.600 273.600 130.400 ;
        RECT 274.800 130.200 275.600 130.400 ;
        RECT 274.200 129.600 275.600 130.200 ;
        RECT 266.200 124.400 267.000 129.600 ;
        RECT 267.800 128.400 268.400 129.600 ;
        RECT 267.600 127.600 268.400 128.400 ;
        RECT 265.200 123.600 267.000 124.400 ;
        RECT 266.200 122.200 267.000 123.600 ;
        RECT 272.600 122.200 273.400 129.600 ;
        RECT 274.200 128.400 274.800 129.600 ;
        RECT 276.400 128.800 277.200 130.400 ;
        RECT 274.000 127.600 274.800 128.400 ;
        RECT 278.000 122.200 278.800 135.800 ;
        RECT 281.200 135.600 282.000 137.200 ;
        RECT 279.600 134.300 280.400 135.200 ;
        RECT 281.200 134.300 282.000 134.400 ;
        RECT 279.600 133.700 282.000 134.300 ;
        RECT 279.600 133.600 280.400 133.700 ;
        RECT 281.200 133.600 282.000 133.700 ;
        RECT 282.800 132.300 283.600 139.800 ;
        RECT 284.400 136.000 285.200 139.800 ;
        RECT 287.600 136.000 288.400 139.800 ;
        RECT 284.400 135.800 288.400 136.000 ;
        RECT 289.200 135.800 290.000 139.800 ;
        RECT 295.600 135.800 296.400 139.800 ;
        RECT 300.000 136.200 301.600 139.800 ;
        RECT 284.600 135.400 288.200 135.800 ;
        RECT 285.200 134.400 286.000 134.800 ;
        RECT 289.200 134.400 289.800 135.800 ;
        RECT 295.600 135.200 298.000 135.800 ;
        RECT 297.200 135.000 298.000 135.200 ;
        RECT 298.600 134.800 299.400 135.600 ;
        RECT 298.600 134.400 299.200 134.800 ;
        RECT 284.400 133.800 286.000 134.400 ;
        RECT 287.400 134.300 290.000 134.400 ;
        RECT 294.000 134.300 294.800 134.400 ;
        RECT 284.400 133.600 285.200 133.800 ;
        RECT 287.400 133.700 294.800 134.300 ;
        RECT 287.400 133.600 290.000 133.700 ;
        RECT 294.000 133.600 294.800 133.700 ;
        RECT 295.600 133.600 297.200 134.400 ;
        RECT 298.400 133.600 299.200 134.400 ;
        RECT 300.000 134.200 300.600 136.200 ;
        RECT 305.200 135.800 306.000 139.800 ;
        RECT 301.200 134.800 302.800 135.600 ;
        RECT 303.400 135.200 306.000 135.800 ;
        RECT 303.400 135.000 304.200 135.200 ;
        RECT 306.800 135.000 307.600 139.800 ;
        RECT 311.200 138.400 312.000 139.800 ;
        RECT 310.000 137.800 312.000 138.400 ;
        RECT 315.600 137.800 316.400 139.800 ;
        RECT 319.800 138.400 321.000 139.800 ;
        RECT 319.600 137.800 321.000 138.400 ;
        RECT 310.000 137.000 310.800 137.800 ;
        RECT 315.600 137.200 316.200 137.800 ;
        RECT 311.600 136.400 312.400 137.200 ;
        RECT 313.400 136.600 316.200 137.200 ;
        RECT 319.600 137.000 320.400 137.800 ;
        RECT 313.400 136.400 314.200 136.600 ;
        RECT 304.400 134.200 306.000 134.400 ;
        RECT 300.000 133.600 301.000 134.200 ;
        RECT 303.800 134.000 306.000 134.200 ;
        RECT 286.000 132.300 286.800 133.200 ;
        RECT 282.800 131.700 286.800 132.300 ;
        RECT 282.800 122.200 283.600 131.700 ;
        RECT 286.000 131.600 286.800 131.700 ;
        RECT 287.400 130.200 288.000 133.600 ;
        RECT 300.400 132.400 301.000 133.600 ;
        RECT 301.600 133.600 306.000 134.000 ;
        RECT 307.600 134.200 309.200 134.400 ;
        RECT 311.800 134.200 312.400 136.400 ;
        RECT 321.400 135.400 322.200 135.600 ;
        RECT 324.400 135.400 325.200 139.800 ;
        RECT 321.400 134.800 325.200 135.400 ;
        RECT 326.000 135.800 326.800 139.800 ;
        RECT 330.400 136.200 332.000 139.800 ;
        RECT 326.000 135.200 328.400 135.800 ;
        RECT 327.600 135.000 328.400 135.200 ;
        RECT 314.800 134.200 315.600 134.400 ;
        RECT 317.400 134.200 318.200 134.400 ;
        RECT 307.600 133.600 318.600 134.200 ;
        RECT 301.600 133.400 304.400 133.600 ;
        RECT 310.600 133.400 311.400 133.600 ;
        RECT 301.600 133.200 302.400 133.400 ;
        RECT 309.000 132.400 309.800 132.600 ;
        RECT 311.600 132.400 312.400 132.600 ;
        RECT 300.400 131.600 301.200 132.400 ;
        RECT 303.000 132.200 303.800 132.400 ;
        RECT 302.200 131.600 303.800 132.200 ;
        RECT 309.000 131.800 314.000 132.400 ;
        RECT 313.200 131.600 314.000 131.800 ;
        RECT 289.200 130.200 290.000 130.400 ;
        RECT 300.400 130.200 301.000 131.600 ;
        RECT 302.200 131.400 303.000 131.600 ;
        RECT 306.800 131.000 312.400 131.200 ;
        RECT 306.800 130.800 312.600 131.000 ;
        RECT 306.800 130.600 316.600 130.800 ;
        RECT 287.000 129.600 288.000 130.200 ;
        RECT 288.600 129.600 290.000 130.200 ;
        RECT 295.600 129.600 298.000 130.200 ;
        RECT 287.000 122.200 287.800 129.600 ;
        RECT 288.600 128.400 289.200 129.600 ;
        RECT 288.400 127.600 289.200 128.400 ;
        RECT 295.600 122.200 296.400 129.600 ;
        RECT 297.200 129.400 298.000 129.600 ;
        RECT 300.000 124.400 301.600 130.200 ;
        RECT 303.400 129.600 306.000 130.200 ;
        RECT 303.400 129.400 304.200 129.600 ;
        RECT 300.000 123.600 302.800 124.400 ;
        RECT 300.000 122.200 301.600 123.600 ;
        RECT 305.200 122.200 306.000 129.600 ;
        RECT 306.800 122.200 307.600 130.600 ;
        RECT 311.800 130.200 316.600 130.600 ;
        RECT 310.000 129.000 315.400 129.600 ;
        RECT 310.000 128.800 310.800 129.000 ;
        RECT 314.600 128.800 315.400 129.000 ;
        RECT 316.000 129.000 316.600 130.200 ;
        RECT 318.000 130.400 318.600 133.600 ;
        RECT 319.600 132.800 320.400 133.000 ;
        RECT 319.600 132.200 323.400 132.800 ;
        RECT 322.600 132.000 323.400 132.200 ;
        RECT 321.000 131.400 321.800 131.600 ;
        RECT 324.400 131.400 325.200 134.800 ;
        RECT 329.000 134.800 329.800 135.600 ;
        RECT 329.000 134.400 329.600 134.800 ;
        RECT 326.000 133.600 327.600 134.400 ;
        RECT 328.800 133.600 329.600 134.400 ;
        RECT 330.400 134.200 331.000 136.200 ;
        RECT 335.600 135.800 336.400 139.800 ;
        RECT 331.600 134.800 333.200 135.600 ;
        RECT 333.800 135.200 336.400 135.800 ;
        RECT 337.200 135.800 338.000 139.800 ;
        RECT 341.600 136.200 343.200 139.800 ;
        RECT 337.200 135.200 339.600 135.800 ;
        RECT 333.800 135.000 334.600 135.200 ;
        RECT 338.800 135.000 339.600 135.200 ;
        RECT 340.200 134.800 341.000 135.600 ;
        RECT 340.200 134.400 340.800 134.800 ;
        RECT 334.800 134.200 336.400 134.400 ;
        RECT 330.400 133.600 331.400 134.200 ;
        RECT 334.200 134.000 336.400 134.200 ;
        RECT 321.000 130.800 325.200 131.400 ;
        RECT 318.000 129.800 320.400 130.400 ;
        RECT 317.400 129.000 318.200 129.200 ;
        RECT 316.000 128.400 318.200 129.000 ;
        RECT 319.800 128.800 320.400 129.800 ;
        RECT 319.800 128.000 321.200 128.800 ;
        RECT 313.400 127.400 314.200 127.600 ;
        RECT 316.200 127.400 317.000 127.600 ;
        RECT 310.000 126.200 310.800 127.000 ;
        RECT 313.400 126.800 317.000 127.400 ;
        RECT 315.600 126.200 316.200 126.800 ;
        RECT 319.600 126.200 320.400 127.000 ;
        RECT 310.000 125.600 312.000 126.200 ;
        RECT 311.200 122.200 312.000 125.600 ;
        RECT 315.600 122.200 316.400 126.200 ;
        RECT 319.800 122.200 321.000 126.200 ;
        RECT 324.400 122.200 325.200 130.800 ;
        RECT 330.800 132.400 331.400 133.600 ;
        RECT 332.000 133.600 336.400 134.000 ;
        RECT 337.200 133.600 338.800 134.400 ;
        RECT 340.000 133.600 340.800 134.400 ;
        RECT 341.600 134.200 342.200 136.200 ;
        RECT 346.800 135.800 347.600 139.800 ;
        RECT 342.800 134.800 344.400 135.600 ;
        RECT 345.000 135.200 347.600 135.800 ;
        RECT 348.400 135.800 349.200 139.800 ;
        RECT 352.800 136.200 354.400 139.800 ;
        RECT 348.400 135.200 350.600 135.800 ;
        RECT 351.600 135.400 353.200 135.600 ;
        RECT 345.000 135.000 345.800 135.200 ;
        RECT 349.800 135.000 350.600 135.200 ;
        RECT 351.200 134.800 353.200 135.400 ;
        RECT 351.200 134.400 351.800 134.800 ;
        RECT 346.000 134.300 347.600 134.400 ;
        RECT 348.400 134.300 351.800 134.400 ;
        RECT 346.000 134.200 351.800 134.300 ;
        RECT 341.600 133.600 342.600 134.200 ;
        RECT 345.400 134.000 351.800 134.200 ;
        RECT 332.000 133.400 334.800 133.600 ;
        RECT 332.000 133.200 332.800 133.400 ;
        RECT 342.000 132.400 342.600 133.600 ;
        RECT 343.200 133.800 351.800 134.000 ;
        RECT 343.200 133.700 350.000 133.800 ;
        RECT 343.200 133.600 347.600 133.700 ;
        RECT 348.400 133.600 350.000 133.700 ;
        RECT 343.200 133.400 346.000 133.600 ;
        RECT 352.400 133.400 353.200 134.200 ;
        RECT 343.200 133.200 344.000 133.400 ;
        RECT 352.400 132.800 353.000 133.400 ;
        RECT 330.800 131.600 331.600 132.400 ;
        RECT 333.400 132.200 334.200 132.400 ;
        RECT 332.600 131.600 334.200 132.200 ;
        RECT 342.000 131.600 342.800 132.400 ;
        RECT 344.600 132.200 345.400 132.400 ;
        RECT 343.800 131.600 345.400 132.200 ;
        RECT 350.400 132.200 353.000 132.800 ;
        RECT 353.800 132.800 354.400 136.200 ;
        RECT 358.000 135.800 358.800 139.800 ;
        RECT 362.200 136.400 363.000 139.800 ;
        RECT 367.000 136.400 367.800 139.800 ;
        RECT 355.000 134.800 355.800 135.600 ;
        RECT 356.400 135.200 358.800 135.800 ;
        RECT 361.200 135.800 363.000 136.400 ;
        RECT 366.000 135.800 367.800 136.400 ;
        RECT 356.400 135.000 357.200 135.200 ;
        RECT 355.200 134.400 355.800 134.800 ;
        RECT 355.200 133.600 356.000 134.400 ;
        RECT 357.200 133.600 358.800 134.400 ;
        RECT 359.600 133.600 360.400 135.200 ;
        RECT 361.200 134.300 362.000 135.800 ;
        RECT 364.400 134.300 365.200 135.200 ;
        RECT 361.200 133.700 365.200 134.300 ;
        RECT 353.800 132.400 354.800 132.800 ;
        RECT 353.800 132.200 355.600 132.400 ;
        RECT 350.400 132.000 351.200 132.200 ;
        RECT 354.200 131.600 355.600 132.200 ;
        RECT 358.000 132.300 358.800 132.400 ;
        RECT 359.700 132.300 360.300 133.600 ;
        RECT 358.000 131.700 360.300 132.300 ;
        RECT 358.000 131.600 358.800 131.700 ;
        RECT 330.800 130.200 331.400 131.600 ;
        RECT 332.600 131.400 333.400 131.600 ;
        RECT 342.000 130.400 342.600 131.600 ;
        RECT 343.800 131.400 344.600 131.600 ;
        RECT 352.600 131.400 353.400 131.600 ;
        RECT 350.000 130.800 353.400 131.400 ;
        RECT 342.000 130.200 344.400 130.400 ;
        RECT 350.000 130.200 350.600 130.800 ;
        RECT 354.200 130.200 354.800 131.600 ;
        RECT 326.000 129.600 328.400 130.200 ;
        RECT 326.000 122.200 326.800 129.600 ;
        RECT 327.600 129.400 328.400 129.600 ;
        RECT 330.400 126.400 332.000 130.200 ;
        RECT 333.800 129.600 336.400 130.200 ;
        RECT 333.800 129.400 334.600 129.600 ;
        RECT 330.400 125.600 333.200 126.400 ;
        RECT 330.400 122.200 332.000 125.600 ;
        RECT 335.600 122.200 336.400 129.600 ;
        RECT 337.200 129.600 339.600 130.200 ;
        RECT 337.200 122.200 338.000 129.600 ;
        RECT 338.800 129.400 339.600 129.600 ;
        RECT 341.600 129.600 344.400 130.200 ;
        RECT 345.000 129.600 347.600 130.200 ;
        RECT 341.600 122.200 343.200 129.600 ;
        RECT 345.000 129.400 345.800 129.600 ;
        RECT 346.800 122.200 347.600 129.600 ;
        RECT 348.400 129.600 350.600 130.200 ;
        RECT 348.400 122.200 349.200 129.600 ;
        RECT 349.800 129.400 350.600 129.600 ;
        RECT 352.800 129.600 354.800 130.200 ;
        RECT 356.400 129.600 358.800 130.200 ;
        RECT 352.800 122.200 354.400 129.600 ;
        RECT 356.400 129.400 357.200 129.600 ;
        RECT 358.000 122.200 358.800 129.600 ;
        RECT 361.200 122.200 362.000 133.700 ;
        RECT 364.400 133.600 365.200 133.700 ;
        RECT 362.800 130.300 363.600 130.400 ;
        RECT 364.400 130.300 365.200 130.400 ;
        RECT 362.800 129.700 365.200 130.300 ;
        RECT 362.800 128.800 363.600 129.700 ;
        RECT 364.400 129.600 365.200 129.700 ;
        RECT 366.000 122.200 366.800 135.800 ;
        RECT 369.200 135.600 370.000 137.200 ;
        RECT 367.600 128.800 368.400 130.400 ;
        RECT 370.800 130.300 371.600 139.800 ;
        RECT 373.000 136.400 373.800 139.800 ;
        RECT 373.000 135.800 374.800 136.400 ;
        RECT 372.400 134.300 373.200 134.400 ;
        RECT 374.000 134.300 374.800 135.800 ;
        RECT 377.200 135.600 378.000 137.200 ;
        RECT 372.400 133.700 374.800 134.300 ;
        RECT 372.400 133.600 373.200 133.700 ;
        RECT 372.400 130.300 373.200 130.400 ;
        RECT 370.800 129.700 373.200 130.300 ;
        RECT 370.800 122.200 371.600 129.700 ;
        RECT 372.400 128.800 373.200 129.700 ;
        RECT 374.000 122.200 374.800 133.700 ;
        RECT 375.600 133.600 376.400 135.200 ;
        RECT 378.800 122.200 379.600 139.800 ;
        RECT 381.000 138.400 381.800 139.800 ;
        RECT 380.400 137.600 381.800 138.400 ;
        RECT 381.000 136.400 381.800 137.600 ;
        RECT 385.800 138.400 386.600 139.800 ;
        RECT 392.600 138.400 393.400 139.800 ;
        RECT 385.800 137.600 387.600 138.400 ;
        RECT 392.600 137.600 394.000 138.400 ;
        RECT 396.400 137.800 397.200 139.800 ;
        RECT 402.200 138.400 403.800 139.800 ;
        RECT 385.800 136.400 386.600 137.600 ;
        RECT 392.600 136.400 393.400 137.600 ;
        RECT 381.000 135.800 382.800 136.400 ;
        RECT 385.800 135.800 387.600 136.400 ;
        RECT 380.400 128.800 381.200 130.400 ;
        RECT 382.000 122.200 382.800 135.800 ;
        RECT 383.600 134.300 384.400 135.200 ;
        RECT 385.200 134.300 386.000 134.400 ;
        RECT 383.600 133.700 386.000 134.300 ;
        RECT 383.600 133.600 384.400 133.700 ;
        RECT 385.200 133.600 386.000 133.700 ;
        RECT 383.600 130.300 384.400 130.400 ;
        RECT 385.200 130.300 386.000 130.400 ;
        RECT 383.600 129.700 386.000 130.300 ;
        RECT 383.600 129.600 384.400 129.700 ;
        RECT 385.200 128.800 386.000 129.700 ;
        RECT 386.800 122.200 387.600 135.800 ;
        RECT 391.600 135.800 393.400 136.400 ;
        RECT 388.400 133.600 389.200 135.200 ;
        RECT 390.000 133.600 390.800 135.200 ;
        RECT 391.600 122.200 392.400 135.800 ;
        RECT 396.400 134.400 397.000 137.800 ;
        RECT 401.200 137.600 403.800 138.400 ;
        RECT 398.000 135.600 398.800 137.200 ;
        RECT 402.200 135.800 403.800 137.600 ;
        RECT 410.600 135.800 412.200 139.800 ;
        RECT 417.200 137.800 418.000 139.800 ;
        RECT 396.400 134.300 397.200 134.400 ;
        RECT 401.200 134.300 402.000 134.400 ;
        RECT 396.400 133.700 402.000 134.300 ;
        RECT 396.400 133.600 397.200 133.700 ;
        RECT 401.200 133.600 402.000 133.700 ;
        RECT 394.800 132.300 395.600 132.400 ;
        RECT 393.300 131.700 395.600 132.300 ;
        RECT 393.300 130.400 393.900 131.700 ;
        RECT 394.800 130.800 395.600 131.700 ;
        RECT 393.200 128.800 394.000 130.400 ;
        RECT 396.400 130.200 397.000 133.600 ;
        RECT 401.400 133.200 402.000 133.600 ;
        RECT 401.400 132.400 402.200 133.200 ;
        RECT 402.800 132.400 403.400 135.800 ;
        RECT 404.400 134.300 405.200 134.400 ;
        RECT 409.200 134.300 410.000 134.400 ;
        RECT 404.400 133.700 410.000 134.300 ;
        RECT 404.400 132.800 405.200 133.700 ;
        RECT 409.200 132.800 410.000 133.700 ;
        RECT 411.000 132.400 411.600 135.800 ;
        RECT 417.200 134.400 417.800 137.800 ;
        RECT 418.800 135.600 419.600 137.200 ;
        RECT 420.400 135.800 421.200 139.800 ;
        RECT 424.800 138.400 426.400 139.800 ;
        RECT 424.800 137.600 427.600 138.400 ;
        RECT 424.800 136.200 426.400 137.600 ;
        RECT 420.400 135.200 422.800 135.800 ;
        RECT 422.000 135.000 422.800 135.200 ;
        RECT 423.400 134.800 424.200 135.600 ;
        RECT 423.400 134.400 424.000 134.800 ;
        RECT 412.400 134.300 413.200 134.400 ;
        RECT 417.200 134.300 418.000 134.400 ;
        RECT 412.400 133.700 418.000 134.300 ;
        RECT 412.400 133.600 413.200 133.700 ;
        RECT 417.200 133.600 418.000 133.700 ;
        RECT 420.400 133.600 422.000 134.400 ;
        RECT 423.200 133.600 424.000 134.400 ;
        RECT 412.400 133.200 413.000 133.600 ;
        RECT 412.200 132.400 413.000 133.200 ;
        RECT 399.600 130.800 400.400 132.400 ;
        RECT 402.800 131.600 403.600 132.400 ;
        RECT 406.000 132.200 406.800 132.400 ;
        RECT 405.200 131.600 406.800 132.200 ;
        RECT 407.600 132.200 408.400 132.400 ;
        RECT 407.600 131.600 409.200 132.200 ;
        RECT 410.800 131.600 411.600 132.400 ;
        RECT 402.800 131.400 403.400 131.600 ;
        RECT 401.400 130.800 403.400 131.400 ;
        RECT 405.200 131.200 406.000 131.600 ;
        RECT 408.400 131.200 409.200 131.600 ;
        RECT 411.000 131.400 411.600 131.600 ;
        RECT 411.000 130.800 413.000 131.400 ;
        RECT 414.000 130.800 414.800 132.400 ;
        RECT 415.600 130.800 416.400 132.400 ;
        RECT 401.400 130.200 402.000 130.800 ;
        RECT 412.400 130.200 413.000 130.800 ;
        RECT 417.200 130.200 417.800 133.600 ;
        RECT 424.800 132.800 425.400 136.200 ;
        RECT 430.000 135.800 430.800 139.800 ;
        RECT 431.600 135.800 432.400 139.800 ;
        RECT 433.200 136.000 434.000 139.800 ;
        RECT 436.400 136.000 437.200 139.800 ;
        RECT 439.600 137.800 440.400 139.800 ;
        RECT 433.200 135.800 437.200 136.000 ;
        RECT 426.000 135.400 427.600 135.600 ;
        RECT 426.000 134.800 428.000 135.400 ;
        RECT 428.600 135.200 430.800 135.800 ;
        RECT 428.600 135.000 429.400 135.200 ;
        RECT 427.400 134.400 428.000 134.800 ;
        RECT 431.800 134.400 432.400 135.800 ;
        RECT 433.400 135.400 437.000 135.800 ;
        RECT 438.000 135.600 438.800 137.200 ;
        RECT 439.800 136.300 440.400 137.800 ;
        RECT 449.200 137.600 450.000 139.800 ;
        RECT 454.000 137.600 454.800 139.800 ;
        RECT 447.600 136.300 448.400 137.200 ;
        RECT 439.700 135.700 448.400 136.300 ;
        RECT 435.600 134.400 436.400 134.800 ;
        RECT 438.100 134.400 438.700 135.600 ;
        RECT 439.800 134.400 440.400 135.700 ;
        RECT 447.600 135.600 448.400 135.700 ;
        RECT 449.400 134.400 450.000 137.600 ;
        RECT 452.400 135.600 453.200 137.200 ;
        RECT 454.200 134.400 454.800 137.600 ;
        RECT 457.200 136.000 458.000 139.800 ;
        RECT 460.400 136.000 461.200 139.800 ;
        RECT 457.200 135.800 461.200 136.000 ;
        RECT 462.000 136.300 462.800 139.800 ;
        RECT 463.600 136.300 464.400 137.200 ;
        RECT 457.400 135.400 461.000 135.800 ;
        RECT 462.000 135.700 464.400 136.300 ;
        RECT 458.000 134.400 458.800 134.800 ;
        RECT 462.000 134.400 462.600 135.700 ;
        RECT 463.600 135.600 464.400 135.700 ;
        RECT 426.000 133.400 426.800 134.200 ;
        RECT 427.400 133.800 430.800 134.400 ;
        RECT 429.200 133.600 430.800 133.800 ;
        RECT 431.600 133.600 434.200 134.400 ;
        RECT 435.600 134.300 437.200 134.400 ;
        RECT 438.000 134.300 438.800 134.400 ;
        RECT 435.600 133.800 438.800 134.300 ;
        RECT 436.400 133.700 438.800 133.800 ;
        RECT 436.400 133.600 437.200 133.700 ;
        RECT 438.000 133.600 438.800 133.700 ;
        RECT 439.600 133.600 440.400 134.400 ;
        RECT 449.200 133.600 450.000 134.400 ;
        RECT 454.000 133.600 454.800 134.400 ;
        RECT 457.200 133.800 458.800 134.400 ;
        RECT 457.200 133.600 458.000 133.800 ;
        RECT 460.200 133.600 462.800 134.400 ;
        RECT 424.400 132.400 425.400 132.800 ;
        RECT 423.600 132.200 425.400 132.400 ;
        RECT 426.200 132.800 426.800 133.400 ;
        RECT 426.200 132.200 428.800 132.800 ;
        RECT 423.600 131.600 425.000 132.200 ;
        RECT 428.000 132.000 428.800 132.200 ;
        RECT 424.400 130.200 425.000 131.600 ;
        RECT 425.800 131.400 426.600 131.600 ;
        RECT 425.800 130.800 429.200 131.400 ;
        RECT 428.600 130.200 429.200 130.800 ;
        RECT 431.600 130.200 432.400 130.400 ;
        RECT 433.600 130.200 434.200 133.600 ;
        RECT 434.800 131.600 435.600 133.200 ;
        RECT 439.800 130.200 440.400 133.600 ;
        RECT 441.200 130.800 442.000 132.400 ;
        RECT 449.400 130.200 450.000 133.600 ;
        RECT 450.800 132.300 451.600 132.400 ;
        RECT 454.200 132.300 454.800 133.600 ;
        RECT 450.800 131.700 454.800 132.300 ;
        RECT 450.800 130.800 451.600 131.700 ;
        RECT 454.200 130.200 454.800 131.700 ;
        RECT 455.600 132.300 456.400 132.400 ;
        RECT 458.800 132.300 459.600 133.200 ;
        RECT 455.600 131.700 459.600 132.300 ;
        RECT 455.600 130.800 456.400 131.700 ;
        RECT 458.800 131.600 459.600 131.700 ;
        RECT 460.200 130.200 460.800 133.600 ;
        RECT 462.000 130.300 462.800 130.400 ;
        RECT 463.600 130.300 464.400 130.400 ;
        RECT 462.000 130.200 464.400 130.300 ;
        RECT 395.400 129.400 397.200 130.200 ;
        RECT 395.400 122.200 396.200 129.400 ;
        RECT 399.600 122.800 400.400 130.200 ;
        RECT 401.200 123.400 402.000 130.200 ;
        RECT 402.800 129.600 406.800 130.200 ;
        RECT 402.800 122.800 403.600 129.600 ;
        RECT 399.600 122.200 403.600 122.800 ;
        RECT 406.000 122.200 406.800 129.600 ;
        RECT 407.600 129.600 411.600 130.200 ;
        RECT 407.600 122.200 408.400 129.600 ;
        RECT 410.800 122.800 411.600 129.600 ;
        RECT 412.400 123.400 413.200 130.200 ;
        RECT 414.000 122.800 414.800 130.200 ;
        RECT 410.800 122.200 414.800 122.800 ;
        RECT 416.200 129.400 418.000 130.200 ;
        RECT 420.400 129.600 422.800 130.200 ;
        RECT 424.400 129.600 426.400 130.200 ;
        RECT 416.200 122.200 417.000 129.400 ;
        RECT 420.400 122.200 421.200 129.600 ;
        RECT 422.000 129.400 422.800 129.600 ;
        RECT 424.800 122.200 426.400 129.600 ;
        RECT 428.600 129.600 430.800 130.200 ;
        RECT 431.600 129.600 433.000 130.200 ;
        RECT 433.600 129.600 434.600 130.200 ;
        RECT 428.600 129.400 429.400 129.600 ;
        RECT 430.000 122.200 430.800 129.600 ;
        RECT 432.400 128.400 433.000 129.600 ;
        RECT 432.400 127.600 433.200 128.400 ;
        RECT 433.800 122.200 434.600 129.600 ;
        RECT 439.600 129.400 441.400 130.200 ;
        RECT 449.200 129.400 451.000 130.200 ;
        RECT 454.000 129.400 455.800 130.200 ;
        RECT 440.600 122.200 441.400 129.400 ;
        RECT 450.200 122.200 451.000 129.400 ;
        RECT 455.000 122.200 455.800 129.400 ;
        RECT 459.800 129.600 460.800 130.200 ;
        RECT 461.400 129.700 464.400 130.200 ;
        RECT 461.400 129.600 462.800 129.700 ;
        RECT 463.600 129.600 464.400 129.700 ;
        RECT 459.800 122.200 460.600 129.600 ;
        RECT 461.400 128.400 462.000 129.600 ;
        RECT 461.200 127.600 462.000 128.400 ;
        RECT 465.200 122.200 466.000 139.800 ;
        RECT 466.800 136.000 467.600 139.800 ;
        RECT 470.000 136.000 470.800 139.800 ;
        RECT 466.800 135.800 470.800 136.000 ;
        RECT 471.600 135.800 472.400 139.800 ;
        RECT 474.800 138.300 475.600 138.400 ;
        RECT 476.800 138.300 477.600 139.800 ;
        RECT 474.800 137.700 477.600 138.300 ;
        RECT 474.800 137.600 475.600 137.700 ;
        RECT 467.000 135.400 470.600 135.800 ;
        RECT 467.600 134.400 468.400 134.800 ;
        RECT 471.600 134.400 472.200 135.800 ;
        RECT 466.800 133.800 468.400 134.400 ;
        RECT 466.800 133.600 467.600 133.800 ;
        RECT 469.800 133.600 472.400 134.400 ;
        RECT 476.800 134.200 477.600 137.700 ;
        RECT 479.600 135.400 480.400 139.800 ;
        RECT 483.800 138.400 485.000 139.800 ;
        RECT 483.800 137.800 485.200 138.400 ;
        RECT 488.400 137.800 489.200 139.800 ;
        RECT 492.800 138.400 493.600 139.800 ;
        RECT 492.800 137.800 494.800 138.400 ;
        RECT 484.400 137.000 485.200 137.800 ;
        RECT 488.600 137.200 489.200 137.800 ;
        RECT 488.600 136.600 491.400 137.200 ;
        RECT 490.600 136.400 491.400 136.600 ;
        RECT 492.400 136.400 493.200 137.200 ;
        RECT 494.000 137.000 494.800 137.800 ;
        RECT 482.600 135.400 483.400 135.600 ;
        RECT 479.600 134.800 483.400 135.400 ;
        RECT 476.800 133.800 478.600 134.200 ;
        RECT 477.000 133.600 478.600 133.800 ;
        RECT 468.400 131.600 469.200 133.200 ;
        RECT 469.800 132.300 470.400 133.600 ;
        RECT 471.600 132.300 472.400 132.400 ;
        RECT 469.800 131.700 472.400 132.300 ;
        RECT 469.800 130.200 470.400 131.700 ;
        RECT 471.600 131.600 472.400 131.700 ;
        RECT 474.800 131.600 476.400 132.400 ;
        RECT 471.600 130.200 472.400 130.400 ;
        RECT 469.400 129.600 470.400 130.200 ;
        RECT 471.000 129.600 472.400 130.200 ;
        RECT 473.200 129.600 474.000 131.200 ;
        RECT 478.000 130.400 478.600 133.600 ;
        RECT 479.600 131.400 480.400 134.800 ;
        RECT 486.600 134.200 487.400 134.400 ;
        RECT 492.400 134.200 493.000 136.400 ;
        RECT 497.200 135.000 498.000 139.800 ;
        RECT 500.400 135.200 501.200 139.800 ;
        RECT 503.600 135.200 504.400 139.800 ;
        RECT 506.800 135.200 507.600 139.800 ;
        RECT 510.000 135.200 510.800 139.800 ;
        RECT 515.800 138.400 516.600 139.800 ;
        RECT 514.800 137.600 516.600 138.400 ;
        RECT 515.800 136.400 516.600 137.600 ;
        RECT 520.600 138.400 521.400 139.800 ;
        RECT 520.600 137.600 522.000 138.400 ;
        RECT 520.600 136.400 521.400 137.600 ;
        RECT 525.400 136.400 526.200 139.800 ;
        RECT 514.800 135.800 516.600 136.400 ;
        RECT 519.600 135.800 521.400 136.400 ;
        RECT 524.400 135.800 526.200 136.400 ;
        RECT 500.400 134.400 502.200 135.200 ;
        RECT 503.600 134.400 505.800 135.200 ;
        RECT 506.800 134.400 509.000 135.200 ;
        RECT 510.000 134.400 512.400 135.200 ;
        RECT 495.600 134.200 497.200 134.400 ;
        RECT 486.200 133.600 497.200 134.200 ;
        RECT 501.400 133.800 502.200 134.400 ;
        RECT 505.000 133.800 505.800 134.400 ;
        RECT 508.200 133.800 509.000 134.400 ;
        RECT 484.400 132.800 485.200 133.000 ;
        RECT 481.400 132.200 485.200 132.800 ;
        RECT 481.400 132.000 482.200 132.200 ;
        RECT 483.000 131.400 483.800 131.600 ;
        RECT 479.600 130.800 483.800 131.400 ;
        RECT 478.000 129.600 478.800 130.400 ;
        RECT 469.400 122.200 470.200 129.600 ;
        RECT 471.000 128.400 471.600 129.600 ;
        RECT 470.800 127.600 471.600 128.400 ;
        RECT 476.400 127.600 477.200 129.200 ;
        RECT 478.000 127.000 478.600 129.600 ;
        RECT 475.000 126.400 478.600 127.000 ;
        RECT 475.000 126.200 475.600 126.400 ;
        RECT 474.800 122.200 475.600 126.200 ;
        RECT 478.000 126.200 478.600 126.400 ;
        RECT 478.000 122.200 478.800 126.200 ;
        RECT 479.600 122.200 480.400 130.800 ;
        RECT 486.200 130.400 486.800 133.600 ;
        RECT 493.400 133.400 494.200 133.600 ;
        RECT 501.400 133.000 504.000 133.800 ;
        RECT 505.000 133.000 507.400 133.800 ;
        RECT 508.200 133.000 510.800 133.800 ;
        RECT 495.000 132.400 495.800 132.600 ;
        RECT 490.800 131.800 495.800 132.400 ;
        RECT 490.800 131.600 491.600 131.800 ;
        RECT 501.400 131.600 502.200 133.000 ;
        RECT 505.000 131.600 505.800 133.000 ;
        RECT 508.200 131.600 509.000 133.000 ;
        RECT 511.600 131.600 512.400 134.400 ;
        RECT 513.200 133.600 514.000 135.200 ;
        RECT 514.800 134.300 515.600 135.800 ;
        RECT 518.000 134.300 518.800 135.200 ;
        RECT 514.800 133.700 518.800 134.300 ;
        RECT 492.400 131.000 498.000 131.200 ;
        RECT 492.200 130.800 498.000 131.000 ;
        RECT 484.400 129.800 486.800 130.400 ;
        RECT 488.200 130.600 498.000 130.800 ;
        RECT 488.200 130.200 493.000 130.600 ;
        RECT 484.400 128.800 485.000 129.800 ;
        RECT 483.600 128.000 485.000 128.800 ;
        RECT 486.600 129.000 487.400 129.200 ;
        RECT 488.200 129.000 488.800 130.200 ;
        RECT 486.600 128.400 488.800 129.000 ;
        RECT 489.400 129.000 494.800 129.600 ;
        RECT 489.400 128.800 490.200 129.000 ;
        RECT 494.000 128.800 494.800 129.000 ;
        RECT 487.800 127.400 488.600 127.600 ;
        RECT 490.600 127.400 491.400 127.600 ;
        RECT 484.400 126.200 485.200 127.000 ;
        RECT 487.800 126.800 491.400 127.400 ;
        RECT 488.600 126.200 489.200 126.800 ;
        RECT 494.000 126.200 494.800 127.000 ;
        RECT 483.800 122.200 485.000 126.200 ;
        RECT 488.400 122.200 489.200 126.200 ;
        RECT 492.800 125.600 494.800 126.200 ;
        RECT 492.800 122.200 493.600 125.600 ;
        RECT 497.200 122.200 498.000 130.600 ;
        RECT 500.400 130.800 502.200 131.600 ;
        RECT 503.600 130.800 505.800 131.600 ;
        RECT 506.800 130.800 509.000 131.600 ;
        RECT 510.000 130.800 512.400 131.600 ;
        RECT 500.400 122.200 501.200 130.800 ;
        RECT 503.600 122.200 504.400 130.800 ;
        RECT 506.800 122.200 507.600 130.800 ;
        RECT 510.000 122.200 510.800 130.800 ;
        RECT 514.800 122.200 515.600 133.700 ;
        RECT 518.000 133.600 518.800 133.700 ;
        RECT 516.400 128.800 517.200 130.400 ;
        RECT 519.600 122.200 520.400 135.800 ;
        RECT 522.800 133.600 523.600 135.200 ;
        RECT 521.200 130.300 522.000 130.400 ;
        RECT 524.400 130.300 525.200 135.800 ;
        RECT 527.600 133.600 528.400 135.200 ;
        RECT 521.200 129.700 525.200 130.300 ;
        RECT 521.200 128.800 522.000 129.700 ;
        RECT 524.400 122.200 525.200 129.700 ;
        RECT 526.000 128.800 526.800 130.400 ;
        RECT 529.200 122.200 530.000 139.800 ;
        RECT 535.000 138.400 535.800 139.800 ;
        RECT 534.000 137.600 535.800 138.400 ;
        RECT 535.000 136.400 535.800 137.600 ;
        RECT 534.000 135.800 535.800 136.400 ;
        RECT 532.400 133.600 533.200 135.200 ;
        RECT 534.000 122.200 534.800 135.800 ;
        RECT 535.600 130.300 536.400 130.400 ;
        RECT 537.200 130.300 538.000 139.800 ;
        RECT 541.000 138.400 541.800 139.800 ;
        RECT 540.400 137.600 541.800 138.400 ;
        RECT 538.800 135.600 539.600 137.200 ;
        RECT 541.000 136.400 541.800 137.600 ;
        RECT 541.000 135.800 542.800 136.400 ;
        RECT 535.600 129.700 538.000 130.300 ;
        RECT 535.600 128.800 536.400 129.700 ;
        RECT 537.200 122.200 538.000 129.700 ;
        RECT 540.400 128.800 541.200 130.400 ;
        RECT 542.000 122.200 542.800 135.800 ;
        RECT 545.200 135.800 546.000 139.800 ;
        RECT 548.400 137.800 549.200 139.800 ;
        RECT 543.600 133.600 544.400 135.200 ;
        RECT 545.200 132.400 545.800 135.800 ;
        RECT 548.400 135.600 549.000 137.800 ;
        RECT 550.000 135.600 550.800 137.200 ;
        RECT 546.600 135.000 549.000 135.600 ;
        RECT 545.200 131.600 546.000 132.400 ;
        RECT 546.600 132.000 547.200 135.000 ;
        RECT 548.200 133.600 549.200 134.400 ;
        RECT 548.000 132.800 548.800 133.600 ;
        RECT 551.600 132.400 552.400 139.800 ;
        RECT 554.800 135.200 555.600 139.800 ;
        RECT 556.400 135.800 557.200 139.800 ;
        RECT 560.800 136.200 562.400 139.800 ;
        RECT 556.400 135.200 558.800 135.800 ;
        RECT 553.400 134.600 555.600 135.200 ;
        RECT 558.000 135.000 558.800 135.200 ;
        RECT 559.400 134.800 560.200 135.600 ;
        RECT 543.600 130.300 544.400 130.400 ;
        RECT 545.200 130.300 545.800 131.600 ;
        RECT 546.600 131.400 547.400 132.000 ;
        RECT 546.600 131.200 550.800 131.400 ;
        RECT 546.800 130.800 550.800 131.200 ;
        RECT 543.600 130.200 545.900 130.300 ;
        RECT 543.600 129.700 546.600 130.200 ;
        RECT 543.600 129.600 544.400 129.700 ;
        RECT 545.200 129.600 546.600 129.700 ;
        RECT 545.800 122.200 546.600 129.600 ;
        RECT 550.000 122.200 550.800 130.800 ;
        RECT 551.600 130.200 552.200 132.400 ;
        RECT 553.400 131.600 554.000 134.600 ;
        RECT 559.400 134.400 560.000 134.800 ;
        RECT 556.400 133.600 558.000 134.400 ;
        RECT 559.200 133.600 560.000 134.400 ;
        RECT 560.800 134.200 561.400 136.200 ;
        RECT 566.000 135.800 566.800 139.800 ;
        RECT 562.000 134.800 563.600 135.600 ;
        RECT 564.200 135.200 566.800 135.800 ;
        RECT 567.600 135.800 568.400 139.800 ;
        RECT 572.000 138.400 573.600 139.800 ;
        RECT 570.800 137.600 573.600 138.400 ;
        RECT 572.000 136.200 573.600 137.600 ;
        RECT 567.600 135.200 570.000 135.800 ;
        RECT 564.200 135.000 565.000 135.200 ;
        RECT 569.200 135.000 570.000 135.200 ;
        RECT 570.600 134.800 571.400 135.600 ;
        RECT 570.600 134.400 571.200 134.800 ;
        RECT 565.200 134.200 566.800 134.400 ;
        RECT 560.800 133.600 561.800 134.200 ;
        RECT 564.600 134.000 566.800 134.200 ;
        RECT 552.800 130.800 554.000 131.600 ;
        RECT 553.400 130.200 554.000 130.800 ;
        RECT 561.200 132.400 561.800 133.600 ;
        RECT 562.400 133.600 566.800 134.000 ;
        RECT 567.600 133.600 569.200 134.400 ;
        RECT 570.400 133.600 571.200 134.400 ;
        RECT 572.000 134.200 572.600 136.200 ;
        RECT 577.200 135.800 578.000 139.800 ;
        RECT 573.200 134.800 574.800 135.600 ;
        RECT 575.400 135.200 578.000 135.800 ;
        RECT 578.800 135.200 579.600 139.800 ;
        RECT 575.400 135.000 576.200 135.200 ;
        RECT 578.800 134.600 581.000 135.200 ;
        RECT 576.400 134.200 578.000 134.400 ;
        RECT 572.000 133.600 573.000 134.200 ;
        RECT 575.800 134.000 578.000 134.200 ;
        RECT 562.400 133.400 565.200 133.600 ;
        RECT 562.400 133.200 563.200 133.400 ;
        RECT 572.400 132.400 573.000 133.600 ;
        RECT 573.600 133.600 578.000 134.000 ;
        RECT 573.600 133.400 576.400 133.600 ;
        RECT 573.600 133.200 574.400 133.400 ;
        RECT 561.200 131.600 562.000 132.400 ;
        RECT 563.800 132.200 564.600 132.400 ;
        RECT 563.000 131.600 564.600 132.200 ;
        RECT 572.400 131.600 573.200 132.400 ;
        RECT 575.000 132.200 575.800 132.400 ;
        RECT 574.200 131.600 575.800 132.200 ;
        RECT 580.400 131.600 581.000 134.600 ;
        RECT 582.000 132.400 582.800 139.800 ;
        RECT 561.200 130.200 561.800 131.600 ;
        RECT 563.000 131.400 563.800 131.600 ;
        RECT 572.400 130.200 573.000 131.600 ;
        RECT 574.200 131.400 575.000 131.600 ;
        RECT 580.400 130.800 581.600 131.600 ;
        RECT 580.400 130.200 581.000 130.800 ;
        RECT 582.200 130.200 582.800 132.400 ;
        RECT 551.600 122.200 552.400 130.200 ;
        RECT 553.400 129.600 555.600 130.200 ;
        RECT 554.800 122.200 555.600 129.600 ;
        RECT 556.400 129.600 558.800 130.200 ;
        RECT 556.400 122.200 557.200 129.600 ;
        RECT 558.000 129.400 558.800 129.600 ;
        RECT 560.800 124.400 562.400 130.200 ;
        RECT 564.200 129.600 566.800 130.200 ;
        RECT 564.200 129.400 565.000 129.600 ;
        RECT 559.600 123.600 562.400 124.400 ;
        RECT 560.800 122.200 562.400 123.600 ;
        RECT 566.000 122.200 566.800 129.600 ;
        RECT 567.600 129.600 570.000 130.200 ;
        RECT 567.600 122.200 568.400 129.600 ;
        RECT 569.200 129.400 570.000 129.600 ;
        RECT 572.000 122.200 573.600 130.200 ;
        RECT 575.400 129.600 578.000 130.200 ;
        RECT 575.400 129.400 576.200 129.600 ;
        RECT 577.200 122.200 578.000 129.600 ;
        RECT 578.800 129.600 581.000 130.200 ;
        RECT 578.800 122.200 579.600 129.600 ;
        RECT 582.000 122.200 582.800 130.200 ;
        RECT 3.800 112.400 4.600 119.800 ;
        RECT 5.200 113.600 6.000 114.400 ;
        RECT 5.400 112.400 6.000 113.600 ;
        RECT 7.600 112.400 8.400 119.800 ;
        RECT 10.800 119.200 14.800 119.800 ;
        RECT 10.800 112.400 11.600 119.200 ;
        RECT 3.800 111.800 4.800 112.400 ;
        RECT 5.400 111.800 6.800 112.400 ;
        RECT 7.600 111.800 11.600 112.400 ;
        RECT 12.400 111.800 13.200 118.600 ;
        RECT 14.000 111.800 14.800 119.200 ;
        RECT 15.600 111.800 16.400 119.800 ;
        RECT 17.200 112.400 18.000 119.800 ;
        RECT 20.400 112.400 21.200 119.800 ;
        RECT 17.200 111.800 21.200 112.400 ;
        RECT 22.000 112.400 22.800 119.800 ;
        RECT 23.400 112.400 24.200 112.600 ;
        RECT 22.000 111.800 24.200 112.400 ;
        RECT 26.400 112.400 28.000 119.800 ;
        RECT 30.000 112.400 30.800 112.600 ;
        RECT 31.600 112.400 32.400 119.800 ;
        RECT 35.800 112.600 36.600 119.800 ;
        RECT 26.400 111.800 28.400 112.400 ;
        RECT 30.000 111.800 32.400 112.400 ;
        RECT 34.800 111.800 36.600 112.600 ;
        RECT 2.800 108.800 3.600 110.400 ;
        RECT 4.200 108.400 4.800 111.800 ;
        RECT 6.000 111.600 6.800 111.800 ;
        RECT 12.400 111.200 13.000 111.800 ;
        RECT 8.400 110.400 9.200 110.800 ;
        RECT 11.000 110.600 13.000 111.200 ;
        RECT 11.000 110.400 11.600 110.600 ;
        RECT 7.600 109.800 9.200 110.400 ;
        RECT 7.600 109.600 8.400 109.800 ;
        RECT 10.800 109.600 11.600 110.400 ;
        RECT 14.000 109.600 14.800 111.200 ;
        RECT 15.800 110.400 16.400 111.800 ;
        RECT 23.600 111.200 24.200 111.800 ;
        RECT 19.600 110.400 20.400 110.800 ;
        RECT 23.600 110.600 27.000 111.200 ;
        RECT 26.200 110.400 27.000 110.600 ;
        RECT 27.800 110.400 28.400 111.800 ;
        RECT 15.600 109.800 18.000 110.400 ;
        RECT 19.600 110.300 21.200 110.400 ;
        RECT 22.000 110.300 22.800 110.400 ;
        RECT 19.600 109.800 22.800 110.300 ;
        RECT 27.800 110.300 29.200 110.400 ;
        RECT 31.600 110.300 32.400 110.400 ;
        RECT 15.600 109.600 16.400 109.800 ;
        RECT 1.200 108.200 2.000 108.400 ;
        RECT 1.200 107.600 2.800 108.200 ;
        RECT 4.200 107.600 6.800 108.400 ;
        RECT 9.200 107.600 10.000 109.200 ;
        RECT 2.000 107.200 2.800 107.600 ;
        RECT 1.400 106.200 5.000 106.600 ;
        RECT 6.000 106.400 6.600 107.600 ;
        RECT 1.200 106.000 5.200 106.200 ;
        RECT 1.200 102.200 2.000 106.000 ;
        RECT 4.400 102.200 5.200 106.000 ;
        RECT 6.000 102.200 6.800 106.400 ;
        RECT 11.000 106.200 11.600 109.600 ;
        RECT 12.200 108.800 13.000 109.600 ;
        RECT 12.400 108.400 13.000 108.800 ;
        RECT 12.400 107.600 13.200 108.400 ;
        RECT 10.600 104.400 12.200 106.200 ;
        RECT 15.600 105.600 16.400 106.400 ;
        RECT 17.400 106.200 18.000 109.800 ;
        RECT 20.400 109.700 22.800 109.800 ;
        RECT 20.400 109.600 21.200 109.700 ;
        RECT 22.000 109.600 22.800 109.700 ;
        RECT 24.000 109.800 24.800 110.000 ;
        RECT 27.800 109.800 32.400 110.300 ;
        RECT 24.000 109.200 26.600 109.800 ;
        RECT 18.800 107.600 19.600 109.200 ;
        RECT 26.000 108.600 26.600 109.200 ;
        RECT 27.400 109.700 32.400 109.800 ;
        RECT 27.400 109.600 29.200 109.700 ;
        RECT 31.600 109.600 32.400 109.700 ;
        RECT 27.400 109.200 28.400 109.600 ;
        RECT 22.000 108.200 23.600 108.400 ;
        RECT 22.000 107.600 25.400 108.200 ;
        RECT 26.000 107.800 26.800 108.600 ;
        RECT 24.800 107.200 25.400 107.600 ;
        RECT 23.400 106.800 24.200 107.000 ;
        RECT 15.800 104.800 16.600 105.600 ;
        RECT 10.600 103.600 13.200 104.400 ;
        RECT 10.600 102.200 12.200 103.600 ;
        RECT 17.200 102.200 18.000 106.200 ;
        RECT 22.000 106.200 24.200 106.800 ;
        RECT 24.800 106.600 26.800 107.200 ;
        RECT 25.200 106.400 26.800 106.600 ;
        RECT 22.000 102.200 22.800 106.200 ;
        RECT 27.400 105.800 28.000 109.200 ;
        RECT 35.000 108.400 35.600 111.800 ;
        RECT 36.400 109.600 37.200 111.200 ;
        RECT 39.600 110.300 40.400 119.800 ;
        RECT 43.800 112.400 44.600 119.800 ;
        RECT 45.200 113.600 46.000 114.400 ;
        RECT 45.400 112.400 46.000 113.600 ;
        RECT 50.200 112.600 51.000 119.800 ;
        RECT 43.800 111.800 44.800 112.400 ;
        RECT 45.400 111.800 46.800 112.400 ;
        RECT 49.200 111.800 51.000 112.600 ;
        RECT 52.400 112.300 53.200 119.800 ;
        RECT 56.400 113.600 57.200 114.400 ;
        RECT 56.400 112.400 57.000 113.600 ;
        RECT 57.800 112.400 58.600 119.800 ;
        RECT 55.600 112.300 57.000 112.400 ;
        RECT 52.400 111.800 57.000 112.300 ;
        RECT 57.600 111.800 58.600 112.400 ;
        RECT 44.200 110.400 44.800 111.800 ;
        RECT 46.000 111.600 46.800 111.800 ;
        RECT 42.800 110.300 43.600 110.400 ;
        RECT 39.600 109.700 43.600 110.300 ;
        RECT 28.800 107.600 29.600 108.400 ;
        RECT 30.800 108.300 32.400 108.400 ;
        RECT 33.200 108.300 34.000 108.400 ;
        RECT 30.800 107.700 34.000 108.300 ;
        RECT 30.800 107.600 32.400 107.700 ;
        RECT 33.200 107.600 34.000 107.700 ;
        RECT 34.800 107.600 35.600 108.400 ;
        RECT 28.800 107.200 29.400 107.600 ;
        RECT 28.600 106.400 29.400 107.200 ;
        RECT 30.000 106.800 30.800 107.000 ;
        RECT 30.000 106.200 32.400 106.800 ;
        RECT 35.000 106.400 35.600 107.600 ;
        RECT 38.000 106.800 38.800 108.400 ;
        RECT 26.400 102.200 28.000 105.800 ;
        RECT 31.600 102.200 32.400 106.200 ;
        RECT 33.200 104.800 34.000 106.400 ;
        RECT 34.800 105.600 35.600 106.400 ;
        RECT 35.000 104.200 35.600 105.600 ;
        RECT 34.800 102.200 35.600 104.200 ;
        RECT 39.600 102.200 40.400 109.700 ;
        RECT 42.800 108.800 43.600 109.700 ;
        RECT 44.200 109.600 45.200 110.400 ;
        RECT 44.200 108.400 44.800 109.600 ;
        RECT 49.400 108.400 50.000 111.800 ;
        RECT 52.400 111.700 56.400 111.800 ;
        RECT 50.800 109.600 51.600 111.200 ;
        RECT 41.200 108.200 42.000 108.400 ;
        RECT 41.200 107.600 42.800 108.200 ;
        RECT 44.200 107.600 46.800 108.400 ;
        RECT 49.200 107.600 50.000 108.400 ;
        RECT 42.000 107.200 42.800 107.600 ;
        RECT 41.400 106.200 45.000 106.600 ;
        RECT 46.000 106.200 46.600 107.600 ;
        RECT 41.200 106.000 45.200 106.200 ;
        RECT 41.200 102.200 42.000 106.000 ;
        RECT 44.400 102.200 45.200 106.000 ;
        RECT 46.000 102.200 46.800 106.200 ;
        RECT 47.600 104.800 48.400 106.400 ;
        RECT 49.400 104.400 50.000 107.600 ;
        RECT 49.200 102.200 50.000 104.400 ;
        RECT 52.400 102.200 53.200 111.700 ;
        RECT 55.600 111.600 56.400 111.700 ;
        RECT 57.600 108.400 58.200 111.800 ;
        RECT 58.800 110.300 59.600 110.400 ;
        RECT 60.400 110.300 61.200 110.400 ;
        RECT 58.800 109.700 61.200 110.300 ;
        RECT 58.800 108.800 59.600 109.700 ;
        RECT 60.400 109.600 61.200 109.700 ;
        RECT 55.600 107.600 58.200 108.400 ;
        RECT 60.400 108.300 61.200 108.400 ;
        RECT 63.600 108.300 64.400 119.800 ;
        RECT 65.200 111.800 66.000 119.800 ;
        RECT 66.800 112.400 67.600 119.800 ;
        RECT 70.000 112.400 70.800 119.800 ;
        RECT 66.800 111.800 70.800 112.400 ;
        RECT 71.600 112.400 72.400 119.800 ;
        RECT 76.000 114.400 77.600 119.800 ;
        RECT 76.000 113.600 78.800 114.400 ;
        RECT 73.200 112.400 74.000 112.600 ;
        RECT 76.000 112.400 77.600 113.600 ;
        RECT 71.600 111.800 74.000 112.400 ;
        RECT 75.600 111.800 77.600 112.400 ;
        RECT 79.800 112.400 80.600 112.600 ;
        RECT 81.200 112.400 82.000 119.800 ;
        RECT 84.400 115.800 85.200 119.800 ;
        RECT 79.800 111.800 82.000 112.400 ;
        RECT 65.400 110.400 66.000 111.800 ;
        RECT 69.200 110.400 70.000 110.800 ;
        RECT 75.600 110.400 76.200 111.800 ;
        RECT 79.800 111.200 80.400 111.800 ;
        RECT 77.000 110.600 80.400 111.200 ;
        RECT 84.600 111.600 85.200 115.800 ;
        RECT 87.600 111.800 88.400 119.800 ;
        RECT 84.600 111.000 87.000 111.600 ;
        RECT 77.000 110.400 77.800 110.600 ;
        RECT 65.200 109.800 67.600 110.400 ;
        RECT 69.200 109.800 70.800 110.400 ;
        RECT 65.200 109.600 66.000 109.800 ;
        RECT 65.200 108.300 66.000 108.400 ;
        RECT 60.400 108.200 62.700 108.300 ;
        RECT 59.600 107.700 62.700 108.200 ;
        RECT 59.600 107.600 61.200 107.700 ;
        RECT 54.000 104.800 54.800 106.400 ;
        RECT 55.800 106.200 56.400 107.600 ;
        RECT 59.600 107.200 60.400 107.600 ;
        RECT 57.400 106.200 61.000 106.600 ;
        RECT 62.100 106.400 62.700 107.700 ;
        RECT 63.600 107.700 66.000 108.300 ;
        RECT 55.600 102.200 56.400 106.200 ;
        RECT 57.200 106.000 61.200 106.200 ;
        RECT 57.200 102.200 58.000 106.000 ;
        RECT 60.400 102.200 61.200 106.000 ;
        RECT 62.000 104.800 62.800 106.400 ;
        RECT 63.600 102.200 64.400 107.700 ;
        RECT 65.200 107.600 66.000 107.700 ;
        RECT 65.200 105.600 66.000 106.400 ;
        RECT 67.000 106.200 67.600 109.800 ;
        RECT 70.000 109.600 70.800 109.800 ;
        RECT 74.800 109.800 76.200 110.400 ;
        RECT 79.200 109.800 80.000 110.000 ;
        RECT 74.800 109.600 76.600 109.800 ;
        RECT 75.600 109.200 76.600 109.600 ;
        RECT 68.400 108.300 69.200 109.200 ;
        RECT 71.600 108.300 73.200 108.400 ;
        RECT 68.400 107.700 73.200 108.300 ;
        RECT 68.400 107.600 69.200 107.700 ;
        RECT 71.600 107.600 73.200 107.700 ;
        RECT 74.400 107.600 75.200 108.400 ;
        RECT 74.600 107.200 75.200 107.600 ;
        RECT 73.200 106.800 74.000 107.000 ;
        RECT 65.400 104.800 66.200 105.600 ;
        RECT 66.800 102.200 67.600 106.200 ;
        RECT 71.600 106.200 74.000 106.800 ;
        RECT 74.600 106.400 75.400 107.200 ;
        RECT 71.600 102.200 72.400 106.200 ;
        RECT 76.000 105.800 76.600 109.200 ;
        RECT 77.400 109.200 80.000 109.800 ;
        RECT 84.400 109.600 85.200 110.400 ;
        RECT 77.400 108.600 78.000 109.200 ;
        RECT 77.200 107.800 78.000 108.600 ;
        RECT 80.400 108.200 82.000 108.400 ;
        RECT 78.600 107.600 82.000 108.200 ;
        RECT 82.800 107.600 83.600 109.200 ;
        RECT 84.600 108.800 85.200 109.600 ;
        RECT 84.600 108.200 85.600 108.800 ;
        RECT 84.800 108.000 85.600 108.200 ;
        RECT 86.400 107.600 87.000 111.000 ;
        RECT 87.800 110.400 88.400 111.800 ;
        RECT 87.600 110.300 88.400 110.400 ;
        RECT 89.200 110.300 90.000 110.400 ;
        RECT 87.600 109.700 90.000 110.300 ;
        RECT 87.600 109.600 88.400 109.700 ;
        RECT 89.200 109.600 90.000 109.700 ;
        RECT 78.600 107.200 79.200 107.600 ;
        RECT 86.400 107.400 87.200 107.600 ;
        RECT 77.200 106.600 79.200 107.200 ;
        RECT 84.200 107.000 87.200 107.400 ;
        RECT 79.800 106.800 80.600 107.000 ;
        RECT 83.000 106.800 87.200 107.000 ;
        RECT 77.200 106.400 78.800 106.600 ;
        RECT 79.800 106.200 82.000 106.800 ;
        RECT 83.000 106.400 84.800 106.800 ;
        RECT 83.000 106.200 83.600 106.400 ;
        RECT 87.800 106.200 88.400 109.600 ;
        RECT 89.200 106.800 90.000 108.400 ;
        RECT 76.000 102.200 77.600 105.800 ;
        RECT 81.200 102.200 82.000 106.200 ;
        RECT 82.800 102.200 83.600 106.200 ;
        RECT 87.000 105.200 88.400 106.200 ;
        RECT 90.800 106.200 91.600 119.800 ;
        RECT 92.400 111.600 93.200 113.200 ;
        RECT 96.600 112.600 97.400 119.800 ;
        RECT 95.600 111.800 97.400 112.600 ;
        RECT 99.400 112.600 100.200 119.800 ;
        RECT 99.400 111.800 101.200 112.600 ;
        RECT 106.200 112.400 107.000 119.800 ;
        RECT 107.600 113.600 108.400 114.400 ;
        RECT 107.800 112.400 108.400 113.600 ;
        RECT 112.600 112.400 113.400 119.800 ;
        RECT 119.000 118.400 119.800 119.800 ;
        RECT 118.000 117.600 119.800 118.400 ;
        RECT 114.000 113.600 114.800 114.400 ;
        RECT 114.200 112.400 114.800 113.600 ;
        RECT 119.000 112.400 119.800 117.600 ;
        RECT 120.400 113.600 121.200 114.400 ;
        RECT 120.600 112.400 121.200 113.600 ;
        RECT 125.400 112.600 126.200 119.800 ;
        RECT 106.200 111.800 107.200 112.400 ;
        RECT 107.800 111.800 109.200 112.400 ;
        RECT 112.600 111.800 113.600 112.400 ;
        RECT 114.200 111.800 115.600 112.400 ;
        RECT 119.000 111.800 120.000 112.400 ;
        RECT 120.600 111.800 122.000 112.400 ;
        RECT 124.400 111.800 126.200 112.600 ;
        RECT 95.800 108.400 96.400 111.800 ;
        RECT 97.200 109.600 98.000 111.200 ;
        RECT 98.800 109.600 99.600 111.200 ;
        RECT 95.600 107.600 96.400 108.400 ;
        RECT 90.800 105.600 92.600 106.200 ;
        RECT 87.000 102.200 87.800 105.200 ;
        RECT 91.800 104.400 92.600 105.600 ;
        RECT 94.000 104.800 94.800 106.400 ;
        RECT 95.800 106.300 96.400 107.600 ;
        RECT 100.400 108.400 101.000 111.800 ;
        RECT 105.200 108.800 106.000 110.400 ;
        RECT 106.600 108.400 107.200 111.800 ;
        RECT 108.400 111.600 109.200 111.800 ;
        RECT 111.600 108.800 112.400 110.400 ;
        RECT 113.000 108.400 113.600 111.800 ;
        RECT 114.800 111.600 115.600 111.800 ;
        RECT 116.400 110.300 117.200 110.400 ;
        RECT 118.000 110.300 118.800 110.400 ;
        RECT 116.400 109.700 118.800 110.300 ;
        RECT 116.400 109.600 117.200 109.700 ;
        RECT 118.000 108.800 118.800 109.700 ;
        RECT 119.400 108.400 120.000 111.800 ;
        RECT 121.200 111.600 122.000 111.800 ;
        RECT 124.600 108.400 125.200 111.800 ;
        RECT 126.000 110.300 126.800 111.200 ;
        RECT 127.600 110.300 128.400 110.400 ;
        RECT 126.000 109.700 128.400 110.300 ;
        RECT 126.000 109.600 126.800 109.700 ;
        RECT 127.600 109.600 128.400 109.700 ;
        RECT 100.400 107.600 101.200 108.400 ;
        RECT 103.600 108.200 104.400 108.400 ;
        RECT 103.600 107.600 105.200 108.200 ;
        RECT 106.600 107.600 109.200 108.400 ;
        RECT 110.000 108.200 110.800 108.400 ;
        RECT 113.000 108.300 115.600 108.400 ;
        RECT 116.400 108.300 117.200 108.400 ;
        RECT 113.000 108.200 117.200 108.300 ;
        RECT 110.000 107.600 111.600 108.200 ;
        RECT 113.000 107.700 118.000 108.200 ;
        RECT 113.000 107.600 115.600 107.700 ;
        RECT 116.400 107.600 118.000 107.700 ;
        RECT 119.400 107.600 122.000 108.400 ;
        RECT 124.400 107.600 125.200 108.400 ;
        RECT 98.800 106.300 99.600 106.400 ;
        RECT 95.700 105.700 99.600 106.300 ;
        RECT 90.800 103.600 92.600 104.400 ;
        RECT 95.800 104.200 96.400 105.700 ;
        RECT 98.800 105.600 99.600 105.700 ;
        RECT 91.800 102.200 92.600 103.600 ;
        RECT 95.600 102.200 96.400 104.200 ;
        RECT 100.400 104.400 101.000 107.600 ;
        RECT 104.400 107.200 105.200 107.600 ;
        RECT 102.000 104.800 102.800 106.400 ;
        RECT 103.800 106.200 107.400 106.600 ;
        RECT 108.400 106.200 109.000 107.600 ;
        RECT 110.800 107.200 111.600 107.600 ;
        RECT 110.200 106.200 113.800 106.600 ;
        RECT 114.800 106.200 115.400 107.600 ;
        RECT 117.200 107.200 118.000 107.600 ;
        RECT 116.600 106.200 120.200 106.600 ;
        RECT 121.200 106.200 121.800 107.600 ;
        RECT 103.600 106.000 107.600 106.200 ;
        RECT 100.400 102.200 101.200 104.400 ;
        RECT 103.600 102.200 104.400 106.000 ;
        RECT 106.800 102.200 107.600 106.000 ;
        RECT 108.400 102.200 109.200 106.200 ;
        RECT 110.000 106.000 114.000 106.200 ;
        RECT 110.000 102.200 110.800 106.000 ;
        RECT 113.200 102.200 114.000 106.000 ;
        RECT 114.800 102.200 115.600 106.200 ;
        RECT 116.400 106.000 120.400 106.200 ;
        RECT 116.400 102.200 117.200 106.000 ;
        RECT 119.600 102.200 120.400 106.000 ;
        RECT 121.200 102.200 122.000 106.200 ;
        RECT 122.800 104.800 123.600 106.400 ;
        RECT 124.600 104.400 125.200 107.600 ;
        RECT 129.200 108.300 130.000 119.800 ;
        RECT 130.800 112.400 131.600 119.800 ;
        RECT 134.000 112.400 134.800 119.800 ;
        RECT 130.800 111.800 134.800 112.400 ;
        RECT 135.600 111.800 136.400 119.800 ;
        RECT 137.200 116.300 138.000 116.400 ;
        RECT 142.000 116.300 142.800 119.800 ;
        RECT 137.200 115.700 142.800 116.300 ;
        RECT 137.200 115.600 138.000 115.700 ;
        RECT 131.600 110.400 132.400 110.800 ;
        RECT 135.600 110.400 136.200 111.800 ;
        RECT 130.800 109.800 132.400 110.400 ;
        RECT 134.000 109.800 136.400 110.400 ;
        RECT 130.800 109.600 131.600 109.800 ;
        RECT 134.000 109.600 134.800 109.800 ;
        RECT 135.600 109.600 136.400 109.800 ;
        RECT 132.400 108.300 133.200 109.200 ;
        RECT 129.200 107.700 133.200 108.300 ;
        RECT 127.600 104.800 128.400 106.400 ;
        RECT 124.400 102.200 125.200 104.400 ;
        RECT 129.200 102.200 130.000 107.700 ;
        RECT 132.400 107.600 133.200 107.700 ;
        RECT 134.000 106.200 134.600 109.600 ;
        RECT 134.000 102.200 134.800 106.200 ;
        RECT 135.600 105.600 136.400 106.400 ;
        RECT 135.400 104.800 136.200 105.600 ;
        RECT 142.000 102.200 142.800 115.700 ;
        RECT 147.800 112.600 148.600 119.800 ;
        RECT 146.800 111.800 148.600 112.600 ;
        RECT 150.000 112.400 150.800 119.800 ;
        RECT 151.800 112.400 152.600 112.600 ;
        RECT 150.000 111.800 152.600 112.400 ;
        RECT 154.400 111.800 156.000 119.800 ;
        RECT 158.000 112.400 158.800 112.600 ;
        RECT 159.600 112.400 160.400 119.800 ;
        RECT 158.000 111.800 160.400 112.400 ;
        RECT 147.000 108.400 147.600 111.800 ;
        RECT 148.400 109.600 149.200 111.200 ;
        RECT 153.000 110.400 153.800 110.600 ;
        RECT 155.000 110.400 155.600 111.800 ;
        RECT 152.200 109.800 153.800 110.400 ;
        RECT 152.200 109.600 153.000 109.800 ;
        RECT 154.800 109.600 155.600 110.400 ;
        RECT 156.400 110.300 157.200 110.400 ;
        RECT 161.200 110.300 162.000 119.800 ;
        RECT 164.400 111.400 165.200 119.800 ;
        RECT 168.800 116.400 169.600 119.800 ;
        RECT 167.600 115.800 169.600 116.400 ;
        RECT 173.200 115.800 174.000 119.800 ;
        RECT 177.400 115.800 178.600 119.800 ;
        RECT 167.600 115.000 168.400 115.800 ;
        RECT 173.200 115.200 173.800 115.800 ;
        RECT 171.000 114.600 174.600 115.200 ;
        RECT 177.200 115.000 178.000 115.800 ;
        RECT 171.000 114.400 171.800 114.600 ;
        RECT 173.800 114.400 174.600 114.600 ;
        RECT 167.600 113.000 168.400 113.200 ;
        RECT 172.200 113.000 173.000 113.200 ;
        RECT 167.600 112.400 173.000 113.000 ;
        RECT 173.600 113.000 175.800 113.600 ;
        RECT 173.600 111.800 174.200 113.000 ;
        RECT 175.000 112.800 175.800 113.000 ;
        RECT 177.400 113.200 178.800 114.000 ;
        RECT 177.400 112.200 178.000 113.200 ;
        RECT 169.400 111.400 174.200 111.800 ;
        RECT 164.400 111.200 174.200 111.400 ;
        RECT 175.600 111.600 178.000 112.200 ;
        RECT 164.400 111.000 170.200 111.200 ;
        RECT 164.400 110.800 170.000 111.000 ;
        RECT 156.400 109.700 162.000 110.300 ;
        RECT 170.800 110.200 171.600 110.400 ;
        RECT 156.400 109.600 157.200 109.700 ;
        RECT 153.600 108.600 154.400 108.800 ;
        RECT 151.600 108.400 154.400 108.600 ;
        RECT 146.800 108.300 147.600 108.400 ;
        RECT 143.700 107.700 147.600 108.300 ;
        RECT 143.700 106.400 144.300 107.700 ;
        RECT 146.800 107.600 147.600 107.700 ;
        RECT 150.000 108.000 154.400 108.400 ;
        RECT 155.000 108.400 155.600 109.600 ;
        RECT 150.000 107.800 152.200 108.000 ;
        RECT 155.000 107.800 156.000 108.400 ;
        RECT 150.000 107.600 151.600 107.800 ;
        RECT 143.600 104.800 144.400 106.400 ;
        RECT 145.200 104.800 146.000 106.400 ;
        RECT 147.000 104.200 147.600 107.600 ;
        RECT 151.800 106.800 152.600 107.000 ;
        RECT 146.800 102.200 147.600 104.200 ;
        RECT 150.000 106.200 152.600 106.800 ;
        RECT 153.200 106.400 154.800 107.200 ;
        RECT 150.000 102.200 150.800 106.200 ;
        RECT 155.400 105.800 156.000 107.800 ;
        RECT 156.800 107.600 157.600 108.400 ;
        RECT 158.800 107.600 160.400 108.400 ;
        RECT 156.800 107.200 157.400 107.600 ;
        RECT 156.600 106.400 157.400 107.200 ;
        RECT 158.000 106.800 158.800 107.000 ;
        RECT 158.000 106.200 160.400 106.800 ;
        RECT 154.400 104.400 156.000 105.800 ;
        RECT 153.200 103.600 156.000 104.400 ;
        RECT 154.400 102.200 156.000 103.600 ;
        RECT 159.600 102.200 160.400 106.200 ;
        RECT 161.200 102.200 162.000 109.700 ;
        RECT 166.600 109.600 171.600 110.200 ;
        RECT 174.000 110.300 174.800 110.400 ;
        RECT 175.600 110.300 176.200 111.600 ;
        RECT 182.000 111.200 182.800 119.800 ;
        RECT 178.600 110.600 182.800 111.200 ;
        RECT 178.600 110.400 179.400 110.600 ;
        RECT 174.000 109.700 176.300 110.300 ;
        RECT 180.200 109.800 181.000 110.000 ;
        RECT 174.000 109.600 174.800 109.700 ;
        RECT 166.600 109.400 167.400 109.600 ;
        RECT 169.200 109.400 170.000 109.600 ;
        RECT 168.200 108.400 169.000 108.600 ;
        RECT 175.600 108.400 176.200 109.700 ;
        RECT 177.200 109.200 181.000 109.800 ;
        RECT 177.200 109.000 178.000 109.200 ;
        RECT 165.200 107.800 176.200 108.400 ;
        RECT 165.200 107.600 166.800 107.800 ;
        RECT 162.800 104.800 163.600 106.400 ;
        RECT 164.400 102.200 165.200 107.000 ;
        RECT 169.400 106.400 170.000 107.800 ;
        RECT 175.000 107.600 175.800 107.800 ;
        RECT 182.000 107.200 182.800 110.600 ;
        RECT 179.000 106.600 182.800 107.200 ;
        RECT 183.600 106.800 184.400 108.400 ;
        RECT 185.200 108.300 186.000 119.800 ;
        RECT 188.400 114.300 189.200 114.400 ;
        RECT 190.000 114.300 190.800 119.800 ;
        RECT 188.400 113.700 190.800 114.300 ;
        RECT 188.400 113.600 189.200 113.700 ;
        RECT 188.400 108.300 189.200 108.400 ;
        RECT 185.200 107.700 189.200 108.300 ;
        RECT 179.000 106.400 179.800 106.600 ;
        RECT 167.600 104.200 168.400 105.000 ;
        RECT 169.200 104.800 170.000 106.400 ;
        RECT 171.000 105.400 171.800 105.600 ;
        RECT 171.000 104.800 173.800 105.400 ;
        RECT 173.200 104.200 173.800 104.800 ;
        RECT 177.200 104.200 178.000 105.000 ;
        RECT 167.600 103.600 169.600 104.200 ;
        RECT 168.800 102.200 169.600 103.600 ;
        RECT 173.200 102.200 174.000 104.200 ;
        RECT 177.200 103.600 178.600 104.200 ;
        RECT 177.400 102.200 178.600 103.600 ;
        RECT 182.000 102.200 182.800 106.600 ;
        RECT 185.200 102.200 186.000 107.700 ;
        RECT 188.400 106.800 189.200 107.700 ;
        RECT 190.000 106.300 190.800 113.700 ;
        RECT 191.600 111.600 192.400 113.200 ;
        RECT 193.200 106.300 194.000 106.400 ;
        RECT 190.000 105.700 194.000 106.300 ;
        RECT 190.000 105.600 191.800 105.700 ;
        RECT 191.000 102.200 191.800 105.600 ;
        RECT 193.200 104.800 194.000 105.700 ;
        RECT 194.800 102.200 195.600 119.800 ;
        RECT 197.200 113.600 198.000 114.400 ;
        RECT 197.200 112.400 197.800 113.600 ;
        RECT 198.600 112.400 199.400 119.800 ;
        RECT 196.400 111.800 197.800 112.400 ;
        RECT 198.400 111.800 199.400 112.400 ;
        RECT 202.800 112.400 203.600 119.800 ;
        RECT 206.000 119.200 210.000 119.800 ;
        RECT 206.000 112.400 206.800 119.200 ;
        RECT 202.800 111.800 206.800 112.400 ;
        RECT 207.600 111.800 208.400 118.600 ;
        RECT 209.200 111.800 210.000 119.200 ;
        RECT 196.400 111.600 197.200 111.800 ;
        RECT 198.400 108.400 199.000 111.800 ;
        RECT 207.600 111.200 208.200 111.800 ;
        RECT 210.800 111.600 211.600 113.200 ;
        RECT 203.600 110.400 204.400 110.800 ;
        RECT 206.200 110.600 208.200 111.200 ;
        RECT 206.200 110.400 206.800 110.600 ;
        RECT 199.600 110.300 200.400 110.400 ;
        RECT 201.200 110.300 202.000 110.400 ;
        RECT 199.600 109.700 202.000 110.300 ;
        RECT 199.600 108.800 200.400 109.700 ;
        RECT 201.200 109.600 202.000 109.700 ;
        RECT 202.800 109.800 204.400 110.400 ;
        RECT 202.800 109.600 203.600 109.800 ;
        RECT 206.000 109.600 206.800 110.400 ;
        RECT 209.200 109.600 210.000 111.200 ;
        RECT 196.400 107.600 199.000 108.400 ;
        RECT 201.200 108.200 202.000 108.400 ;
        RECT 200.400 107.600 202.000 108.200 ;
        RECT 204.400 107.600 205.200 109.200 ;
        RECT 196.600 106.200 197.200 107.600 ;
        RECT 200.400 107.200 201.200 107.600 ;
        RECT 198.200 106.200 201.800 106.600 ;
        RECT 206.200 106.200 206.800 109.600 ;
        RECT 207.400 108.800 208.200 109.600 ;
        RECT 207.600 108.400 208.200 108.800 ;
        RECT 207.600 107.600 208.400 108.400 ;
        RECT 209.200 108.300 210.000 108.400 ;
        RECT 212.400 108.300 213.200 119.800 ;
        RECT 215.600 111.800 216.400 119.800 ;
        RECT 217.200 112.400 218.000 119.800 ;
        RECT 220.400 112.400 221.200 119.800 ;
        RECT 217.200 111.800 221.200 112.400 ;
        RECT 222.000 112.400 222.800 119.800 ;
        RECT 225.200 119.200 229.200 119.800 ;
        RECT 225.200 112.400 226.000 119.200 ;
        RECT 222.000 111.800 226.000 112.400 ;
        RECT 226.800 111.800 227.600 118.600 ;
        RECT 228.400 111.800 229.200 119.200 ;
        RECT 230.800 113.600 231.600 114.400 ;
        RECT 230.800 112.400 231.400 113.600 ;
        RECT 232.200 112.400 233.000 119.800 ;
        RECT 240.200 112.800 241.000 119.800 ;
        RECT 244.400 115.000 245.200 119.000 ;
        RECT 230.000 111.800 231.400 112.400 ;
        RECT 215.800 110.400 216.400 111.800 ;
        RECT 226.800 111.200 227.400 111.800 ;
        RECT 230.000 111.600 230.800 111.800 ;
        RECT 232.000 111.600 234.000 112.400 ;
        RECT 239.400 112.200 241.000 112.800 ;
        RECT 219.600 110.400 220.400 110.800 ;
        RECT 222.800 110.400 223.600 110.800 ;
        RECT 225.400 110.600 227.400 111.200 ;
        RECT 225.400 110.400 226.000 110.600 ;
        RECT 215.600 109.800 218.000 110.400 ;
        RECT 219.600 109.800 221.200 110.400 ;
        RECT 215.600 109.600 216.400 109.800 ;
        RECT 217.200 109.600 218.000 109.800 ;
        RECT 220.400 109.600 221.200 109.800 ;
        RECT 222.000 109.800 223.600 110.400 ;
        RECT 222.000 109.600 222.800 109.800 ;
        RECT 225.200 109.600 226.000 110.400 ;
        RECT 228.400 109.600 229.200 111.200 ;
        RECT 209.200 107.700 213.200 108.300 ;
        RECT 209.200 107.600 210.000 107.700 ;
        RECT 212.400 106.200 213.200 107.700 ;
        RECT 214.000 106.800 214.800 108.400 ;
        RECT 196.400 102.200 197.200 106.200 ;
        RECT 198.000 106.000 202.000 106.200 ;
        RECT 198.000 102.200 198.800 106.000 ;
        RECT 201.200 102.200 202.000 106.000 ;
        RECT 205.800 102.200 207.400 106.200 ;
        RECT 211.400 105.600 213.200 106.200 ;
        RECT 215.600 105.600 216.400 106.400 ;
        RECT 217.400 106.200 218.000 109.600 ;
        RECT 218.800 107.600 219.600 109.200 ;
        RECT 223.600 107.600 224.400 109.200 ;
        RECT 225.400 108.400 226.000 109.600 ;
        RECT 226.600 108.800 227.400 109.600 ;
        RECT 225.200 107.600 226.000 108.400 ;
        RECT 226.800 108.400 227.400 108.800 ;
        RECT 232.000 108.400 232.600 111.600 ;
        RECT 233.200 108.800 234.000 110.400 ;
        RECT 234.800 110.300 235.600 110.400 ;
        RECT 238.000 110.300 238.800 111.200 ;
        RECT 234.800 109.700 238.800 110.300 ;
        RECT 234.800 109.600 235.600 109.700 ;
        RECT 238.000 109.600 238.800 109.700 ;
        RECT 239.400 108.400 240.000 112.200 ;
        RECT 244.600 111.600 245.200 115.000 ;
        RECT 246.000 112.400 246.800 119.800 ;
        RECT 250.400 118.400 252.000 119.800 ;
        RECT 250.400 117.600 253.200 118.400 ;
        RECT 247.600 112.400 248.400 112.600 ;
        RECT 246.000 111.800 248.400 112.400 ;
        RECT 250.400 111.800 252.000 117.600 ;
        RECT 253.800 112.400 254.600 112.600 ;
        RECT 255.600 112.400 256.400 119.800 ;
        RECT 253.800 111.800 256.400 112.400 ;
        RECT 241.400 111.000 245.200 111.600 ;
        RECT 241.400 109.000 242.000 111.000 ;
        RECT 250.800 110.400 251.400 111.800 ;
        RECT 252.600 110.400 253.400 110.600 ;
        RECT 226.800 107.600 227.600 108.400 ;
        RECT 230.000 107.600 232.600 108.400 ;
        RECT 234.800 108.200 235.600 108.400 ;
        RECT 234.000 107.600 235.600 108.200 ;
        RECT 238.000 107.600 240.000 108.400 ;
        RECT 240.600 108.200 242.000 109.000 ;
        RECT 242.800 108.800 243.600 110.400 ;
        RECT 244.400 108.800 245.200 110.400 ;
        RECT 250.800 109.600 251.600 110.400 ;
        RECT 252.600 109.800 254.200 110.400 ;
        RECT 253.400 109.600 254.200 109.800 ;
        RECT 250.800 108.400 251.400 109.600 ;
        RECT 225.400 106.200 226.000 107.600 ;
        RECT 230.200 106.200 230.800 107.600 ;
        RECT 234.000 107.200 234.800 107.600 ;
        RECT 239.400 107.000 240.000 107.600 ;
        RECT 241.000 107.800 242.000 108.200 ;
        RECT 241.000 107.200 245.200 107.800 ;
        RECT 246.000 107.600 247.600 108.400 ;
        RECT 248.800 107.600 249.600 108.400 ;
        RECT 239.400 106.600 240.200 107.000 ;
        RECT 231.800 106.200 235.400 106.600 ;
        RECT 211.400 102.200 212.200 105.600 ;
        RECT 215.800 104.800 216.600 105.600 ;
        RECT 217.200 102.200 218.000 106.200 ;
        RECT 225.000 102.200 226.600 106.200 ;
        RECT 230.000 102.200 230.800 106.200 ;
        RECT 231.600 106.000 235.600 106.200 ;
        RECT 239.400 106.000 241.000 106.600 ;
        RECT 231.600 102.200 232.400 106.000 ;
        RECT 234.800 102.200 235.600 106.000 ;
        RECT 239.600 105.600 241.000 106.000 ;
        RECT 240.200 103.000 241.000 105.600 ;
        RECT 244.600 105.000 245.200 107.200 ;
        RECT 249.000 107.200 249.600 107.600 ;
        RECT 250.400 107.800 251.400 108.400 ;
        RECT 252.000 108.600 252.800 108.800 ;
        RECT 252.000 108.400 254.800 108.600 ;
        RECT 252.000 108.000 256.400 108.400 ;
        RECT 254.200 107.800 256.400 108.000 ;
        RECT 247.600 106.800 248.400 107.000 ;
        RECT 244.400 103.000 245.200 105.000 ;
        RECT 246.000 106.200 248.400 106.800 ;
        RECT 249.000 106.400 249.800 107.200 ;
        RECT 246.000 102.200 246.800 106.200 ;
        RECT 250.400 105.800 251.000 107.800 ;
        RECT 254.800 107.600 256.400 107.800 ;
        RECT 251.600 106.400 253.200 107.200 ;
        RECT 253.800 106.800 254.600 107.000 ;
        RECT 253.800 106.200 256.400 106.800 ;
        RECT 250.400 102.200 252.000 105.800 ;
        RECT 255.600 102.200 256.400 106.200 ;
        RECT 257.200 104.800 258.000 106.400 ;
        RECT 258.800 102.200 259.600 119.800 ;
        RECT 260.400 111.600 261.200 113.200 ;
        RECT 262.000 112.300 262.800 119.800 ;
        RECT 266.000 113.600 266.800 114.400 ;
        RECT 266.000 112.400 266.600 113.600 ;
        RECT 267.400 112.400 268.200 119.800 ;
        RECT 265.200 112.300 266.600 112.400 ;
        RECT 262.000 111.800 266.600 112.300 ;
        RECT 267.200 111.800 268.200 112.400 ;
        RECT 262.000 111.700 266.000 111.800 ;
        RECT 262.000 106.200 262.800 111.700 ;
        RECT 265.200 111.600 266.000 111.700 ;
        RECT 267.200 108.400 267.800 111.800 ;
        RECT 268.400 108.800 269.200 110.400 ;
        RECT 263.600 106.800 264.400 108.400 ;
        RECT 265.200 107.600 267.800 108.400 ;
        RECT 270.000 108.300 270.800 108.400 ;
        RECT 271.600 108.300 272.400 108.400 ;
        RECT 270.000 108.200 272.400 108.300 ;
        RECT 269.200 107.700 272.400 108.200 ;
        RECT 269.200 107.600 270.800 107.700 ;
        RECT 265.400 106.200 266.000 107.600 ;
        RECT 269.200 107.200 270.000 107.600 ;
        RECT 271.600 106.800 272.400 107.700 ;
        RECT 267.000 106.200 270.600 106.600 ;
        RECT 273.200 106.200 274.000 119.800 ;
        RECT 274.800 111.600 275.600 113.200 ;
        RECT 279.000 112.400 279.800 119.800 ;
        RECT 280.400 113.600 281.200 114.400 ;
        RECT 280.600 112.400 281.200 113.600 ;
        RECT 282.800 112.400 283.600 119.800 ;
        RECT 287.200 114.400 288.800 119.800 ;
        RECT 287.200 113.600 290.000 114.400 ;
        RECT 284.400 112.400 285.200 112.600 ;
        RECT 287.200 112.400 288.800 113.600 ;
        RECT 279.000 111.800 280.000 112.400 ;
        RECT 280.600 111.800 282.000 112.400 ;
        RECT 282.800 111.800 285.200 112.400 ;
        RECT 286.800 111.800 288.800 112.400 ;
        RECT 291.000 112.400 291.800 112.600 ;
        RECT 292.400 112.400 293.200 119.800 ;
        RECT 291.000 111.800 293.200 112.400 ;
        RECT 279.400 110.400 280.000 111.800 ;
        RECT 281.200 111.600 282.000 111.800 ;
        RECT 286.800 110.400 287.400 111.800 ;
        RECT 291.000 111.200 291.600 111.800 ;
        RECT 288.200 110.600 291.600 111.200 ;
        RECT 288.200 110.400 289.000 110.600 ;
        RECT 278.000 108.800 278.800 110.400 ;
        RECT 279.400 109.600 280.400 110.400 ;
        RECT 286.000 109.800 287.400 110.400 ;
        RECT 300.400 110.300 301.200 119.800 ;
        RECT 303.600 112.400 304.400 119.800 ;
        RECT 303.600 111.800 305.800 112.400 ;
        RECT 306.800 111.800 307.600 119.800 ;
        RECT 305.200 111.200 305.800 111.800 ;
        RECT 305.200 110.400 306.400 111.200 ;
        RECT 303.600 110.300 304.400 110.400 ;
        RECT 290.400 109.800 291.200 110.000 ;
        RECT 286.000 109.600 287.800 109.800 ;
        RECT 279.400 108.400 280.000 109.600 ;
        RECT 286.800 109.200 287.800 109.600 ;
        RECT 276.400 108.200 277.200 108.400 ;
        RECT 276.400 107.600 278.000 108.200 ;
        RECT 279.400 107.600 282.000 108.400 ;
        RECT 282.800 107.600 284.400 108.400 ;
        RECT 285.600 107.600 286.400 108.400 ;
        RECT 277.200 107.200 278.000 107.600 ;
        RECT 276.600 106.200 280.200 106.600 ;
        RECT 281.200 106.200 281.800 107.600 ;
        RECT 285.800 107.200 286.400 107.600 ;
        RECT 284.400 106.800 285.200 107.000 ;
        RECT 282.800 106.200 285.200 106.800 ;
        RECT 285.800 106.400 286.600 107.200 ;
        RECT 261.000 105.600 262.800 106.200 ;
        RECT 261.000 102.200 261.800 105.600 ;
        RECT 265.200 102.200 266.000 106.200 ;
        RECT 266.800 106.000 270.800 106.200 ;
        RECT 266.800 102.200 267.600 106.000 ;
        RECT 270.000 102.200 270.800 106.000 ;
        RECT 273.200 105.600 275.000 106.200 ;
        RECT 274.200 102.200 275.000 105.600 ;
        RECT 276.400 106.000 280.400 106.200 ;
        RECT 276.400 102.200 277.200 106.000 ;
        RECT 279.600 102.200 280.400 106.000 ;
        RECT 281.200 102.200 282.000 106.200 ;
        RECT 282.800 102.200 283.600 106.200 ;
        RECT 287.200 105.800 287.800 109.200 ;
        RECT 288.600 109.200 291.200 109.800 ;
        RECT 300.400 109.700 304.400 110.300 ;
        RECT 288.600 108.600 289.200 109.200 ;
        RECT 288.400 107.800 289.200 108.600 ;
        RECT 291.600 108.200 293.200 108.400 ;
        RECT 289.800 107.600 293.200 108.200 ;
        RECT 289.800 107.200 290.400 107.600 ;
        RECT 288.400 106.600 290.400 107.200 ;
        RECT 291.000 106.800 291.800 107.000 ;
        RECT 298.800 106.800 299.600 108.400 ;
        RECT 288.400 106.400 290.000 106.600 ;
        RECT 291.000 106.200 293.200 106.800 ;
        RECT 287.200 102.200 288.800 105.800 ;
        RECT 292.400 102.200 293.200 106.200 ;
        RECT 300.400 102.200 301.200 109.700 ;
        RECT 303.600 108.800 304.400 109.700 ;
        RECT 305.200 107.400 305.800 110.400 ;
        RECT 307.000 109.600 307.600 111.800 ;
        RECT 308.400 111.400 309.200 119.800 ;
        RECT 312.800 116.400 313.600 119.800 ;
        RECT 311.600 115.800 313.600 116.400 ;
        RECT 317.200 115.800 318.000 119.800 ;
        RECT 321.400 115.800 322.600 119.800 ;
        RECT 311.600 115.000 312.400 115.800 ;
        RECT 317.200 115.200 317.800 115.800 ;
        RECT 315.000 114.600 318.600 115.200 ;
        RECT 321.200 115.000 322.000 115.800 ;
        RECT 315.000 114.400 315.800 114.600 ;
        RECT 317.800 114.400 318.600 114.600 ;
        RECT 311.600 113.000 312.400 113.200 ;
        RECT 316.200 113.000 317.000 113.200 ;
        RECT 311.600 112.400 317.000 113.000 ;
        RECT 317.600 113.000 319.800 113.600 ;
        RECT 317.600 111.800 318.200 113.000 ;
        RECT 319.000 112.800 319.800 113.000 ;
        RECT 321.400 113.200 322.800 114.000 ;
        RECT 321.400 112.200 322.000 113.200 ;
        RECT 313.400 111.400 318.200 111.800 ;
        RECT 308.400 111.200 318.200 111.400 ;
        RECT 319.600 111.600 322.000 112.200 ;
        RECT 308.400 111.000 314.200 111.200 ;
        RECT 308.400 110.800 314.000 111.000 ;
        RECT 314.800 110.200 315.600 110.400 ;
        RECT 303.600 106.800 305.800 107.400 ;
        RECT 303.600 102.200 304.400 106.800 ;
        RECT 306.800 102.200 307.600 109.600 ;
        RECT 310.600 109.600 315.600 110.200 ;
        RECT 310.600 109.400 311.400 109.600 ;
        RECT 313.200 109.400 314.000 109.600 ;
        RECT 312.200 108.400 313.000 108.600 ;
        RECT 319.600 108.400 320.200 111.600 ;
        RECT 326.000 111.200 326.800 119.800 ;
        RECT 322.600 110.600 326.800 111.200 ;
        RECT 327.600 111.400 328.400 119.800 ;
        RECT 332.000 116.400 332.800 119.800 ;
        RECT 330.800 115.800 332.800 116.400 ;
        RECT 336.400 115.800 337.200 119.800 ;
        RECT 340.600 115.800 341.800 119.800 ;
        RECT 330.800 115.000 331.600 115.800 ;
        RECT 336.400 115.200 337.000 115.800 ;
        RECT 334.200 114.600 337.800 115.200 ;
        RECT 340.400 115.000 341.200 115.800 ;
        RECT 334.200 114.400 335.000 114.600 ;
        RECT 337.000 114.400 337.800 114.600 ;
        RECT 330.800 113.000 331.600 113.200 ;
        RECT 335.400 113.000 336.200 113.200 ;
        RECT 330.800 112.400 336.200 113.000 ;
        RECT 336.800 113.000 339.000 113.600 ;
        RECT 336.800 111.800 337.400 113.000 ;
        RECT 338.200 112.800 339.000 113.000 ;
        RECT 340.600 113.200 342.000 114.000 ;
        RECT 340.600 112.200 341.200 113.200 ;
        RECT 332.600 111.400 337.400 111.800 ;
        RECT 327.600 111.200 337.400 111.400 ;
        RECT 338.800 111.600 341.200 112.200 ;
        RECT 327.600 111.000 333.400 111.200 ;
        RECT 327.600 110.800 333.200 111.000 ;
        RECT 322.600 110.400 323.400 110.600 ;
        RECT 324.200 109.800 325.000 110.000 ;
        RECT 321.200 109.200 325.000 109.800 ;
        RECT 321.200 109.000 322.000 109.200 ;
        RECT 309.200 107.800 320.200 108.400 ;
        RECT 309.200 107.600 310.800 107.800 ;
        RECT 308.400 102.200 309.200 107.000 ;
        RECT 313.400 105.600 314.000 107.800 ;
        RECT 314.800 107.600 315.600 107.800 ;
        RECT 319.000 107.600 319.800 107.800 ;
        RECT 326.000 107.200 326.800 110.600 ;
        RECT 334.000 110.200 334.800 110.400 ;
        RECT 329.800 109.600 334.800 110.200 ;
        RECT 329.800 109.400 330.600 109.600 ;
        RECT 332.400 109.400 333.200 109.600 ;
        RECT 331.400 108.400 332.200 108.600 ;
        RECT 338.800 108.400 339.400 111.600 ;
        RECT 345.200 111.200 346.000 119.800 ;
        RECT 348.400 112.800 349.200 119.800 ;
        RECT 341.800 110.600 346.000 111.200 ;
        RECT 341.800 110.400 342.600 110.600 ;
        RECT 343.400 109.800 344.200 110.000 ;
        RECT 340.400 109.200 344.200 109.800 ;
        RECT 340.400 109.000 341.200 109.200 ;
        RECT 328.400 107.800 339.400 108.400 ;
        RECT 328.400 107.600 330.000 107.800 ;
        RECT 323.000 106.600 326.800 107.200 ;
        RECT 323.000 106.400 323.800 106.600 ;
        RECT 311.600 104.200 312.400 105.000 ;
        RECT 313.200 104.800 314.000 105.600 ;
        RECT 315.000 105.400 315.800 105.600 ;
        RECT 315.000 104.800 317.800 105.400 ;
        RECT 317.200 104.200 317.800 104.800 ;
        RECT 321.200 104.200 322.000 105.000 ;
        RECT 311.600 103.600 313.600 104.200 ;
        RECT 312.800 102.200 313.600 103.600 ;
        RECT 317.200 102.200 318.000 104.200 ;
        RECT 321.200 103.600 322.600 104.200 ;
        RECT 321.400 102.200 322.600 103.600 ;
        RECT 326.000 102.200 326.800 106.600 ;
        RECT 327.600 102.200 328.400 107.000 ;
        RECT 332.600 105.600 333.200 107.800 ;
        RECT 338.200 107.600 339.000 107.800 ;
        RECT 345.200 107.200 346.000 110.600 ;
        RECT 342.200 106.600 346.000 107.200 ;
        RECT 342.200 106.400 343.000 106.600 ;
        RECT 330.800 104.200 331.600 105.000 ;
        RECT 332.400 104.800 333.200 105.600 ;
        RECT 334.200 105.400 335.000 105.600 ;
        RECT 334.200 104.800 337.000 105.400 ;
        RECT 336.400 104.200 337.000 104.800 ;
        RECT 340.400 104.200 341.200 105.000 ;
        RECT 330.800 103.600 332.800 104.200 ;
        RECT 332.000 102.200 332.800 103.600 ;
        RECT 336.400 102.200 337.200 104.200 ;
        RECT 340.400 103.600 341.800 104.200 ;
        RECT 340.600 102.200 341.800 103.600 ;
        RECT 345.200 102.200 346.000 106.600 ;
        RECT 348.200 111.800 349.200 112.800 ;
        RECT 351.600 112.400 352.400 119.800 ;
        RECT 349.800 111.800 352.400 112.400 ;
        RECT 353.200 112.400 354.000 119.800 ;
        RECT 356.400 112.800 357.200 119.800 ;
        RECT 353.200 111.800 355.800 112.400 ;
        RECT 356.400 111.800 357.400 112.800 ;
        RECT 359.600 112.400 360.400 119.800 ;
        RECT 362.800 112.800 363.600 119.800 ;
        RECT 359.600 111.800 362.200 112.400 ;
        RECT 362.800 111.800 363.800 112.800 ;
        RECT 368.600 112.400 369.400 119.800 ;
        RECT 370.000 113.600 370.800 114.400 ;
        RECT 370.200 112.400 370.800 113.600 ;
        RECT 376.200 112.800 377.000 119.800 ;
        RECT 380.400 115.000 381.200 119.000 ;
        RECT 368.600 111.800 369.600 112.400 ;
        RECT 370.200 111.800 371.600 112.400 ;
        RECT 348.200 108.400 348.800 111.800 ;
        RECT 349.800 109.800 350.400 111.800 ;
        RECT 349.400 109.000 350.400 109.800 ;
        RECT 348.200 107.600 349.200 108.400 ;
        RECT 348.200 106.200 348.800 107.600 ;
        RECT 349.800 107.400 350.400 109.000 ;
        RECT 351.400 110.300 352.400 110.400 ;
        RECT 353.200 110.300 354.200 110.400 ;
        RECT 351.400 109.700 354.200 110.300 ;
        RECT 351.400 109.600 352.400 109.700 ;
        RECT 353.200 109.600 354.200 109.700 ;
        RECT 351.400 108.800 352.200 109.600 ;
        RECT 353.400 108.800 354.200 109.600 ;
        RECT 355.200 109.800 355.800 111.800 ;
        RECT 355.200 109.000 356.200 109.800 ;
        RECT 355.200 107.400 355.800 109.000 ;
        RECT 356.800 108.400 357.400 111.800 ;
        RECT 359.600 109.600 360.600 110.400 ;
        RECT 359.800 108.800 360.600 109.600 ;
        RECT 361.600 109.800 362.200 111.800 ;
        RECT 361.600 109.000 362.600 109.800 ;
        RECT 356.400 107.600 357.400 108.400 ;
        RECT 349.800 106.800 352.400 107.400 ;
        RECT 348.200 105.600 349.200 106.200 ;
        RECT 348.400 102.200 349.200 105.600 ;
        RECT 351.600 102.200 352.400 106.800 ;
        RECT 353.200 106.800 355.800 107.400 ;
        RECT 353.200 102.200 354.000 106.800 ;
        RECT 356.800 106.200 357.400 107.600 ;
        RECT 361.600 107.400 362.200 109.000 ;
        RECT 363.200 108.400 363.800 111.800 ;
        RECT 367.600 108.800 368.400 110.400 ;
        RECT 369.000 110.300 369.600 111.800 ;
        RECT 370.800 111.600 371.600 111.800 ;
        RECT 375.400 112.200 377.000 112.800 ;
        RECT 374.000 110.300 374.800 111.200 ;
        RECT 369.000 109.700 374.800 110.300 ;
        RECT 369.000 108.400 369.600 109.700 ;
        RECT 374.000 109.600 374.800 109.700 ;
        RECT 375.400 110.400 376.000 112.200 ;
        RECT 380.600 111.600 381.200 115.000 ;
        RECT 382.800 113.600 383.600 114.400 ;
        RECT 382.800 112.400 383.400 113.600 ;
        RECT 384.200 112.400 385.000 119.800 ;
        RECT 391.000 112.400 391.800 119.800 ;
        RECT 392.400 113.600 393.200 114.400 ;
        RECT 392.600 112.400 393.200 113.600 ;
        RECT 382.000 111.800 383.400 112.400 ;
        RECT 384.000 111.800 385.000 112.400 ;
        RECT 382.000 111.600 382.800 111.800 ;
        RECT 377.400 111.000 381.200 111.600 ;
        RECT 375.400 109.600 376.400 110.400 ;
        RECT 375.400 108.400 376.000 109.600 ;
        RECT 377.400 109.000 378.000 111.000 ;
        RECT 362.800 107.600 363.800 108.400 ;
        RECT 366.000 108.200 366.800 108.400 ;
        RECT 366.000 107.600 367.600 108.200 ;
        RECT 369.000 107.600 371.600 108.400 ;
        RECT 374.000 107.600 376.000 108.400 ;
        RECT 376.600 108.200 378.000 109.000 ;
        RECT 378.800 108.800 379.600 110.400 ;
        RECT 380.400 108.800 381.200 110.400 ;
        RECT 384.000 108.400 384.600 111.800 ;
        RECT 390.000 111.600 392.000 112.400 ;
        RECT 392.600 111.800 394.000 112.400 ;
        RECT 393.200 111.600 394.000 111.800 ;
        RECT 394.800 111.600 395.600 113.200 ;
        RECT 385.200 110.300 386.000 110.400 ;
        RECT 386.800 110.300 387.600 110.400 ;
        RECT 390.000 110.300 390.800 110.400 ;
        RECT 385.200 109.700 390.800 110.300 ;
        RECT 385.200 108.800 386.000 109.700 ;
        RECT 386.800 109.600 387.600 109.700 ;
        RECT 390.000 108.800 390.800 109.700 ;
        RECT 391.400 108.400 392.000 111.600 ;
        RECT 356.400 105.600 357.400 106.200 ;
        RECT 359.600 106.800 362.200 107.400 ;
        RECT 356.400 102.200 357.200 105.600 ;
        RECT 359.600 102.200 360.400 106.800 ;
        RECT 363.200 106.200 363.800 107.600 ;
        RECT 366.800 107.200 367.600 107.600 ;
        RECT 366.200 106.200 369.800 106.600 ;
        RECT 370.800 106.200 371.400 107.600 ;
        RECT 375.400 107.000 376.000 107.600 ;
        RECT 377.000 107.800 378.000 108.200 ;
        RECT 377.000 107.200 381.200 107.800 ;
        RECT 382.000 107.600 384.600 108.400 ;
        RECT 386.800 108.200 387.600 108.400 ;
        RECT 386.000 107.600 387.600 108.200 ;
        RECT 388.400 108.200 389.200 108.400 ;
        RECT 388.400 107.600 390.000 108.200 ;
        RECT 391.400 107.600 394.000 108.400 ;
        RECT 375.400 106.600 376.200 107.000 ;
        RECT 362.800 105.600 363.800 106.200 ;
        RECT 366.000 106.000 370.000 106.200 ;
        RECT 362.800 102.200 363.600 105.600 ;
        RECT 366.000 102.200 366.800 106.000 ;
        RECT 369.200 102.200 370.000 106.000 ;
        RECT 370.800 102.200 371.600 106.200 ;
        RECT 375.400 106.000 377.000 106.600 ;
        RECT 376.200 103.000 377.000 106.000 ;
        RECT 380.600 105.000 381.200 107.200 ;
        RECT 382.200 106.400 382.800 107.600 ;
        RECT 386.000 107.200 386.800 107.600 ;
        RECT 389.200 107.200 390.000 107.600 ;
        RECT 380.400 103.000 381.200 105.000 ;
        RECT 382.000 102.200 382.800 106.400 ;
        RECT 383.800 106.200 387.400 106.600 ;
        RECT 388.600 106.200 392.200 106.600 ;
        RECT 393.200 106.200 393.800 107.600 ;
        RECT 396.400 106.200 397.200 119.800 ;
        RECT 402.200 112.600 403.000 119.800 ;
        RECT 401.200 111.800 403.000 112.600 ;
        RECT 401.400 108.400 402.000 111.800 ;
        RECT 402.800 110.300 403.600 111.200 ;
        RECT 404.400 110.300 405.200 119.800 ;
        RECT 410.200 112.400 411.000 119.800 ;
        RECT 416.200 118.400 417.000 119.800 ;
        RECT 416.200 117.600 418.000 118.400 ;
        RECT 411.600 113.600 412.400 114.400 ;
        RECT 411.800 112.400 412.400 113.600 ;
        RECT 414.800 113.600 415.600 114.400 ;
        RECT 414.800 112.400 415.400 113.600 ;
        RECT 416.200 112.400 417.000 117.600 ;
        RECT 410.200 111.800 411.200 112.400 ;
        RECT 411.800 111.800 413.200 112.400 ;
        RECT 402.800 109.700 405.200 110.300 ;
        RECT 402.800 109.600 403.600 109.700 ;
        RECT 398.000 106.800 398.800 108.400 ;
        RECT 401.200 107.600 402.000 108.400 ;
        RECT 383.600 106.000 387.600 106.200 ;
        RECT 383.600 102.200 384.400 106.000 ;
        RECT 386.800 102.200 387.600 106.000 ;
        RECT 388.400 106.000 392.400 106.200 ;
        RECT 388.400 102.200 389.200 106.000 ;
        RECT 391.600 102.200 392.400 106.000 ;
        RECT 393.200 102.200 394.000 106.200 ;
        RECT 395.400 105.600 397.200 106.200 ;
        RECT 395.400 104.400 396.200 105.600 ;
        RECT 399.600 104.800 400.400 106.400 ;
        RECT 401.400 104.400 402.000 107.600 ;
        RECT 394.800 103.600 396.200 104.400 ;
        RECT 395.400 102.200 396.200 103.600 ;
        RECT 401.200 102.200 402.000 104.400 ;
        RECT 404.400 108.300 405.200 109.700 ;
        RECT 406.000 110.300 406.800 110.400 ;
        RECT 409.200 110.300 410.000 110.400 ;
        RECT 406.000 109.700 410.000 110.300 ;
        RECT 406.000 109.600 406.800 109.700 ;
        RECT 409.200 108.800 410.000 109.700 ;
        RECT 410.600 110.300 411.200 111.800 ;
        RECT 412.400 111.600 413.200 111.800 ;
        RECT 414.000 111.800 415.400 112.400 ;
        RECT 416.000 111.800 417.000 112.400 ;
        RECT 420.400 112.400 421.200 119.800 ;
        RECT 422.000 112.400 422.800 112.600 ;
        RECT 424.800 112.400 426.400 119.800 ;
        RECT 420.400 111.800 422.800 112.400 ;
        RECT 424.400 111.800 426.400 112.400 ;
        RECT 428.600 112.400 429.400 112.600 ;
        RECT 430.000 112.400 430.800 119.800 ;
        RECT 428.600 111.800 430.800 112.400 ;
        RECT 414.000 111.600 414.800 111.800 ;
        RECT 412.400 110.300 413.200 110.400 ;
        RECT 410.600 109.700 413.200 110.300 ;
        RECT 410.600 108.400 411.200 109.700 ;
        RECT 412.400 109.600 413.200 109.700 ;
        RECT 416.000 108.400 416.600 111.800 ;
        RECT 424.400 110.400 425.000 111.800 ;
        RECT 428.600 111.200 429.200 111.800 ;
        RECT 425.800 110.600 429.200 111.200 ;
        RECT 431.600 111.400 432.400 119.800 ;
        RECT 436.000 116.400 436.800 119.800 ;
        RECT 434.800 115.800 436.800 116.400 ;
        RECT 440.400 115.800 441.200 119.800 ;
        RECT 444.600 115.800 445.800 119.800 ;
        RECT 434.800 115.000 435.600 115.800 ;
        RECT 440.400 115.200 441.000 115.800 ;
        RECT 438.200 114.600 441.800 115.200 ;
        RECT 444.400 115.000 445.200 115.800 ;
        RECT 438.200 114.400 439.000 114.600 ;
        RECT 441.000 114.400 441.800 114.600 ;
        RECT 434.800 113.000 435.600 113.200 ;
        RECT 439.400 113.000 440.200 113.200 ;
        RECT 434.800 112.400 440.200 113.000 ;
        RECT 440.800 113.000 443.000 113.600 ;
        RECT 440.800 111.800 441.400 113.000 ;
        RECT 442.200 112.800 443.000 113.000 ;
        RECT 444.600 113.200 446.000 114.000 ;
        RECT 444.600 112.200 445.200 113.200 ;
        RECT 436.600 111.400 441.400 111.800 ;
        RECT 431.600 111.200 441.400 111.400 ;
        RECT 442.800 111.600 445.200 112.200 ;
        RECT 431.600 111.000 437.400 111.200 ;
        RECT 431.600 110.800 437.200 111.000 ;
        RECT 425.800 110.400 426.600 110.600 ;
        RECT 417.200 108.800 418.000 110.400 ;
        RECT 423.600 109.800 425.000 110.400 ;
        RECT 438.000 110.200 438.800 110.400 ;
        RECT 428.000 109.800 428.800 110.000 ;
        RECT 423.600 109.600 425.400 109.800 ;
        RECT 424.400 109.200 425.400 109.600 ;
        RECT 407.600 108.300 408.400 108.400 ;
        RECT 404.400 108.200 408.400 108.300 ;
        RECT 404.400 107.700 409.200 108.200 ;
        RECT 404.400 102.200 405.200 107.700 ;
        RECT 407.600 107.600 409.200 107.700 ;
        RECT 410.600 107.600 413.200 108.400 ;
        RECT 414.000 107.600 416.600 108.400 ;
        RECT 418.800 108.200 419.600 108.400 ;
        RECT 418.000 107.600 419.600 108.200 ;
        RECT 420.400 107.600 422.000 108.400 ;
        RECT 423.200 107.600 424.000 108.400 ;
        RECT 408.400 107.200 409.200 107.600 ;
        RECT 406.000 104.800 406.800 106.400 ;
        RECT 407.800 106.200 411.400 106.600 ;
        RECT 412.400 106.200 413.000 107.600 ;
        RECT 414.200 106.200 414.800 107.600 ;
        RECT 418.000 107.200 418.800 107.600 ;
        RECT 423.400 107.200 424.000 107.600 ;
        RECT 422.000 106.800 422.800 107.000 ;
        RECT 415.800 106.200 419.400 106.600 ;
        RECT 420.400 106.200 422.800 106.800 ;
        RECT 423.400 106.400 424.200 107.200 ;
        RECT 407.600 106.000 411.600 106.200 ;
        RECT 407.600 102.200 408.400 106.000 ;
        RECT 410.800 102.200 411.600 106.000 ;
        RECT 412.400 102.200 413.200 106.200 ;
        RECT 414.000 102.200 414.800 106.200 ;
        RECT 415.600 106.000 419.600 106.200 ;
        RECT 415.600 102.200 416.400 106.000 ;
        RECT 418.800 102.200 419.600 106.000 ;
        RECT 420.400 102.200 421.200 106.200 ;
        RECT 424.800 105.800 425.400 109.200 ;
        RECT 426.200 109.200 428.800 109.800 ;
        RECT 433.800 109.600 438.800 110.200 ;
        RECT 433.800 109.400 434.600 109.600 ;
        RECT 436.400 109.400 437.200 109.600 ;
        RECT 426.200 108.600 426.800 109.200 ;
        RECT 426.000 107.800 426.800 108.600 ;
        RECT 435.400 108.400 436.200 108.600 ;
        RECT 442.800 108.400 443.400 111.600 ;
        RECT 449.200 111.200 450.000 119.800 ;
        RECT 445.800 110.600 450.000 111.200 ;
        RECT 445.800 110.400 446.600 110.600 ;
        RECT 447.400 109.800 448.200 110.000 ;
        RECT 444.400 109.200 448.200 109.800 ;
        RECT 444.400 109.000 445.200 109.200 ;
        RECT 429.200 108.200 430.800 108.400 ;
        RECT 427.400 107.600 430.800 108.200 ;
        RECT 432.400 107.800 443.400 108.400 ;
        RECT 432.400 107.600 434.000 107.800 ;
        RECT 427.400 107.200 428.000 107.600 ;
        RECT 426.000 106.600 428.000 107.200 ;
        RECT 428.600 106.800 429.400 107.000 ;
        RECT 426.000 106.400 427.600 106.600 ;
        RECT 428.600 106.200 430.800 106.800 ;
        RECT 424.800 102.200 426.400 105.800 ;
        RECT 430.000 102.200 430.800 106.200 ;
        RECT 431.600 102.200 432.400 107.000 ;
        RECT 436.600 105.600 437.200 107.800 ;
        RECT 442.200 107.600 443.000 107.800 ;
        RECT 449.200 107.200 450.000 110.600 ;
        RECT 446.200 106.600 450.000 107.200 ;
        RECT 446.200 106.400 447.000 106.600 ;
        RECT 434.800 104.200 435.600 105.000 ;
        RECT 436.400 104.800 437.200 105.600 ;
        RECT 438.200 105.400 439.000 105.600 ;
        RECT 438.200 104.800 441.000 105.400 ;
        RECT 440.400 104.200 441.000 104.800 ;
        RECT 444.400 104.200 445.200 105.000 ;
        RECT 434.800 103.600 436.800 104.200 ;
        RECT 436.000 102.200 436.800 103.600 ;
        RECT 440.400 102.200 441.200 104.200 ;
        RECT 444.400 103.600 445.800 104.200 ;
        RECT 444.600 102.200 445.800 103.600 ;
        RECT 449.200 102.200 450.000 106.600 ;
        RECT 457.200 102.200 458.000 119.800 ;
        RECT 458.800 110.300 459.600 110.400 ;
        RECT 460.400 110.300 461.200 119.800 ;
        RECT 458.800 109.700 461.200 110.300 ;
        RECT 458.800 109.600 459.600 109.700 ;
        RECT 458.800 106.800 459.600 108.400 ;
        RECT 460.400 102.200 461.200 109.700 ;
        RECT 463.600 111.800 464.400 119.800 ;
        RECT 466.800 112.400 467.600 119.800 ;
        RECT 465.400 111.800 467.600 112.400 ;
        RECT 468.400 112.400 469.200 119.800 ;
        RECT 470.000 112.400 470.800 112.600 ;
        RECT 468.400 111.800 470.800 112.400 ;
        RECT 472.800 111.800 474.400 119.800 ;
        RECT 476.200 112.400 477.000 112.600 ;
        RECT 478.000 112.400 478.800 119.800 ;
        RECT 476.200 111.800 478.800 112.400 ;
        RECT 463.600 109.600 464.200 111.800 ;
        RECT 465.400 111.200 466.000 111.800 ;
        RECT 464.800 110.400 466.000 111.200 ;
        RECT 473.200 110.400 473.800 111.800 ;
        RECT 475.000 110.400 475.800 110.600 ;
        RECT 462.000 106.800 462.800 108.400 ;
        RECT 463.600 102.200 464.400 109.600 ;
        RECT 465.400 107.400 466.000 110.400 ;
        RECT 466.800 108.800 467.600 110.400 ;
        RECT 473.200 109.600 474.000 110.400 ;
        RECT 475.000 109.800 476.600 110.400 ;
        RECT 475.800 109.600 476.600 109.800 ;
        RECT 473.200 108.400 473.800 109.600 ;
        RECT 468.400 107.600 470.000 108.400 ;
        RECT 471.200 107.600 472.000 108.400 ;
        RECT 465.400 106.800 467.600 107.400 ;
        RECT 471.400 107.200 472.000 107.600 ;
        RECT 472.800 107.800 473.800 108.400 ;
        RECT 474.400 108.600 475.200 108.800 ;
        RECT 474.400 108.400 477.200 108.600 ;
        RECT 474.400 108.000 478.800 108.400 ;
        RECT 476.600 107.800 478.800 108.000 ;
        RECT 470.000 106.800 470.800 107.000 ;
        RECT 466.800 102.200 467.600 106.800 ;
        RECT 468.400 106.200 470.800 106.800 ;
        RECT 471.400 106.400 472.200 107.200 ;
        RECT 468.400 102.200 469.200 106.200 ;
        RECT 472.800 105.800 473.400 107.800 ;
        RECT 477.200 107.600 478.800 107.800 ;
        RECT 474.000 106.400 475.600 107.200 ;
        RECT 476.200 106.800 477.000 107.000 ;
        RECT 479.600 106.800 480.400 108.400 ;
        RECT 476.200 106.200 478.800 106.800 ;
        RECT 472.800 102.200 474.400 105.800 ;
        RECT 478.000 102.200 478.800 106.200 ;
        RECT 481.200 102.200 482.000 119.800 ;
        RECT 484.400 111.400 485.200 119.800 ;
        RECT 488.800 116.400 489.600 119.800 ;
        RECT 487.600 115.800 489.600 116.400 ;
        RECT 493.200 115.800 494.000 119.800 ;
        RECT 497.400 115.800 498.600 119.800 ;
        RECT 487.600 115.000 488.400 115.800 ;
        RECT 493.200 115.200 493.800 115.800 ;
        RECT 491.000 114.600 494.600 115.200 ;
        RECT 497.200 115.000 498.000 115.800 ;
        RECT 491.000 114.400 491.800 114.600 ;
        RECT 493.800 114.400 494.600 114.600 ;
        RECT 487.600 113.000 488.400 113.200 ;
        RECT 492.200 113.000 493.000 113.200 ;
        RECT 487.600 112.400 493.000 113.000 ;
        RECT 493.600 113.000 495.800 113.600 ;
        RECT 493.600 111.800 494.200 113.000 ;
        RECT 495.000 112.800 495.800 113.000 ;
        RECT 497.400 113.200 498.800 114.000 ;
        RECT 497.400 112.200 498.000 113.200 ;
        RECT 489.400 111.400 494.200 111.800 ;
        RECT 484.400 111.200 494.200 111.400 ;
        RECT 495.600 111.600 498.000 112.200 ;
        RECT 484.400 111.000 490.200 111.200 ;
        RECT 484.400 110.800 490.000 111.000 ;
        RECT 495.600 110.400 496.200 111.600 ;
        RECT 502.000 111.200 502.800 119.800 ;
        RECT 498.600 110.600 502.800 111.200 ;
        RECT 503.600 111.400 504.400 119.800 ;
        RECT 508.000 116.400 508.800 119.800 ;
        RECT 506.800 115.800 508.800 116.400 ;
        RECT 512.400 115.800 513.200 119.800 ;
        RECT 516.600 115.800 517.800 119.800 ;
        RECT 506.800 115.000 507.600 115.800 ;
        RECT 512.400 115.200 513.000 115.800 ;
        RECT 510.200 114.600 513.800 115.200 ;
        RECT 516.400 115.000 517.200 115.800 ;
        RECT 510.200 114.400 511.000 114.600 ;
        RECT 513.000 114.400 513.800 114.600 ;
        RECT 517.400 114.000 518.800 114.400 ;
        RECT 516.600 113.600 518.800 114.000 ;
        RECT 506.800 113.000 507.600 113.200 ;
        RECT 511.400 113.000 512.200 113.200 ;
        RECT 506.800 112.400 512.200 113.000 ;
        RECT 512.800 113.000 515.000 113.600 ;
        RECT 512.800 111.800 513.400 113.000 ;
        RECT 514.200 112.800 515.000 113.000 ;
        RECT 516.600 113.200 518.000 113.600 ;
        RECT 516.600 112.200 517.200 113.200 ;
        RECT 508.600 111.400 513.400 111.800 ;
        RECT 503.600 111.200 513.400 111.400 ;
        RECT 514.800 111.600 517.200 112.200 ;
        RECT 503.600 111.000 509.400 111.200 ;
        RECT 503.600 110.800 509.200 111.000 ;
        RECT 498.600 110.400 499.400 110.600 ;
        RECT 490.800 110.200 491.600 110.400 ;
        RECT 486.600 109.600 491.600 110.200 ;
        RECT 495.600 109.600 496.400 110.400 ;
        RECT 500.200 109.800 501.000 110.000 ;
        RECT 486.600 109.400 487.400 109.600 ;
        RECT 489.200 109.400 490.000 109.600 ;
        RECT 488.200 108.400 489.000 108.600 ;
        RECT 495.600 108.400 496.200 109.600 ;
        RECT 497.200 109.200 501.000 109.800 ;
        RECT 497.200 109.000 498.000 109.200 ;
        RECT 485.200 107.800 496.200 108.400 ;
        RECT 485.200 107.600 486.800 107.800 ;
        RECT 484.400 102.200 485.200 107.000 ;
        RECT 489.400 105.600 490.000 107.800 ;
        RECT 495.000 107.600 495.800 107.800 ;
        RECT 502.000 107.200 502.800 110.600 ;
        RECT 510.000 110.200 510.800 110.400 ;
        RECT 505.800 109.600 510.800 110.200 ;
        RECT 505.800 109.400 506.600 109.600 ;
        RECT 508.400 109.400 509.200 109.600 ;
        RECT 507.400 108.400 508.200 108.600 ;
        RECT 514.800 108.400 515.400 111.600 ;
        RECT 521.200 111.200 522.000 119.800 ;
        RECT 522.800 112.400 523.600 119.800 ;
        RECT 524.200 112.400 525.000 112.600 ;
        RECT 522.800 111.800 525.000 112.400 ;
        RECT 527.200 112.400 528.800 119.800 ;
        RECT 530.800 112.400 531.600 112.600 ;
        RECT 532.400 112.400 533.200 119.800 ;
        RECT 527.200 111.800 529.200 112.400 ;
        RECT 530.800 111.800 533.200 112.400 ;
        RECT 534.000 112.400 534.800 119.800 ;
        RECT 535.400 112.400 536.200 112.600 ;
        RECT 534.000 111.800 536.200 112.400 ;
        RECT 538.400 112.400 540.000 119.800 ;
        RECT 542.000 112.400 542.800 112.600 ;
        RECT 543.600 112.400 544.400 119.800 ;
        RECT 538.400 111.800 540.400 112.400 ;
        RECT 542.000 111.800 544.400 112.400 ;
        RECT 517.800 110.600 522.000 111.200 ;
        RECT 524.400 111.200 525.000 111.800 ;
        RECT 524.400 110.600 527.800 111.200 ;
        RECT 517.800 110.400 518.600 110.600 ;
        RECT 519.400 109.800 520.200 110.000 ;
        RECT 516.400 109.200 520.200 109.800 ;
        RECT 516.400 109.000 517.200 109.200 ;
        RECT 504.400 107.800 515.400 108.400 ;
        RECT 504.400 107.600 506.000 107.800 ;
        RECT 499.000 106.600 502.800 107.200 ;
        RECT 499.000 106.400 499.800 106.600 ;
        RECT 487.600 104.200 488.400 105.000 ;
        RECT 489.200 104.800 490.000 105.600 ;
        RECT 491.000 105.400 491.800 105.600 ;
        RECT 491.000 104.800 493.800 105.400 ;
        RECT 493.200 104.200 493.800 104.800 ;
        RECT 497.200 104.200 498.000 105.000 ;
        RECT 487.600 103.600 489.600 104.200 ;
        RECT 488.800 102.200 489.600 103.600 ;
        RECT 493.200 102.200 494.000 104.200 ;
        RECT 497.200 103.600 498.600 104.200 ;
        RECT 497.400 102.200 498.600 103.600 ;
        RECT 502.000 102.200 502.800 106.600 ;
        RECT 503.600 102.200 504.400 107.000 ;
        RECT 508.600 105.600 509.200 107.800 ;
        RECT 510.000 107.600 510.800 107.800 ;
        RECT 514.200 107.600 515.000 107.800 ;
        RECT 521.200 107.200 522.000 110.600 ;
        RECT 527.000 110.400 527.800 110.600 ;
        RECT 528.600 110.400 529.200 111.800 ;
        RECT 535.600 111.200 536.200 111.800 ;
        RECT 535.600 110.600 539.000 111.200 ;
        RECT 538.200 110.400 539.000 110.600 ;
        RECT 539.800 110.400 540.400 111.800 ;
        RECT 545.200 111.400 546.000 119.800 ;
        RECT 549.600 116.400 550.400 119.800 ;
        RECT 548.400 115.800 550.400 116.400 ;
        RECT 554.000 115.800 554.800 119.800 ;
        RECT 558.200 115.800 559.400 119.800 ;
        RECT 548.400 115.000 549.200 115.800 ;
        RECT 554.000 115.200 554.600 115.800 ;
        RECT 551.800 114.600 555.400 115.200 ;
        RECT 558.000 115.000 558.800 115.800 ;
        RECT 551.800 114.400 552.600 114.600 ;
        RECT 554.600 114.400 555.400 114.600 ;
        RECT 548.400 113.000 549.200 113.200 ;
        RECT 553.000 113.000 553.800 113.200 ;
        RECT 548.400 112.400 553.800 113.000 ;
        RECT 554.400 113.000 556.600 113.600 ;
        RECT 554.400 111.800 555.000 113.000 ;
        RECT 555.800 112.800 556.600 113.000 ;
        RECT 558.200 113.200 559.600 114.000 ;
        RECT 558.200 112.200 558.800 113.200 ;
        RECT 550.200 111.400 555.000 111.800 ;
        RECT 545.200 111.200 555.000 111.400 ;
        RECT 556.400 111.600 558.800 112.200 ;
        RECT 545.200 111.000 551.000 111.200 ;
        RECT 545.200 110.800 550.800 111.000 ;
        RECT 524.800 109.800 525.600 110.000 ;
        RECT 528.600 109.800 530.000 110.400 ;
        RECT 524.800 109.200 527.400 109.800 ;
        RECT 526.800 108.600 527.400 109.200 ;
        RECT 528.200 109.600 530.000 109.800 ;
        RECT 536.000 109.800 536.800 110.000 ;
        RECT 539.800 109.800 541.200 110.400 ;
        RECT 551.600 110.200 552.400 110.400 ;
        RECT 528.200 109.200 529.200 109.600 ;
        RECT 536.000 109.200 538.600 109.800 ;
        RECT 522.800 108.200 524.400 108.400 ;
        RECT 522.800 107.600 526.200 108.200 ;
        RECT 526.800 107.800 527.600 108.600 ;
        RECT 518.200 106.600 522.000 107.200 ;
        RECT 525.600 107.200 526.200 107.600 ;
        RECT 524.200 106.800 525.000 107.000 ;
        RECT 518.200 106.400 519.000 106.600 ;
        RECT 506.800 104.200 507.600 105.000 ;
        RECT 508.400 104.800 509.200 105.600 ;
        RECT 510.200 105.400 511.000 105.600 ;
        RECT 510.200 104.800 513.000 105.400 ;
        RECT 512.400 104.200 513.000 104.800 ;
        RECT 516.400 104.200 517.200 105.000 ;
        RECT 506.800 103.600 508.800 104.200 ;
        RECT 508.000 102.200 508.800 103.600 ;
        RECT 512.400 102.200 513.200 104.200 ;
        RECT 516.400 103.600 517.800 104.200 ;
        RECT 516.600 102.200 517.800 103.600 ;
        RECT 521.200 102.200 522.000 106.600 ;
        RECT 522.800 106.200 525.000 106.800 ;
        RECT 525.600 106.600 527.600 107.200 ;
        RECT 526.000 106.400 527.600 106.600 ;
        RECT 522.800 102.200 523.600 106.200 ;
        RECT 528.200 105.800 528.800 109.200 ;
        RECT 538.000 108.600 538.600 109.200 ;
        RECT 539.400 109.600 541.200 109.800 ;
        RECT 547.400 109.600 552.400 110.200 ;
        RECT 554.800 110.300 555.600 110.400 ;
        RECT 556.400 110.300 557.000 111.600 ;
        RECT 562.800 111.200 563.600 119.800 ;
        RECT 559.400 110.600 563.600 111.200 ;
        RECT 564.400 111.400 565.200 119.800 ;
        RECT 568.800 116.400 569.600 119.800 ;
        RECT 567.600 115.800 569.600 116.400 ;
        RECT 573.200 115.800 574.000 119.800 ;
        RECT 577.400 115.800 578.600 119.800 ;
        RECT 567.600 115.000 568.400 115.800 ;
        RECT 573.200 115.200 573.800 115.800 ;
        RECT 571.000 114.600 574.600 115.200 ;
        RECT 577.200 115.000 578.000 115.800 ;
        RECT 571.000 114.400 571.800 114.600 ;
        RECT 573.800 114.400 574.600 114.600 ;
        RECT 567.600 113.000 568.400 113.200 ;
        RECT 572.200 113.000 573.000 113.200 ;
        RECT 567.600 112.400 573.000 113.000 ;
        RECT 573.600 113.000 575.800 113.600 ;
        RECT 573.600 111.800 574.200 113.000 ;
        RECT 575.000 112.800 575.800 113.000 ;
        RECT 577.400 113.200 578.800 114.000 ;
        RECT 577.400 112.200 578.000 113.200 ;
        RECT 569.400 111.400 574.200 111.800 ;
        RECT 564.400 111.200 574.200 111.400 ;
        RECT 575.600 111.600 578.000 112.200 ;
        RECT 564.400 111.000 570.200 111.200 ;
        RECT 564.400 110.800 570.000 111.000 ;
        RECT 559.400 110.400 560.200 110.600 ;
        RECT 554.800 109.700 557.100 110.300 ;
        RECT 561.000 109.800 561.800 110.000 ;
        RECT 554.800 109.600 555.600 109.700 ;
        RECT 539.400 109.200 540.400 109.600 ;
        RECT 547.400 109.400 548.200 109.600 ;
        RECT 529.600 107.600 530.400 108.400 ;
        RECT 531.600 107.600 533.200 108.400 ;
        RECT 534.000 108.200 535.600 108.400 ;
        RECT 534.000 107.600 537.400 108.200 ;
        RECT 538.000 107.800 538.800 108.600 ;
        RECT 529.600 107.200 530.200 107.600 ;
        RECT 529.400 106.400 530.200 107.200 ;
        RECT 536.800 107.200 537.400 107.600 ;
        RECT 530.800 106.800 531.600 107.000 ;
        RECT 535.400 106.800 536.200 107.000 ;
        RECT 530.800 106.200 533.200 106.800 ;
        RECT 527.200 104.400 528.800 105.800 ;
        RECT 527.200 103.600 530.000 104.400 ;
        RECT 527.200 102.200 528.800 103.600 ;
        RECT 532.400 102.200 533.200 106.200 ;
        RECT 534.000 106.200 536.200 106.800 ;
        RECT 536.800 106.600 538.800 107.200 ;
        RECT 537.200 106.400 538.800 106.600 ;
        RECT 534.000 102.200 534.800 106.200 ;
        RECT 539.400 105.800 540.000 109.200 ;
        RECT 549.000 108.400 549.800 108.600 ;
        RECT 556.400 108.400 557.000 109.700 ;
        RECT 558.000 109.200 561.800 109.800 ;
        RECT 558.000 109.000 558.800 109.200 ;
        RECT 540.800 107.600 541.600 108.400 ;
        RECT 542.800 107.600 544.400 108.400 ;
        RECT 546.000 107.800 557.000 108.400 ;
        RECT 546.000 107.600 547.600 107.800 ;
        RECT 540.800 107.200 541.400 107.600 ;
        RECT 540.600 106.400 541.400 107.200 ;
        RECT 542.000 106.800 542.800 107.000 ;
        RECT 542.000 106.200 544.400 106.800 ;
        RECT 538.400 104.400 540.000 105.800 ;
        RECT 538.400 103.600 541.200 104.400 ;
        RECT 538.400 102.200 540.000 103.600 ;
        RECT 543.600 102.200 544.400 106.200 ;
        RECT 545.200 102.200 546.000 107.000 ;
        RECT 550.200 105.600 550.800 107.800 ;
        RECT 555.800 107.600 556.600 107.800 ;
        RECT 562.800 107.200 563.600 110.600 ;
        RECT 570.800 110.200 571.600 110.400 ;
        RECT 566.600 109.600 571.600 110.200 ;
        RECT 566.600 109.400 567.400 109.600 ;
        RECT 569.200 109.400 570.000 109.600 ;
        RECT 568.200 108.400 569.000 108.600 ;
        RECT 575.600 108.400 576.200 111.600 ;
        RECT 582.000 111.200 582.800 119.800 ;
        RECT 578.600 110.600 582.800 111.200 ;
        RECT 578.600 110.400 579.400 110.600 ;
        RECT 580.200 109.800 581.000 110.000 ;
        RECT 577.200 109.200 581.000 109.800 ;
        RECT 577.200 109.000 578.000 109.200 ;
        RECT 565.200 107.800 576.200 108.400 ;
        RECT 565.200 107.600 566.800 107.800 ;
        RECT 559.800 106.600 563.600 107.200 ;
        RECT 559.800 106.400 560.600 106.600 ;
        RECT 548.400 104.200 549.200 105.000 ;
        RECT 550.000 104.800 550.800 105.600 ;
        RECT 551.800 105.400 552.600 105.600 ;
        RECT 551.800 104.800 554.600 105.400 ;
        RECT 554.000 104.200 554.600 104.800 ;
        RECT 558.000 104.200 558.800 105.000 ;
        RECT 548.400 103.600 550.400 104.200 ;
        RECT 549.600 102.200 550.400 103.600 ;
        RECT 554.000 102.200 554.800 104.200 ;
        RECT 558.000 103.600 559.400 104.200 ;
        RECT 558.200 102.200 559.400 103.600 ;
        RECT 562.800 102.200 563.600 106.600 ;
        RECT 564.400 102.200 565.200 107.000 ;
        RECT 569.400 105.600 570.000 107.800 ;
        RECT 575.000 107.600 575.800 107.800 ;
        RECT 582.000 107.200 582.800 110.600 ;
        RECT 579.000 106.600 582.800 107.200 ;
        RECT 579.000 106.400 579.800 106.600 ;
        RECT 567.600 104.200 568.400 105.000 ;
        RECT 569.200 104.800 570.000 105.600 ;
        RECT 571.000 105.400 571.800 105.600 ;
        RECT 571.000 104.800 573.800 105.400 ;
        RECT 573.200 104.200 573.800 104.800 ;
        RECT 577.200 104.200 578.000 105.000 ;
        RECT 567.600 103.600 569.600 104.200 ;
        RECT 568.800 102.200 569.600 103.600 ;
        RECT 573.200 102.200 574.000 104.200 ;
        RECT 577.200 103.600 578.600 104.200 ;
        RECT 577.400 102.200 578.600 103.600 ;
        RECT 582.000 102.200 582.800 106.600 ;
        RECT 1.200 93.600 2.000 95.200 ;
        RECT 2.800 82.200 3.600 99.800 ;
        RECT 4.400 95.600 5.200 97.200 ;
        RECT 6.000 90.300 6.800 99.800 ;
        RECT 11.200 94.200 12.000 99.800 ;
        RECT 14.000 96.000 14.800 99.800 ;
        RECT 17.200 96.000 18.000 99.800 ;
        RECT 14.000 95.800 18.000 96.000 ;
        RECT 18.800 95.800 19.600 99.800 ;
        RECT 22.000 96.400 22.800 99.800 ;
        RECT 21.800 95.800 22.800 96.400 ;
        RECT 14.200 95.400 17.800 95.800 ;
        RECT 14.800 94.400 15.600 94.800 ;
        RECT 18.800 94.400 19.400 95.800 ;
        RECT 21.800 94.400 22.400 95.800 ;
        RECT 25.200 95.200 26.000 99.800 ;
        RECT 28.400 97.600 29.200 99.800 ;
        RECT 26.800 95.600 27.600 97.200 ;
        RECT 23.400 94.600 26.000 95.200 ;
        RECT 11.200 93.800 13.000 94.200 ;
        RECT 11.400 93.600 13.000 93.800 ;
        RECT 14.000 93.800 15.600 94.400 ;
        RECT 14.000 93.600 14.800 93.800 ;
        RECT 17.000 93.600 19.600 94.400 ;
        RECT 21.800 93.600 22.800 94.400 ;
        RECT 9.200 91.600 10.800 92.400 ;
        RECT 7.600 90.300 8.400 91.200 ;
        RECT 6.000 89.700 8.400 90.300 ;
        RECT 6.000 82.200 6.800 89.700 ;
        RECT 7.600 89.600 8.400 89.700 ;
        RECT 12.400 90.400 13.000 93.600 ;
        RECT 14.000 92.300 14.800 92.400 ;
        RECT 15.600 92.300 16.400 93.200 ;
        RECT 14.000 91.700 16.400 92.300 ;
        RECT 14.000 91.600 14.800 91.700 ;
        RECT 15.600 91.600 16.400 91.700 ;
        RECT 17.000 92.300 17.600 93.600 ;
        RECT 20.400 92.300 21.200 92.400 ;
        RECT 17.000 91.700 21.200 92.300 ;
        RECT 12.400 89.600 13.200 90.400 ;
        RECT 17.000 90.200 17.600 91.700 ;
        RECT 20.400 91.600 21.200 91.700 ;
        RECT 18.800 90.200 19.600 90.400 ;
        RECT 16.600 89.600 17.600 90.200 ;
        RECT 18.200 89.600 19.600 90.200 ;
        RECT 21.800 90.200 22.400 93.600 ;
        RECT 23.400 93.000 24.000 94.600 ;
        RECT 28.600 94.400 29.200 97.600 ;
        RECT 31.600 95.600 32.400 97.200 ;
        RECT 28.400 93.600 29.200 94.400 ;
        RECT 23.000 92.200 24.000 93.000 ;
        RECT 23.400 90.200 24.000 92.200 ;
        RECT 25.000 92.400 25.800 93.200 ;
        RECT 25.000 91.600 26.000 92.400 ;
        RECT 28.600 90.200 29.200 93.600 ;
        RECT 30.000 90.800 30.800 92.400 ;
        RECT 10.800 87.600 11.600 89.200 ;
        RECT 12.400 87.000 13.000 89.600 ;
        RECT 9.400 86.400 13.000 87.000 ;
        RECT 9.400 86.200 10.000 86.400 ;
        RECT 9.200 82.200 10.000 86.200 ;
        RECT 12.400 86.200 13.000 86.400 ;
        RECT 12.400 82.200 13.200 86.200 ;
        RECT 16.600 82.200 17.400 89.600 ;
        RECT 18.200 88.400 18.800 89.600 ;
        RECT 21.800 89.200 22.800 90.200 ;
        RECT 23.400 89.600 26.000 90.200 ;
        RECT 18.000 87.600 18.800 88.400 ;
        RECT 22.000 82.200 22.800 89.200 ;
        RECT 25.200 82.200 26.000 89.600 ;
        RECT 28.400 89.400 30.200 90.200 ;
        RECT 29.400 82.200 30.200 89.400 ;
        RECT 33.200 82.200 34.000 99.800 ;
        RECT 34.800 96.000 35.600 99.800 ;
        RECT 38.000 96.000 38.800 99.800 ;
        RECT 34.800 95.800 38.800 96.000 ;
        RECT 39.600 96.300 40.400 99.800 ;
        RECT 41.200 96.300 42.000 97.200 ;
        RECT 35.000 95.400 38.600 95.800 ;
        RECT 39.600 95.700 42.000 96.300 ;
        RECT 35.600 94.400 36.400 94.800 ;
        RECT 39.600 94.400 40.200 95.700 ;
        RECT 41.200 95.600 42.000 95.700 ;
        RECT 34.800 93.800 36.400 94.400 ;
        RECT 37.800 94.300 40.400 94.400 ;
        RECT 41.200 94.300 42.000 94.400 ;
        RECT 34.800 93.600 35.600 93.800 ;
        RECT 37.800 93.700 42.000 94.300 ;
        RECT 37.800 93.600 40.400 93.700 ;
        RECT 41.200 93.600 42.000 93.700 ;
        RECT 36.400 91.600 37.200 93.200 ;
        RECT 37.800 90.200 38.400 93.600 ;
        RECT 39.600 90.200 40.400 90.400 ;
        RECT 37.400 89.600 38.400 90.200 ;
        RECT 39.000 89.600 40.400 90.200 ;
        RECT 42.800 90.300 43.600 99.800 ;
        RECT 44.400 95.800 45.200 99.800 ;
        RECT 46.000 96.000 46.800 99.800 ;
        RECT 49.200 96.000 50.000 99.800 ;
        RECT 46.000 95.800 50.000 96.000 ;
        RECT 44.600 94.400 45.200 95.800 ;
        RECT 46.200 95.400 49.800 95.800 ;
        RECT 50.800 95.600 51.600 97.200 ;
        RECT 48.400 94.400 49.200 94.800 ;
        RECT 44.400 93.600 47.000 94.400 ;
        RECT 48.400 94.300 50.000 94.400 ;
        RECT 50.900 94.300 51.500 95.600 ;
        RECT 48.400 93.800 51.500 94.300 ;
        RECT 49.200 93.700 51.500 93.800 ;
        RECT 49.200 93.600 50.000 93.700 ;
        RECT 44.400 90.300 45.200 90.400 ;
        RECT 42.800 90.200 45.200 90.300 ;
        RECT 46.400 90.200 47.000 93.600 ;
        RECT 47.600 92.300 48.400 93.200 ;
        RECT 50.800 92.300 51.600 92.400 ;
        RECT 47.600 91.700 51.600 92.300 ;
        RECT 47.600 91.600 48.400 91.700 ;
        RECT 50.800 91.600 51.600 91.700 ;
        RECT 42.800 89.700 45.800 90.200 ;
        RECT 37.400 82.200 38.200 89.600 ;
        RECT 39.000 88.400 39.600 89.600 ;
        RECT 38.800 87.600 39.600 88.400 ;
        RECT 42.800 82.200 43.600 89.700 ;
        RECT 44.400 89.600 45.800 89.700 ;
        RECT 46.400 89.600 47.400 90.200 ;
        RECT 45.200 88.400 45.800 89.600 ;
        RECT 45.200 87.600 46.000 88.400 ;
        RECT 46.600 86.400 47.400 89.600 ;
        RECT 46.600 85.600 48.400 86.400 ;
        RECT 46.600 82.200 47.400 85.600 ;
        RECT 52.400 82.200 53.200 99.800 ;
        RECT 57.600 96.400 58.400 99.800 ;
        RECT 60.600 96.400 61.400 97.200 ;
        RECT 57.600 95.600 59.600 96.400 ;
        RECT 60.400 95.600 61.200 96.400 ;
        RECT 62.000 95.800 62.800 99.800 ;
        RECT 66.800 96.000 67.600 99.800 ;
        RECT 70.000 96.000 70.800 99.800 ;
        RECT 66.800 95.800 70.800 96.000 ;
        RECT 71.600 95.800 72.400 99.800 ;
        RECT 75.800 96.400 76.600 99.800 ;
        RECT 80.600 96.400 81.400 99.800 ;
        RECT 74.800 95.800 76.600 96.400 ;
        RECT 79.600 95.800 81.400 96.400 ;
        RECT 57.600 94.200 58.400 95.600 ;
        RECT 57.600 93.800 59.400 94.200 ;
        RECT 57.800 93.600 59.400 93.800 ;
        RECT 55.600 91.600 57.200 92.400 ;
        RECT 54.000 89.600 54.800 91.200 ;
        RECT 58.800 90.400 59.400 93.600 ;
        RECT 62.200 92.400 62.800 95.800 ;
        RECT 67.000 95.400 70.600 95.800 ;
        RECT 67.600 94.400 68.400 94.800 ;
        RECT 71.600 94.400 72.200 95.800 ;
        RECT 63.600 92.800 64.400 94.400 ;
        RECT 66.800 93.800 68.400 94.400 ;
        RECT 66.800 93.600 67.600 93.800 ;
        RECT 69.800 93.600 72.400 94.400 ;
        RECT 73.200 93.600 74.000 95.200 ;
        RECT 60.400 92.200 61.200 92.400 ;
        RECT 62.000 92.200 62.800 92.400 ;
        RECT 65.200 92.200 66.000 92.400 ;
        RECT 60.400 91.600 62.800 92.200 ;
        RECT 64.400 91.600 66.000 92.200 ;
        RECT 68.400 91.600 69.200 93.200 ;
        RECT 69.800 92.300 70.400 93.600 ;
        RECT 73.200 92.300 74.000 92.400 ;
        RECT 69.800 91.700 74.000 92.300 ;
        RECT 58.800 89.600 59.600 90.400 ;
        RECT 60.600 90.200 61.200 91.600 ;
        RECT 64.400 91.200 65.200 91.600 ;
        RECT 69.800 90.200 70.400 91.700 ;
        RECT 73.200 91.600 74.000 91.700 ;
        RECT 71.600 90.200 72.400 90.400 ;
        RECT 57.200 87.600 58.000 89.200 ;
        RECT 58.800 87.000 59.400 89.600 ;
        RECT 55.800 86.400 59.400 87.000 ;
        RECT 55.800 86.200 56.400 86.400 ;
        RECT 55.600 82.200 56.400 86.200 ;
        RECT 58.800 86.200 59.400 86.400 ;
        RECT 58.800 82.200 59.600 86.200 ;
        RECT 60.400 82.200 61.200 90.200 ;
        RECT 62.000 89.600 66.000 90.200 ;
        RECT 62.000 82.200 62.800 89.600 ;
        RECT 65.200 82.200 66.000 89.600 ;
        RECT 69.400 89.600 70.400 90.200 ;
        RECT 71.000 89.600 72.400 90.200 ;
        RECT 69.400 82.200 70.200 89.600 ;
        RECT 71.000 88.400 71.600 89.600 ;
        RECT 70.800 87.600 71.600 88.400 ;
        RECT 74.800 82.200 75.600 95.800 ;
        RECT 78.000 93.600 78.800 95.200 ;
        RECT 79.600 92.300 80.400 95.800 ;
        RECT 81.200 92.300 82.000 92.400 ;
        RECT 79.600 91.700 82.000 92.300 ;
        RECT 76.400 88.800 77.200 90.400 ;
        RECT 79.600 82.200 80.400 91.700 ;
        RECT 81.200 91.600 82.000 91.700 ;
        RECT 81.200 90.300 82.000 90.400 ;
        RECT 82.800 90.300 83.600 99.800 ;
        RECT 86.600 98.400 87.400 99.800 ;
        RECT 86.600 97.600 88.400 98.400 ;
        RECT 84.400 95.600 85.200 97.200 ;
        RECT 86.600 96.400 87.400 97.600 ;
        RECT 93.400 96.400 94.200 99.800 ;
        RECT 86.600 95.800 88.400 96.400 ;
        RECT 81.200 89.700 83.600 90.300 ;
        RECT 81.200 88.800 82.000 89.700 ;
        RECT 82.800 82.200 83.600 89.700 ;
        RECT 84.400 90.300 85.200 90.400 ;
        RECT 86.000 90.300 86.800 90.400 ;
        RECT 84.400 89.700 86.800 90.300 ;
        RECT 84.400 89.600 85.200 89.700 ;
        RECT 86.000 88.800 86.800 89.700 ;
        RECT 87.600 82.200 88.400 95.800 ;
        RECT 92.400 95.600 94.800 96.400 ;
        RECT 98.800 95.800 99.600 99.800 ;
        RECT 100.200 96.400 101.000 97.200 ;
        RECT 89.200 93.600 90.000 95.200 ;
        RECT 90.800 93.600 91.600 95.200 ;
        RECT 92.400 82.200 93.200 95.600 ;
        RECT 97.200 92.800 98.000 94.400 ;
        RECT 98.800 94.300 99.400 95.800 ;
        RECT 100.400 95.600 101.200 96.400 ;
        RECT 105.200 95.800 106.000 99.800 ;
        RECT 106.600 96.400 107.400 97.200 ;
        RECT 103.600 94.300 104.400 94.400 ;
        RECT 98.800 93.700 104.400 94.300 ;
        RECT 95.600 92.300 96.400 92.400 ;
        RECT 94.100 92.200 96.400 92.300 ;
        RECT 98.800 92.200 99.400 93.700 ;
        RECT 103.600 92.800 104.400 93.700 ;
        RECT 100.400 92.200 101.200 92.400 ;
        RECT 94.100 91.700 97.200 92.200 ;
        RECT 94.100 90.400 94.700 91.700 ;
        RECT 95.600 91.600 97.200 91.700 ;
        RECT 98.800 91.600 101.200 92.200 ;
        RECT 102.000 92.200 102.800 92.400 ;
        RECT 105.200 92.200 105.800 95.800 ;
        RECT 106.800 95.600 107.600 96.400 ;
        RECT 111.600 95.800 112.400 99.800 ;
        RECT 113.000 96.400 113.800 97.200 ;
        RECT 113.200 96.300 114.000 96.400 ;
        RECT 114.800 96.300 115.600 97.200 ;
        RECT 110.000 92.800 110.800 94.400 ;
        RECT 106.800 92.200 107.600 92.400 ;
        RECT 102.000 91.600 103.600 92.200 ;
        RECT 105.200 91.600 107.600 92.200 ;
        RECT 108.400 92.200 109.200 92.400 ;
        RECT 111.600 92.200 112.200 95.800 ;
        RECT 113.200 95.700 115.600 96.300 ;
        RECT 113.200 95.600 114.000 95.700 ;
        RECT 114.800 95.600 115.600 95.700 ;
        RECT 113.200 92.200 114.000 92.400 ;
        RECT 108.400 91.600 110.000 92.200 ;
        RECT 111.600 91.600 114.000 92.200 ;
        RECT 96.400 91.200 97.200 91.600 ;
        RECT 94.000 88.800 94.800 90.400 ;
        RECT 100.400 90.200 101.000 91.600 ;
        RECT 102.800 91.200 103.600 91.600 ;
        RECT 106.800 90.200 107.400 91.600 ;
        RECT 109.200 91.200 110.000 91.600 ;
        RECT 113.200 90.200 113.800 91.600 ;
        RECT 116.400 90.300 117.200 99.800 ;
        RECT 118.000 95.800 118.800 99.800 ;
        RECT 119.600 96.000 120.400 99.800 ;
        RECT 122.800 96.000 123.600 99.800 ;
        RECT 124.600 96.400 125.400 97.200 ;
        RECT 119.600 95.800 123.600 96.000 ;
        RECT 118.200 94.400 118.800 95.800 ;
        RECT 119.800 95.400 123.400 95.800 ;
        RECT 124.400 95.600 125.200 96.400 ;
        RECT 126.000 95.800 126.800 99.800 ;
        RECT 132.400 97.800 133.200 99.800 ;
        RECT 122.000 94.400 122.800 94.800 ;
        RECT 118.000 93.600 120.600 94.400 ;
        RECT 122.000 93.800 123.600 94.400 ;
        RECT 122.800 93.600 123.600 93.800 ;
        RECT 118.000 90.300 118.800 90.400 ;
        RECT 116.400 90.200 118.800 90.300 ;
        RECT 120.000 90.200 120.600 93.600 ;
        RECT 121.200 91.600 122.000 93.200 ;
        RECT 124.400 92.200 125.200 92.400 ;
        RECT 126.200 92.200 126.800 95.800 ;
        RECT 130.800 95.600 131.600 97.200 ;
        RECT 132.600 94.400 133.200 97.800 ;
        RECT 140.400 95.800 141.200 99.800 ;
        RECT 142.000 96.000 142.800 99.800 ;
        RECT 145.200 96.000 146.000 99.800 ;
        RECT 142.000 95.800 146.000 96.000 ;
        RECT 146.800 95.800 147.600 99.800 ;
        RECT 148.400 96.000 149.200 99.800 ;
        RECT 151.600 96.000 152.400 99.800 ;
        RECT 148.400 95.800 152.400 96.000 ;
        RECT 153.800 96.400 154.600 99.800 ;
        RECT 153.800 95.800 155.600 96.400 ;
        RECT 140.600 94.400 141.200 95.800 ;
        RECT 142.200 95.400 145.800 95.800 ;
        RECT 144.400 94.400 145.200 94.800 ;
        RECT 147.000 94.400 147.600 95.800 ;
        RECT 148.600 95.400 152.200 95.800 ;
        RECT 150.800 94.400 151.600 94.800 ;
        RECT 127.600 94.300 128.400 94.400 ;
        RECT 132.400 94.300 133.200 94.400 ;
        RECT 127.600 93.700 133.200 94.300 ;
        RECT 127.600 92.800 128.400 93.700 ;
        RECT 132.400 93.600 133.200 93.700 ;
        RECT 140.400 93.600 143.000 94.400 ;
        RECT 144.400 93.800 146.000 94.400 ;
        RECT 145.200 93.600 146.000 93.800 ;
        RECT 146.800 93.600 149.400 94.400 ;
        RECT 150.800 94.300 152.400 94.400 ;
        RECT 154.800 94.300 155.600 95.800 ;
        RECT 150.800 93.800 155.600 94.300 ;
        RECT 151.600 93.700 155.600 93.800 ;
        RECT 151.600 93.600 152.400 93.700 ;
        RECT 129.200 92.200 130.000 92.400 ;
        RECT 124.400 91.600 126.800 92.200 ;
        RECT 128.400 91.600 130.000 92.200 ;
        RECT 124.600 90.200 125.200 91.600 ;
        RECT 128.400 91.200 129.200 91.600 ;
        RECT 132.600 90.200 133.200 93.600 ;
        RECT 134.000 90.800 134.800 92.400 ;
        RECT 140.400 90.200 141.200 90.400 ;
        RECT 142.400 90.200 143.000 93.600 ;
        RECT 143.600 92.300 144.400 93.200 ;
        RECT 145.200 92.300 146.000 92.400 ;
        RECT 143.600 91.700 146.000 92.300 ;
        RECT 143.600 91.600 144.400 91.700 ;
        RECT 145.200 91.600 146.000 91.700 ;
        RECT 146.800 90.200 147.600 90.400 ;
        RECT 148.800 90.200 149.400 93.600 ;
        RECT 150.000 91.600 150.800 93.200 ;
        RECT 95.600 89.600 99.600 90.200 ;
        RECT 95.600 82.200 96.400 89.600 ;
        RECT 98.800 82.200 99.600 89.600 ;
        RECT 100.400 82.200 101.200 90.200 ;
        RECT 102.000 89.600 106.000 90.200 ;
        RECT 102.000 82.200 102.800 89.600 ;
        RECT 105.200 82.200 106.000 89.600 ;
        RECT 106.800 82.200 107.600 90.200 ;
        RECT 108.400 89.600 112.400 90.200 ;
        RECT 108.400 82.200 109.200 89.600 ;
        RECT 111.600 82.200 112.400 89.600 ;
        RECT 113.200 88.300 114.000 90.200 ;
        RECT 116.400 89.700 119.400 90.200 ;
        RECT 114.800 88.300 115.600 88.400 ;
        RECT 113.200 87.700 115.600 88.300 ;
        RECT 113.200 82.200 114.000 87.700 ;
        RECT 114.800 87.600 115.600 87.700 ;
        RECT 116.400 82.200 117.200 89.700 ;
        RECT 118.000 89.600 119.400 89.700 ;
        RECT 120.000 89.600 121.000 90.200 ;
        RECT 118.800 88.400 119.400 89.600 ;
        RECT 118.800 87.600 119.600 88.400 ;
        RECT 120.200 82.200 121.000 89.600 ;
        RECT 124.400 82.200 125.200 90.200 ;
        RECT 126.000 89.600 130.000 90.200 ;
        RECT 126.000 82.200 126.800 89.600 ;
        RECT 129.200 82.200 130.000 89.600 ;
        RECT 132.400 89.400 134.200 90.200 ;
        RECT 140.400 89.600 141.800 90.200 ;
        RECT 142.400 89.600 143.400 90.200 ;
        RECT 146.800 89.600 148.200 90.200 ;
        RECT 148.800 89.600 149.800 90.200 ;
        RECT 133.400 82.200 134.200 89.400 ;
        RECT 141.200 88.400 141.800 89.600 ;
        RECT 141.200 87.600 142.000 88.400 ;
        RECT 142.600 84.400 143.400 89.600 ;
        RECT 147.600 88.400 148.200 89.600 ;
        RECT 147.600 87.600 148.400 88.400 ;
        RECT 142.600 83.600 144.400 84.400 ;
        RECT 142.600 82.200 143.400 83.600 ;
        RECT 149.000 82.200 149.800 89.600 ;
        RECT 153.200 88.800 154.000 90.400 ;
        RECT 154.800 82.200 155.600 93.700 ;
        RECT 156.400 93.600 157.200 95.200 ;
        RECT 158.000 95.000 158.800 99.800 ;
        RECT 162.400 98.400 163.200 99.800 ;
        RECT 161.200 97.800 163.200 98.400 ;
        RECT 166.800 97.800 167.600 99.800 ;
        RECT 171.000 98.400 172.200 99.800 ;
        RECT 170.800 97.800 172.200 98.400 ;
        RECT 161.200 97.000 162.000 97.800 ;
        RECT 166.800 97.200 167.400 97.800 ;
        RECT 162.800 96.400 163.600 97.200 ;
        RECT 164.600 96.600 167.400 97.200 ;
        RECT 170.800 97.000 171.600 97.800 ;
        RECT 164.600 96.400 165.400 96.600 ;
        RECT 158.800 94.200 160.400 94.400 ;
        RECT 163.000 94.200 163.600 96.400 ;
        RECT 172.600 95.400 173.400 95.600 ;
        RECT 175.600 95.400 176.400 99.800 ;
        RECT 172.600 94.800 176.400 95.400 ;
        RECT 166.000 94.200 166.800 94.400 ;
        RECT 168.600 94.200 169.400 94.400 ;
        RECT 158.800 93.600 169.800 94.200 ;
        RECT 161.800 93.400 162.600 93.600 ;
        RECT 160.200 92.400 161.000 92.600 ;
        RECT 162.800 92.400 163.600 92.600 ;
        RECT 169.200 92.400 169.800 93.600 ;
        RECT 170.800 92.800 171.600 93.000 ;
        RECT 160.200 91.800 165.200 92.400 ;
        RECT 164.400 91.600 165.200 91.800 ;
        RECT 169.200 91.600 170.000 92.400 ;
        RECT 170.800 92.200 174.600 92.800 ;
        RECT 173.800 92.000 174.600 92.200 ;
        RECT 158.000 91.000 163.600 91.200 ;
        RECT 158.000 90.800 163.800 91.000 ;
        RECT 158.000 90.600 167.800 90.800 ;
        RECT 158.000 82.200 158.800 90.600 ;
        RECT 163.000 90.200 167.800 90.600 ;
        RECT 161.200 89.000 166.600 89.600 ;
        RECT 161.200 88.800 162.000 89.000 ;
        RECT 165.800 88.800 166.600 89.000 ;
        RECT 167.200 89.000 167.800 90.200 ;
        RECT 169.200 90.400 169.800 91.600 ;
        RECT 172.200 91.400 173.000 91.600 ;
        RECT 175.600 91.400 176.400 94.800 ;
        RECT 178.800 97.800 179.600 99.800 ;
        RECT 183.600 97.800 184.400 99.800 ;
        RECT 178.800 94.400 179.400 97.800 ;
        RECT 180.400 95.600 181.200 97.200 ;
        RECT 182.000 95.600 182.800 97.200 ;
        RECT 183.800 96.300 184.400 97.800 ;
        RECT 188.400 97.800 189.200 99.800 ;
        RECT 193.200 97.800 194.000 99.800 ;
        RECT 186.800 96.300 187.600 96.400 ;
        RECT 183.700 95.700 187.600 96.300 ;
        RECT 178.800 94.300 179.600 94.400 ;
        RECT 182.100 94.300 182.700 95.600 ;
        RECT 183.800 94.400 184.400 95.700 ;
        RECT 186.800 95.600 187.600 95.700 ;
        RECT 178.800 93.700 182.700 94.300 ;
        RECT 178.800 93.600 179.600 93.700 ;
        RECT 183.600 93.600 184.400 94.400 ;
        RECT 172.200 90.800 176.400 91.400 ;
        RECT 177.200 90.800 178.000 92.400 ;
        RECT 169.200 89.800 171.600 90.400 ;
        RECT 168.600 89.000 169.400 89.200 ;
        RECT 167.200 88.400 169.400 89.000 ;
        RECT 171.000 88.800 171.600 89.800 ;
        RECT 171.000 88.000 172.400 88.800 ;
        RECT 164.600 87.400 165.400 87.600 ;
        RECT 167.400 87.400 168.200 87.600 ;
        RECT 161.200 86.200 162.000 87.000 ;
        RECT 164.600 86.800 168.200 87.400 ;
        RECT 166.800 86.200 167.400 86.800 ;
        RECT 170.800 86.200 171.600 87.000 ;
        RECT 161.200 85.600 163.200 86.200 ;
        RECT 162.400 82.200 163.200 85.600 ;
        RECT 166.800 82.200 167.600 86.200 ;
        RECT 171.000 82.200 172.200 86.200 ;
        RECT 175.600 82.200 176.400 90.800 ;
        RECT 178.800 90.200 179.400 93.600 ;
        RECT 183.800 90.200 184.400 93.600 ;
        RECT 188.400 94.400 189.000 97.800 ;
        RECT 190.000 95.600 190.800 97.200 ;
        RECT 191.600 95.600 192.400 97.200 ;
        RECT 188.400 94.300 189.200 94.400 ;
        RECT 191.700 94.300 192.300 95.600 ;
        RECT 193.400 94.400 194.000 97.800 ;
        RECT 196.400 96.000 197.200 99.800 ;
        RECT 199.600 96.000 200.400 99.800 ;
        RECT 196.400 95.800 200.400 96.000 ;
        RECT 201.200 95.800 202.000 99.800 ;
        RECT 202.800 95.800 203.600 99.800 ;
        RECT 204.400 96.000 205.200 99.800 ;
        RECT 207.600 96.000 208.400 99.800 ;
        RECT 204.400 95.800 208.400 96.000 ;
        RECT 196.600 95.400 200.200 95.800 ;
        RECT 197.200 94.400 198.000 94.800 ;
        RECT 201.200 94.400 201.800 95.800 ;
        RECT 203.000 94.400 203.600 95.800 ;
        RECT 204.600 95.400 208.200 95.800 ;
        RECT 209.200 95.600 210.000 97.200 ;
        RECT 206.800 94.400 207.600 94.800 ;
        RECT 188.400 93.700 192.300 94.300 ;
        RECT 193.200 94.300 194.000 94.400 ;
        RECT 194.800 94.300 195.600 94.400 ;
        RECT 193.200 93.700 195.600 94.300 ;
        RECT 188.400 93.600 189.200 93.700 ;
        RECT 193.200 93.600 194.000 93.700 ;
        RECT 194.800 93.600 195.600 93.700 ;
        RECT 196.400 93.800 198.000 94.400 ;
        RECT 196.400 93.600 197.200 93.800 ;
        RECT 199.400 93.600 202.000 94.400 ;
        RECT 202.800 93.600 205.400 94.400 ;
        RECT 206.800 94.300 208.400 94.400 ;
        RECT 209.300 94.300 209.900 95.600 ;
        RECT 206.800 93.800 209.900 94.300 ;
        RECT 207.600 93.700 209.900 93.800 ;
        RECT 210.800 94.300 211.600 99.800 ;
        RECT 215.000 95.800 216.600 99.800 ;
        RECT 223.000 98.400 223.800 99.800 ;
        RECT 223.000 97.600 224.400 98.400 ;
        RECT 223.000 96.400 223.800 97.600 ;
        RECT 222.000 95.800 223.800 96.400 ;
        RECT 225.200 95.800 226.000 99.800 ;
        RECT 226.800 96.000 227.600 99.800 ;
        RECT 230.000 96.000 230.800 99.800 ;
        RECT 226.800 95.800 230.800 96.000 ;
        RECT 214.000 94.300 214.800 94.400 ;
        RECT 210.800 93.700 214.800 94.300 ;
        RECT 207.600 93.600 208.400 93.700 ;
        RECT 185.200 90.800 186.000 92.400 ;
        RECT 186.800 90.800 187.600 92.400 ;
        RECT 188.400 90.200 189.000 93.600 ;
        RECT 193.400 90.200 194.000 93.600 ;
        RECT 194.800 90.800 195.600 92.400 ;
        RECT 198.000 91.600 198.800 93.200 ;
        RECT 199.400 92.300 200.000 93.600 ;
        RECT 202.800 92.300 203.600 92.400 ;
        RECT 199.400 91.700 203.600 92.300 ;
        RECT 199.400 90.200 200.000 91.700 ;
        RECT 202.800 91.600 203.600 91.700 ;
        RECT 201.200 90.200 202.000 90.400 ;
        RECT 177.800 89.400 179.600 90.200 ;
        RECT 183.600 89.400 185.400 90.200 ;
        RECT 177.800 82.200 178.600 89.400 ;
        RECT 184.600 82.200 185.400 89.400 ;
        RECT 187.400 89.400 189.200 90.200 ;
        RECT 193.200 89.400 195.000 90.200 ;
        RECT 187.400 82.200 188.200 89.400 ;
        RECT 194.200 82.200 195.000 89.400 ;
        RECT 199.000 89.600 200.000 90.200 ;
        RECT 200.600 89.600 202.000 90.200 ;
        RECT 202.800 90.200 203.600 90.400 ;
        RECT 204.800 90.200 205.400 93.600 ;
        RECT 206.000 91.600 206.800 93.200 ;
        RECT 202.800 89.600 204.200 90.200 ;
        RECT 204.800 89.600 205.800 90.200 ;
        RECT 199.000 82.200 199.800 89.600 ;
        RECT 200.600 88.400 201.200 89.600 ;
        RECT 200.400 87.600 201.200 88.400 ;
        RECT 203.600 88.400 204.200 89.600 ;
        RECT 203.600 87.600 204.400 88.400 ;
        RECT 205.000 84.400 205.800 89.600 ;
        RECT 205.000 83.600 206.800 84.400 ;
        RECT 205.000 82.200 205.800 83.600 ;
        RECT 210.800 82.200 211.600 93.700 ;
        RECT 214.000 93.600 214.800 93.700 ;
        RECT 214.200 93.200 214.800 93.600 ;
        RECT 214.200 92.400 215.000 93.200 ;
        RECT 215.600 92.400 216.200 95.800 ;
        RECT 217.200 92.800 218.000 94.400 ;
        RECT 220.400 93.600 221.200 95.200 ;
        RECT 212.400 90.800 213.200 92.400 ;
        RECT 215.600 91.600 216.400 92.400 ;
        RECT 218.800 92.200 219.600 92.400 ;
        RECT 218.000 91.600 219.600 92.200 ;
        RECT 215.600 91.400 216.200 91.600 ;
        RECT 214.200 90.800 216.200 91.400 ;
        RECT 218.000 91.200 218.800 91.600 ;
        RECT 214.200 90.200 214.800 90.800 ;
        RECT 212.400 82.800 213.200 90.200 ;
        RECT 214.000 83.400 214.800 90.200 ;
        RECT 215.600 89.600 219.600 90.200 ;
        RECT 215.600 82.800 216.400 89.600 ;
        RECT 212.400 82.200 216.400 82.800 ;
        RECT 218.800 82.200 219.600 89.600 ;
        RECT 222.000 82.200 222.800 95.800 ;
        RECT 225.400 94.400 226.000 95.800 ;
        RECT 227.000 95.400 230.600 95.800 ;
        RECT 229.200 94.400 230.000 94.800 ;
        RECT 225.200 93.600 227.800 94.400 ;
        RECT 229.200 93.800 230.800 94.400 ;
        RECT 230.000 93.600 230.800 93.800 ;
        RECT 227.200 92.400 227.800 93.600 ;
        RECT 226.800 91.600 227.800 92.400 ;
        RECT 228.400 92.300 229.200 93.200 ;
        RECT 231.600 92.300 232.400 99.800 ;
        RECT 233.200 95.600 234.000 97.200 ;
        RECT 237.800 95.800 239.400 99.800 ;
        RECT 244.400 97.800 245.200 99.800 ;
        RECT 236.400 92.800 237.200 94.400 ;
        RECT 238.200 92.400 238.800 95.800 ;
        RECT 242.800 95.600 243.600 97.200 ;
        RECT 244.600 94.400 245.200 97.800 ;
        RECT 239.600 94.300 240.400 94.400 ;
        RECT 241.200 94.300 242.000 94.400 ;
        RECT 239.600 93.700 242.000 94.300 ;
        RECT 239.600 93.600 240.400 93.700 ;
        RECT 241.200 93.600 242.000 93.700 ;
        RECT 244.400 93.600 245.200 94.400 ;
        RECT 247.600 97.000 248.400 99.000 ;
        RECT 247.600 94.800 248.200 97.000 ;
        RECT 251.800 96.000 252.600 99.000 ;
        RECT 251.800 95.400 253.400 96.000 ;
        RECT 252.600 95.000 253.400 95.400 ;
        RECT 257.200 95.800 258.000 99.800 ;
        RECT 261.600 96.200 263.200 99.800 ;
        RECT 257.200 95.200 259.600 95.800 ;
        RECT 258.800 95.000 259.600 95.200 ;
        RECT 247.600 94.200 251.800 94.800 ;
        RECT 239.600 93.200 240.200 93.600 ;
        RECT 239.400 92.400 240.200 93.200 ;
        RECT 228.400 91.700 232.400 92.300 ;
        RECT 228.400 91.600 229.200 91.700 ;
        RECT 223.600 88.800 224.400 90.400 ;
        RECT 225.200 90.200 226.000 90.400 ;
        RECT 227.200 90.200 227.800 91.600 ;
        RECT 225.200 89.600 226.600 90.200 ;
        RECT 227.200 89.600 228.200 90.200 ;
        RECT 226.000 88.400 226.600 89.600 ;
        RECT 226.000 87.600 226.800 88.400 ;
        RECT 227.400 82.200 228.200 89.600 ;
        RECT 231.600 82.200 232.400 91.700 ;
        RECT 234.800 92.200 235.600 92.400 ;
        RECT 234.800 91.600 236.400 92.200 ;
        RECT 238.000 91.600 238.800 92.400 ;
        RECT 235.600 91.200 236.400 91.600 ;
        RECT 238.200 91.400 238.800 91.600 ;
        RECT 241.200 92.300 242.000 92.400 ;
        RECT 244.600 92.300 245.200 93.600 ;
        RECT 250.800 93.800 251.800 94.200 ;
        RECT 252.800 94.400 253.400 95.000 ;
        RECT 260.200 94.800 261.000 95.600 ;
        RECT 260.200 94.400 260.800 94.800 ;
        RECT 252.800 94.300 254.800 94.400 ;
        RECT 255.600 94.300 256.400 94.400 ;
        RECT 241.200 91.700 245.200 92.300 ;
        RECT 238.200 90.800 240.200 91.400 ;
        RECT 241.200 90.800 242.000 91.700 ;
        RECT 239.600 90.200 240.200 90.800 ;
        RECT 244.600 90.200 245.200 91.700 ;
        RECT 246.000 90.800 246.800 92.400 ;
        RECT 247.600 91.600 248.400 93.200 ;
        RECT 249.200 91.600 250.000 93.200 ;
        RECT 250.800 93.000 252.200 93.800 ;
        RECT 252.800 93.700 256.400 94.300 ;
        RECT 252.800 93.600 254.800 93.700 ;
        RECT 255.600 93.600 256.400 93.700 ;
        RECT 257.200 93.600 258.800 94.400 ;
        RECT 260.000 93.600 260.800 94.400 ;
        RECT 250.800 91.000 251.400 93.000 ;
        RECT 247.600 90.400 251.400 91.000 ;
        RECT 234.800 89.600 238.800 90.200 ;
        RECT 234.800 82.200 235.600 89.600 ;
        RECT 238.000 82.800 238.800 89.600 ;
        RECT 239.600 83.400 240.400 90.200 ;
        RECT 241.200 82.800 242.000 90.200 ;
        RECT 244.400 89.400 246.200 90.200 ;
        RECT 238.000 82.200 242.000 82.800 ;
        RECT 245.400 82.200 246.200 89.400 ;
        RECT 247.600 87.000 248.200 90.400 ;
        RECT 252.800 89.800 253.400 93.600 ;
        RECT 261.600 92.800 262.200 96.200 ;
        RECT 266.800 95.800 267.600 99.800 ;
        RECT 271.000 98.400 271.800 99.800 ;
        RECT 270.000 97.600 271.800 98.400 ;
        RECT 271.000 96.400 271.800 97.600 ;
        RECT 262.800 95.400 264.400 95.600 ;
        RECT 262.800 94.800 264.800 95.400 ;
        RECT 265.400 95.200 267.600 95.800 ;
        RECT 270.000 95.800 271.800 96.400 ;
        RECT 265.400 95.000 266.200 95.200 ;
        RECT 264.200 94.400 264.800 94.800 ;
        RECT 262.800 93.400 263.600 94.200 ;
        RECT 264.200 93.800 267.600 94.400 ;
        RECT 266.000 93.600 267.600 93.800 ;
        RECT 268.400 93.600 269.200 95.200 ;
        RECT 261.200 92.400 262.200 92.800 ;
        RECT 254.000 90.800 254.800 92.400 ;
        RECT 260.400 92.200 262.200 92.400 ;
        RECT 263.000 92.800 263.600 93.400 ;
        RECT 263.000 92.200 265.600 92.800 ;
        RECT 260.400 91.600 261.800 92.200 ;
        RECT 264.800 92.000 265.600 92.200 ;
        RECT 261.200 90.400 261.800 91.600 ;
        RECT 262.600 91.400 263.400 91.600 ;
        RECT 262.600 90.800 266.000 91.400 ;
        RECT 260.400 90.200 261.800 90.400 ;
        RECT 265.400 90.200 266.000 90.800 ;
        RECT 251.800 89.200 253.400 89.800 ;
        RECT 257.200 89.600 259.600 90.200 ;
        RECT 260.400 89.600 263.200 90.200 ;
        RECT 247.600 83.000 248.400 87.000 ;
        RECT 251.800 82.200 252.600 89.200 ;
        RECT 257.200 82.200 258.000 89.600 ;
        RECT 258.800 89.400 259.600 89.600 ;
        RECT 261.600 82.200 263.200 89.600 ;
        RECT 265.400 89.600 267.600 90.200 ;
        RECT 265.400 89.400 266.200 89.600 ;
        RECT 266.800 82.200 267.600 89.600 ;
        RECT 270.000 82.200 270.800 95.800 ;
        RECT 271.600 90.300 272.400 90.400 ;
        RECT 273.200 90.300 274.000 99.800 ;
        RECT 274.800 95.600 275.600 97.200 ;
        RECT 278.000 96.400 278.800 99.800 ;
        RECT 277.800 95.800 278.800 96.400 ;
        RECT 277.800 94.400 278.400 95.800 ;
        RECT 281.200 95.200 282.000 99.800 ;
        RECT 283.400 96.400 284.200 99.800 ;
        RECT 287.600 98.300 288.400 98.400 ;
        RECT 292.400 98.300 293.200 99.800 ;
        RECT 287.600 97.700 293.200 98.300 ;
        RECT 287.600 97.600 288.400 97.700 ;
        RECT 283.400 95.800 285.200 96.400 ;
        RECT 292.400 95.800 293.200 97.700 ;
        RECT 294.000 96.000 294.800 99.800 ;
        RECT 297.200 96.000 298.000 99.800 ;
        RECT 301.400 96.400 302.200 99.800 ;
        RECT 294.000 95.800 298.000 96.000 ;
        RECT 300.400 95.800 302.200 96.400 ;
        RECT 279.400 94.600 282.000 95.200 ;
        RECT 276.400 94.300 277.200 94.400 ;
        RECT 277.800 94.300 278.800 94.400 ;
        RECT 276.400 93.700 278.800 94.300 ;
        RECT 276.400 93.600 277.200 93.700 ;
        RECT 277.800 93.600 278.800 93.700 ;
        RECT 271.600 89.700 274.000 90.300 ;
        RECT 271.600 88.800 272.400 89.700 ;
        RECT 273.200 82.200 274.000 89.700 ;
        RECT 277.800 90.200 278.400 93.600 ;
        RECT 279.400 93.000 280.000 94.600 ;
        RECT 279.000 92.200 280.000 93.000 ;
        RECT 279.400 90.200 280.000 92.200 ;
        RECT 281.000 92.400 281.800 93.200 ;
        RECT 281.000 92.300 282.000 92.400 ;
        RECT 282.800 92.300 283.600 92.400 ;
        RECT 281.000 91.700 283.600 92.300 ;
        RECT 281.000 91.600 282.000 91.700 ;
        RECT 282.800 91.600 283.600 91.700 ;
        RECT 277.800 89.200 278.800 90.200 ;
        RECT 279.400 89.600 282.000 90.200 ;
        RECT 278.000 82.200 278.800 89.200 ;
        RECT 281.200 82.200 282.000 89.600 ;
        RECT 282.800 88.800 283.600 90.400 ;
        RECT 284.400 88.300 285.200 95.800 ;
        RECT 286.000 93.600 286.800 95.200 ;
        RECT 292.600 94.400 293.200 95.800 ;
        RECT 294.200 95.400 297.800 95.800 ;
        RECT 296.400 94.400 297.200 94.800 ;
        RECT 292.400 93.600 295.000 94.400 ;
        RECT 296.400 94.300 298.000 94.400 ;
        RECT 298.800 94.300 299.600 95.200 ;
        RECT 296.400 93.800 299.600 94.300 ;
        RECT 297.200 93.700 299.600 93.800 ;
        RECT 297.200 93.600 298.000 93.700 ;
        RECT 298.800 93.600 299.600 93.700 ;
        RECT 300.400 94.300 301.200 95.800 ;
        RECT 303.600 95.600 304.400 97.200 ;
        RECT 302.000 94.300 302.800 94.400 ;
        RECT 300.400 93.700 302.800 94.300 ;
        RECT 292.400 90.200 293.200 90.400 ;
        RECT 294.400 90.200 295.000 93.600 ;
        RECT 295.600 91.600 296.400 93.200 ;
        RECT 292.400 89.600 293.800 90.200 ;
        RECT 294.400 89.600 295.400 90.200 ;
        RECT 293.200 88.400 293.800 89.600 ;
        RECT 290.800 88.300 291.600 88.400 ;
        RECT 284.400 87.700 291.600 88.300 ;
        RECT 284.400 82.200 285.200 87.700 ;
        RECT 290.800 87.600 291.600 87.700 ;
        RECT 293.200 87.600 294.000 88.400 ;
        RECT 294.600 82.200 295.400 89.600 ;
        RECT 300.400 82.200 301.200 93.700 ;
        RECT 302.000 93.600 302.800 93.700 ;
        RECT 302.000 90.300 302.800 90.400 ;
        RECT 305.200 90.300 306.000 99.800 ;
        RECT 309.400 96.400 310.200 99.800 ;
        RECT 308.400 95.800 310.200 96.400 ;
        RECT 306.800 93.600 307.600 95.200 ;
        RECT 302.000 89.700 306.000 90.300 ;
        RECT 302.000 88.800 302.800 89.700 ;
        RECT 305.200 82.200 306.000 89.700 ;
        RECT 308.400 82.200 309.200 95.800 ;
        RECT 311.600 95.000 312.400 99.800 ;
        RECT 316.000 98.400 316.800 99.800 ;
        RECT 314.800 97.800 316.800 98.400 ;
        RECT 320.400 97.800 321.200 99.800 ;
        RECT 324.600 98.400 325.800 99.800 ;
        RECT 324.400 97.800 325.800 98.400 ;
        RECT 314.800 97.000 315.600 97.800 ;
        RECT 320.400 97.200 321.000 97.800 ;
        RECT 316.400 96.400 317.200 97.200 ;
        RECT 318.200 96.600 321.000 97.200 ;
        RECT 324.400 97.000 325.200 97.800 ;
        RECT 318.200 96.400 319.000 96.600 ;
        RECT 312.400 94.200 314.000 94.400 ;
        RECT 316.600 94.200 317.200 96.400 ;
        RECT 326.200 95.400 327.000 95.600 ;
        RECT 329.200 95.400 330.000 99.800 ;
        RECT 326.200 94.800 330.000 95.400 ;
        RECT 330.800 95.000 331.600 99.800 ;
        RECT 335.200 98.400 336.000 99.800 ;
        RECT 334.000 97.800 336.000 98.400 ;
        RECT 339.600 97.800 340.400 99.800 ;
        RECT 343.800 98.400 345.000 99.800 ;
        RECT 343.600 97.800 345.000 98.400 ;
        RECT 334.000 97.000 334.800 97.800 ;
        RECT 339.600 97.200 340.200 97.800 ;
        RECT 335.600 96.400 336.400 97.200 ;
        RECT 337.400 96.600 340.200 97.200 ;
        RECT 343.600 97.000 344.400 97.800 ;
        RECT 337.400 96.400 338.200 96.600 ;
        RECT 322.200 94.200 323.000 94.400 ;
        RECT 312.400 93.600 323.400 94.200 ;
        RECT 315.400 93.400 316.200 93.600 ;
        RECT 313.800 92.400 314.600 92.600 ;
        RECT 316.400 92.400 317.200 92.600 ;
        RECT 322.800 92.400 323.400 93.600 ;
        RECT 324.400 92.800 325.200 93.000 ;
        RECT 313.800 91.800 318.800 92.400 ;
        RECT 318.000 91.600 318.800 91.800 ;
        RECT 322.800 91.600 323.600 92.400 ;
        RECT 324.400 92.200 328.200 92.800 ;
        RECT 327.400 92.000 328.200 92.200 ;
        RECT 311.600 91.000 317.200 91.200 ;
        RECT 311.600 90.800 317.400 91.000 ;
        RECT 311.600 90.600 321.400 90.800 ;
        RECT 310.000 88.800 310.800 90.400 ;
        RECT 311.600 82.200 312.400 90.600 ;
        RECT 316.600 90.200 321.400 90.600 ;
        RECT 314.800 89.000 320.200 89.600 ;
        RECT 314.800 88.800 315.600 89.000 ;
        RECT 319.400 88.800 320.200 89.000 ;
        RECT 320.800 89.000 321.400 90.200 ;
        RECT 322.800 90.400 323.400 91.600 ;
        RECT 325.800 91.400 326.600 91.600 ;
        RECT 329.200 91.400 330.000 94.800 ;
        RECT 331.600 94.200 333.200 94.400 ;
        RECT 335.800 94.200 336.400 96.400 ;
        RECT 345.400 95.400 346.200 95.600 ;
        RECT 348.400 95.400 349.200 99.800 ;
        RECT 345.400 94.800 349.200 95.400 ;
        RECT 341.400 94.200 342.200 94.400 ;
        RECT 331.600 93.600 342.600 94.200 ;
        RECT 334.600 93.400 335.400 93.600 ;
        RECT 333.000 92.400 333.800 92.600 ;
        RECT 335.600 92.400 336.400 92.600 ;
        RECT 342.000 92.400 342.600 93.600 ;
        RECT 343.600 92.800 344.400 93.000 ;
        RECT 333.000 91.800 338.000 92.400 ;
        RECT 337.200 91.600 338.000 91.800 ;
        RECT 342.000 91.600 342.800 92.400 ;
        RECT 343.600 92.200 347.400 92.800 ;
        RECT 346.600 92.000 347.400 92.200 ;
        RECT 325.800 90.800 330.000 91.400 ;
        RECT 322.800 89.800 325.200 90.400 ;
        RECT 322.200 89.000 323.000 89.200 ;
        RECT 320.800 88.400 323.000 89.000 ;
        RECT 324.600 88.800 325.200 89.800 ;
        RECT 324.600 88.000 326.000 88.800 ;
        RECT 318.200 87.400 319.000 87.600 ;
        RECT 321.000 87.400 321.800 87.600 ;
        RECT 314.800 86.200 315.600 87.000 ;
        RECT 318.200 86.800 321.800 87.400 ;
        RECT 320.400 86.200 321.000 86.800 ;
        RECT 324.400 86.200 325.200 87.000 ;
        RECT 314.800 85.600 316.800 86.200 ;
        RECT 316.000 82.200 316.800 85.600 ;
        RECT 320.400 82.200 321.200 86.200 ;
        RECT 324.600 82.200 325.800 86.200 ;
        RECT 329.200 82.200 330.000 90.800 ;
        RECT 330.800 91.000 336.400 91.200 ;
        RECT 330.800 90.800 336.600 91.000 ;
        RECT 330.800 90.600 340.600 90.800 ;
        RECT 330.800 82.200 331.600 90.600 ;
        RECT 335.800 90.200 340.600 90.600 ;
        RECT 334.000 89.000 339.400 89.600 ;
        RECT 334.000 88.800 334.800 89.000 ;
        RECT 338.600 88.800 339.400 89.000 ;
        RECT 340.000 89.000 340.600 90.200 ;
        RECT 342.000 90.400 342.600 91.600 ;
        RECT 345.000 91.400 345.800 91.600 ;
        RECT 348.400 91.400 349.200 94.800 ;
        RECT 350.000 95.200 350.800 99.800 ;
        RECT 353.200 96.400 354.000 99.800 ;
        RECT 358.000 97.800 358.800 99.800 ;
        RECT 353.200 95.800 354.200 96.400 ;
        RECT 350.000 94.600 352.600 95.200 ;
        RECT 350.200 92.400 351.000 93.200 ;
        RECT 350.000 91.600 351.000 92.400 ;
        RECT 352.000 93.000 352.600 94.600 ;
        RECT 353.600 94.400 354.200 95.800 ;
        RECT 356.400 95.600 357.200 97.200 ;
        RECT 358.200 95.600 358.800 97.800 ;
        RECT 361.200 95.800 362.000 99.800 ;
        RECT 363.400 96.400 364.200 99.800 ;
        RECT 363.400 95.800 365.200 96.400 ;
        RECT 358.200 95.000 360.600 95.600 ;
        RECT 353.200 94.300 354.200 94.400 ;
        RECT 358.000 94.300 359.000 94.400 ;
        RECT 353.200 93.700 359.000 94.300 ;
        RECT 353.200 93.600 354.200 93.700 ;
        RECT 358.000 93.600 359.000 93.700 ;
        RECT 352.000 92.200 353.000 93.000 ;
        RECT 345.000 90.800 349.200 91.400 ;
        RECT 342.000 89.800 344.400 90.400 ;
        RECT 341.400 89.000 342.200 89.200 ;
        RECT 340.000 88.400 342.200 89.000 ;
        RECT 343.800 88.800 344.400 89.800 ;
        RECT 343.800 88.400 345.200 88.800 ;
        RECT 343.800 88.000 346.000 88.400 ;
        RECT 344.600 87.600 346.000 88.000 ;
        RECT 337.400 87.400 338.200 87.600 ;
        RECT 340.200 87.400 341.000 87.600 ;
        RECT 334.000 86.200 334.800 87.000 ;
        RECT 337.400 86.800 341.000 87.400 ;
        RECT 339.600 86.200 340.200 86.800 ;
        RECT 343.600 86.200 344.400 87.000 ;
        RECT 334.000 85.600 336.000 86.200 ;
        RECT 335.200 82.200 336.000 85.600 ;
        RECT 339.600 82.200 340.400 86.200 ;
        RECT 343.800 82.200 345.000 86.200 ;
        RECT 348.400 82.200 349.200 90.800 ;
        RECT 352.000 90.200 352.600 92.200 ;
        RECT 353.600 90.200 354.200 93.600 ;
        RECT 358.400 92.800 359.200 93.600 ;
        RECT 360.000 92.000 360.600 95.000 ;
        RECT 361.400 92.400 362.000 95.800 ;
        RECT 359.800 91.400 360.600 92.000 ;
        RECT 361.200 91.600 362.000 92.400 ;
        RECT 350.000 89.600 352.600 90.200 ;
        RECT 350.000 82.200 350.800 89.600 ;
        RECT 353.200 89.200 354.200 90.200 ;
        RECT 356.400 91.200 360.600 91.400 ;
        RECT 356.400 90.800 360.400 91.200 ;
        RECT 353.200 82.200 354.000 89.200 ;
        RECT 356.400 82.200 357.200 90.800 ;
        RECT 361.400 90.300 362.000 91.600 ;
        RECT 364.400 92.300 365.200 95.800 ;
        RECT 367.600 95.800 368.400 99.800 ;
        RECT 372.000 98.400 373.600 99.800 ;
        RECT 372.000 97.600 374.800 98.400 ;
        RECT 372.000 96.200 373.600 97.600 ;
        RECT 367.600 95.200 370.000 95.800 ;
        RECT 366.000 93.600 366.800 95.200 ;
        RECT 369.200 95.000 370.000 95.200 ;
        RECT 370.600 94.800 371.400 95.600 ;
        RECT 370.600 94.400 371.200 94.800 ;
        RECT 367.600 93.600 369.200 94.400 ;
        RECT 370.400 93.600 371.200 94.400 ;
        RECT 372.000 94.200 372.600 96.200 ;
        RECT 377.200 95.800 378.000 99.800 ;
        RECT 380.400 97.800 381.200 99.800 ;
        RECT 373.200 94.800 374.800 95.600 ;
        RECT 375.400 95.200 378.000 95.800 ;
        RECT 378.800 95.600 379.600 97.200 ;
        RECT 375.400 95.000 376.200 95.200 ;
        RECT 380.600 94.400 381.200 97.800 ;
        RECT 383.600 96.000 384.400 99.800 ;
        RECT 386.800 96.000 387.600 99.800 ;
        RECT 383.600 95.800 387.600 96.000 ;
        RECT 388.400 95.800 389.200 99.800 ;
        RECT 393.200 95.800 394.000 99.800 ;
        RECT 394.600 96.400 395.400 97.200 ;
        RECT 383.800 95.400 387.400 95.800 ;
        RECT 384.400 94.400 385.200 94.800 ;
        RECT 388.400 94.400 389.000 95.800 ;
        RECT 376.400 94.200 378.000 94.400 ;
        RECT 372.000 93.600 373.000 94.200 ;
        RECT 375.800 94.000 378.000 94.200 ;
        RECT 367.700 92.400 368.300 93.600 ;
        RECT 372.400 92.400 373.000 93.600 ;
        RECT 373.600 93.600 378.000 94.000 ;
        RECT 380.400 93.600 381.200 94.400 ;
        RECT 383.600 93.800 385.200 94.400 ;
        RECT 386.600 94.300 389.200 94.400 ;
        RECT 390.000 94.300 390.800 94.400 ;
        RECT 383.600 93.600 384.400 93.800 ;
        RECT 386.600 93.700 390.800 94.300 ;
        RECT 386.600 93.600 389.200 93.700 ;
        RECT 390.000 93.600 390.800 93.700 ;
        RECT 373.600 93.400 376.400 93.600 ;
        RECT 373.600 93.200 374.400 93.400 ;
        RECT 367.600 92.300 368.400 92.400 ;
        RECT 364.400 91.700 368.400 92.300 ;
        RECT 362.800 90.300 363.600 90.400 ;
        RECT 361.300 90.200 363.600 90.300 ;
        RECT 360.600 89.700 363.600 90.200 ;
        RECT 360.600 89.600 362.000 89.700 ;
        RECT 360.600 82.200 361.400 89.600 ;
        RECT 362.800 88.800 363.600 89.700 ;
        RECT 364.400 82.200 365.200 91.700 ;
        RECT 367.600 91.600 368.400 91.700 ;
        RECT 372.400 91.600 373.200 92.400 ;
        RECT 375.000 92.200 375.800 92.400 ;
        RECT 374.200 91.600 375.800 92.200 ;
        RECT 372.400 90.200 373.000 91.600 ;
        RECT 374.200 91.400 375.000 91.600 ;
        RECT 380.600 90.200 381.200 93.600 ;
        RECT 382.000 90.800 382.800 92.400 ;
        RECT 385.200 91.600 386.000 93.200 ;
        RECT 386.600 90.200 387.200 93.600 ;
        RECT 391.600 92.800 392.400 94.400 ;
        RECT 390.000 92.200 390.800 92.400 ;
        RECT 393.200 92.200 393.800 95.800 ;
        RECT 394.800 95.600 395.600 96.400 ;
        RECT 396.400 95.800 397.200 99.800 ;
        RECT 400.600 96.800 401.400 99.800 ;
        RECT 400.600 95.800 402.000 96.800 ;
        RECT 402.800 96.000 403.600 99.800 ;
        RECT 406.000 96.000 406.800 99.800 ;
        RECT 402.800 95.800 406.800 96.000 ;
        RECT 407.600 95.800 408.400 99.800 ;
        RECT 409.800 98.400 410.600 99.800 ;
        RECT 409.800 97.600 411.600 98.400 ;
        RECT 409.800 96.400 410.600 97.600 ;
        RECT 409.800 95.800 411.600 96.400 ;
        RECT 396.600 95.600 397.200 95.800 ;
        RECT 396.600 95.200 398.400 95.600 ;
        RECT 396.600 95.000 400.800 95.200 ;
        RECT 397.800 94.600 400.800 95.000 ;
        RECT 400.000 94.400 400.800 94.600 ;
        RECT 396.400 92.800 397.200 94.400 ;
        RECT 398.400 93.800 399.200 94.000 ;
        RECT 398.200 93.200 399.200 93.800 ;
        RECT 398.200 92.400 398.800 93.200 ;
        RECT 394.800 92.200 395.600 92.400 ;
        RECT 390.000 91.600 391.600 92.200 ;
        RECT 393.200 91.600 395.600 92.200 ;
        RECT 398.000 91.600 398.800 92.400 ;
        RECT 390.800 91.200 391.600 91.600 ;
        RECT 388.400 90.200 389.200 90.400 ;
        RECT 394.800 90.200 395.400 91.600 ;
        RECT 400.000 91.000 400.600 94.400 ;
        RECT 401.400 92.400 402.000 95.800 ;
        RECT 403.000 95.400 406.600 95.800 ;
        RECT 403.600 94.400 404.400 94.800 ;
        RECT 407.600 94.400 408.200 95.800 ;
        RECT 402.800 93.800 404.400 94.400 ;
        RECT 402.800 93.600 403.600 93.800 ;
        RECT 405.800 93.600 408.400 94.400 ;
        RECT 401.200 92.300 402.000 92.400 ;
        RECT 404.400 92.300 405.200 93.200 ;
        RECT 401.200 91.700 405.200 92.300 ;
        RECT 401.200 91.600 402.000 91.700 ;
        RECT 404.400 91.600 405.200 91.700 ;
        RECT 398.200 90.400 400.600 91.000 ;
        RECT 367.600 89.600 370.000 90.200 ;
        RECT 367.600 82.200 368.400 89.600 ;
        RECT 369.200 89.400 370.000 89.600 ;
        RECT 372.000 82.200 373.600 90.200 ;
        RECT 375.400 89.600 378.000 90.200 ;
        RECT 375.400 89.400 376.200 89.600 ;
        RECT 377.200 82.200 378.000 89.600 ;
        RECT 380.400 89.400 382.200 90.200 ;
        RECT 381.400 88.400 382.200 89.400 ;
        RECT 386.200 89.600 387.200 90.200 ;
        RECT 387.800 89.600 389.200 90.200 ;
        RECT 390.000 89.600 394.000 90.200 ;
        RECT 381.400 87.600 382.800 88.400 ;
        RECT 381.400 82.200 382.200 87.600 ;
        RECT 386.200 82.200 387.000 89.600 ;
        RECT 387.800 88.400 388.400 89.600 ;
        RECT 387.600 87.600 388.400 88.400 ;
        RECT 390.000 82.200 390.800 89.600 ;
        RECT 393.200 82.200 394.000 89.600 ;
        RECT 394.800 82.200 395.600 90.200 ;
        RECT 398.200 86.200 398.800 90.400 ;
        RECT 401.400 90.200 402.000 91.600 ;
        RECT 405.800 90.200 406.400 93.600 ;
        RECT 407.600 90.200 408.400 90.400 ;
        RECT 398.000 82.200 398.800 86.200 ;
        RECT 401.200 82.200 402.000 90.200 ;
        RECT 405.400 89.600 406.400 90.200 ;
        RECT 407.000 89.600 408.400 90.200 ;
        RECT 405.400 82.200 406.200 89.600 ;
        RECT 407.000 88.400 407.600 89.600 ;
        RECT 409.200 88.800 410.000 90.400 ;
        RECT 406.800 87.600 407.600 88.400 ;
        RECT 410.800 82.200 411.600 95.800 ;
        RECT 412.400 94.300 413.200 95.200 ;
        RECT 414.000 94.300 414.800 99.800 ;
        RECT 417.200 95.200 418.000 99.800 ;
        RECT 418.800 95.800 419.600 99.800 ;
        RECT 420.400 96.000 421.200 99.800 ;
        RECT 423.600 96.000 424.400 99.800 ;
        RECT 420.400 95.800 424.400 96.000 ;
        RECT 425.200 95.800 426.000 99.800 ;
        RECT 426.800 96.000 427.600 99.800 ;
        RECT 430.000 96.000 430.800 99.800 ;
        RECT 426.800 95.800 430.800 96.000 ;
        RECT 412.400 93.700 414.800 94.300 ;
        RECT 412.400 93.600 413.200 93.700 ;
        RECT 414.000 92.400 414.800 93.700 ;
        RECT 415.800 94.600 418.000 95.200 ;
        RECT 414.000 90.200 414.600 92.400 ;
        RECT 415.800 91.600 416.400 94.600 ;
        RECT 419.000 94.400 419.600 95.800 ;
        RECT 420.600 95.400 424.200 95.800 ;
        RECT 422.800 94.400 423.600 94.800 ;
        RECT 425.400 94.400 426.000 95.800 ;
        RECT 427.000 95.400 430.600 95.800 ;
        RECT 431.600 95.000 432.400 99.800 ;
        RECT 436.000 98.400 436.800 99.800 ;
        RECT 434.800 97.800 436.800 98.400 ;
        RECT 440.400 97.800 441.200 99.800 ;
        RECT 444.600 98.400 445.800 99.800 ;
        RECT 444.400 97.800 445.800 98.400 ;
        RECT 449.200 98.300 450.000 99.800 ;
        RECT 450.800 98.300 451.600 98.400 ;
        RECT 434.800 97.000 435.600 97.800 ;
        RECT 440.400 97.200 441.000 97.800 ;
        RECT 436.400 96.400 437.200 97.200 ;
        RECT 438.200 96.600 441.000 97.200 ;
        RECT 444.400 97.000 445.200 97.800 ;
        RECT 449.200 97.700 451.600 98.300 ;
        RECT 438.200 96.400 439.000 96.600 ;
        RECT 429.200 94.400 430.000 94.800 ;
        RECT 418.800 93.600 421.400 94.400 ;
        RECT 422.800 93.800 424.400 94.400 ;
        RECT 423.600 93.600 424.400 93.800 ;
        RECT 425.200 93.600 427.800 94.400 ;
        RECT 429.200 93.800 430.800 94.400 ;
        RECT 430.000 93.600 430.800 93.800 ;
        RECT 432.400 94.200 434.000 94.400 ;
        RECT 436.600 94.200 437.200 96.400 ;
        RECT 446.200 95.400 447.000 95.600 ;
        RECT 449.200 95.400 450.000 97.700 ;
        RECT 450.800 97.600 451.600 97.700 ;
        RECT 446.200 94.800 450.000 95.400 ;
        RECT 455.600 95.800 456.400 99.800 ;
        RECT 460.000 98.400 461.600 99.800 ;
        RECT 460.000 97.600 462.800 98.400 ;
        RECT 460.000 96.200 461.600 97.600 ;
        RECT 455.600 95.200 458.000 95.800 ;
        RECT 457.200 95.000 458.000 95.200 ;
        RECT 442.200 94.200 443.000 94.400 ;
        RECT 432.400 93.600 443.400 94.200 ;
        RECT 417.200 91.600 418.000 93.200 ;
        RECT 415.200 90.800 416.400 91.600 ;
        RECT 415.800 90.200 416.400 90.800 ;
        RECT 420.800 90.400 421.400 93.600 ;
        RECT 422.000 91.600 422.800 93.200 ;
        RECT 418.800 90.200 419.600 90.400 ;
        RECT 414.000 82.200 414.800 90.200 ;
        RECT 415.800 89.600 418.000 90.200 ;
        RECT 418.800 89.600 420.200 90.200 ;
        RECT 420.800 89.600 422.800 90.400 ;
        RECT 425.200 90.200 426.000 90.400 ;
        RECT 427.200 90.200 427.800 93.600 ;
        RECT 435.400 93.400 436.200 93.600 ;
        RECT 428.400 91.600 429.200 93.200 ;
        RECT 433.800 92.400 434.600 92.600 ;
        RECT 436.400 92.400 437.200 92.600 ;
        RECT 433.800 91.800 438.800 92.400 ;
        RECT 438.000 91.600 438.800 91.800 ;
        RECT 431.600 91.000 437.200 91.200 ;
        RECT 431.600 90.800 437.400 91.000 ;
        RECT 431.600 90.600 441.400 90.800 ;
        RECT 425.200 89.600 426.600 90.200 ;
        RECT 427.200 89.600 428.200 90.200 ;
        RECT 417.200 82.200 418.000 89.600 ;
        RECT 419.600 88.400 420.200 89.600 ;
        RECT 419.600 87.600 420.400 88.400 ;
        RECT 421.000 82.200 421.800 89.600 ;
        RECT 426.000 88.400 426.600 89.600 ;
        RECT 426.000 87.600 426.800 88.400 ;
        RECT 427.400 82.200 428.200 89.600 ;
        RECT 431.600 82.200 432.400 90.600 ;
        RECT 436.600 90.200 441.400 90.600 ;
        RECT 434.800 89.000 440.200 89.600 ;
        RECT 434.800 88.800 435.600 89.000 ;
        RECT 439.400 88.800 440.200 89.000 ;
        RECT 440.800 89.000 441.400 90.200 ;
        RECT 442.800 90.400 443.400 93.600 ;
        RECT 444.400 92.800 445.200 93.000 ;
        RECT 444.400 92.200 448.200 92.800 ;
        RECT 447.400 92.000 448.200 92.200 ;
        RECT 445.800 91.400 446.600 91.600 ;
        RECT 449.200 91.400 450.000 94.800 ;
        RECT 458.600 94.800 459.400 95.600 ;
        RECT 458.600 94.400 459.200 94.800 ;
        RECT 452.400 94.300 453.200 94.400 ;
        RECT 455.600 94.300 457.200 94.400 ;
        RECT 452.400 93.700 457.200 94.300 ;
        RECT 452.400 93.600 453.200 93.700 ;
        RECT 455.600 93.600 457.200 93.700 ;
        RECT 458.400 93.600 459.200 94.400 ;
        RECT 460.000 92.800 460.600 96.200 ;
        RECT 465.200 95.800 466.000 99.800 ;
        RECT 461.200 95.400 462.800 95.600 ;
        RECT 461.200 94.800 463.200 95.400 ;
        RECT 463.800 95.200 466.000 95.800 ;
        RECT 466.800 95.800 467.600 99.800 ;
        RECT 471.200 96.200 472.800 99.800 ;
        RECT 466.800 95.200 469.000 95.800 ;
        RECT 470.000 95.400 471.600 95.600 ;
        RECT 463.800 95.000 464.600 95.200 ;
        RECT 468.200 95.000 469.000 95.200 ;
        RECT 462.600 94.400 463.200 94.800 ;
        RECT 469.600 94.800 471.600 95.400 ;
        RECT 469.600 94.400 470.200 94.800 ;
        RECT 461.200 93.400 462.000 94.200 ;
        RECT 462.600 93.800 466.000 94.400 ;
        RECT 464.400 93.600 466.000 93.800 ;
        RECT 466.800 93.800 470.200 94.400 ;
        RECT 466.800 93.600 468.400 93.800 ;
        RECT 459.600 92.400 460.600 92.800 ;
        RECT 458.800 92.200 460.600 92.400 ;
        RECT 461.400 92.800 462.000 93.400 ;
        RECT 470.800 93.400 471.600 94.200 ;
        RECT 470.800 92.800 471.400 93.400 ;
        RECT 461.400 92.200 464.000 92.800 ;
        RECT 458.800 91.600 460.200 92.200 ;
        RECT 463.200 92.000 464.000 92.200 ;
        RECT 468.800 92.200 471.400 92.800 ;
        RECT 472.200 92.800 472.800 96.200 ;
        RECT 476.400 95.800 477.200 99.800 ;
        RECT 473.400 94.800 474.200 95.600 ;
        RECT 474.800 95.200 477.200 95.800 ;
        RECT 478.000 95.600 478.800 97.200 ;
        RECT 474.800 95.000 475.600 95.200 ;
        RECT 473.600 94.400 474.200 94.800 ;
        RECT 473.600 93.600 474.400 94.400 ;
        RECT 475.600 93.600 477.200 94.400 ;
        RECT 472.200 92.400 473.200 92.800 ;
        RECT 472.200 92.300 474.000 92.400 ;
        RECT 478.000 92.300 478.800 92.400 ;
        RECT 472.200 92.200 478.800 92.300 ;
        RECT 468.800 92.000 469.600 92.200 ;
        RECT 472.600 91.700 478.800 92.200 ;
        RECT 472.600 91.600 474.000 91.700 ;
        RECT 478.000 91.600 478.800 91.700 ;
        RECT 445.800 90.800 450.000 91.400 ;
        RECT 442.800 89.800 445.200 90.400 ;
        RECT 442.200 89.000 443.000 89.200 ;
        RECT 440.800 88.400 443.000 89.000 ;
        RECT 444.600 88.800 445.200 89.800 ;
        RECT 444.600 88.000 446.000 88.800 ;
        RECT 438.200 87.400 439.000 87.600 ;
        RECT 441.000 87.400 441.800 87.600 ;
        RECT 434.800 86.200 435.600 87.000 ;
        RECT 438.200 86.800 441.800 87.400 ;
        RECT 440.400 86.200 441.000 86.800 ;
        RECT 444.400 86.200 445.200 87.000 ;
        RECT 434.800 85.600 436.800 86.200 ;
        RECT 436.000 82.200 436.800 85.600 ;
        RECT 440.400 82.200 441.200 86.200 ;
        RECT 444.600 82.200 445.800 86.200 ;
        RECT 449.200 82.200 450.000 90.800 ;
        RECT 459.600 90.200 460.200 91.600 ;
        RECT 461.000 91.400 461.800 91.600 ;
        RECT 471.000 91.400 471.800 91.600 ;
        RECT 461.000 90.800 464.400 91.400 ;
        RECT 463.800 90.200 464.400 90.800 ;
        RECT 468.400 90.800 471.800 91.400 ;
        RECT 468.400 90.200 469.000 90.800 ;
        RECT 472.600 90.200 473.200 91.600 ;
        RECT 479.600 90.300 480.400 99.800 ;
        RECT 484.800 94.300 485.600 99.800 ;
        RECT 490.200 98.400 491.000 99.800 ;
        RECT 490.200 97.600 491.600 98.400 ;
        RECT 490.200 96.400 491.000 97.600 ;
        RECT 489.200 95.800 491.000 96.400 ;
        RECT 487.600 94.300 488.400 95.200 ;
        RECT 484.800 93.800 488.400 94.300 ;
        RECT 485.000 93.700 488.400 93.800 ;
        RECT 485.000 93.600 486.600 93.700 ;
        RECT 487.600 93.600 488.400 93.700 ;
        RECT 482.800 91.600 484.400 92.400 ;
        RECT 481.200 90.300 482.000 91.200 ;
        RECT 455.600 89.600 458.000 90.200 ;
        RECT 459.600 89.600 461.600 90.200 ;
        RECT 455.600 82.200 456.400 89.600 ;
        RECT 457.200 89.400 458.000 89.600 ;
        RECT 460.000 82.200 461.600 89.600 ;
        RECT 463.800 89.600 466.000 90.200 ;
        RECT 463.800 89.400 464.600 89.600 ;
        RECT 465.200 82.200 466.000 89.600 ;
        RECT 466.800 89.600 469.000 90.200 ;
        RECT 466.800 82.200 467.600 89.600 ;
        RECT 468.200 89.400 469.000 89.600 ;
        RECT 471.200 89.600 473.200 90.200 ;
        RECT 474.800 89.600 477.200 90.200 ;
        RECT 471.200 82.200 472.800 89.600 ;
        RECT 474.800 89.400 475.600 89.600 ;
        RECT 476.400 82.200 477.200 89.600 ;
        RECT 479.600 89.700 482.000 90.300 ;
        RECT 479.600 82.200 480.400 89.700 ;
        RECT 481.200 89.600 482.000 89.700 ;
        RECT 486.000 90.400 486.600 93.600 ;
        RECT 486.000 89.600 486.800 90.400 ;
        RECT 484.400 87.600 485.200 89.200 ;
        RECT 486.000 87.000 486.600 89.600 ;
        RECT 483.000 86.400 486.600 87.000 ;
        RECT 483.000 86.200 483.600 86.400 ;
        RECT 482.800 82.200 483.600 86.200 ;
        RECT 486.000 86.200 486.600 86.400 ;
        RECT 486.000 82.200 486.800 86.200 ;
        RECT 489.200 82.200 490.000 95.800 ;
        RECT 492.400 95.000 493.200 99.800 ;
        RECT 496.800 98.400 497.600 99.800 ;
        RECT 495.600 97.800 497.600 98.400 ;
        RECT 501.200 97.800 502.000 99.800 ;
        RECT 505.400 98.400 506.600 99.800 ;
        RECT 505.200 97.800 506.600 98.400 ;
        RECT 495.600 97.000 496.400 97.800 ;
        RECT 501.200 97.200 501.800 97.800 ;
        RECT 497.200 96.400 498.000 97.200 ;
        RECT 499.000 96.600 501.800 97.200 ;
        RECT 505.200 97.000 506.000 97.800 ;
        RECT 499.000 96.400 499.800 96.600 ;
        RECT 493.200 94.200 494.800 94.400 ;
        RECT 497.400 94.200 498.000 96.400 ;
        RECT 507.000 95.400 507.800 95.600 ;
        RECT 510.000 95.400 510.800 99.800 ;
        RECT 507.000 94.800 510.800 95.400 ;
        RECT 503.000 94.200 503.800 94.400 ;
        RECT 493.200 93.600 504.200 94.200 ;
        RECT 496.200 93.400 497.000 93.600 ;
        RECT 494.600 92.400 495.400 92.600 ;
        RECT 497.200 92.400 498.000 92.600 ;
        RECT 503.600 92.400 504.200 93.600 ;
        RECT 505.200 92.800 506.000 93.000 ;
        RECT 494.600 91.800 499.600 92.400 ;
        RECT 498.800 91.600 499.600 91.800 ;
        RECT 503.600 91.600 504.400 92.400 ;
        RECT 505.200 92.200 509.000 92.800 ;
        RECT 508.200 92.000 509.000 92.200 ;
        RECT 492.400 91.000 498.000 91.200 ;
        RECT 492.400 90.800 498.200 91.000 ;
        RECT 492.400 90.600 502.200 90.800 ;
        RECT 490.800 88.800 491.600 90.400 ;
        RECT 492.400 82.200 493.200 90.600 ;
        RECT 497.400 90.200 502.200 90.600 ;
        RECT 495.600 89.000 501.000 89.600 ;
        RECT 495.600 88.800 496.400 89.000 ;
        RECT 500.200 88.800 501.000 89.000 ;
        RECT 501.600 89.000 502.200 90.200 ;
        RECT 503.600 90.400 504.200 91.600 ;
        RECT 506.600 91.400 507.400 91.600 ;
        RECT 510.000 91.400 510.800 94.800 ;
        RECT 506.600 90.800 510.800 91.400 ;
        RECT 503.600 89.800 506.000 90.400 ;
        RECT 503.000 89.000 503.800 89.200 ;
        RECT 501.600 88.400 503.800 89.000 ;
        RECT 505.400 88.800 506.000 89.800 ;
        RECT 505.400 88.000 506.800 88.800 ;
        RECT 499.000 87.400 499.800 87.600 ;
        RECT 501.800 87.400 502.600 87.600 ;
        RECT 495.600 86.200 496.400 87.000 ;
        RECT 499.000 86.800 502.600 87.400 ;
        RECT 501.200 86.200 501.800 86.800 ;
        RECT 505.200 86.200 506.000 87.000 ;
        RECT 495.600 85.600 497.600 86.200 ;
        RECT 496.800 82.200 497.600 85.600 ;
        RECT 501.200 82.200 502.000 86.200 ;
        RECT 505.400 82.200 506.600 86.200 ;
        RECT 510.000 82.200 510.800 90.800 ;
        RECT 511.600 95.400 512.400 99.800 ;
        RECT 515.800 98.400 517.000 99.800 ;
        RECT 515.800 97.800 517.200 98.400 ;
        RECT 520.400 97.800 521.200 99.800 ;
        RECT 524.800 98.400 525.600 99.800 ;
        RECT 524.800 97.800 526.800 98.400 ;
        RECT 516.400 97.000 517.200 97.800 ;
        RECT 520.600 97.200 521.200 97.800 ;
        RECT 520.600 96.600 523.400 97.200 ;
        RECT 522.600 96.400 523.400 96.600 ;
        RECT 524.400 96.400 525.200 97.200 ;
        RECT 526.000 97.000 526.800 97.800 ;
        RECT 514.600 95.400 515.400 95.600 ;
        RECT 511.600 94.800 515.400 95.400 ;
        RECT 511.600 91.400 512.400 94.800 ;
        RECT 518.600 94.200 519.400 94.400 ;
        RECT 524.400 94.200 525.000 96.400 ;
        RECT 529.200 95.000 530.000 99.800 ;
        RECT 530.800 95.000 531.600 99.800 ;
        RECT 535.200 98.400 536.000 99.800 ;
        RECT 534.000 97.800 536.000 98.400 ;
        RECT 539.600 97.800 540.400 99.800 ;
        RECT 543.800 98.400 545.000 99.800 ;
        RECT 543.600 97.800 545.000 98.400 ;
        RECT 534.000 97.000 534.800 97.800 ;
        RECT 539.600 97.200 540.200 97.800 ;
        RECT 535.600 96.400 536.400 97.200 ;
        RECT 537.400 96.600 540.200 97.200 ;
        RECT 543.600 97.000 544.400 97.800 ;
        RECT 537.400 96.400 538.200 96.600 ;
        RECT 527.600 94.300 529.200 94.400 ;
        RECT 531.600 94.300 533.200 94.400 ;
        RECT 527.600 94.200 533.200 94.300 ;
        RECT 535.800 94.200 536.400 96.400 ;
        RECT 545.400 95.400 546.200 95.600 ;
        RECT 548.400 95.400 549.200 99.800 ;
        RECT 545.400 94.800 549.200 95.400 ;
        RECT 541.400 94.200 542.800 94.400 ;
        RECT 518.200 93.700 542.800 94.200 ;
        RECT 518.200 93.600 529.200 93.700 ;
        RECT 531.600 93.600 542.800 93.700 ;
        RECT 516.400 92.800 517.200 93.000 ;
        RECT 513.400 92.200 517.200 92.800 ;
        RECT 518.200 92.400 518.800 93.600 ;
        RECT 525.400 93.400 526.200 93.600 ;
        RECT 534.600 93.400 535.400 93.600 ;
        RECT 524.400 92.400 525.200 92.600 ;
        RECT 527.000 92.400 527.800 92.600 ;
        RECT 513.400 92.000 514.200 92.200 ;
        RECT 518.000 91.600 518.800 92.400 ;
        RECT 522.800 91.800 527.800 92.400 ;
        RECT 533.000 92.400 533.800 92.600 ;
        RECT 533.000 91.800 538.000 92.400 ;
        RECT 522.800 91.600 523.600 91.800 ;
        RECT 537.200 91.600 538.000 91.800 ;
        RECT 515.000 91.400 515.800 91.600 ;
        RECT 511.600 90.800 515.800 91.400 ;
        RECT 511.600 82.200 512.400 90.800 ;
        RECT 518.200 90.400 518.800 91.600 ;
        RECT 524.400 91.000 530.000 91.200 ;
        RECT 524.200 90.800 530.000 91.000 ;
        RECT 516.400 89.800 518.800 90.400 ;
        RECT 520.200 90.600 530.000 90.800 ;
        RECT 520.200 90.200 525.000 90.600 ;
        RECT 516.400 88.800 517.000 89.800 ;
        RECT 515.600 88.000 517.000 88.800 ;
        RECT 518.600 89.000 519.400 89.200 ;
        RECT 520.200 89.000 520.800 90.200 ;
        RECT 518.600 88.400 520.800 89.000 ;
        RECT 521.400 89.000 526.800 89.600 ;
        RECT 521.400 88.800 522.200 89.000 ;
        RECT 526.000 88.800 526.800 89.000 ;
        RECT 519.800 87.400 520.600 87.600 ;
        RECT 522.600 87.400 523.400 87.600 ;
        RECT 516.400 86.200 517.200 87.000 ;
        RECT 519.800 86.800 523.400 87.400 ;
        RECT 520.600 86.200 521.200 86.800 ;
        RECT 526.000 86.200 526.800 87.000 ;
        RECT 515.800 82.200 517.000 86.200 ;
        RECT 520.400 82.200 521.200 86.200 ;
        RECT 524.800 85.600 526.800 86.200 ;
        RECT 524.800 82.200 525.600 85.600 ;
        RECT 529.200 82.200 530.000 90.600 ;
        RECT 530.800 91.000 536.400 91.200 ;
        RECT 530.800 90.800 536.600 91.000 ;
        RECT 530.800 90.600 540.600 90.800 ;
        RECT 530.800 82.200 531.600 90.600 ;
        RECT 535.800 90.200 540.600 90.600 ;
        RECT 534.000 89.000 539.400 89.600 ;
        RECT 534.000 88.800 534.800 89.000 ;
        RECT 538.600 88.800 539.400 89.000 ;
        RECT 540.000 89.000 540.600 90.200 ;
        RECT 542.000 90.400 542.600 93.600 ;
        RECT 543.600 92.800 544.400 93.000 ;
        RECT 543.600 92.200 547.400 92.800 ;
        RECT 546.600 92.000 547.400 92.200 ;
        RECT 545.000 91.400 545.800 91.600 ;
        RECT 548.400 91.400 549.200 94.800 ;
        RECT 545.000 90.800 549.200 91.400 ;
        RECT 542.000 89.800 544.400 90.400 ;
        RECT 541.400 89.000 542.200 89.200 ;
        RECT 540.000 88.400 542.200 89.000 ;
        RECT 543.800 88.800 544.400 89.800 ;
        RECT 543.800 88.000 545.200 88.800 ;
        RECT 537.400 87.400 538.200 87.600 ;
        RECT 540.200 87.400 541.000 87.600 ;
        RECT 534.000 86.200 534.800 87.000 ;
        RECT 537.400 86.800 541.000 87.400 ;
        RECT 539.600 86.200 540.200 86.800 ;
        RECT 543.600 86.200 544.400 87.000 ;
        RECT 534.000 85.600 536.000 86.200 ;
        RECT 535.200 82.200 536.000 85.600 ;
        RECT 539.600 82.200 540.400 86.200 ;
        RECT 543.800 82.200 545.000 86.200 ;
        RECT 548.400 82.200 549.200 90.800 ;
        RECT 550.000 82.200 550.800 99.800 ;
        RECT 551.600 93.600 552.400 95.200 ;
        RECT 553.200 95.000 554.000 99.800 ;
        RECT 557.600 98.400 558.400 99.800 ;
        RECT 556.400 97.800 558.400 98.400 ;
        RECT 562.000 97.800 562.800 99.800 ;
        RECT 566.200 98.400 567.400 99.800 ;
        RECT 566.000 97.800 567.400 98.400 ;
        RECT 556.400 97.000 557.200 97.800 ;
        RECT 562.000 97.200 562.600 97.800 ;
        RECT 558.000 96.400 558.800 97.200 ;
        RECT 559.800 96.600 562.600 97.200 ;
        RECT 566.000 97.000 566.800 97.800 ;
        RECT 559.800 96.400 560.600 96.600 ;
        RECT 554.000 94.200 555.600 94.400 ;
        RECT 558.200 94.200 558.800 96.400 ;
        RECT 567.800 95.400 568.600 95.600 ;
        RECT 570.800 95.400 571.600 99.800 ;
        RECT 567.800 94.800 571.600 95.400 ;
        RECT 563.800 94.200 564.600 94.400 ;
        RECT 554.000 93.600 565.000 94.200 ;
        RECT 557.000 93.400 557.800 93.600 ;
        RECT 555.400 92.400 556.200 92.600 ;
        RECT 558.000 92.400 558.800 92.600 ;
        RECT 555.400 91.800 560.400 92.400 ;
        RECT 559.600 91.600 560.400 91.800 ;
        RECT 553.200 91.000 558.800 91.200 ;
        RECT 553.200 90.800 559.000 91.000 ;
        RECT 553.200 90.600 563.000 90.800 ;
        RECT 553.200 82.200 554.000 90.600 ;
        RECT 558.200 90.200 563.000 90.600 ;
        RECT 556.400 89.000 561.800 89.600 ;
        RECT 556.400 88.800 557.200 89.000 ;
        RECT 561.000 88.800 561.800 89.000 ;
        RECT 562.400 89.000 563.000 90.200 ;
        RECT 564.400 90.400 565.000 93.600 ;
        RECT 566.000 92.800 566.800 93.000 ;
        RECT 566.000 92.200 569.800 92.800 ;
        RECT 569.000 92.000 569.800 92.200 ;
        RECT 567.400 91.400 568.200 91.600 ;
        RECT 570.800 91.400 571.600 94.800 ;
        RECT 572.400 95.200 573.200 99.800 ;
        RECT 577.200 95.200 578.000 99.800 ;
        RECT 572.400 94.600 574.600 95.200 ;
        RECT 577.200 94.600 579.400 95.200 ;
        RECT 572.400 91.600 573.200 93.200 ;
        RECT 574.000 91.600 574.600 94.600 ;
        RECT 577.200 91.600 578.000 93.200 ;
        RECT 578.800 91.600 579.400 94.600 ;
        RECT 567.400 90.800 571.600 91.400 ;
        RECT 564.400 89.800 566.800 90.400 ;
        RECT 563.800 89.000 564.600 89.200 ;
        RECT 562.400 88.400 564.600 89.000 ;
        RECT 566.200 88.800 566.800 89.800 ;
        RECT 566.200 88.400 567.600 88.800 ;
        RECT 566.200 88.000 568.400 88.400 ;
        RECT 567.000 87.600 568.400 88.000 ;
        RECT 559.800 87.400 560.600 87.600 ;
        RECT 562.600 87.400 563.400 87.600 ;
        RECT 556.400 86.200 557.200 87.000 ;
        RECT 559.800 86.800 563.400 87.400 ;
        RECT 562.000 86.200 562.600 86.800 ;
        RECT 566.000 86.200 566.800 87.000 ;
        RECT 556.400 85.600 558.400 86.200 ;
        RECT 557.600 82.200 558.400 85.600 ;
        RECT 562.000 82.200 562.800 86.200 ;
        RECT 566.200 82.200 567.400 86.200 ;
        RECT 570.800 82.200 571.600 90.800 ;
        RECT 574.000 90.800 575.200 91.600 ;
        RECT 578.800 90.800 580.000 91.600 ;
        RECT 574.000 90.200 574.600 90.800 ;
        RECT 578.800 90.200 579.400 90.800 ;
        RECT 572.400 89.600 574.600 90.200 ;
        RECT 577.200 89.600 579.400 90.200 ;
        RECT 572.400 82.200 573.200 89.600 ;
        RECT 577.200 82.200 578.000 89.600 ;
        RECT 1.200 72.400 2.000 79.800 ;
        RECT 2.600 72.400 3.400 72.600 ;
        RECT 1.200 71.800 3.400 72.400 ;
        RECT 5.600 72.400 7.200 79.800 ;
        RECT 9.200 72.400 10.000 72.600 ;
        RECT 10.800 72.400 11.600 79.800 ;
        RECT 5.600 71.800 7.600 72.400 ;
        RECT 9.200 71.800 11.600 72.400 ;
        RECT 2.800 71.200 3.400 71.800 ;
        RECT 2.800 70.600 6.200 71.200 ;
        RECT 5.400 70.400 6.200 70.600 ;
        RECT 7.000 70.400 7.600 71.800 ;
        RECT 12.400 71.600 13.200 73.200 ;
        RECT 3.200 69.800 4.000 70.000 ;
        RECT 7.000 69.800 8.400 70.400 ;
        RECT 3.200 69.200 5.800 69.800 ;
        RECT 5.200 68.600 5.800 69.200 ;
        RECT 6.600 69.600 8.400 69.800 ;
        RECT 6.600 69.200 7.600 69.600 ;
        RECT 1.200 68.200 2.800 68.400 ;
        RECT 1.200 67.600 4.600 68.200 ;
        RECT 5.200 67.800 6.000 68.600 ;
        RECT 4.000 67.200 4.600 67.600 ;
        RECT 2.600 66.800 3.400 67.000 ;
        RECT 1.200 66.200 3.400 66.800 ;
        RECT 4.000 66.600 6.000 67.200 ;
        RECT 4.400 66.400 6.000 66.600 ;
        RECT 1.200 62.200 2.000 66.200 ;
        RECT 6.600 65.800 7.200 69.200 ;
        RECT 8.000 67.600 8.800 68.400 ;
        RECT 10.000 68.300 11.600 68.400 ;
        RECT 12.400 68.300 13.200 68.400 ;
        RECT 10.000 67.700 13.200 68.300 ;
        RECT 10.000 67.600 11.600 67.700 ;
        RECT 12.400 67.600 13.200 67.700 ;
        RECT 8.000 67.200 8.600 67.600 ;
        RECT 7.800 66.400 8.600 67.200 ;
        RECT 9.200 66.800 10.000 67.000 ;
        RECT 9.200 66.200 11.600 66.800 ;
        RECT 14.000 66.200 14.800 79.800 ;
        RECT 19.800 72.400 20.600 79.800 ;
        RECT 21.200 73.600 22.000 74.400 ;
        RECT 21.400 72.400 22.000 73.600 ;
        RECT 19.800 71.800 20.800 72.400 ;
        RECT 21.400 71.800 22.800 72.400 ;
        RECT 18.800 68.800 19.600 70.400 ;
        RECT 20.200 68.400 20.800 71.800 ;
        RECT 22.000 71.600 22.800 71.800 ;
        RECT 15.600 66.800 16.400 68.400 ;
        RECT 17.200 68.200 18.000 68.400 ;
        RECT 20.200 68.300 22.800 68.400 ;
        RECT 23.600 68.300 24.400 68.400 ;
        RECT 17.200 67.600 18.800 68.200 ;
        RECT 20.200 67.700 24.400 68.300 ;
        RECT 20.200 67.600 22.800 67.700 ;
        RECT 18.000 67.200 18.800 67.600 ;
        RECT 17.400 66.200 21.000 66.600 ;
        RECT 22.000 66.200 22.600 67.600 ;
        RECT 23.600 66.800 24.400 67.700 ;
        RECT 25.200 66.200 26.000 79.800 ;
        RECT 29.200 73.600 30.000 74.400 ;
        RECT 26.800 71.600 27.600 73.200 ;
        RECT 29.200 72.400 29.800 73.600 ;
        RECT 30.600 72.400 31.400 79.800 ;
        RECT 28.400 71.800 29.800 72.400 ;
        RECT 28.400 71.600 29.200 71.800 ;
        RECT 30.400 71.600 32.400 72.400 ;
        RECT 30.400 68.400 31.000 71.600 ;
        RECT 31.600 68.800 32.400 70.400 ;
        RECT 28.400 67.600 31.000 68.400 ;
        RECT 33.200 68.200 34.000 68.400 ;
        RECT 32.400 67.600 34.000 68.200 ;
        RECT 28.600 66.200 29.200 67.600 ;
        RECT 32.400 67.200 33.200 67.600 ;
        RECT 30.200 66.200 33.800 66.600 ;
        RECT 5.600 64.400 7.200 65.800 ;
        RECT 4.400 63.600 7.200 64.400 ;
        RECT 5.600 62.200 7.200 63.600 ;
        RECT 10.800 62.200 11.600 66.200 ;
        RECT 13.000 65.600 14.800 66.200 ;
        RECT 17.200 66.000 21.200 66.200 ;
        RECT 13.000 64.400 13.800 65.600 ;
        RECT 12.400 63.600 13.800 64.400 ;
        RECT 13.000 62.200 13.800 63.600 ;
        RECT 17.200 62.200 18.000 66.000 ;
        RECT 20.400 62.200 21.200 66.000 ;
        RECT 22.000 62.200 22.800 66.200 ;
        RECT 25.200 65.600 27.000 66.200 ;
        RECT 26.200 64.400 27.000 65.600 ;
        RECT 26.200 63.600 27.600 64.400 ;
        RECT 26.200 62.200 27.000 63.600 ;
        RECT 28.400 62.200 29.200 66.200 ;
        RECT 30.000 66.000 34.000 66.200 ;
        RECT 30.000 62.200 30.800 66.000 ;
        RECT 33.200 62.200 34.000 66.000 ;
        RECT 34.800 62.200 35.600 79.800 ;
        RECT 40.600 72.600 41.400 79.800 ;
        RECT 39.600 71.800 41.400 72.600 ;
        RECT 45.400 72.400 46.200 79.800 ;
        RECT 46.800 73.600 47.600 74.400 ;
        RECT 47.000 72.400 47.600 73.600 ;
        RECT 45.400 71.800 46.400 72.400 ;
        RECT 47.000 72.300 48.400 72.400 ;
        RECT 49.200 72.300 50.000 79.800 ;
        RECT 47.000 71.800 50.000 72.300 ;
        RECT 53.000 72.600 53.800 79.800 ;
        RECT 57.800 72.600 58.600 79.800 ;
        RECT 53.000 71.800 54.800 72.600 ;
        RECT 57.800 71.800 59.600 72.600 ;
        RECT 64.600 72.400 65.400 79.800 ;
        RECT 66.000 73.600 66.800 74.400 ;
        RECT 66.200 72.400 66.800 73.600 ;
        RECT 39.800 68.400 40.400 71.800 ;
        RECT 41.200 69.600 42.000 71.200 ;
        RECT 44.400 68.800 45.200 70.400 ;
        RECT 45.800 68.400 46.400 71.800 ;
        RECT 47.600 71.700 50.000 71.800 ;
        RECT 47.600 71.600 48.400 71.700 ;
        RECT 36.400 66.800 37.200 68.400 ;
        RECT 39.600 68.300 40.400 68.400 ;
        RECT 42.800 68.300 43.600 68.400 ;
        RECT 39.600 68.200 43.600 68.300 ;
        RECT 39.600 67.700 44.400 68.200 ;
        RECT 39.600 67.600 40.400 67.700 ;
        RECT 42.800 67.600 44.400 67.700 ;
        RECT 45.800 67.600 48.400 68.400 ;
        RECT 38.000 64.800 38.800 66.400 ;
        RECT 39.800 64.200 40.400 67.600 ;
        RECT 43.600 67.200 44.400 67.600 ;
        RECT 43.000 66.200 46.600 66.600 ;
        RECT 47.600 66.200 48.200 67.600 ;
        RECT 39.600 62.200 40.400 64.200 ;
        RECT 42.800 66.000 46.800 66.200 ;
        RECT 42.800 62.200 43.600 66.000 ;
        RECT 46.000 62.200 46.800 66.000 ;
        RECT 47.600 62.200 48.400 66.200 ;
        RECT 49.200 62.200 50.000 71.700 ;
        RECT 50.800 70.300 51.600 70.400 ;
        RECT 52.400 70.300 53.200 71.200 ;
        RECT 50.800 69.700 53.200 70.300 ;
        RECT 50.800 69.600 51.600 69.700 ;
        RECT 52.400 69.600 53.200 69.700 ;
        RECT 54.000 68.400 54.600 71.800 ;
        RECT 55.600 70.300 56.400 70.400 ;
        RECT 57.200 70.300 58.000 71.200 ;
        RECT 55.600 69.700 58.000 70.300 ;
        RECT 55.600 69.600 56.400 69.700 ;
        RECT 57.200 69.600 58.000 69.700 ;
        RECT 58.800 68.400 59.400 71.800 ;
        RECT 63.600 71.600 65.600 72.400 ;
        RECT 66.200 71.800 67.600 72.400 ;
        RECT 66.800 71.600 67.600 71.800 ;
        RECT 62.000 70.300 62.800 70.400 ;
        RECT 63.600 70.300 64.400 70.400 ;
        RECT 62.000 69.700 64.400 70.300 ;
        RECT 62.000 69.600 62.800 69.700 ;
        RECT 63.600 68.800 64.400 69.700 ;
        RECT 65.000 68.400 65.600 71.600 ;
        RECT 70.000 71.200 70.800 79.800 ;
        RECT 73.200 71.200 74.000 79.800 ;
        RECT 70.000 70.400 74.000 71.200 ;
        RECT 54.000 68.300 54.800 68.400 ;
        RECT 57.200 68.300 58.000 68.400 ;
        RECT 54.000 67.700 58.000 68.300 ;
        RECT 54.000 67.600 54.800 67.700 ;
        RECT 57.200 67.600 58.000 67.700 ;
        RECT 58.800 67.600 59.600 68.400 ;
        RECT 62.000 68.300 62.800 68.400 ;
        RECT 60.500 68.200 62.800 68.300 ;
        RECT 60.500 67.700 63.600 68.200 ;
        RECT 50.800 64.800 51.600 66.400 ;
        RECT 54.000 64.200 54.600 67.600 ;
        RECT 55.600 66.300 56.400 66.400 ;
        RECT 58.800 66.300 59.400 67.600 ;
        RECT 60.500 66.400 61.100 67.700 ;
        RECT 62.000 67.600 63.600 67.700 ;
        RECT 65.000 67.600 67.600 68.400 ;
        RECT 70.000 67.600 70.800 70.400 ;
        RECT 62.800 67.200 63.600 67.600 ;
        RECT 55.600 65.700 59.500 66.300 ;
        RECT 55.600 64.800 56.400 65.700 ;
        RECT 58.800 64.200 59.400 65.700 ;
        RECT 60.400 64.800 61.200 66.400 ;
        RECT 62.200 66.200 65.800 66.600 ;
        RECT 66.800 66.200 67.400 67.600 ;
        RECT 70.000 66.800 74.000 67.600 ;
        RECT 74.800 66.800 75.600 68.400 ;
        RECT 62.000 66.000 66.000 66.200 ;
        RECT 54.000 62.200 54.800 64.200 ;
        RECT 58.800 62.200 59.600 64.200 ;
        RECT 62.000 62.200 62.800 66.000 ;
        RECT 65.200 62.200 66.000 66.000 ;
        RECT 66.800 62.200 67.600 66.200 ;
        RECT 70.000 62.200 70.800 66.800 ;
        RECT 73.200 62.200 74.000 66.800 ;
        RECT 76.400 64.800 77.200 66.400 ;
        RECT 78.000 62.200 78.800 79.800 ;
        RECT 79.600 72.400 80.400 79.800 ;
        RECT 82.800 72.800 83.600 79.800 ;
        RECT 79.600 71.800 82.200 72.400 ;
        RECT 82.800 71.800 83.800 72.800 ;
        RECT 79.600 69.600 80.600 70.400 ;
        RECT 79.800 68.800 80.600 69.600 ;
        RECT 81.600 69.800 82.200 71.800 ;
        RECT 81.600 69.000 82.600 69.800 ;
        RECT 81.600 67.400 82.200 69.000 ;
        RECT 83.200 68.400 83.800 71.800 ;
        RECT 82.800 67.600 83.800 68.400 ;
        RECT 79.600 66.800 82.200 67.400 ;
        RECT 79.600 62.200 80.400 66.800 ;
        RECT 83.200 66.200 83.800 67.600 ;
        RECT 86.000 66.800 86.800 68.400 ;
        RECT 82.800 65.600 83.800 66.200 ;
        RECT 87.600 66.200 88.400 79.800 ;
        RECT 89.200 72.300 90.000 73.200 ;
        RECT 90.800 72.300 91.600 79.800 ;
        RECT 89.200 71.700 91.600 72.300 ;
        RECT 89.200 71.600 90.000 71.700 ;
        RECT 87.600 65.600 89.400 66.200 ;
        RECT 82.800 62.200 83.600 65.600 ;
        RECT 88.600 64.400 89.400 65.600 ;
        RECT 88.600 63.600 90.000 64.400 ;
        RECT 88.600 62.200 89.400 63.600 ;
        RECT 90.800 62.200 91.600 71.700 ;
        RECT 94.000 66.800 94.800 68.400 ;
        RECT 92.400 64.800 93.200 66.400 ;
        RECT 95.600 66.200 96.400 79.800 ;
        RECT 97.200 71.600 98.000 73.200 ;
        RECT 98.800 66.800 99.600 68.400 ;
        RECT 100.400 66.200 101.200 79.800 ;
        RECT 102.000 71.600 102.800 73.200 ;
        RECT 106.200 72.400 107.000 79.800 ;
        RECT 107.600 73.600 108.400 74.400 ;
        RECT 107.800 72.400 108.400 73.600 ;
        RECT 110.600 72.600 111.400 79.800 ;
        RECT 105.200 71.600 107.200 72.400 ;
        RECT 107.800 71.800 109.200 72.400 ;
        RECT 110.600 71.800 112.400 72.600 ;
        RECT 114.800 71.800 115.600 79.800 ;
        RECT 116.400 72.400 117.200 79.800 ;
        RECT 119.600 72.400 120.400 79.800 ;
        RECT 116.400 71.800 120.400 72.400 ;
        RECT 123.800 72.400 124.600 79.800 ;
        RECT 125.200 73.600 126.000 74.400 ;
        RECT 125.400 72.400 126.000 73.600 ;
        RECT 123.800 71.800 124.800 72.400 ;
        RECT 125.400 71.800 126.800 72.400 ;
        RECT 108.400 71.600 109.200 71.800 ;
        RECT 105.200 68.800 106.000 70.400 ;
        RECT 106.600 68.400 107.200 71.600 ;
        RECT 110.000 69.600 110.800 71.200 ;
        RECT 111.600 68.400 112.200 71.800 ;
        RECT 115.000 70.400 115.600 71.800 ;
        RECT 118.800 70.400 119.600 70.800 ;
        RECT 114.800 69.800 117.200 70.400 ;
        RECT 118.800 69.800 120.400 70.400 ;
        RECT 114.800 69.600 115.600 69.800 ;
        RECT 116.400 69.600 117.200 69.800 ;
        RECT 119.600 69.600 120.400 69.800 ;
        RECT 103.600 68.200 104.400 68.400 ;
        RECT 103.600 67.600 105.200 68.200 ;
        RECT 106.600 67.600 109.200 68.400 ;
        RECT 111.600 68.300 112.400 68.400 ;
        RECT 111.600 67.700 115.500 68.300 ;
        RECT 111.600 67.600 112.400 67.700 ;
        RECT 104.400 67.200 105.200 67.600 ;
        RECT 103.800 66.200 107.400 66.600 ;
        RECT 108.400 66.200 109.000 67.600 ;
        RECT 95.600 65.600 97.400 66.200 ;
        RECT 100.400 65.600 102.200 66.200 ;
        RECT 96.600 64.400 97.400 65.600 ;
        RECT 101.400 64.400 102.200 65.600 ;
        RECT 96.600 63.600 98.000 64.400 ;
        RECT 100.400 63.600 102.200 64.400 ;
        RECT 96.600 62.200 97.400 63.600 ;
        RECT 101.400 62.200 102.200 63.600 ;
        RECT 103.600 66.000 107.600 66.200 ;
        RECT 103.600 62.200 104.400 66.000 ;
        RECT 106.800 62.200 107.600 66.000 ;
        RECT 108.400 62.200 109.200 66.200 ;
        RECT 111.600 64.200 112.200 67.600 ;
        RECT 114.900 66.400 115.500 67.700 ;
        RECT 113.200 64.800 114.000 66.400 ;
        RECT 114.800 65.600 115.600 66.400 ;
        RECT 116.600 66.200 117.200 69.600 ;
        RECT 118.000 67.600 118.800 69.200 ;
        RECT 122.800 68.800 123.600 70.400 ;
        RECT 124.200 70.300 124.800 71.800 ;
        RECT 126.000 71.600 126.800 71.800 ;
        RECT 127.600 71.600 128.400 73.200 ;
        RECT 129.200 72.300 130.000 79.800 ;
        RECT 133.200 73.600 134.000 74.400 ;
        RECT 133.200 72.400 133.800 73.600 ;
        RECT 134.600 72.400 135.400 79.800 ;
        RECT 132.400 72.300 133.800 72.400 ;
        RECT 129.200 71.800 133.800 72.300 ;
        RECT 134.400 71.800 135.400 72.400 ;
        RECT 143.600 72.400 144.400 79.800 ;
        RECT 145.200 72.400 146.000 72.600 ;
        RECT 148.000 72.400 149.600 79.800 ;
        RECT 143.600 71.800 146.000 72.400 ;
        RECT 147.600 71.800 149.600 72.400 ;
        RECT 151.800 72.400 152.600 72.600 ;
        RECT 153.200 72.400 154.000 79.800 ;
        RECT 151.800 71.800 154.000 72.400 ;
        RECT 129.200 71.700 133.200 71.800 ;
        RECT 127.700 70.300 128.300 71.600 ;
        RECT 124.200 69.700 128.300 70.300 ;
        RECT 124.200 68.400 124.800 69.700 ;
        RECT 121.200 68.200 122.000 68.400 ;
        RECT 121.200 67.600 122.800 68.200 ;
        RECT 124.200 67.600 126.800 68.400 ;
        RECT 122.000 67.200 122.800 67.600 ;
        RECT 121.400 66.200 125.000 66.600 ;
        RECT 126.000 66.200 126.600 67.600 ;
        RECT 129.200 66.200 130.000 71.700 ;
        RECT 132.400 71.600 133.200 71.700 ;
        RECT 134.400 68.400 135.000 71.800 ;
        RECT 147.600 70.400 148.200 71.800 ;
        RECT 151.800 71.200 152.400 71.800 ;
        RECT 149.000 70.600 152.400 71.200 ;
        RECT 154.800 71.400 155.600 79.800 ;
        RECT 159.200 76.400 160.000 79.800 ;
        RECT 158.000 75.800 160.000 76.400 ;
        RECT 163.600 75.800 164.400 79.800 ;
        RECT 167.800 75.800 169.000 79.800 ;
        RECT 158.000 75.000 158.800 75.800 ;
        RECT 163.600 75.200 164.200 75.800 ;
        RECT 161.400 74.600 165.000 75.200 ;
        RECT 167.600 75.000 168.400 75.800 ;
        RECT 161.400 74.400 162.200 74.600 ;
        RECT 164.200 74.400 165.000 74.600 ;
        RECT 158.000 73.000 158.800 73.200 ;
        RECT 162.600 73.000 163.400 73.200 ;
        RECT 158.000 72.400 163.400 73.000 ;
        RECT 164.000 73.000 166.200 73.600 ;
        RECT 164.000 71.800 164.600 73.000 ;
        RECT 165.400 72.800 166.200 73.000 ;
        RECT 167.800 73.200 169.200 74.000 ;
        RECT 167.800 72.200 168.400 73.200 ;
        RECT 159.800 71.400 164.600 71.800 ;
        RECT 154.800 71.200 164.600 71.400 ;
        RECT 166.000 71.600 168.400 72.200 ;
        RECT 154.800 71.000 160.600 71.200 ;
        RECT 154.800 70.800 160.400 71.000 ;
        RECT 149.000 70.400 149.800 70.600 ;
        RECT 166.000 70.400 166.600 71.600 ;
        RECT 172.400 71.200 173.200 79.800 ;
        RECT 176.600 78.400 177.400 79.800 ;
        RECT 175.600 77.600 177.400 78.400 ;
        RECT 176.600 72.400 177.400 77.600 ;
        RECT 178.000 73.600 178.800 74.400 ;
        RECT 178.200 72.400 178.800 73.600 ;
        RECT 176.600 71.800 177.600 72.400 ;
        RECT 178.200 72.300 179.600 72.400 ;
        RECT 180.400 72.300 181.200 72.400 ;
        RECT 178.200 71.800 181.200 72.300 ;
        RECT 169.000 70.600 173.200 71.200 ;
        RECT 169.000 70.400 169.800 70.600 ;
        RECT 135.600 70.300 136.400 70.400 ;
        RECT 143.600 70.300 144.400 70.400 ;
        RECT 135.600 69.700 144.400 70.300 ;
        RECT 135.600 68.800 136.400 69.700 ;
        RECT 143.600 69.600 144.400 69.700 ;
        RECT 146.800 69.800 148.200 70.400 ;
        RECT 161.200 70.200 162.000 70.400 ;
        RECT 151.200 69.800 152.000 70.000 ;
        RECT 146.800 69.600 148.600 69.800 ;
        RECT 147.600 69.200 148.600 69.600 ;
        RECT 130.800 66.800 131.600 68.400 ;
        RECT 132.400 67.600 135.000 68.400 ;
        RECT 137.200 68.200 138.000 68.400 ;
        RECT 136.400 67.600 138.000 68.200 ;
        RECT 143.600 67.600 145.200 68.400 ;
        RECT 146.400 67.600 147.200 68.400 ;
        RECT 132.600 66.200 133.200 67.600 ;
        RECT 136.400 67.200 137.200 67.600 ;
        RECT 146.600 67.200 147.200 67.600 ;
        RECT 145.200 66.800 146.000 67.000 ;
        RECT 134.200 66.200 137.800 66.600 ;
        RECT 143.600 66.200 146.000 66.800 ;
        RECT 146.600 66.400 147.400 67.200 ;
        RECT 115.000 64.800 115.800 65.600 ;
        RECT 111.600 62.200 112.400 64.200 ;
        RECT 116.400 62.200 117.200 66.200 ;
        RECT 121.200 66.000 125.200 66.200 ;
        RECT 121.200 62.200 122.000 66.000 ;
        RECT 124.400 62.200 125.200 66.000 ;
        RECT 126.000 62.200 126.800 66.200 ;
        RECT 128.200 65.600 130.000 66.200 ;
        RECT 128.200 62.200 129.000 65.600 ;
        RECT 132.400 62.200 133.200 66.200 ;
        RECT 134.000 66.000 138.000 66.200 ;
        RECT 134.000 62.200 134.800 66.000 ;
        RECT 137.200 62.200 138.000 66.000 ;
        RECT 143.600 62.200 144.400 66.200 ;
        RECT 148.000 65.800 148.600 69.200 ;
        RECT 149.400 69.200 152.000 69.800 ;
        RECT 157.000 69.600 162.000 70.200 ;
        RECT 166.000 69.600 166.800 70.400 ;
        RECT 170.600 69.800 171.400 70.000 ;
        RECT 157.000 69.400 157.800 69.600 ;
        RECT 159.600 69.400 160.400 69.600 ;
        RECT 149.400 68.600 150.000 69.200 ;
        RECT 149.200 67.800 150.000 68.600 ;
        RECT 158.600 68.400 159.400 68.600 ;
        RECT 166.000 68.400 166.600 69.600 ;
        RECT 167.600 69.200 171.400 69.800 ;
        RECT 167.600 69.000 168.400 69.200 ;
        RECT 152.400 68.200 154.000 68.400 ;
        RECT 150.600 67.600 154.000 68.200 ;
        RECT 155.600 67.800 166.600 68.400 ;
        RECT 155.600 67.600 157.200 67.800 ;
        RECT 150.600 67.200 151.200 67.600 ;
        RECT 149.200 66.600 151.200 67.200 ;
        RECT 151.800 66.800 152.600 67.000 ;
        RECT 149.200 66.400 150.800 66.600 ;
        RECT 151.800 66.200 154.000 66.800 ;
        RECT 148.000 64.400 149.600 65.800 ;
        RECT 146.800 63.600 149.600 64.400 ;
        RECT 148.000 62.200 149.600 63.600 ;
        RECT 153.200 62.200 154.000 66.200 ;
        RECT 154.800 62.200 155.600 67.000 ;
        RECT 159.800 65.600 160.400 67.800 ;
        RECT 165.400 67.600 166.200 67.800 ;
        RECT 172.400 67.200 173.200 70.600 ;
        RECT 175.600 68.800 176.400 70.400 ;
        RECT 177.000 68.400 177.600 71.800 ;
        RECT 178.800 71.700 181.200 71.800 ;
        RECT 178.800 71.600 179.600 71.700 ;
        RECT 180.400 71.600 181.200 71.700 ;
        RECT 174.000 68.200 174.800 68.400 ;
        RECT 174.000 67.600 175.600 68.200 ;
        RECT 177.000 67.600 179.600 68.400 ;
        RECT 174.800 67.200 175.600 67.600 ;
        RECT 169.400 66.600 173.200 67.200 ;
        RECT 169.400 66.400 170.200 66.600 ;
        RECT 158.000 64.200 158.800 65.000 ;
        RECT 159.600 64.800 160.400 65.600 ;
        RECT 161.400 65.400 162.200 65.600 ;
        RECT 161.400 64.800 164.200 65.400 ;
        RECT 163.600 64.200 164.200 64.800 ;
        RECT 167.600 64.200 168.400 65.000 ;
        RECT 158.000 63.600 160.000 64.200 ;
        RECT 159.200 62.200 160.000 63.600 ;
        RECT 163.600 62.200 164.400 64.200 ;
        RECT 167.600 63.600 169.000 64.200 ;
        RECT 167.800 62.200 169.000 63.600 ;
        RECT 172.400 62.200 173.200 66.600 ;
        RECT 174.200 66.200 177.800 66.600 ;
        RECT 178.800 66.200 179.400 67.600 ;
        RECT 174.000 66.000 178.000 66.200 ;
        RECT 174.000 62.200 174.800 66.000 ;
        RECT 177.200 62.200 178.000 66.000 ;
        RECT 178.800 62.200 179.600 66.200 ;
        RECT 180.400 64.800 181.200 66.400 ;
        RECT 182.000 62.200 182.800 79.800 ;
        RECT 184.200 78.400 185.000 79.800 ;
        RECT 184.200 77.600 186.000 78.400 ;
        RECT 184.200 72.600 185.000 77.600 ;
        RECT 184.200 71.800 186.000 72.600 ;
        RECT 183.600 69.600 184.400 71.200 ;
        RECT 185.200 68.400 185.800 71.800 ;
        RECT 185.200 67.600 186.000 68.400 ;
        RECT 185.200 64.200 185.800 67.600 ;
        RECT 188.400 66.800 189.200 68.400 ;
        RECT 186.800 64.800 187.600 66.400 ;
        RECT 190.000 66.200 190.800 79.800 ;
        RECT 193.800 78.400 194.600 79.800 ;
        RECT 200.600 78.400 201.400 79.800 ;
        RECT 193.800 77.600 195.600 78.400 ;
        RECT 199.600 77.600 201.400 78.400 ;
        RECT 191.600 71.600 192.400 73.200 ;
        RECT 193.800 72.600 194.600 77.600 ;
        RECT 193.800 71.800 195.600 72.600 ;
        RECT 200.600 72.400 201.400 77.600 ;
        RECT 202.000 73.600 202.800 74.400 ;
        RECT 202.200 72.400 202.800 73.600 ;
        RECT 200.600 71.800 201.600 72.400 ;
        RECT 202.200 71.800 203.600 72.400 ;
        RECT 193.200 69.600 194.000 71.200 ;
        RECT 194.800 68.400 195.400 71.800 ;
        RECT 199.600 68.800 200.400 70.400 ;
        RECT 201.000 68.400 201.600 71.800 ;
        RECT 202.800 71.600 203.600 71.800 ;
        RECT 204.400 72.300 205.200 79.800 ;
        RECT 208.400 73.600 209.200 74.400 ;
        RECT 208.400 72.400 209.000 73.600 ;
        RECT 209.800 72.400 210.600 79.800 ;
        RECT 207.600 72.300 209.000 72.400 ;
        RECT 204.400 71.800 209.000 72.300 ;
        RECT 204.400 71.700 208.400 71.800 ;
        RECT 194.800 67.600 195.600 68.400 ;
        RECT 198.000 68.200 198.800 68.400 ;
        RECT 198.000 67.600 199.600 68.200 ;
        RECT 201.000 67.600 203.600 68.400 ;
        RECT 190.000 65.600 191.800 66.200 ;
        RECT 185.200 62.200 186.000 64.200 ;
        RECT 191.000 62.200 191.800 65.600 ;
        RECT 194.800 64.200 195.400 67.600 ;
        RECT 198.800 67.200 199.600 67.600 ;
        RECT 196.400 64.800 197.200 66.400 ;
        RECT 198.200 66.200 201.800 66.600 ;
        RECT 202.800 66.200 203.400 67.600 ;
        RECT 198.000 66.000 202.000 66.200 ;
        RECT 194.800 62.200 195.600 64.200 ;
        RECT 198.000 62.200 198.800 66.000 ;
        RECT 201.200 62.200 202.000 66.000 ;
        RECT 202.800 62.200 203.600 66.200 ;
        RECT 204.400 62.200 205.200 71.700 ;
        RECT 207.600 71.600 208.400 71.700 ;
        RECT 209.600 71.600 211.600 72.400 ;
        RECT 214.000 71.800 214.800 79.800 ;
        RECT 215.600 72.400 216.400 79.800 ;
        RECT 218.800 72.400 219.600 79.800 ;
        RECT 215.600 71.800 219.600 72.400 ;
        RECT 209.600 68.400 210.200 71.600 ;
        RECT 214.200 70.400 214.800 71.800 ;
        RECT 218.000 70.400 218.800 70.800 ;
        RECT 210.800 70.300 211.600 70.400 ;
        RECT 212.400 70.300 213.200 70.400 ;
        RECT 210.800 69.700 213.200 70.300 ;
        RECT 210.800 68.800 211.600 69.700 ;
        RECT 212.400 69.600 213.200 69.700 ;
        RECT 214.000 69.800 216.400 70.400 ;
        RECT 218.000 69.800 219.600 70.400 ;
        RECT 214.000 69.600 214.800 69.800 ;
        RECT 207.600 67.600 210.200 68.400 ;
        RECT 212.400 68.200 213.200 68.400 ;
        RECT 211.600 67.600 213.200 68.200 ;
        RECT 206.000 64.800 206.800 66.400 ;
        RECT 207.800 66.200 208.400 67.600 ;
        RECT 211.600 67.200 212.400 67.600 ;
        RECT 209.400 66.200 213.000 66.600 ;
        RECT 215.800 66.400 216.400 69.800 ;
        RECT 218.800 69.600 219.600 69.800 ;
        RECT 217.200 68.300 218.000 69.200 ;
        RECT 222.000 68.300 222.800 79.800 ;
        RECT 217.200 67.700 222.800 68.300 ;
        RECT 217.200 67.600 218.000 67.700 ;
        RECT 207.600 62.200 208.400 66.200 ;
        RECT 209.200 66.000 213.200 66.200 ;
        RECT 209.200 62.200 210.000 66.000 ;
        RECT 212.400 62.200 213.200 66.000 ;
        RECT 214.000 65.600 214.800 66.400 ;
        RECT 214.200 64.800 215.000 65.600 ;
        RECT 215.600 62.200 216.400 66.400 ;
        RECT 220.400 64.800 221.200 66.400 ;
        RECT 222.000 62.200 222.800 67.700 ;
        RECT 223.600 64.800 224.400 66.400 ;
        RECT 225.200 62.200 226.000 79.800 ;
        RECT 229.400 74.400 230.200 79.800 ;
        RECT 228.400 73.600 230.200 74.400 ;
        RECT 230.800 73.600 231.600 74.400 ;
        RECT 229.400 72.400 230.200 73.600 ;
        RECT 231.000 72.400 231.600 73.600 ;
        RECT 229.400 71.800 230.400 72.400 ;
        RECT 231.000 72.300 232.400 72.400 ;
        RECT 233.200 72.300 234.000 79.800 ;
        RECT 231.000 71.800 234.000 72.300 ;
        RECT 236.400 71.800 237.200 79.800 ;
        RECT 238.000 72.400 238.800 79.800 ;
        RECT 241.200 72.400 242.000 79.800 ;
        RECT 242.800 75.800 243.600 79.800 ;
        RECT 243.000 75.600 243.600 75.800 ;
        RECT 246.000 75.800 246.800 79.800 ;
        RECT 246.000 75.600 246.600 75.800 ;
        RECT 243.000 75.000 246.600 75.600 ;
        RECT 243.000 72.400 243.600 75.000 ;
        RECT 244.400 72.800 245.200 74.400 ;
        RECT 251.800 72.400 252.600 79.800 ;
        RECT 253.200 73.600 254.000 74.400 ;
        RECT 253.400 72.400 254.000 73.600 ;
        RECT 238.000 71.800 242.000 72.400 ;
        RECT 226.800 70.300 227.600 70.400 ;
        RECT 228.400 70.300 229.200 70.400 ;
        RECT 226.800 69.700 229.200 70.300 ;
        RECT 226.800 69.600 227.600 69.700 ;
        RECT 228.400 68.800 229.200 69.700 ;
        RECT 229.800 68.400 230.400 71.800 ;
        RECT 231.600 71.700 234.000 71.800 ;
        RECT 231.600 71.600 232.400 71.700 ;
        RECT 226.800 68.200 227.600 68.400 ;
        RECT 226.800 67.600 228.400 68.200 ;
        RECT 229.800 67.600 232.400 68.400 ;
        RECT 227.600 67.200 228.400 67.600 ;
        RECT 227.000 66.200 230.600 66.600 ;
        RECT 231.600 66.200 232.200 67.600 ;
        RECT 226.800 66.000 230.800 66.200 ;
        RECT 226.800 62.200 227.600 66.000 ;
        RECT 230.000 62.200 230.800 66.000 ;
        RECT 231.600 62.200 232.400 66.200 ;
        RECT 233.200 62.200 234.000 71.700 ;
        RECT 236.600 70.400 237.200 71.800 ;
        RECT 242.800 71.600 243.600 72.400 ;
        RECT 240.400 70.400 241.200 70.800 ;
        RECT 236.400 69.800 238.800 70.400 ;
        RECT 240.400 69.800 242.000 70.400 ;
        RECT 236.400 69.600 237.200 69.800 ;
        RECT 234.800 66.300 235.600 66.400 ;
        RECT 236.400 66.300 237.200 66.400 ;
        RECT 234.800 65.700 237.200 66.300 ;
        RECT 238.200 66.200 238.800 69.800 ;
        RECT 241.200 69.600 242.000 69.800 ;
        RECT 239.600 67.600 240.400 69.200 ;
        RECT 243.000 68.400 243.600 71.600 ;
        RECT 247.600 70.800 248.400 72.400 ;
        RECT 251.800 71.800 252.800 72.400 ;
        RECT 253.400 71.800 254.800 72.400 ;
        RECT 245.200 69.600 246.800 70.400 ;
        RECT 250.800 68.800 251.600 70.400 ;
        RECT 252.200 68.400 252.800 71.800 ;
        RECT 254.000 71.600 254.800 71.800 ;
        RECT 243.000 68.200 244.600 68.400 ;
        RECT 249.200 68.200 250.000 68.400 ;
        RECT 243.000 67.800 244.800 68.200 ;
        RECT 234.800 64.800 235.600 65.700 ;
        RECT 236.400 65.600 237.200 65.700 ;
        RECT 236.600 64.800 237.400 65.600 ;
        RECT 238.000 62.200 238.800 66.200 ;
        RECT 244.000 66.300 244.800 67.800 ;
        RECT 249.200 67.600 250.800 68.200 ;
        RECT 252.200 67.600 254.800 68.400 ;
        RECT 250.000 67.200 250.800 67.600 ;
        RECT 246.000 66.300 246.800 66.400 ;
        RECT 244.000 65.700 246.800 66.300 ;
        RECT 249.400 66.200 253.000 66.600 ;
        RECT 254.000 66.200 254.600 67.600 ;
        RECT 255.600 66.800 256.400 68.400 ;
        RECT 257.200 66.200 258.000 79.800 ;
        RECT 258.800 71.600 259.600 73.200 ;
        RECT 244.000 62.200 244.800 65.700 ;
        RECT 246.000 65.600 246.800 65.700 ;
        RECT 249.200 66.000 253.200 66.200 ;
        RECT 249.200 62.200 250.000 66.000 ;
        RECT 252.400 62.200 253.200 66.000 ;
        RECT 254.000 62.200 254.800 66.200 ;
        RECT 257.200 65.600 259.000 66.200 ;
        RECT 258.200 64.400 259.000 65.600 ;
        RECT 258.200 63.600 259.600 64.400 ;
        RECT 258.200 62.200 259.000 63.600 ;
        RECT 260.400 62.200 261.200 79.800 ;
        RECT 265.200 70.300 266.000 79.800 ;
        RECT 269.400 72.400 270.200 79.800 ;
        RECT 275.400 78.400 276.200 79.800 ;
        RECT 275.400 77.600 277.200 78.400 ;
        RECT 270.800 73.600 271.600 74.400 ;
        RECT 271.000 72.400 271.600 73.600 ;
        RECT 274.000 73.600 274.800 74.400 ;
        RECT 274.000 72.400 274.600 73.600 ;
        RECT 275.400 72.400 276.200 77.600 ;
        RECT 282.200 72.600 283.000 79.800 ;
        RECT 286.000 75.800 286.800 79.800 ;
        RECT 286.200 75.600 286.800 75.800 ;
        RECT 289.200 75.800 290.000 79.800 ;
        RECT 289.200 75.600 289.800 75.800 ;
        RECT 286.200 75.000 289.800 75.600 ;
        RECT 287.600 72.800 288.400 74.400 ;
        RECT 269.400 71.800 270.400 72.400 ;
        RECT 271.000 71.800 272.400 72.400 ;
        RECT 269.800 70.400 270.400 71.800 ;
        RECT 271.600 71.600 272.400 71.800 ;
        RECT 273.200 71.800 274.600 72.400 ;
        RECT 275.200 71.800 276.200 72.400 ;
        RECT 281.200 71.800 283.000 72.600 ;
        RECT 289.200 72.400 289.800 75.000 ;
        RECT 273.200 71.600 274.000 71.800 ;
        RECT 268.400 70.300 269.200 70.400 ;
        RECT 265.200 69.700 269.200 70.300 ;
        RECT 262.000 64.800 262.800 66.400 ;
        RECT 263.600 64.800 264.400 66.400 ;
        RECT 265.200 62.200 266.000 69.700 ;
        RECT 268.400 68.800 269.200 69.700 ;
        RECT 269.800 69.600 270.800 70.400 ;
        RECT 269.800 68.400 270.400 69.600 ;
        RECT 275.200 68.400 275.800 71.800 ;
        RECT 276.400 68.800 277.200 70.400 ;
        RECT 281.400 68.400 282.000 71.800 ;
        RECT 282.800 69.600 283.600 71.200 ;
        RECT 284.400 70.800 285.200 72.400 ;
        RECT 289.200 71.600 290.000 72.400 ;
        RECT 297.200 72.300 298.000 79.800 ;
        RECT 299.600 73.600 300.400 74.400 ;
        RECT 299.600 72.400 300.200 73.600 ;
        RECT 301.000 72.400 301.800 79.800 ;
        RECT 298.800 72.300 300.200 72.400 ;
        RECT 297.200 71.800 300.200 72.300 ;
        RECT 300.800 71.800 301.800 72.400 ;
        RECT 297.200 71.700 299.600 71.800 ;
        RECT 286.000 69.600 287.600 70.400 ;
        RECT 289.200 68.400 289.800 71.600 ;
        RECT 266.800 68.200 267.600 68.400 ;
        RECT 266.800 67.600 268.400 68.200 ;
        RECT 269.800 67.600 272.400 68.400 ;
        RECT 273.200 67.600 275.800 68.400 ;
        RECT 278.000 68.300 278.800 68.400 ;
        RECT 279.600 68.300 280.400 68.400 ;
        RECT 278.000 68.200 280.400 68.300 ;
        RECT 277.200 67.700 280.400 68.200 ;
        RECT 277.200 67.600 278.800 67.700 ;
        RECT 279.600 67.600 280.400 67.700 ;
        RECT 281.200 68.300 282.000 68.400 ;
        RECT 282.800 68.300 283.600 68.400 ;
        RECT 281.200 67.700 283.600 68.300 ;
        RECT 288.200 68.200 289.800 68.400 ;
        RECT 281.200 67.600 282.000 67.700 ;
        RECT 282.800 67.600 283.600 67.700 ;
        RECT 288.000 67.800 289.800 68.200 ;
        RECT 290.800 68.300 291.600 68.400 ;
        RECT 295.600 68.300 296.400 68.400 ;
        RECT 267.600 67.200 268.400 67.600 ;
        RECT 267.000 66.200 270.600 66.600 ;
        RECT 271.600 66.200 272.200 67.600 ;
        RECT 273.400 66.200 274.000 67.600 ;
        RECT 277.200 67.200 278.000 67.600 ;
        RECT 275.000 66.200 278.600 66.600 ;
        RECT 266.800 66.000 270.800 66.200 ;
        RECT 266.800 62.200 267.600 66.000 ;
        RECT 270.000 62.200 270.800 66.000 ;
        RECT 271.600 62.200 272.400 66.200 ;
        RECT 273.200 62.200 274.000 66.200 ;
        RECT 274.800 66.000 278.800 66.200 ;
        RECT 274.800 62.200 275.600 66.000 ;
        RECT 278.000 62.200 278.800 66.000 ;
        RECT 279.600 64.800 280.400 66.400 ;
        RECT 281.400 64.200 282.000 67.600 ;
        RECT 281.200 62.200 282.000 64.200 ;
        RECT 288.000 62.200 288.800 67.800 ;
        RECT 290.800 67.700 296.400 68.300 ;
        RECT 290.800 67.600 291.600 67.700 ;
        RECT 295.600 67.600 296.400 67.700 ;
        RECT 295.600 64.800 296.400 66.400 ;
        RECT 297.200 62.200 298.000 71.700 ;
        RECT 298.800 71.600 299.600 71.700 ;
        RECT 298.800 70.300 299.600 70.400 ;
        RECT 300.800 70.300 301.400 71.800 ;
        RECT 298.800 69.700 301.400 70.300 ;
        RECT 298.800 69.600 299.600 69.700 ;
        RECT 300.800 68.400 301.400 69.700 ;
        RECT 302.000 68.800 302.800 70.400 ;
        RECT 298.800 67.600 301.400 68.400 ;
        RECT 303.600 68.200 304.400 68.400 ;
        RECT 302.800 67.600 304.400 68.200 ;
        RECT 299.000 66.200 299.600 67.600 ;
        RECT 302.800 67.200 303.600 67.600 ;
        RECT 300.600 66.200 304.200 66.600 ;
        RECT 298.800 62.200 299.600 66.200 ;
        RECT 300.400 66.000 304.400 66.200 ;
        RECT 300.400 62.200 301.200 66.000 ;
        RECT 303.600 62.200 304.400 66.000 ;
        RECT 305.200 62.200 306.000 79.800 ;
        RECT 311.000 72.400 311.800 79.800 ;
        RECT 312.400 73.600 313.200 74.400 ;
        RECT 312.600 72.400 313.200 73.600 ;
        RECT 311.000 71.800 312.000 72.400 ;
        RECT 312.600 72.300 314.000 72.400 ;
        RECT 314.800 72.300 315.600 79.800 ;
        RECT 312.600 71.800 315.600 72.300 ;
        RECT 318.000 71.800 318.800 79.800 ;
        RECT 319.600 72.400 320.400 79.800 ;
        RECT 322.800 72.400 323.600 79.800 ;
        RECT 319.600 71.800 323.600 72.400 ;
        RECT 325.000 72.600 325.800 79.800 ;
        RECT 325.000 71.800 326.800 72.600 ;
        RECT 311.400 70.400 312.000 71.800 ;
        RECT 313.200 71.700 315.600 71.800 ;
        RECT 313.200 71.600 314.000 71.700 ;
        RECT 310.000 68.800 310.800 70.400 ;
        RECT 311.400 69.600 312.400 70.400 ;
        RECT 311.400 68.400 312.000 69.600 ;
        RECT 308.400 68.200 309.200 68.400 ;
        RECT 308.400 67.600 310.000 68.200 ;
        RECT 311.400 67.600 314.000 68.400 ;
        RECT 309.200 67.200 310.000 67.600 ;
        RECT 306.800 64.800 307.600 66.400 ;
        RECT 308.600 66.200 312.200 66.600 ;
        RECT 313.200 66.200 313.800 67.600 ;
        RECT 308.400 66.000 312.400 66.200 ;
        RECT 308.400 62.200 309.200 66.000 ;
        RECT 311.600 62.200 312.400 66.000 ;
        RECT 313.200 62.200 314.000 66.200 ;
        RECT 314.800 62.200 315.600 71.700 ;
        RECT 318.200 70.400 318.800 71.800 ;
        RECT 322.000 70.400 322.800 70.800 ;
        RECT 318.000 69.800 320.400 70.400 ;
        RECT 322.000 69.800 323.600 70.400 ;
        RECT 318.000 69.600 318.800 69.800 ;
        RECT 319.800 66.400 320.400 69.800 ;
        RECT 322.800 69.600 323.600 69.800 ;
        RECT 324.400 69.600 325.200 71.200 ;
        RECT 321.200 67.600 322.000 69.200 ;
        RECT 326.000 68.400 326.600 71.800 ;
        RECT 326.000 67.600 326.800 68.400 ;
        RECT 316.400 66.300 317.200 66.400 ;
        RECT 318.000 66.300 318.800 66.400 ;
        RECT 316.400 65.700 318.800 66.300 ;
        RECT 316.400 64.800 317.200 65.700 ;
        RECT 318.000 65.600 318.800 65.700 ;
        RECT 318.200 64.800 319.000 65.600 ;
        RECT 319.600 62.200 320.400 66.400 ;
        RECT 326.000 64.400 326.600 67.600 ;
        RECT 327.600 66.300 328.400 66.400 ;
        RECT 329.200 66.300 330.000 79.800 ;
        RECT 332.400 72.400 333.200 79.800 ;
        RECT 334.000 72.400 334.800 72.600 ;
        RECT 336.800 72.400 338.400 79.800 ;
        RECT 332.400 71.800 334.800 72.400 ;
        RECT 336.400 71.800 338.400 72.400 ;
        RECT 340.600 72.400 341.400 72.600 ;
        RECT 342.000 72.400 342.800 79.800 ;
        RECT 340.600 71.800 342.800 72.400 ;
        RECT 336.400 70.400 337.000 71.800 ;
        RECT 340.600 71.200 341.200 71.800 ;
        RECT 337.800 70.600 341.200 71.200 ;
        RECT 343.600 71.400 344.400 79.800 ;
        RECT 348.000 76.400 348.800 79.800 ;
        RECT 346.800 75.800 348.800 76.400 ;
        RECT 352.400 75.800 353.200 79.800 ;
        RECT 356.600 75.800 357.800 79.800 ;
        RECT 346.800 75.000 347.600 75.800 ;
        RECT 352.400 75.200 353.000 75.800 ;
        RECT 350.200 74.600 353.800 75.200 ;
        RECT 356.400 75.000 357.200 75.800 ;
        RECT 350.200 74.400 351.000 74.600 ;
        RECT 353.000 74.400 353.800 74.600 ;
        RECT 346.800 73.000 347.600 73.200 ;
        RECT 351.400 73.000 352.200 73.200 ;
        RECT 346.800 72.400 352.200 73.000 ;
        RECT 352.800 73.000 355.000 73.600 ;
        RECT 352.800 71.800 353.400 73.000 ;
        RECT 354.200 72.800 355.000 73.000 ;
        RECT 356.600 73.200 358.000 74.000 ;
        RECT 356.600 72.200 357.200 73.200 ;
        RECT 348.600 71.400 353.400 71.800 ;
        RECT 343.600 71.200 353.400 71.400 ;
        RECT 354.800 71.600 357.200 72.200 ;
        RECT 343.600 71.000 349.400 71.200 ;
        RECT 343.600 70.800 349.200 71.000 ;
        RECT 337.800 70.400 338.600 70.600 ;
        RECT 335.600 69.800 337.000 70.400 ;
        RECT 350.000 70.200 350.800 70.400 ;
        RECT 340.000 69.800 340.800 70.000 ;
        RECT 335.600 69.600 337.400 69.800 ;
        RECT 336.400 69.200 337.400 69.600 ;
        RECT 332.400 68.300 334.000 68.400 ;
        RECT 330.900 67.700 334.000 68.300 ;
        RECT 330.900 66.400 331.500 67.700 ;
        RECT 332.400 67.600 334.000 67.700 ;
        RECT 335.200 67.600 336.000 68.400 ;
        RECT 335.400 67.200 336.000 67.600 ;
        RECT 334.000 66.800 334.800 67.000 ;
        RECT 327.600 65.700 330.000 66.300 ;
        RECT 327.600 64.800 328.400 65.700 ;
        RECT 326.000 62.200 326.800 64.400 ;
        RECT 329.200 62.200 330.000 65.700 ;
        RECT 330.800 64.800 331.600 66.400 ;
        RECT 332.400 66.200 334.800 66.800 ;
        RECT 335.400 66.400 336.200 67.200 ;
        RECT 332.400 62.200 333.200 66.200 ;
        RECT 336.800 65.800 337.400 69.200 ;
        RECT 338.200 69.200 340.800 69.800 ;
        RECT 345.800 69.600 350.800 70.200 ;
        RECT 345.800 69.400 346.600 69.600 ;
        RECT 348.400 69.400 349.200 69.600 ;
        RECT 338.200 68.600 338.800 69.200 ;
        RECT 338.000 67.800 338.800 68.600 ;
        RECT 347.400 68.400 348.200 68.600 ;
        RECT 354.800 68.400 355.400 71.600 ;
        RECT 361.200 71.200 362.000 79.800 ;
        RECT 357.800 70.600 362.000 71.200 ;
        RECT 362.800 71.400 363.600 79.800 ;
        RECT 367.200 76.400 368.000 79.800 ;
        RECT 366.000 75.800 368.000 76.400 ;
        RECT 371.600 75.800 372.400 79.800 ;
        RECT 375.800 75.800 377.000 79.800 ;
        RECT 366.000 75.000 366.800 75.800 ;
        RECT 371.600 75.200 372.200 75.800 ;
        RECT 369.400 74.600 373.000 75.200 ;
        RECT 375.600 75.000 376.400 75.800 ;
        RECT 369.400 74.400 370.200 74.600 ;
        RECT 372.200 74.400 373.000 74.600 ;
        RECT 366.000 73.000 366.800 73.200 ;
        RECT 370.600 73.000 371.400 73.200 ;
        RECT 366.000 72.400 371.400 73.000 ;
        RECT 372.000 73.000 374.200 73.600 ;
        RECT 372.000 71.800 372.600 73.000 ;
        RECT 373.400 72.800 374.200 73.000 ;
        RECT 375.800 73.200 377.200 74.000 ;
        RECT 375.800 72.200 376.400 73.200 ;
        RECT 367.800 71.400 372.600 71.800 ;
        RECT 362.800 71.200 372.600 71.400 ;
        RECT 374.000 71.600 376.400 72.200 ;
        RECT 362.800 71.000 368.600 71.200 ;
        RECT 362.800 70.800 368.400 71.000 ;
        RECT 357.800 70.400 358.600 70.600 ;
        RECT 359.400 69.800 360.200 70.000 ;
        RECT 356.400 69.200 360.200 69.800 ;
        RECT 356.400 69.000 357.200 69.200 ;
        RECT 341.200 68.200 342.800 68.400 ;
        RECT 339.400 67.600 342.800 68.200 ;
        RECT 344.400 67.800 355.400 68.400 ;
        RECT 344.400 67.600 346.000 67.800 ;
        RECT 339.400 67.200 340.000 67.600 ;
        RECT 338.000 66.600 340.000 67.200 ;
        RECT 340.600 66.800 341.400 67.000 ;
        RECT 338.000 66.400 339.600 66.600 ;
        RECT 340.600 66.200 342.800 66.800 ;
        RECT 336.800 64.400 338.400 65.800 ;
        RECT 336.800 63.600 339.600 64.400 ;
        RECT 336.800 62.200 338.400 63.600 ;
        RECT 342.000 62.200 342.800 66.200 ;
        RECT 343.600 62.200 344.400 67.000 ;
        RECT 348.600 65.600 349.200 67.800 ;
        RECT 353.200 67.600 355.000 67.800 ;
        RECT 361.200 67.200 362.000 70.600 ;
        RECT 369.200 70.200 370.000 70.400 ;
        RECT 365.000 69.600 370.000 70.200 ;
        RECT 365.000 69.400 365.800 69.600 ;
        RECT 367.600 69.400 368.400 69.600 ;
        RECT 366.600 68.400 367.400 68.600 ;
        RECT 374.000 68.400 374.600 71.600 ;
        RECT 380.400 71.200 381.200 79.800 ;
        RECT 377.000 70.600 381.200 71.200 ;
        RECT 377.000 70.400 377.800 70.600 ;
        RECT 378.600 69.800 379.400 70.000 ;
        RECT 375.600 69.200 379.400 69.800 ;
        RECT 375.600 69.000 376.400 69.200 ;
        RECT 363.600 67.800 374.600 68.400 ;
        RECT 380.400 68.300 381.200 70.600 ;
        RECT 382.000 68.300 382.800 68.400 ;
        RECT 363.600 67.600 365.200 67.800 ;
        RECT 358.200 66.600 362.000 67.200 ;
        RECT 358.200 66.400 359.000 66.600 ;
        RECT 346.800 64.200 347.600 65.000 ;
        RECT 348.400 64.800 349.200 65.600 ;
        RECT 350.200 65.400 351.000 65.600 ;
        RECT 350.200 64.800 353.000 65.400 ;
        RECT 352.400 64.200 353.000 64.800 ;
        RECT 356.400 64.200 357.200 65.000 ;
        RECT 346.800 63.600 348.800 64.200 ;
        RECT 348.000 62.200 348.800 63.600 ;
        RECT 352.400 62.200 353.200 64.200 ;
        RECT 356.400 63.600 357.800 64.200 ;
        RECT 356.600 62.200 357.800 63.600 ;
        RECT 361.200 62.200 362.000 66.600 ;
        RECT 362.800 62.200 363.600 67.000 ;
        RECT 367.800 65.600 368.400 67.800 ;
        RECT 372.400 67.600 374.200 67.800 ;
        RECT 380.400 67.700 382.800 68.300 ;
        RECT 380.400 67.200 381.200 67.700 ;
        RECT 377.400 66.600 381.200 67.200 ;
        RECT 382.000 66.800 382.800 67.700 ;
        RECT 377.400 66.400 378.200 66.600 ;
        RECT 366.000 64.200 366.800 65.000 ;
        RECT 367.600 64.800 368.400 65.600 ;
        RECT 369.400 65.400 370.200 65.600 ;
        RECT 369.400 64.800 372.200 65.400 ;
        RECT 371.600 64.200 372.200 64.800 ;
        RECT 375.600 64.200 376.400 65.000 ;
        RECT 366.000 63.600 368.000 64.200 ;
        RECT 367.200 62.200 368.000 63.600 ;
        RECT 371.600 62.200 372.400 64.200 ;
        RECT 375.600 63.600 377.000 64.200 ;
        RECT 375.800 62.200 377.000 63.600 ;
        RECT 380.400 62.200 381.200 66.600 ;
        RECT 383.600 66.300 384.400 79.800 ;
        RECT 385.200 71.600 386.000 73.200 ;
        RECT 388.400 70.300 389.200 79.800 ;
        RECT 392.600 78.400 393.400 79.800 ;
        RECT 391.600 77.600 393.400 78.400 ;
        RECT 392.600 72.400 393.400 77.600 ;
        RECT 394.000 73.600 394.800 74.400 ;
        RECT 394.200 72.400 394.800 73.600 ;
        RECT 397.200 73.600 398.000 74.400 ;
        RECT 397.200 72.400 397.800 73.600 ;
        RECT 398.600 72.400 399.400 79.800 ;
        RECT 392.600 71.800 393.600 72.400 ;
        RECT 394.200 71.800 395.600 72.400 ;
        RECT 391.600 70.300 392.400 70.400 ;
        RECT 388.400 69.700 392.400 70.300 ;
        RECT 386.800 66.300 387.600 66.400 ;
        RECT 383.600 65.700 387.600 66.300 ;
        RECT 383.600 65.600 385.400 65.700 ;
        RECT 384.600 62.200 385.400 65.600 ;
        RECT 386.800 64.800 387.600 65.700 ;
        RECT 388.400 62.200 389.200 69.700 ;
        RECT 391.600 68.800 392.400 69.700 ;
        RECT 393.000 68.400 393.600 71.800 ;
        RECT 394.800 71.600 395.600 71.800 ;
        RECT 396.400 71.800 397.800 72.400 ;
        RECT 398.400 71.800 399.400 72.400 ;
        RECT 396.400 71.600 397.200 71.800 ;
        RECT 394.900 70.300 395.500 71.600 ;
        RECT 398.400 70.300 399.000 71.800 ;
        RECT 394.900 69.700 399.000 70.300 ;
        RECT 398.400 68.400 399.000 69.700 ;
        RECT 399.600 68.800 400.400 70.400 ;
        RECT 390.000 68.200 390.800 68.400 ;
        RECT 390.000 67.600 391.600 68.200 ;
        RECT 393.000 67.600 395.600 68.400 ;
        RECT 396.400 67.600 399.000 68.400 ;
        RECT 401.200 68.300 402.000 68.400 ;
        RECT 402.800 68.300 403.600 68.400 ;
        RECT 401.200 68.200 403.600 68.300 ;
        RECT 400.400 67.700 403.600 68.200 ;
        RECT 400.400 67.600 402.000 67.700 ;
        RECT 390.800 67.200 391.600 67.600 ;
        RECT 390.200 66.200 393.800 66.600 ;
        RECT 394.800 66.200 395.400 67.600 ;
        RECT 396.600 66.200 397.200 67.600 ;
        RECT 400.400 67.200 401.200 67.600 ;
        RECT 402.800 66.800 403.600 67.700 ;
        RECT 404.400 68.300 405.200 79.800 ;
        RECT 406.000 71.600 406.800 73.200 ;
        RECT 409.200 70.300 410.000 79.800 ;
        RECT 410.800 71.600 411.600 73.200 ;
        RECT 412.400 70.300 413.200 70.400 ;
        RECT 409.200 69.700 413.200 70.300 ;
        RECT 407.600 68.300 408.400 68.400 ;
        RECT 404.400 67.700 408.400 68.300 ;
        RECT 398.200 66.200 401.800 66.600 ;
        RECT 404.400 66.200 405.200 67.700 ;
        RECT 407.600 66.800 408.400 67.700 ;
        RECT 409.200 66.200 410.000 69.700 ;
        RECT 412.400 69.600 413.200 69.700 ;
        RECT 412.400 66.800 413.200 68.400 ;
        RECT 390.000 66.000 394.000 66.200 ;
        RECT 390.000 62.200 390.800 66.000 ;
        RECT 393.200 62.200 394.000 66.000 ;
        RECT 394.800 62.200 395.600 66.200 ;
        RECT 396.400 62.200 397.200 66.200 ;
        RECT 398.000 66.000 402.000 66.200 ;
        RECT 398.000 62.200 398.800 66.000 ;
        RECT 401.200 62.200 402.000 66.000 ;
        RECT 404.400 65.600 406.200 66.200 ;
        RECT 409.200 65.600 411.000 66.200 ;
        RECT 405.400 62.200 406.200 65.600 ;
        RECT 410.200 62.200 411.000 65.600 ;
        RECT 414.000 62.200 414.800 79.800 ;
        RECT 417.200 70.300 418.000 79.800 ;
        RECT 419.400 72.600 420.200 79.800 ;
        RECT 419.400 71.800 421.200 72.600 ;
        RECT 418.800 70.300 419.600 71.200 ;
        RECT 417.200 69.700 419.600 70.300 ;
        RECT 415.600 64.800 416.400 66.400 ;
        RECT 417.200 62.200 418.000 69.700 ;
        RECT 418.800 69.600 419.600 69.700 ;
        RECT 420.400 68.400 421.000 71.800 ;
        RECT 420.400 67.600 421.200 68.400 ;
        RECT 420.400 64.400 421.000 67.600 ;
        RECT 423.600 66.800 424.400 68.400 ;
        RECT 425.200 66.400 426.000 79.800 ;
        RECT 426.800 71.600 427.600 73.200 ;
        RECT 428.400 68.300 429.200 79.800 ;
        RECT 431.600 72.400 432.400 79.800 ;
        RECT 434.800 72.400 435.600 79.800 ;
        RECT 431.600 71.800 435.600 72.400 ;
        RECT 436.400 71.800 437.200 79.800 ;
        RECT 438.000 72.400 438.800 79.800 ;
        RECT 439.600 72.400 440.400 72.600 ;
        RECT 438.000 71.800 440.400 72.400 ;
        RECT 442.400 71.800 444.000 79.800 ;
        RECT 445.800 72.400 446.600 72.600 ;
        RECT 447.600 72.400 448.400 79.800 ;
        RECT 445.800 71.800 448.400 72.400 ;
        RECT 456.600 71.800 458.600 79.800 ;
        RECT 462.000 72.400 462.800 79.800 ;
        RECT 466.400 78.400 468.000 79.800 ;
        RECT 466.400 77.600 469.200 78.400 ;
        RECT 463.400 72.400 464.200 72.600 ;
        RECT 462.000 71.800 464.200 72.400 ;
        RECT 466.400 72.400 468.000 77.600 ;
        RECT 470.000 72.400 470.800 72.600 ;
        RECT 471.600 72.400 472.400 79.800 ;
        RECT 466.400 71.800 468.400 72.400 ;
        RECT 470.000 71.800 472.400 72.400 ;
        RECT 475.800 72.400 476.600 79.800 ;
        RECT 477.200 73.600 478.000 74.400 ;
        RECT 477.400 72.400 478.000 73.600 ;
        RECT 482.200 72.600 483.000 79.800 ;
        RECT 475.800 71.800 476.800 72.400 ;
        RECT 477.400 71.800 478.800 72.400 ;
        RECT 481.200 71.800 483.000 72.600 ;
        RECT 486.000 72.300 486.800 79.800 ;
        RECT 488.400 73.600 489.200 74.400 ;
        RECT 488.400 72.400 489.000 73.600 ;
        RECT 489.800 72.400 490.600 79.800 ;
        RECT 494.800 73.600 495.600 74.400 ;
        RECT 494.800 72.400 495.400 73.600 ;
        RECT 496.200 72.400 497.000 79.800 ;
        RECT 487.600 72.300 489.000 72.400 ;
        RECT 486.000 71.800 489.000 72.300 ;
        RECT 489.600 71.800 490.600 72.400 ;
        RECT 494.000 71.800 495.400 72.400 ;
        RECT 496.000 71.800 497.000 72.400 ;
        RECT 502.000 72.300 502.800 79.800 ;
        RECT 504.400 73.600 505.200 74.400 ;
        RECT 504.400 72.400 505.000 73.600 ;
        RECT 505.800 72.400 506.600 79.800 ;
        RECT 503.600 72.300 505.000 72.400 ;
        RECT 502.000 71.800 505.000 72.300 ;
        RECT 505.600 71.800 506.600 72.400 ;
        RECT 510.600 72.600 511.400 79.800 ;
        RECT 517.400 74.400 518.200 79.800 ;
        RECT 517.400 73.600 518.800 74.400 ;
        RECT 517.400 72.600 518.200 73.600 ;
        RECT 510.600 71.800 512.400 72.600 ;
        RECT 516.400 71.800 518.200 72.600 ;
        RECT 522.200 72.400 523.000 79.800 ;
        RECT 528.200 78.400 529.000 79.800 ;
        RECT 528.200 77.600 530.000 78.400 ;
        RECT 523.600 73.600 524.400 74.400 ;
        RECT 523.800 72.400 524.400 73.600 ;
        RECT 526.800 73.600 527.600 74.400 ;
        RECT 526.800 72.400 527.400 73.600 ;
        RECT 528.200 72.400 529.000 77.600 ;
        RECT 522.200 71.800 523.200 72.400 ;
        RECT 523.800 71.800 525.200 72.400 ;
        RECT 432.400 70.400 433.200 70.800 ;
        RECT 436.400 70.400 437.000 71.800 ;
        RECT 442.800 70.400 443.400 71.800 ;
        RECT 444.600 70.400 445.400 70.600 ;
        RECT 431.600 69.800 433.200 70.400 ;
        RECT 434.800 69.800 437.200 70.400 ;
        RECT 431.600 69.600 432.400 69.800 ;
        RECT 433.200 68.300 434.000 69.200 ;
        RECT 428.400 67.700 434.000 68.300 ;
        RECT 422.000 64.800 422.800 66.400 ;
        RECT 425.200 65.600 427.600 66.400 ;
        RECT 420.400 62.200 421.200 64.400 ;
        RECT 426.200 62.200 427.000 65.600 ;
        RECT 428.400 62.200 429.200 67.700 ;
        RECT 433.200 67.600 434.000 67.700 ;
        RECT 430.000 64.800 430.800 66.400 ;
        RECT 434.800 66.200 435.400 69.800 ;
        RECT 436.400 69.600 437.200 69.800 ;
        RECT 438.000 70.300 438.800 70.400 ;
        RECT 442.800 70.300 443.600 70.400 ;
        RECT 438.000 69.700 443.600 70.300 ;
        RECT 444.600 69.800 446.200 70.400 ;
        RECT 438.000 69.600 438.800 69.700 ;
        RECT 442.800 69.600 443.600 69.700 ;
        RECT 445.400 69.600 446.200 69.800 ;
        RECT 442.800 68.400 443.400 69.600 ;
        RECT 438.000 67.600 439.600 68.400 ;
        RECT 440.800 67.600 441.600 68.400 ;
        RECT 441.000 67.200 441.600 67.600 ;
        RECT 442.400 67.800 443.400 68.400 ;
        RECT 444.000 68.600 444.800 68.800 ;
        RECT 444.000 68.400 446.800 68.600 ;
        RECT 444.000 68.000 448.400 68.400 ;
        RECT 446.200 67.800 448.400 68.000 ;
        RECT 439.600 66.800 440.400 67.000 ;
        RECT 434.800 62.200 435.600 66.200 ;
        RECT 436.400 65.600 437.200 66.400 ;
        RECT 438.000 66.200 440.400 66.800 ;
        RECT 441.000 66.400 441.800 67.200 ;
        RECT 436.200 64.800 437.000 65.600 ;
        RECT 438.000 62.200 438.800 66.200 ;
        RECT 442.400 65.800 443.000 67.800 ;
        RECT 446.800 67.600 448.400 67.800 ;
        RECT 450.800 68.300 451.600 68.400 ;
        RECT 454.000 68.300 454.800 69.200 ;
        RECT 455.600 68.800 456.400 70.400 ;
        RECT 457.400 68.400 458.000 71.800 ;
        RECT 463.600 71.200 464.200 71.800 ;
        RECT 463.600 70.600 467.000 71.200 ;
        RECT 466.200 70.400 467.000 70.600 ;
        RECT 467.800 70.400 468.400 71.800 ;
        RECT 458.800 68.800 459.600 70.400 ;
        RECT 464.000 69.800 464.800 70.000 ;
        RECT 467.800 69.800 469.200 70.400 ;
        RECT 464.000 69.200 466.600 69.800 ;
        RECT 466.000 68.600 466.600 69.200 ;
        RECT 467.400 69.600 469.200 69.800 ;
        RECT 467.400 69.200 468.400 69.600 ;
        RECT 450.800 67.700 454.800 68.300 ;
        RECT 457.200 68.200 458.000 68.400 ;
        RECT 460.400 68.200 461.200 68.400 ;
        RECT 450.800 67.600 451.600 67.700 ;
        RECT 454.000 67.600 454.800 67.700 ;
        RECT 455.600 67.600 458.000 68.200 ;
        RECT 459.600 67.600 461.200 68.200 ;
        RECT 462.000 68.200 463.600 68.400 ;
        RECT 462.000 67.600 465.400 68.200 ;
        RECT 466.000 67.800 466.800 68.600 ;
        RECT 443.600 66.400 445.200 67.200 ;
        RECT 445.800 66.800 446.600 67.000 ;
        RECT 445.800 66.200 448.400 66.800 ;
        RECT 455.600 66.200 456.200 67.600 ;
        RECT 459.600 67.200 460.400 67.600 ;
        RECT 464.800 67.200 465.400 67.600 ;
        RECT 463.400 66.800 464.200 67.000 ;
        RECT 457.400 66.200 461.000 66.600 ;
        RECT 462.000 66.200 464.200 66.800 ;
        RECT 464.800 66.600 466.800 67.200 ;
        RECT 465.200 66.400 466.800 66.600 ;
        RECT 442.400 62.200 444.000 65.800 ;
        RECT 447.600 62.200 448.400 66.200 ;
        RECT 454.000 62.800 454.800 66.200 ;
        RECT 455.600 63.400 456.400 66.200 ;
        RECT 457.200 66.000 461.200 66.200 ;
        RECT 457.200 62.800 458.000 66.000 ;
        RECT 454.000 62.200 458.000 62.800 ;
        RECT 460.400 62.200 461.200 66.000 ;
        RECT 462.000 62.200 462.800 66.200 ;
        RECT 467.400 65.800 468.000 69.200 ;
        RECT 474.800 68.800 475.600 70.400 ;
        RECT 476.200 68.400 476.800 71.800 ;
        RECT 478.000 71.600 478.800 71.800 ;
        RECT 481.400 68.400 482.000 71.800 ;
        RECT 486.000 71.700 488.400 71.800 ;
        RECT 482.800 70.300 483.600 71.200 ;
        RECT 484.400 70.300 485.200 70.400 ;
        RECT 482.800 69.700 485.200 70.300 ;
        RECT 482.800 69.600 483.600 69.700 ;
        RECT 484.400 69.600 485.200 69.700 ;
        RECT 468.800 67.600 469.600 68.400 ;
        RECT 470.800 67.600 472.400 68.400 ;
        RECT 473.200 68.200 474.000 68.400 ;
        RECT 473.200 67.600 474.800 68.200 ;
        RECT 476.200 67.600 478.800 68.400 ;
        RECT 481.200 68.300 482.000 68.400 ;
        RECT 484.400 68.300 485.200 68.400 ;
        RECT 481.200 67.700 485.200 68.300 ;
        RECT 481.200 67.600 482.000 67.700 ;
        RECT 484.400 67.600 485.200 67.700 ;
        RECT 468.800 67.200 469.400 67.600 ;
        RECT 474.000 67.200 474.800 67.600 ;
        RECT 468.600 66.400 469.400 67.200 ;
        RECT 470.000 66.800 470.800 67.000 ;
        RECT 470.000 66.200 472.400 66.800 ;
        RECT 473.400 66.200 477.000 66.600 ;
        RECT 478.000 66.400 478.600 67.600 ;
        RECT 466.400 62.200 468.000 65.800 ;
        RECT 471.600 62.200 472.400 66.200 ;
        RECT 473.200 66.000 477.200 66.200 ;
        RECT 473.200 62.200 474.000 66.000 ;
        RECT 476.400 62.200 477.200 66.000 ;
        RECT 478.000 62.200 478.800 66.400 ;
        RECT 479.600 64.800 480.400 66.400 ;
        RECT 481.400 64.200 482.000 67.600 ;
        RECT 484.400 64.800 485.200 66.400 ;
        RECT 481.200 62.200 482.000 64.200 ;
        RECT 486.000 62.200 486.800 71.700 ;
        RECT 487.600 71.600 488.400 71.700 ;
        RECT 487.600 70.300 488.400 70.400 ;
        RECT 489.600 70.300 490.200 71.800 ;
        RECT 494.000 71.600 494.800 71.800 ;
        RECT 487.600 69.700 490.200 70.300 ;
        RECT 487.600 69.600 488.400 69.700 ;
        RECT 489.600 68.400 490.200 69.700 ;
        RECT 490.800 68.800 491.600 70.400 ;
        RECT 492.400 70.300 493.200 70.400 ;
        RECT 496.000 70.300 496.600 71.800 ;
        RECT 502.000 71.700 504.400 71.800 ;
        RECT 492.400 69.700 496.600 70.300 ;
        RECT 492.400 69.600 493.200 69.700 ;
        RECT 496.000 68.400 496.600 69.700 ;
        RECT 497.200 68.800 498.000 70.400 ;
        RECT 487.600 67.600 490.200 68.400 ;
        RECT 492.400 68.200 493.200 68.400 ;
        RECT 491.600 67.600 493.200 68.200 ;
        RECT 494.000 67.600 496.600 68.400 ;
        RECT 498.800 68.200 499.600 68.400 ;
        RECT 498.000 67.600 499.600 68.200 ;
        RECT 487.800 66.200 488.400 67.600 ;
        RECT 491.600 67.200 492.400 67.600 ;
        RECT 489.400 66.200 493.000 66.600 ;
        RECT 494.200 66.200 494.800 67.600 ;
        RECT 498.000 67.200 498.800 67.600 ;
        RECT 495.800 66.200 499.400 66.600 ;
        RECT 487.600 62.200 488.400 66.200 ;
        RECT 489.200 66.000 493.200 66.200 ;
        RECT 489.200 62.200 490.000 66.000 ;
        RECT 492.400 62.200 493.200 66.000 ;
        RECT 494.000 62.200 494.800 66.200 ;
        RECT 495.600 66.000 499.600 66.200 ;
        RECT 495.600 62.200 496.400 66.000 ;
        RECT 498.800 62.200 499.600 66.000 ;
        RECT 500.400 64.800 501.200 66.400 ;
        RECT 502.000 62.200 502.800 71.700 ;
        RECT 503.600 71.600 504.400 71.700 ;
        RECT 503.600 70.300 504.400 70.400 ;
        RECT 505.600 70.300 506.200 71.800 ;
        RECT 503.600 69.700 506.200 70.300 ;
        RECT 503.600 69.600 504.400 69.700 ;
        RECT 505.600 68.400 506.200 69.700 ;
        RECT 506.800 68.800 507.600 70.400 ;
        RECT 510.000 69.600 510.800 71.200 ;
        RECT 511.600 68.400 512.200 71.800 ;
        RECT 516.600 68.400 517.200 71.800 ;
        RECT 518.000 69.600 518.800 71.200 ;
        RECT 519.600 70.300 520.400 70.400 ;
        RECT 521.200 70.300 522.000 70.400 ;
        RECT 519.600 69.700 522.000 70.300 ;
        RECT 519.600 69.600 520.400 69.700 ;
        RECT 521.200 68.800 522.000 69.700 ;
        RECT 522.600 70.300 523.200 71.800 ;
        RECT 524.400 71.600 525.200 71.800 ;
        RECT 526.000 71.800 527.400 72.400 ;
        RECT 528.000 71.800 529.000 72.400 ;
        RECT 532.400 71.800 533.200 79.800 ;
        RECT 535.600 72.400 536.400 79.800 ;
        RECT 534.200 71.800 536.400 72.400 ;
        RECT 537.200 72.400 538.000 79.800 ;
        RECT 537.200 71.800 539.400 72.400 ;
        RECT 540.400 71.800 541.200 79.800 ;
        RECT 526.000 71.600 526.800 71.800 ;
        RECT 526.100 70.300 526.700 71.600 ;
        RECT 522.600 69.700 526.700 70.300 ;
        RECT 522.600 68.400 523.200 69.700 ;
        RECT 528.000 68.400 528.600 71.800 ;
        RECT 529.200 68.800 530.000 70.400 ;
        RECT 532.400 69.600 533.000 71.800 ;
        RECT 534.200 71.200 534.800 71.800 ;
        RECT 533.600 70.400 534.800 71.200 ;
        RECT 538.800 71.200 539.400 71.800 ;
        RECT 538.800 70.400 540.000 71.200 ;
        RECT 503.600 67.600 506.200 68.400 ;
        RECT 508.400 68.200 509.200 68.400 ;
        RECT 507.600 67.600 509.200 68.200 ;
        RECT 511.600 68.300 512.400 68.400 ;
        RECT 514.800 68.300 515.600 68.400 ;
        RECT 511.600 67.700 515.600 68.300 ;
        RECT 511.600 67.600 512.400 67.700 ;
        RECT 514.800 67.600 515.600 67.700 ;
        RECT 516.400 67.600 517.200 68.400 ;
        RECT 519.600 68.200 520.400 68.400 ;
        RECT 519.600 67.600 521.200 68.200 ;
        RECT 522.600 67.600 525.200 68.400 ;
        RECT 526.000 67.600 528.600 68.400 ;
        RECT 530.800 68.200 531.600 68.400 ;
        RECT 530.000 67.600 531.600 68.200 ;
        RECT 503.800 66.200 504.400 67.600 ;
        RECT 507.600 67.200 508.400 67.600 ;
        RECT 505.400 66.200 509.000 66.600 ;
        RECT 503.600 62.200 504.400 66.200 ;
        RECT 505.200 66.000 509.200 66.200 ;
        RECT 505.200 62.200 506.000 66.000 ;
        RECT 508.400 62.200 509.200 66.000 ;
        RECT 511.600 64.200 512.200 67.600 ;
        RECT 513.200 64.800 514.000 66.400 ;
        RECT 514.800 64.800 515.600 66.400 ;
        RECT 516.600 64.200 517.200 67.600 ;
        RECT 520.400 67.200 521.200 67.600 ;
        RECT 519.800 66.200 523.400 66.600 ;
        RECT 524.400 66.200 525.000 67.600 ;
        RECT 526.200 66.200 526.800 67.600 ;
        RECT 530.000 67.200 530.800 67.600 ;
        RECT 527.800 66.200 531.400 66.600 ;
        RECT 511.600 62.200 512.400 64.200 ;
        RECT 516.400 62.200 517.200 64.200 ;
        RECT 519.600 66.000 523.600 66.200 ;
        RECT 519.600 62.200 520.400 66.000 ;
        RECT 522.800 62.200 523.600 66.000 ;
        RECT 524.400 62.200 525.200 66.200 ;
        RECT 526.000 62.200 526.800 66.200 ;
        RECT 527.600 66.000 531.600 66.200 ;
        RECT 527.600 62.200 528.400 66.000 ;
        RECT 530.800 62.200 531.600 66.000 ;
        RECT 532.400 62.200 533.200 69.600 ;
        RECT 534.200 67.400 534.800 70.400 ;
        RECT 535.600 70.300 536.400 70.400 ;
        RECT 537.200 70.300 538.000 70.400 ;
        RECT 535.600 69.700 538.000 70.300 ;
        RECT 535.600 68.800 536.400 69.700 ;
        RECT 537.200 68.800 538.000 69.700 ;
        RECT 538.800 67.400 539.400 70.400 ;
        RECT 540.600 69.600 541.200 71.800 ;
        RECT 542.000 71.400 542.800 79.800 ;
        RECT 546.400 76.400 547.200 79.800 ;
        RECT 545.200 75.800 547.200 76.400 ;
        RECT 550.800 75.800 551.600 79.800 ;
        RECT 555.000 75.800 556.200 79.800 ;
        RECT 545.200 75.000 546.000 75.800 ;
        RECT 550.800 75.200 551.400 75.800 ;
        RECT 548.600 74.600 552.200 75.200 ;
        RECT 554.800 75.000 555.600 75.800 ;
        RECT 548.600 74.400 549.400 74.600 ;
        RECT 551.400 74.400 552.200 74.600 ;
        RECT 545.200 73.000 546.000 73.200 ;
        RECT 549.800 73.000 550.600 73.200 ;
        RECT 545.200 72.400 550.600 73.000 ;
        RECT 551.200 73.000 553.400 73.600 ;
        RECT 551.200 71.800 551.800 73.000 ;
        RECT 552.600 72.800 553.400 73.000 ;
        RECT 555.000 73.200 556.400 74.000 ;
        RECT 555.000 72.200 555.600 73.200 ;
        RECT 547.000 71.400 551.800 71.800 ;
        RECT 542.000 71.200 551.800 71.400 ;
        RECT 553.200 71.600 555.600 72.200 ;
        RECT 542.000 71.000 547.800 71.200 ;
        RECT 542.000 70.800 547.600 71.000 ;
        RECT 548.400 70.200 549.200 70.400 ;
        RECT 534.200 66.800 536.400 67.400 ;
        RECT 535.600 62.200 536.400 66.800 ;
        RECT 537.200 66.800 539.400 67.400 ;
        RECT 537.200 62.200 538.000 66.800 ;
        RECT 540.400 62.200 541.200 69.600 ;
        RECT 544.200 69.600 549.200 70.200 ;
        RECT 544.200 69.400 545.000 69.600 ;
        RECT 546.800 69.400 547.600 69.600 ;
        RECT 545.800 68.400 546.600 68.600 ;
        RECT 553.200 68.400 553.800 71.600 ;
        RECT 559.600 71.200 560.400 79.800 ;
        RECT 556.200 70.600 560.400 71.200 ;
        RECT 561.200 71.400 562.000 79.800 ;
        RECT 565.600 76.400 566.400 79.800 ;
        RECT 564.400 75.800 566.400 76.400 ;
        RECT 570.000 75.800 570.800 79.800 ;
        RECT 574.200 75.800 575.400 79.800 ;
        RECT 564.400 75.000 565.200 75.800 ;
        RECT 570.000 75.200 570.600 75.800 ;
        RECT 567.800 74.600 571.400 75.200 ;
        RECT 574.000 75.000 574.800 75.800 ;
        RECT 567.800 74.400 568.600 74.600 ;
        RECT 570.600 74.400 571.400 74.600 ;
        RECT 564.400 73.000 565.200 73.200 ;
        RECT 569.000 73.000 569.800 73.200 ;
        RECT 564.400 72.400 569.800 73.000 ;
        RECT 570.400 73.000 572.600 73.600 ;
        RECT 570.400 71.800 571.000 73.000 ;
        RECT 571.800 72.800 572.600 73.000 ;
        RECT 574.200 73.200 575.600 74.000 ;
        RECT 574.200 72.200 574.800 73.200 ;
        RECT 566.200 71.400 571.000 71.800 ;
        RECT 561.200 71.200 571.000 71.400 ;
        RECT 572.400 71.600 574.800 72.200 ;
        RECT 561.200 71.000 567.000 71.200 ;
        RECT 561.200 70.800 566.800 71.000 ;
        RECT 556.200 70.400 557.000 70.600 ;
        RECT 557.800 69.800 558.600 70.000 ;
        RECT 554.800 69.200 558.600 69.800 ;
        RECT 554.800 69.000 555.600 69.200 ;
        RECT 542.800 67.800 553.800 68.400 ;
        RECT 542.800 67.600 544.400 67.800 ;
        RECT 542.000 62.200 542.800 67.000 ;
        RECT 547.000 65.600 547.600 67.800 ;
        RECT 550.000 67.600 550.800 67.800 ;
        RECT 552.600 67.600 553.400 67.800 ;
        RECT 559.600 67.200 560.400 70.600 ;
        RECT 567.600 70.200 568.400 70.400 ;
        RECT 563.400 69.600 568.400 70.200 ;
        RECT 563.400 69.400 564.200 69.600 ;
        RECT 566.000 69.400 566.800 69.600 ;
        RECT 565.000 68.400 565.800 68.600 ;
        RECT 572.400 68.400 573.000 71.600 ;
        RECT 578.800 71.200 579.600 79.800 ;
        RECT 580.400 72.400 581.200 79.800 ;
        RECT 580.400 71.800 582.600 72.400 ;
        RECT 575.400 70.600 579.600 71.200 ;
        RECT 575.400 70.400 576.200 70.600 ;
        RECT 577.000 69.800 577.800 70.000 ;
        RECT 574.000 69.200 577.800 69.800 ;
        RECT 574.000 69.000 574.800 69.200 ;
        RECT 562.000 67.800 573.200 68.400 ;
        RECT 562.000 67.600 563.600 67.800 ;
        RECT 556.600 66.600 560.400 67.200 ;
        RECT 556.600 66.400 557.400 66.600 ;
        RECT 545.200 64.200 546.000 65.000 ;
        RECT 546.800 64.800 547.600 65.600 ;
        RECT 548.600 65.400 549.400 65.600 ;
        RECT 548.600 64.800 551.400 65.400 ;
        RECT 550.800 64.200 551.400 64.800 ;
        RECT 554.800 64.200 555.600 65.000 ;
        RECT 545.200 63.600 547.200 64.200 ;
        RECT 546.400 62.200 547.200 63.600 ;
        RECT 550.800 62.200 551.600 64.200 ;
        RECT 554.800 63.600 556.200 64.200 ;
        RECT 555.000 62.200 556.200 63.600 ;
        RECT 559.600 62.200 560.400 66.600 ;
        RECT 561.200 62.200 562.000 67.000 ;
        RECT 566.200 65.600 566.800 67.800 ;
        RECT 567.600 67.600 568.400 67.800 ;
        RECT 571.800 67.600 573.200 67.800 ;
        RECT 578.800 67.200 579.600 70.600 ;
        RECT 582.000 71.200 582.600 71.800 ;
        RECT 582.000 70.400 583.200 71.200 ;
        RECT 580.400 68.800 581.200 70.400 ;
        RECT 582.000 67.400 582.600 70.400 ;
        RECT 575.800 66.600 579.600 67.200 ;
        RECT 575.800 66.400 576.600 66.600 ;
        RECT 564.400 64.200 565.200 65.000 ;
        RECT 566.000 64.800 566.800 65.600 ;
        RECT 567.800 65.400 568.600 65.600 ;
        RECT 567.800 64.800 570.600 65.400 ;
        RECT 570.000 64.200 570.600 64.800 ;
        RECT 574.000 64.200 574.800 65.000 ;
        RECT 564.400 63.600 566.400 64.200 ;
        RECT 565.600 62.200 566.400 63.600 ;
        RECT 570.000 62.200 570.800 64.200 ;
        RECT 574.000 63.600 575.400 64.200 ;
        RECT 574.200 62.200 575.400 63.600 ;
        RECT 578.800 62.200 579.600 66.600 ;
        RECT 580.400 66.800 582.600 67.400 ;
        RECT 580.400 62.200 581.200 66.800 ;
        RECT 2.800 57.600 3.600 59.800 ;
        RECT 8.600 58.400 9.400 59.800 ;
        RECT 8.600 57.600 10.000 58.400 ;
        RECT 2.800 54.400 3.400 57.600 ;
        RECT 4.400 55.600 5.200 57.200 ;
        RECT 8.600 56.400 9.400 57.600 ;
        RECT 13.400 56.400 14.200 59.800 ;
        RECT 17.200 57.800 18.000 59.800 ;
        RECT 7.600 55.800 9.400 56.400 ;
        RECT 12.400 55.800 14.200 56.400 ;
        RECT 2.800 53.600 3.600 54.400 ;
        RECT 4.500 54.300 5.100 55.600 ;
        RECT 6.000 54.300 6.800 55.200 ;
        RECT 4.500 53.700 6.800 54.300 ;
        RECT 6.000 53.600 6.800 53.700 ;
        RECT 1.200 50.800 2.000 52.400 ;
        RECT 2.800 50.200 3.400 53.600 ;
        RECT 1.800 49.400 3.600 50.200 ;
        RECT 1.800 42.200 2.600 49.400 ;
        RECT 7.600 42.200 8.400 55.800 ;
        RECT 10.800 53.600 11.600 55.200 ;
        RECT 9.200 50.300 10.000 50.400 ;
        RECT 12.400 50.300 13.200 55.800 ;
        RECT 15.600 55.600 16.400 57.200 ;
        RECT 17.400 54.400 18.000 57.800 ;
        RECT 23.000 56.400 23.800 59.800 ;
        RECT 22.000 55.800 23.800 56.400 ;
        RECT 27.800 55.800 29.400 59.800 ;
        RECT 17.200 53.600 18.000 54.400 ;
        RECT 20.400 53.600 21.200 55.200 ;
        RECT 9.200 49.700 13.200 50.300 ;
        RECT 9.200 48.800 10.000 49.700 ;
        RECT 12.400 42.200 13.200 49.700 ;
        RECT 14.000 48.800 14.800 50.400 ;
        RECT 17.400 50.200 18.000 53.600 ;
        RECT 18.800 50.800 19.600 52.400 ;
        RECT 20.400 52.300 21.200 52.400 ;
        RECT 22.000 52.300 22.800 55.800 ;
        RECT 23.600 54.300 24.400 54.400 ;
        RECT 26.800 54.300 27.600 54.400 ;
        RECT 23.600 53.700 27.600 54.300 ;
        RECT 23.600 53.600 24.400 53.700 ;
        RECT 26.800 53.600 27.600 53.700 ;
        RECT 27.000 53.200 27.600 53.600 ;
        RECT 27.000 52.400 27.800 53.200 ;
        RECT 28.400 52.400 29.000 55.800 ;
        RECT 33.200 55.600 34.000 57.200 ;
        RECT 30.000 52.800 30.800 54.400 ;
        RECT 20.400 51.700 22.800 52.300 ;
        RECT 20.400 51.600 21.200 51.700 ;
        RECT 17.200 49.400 19.000 50.200 ;
        RECT 18.200 44.400 19.000 49.400 ;
        RECT 17.200 43.600 19.000 44.400 ;
        RECT 18.200 42.200 19.000 43.600 ;
        RECT 22.000 42.200 22.800 51.700 ;
        RECT 25.200 50.800 26.000 52.400 ;
        RECT 28.400 51.600 29.200 52.400 ;
        RECT 31.600 52.200 32.400 52.400 ;
        RECT 30.800 51.600 32.400 52.200 ;
        RECT 34.800 52.300 35.600 59.800 ;
        RECT 39.000 55.800 40.600 59.800 ;
        RECT 36.400 54.300 37.200 54.400 ;
        RECT 38.000 54.300 38.800 54.400 ;
        RECT 36.400 53.700 38.800 54.300 ;
        RECT 36.400 53.600 37.200 53.700 ;
        RECT 38.000 53.600 38.800 53.700 ;
        RECT 38.200 53.200 38.800 53.600 ;
        RECT 38.200 52.400 39.000 53.200 ;
        RECT 39.600 52.400 40.200 55.800 ;
        RECT 41.200 52.800 42.000 54.400 ;
        RECT 45.600 54.200 46.400 59.800 ;
        RECT 50.800 55.800 51.600 59.800 ;
        RECT 52.400 56.000 53.200 59.800 ;
        RECT 55.600 56.000 56.400 59.800 ;
        RECT 52.400 55.800 56.400 56.000 ;
        RECT 51.000 54.400 51.600 55.800 ;
        RECT 52.600 55.400 56.200 55.800 ;
        RECT 57.200 55.600 58.000 57.200 ;
        RECT 54.800 54.400 55.600 54.800 ;
        RECT 44.600 53.800 46.400 54.200 ;
        RECT 44.600 53.600 46.200 53.800 ;
        RECT 50.800 53.600 53.400 54.400 ;
        RECT 54.800 54.300 56.400 54.400 ;
        RECT 57.300 54.300 57.900 55.600 ;
        RECT 54.800 53.800 57.900 54.300 ;
        RECT 55.600 53.700 57.900 53.800 ;
        RECT 55.600 53.600 56.400 53.700 ;
        RECT 36.400 52.300 37.200 52.400 ;
        RECT 34.800 51.700 37.200 52.300 ;
        RECT 28.400 51.400 29.000 51.600 ;
        RECT 27.000 50.800 29.000 51.400 ;
        RECT 30.800 51.200 31.600 51.600 ;
        RECT 23.600 48.800 24.400 50.400 ;
        RECT 27.000 50.200 27.600 50.800 ;
        RECT 25.200 42.800 26.000 50.200 ;
        RECT 26.800 43.400 27.600 50.200 ;
        RECT 28.400 49.600 32.400 50.200 ;
        RECT 28.400 42.800 29.200 49.600 ;
        RECT 25.200 42.200 29.200 42.800 ;
        RECT 31.600 42.200 32.400 49.600 ;
        RECT 34.800 42.200 35.600 51.700 ;
        RECT 36.400 50.800 37.200 51.700 ;
        RECT 39.600 51.600 40.400 52.400 ;
        RECT 42.800 52.200 43.600 52.400 ;
        RECT 42.000 51.600 43.600 52.200 ;
        RECT 39.600 51.400 40.200 51.600 ;
        RECT 38.200 50.800 40.200 51.400 ;
        RECT 42.000 51.200 42.800 51.600 ;
        RECT 38.200 50.200 38.800 50.800 ;
        RECT 44.600 50.400 45.200 53.600 ;
        RECT 46.800 51.600 48.400 52.400 ;
        RECT 36.400 42.800 37.200 50.200 ;
        RECT 38.000 43.400 38.800 50.200 ;
        RECT 39.600 49.600 43.600 50.200 ;
        RECT 44.400 49.600 45.200 50.400 ;
        RECT 49.200 49.600 50.000 51.200 ;
        RECT 50.800 50.200 51.600 50.400 ;
        RECT 52.800 50.200 53.400 53.600 ;
        RECT 54.000 51.600 54.800 53.200 ;
        RECT 50.800 49.600 52.200 50.200 ;
        RECT 52.800 49.600 53.800 50.200 ;
        RECT 39.600 42.800 40.400 49.600 ;
        RECT 36.400 42.200 40.400 42.800 ;
        RECT 42.800 42.200 43.600 49.600 ;
        RECT 44.600 47.000 45.200 49.600 ;
        RECT 46.000 47.600 46.800 49.200 ;
        RECT 51.600 48.400 52.200 49.600 ;
        RECT 51.600 47.600 52.400 48.400 ;
        RECT 44.600 46.400 48.200 47.000 ;
        RECT 44.600 46.200 45.200 46.400 ;
        RECT 44.400 42.200 45.200 46.200 ;
        RECT 47.600 46.200 48.200 46.400 ;
        RECT 47.600 42.200 48.400 46.200 ;
        RECT 53.000 42.200 53.800 49.600 ;
        RECT 58.800 42.200 59.600 59.800 ;
        RECT 60.400 55.600 61.200 57.200 ;
        RECT 62.000 42.200 62.800 59.800 ;
        RECT 63.800 56.400 64.600 57.200 ;
        RECT 63.600 55.600 64.400 56.400 ;
        RECT 65.200 55.800 66.000 59.800 ;
        RECT 73.800 56.000 74.600 59.000 ;
        RECT 78.000 57.000 78.800 59.000 ;
        RECT 63.600 52.200 64.400 52.400 ;
        RECT 65.400 52.200 66.000 55.800 ;
        RECT 73.000 55.400 74.600 56.000 ;
        RECT 73.000 55.000 73.800 55.400 ;
        RECT 73.000 54.400 73.600 55.000 ;
        RECT 78.200 54.800 78.800 57.000 ;
        RECT 79.600 56.000 80.400 59.800 ;
        RECT 82.800 56.000 83.600 59.800 ;
        RECT 79.600 55.800 83.600 56.000 ;
        RECT 84.400 55.800 85.200 59.800 ;
        RECT 86.600 58.400 87.400 59.800 ;
        RECT 86.000 57.600 87.400 58.400 ;
        RECT 86.600 56.400 87.400 57.600 ;
        RECT 91.400 56.400 92.200 59.800 ;
        RECT 96.200 56.400 97.000 59.800 ;
        RECT 86.600 55.800 88.400 56.400 ;
        RECT 91.400 55.800 93.200 56.400 ;
        RECT 96.200 55.800 98.000 56.400 ;
        RECT 100.400 56.000 101.200 59.800 ;
        RECT 103.600 56.000 104.400 59.800 ;
        RECT 100.400 55.800 104.400 56.000 ;
        RECT 105.200 55.800 106.000 59.800 ;
        RECT 79.800 55.400 83.400 55.800 ;
        RECT 66.800 52.800 67.600 54.400 ;
        RECT 71.600 53.600 73.600 54.400 ;
        RECT 74.600 54.200 78.800 54.800 ;
        RECT 80.400 54.400 81.200 54.800 ;
        RECT 84.400 54.400 85.000 55.800 ;
        RECT 74.600 53.800 75.600 54.200 ;
        RECT 68.400 52.300 69.200 52.400 ;
        RECT 71.600 52.300 72.400 52.400 ;
        RECT 68.400 52.200 72.400 52.300 ;
        RECT 63.600 51.600 66.000 52.200 ;
        RECT 67.600 51.700 72.400 52.200 ;
        RECT 67.600 51.600 69.200 51.700 ;
        RECT 63.800 50.200 64.400 51.600 ;
        RECT 67.600 51.200 68.400 51.600 ;
        RECT 71.600 50.800 72.400 51.700 ;
        RECT 63.600 42.200 64.400 50.200 ;
        RECT 65.200 49.600 69.200 50.200 ;
        RECT 65.200 42.200 66.000 49.600 ;
        RECT 68.400 42.200 69.200 49.600 ;
        RECT 73.000 49.800 73.600 53.600 ;
        RECT 74.200 53.000 75.600 53.800 ;
        RECT 79.600 53.800 81.200 54.400 ;
        RECT 79.600 53.600 80.400 53.800 ;
        RECT 82.600 53.600 85.200 54.400 ;
        RECT 75.000 51.000 75.600 53.000 ;
        RECT 76.400 51.600 77.200 53.200 ;
        RECT 78.000 51.600 78.800 53.200 ;
        RECT 81.200 51.600 82.000 53.200 ;
        RECT 75.000 50.400 78.800 51.000 ;
        RECT 73.000 49.200 74.600 49.800 ;
        RECT 73.800 44.400 74.600 49.200 ;
        RECT 78.200 47.000 78.800 50.400 ;
        RECT 82.600 50.200 83.200 53.600 ;
        RECT 84.400 50.200 85.200 50.400 ;
        RECT 73.200 43.600 74.600 44.400 ;
        RECT 73.800 42.200 74.600 43.600 ;
        RECT 78.000 43.000 78.800 47.000 ;
        RECT 82.200 49.600 83.200 50.200 ;
        RECT 83.800 49.600 85.200 50.200 ;
        RECT 82.200 44.400 83.000 49.600 ;
        RECT 83.800 48.400 84.400 49.600 ;
        RECT 86.000 48.800 86.800 50.400 ;
        RECT 83.600 47.600 84.400 48.400 ;
        RECT 81.200 43.600 83.000 44.400 ;
        RECT 82.200 42.200 83.000 43.600 ;
        RECT 87.600 42.200 88.400 55.800 ;
        RECT 89.200 53.600 90.000 55.200 ;
        RECT 90.800 48.800 91.600 50.400 ;
        RECT 92.400 42.200 93.200 55.800 ;
        RECT 94.000 54.300 94.800 55.200 ;
        RECT 97.200 54.300 98.000 55.800 ;
        RECT 100.600 55.400 104.200 55.800 ;
        RECT 94.000 53.700 98.000 54.300 ;
        RECT 94.000 53.600 94.800 53.700 ;
        RECT 95.600 48.800 96.400 50.400 ;
        RECT 97.200 42.200 98.000 53.700 ;
        RECT 98.800 54.300 99.600 55.200 ;
        RECT 101.200 54.400 102.000 54.800 ;
        RECT 105.200 54.400 105.800 55.800 ;
        RECT 106.800 55.600 107.600 57.200 ;
        RECT 100.400 54.300 102.000 54.400 ;
        RECT 98.800 53.800 102.000 54.300 ;
        RECT 98.800 53.700 101.200 53.800 ;
        RECT 98.800 53.600 99.600 53.700 ;
        RECT 100.400 53.600 101.200 53.700 ;
        RECT 103.400 53.600 106.000 54.400 ;
        RECT 108.400 54.300 109.200 59.800 ;
        RECT 110.000 56.000 110.800 59.800 ;
        RECT 113.200 56.000 114.000 59.800 ;
        RECT 110.000 55.800 114.000 56.000 ;
        RECT 114.800 55.800 115.600 59.800 ;
        RECT 118.000 57.800 118.800 59.800 ;
        RECT 110.200 55.400 113.800 55.800 ;
        RECT 110.800 54.400 111.600 54.800 ;
        RECT 114.800 54.400 115.400 55.800 ;
        RECT 116.400 55.600 117.200 57.200 ;
        RECT 118.200 54.400 118.800 57.800 ;
        RECT 110.000 54.300 111.600 54.400 ;
        RECT 108.400 53.800 111.600 54.300 ;
        RECT 108.400 53.700 110.800 53.800 ;
        RECT 102.000 51.600 102.800 53.200 ;
        RECT 103.400 50.200 104.000 53.600 ;
        RECT 105.200 50.200 106.000 50.400 ;
        RECT 103.000 49.600 104.000 50.200 ;
        RECT 104.600 49.600 106.000 50.200 ;
        RECT 103.000 44.400 103.800 49.600 ;
        RECT 104.600 48.400 105.200 49.600 ;
        RECT 104.400 47.600 105.200 48.400 ;
        RECT 102.000 43.600 103.800 44.400 ;
        RECT 103.000 42.200 103.800 43.600 ;
        RECT 108.400 42.200 109.200 53.700 ;
        RECT 110.000 53.600 110.800 53.700 ;
        RECT 113.000 53.600 115.600 54.400 ;
        RECT 118.000 53.600 118.800 54.400 ;
        RECT 111.600 51.600 112.400 53.200 ;
        RECT 113.000 50.200 113.600 53.600 ;
        RECT 118.200 52.400 118.800 53.600 ;
        RECT 118.000 51.600 118.800 52.400 ;
        RECT 114.800 50.200 115.600 50.400 ;
        RECT 118.200 50.200 118.800 51.600 ;
        RECT 119.600 52.300 120.400 52.400 ;
        RECT 121.200 52.300 122.000 59.800 ;
        RECT 122.800 55.600 123.600 57.200 ;
        RECT 124.400 55.800 125.200 59.800 ;
        RECT 126.000 56.000 126.800 59.800 ;
        RECT 129.200 56.000 130.000 59.800 ;
        RECT 126.000 55.800 130.000 56.000 ;
        RECT 124.600 54.400 125.200 55.800 ;
        RECT 126.200 55.400 129.800 55.800 ;
        RECT 128.400 54.400 129.200 54.800 ;
        RECT 124.400 53.600 127.000 54.400 ;
        RECT 128.400 53.800 130.000 54.400 ;
        RECT 129.200 53.600 130.000 53.800 ;
        RECT 119.600 51.700 122.000 52.300 ;
        RECT 119.600 50.800 120.400 51.700 ;
        RECT 112.600 49.600 113.600 50.200 ;
        RECT 114.200 49.600 115.600 50.200 ;
        RECT 112.600 42.200 113.400 49.600 ;
        RECT 114.200 48.400 114.800 49.600 ;
        RECT 118.000 49.400 119.800 50.200 ;
        RECT 114.000 47.600 114.800 48.400 ;
        RECT 119.000 42.200 119.800 49.400 ;
        RECT 121.200 42.200 122.000 51.700 ;
        RECT 124.400 50.200 125.200 50.400 ;
        RECT 126.400 50.200 127.000 53.600 ;
        RECT 127.600 51.600 128.400 53.200 ;
        RECT 124.400 49.600 125.800 50.200 ;
        RECT 126.400 49.600 127.400 50.200 ;
        RECT 125.200 48.400 125.800 49.600 ;
        RECT 125.200 47.600 126.000 48.400 ;
        RECT 126.600 42.200 127.400 49.600 ;
        RECT 130.800 42.200 131.600 59.800 ;
        RECT 132.400 55.600 133.200 57.200 ;
        RECT 138.800 56.000 139.600 59.800 ;
        RECT 142.000 56.000 142.800 59.800 ;
        RECT 138.800 55.800 142.800 56.000 ;
        RECT 143.600 55.800 144.400 59.800 ;
        RECT 132.500 54.300 133.100 55.600 ;
        RECT 139.000 55.400 142.600 55.800 ;
        RECT 139.600 54.400 140.400 54.800 ;
        RECT 143.600 54.400 144.200 55.800 ;
        RECT 138.800 54.300 140.400 54.400 ;
        RECT 132.500 53.800 140.400 54.300 ;
        RECT 132.500 53.700 139.600 53.800 ;
        RECT 138.800 53.600 139.600 53.700 ;
        RECT 141.800 53.600 144.400 54.400 ;
        RECT 140.400 51.600 141.200 53.200 ;
        RECT 141.800 50.200 142.400 53.600 ;
        RECT 143.600 50.300 144.400 50.400 ;
        RECT 145.200 50.300 146.000 59.800 ;
        RECT 146.800 56.300 147.600 57.200 ;
        RECT 148.600 56.400 149.400 57.200 ;
        RECT 148.400 56.300 149.200 56.400 ;
        RECT 146.800 55.700 149.200 56.300 ;
        RECT 150.000 55.800 150.800 59.800 ;
        RECT 146.800 55.600 147.600 55.700 ;
        RECT 148.400 55.600 149.200 55.700 ;
        RECT 148.400 52.200 149.200 52.400 ;
        RECT 150.200 52.200 150.800 55.800 ;
        RECT 154.800 55.800 155.600 59.800 ;
        RECT 159.200 56.200 160.800 59.800 ;
        RECT 154.800 55.200 157.200 55.800 ;
        RECT 156.400 55.000 157.200 55.200 ;
        RECT 157.800 54.800 158.600 55.600 ;
        RECT 157.800 54.400 158.400 54.800 ;
        RECT 151.600 52.800 152.400 54.400 ;
        RECT 153.200 54.300 154.000 54.400 ;
        RECT 154.800 54.300 156.400 54.400 ;
        RECT 153.200 53.700 156.400 54.300 ;
        RECT 153.200 53.600 154.000 53.700 ;
        RECT 154.800 53.600 156.400 53.700 ;
        RECT 157.600 53.600 158.400 54.400 ;
        RECT 159.200 54.200 159.800 56.200 ;
        RECT 164.400 55.800 165.200 59.800 ;
        RECT 160.400 54.800 162.000 55.600 ;
        RECT 162.600 55.200 165.200 55.800 ;
        RECT 166.000 55.800 166.800 59.800 ;
        RECT 170.400 56.200 172.000 59.800 ;
        RECT 166.000 55.200 168.400 55.800 ;
        RECT 162.600 55.000 163.400 55.200 ;
        RECT 167.600 55.000 168.400 55.200 ;
        RECT 169.000 54.800 169.800 55.600 ;
        RECT 169.000 54.400 169.600 54.800 ;
        RECT 163.600 54.200 165.200 54.400 ;
        RECT 159.200 53.600 160.200 54.200 ;
        RECT 163.000 54.000 165.200 54.200 ;
        RECT 159.600 52.400 160.200 53.600 ;
        RECT 160.800 53.600 165.200 54.000 ;
        RECT 166.000 53.600 167.600 54.400 ;
        RECT 168.800 53.600 169.600 54.400 ;
        RECT 160.800 53.400 163.600 53.600 ;
        RECT 160.800 53.200 161.600 53.400 ;
        RECT 170.400 52.800 171.000 56.200 ;
        RECT 175.600 55.800 176.400 59.800 ;
        RECT 171.600 55.400 173.200 55.600 ;
        RECT 171.600 54.800 173.600 55.400 ;
        RECT 174.200 55.200 176.400 55.800 ;
        RECT 174.200 55.000 175.000 55.200 ;
        RECT 177.200 55.000 178.000 59.800 ;
        RECT 181.600 58.400 182.400 59.800 ;
        RECT 180.400 57.800 182.400 58.400 ;
        RECT 186.000 57.800 186.800 59.800 ;
        RECT 190.200 58.400 191.400 59.800 ;
        RECT 190.000 57.800 191.400 58.400 ;
        RECT 180.400 57.000 181.200 57.800 ;
        RECT 186.000 57.200 186.600 57.800 ;
        RECT 182.000 56.400 182.800 57.200 ;
        RECT 183.800 56.600 186.600 57.200 ;
        RECT 190.000 57.000 190.800 57.800 ;
        RECT 183.800 56.400 184.600 56.600 ;
        RECT 173.000 54.400 173.600 54.800 ;
        RECT 171.600 53.400 172.400 54.200 ;
        RECT 173.000 53.800 176.400 54.400 ;
        RECT 174.800 53.600 176.400 53.800 ;
        RECT 178.000 54.200 179.600 54.400 ;
        RECT 182.200 54.200 182.800 56.400 ;
        RECT 191.800 55.400 192.600 55.600 ;
        RECT 194.800 55.400 195.600 59.800 ;
        RECT 191.800 54.800 195.600 55.400 ;
        RECT 187.800 54.200 188.600 54.400 ;
        RECT 178.000 53.600 189.000 54.200 ;
        RECT 181.000 53.400 181.800 53.600 ;
        RECT 170.000 52.400 171.000 52.800 ;
        RECT 153.200 52.300 154.000 52.400 ;
        RECT 159.600 52.300 160.400 52.400 ;
        RECT 153.200 52.200 160.400 52.300 ;
        RECT 162.200 52.200 163.000 52.400 ;
        RECT 148.400 51.600 150.800 52.200 ;
        RECT 152.400 51.700 160.400 52.200 ;
        RECT 152.400 51.600 154.000 51.700 ;
        RECT 159.600 51.600 160.400 51.700 ;
        RECT 161.400 51.600 163.000 52.200 ;
        RECT 169.200 52.200 171.000 52.400 ;
        RECT 171.800 52.800 172.400 53.400 ;
        RECT 171.800 52.200 174.400 52.800 ;
        RECT 169.200 51.600 170.600 52.200 ;
        RECT 173.600 52.000 174.400 52.200 ;
        RECT 179.400 52.400 180.200 52.600 ;
        RECT 182.000 52.400 182.800 52.600 ;
        RECT 179.400 51.800 184.400 52.400 ;
        RECT 183.600 51.600 184.400 51.800 ;
        RECT 143.600 50.200 146.000 50.300 ;
        RECT 148.600 50.200 149.200 51.600 ;
        RECT 152.400 51.200 153.200 51.600 ;
        RECT 159.600 50.200 160.200 51.600 ;
        RECT 161.400 51.400 162.200 51.600 ;
        RECT 170.000 50.200 170.600 51.600 ;
        RECT 171.400 51.400 172.200 51.600 ;
        RECT 171.400 50.800 174.800 51.400 ;
        RECT 174.200 50.200 174.800 50.800 ;
        RECT 177.200 51.000 182.800 51.200 ;
        RECT 177.200 50.800 183.000 51.000 ;
        RECT 177.200 50.600 187.000 50.800 ;
        RECT 141.400 49.600 142.400 50.200 ;
        RECT 143.000 49.700 146.000 50.200 ;
        RECT 143.000 49.600 144.400 49.700 ;
        RECT 141.400 42.200 142.200 49.600 ;
        RECT 143.000 48.400 143.600 49.600 ;
        RECT 142.800 47.600 143.600 48.400 ;
        RECT 145.200 42.200 146.000 49.700 ;
        RECT 148.400 42.200 149.200 50.200 ;
        RECT 150.000 49.600 154.000 50.200 ;
        RECT 150.000 42.200 150.800 49.600 ;
        RECT 153.200 42.200 154.000 49.600 ;
        RECT 154.800 49.600 157.200 50.200 ;
        RECT 154.800 42.200 155.600 49.600 ;
        RECT 156.400 49.400 157.200 49.600 ;
        RECT 159.200 44.400 160.800 50.200 ;
        RECT 162.600 49.600 165.200 50.200 ;
        RECT 162.600 49.400 163.400 49.600 ;
        RECT 158.000 43.600 160.800 44.400 ;
        RECT 159.200 42.200 160.800 43.600 ;
        RECT 164.400 42.200 165.200 49.600 ;
        RECT 166.000 49.600 168.400 50.200 ;
        RECT 170.000 49.600 172.000 50.200 ;
        RECT 166.000 42.200 166.800 49.600 ;
        RECT 167.600 49.400 168.400 49.600 ;
        RECT 170.400 48.400 172.000 49.600 ;
        RECT 174.200 49.600 176.400 50.200 ;
        RECT 174.200 49.400 175.000 49.600 ;
        RECT 170.400 47.600 173.200 48.400 ;
        RECT 170.400 42.200 172.000 47.600 ;
        RECT 175.600 42.200 176.400 49.600 ;
        RECT 177.200 42.200 178.000 50.600 ;
        RECT 182.200 50.200 187.000 50.600 ;
        RECT 180.400 49.000 185.800 49.600 ;
        RECT 180.400 48.800 181.200 49.000 ;
        RECT 185.000 48.800 185.800 49.000 ;
        RECT 186.400 49.000 187.000 50.200 ;
        RECT 188.400 50.400 189.000 53.600 ;
        RECT 190.000 52.800 190.800 53.000 ;
        RECT 190.000 52.200 193.800 52.800 ;
        RECT 193.000 52.000 193.800 52.200 ;
        RECT 191.400 51.400 192.200 51.600 ;
        RECT 194.800 51.400 195.600 54.800 ;
        RECT 191.400 50.800 195.600 51.400 ;
        RECT 188.400 49.800 190.800 50.400 ;
        RECT 187.800 49.000 188.600 49.200 ;
        RECT 186.400 48.400 188.600 49.000 ;
        RECT 190.200 48.800 190.800 49.800 ;
        RECT 190.200 48.000 191.600 48.800 ;
        RECT 183.800 47.400 184.600 47.600 ;
        RECT 186.600 47.400 187.400 47.600 ;
        RECT 180.400 46.200 181.200 47.000 ;
        RECT 183.800 46.800 187.400 47.400 ;
        RECT 186.000 46.200 186.600 46.800 ;
        RECT 190.000 46.200 190.800 47.000 ;
        RECT 180.400 45.600 182.400 46.200 ;
        RECT 181.600 42.200 182.400 45.600 ;
        RECT 186.000 42.200 186.800 46.200 ;
        RECT 190.200 42.200 191.400 46.200 ;
        RECT 194.800 42.200 195.600 50.800 ;
        RECT 196.400 42.200 197.200 59.800 ;
        RECT 199.600 55.800 200.400 59.800 ;
        RECT 204.000 58.400 205.600 59.800 ;
        RECT 204.000 57.600 206.800 58.400 ;
        RECT 204.000 56.200 205.600 57.600 ;
        RECT 199.600 55.200 202.000 55.800 ;
        RECT 198.000 53.600 198.800 55.200 ;
        RECT 201.200 55.000 202.000 55.200 ;
        RECT 202.600 54.800 203.400 55.600 ;
        RECT 202.600 54.400 203.200 54.800 ;
        RECT 199.600 53.600 201.200 54.400 ;
        RECT 202.400 53.600 203.200 54.400 ;
        RECT 204.000 54.200 204.600 56.200 ;
        RECT 209.200 55.800 210.000 59.800 ;
        RECT 210.800 55.800 211.600 59.800 ;
        RECT 212.400 56.000 213.200 59.800 ;
        RECT 215.600 56.000 216.400 59.800 ;
        RECT 212.400 55.800 216.400 56.000 ;
        RECT 205.200 54.800 206.800 55.600 ;
        RECT 207.400 55.200 210.000 55.800 ;
        RECT 207.400 55.000 208.200 55.200 ;
        RECT 211.000 54.400 211.600 55.800 ;
        RECT 212.600 55.400 216.200 55.800 ;
        RECT 214.800 54.400 215.600 54.800 ;
        RECT 208.400 54.200 210.000 54.400 ;
        RECT 204.000 53.600 205.000 54.200 ;
        RECT 207.800 54.000 210.000 54.200 ;
        RECT 204.400 52.400 205.000 53.600 ;
        RECT 205.600 53.600 210.000 54.000 ;
        RECT 210.800 53.600 213.400 54.400 ;
        RECT 214.800 53.800 216.400 54.400 ;
        RECT 215.600 53.600 216.400 53.800 ;
        RECT 217.200 53.600 218.000 55.200 ;
        RECT 205.600 53.400 208.400 53.600 ;
        RECT 205.600 53.200 206.400 53.400 ;
        RECT 204.400 51.600 205.200 52.400 ;
        RECT 207.000 52.200 207.800 52.400 ;
        RECT 206.200 51.600 207.800 52.200 ;
        RECT 204.400 50.200 205.000 51.600 ;
        RECT 206.200 51.400 207.000 51.600 ;
        RECT 210.800 50.200 211.600 50.400 ;
        RECT 212.800 50.200 213.400 53.600 ;
        RECT 214.000 52.300 214.800 53.200 ;
        RECT 218.800 52.300 219.600 59.800 ;
        RECT 222.000 57.600 222.800 59.800 ;
        RECT 226.800 57.600 227.600 59.800 ;
        RECT 231.600 57.800 232.400 59.800 ;
        RECT 222.000 54.400 222.600 57.600 ;
        RECT 223.600 55.600 224.400 57.200 ;
        RECT 226.800 54.400 227.400 57.600 ;
        RECT 228.400 55.600 229.200 57.200 ;
        RECT 230.000 55.600 230.800 57.200 ;
        RECT 222.000 53.600 222.800 54.400 ;
        RECT 226.800 53.600 227.600 54.400 ;
        RECT 228.500 54.300 229.100 55.600 ;
        RECT 231.800 54.400 232.400 57.800 ;
        RECT 234.800 56.000 235.600 59.800 ;
        RECT 238.000 56.000 238.800 59.800 ;
        RECT 234.800 55.800 238.800 56.000 ;
        RECT 239.600 55.800 240.400 59.800 ;
        RECT 241.200 55.800 242.000 59.800 ;
        RECT 245.600 58.400 247.200 59.800 ;
        RECT 245.600 57.600 248.400 58.400 ;
        RECT 245.600 56.200 247.200 57.600 ;
        RECT 235.000 55.400 238.600 55.800 ;
        RECT 235.600 54.400 236.400 54.800 ;
        RECT 239.600 54.400 240.200 55.800 ;
        RECT 241.200 55.200 243.400 55.800 ;
        RECT 244.400 55.400 246.000 55.600 ;
        RECT 242.600 55.000 243.400 55.200 ;
        RECT 244.000 54.800 246.000 55.400 ;
        RECT 244.000 54.400 244.600 54.800 ;
        RECT 231.600 54.300 232.400 54.400 ;
        RECT 228.500 53.700 232.400 54.300 ;
        RECT 231.600 53.600 232.400 53.700 ;
        RECT 234.800 53.800 236.400 54.400 ;
        RECT 234.800 53.600 235.600 53.800 ;
        RECT 237.800 53.600 240.400 54.400 ;
        RECT 241.200 53.800 244.600 54.400 ;
        RECT 241.200 53.600 242.800 53.800 ;
        RECT 220.400 52.300 221.200 52.400 ;
        RECT 214.000 51.700 221.200 52.300 ;
        RECT 214.000 51.600 214.800 51.700 ;
        RECT 199.600 49.600 202.000 50.200 ;
        RECT 199.600 42.200 200.400 49.600 ;
        RECT 201.200 49.400 202.000 49.600 ;
        RECT 204.000 42.200 205.600 50.200 ;
        RECT 207.400 49.600 210.000 50.200 ;
        RECT 210.800 49.600 212.200 50.200 ;
        RECT 212.800 49.600 213.800 50.200 ;
        RECT 207.400 49.400 208.200 49.600 ;
        RECT 209.200 42.200 210.000 49.600 ;
        RECT 211.600 48.400 212.200 49.600 ;
        RECT 211.600 47.600 212.400 48.400 ;
        RECT 213.000 42.200 213.800 49.600 ;
        RECT 218.800 42.200 219.600 51.700 ;
        RECT 220.400 50.800 221.200 51.700 ;
        RECT 222.000 52.300 222.600 53.600 ;
        RECT 225.200 52.300 226.000 52.400 ;
        RECT 222.000 51.700 226.000 52.300 ;
        RECT 222.000 50.200 222.600 51.700 ;
        RECT 225.200 50.800 226.000 51.700 ;
        RECT 226.800 50.200 227.400 53.600 ;
        RECT 231.800 50.200 232.400 53.600 ;
        RECT 233.200 52.300 234.000 52.400 ;
        RECT 236.400 52.300 237.200 53.200 ;
        RECT 233.200 51.700 237.200 52.300 ;
        RECT 233.200 50.800 234.000 51.700 ;
        RECT 236.400 51.600 237.200 51.700 ;
        RECT 237.800 50.400 238.400 53.600 ;
        RECT 245.200 53.400 246.000 54.200 ;
        RECT 245.200 52.800 245.800 53.400 ;
        RECT 243.200 52.200 245.800 52.800 ;
        RECT 246.600 52.800 247.200 56.200 ;
        RECT 250.800 55.800 251.600 59.800 ;
        RECT 247.800 54.800 248.600 55.600 ;
        RECT 249.200 55.200 251.600 55.800 ;
        RECT 252.400 55.200 253.200 59.800 ;
        RECT 255.600 56.400 256.400 59.800 ;
        RECT 255.600 55.800 256.600 56.400 ;
        RECT 249.200 55.000 250.000 55.200 ;
        RECT 248.000 54.400 248.600 54.800 ;
        RECT 252.400 54.600 255.000 55.200 ;
        RECT 248.000 53.600 248.800 54.400 ;
        RECT 250.000 53.600 251.600 54.400 ;
        RECT 246.600 52.400 247.600 52.800 ;
        RECT 252.600 52.400 253.400 53.200 ;
        RECT 246.600 52.200 248.400 52.400 ;
        RECT 243.200 52.000 244.000 52.200 ;
        RECT 247.000 51.600 248.400 52.200 ;
        RECT 252.400 51.600 253.400 52.400 ;
        RECT 254.400 53.000 255.000 54.600 ;
        RECT 256.000 54.400 256.600 55.800 ;
        RECT 258.800 55.200 259.600 59.800 ;
        RECT 258.800 54.600 261.000 55.200 ;
        RECT 255.600 53.600 256.600 54.400 ;
        RECT 254.400 52.200 255.400 53.000 ;
        RECT 245.400 51.400 246.200 51.600 ;
        RECT 242.800 50.800 246.200 51.400 ;
        RECT 221.000 49.400 222.800 50.200 ;
        RECT 225.800 49.400 227.600 50.200 ;
        RECT 231.600 49.400 233.400 50.200 ;
        RECT 236.400 49.600 238.400 50.400 ;
        RECT 239.600 50.200 240.400 50.400 ;
        RECT 242.800 50.200 243.400 50.800 ;
        RECT 247.000 50.200 247.600 51.600 ;
        RECT 254.400 50.200 255.000 52.200 ;
        RECT 256.000 50.200 256.600 53.600 ;
        RECT 258.800 51.600 259.600 53.200 ;
        RECT 260.400 51.600 261.000 54.600 ;
        RECT 262.000 52.400 262.800 59.800 ;
        RECT 263.600 55.200 264.400 59.800 ;
        RECT 266.800 56.400 267.600 59.800 ;
        RECT 266.800 55.800 267.800 56.400 ;
        RECT 263.600 54.600 266.200 55.200 ;
        RECT 263.800 52.400 264.600 53.200 ;
        RECT 260.400 50.800 261.600 51.600 ;
        RECT 260.400 50.200 261.000 50.800 ;
        RECT 262.200 50.200 262.800 52.400 ;
        RECT 263.600 51.600 264.600 52.400 ;
        RECT 265.600 53.000 266.200 54.600 ;
        RECT 267.200 54.400 267.800 55.800 ;
        RECT 266.800 53.600 267.800 54.400 ;
        RECT 265.600 52.200 266.600 53.000 ;
        RECT 265.600 50.200 266.200 52.200 ;
        RECT 267.200 50.200 267.800 53.600 ;
        RECT 239.000 49.600 240.400 50.200 ;
        RECT 241.200 49.600 243.400 50.200 ;
        RECT 221.000 42.200 221.800 49.400 ;
        RECT 225.800 42.200 226.600 49.400 ;
        RECT 232.600 42.200 233.400 49.400 ;
        RECT 237.400 42.200 238.200 49.600 ;
        RECT 239.000 48.400 239.600 49.600 ;
        RECT 238.800 47.600 239.600 48.400 ;
        RECT 241.200 42.200 242.000 49.600 ;
        RECT 242.600 49.400 243.400 49.600 ;
        RECT 245.600 49.600 247.600 50.200 ;
        RECT 249.200 49.600 251.600 50.200 ;
        RECT 245.600 42.200 247.200 49.600 ;
        RECT 249.200 49.400 250.000 49.600 ;
        RECT 250.800 42.200 251.600 49.600 ;
        RECT 252.400 49.600 255.000 50.200 ;
        RECT 252.400 42.200 253.200 49.600 ;
        RECT 255.600 49.200 256.600 50.200 ;
        RECT 258.800 49.600 261.000 50.200 ;
        RECT 255.600 42.200 256.400 49.200 ;
        RECT 258.800 42.200 259.600 49.600 ;
        RECT 262.000 42.200 262.800 50.200 ;
        RECT 263.600 49.600 266.200 50.200 ;
        RECT 263.600 42.200 264.400 49.600 ;
        RECT 266.800 49.200 267.800 50.200 ;
        RECT 270.000 52.400 270.800 59.800 ;
        RECT 273.200 55.200 274.000 59.800 ;
        RECT 271.800 54.600 274.000 55.200 ;
        RECT 270.000 50.200 270.600 52.400 ;
        RECT 271.800 51.600 272.400 54.600 ;
        RECT 273.200 51.600 274.000 53.200 ;
        RECT 274.800 52.300 275.600 59.800 ;
        RECT 279.600 57.600 280.400 59.800 ;
        RECT 284.400 57.600 285.200 59.800 ;
        RECT 276.400 54.300 277.200 55.200 ;
        RECT 279.600 54.400 280.200 57.600 ;
        RECT 281.200 56.300 282.000 57.200 ;
        RECT 282.800 56.300 283.600 56.400 ;
        RECT 281.200 55.700 283.600 56.300 ;
        RECT 281.200 55.600 282.000 55.700 ;
        RECT 282.800 55.600 283.600 55.700 ;
        RECT 284.400 54.400 285.000 57.600 ;
        RECT 286.000 55.600 286.800 57.200 ;
        RECT 292.400 56.000 293.200 59.800 ;
        RECT 295.600 56.000 296.400 59.800 ;
        RECT 292.400 55.800 296.400 56.000 ;
        RECT 297.200 56.300 298.000 59.800 ;
        RECT 299.000 56.400 299.800 57.200 ;
        RECT 298.800 56.300 299.600 56.400 ;
        RECT 292.600 55.400 296.200 55.800 ;
        RECT 297.200 55.700 299.600 56.300 ;
        RECT 293.200 54.400 294.000 54.800 ;
        RECT 297.200 54.400 297.800 55.700 ;
        RECT 298.800 55.600 299.600 55.700 ;
        RECT 300.400 55.600 301.200 59.800 ;
        RECT 307.800 56.400 308.600 59.800 ;
        RECT 278.000 54.300 278.800 54.400 ;
        RECT 276.400 53.700 278.800 54.300 ;
        RECT 276.400 53.600 277.200 53.700 ;
        RECT 278.000 53.600 278.800 53.700 ;
        RECT 279.600 53.600 280.400 54.400 ;
        RECT 284.400 53.600 285.200 54.400 ;
        RECT 292.400 53.800 294.000 54.400 ;
        RECT 292.400 53.600 293.200 53.800 ;
        RECT 295.400 53.600 298.000 54.400 ;
        RECT 276.400 52.300 277.200 52.400 ;
        RECT 274.800 51.700 277.200 52.300 ;
        RECT 271.200 50.800 272.400 51.600 ;
        RECT 271.800 50.200 272.400 50.800 ;
        RECT 266.800 42.200 267.600 49.200 ;
        RECT 270.000 42.200 270.800 50.200 ;
        RECT 271.800 49.600 274.000 50.200 ;
        RECT 273.200 42.200 274.000 49.600 ;
        RECT 274.800 42.200 275.600 51.700 ;
        RECT 276.400 51.600 277.200 51.700 ;
        RECT 278.000 50.800 278.800 52.400 ;
        RECT 279.600 50.200 280.200 53.600 ;
        RECT 282.800 50.800 283.600 52.400 ;
        RECT 284.400 50.200 285.000 53.600 ;
        RECT 294.000 51.600 294.800 53.200 ;
        RECT 295.400 50.200 296.000 53.600 ;
        RECT 298.800 52.200 299.600 52.400 ;
        RECT 300.600 52.200 301.200 55.600 ;
        RECT 306.800 55.800 308.600 56.400 ;
        RECT 302.000 54.300 302.800 54.400 ;
        RECT 303.600 54.300 304.400 54.400 ;
        RECT 302.000 53.700 304.400 54.300 ;
        RECT 302.000 52.800 302.800 53.700 ;
        RECT 303.600 53.600 304.400 53.700 ;
        RECT 305.200 53.600 306.000 55.200 ;
        RECT 306.800 54.300 307.600 55.800 ;
        RECT 308.400 54.300 309.200 54.400 ;
        RECT 306.800 53.700 309.200 54.300 ;
        RECT 303.600 52.300 304.400 52.400 ;
        RECT 305.200 52.300 306.000 52.400 ;
        RECT 303.600 52.200 306.000 52.300 ;
        RECT 298.800 51.600 301.200 52.200 ;
        RECT 302.800 51.700 306.000 52.200 ;
        RECT 302.800 51.600 304.400 51.700 ;
        RECT 305.200 51.600 306.000 51.700 ;
        RECT 297.200 50.200 298.000 50.400 ;
        RECT 299.000 50.200 299.600 51.600 ;
        RECT 302.800 51.200 303.600 51.600 ;
        RECT 278.600 49.400 280.400 50.200 ;
        RECT 283.400 49.400 285.200 50.200 ;
        RECT 295.000 49.600 296.000 50.200 ;
        RECT 296.600 49.600 298.000 50.200 ;
        RECT 278.600 42.200 279.400 49.400 ;
        RECT 283.400 42.200 284.200 49.400 ;
        RECT 295.000 42.200 295.800 49.600 ;
        RECT 296.600 48.400 297.200 49.600 ;
        RECT 296.400 47.600 297.200 48.400 ;
        RECT 298.800 42.200 299.600 50.200 ;
        RECT 300.400 49.600 304.400 50.200 ;
        RECT 300.400 42.200 301.200 49.600 ;
        RECT 303.600 42.200 304.400 49.600 ;
        RECT 306.800 42.200 307.600 53.700 ;
        RECT 308.400 53.600 309.200 53.700 ;
        RECT 308.400 50.300 309.200 50.400 ;
        RECT 310.000 50.300 310.800 59.800 ;
        RECT 311.600 55.600 312.400 57.200 ;
        RECT 316.200 55.800 317.800 59.800 ;
        RECT 324.200 55.800 325.800 59.800 ;
        RECT 330.800 57.800 331.600 59.800 ;
        RECT 316.400 55.600 317.200 55.800 ;
        RECT 314.800 52.800 315.600 54.400 ;
        RECT 316.600 52.400 317.200 55.600 ;
        RECT 318.000 53.600 318.800 54.400 ;
        RECT 318.000 53.200 318.600 53.600 ;
        RECT 317.800 52.400 318.600 53.200 ;
        RECT 322.800 52.800 323.600 54.400 ;
        RECT 324.600 52.400 325.200 55.800 ;
        RECT 330.800 54.400 331.400 57.800 ;
        RECT 332.400 55.600 333.200 57.200 ;
        RECT 334.000 55.200 334.800 59.800 ;
        RECT 334.000 54.600 336.200 55.200 ;
        RECT 326.000 53.600 326.800 54.400 ;
        RECT 330.800 53.600 331.600 54.400 ;
        RECT 326.000 53.200 326.600 53.600 ;
        RECT 325.800 52.400 326.600 53.200 ;
        RECT 313.200 52.200 314.000 52.400 ;
        RECT 313.200 51.600 314.800 52.200 ;
        RECT 316.400 51.600 317.200 52.400 ;
        RECT 314.000 51.200 314.800 51.600 ;
        RECT 316.600 51.400 317.200 51.600 ;
        RECT 316.600 50.800 318.600 51.400 ;
        RECT 319.600 50.800 320.400 52.400 ;
        RECT 321.200 52.200 322.000 52.400 ;
        RECT 321.200 51.600 322.800 52.200 ;
        RECT 324.400 51.600 325.200 52.400 ;
        RECT 322.000 51.200 322.800 51.600 ;
        RECT 324.600 51.400 325.200 51.600 ;
        RECT 324.600 50.800 326.600 51.400 ;
        RECT 327.600 50.800 328.400 52.400 ;
        RECT 329.200 50.800 330.000 52.400 ;
        RECT 330.800 52.300 331.400 53.600 ;
        RECT 332.400 52.300 333.200 52.400 ;
        RECT 330.800 51.700 333.200 52.300 ;
        RECT 308.400 49.700 310.800 50.300 ;
        RECT 318.000 50.200 318.600 50.800 ;
        RECT 326.000 50.200 326.600 50.800 ;
        RECT 330.800 50.200 331.400 51.700 ;
        RECT 332.400 51.600 333.200 51.700 ;
        RECT 334.000 51.600 334.800 53.200 ;
        RECT 335.600 51.600 336.200 54.600 ;
        RECT 337.200 52.400 338.000 59.800 ;
        RECT 338.800 56.000 339.600 59.800 ;
        RECT 342.000 56.000 342.800 59.800 ;
        RECT 338.800 55.800 342.800 56.000 ;
        RECT 343.600 55.800 344.400 59.800 ;
        RECT 345.200 55.800 346.000 59.800 ;
        RECT 346.800 56.000 347.600 59.800 ;
        RECT 350.000 56.000 350.800 59.800 ;
        RECT 346.800 55.800 350.800 56.000 ;
        RECT 339.000 55.400 342.600 55.800 ;
        RECT 339.600 54.400 340.400 54.800 ;
        RECT 343.600 54.400 344.200 55.800 ;
        RECT 345.400 54.400 346.000 55.800 ;
        RECT 347.000 55.400 350.600 55.800 ;
        RECT 351.600 55.000 352.400 59.800 ;
        RECT 356.000 58.400 356.800 59.800 ;
        RECT 354.800 57.800 356.800 58.400 ;
        RECT 360.400 57.800 361.200 59.800 ;
        RECT 364.600 58.400 365.800 59.800 ;
        RECT 364.400 57.800 365.800 58.400 ;
        RECT 354.800 57.000 355.600 57.800 ;
        RECT 360.400 57.200 361.000 57.800 ;
        RECT 356.400 56.400 357.200 57.200 ;
        RECT 358.200 56.600 361.000 57.200 ;
        RECT 364.400 57.000 365.200 57.800 ;
        RECT 358.200 56.400 359.000 56.600 ;
        RECT 349.200 54.400 350.000 54.800 ;
        RECT 338.800 53.800 340.400 54.400 ;
        RECT 338.800 53.600 339.600 53.800 ;
        RECT 341.800 53.600 344.400 54.400 ;
        RECT 345.200 53.600 347.800 54.400 ;
        RECT 349.200 53.800 350.800 54.400 ;
        RECT 350.000 53.600 350.800 53.800 ;
        RECT 352.400 54.200 354.000 54.400 ;
        RECT 356.600 54.200 357.200 56.400 ;
        RECT 366.200 55.400 367.000 55.600 ;
        RECT 369.200 55.400 370.000 59.800 ;
        RECT 366.200 54.800 370.000 55.400 ;
        RECT 370.800 55.000 371.600 59.800 ;
        RECT 375.200 58.400 376.000 59.800 ;
        RECT 374.000 57.800 376.000 58.400 ;
        RECT 379.600 57.800 380.400 59.800 ;
        RECT 383.800 58.400 385.000 59.800 ;
        RECT 383.600 57.800 385.000 58.400 ;
        RECT 374.000 57.000 374.800 57.800 ;
        RECT 379.600 57.200 380.200 57.800 ;
        RECT 375.600 56.400 376.400 57.200 ;
        RECT 377.400 56.600 380.200 57.200 ;
        RECT 383.600 57.000 384.400 57.800 ;
        RECT 377.400 56.400 378.200 56.600 ;
        RECT 362.200 54.200 363.000 54.400 ;
        RECT 352.400 53.600 363.400 54.200 ;
        RECT 335.600 50.800 336.800 51.600 ;
        RECT 335.600 50.200 336.200 50.800 ;
        RECT 337.400 50.200 338.000 52.400 ;
        RECT 340.400 51.600 341.200 53.200 ;
        RECT 341.800 52.300 342.400 53.600 ;
        RECT 347.200 52.400 347.800 53.600 ;
        RECT 355.400 53.400 356.200 53.600 ;
        RECT 341.800 51.700 345.900 52.300 ;
        RECT 341.800 50.200 342.400 51.700 ;
        RECT 345.300 50.400 345.900 51.700 ;
        RECT 346.800 51.600 347.800 52.400 ;
        RECT 348.400 51.600 349.200 53.200 ;
        RECT 353.800 52.400 354.600 52.600 ;
        RECT 356.400 52.400 357.200 52.600 ;
        RECT 353.800 51.800 358.800 52.400 ;
        RECT 358.000 51.600 358.800 51.800 ;
        RECT 343.600 50.200 344.400 50.400 ;
        RECT 308.400 47.600 309.200 49.700 ;
        RECT 310.000 42.200 310.800 49.700 ;
        RECT 313.200 49.600 317.200 50.200 ;
        RECT 313.200 42.200 314.000 49.600 ;
        RECT 316.400 42.800 317.200 49.600 ;
        RECT 318.000 43.400 318.800 50.200 ;
        RECT 319.600 42.800 320.400 50.200 ;
        RECT 316.400 42.200 320.400 42.800 ;
        RECT 321.200 49.600 325.200 50.200 ;
        RECT 321.200 42.200 322.000 49.600 ;
        RECT 324.400 42.800 325.200 49.600 ;
        RECT 326.000 43.400 326.800 50.200 ;
        RECT 327.600 42.800 328.400 50.200 ;
        RECT 324.400 42.200 328.400 42.800 ;
        RECT 329.800 49.400 331.600 50.200 ;
        RECT 334.000 49.600 336.200 50.200 ;
        RECT 329.800 42.200 330.600 49.400 ;
        RECT 334.000 42.200 334.800 49.600 ;
        RECT 337.200 42.200 338.000 50.200 ;
        RECT 341.400 49.600 342.400 50.200 ;
        RECT 343.000 49.600 344.400 50.200 ;
        RECT 345.200 50.200 346.000 50.400 ;
        RECT 347.200 50.200 347.800 51.600 ;
        RECT 351.600 51.000 357.200 51.200 ;
        RECT 351.600 50.800 357.400 51.000 ;
        RECT 351.600 50.600 361.400 50.800 ;
        RECT 345.200 49.600 346.600 50.200 ;
        RECT 347.200 49.600 348.200 50.200 ;
        RECT 341.400 42.200 342.200 49.600 ;
        RECT 343.000 48.400 343.600 49.600 ;
        RECT 342.800 47.600 343.600 48.400 ;
        RECT 346.000 48.400 346.600 49.600 ;
        RECT 346.000 47.600 346.800 48.400 ;
        RECT 347.400 42.200 348.200 49.600 ;
        RECT 351.600 42.200 352.400 50.600 ;
        RECT 356.600 50.200 361.400 50.600 ;
        RECT 354.800 49.000 360.200 49.600 ;
        RECT 354.800 48.800 355.600 49.000 ;
        RECT 359.400 48.800 360.200 49.000 ;
        RECT 360.800 49.000 361.400 50.200 ;
        RECT 362.800 50.400 363.400 53.600 ;
        RECT 364.400 52.800 365.200 53.000 ;
        RECT 364.400 52.200 368.200 52.800 ;
        RECT 367.400 52.000 368.200 52.200 ;
        RECT 365.800 51.400 366.600 51.600 ;
        RECT 369.200 51.400 370.000 54.800 ;
        RECT 371.600 54.200 373.200 54.400 ;
        RECT 375.800 54.200 376.400 56.400 ;
        RECT 385.400 55.400 386.200 55.600 ;
        RECT 388.400 55.400 389.200 59.800 ;
        RECT 390.000 55.600 390.800 57.200 ;
        RECT 385.400 54.800 389.200 55.400 ;
        RECT 381.400 54.200 382.200 54.400 ;
        RECT 371.600 53.600 382.600 54.200 ;
        RECT 374.600 53.400 375.400 53.600 ;
        RECT 373.000 52.400 373.800 52.600 ;
        RECT 375.600 52.400 376.400 52.600 ;
        RECT 373.000 51.800 378.000 52.400 ;
        RECT 377.200 51.600 378.000 51.800 ;
        RECT 365.800 50.800 370.000 51.400 ;
        RECT 362.800 49.800 365.200 50.400 ;
        RECT 362.200 49.000 363.000 49.200 ;
        RECT 360.800 48.400 363.000 49.000 ;
        RECT 364.600 48.800 365.200 49.800 ;
        RECT 364.600 48.000 366.000 48.800 ;
        RECT 358.200 47.400 359.000 47.600 ;
        RECT 361.000 47.400 361.800 47.600 ;
        RECT 354.800 46.200 355.600 47.000 ;
        RECT 358.200 46.800 361.800 47.400 ;
        RECT 360.400 46.200 361.000 46.800 ;
        RECT 364.400 46.200 365.200 47.000 ;
        RECT 354.800 45.600 356.800 46.200 ;
        RECT 356.000 42.200 356.800 45.600 ;
        RECT 360.400 42.200 361.200 46.200 ;
        RECT 364.600 42.200 365.800 46.200 ;
        RECT 369.200 42.200 370.000 50.800 ;
        RECT 370.800 51.000 376.400 51.200 ;
        RECT 370.800 50.800 376.600 51.000 ;
        RECT 370.800 50.600 380.600 50.800 ;
        RECT 370.800 42.200 371.600 50.600 ;
        RECT 375.800 50.200 380.600 50.600 ;
        RECT 374.000 49.000 379.400 49.600 ;
        RECT 374.000 48.800 374.800 49.000 ;
        RECT 378.600 48.800 379.400 49.000 ;
        RECT 380.000 49.000 380.600 50.200 ;
        RECT 382.000 50.400 382.600 53.600 ;
        RECT 383.600 52.800 384.400 53.000 ;
        RECT 383.600 52.200 387.400 52.800 ;
        RECT 386.600 52.000 387.400 52.200 ;
        RECT 385.000 51.400 385.800 51.600 ;
        RECT 388.400 51.400 389.200 54.800 ;
        RECT 385.000 50.800 389.200 51.400 ;
        RECT 382.000 49.800 384.400 50.400 ;
        RECT 381.400 49.000 382.200 49.200 ;
        RECT 380.000 48.400 382.200 49.000 ;
        RECT 383.800 48.800 384.400 49.800 ;
        RECT 383.800 48.400 385.200 48.800 ;
        RECT 383.800 48.000 386.000 48.400 ;
        RECT 384.600 47.600 386.000 48.000 ;
        RECT 377.400 47.400 378.200 47.600 ;
        RECT 380.200 47.400 381.000 47.600 ;
        RECT 374.000 46.200 374.800 47.000 ;
        RECT 377.400 46.800 381.000 47.400 ;
        RECT 379.600 46.200 380.200 46.800 ;
        RECT 383.600 46.200 384.400 47.000 ;
        RECT 374.000 45.600 376.000 46.200 ;
        RECT 375.200 42.200 376.000 45.600 ;
        RECT 379.600 42.200 380.400 46.200 ;
        RECT 383.800 42.200 385.000 46.200 ;
        RECT 388.400 42.200 389.200 50.800 ;
        RECT 391.600 50.300 392.400 59.800 ;
        RECT 393.800 58.400 394.600 59.800 ;
        RECT 393.800 57.600 395.600 58.400 ;
        RECT 393.800 56.400 394.600 57.600 ;
        RECT 393.800 55.800 395.600 56.400 ;
        RECT 393.200 50.300 394.000 50.400 ;
        RECT 391.600 49.700 394.000 50.300 ;
        RECT 391.600 42.200 392.400 49.700 ;
        RECT 393.200 48.800 394.000 49.700 ;
        RECT 394.800 42.200 395.600 55.800 ;
        RECT 396.400 53.600 397.200 55.200 ;
        RECT 398.000 55.000 398.800 59.800 ;
        RECT 402.400 58.400 403.200 59.800 ;
        RECT 401.200 57.800 403.200 58.400 ;
        RECT 406.800 57.800 407.600 59.800 ;
        RECT 411.000 58.400 412.200 59.800 ;
        RECT 410.800 57.800 412.200 58.400 ;
        RECT 401.200 57.000 402.000 57.800 ;
        RECT 406.800 57.200 407.400 57.800 ;
        RECT 402.800 56.400 403.600 57.200 ;
        RECT 404.600 56.600 407.400 57.200 ;
        RECT 410.800 57.000 411.600 57.800 ;
        RECT 404.600 56.400 405.400 56.600 ;
        RECT 398.800 54.200 400.400 54.400 ;
        RECT 403.000 54.200 403.600 56.400 ;
        RECT 412.600 55.400 413.400 55.600 ;
        RECT 415.600 55.400 416.400 59.800 ;
        RECT 412.600 54.800 416.400 55.400 ;
        RECT 408.600 54.200 410.000 54.400 ;
        RECT 398.800 53.600 410.000 54.200 ;
        RECT 401.800 53.400 402.600 53.600 ;
        RECT 400.200 52.400 401.000 52.600 ;
        RECT 402.800 52.400 403.600 52.600 ;
        RECT 400.200 51.800 405.200 52.400 ;
        RECT 404.400 51.600 405.200 51.800 ;
        RECT 398.000 51.000 403.600 51.200 ;
        RECT 398.000 50.800 403.800 51.000 ;
        RECT 398.000 50.600 407.800 50.800 ;
        RECT 398.000 42.200 398.800 50.600 ;
        RECT 403.000 50.200 407.800 50.600 ;
        RECT 401.200 49.000 406.600 49.600 ;
        RECT 401.200 48.800 402.000 49.000 ;
        RECT 405.800 48.800 406.600 49.000 ;
        RECT 407.200 49.000 407.800 50.200 ;
        RECT 409.200 50.400 409.800 53.600 ;
        RECT 410.800 52.800 411.600 53.000 ;
        RECT 410.800 52.200 414.600 52.800 ;
        RECT 413.800 52.000 414.600 52.200 ;
        RECT 412.200 51.400 413.000 51.600 ;
        RECT 415.600 51.400 416.400 54.800 ;
        RECT 417.200 55.200 418.000 59.800 ;
        RECT 420.400 56.400 421.200 59.800 ;
        RECT 420.400 55.800 421.400 56.400 ;
        RECT 417.200 54.600 419.800 55.200 ;
        RECT 417.400 52.400 418.200 53.200 ;
        RECT 417.200 51.600 418.200 52.400 ;
        RECT 419.200 53.000 419.800 54.600 ;
        RECT 420.800 54.400 421.400 55.800 ;
        RECT 423.600 55.800 424.400 59.800 ;
        RECT 428.000 56.200 429.600 59.800 ;
        RECT 423.600 55.200 425.800 55.800 ;
        RECT 426.800 55.400 428.400 55.600 ;
        RECT 425.000 55.000 425.800 55.200 ;
        RECT 426.400 54.800 428.400 55.400 ;
        RECT 426.400 54.400 427.000 54.800 ;
        RECT 420.400 54.300 421.400 54.400 ;
        RECT 422.000 54.300 422.800 54.400 ;
        RECT 423.600 54.300 427.000 54.400 ;
        RECT 420.400 53.800 427.000 54.300 ;
        RECT 420.400 53.700 425.200 53.800 ;
        RECT 420.400 53.600 421.400 53.700 ;
        RECT 422.000 53.600 422.800 53.700 ;
        RECT 423.600 53.600 425.200 53.700 ;
        RECT 419.200 52.200 420.200 53.000 ;
        RECT 412.200 50.800 416.400 51.400 ;
        RECT 409.200 49.800 411.600 50.400 ;
        RECT 408.600 49.000 409.400 49.200 ;
        RECT 407.200 48.400 409.400 49.000 ;
        RECT 411.000 48.800 411.600 49.800 ;
        RECT 411.000 48.000 412.400 48.800 ;
        RECT 404.600 47.400 405.400 47.600 ;
        RECT 407.400 47.400 408.200 47.600 ;
        RECT 401.200 46.200 402.000 47.000 ;
        RECT 404.600 46.800 408.200 47.400 ;
        RECT 406.800 46.200 407.400 46.800 ;
        RECT 410.800 46.200 411.600 47.000 ;
        RECT 401.200 45.600 403.200 46.200 ;
        RECT 402.400 42.200 403.200 45.600 ;
        RECT 406.800 42.200 407.600 46.200 ;
        RECT 411.000 42.200 412.200 46.200 ;
        RECT 415.600 42.200 416.400 50.800 ;
        RECT 419.200 50.200 419.800 52.200 ;
        RECT 420.800 50.200 421.400 53.600 ;
        RECT 427.600 53.400 428.400 54.200 ;
        RECT 427.600 52.800 428.200 53.400 ;
        RECT 425.600 52.200 428.200 52.800 ;
        RECT 429.000 52.800 429.600 56.200 ;
        RECT 433.200 55.800 434.000 59.800 ;
        RECT 434.800 56.000 435.600 59.800 ;
        RECT 438.000 56.000 438.800 59.800 ;
        RECT 434.800 55.800 438.800 56.000 ;
        RECT 439.600 55.800 440.400 59.800 ;
        RECT 430.200 54.800 431.000 55.600 ;
        RECT 431.600 55.200 434.000 55.800 ;
        RECT 435.000 55.400 438.600 55.800 ;
        RECT 431.600 55.000 432.400 55.200 ;
        RECT 430.400 54.400 431.000 54.800 ;
        RECT 435.600 54.400 436.400 54.800 ;
        RECT 439.600 54.400 440.200 55.800 ;
        RECT 441.200 55.600 442.000 57.200 ;
        RECT 430.400 53.600 431.200 54.400 ;
        RECT 432.400 53.600 434.000 54.400 ;
        RECT 434.800 53.800 436.400 54.400 ;
        RECT 434.800 53.600 435.600 53.800 ;
        RECT 437.800 53.600 440.400 54.400 ;
        RECT 429.000 52.400 430.000 52.800 ;
        RECT 429.000 52.300 430.800 52.400 ;
        RECT 436.400 52.300 437.200 53.200 ;
        RECT 429.000 52.200 437.200 52.300 ;
        RECT 425.600 52.000 426.400 52.200 ;
        RECT 429.400 51.700 437.200 52.200 ;
        RECT 429.400 51.600 430.800 51.700 ;
        RECT 436.400 51.600 437.200 51.700 ;
        RECT 427.800 51.400 428.600 51.600 ;
        RECT 425.200 50.800 428.600 51.400 ;
        RECT 425.200 50.200 425.800 50.800 ;
        RECT 429.400 50.200 430.000 51.600 ;
        RECT 437.800 50.200 438.400 53.600 ;
        RECT 439.600 50.300 440.400 50.400 ;
        RECT 442.800 50.300 443.600 59.800 ;
        RECT 451.800 56.400 452.600 59.800 ;
        RECT 450.800 55.800 452.600 56.400 ;
        RECT 454.000 55.800 454.800 59.800 ;
        RECT 455.600 56.000 456.400 59.800 ;
        RECT 458.800 56.000 459.600 59.800 ;
        RECT 463.000 56.400 463.800 59.800 ;
        RECT 465.800 56.800 466.600 59.800 ;
        RECT 455.600 55.800 459.600 56.000 ;
        RECT 462.000 55.800 463.800 56.400 ;
        RECT 465.200 55.800 466.600 56.800 ;
        RECT 470.000 55.800 470.800 59.800 ;
        RECT 474.800 55.800 475.600 59.800 ;
        RECT 479.600 57.800 480.400 59.800 ;
        RECT 484.400 57.800 485.200 59.800 ;
        RECT 476.200 56.400 477.000 57.200 ;
        RECT 449.200 53.600 450.000 55.200 ;
        RECT 439.600 50.200 443.600 50.300 ;
        RECT 417.200 49.600 419.800 50.200 ;
        RECT 417.200 42.200 418.000 49.600 ;
        RECT 420.400 49.200 421.400 50.200 ;
        RECT 423.600 49.600 425.800 50.200 ;
        RECT 420.400 42.200 421.200 49.200 ;
        RECT 423.600 42.200 424.400 49.600 ;
        RECT 425.000 49.400 425.800 49.600 ;
        RECT 428.000 49.600 430.000 50.200 ;
        RECT 431.600 49.600 434.000 50.200 ;
        RECT 428.000 42.200 429.600 49.600 ;
        RECT 431.600 49.400 432.400 49.600 ;
        RECT 433.200 42.200 434.000 49.600 ;
        RECT 437.400 49.600 438.400 50.200 ;
        RECT 439.000 49.700 443.600 50.200 ;
        RECT 439.000 49.600 440.400 49.700 ;
        RECT 437.400 44.400 438.200 49.600 ;
        RECT 439.000 48.400 439.600 49.600 ;
        RECT 438.800 47.600 439.600 48.400 ;
        RECT 436.400 43.600 438.200 44.400 ;
        RECT 437.400 42.200 438.200 43.600 ;
        RECT 442.800 42.200 443.600 49.700 ;
        RECT 450.800 52.300 451.600 55.800 ;
        RECT 454.200 54.400 454.800 55.800 ;
        RECT 455.800 55.400 459.400 55.800 ;
        RECT 458.000 54.400 458.800 54.800 ;
        RECT 454.000 53.600 456.600 54.400 ;
        RECT 458.000 53.800 459.600 54.400 ;
        RECT 458.800 53.600 459.600 53.800 ;
        RECT 460.400 53.600 461.200 55.200 ;
        RECT 462.000 54.300 462.800 55.800 ;
        RECT 463.600 54.300 464.400 54.400 ;
        RECT 462.000 53.700 464.400 54.300 ;
        RECT 450.800 51.700 454.700 52.300 ;
        RECT 450.800 42.200 451.600 51.700 ;
        RECT 454.100 50.400 454.700 51.700 ;
        RECT 452.400 48.800 453.200 50.400 ;
        RECT 454.000 50.200 454.800 50.400 ;
        RECT 456.000 50.200 456.600 53.600 ;
        RECT 457.200 51.600 458.000 53.200 ;
        RECT 454.000 49.600 455.400 50.200 ;
        RECT 456.000 49.600 457.000 50.200 ;
        RECT 454.800 48.400 455.400 49.600 ;
        RECT 454.800 47.600 455.600 48.400 ;
        RECT 456.200 42.200 457.000 49.600 ;
        RECT 462.000 42.200 462.800 53.700 ;
        RECT 463.600 53.600 464.400 53.700 ;
        RECT 465.200 52.400 465.800 55.800 ;
        RECT 470.000 55.600 470.600 55.800 ;
        RECT 468.800 55.200 470.600 55.600 ;
        RECT 466.400 55.000 470.600 55.200 ;
        RECT 466.400 54.600 469.400 55.000 ;
        RECT 466.400 54.400 467.200 54.600 ;
        RECT 465.200 51.600 466.000 52.400 ;
        RECT 465.200 50.400 465.800 51.600 ;
        RECT 466.600 51.000 467.200 54.400 ;
        RECT 470.000 54.300 470.800 54.400 ;
        RECT 473.200 54.300 474.000 54.400 ;
        RECT 468.000 53.800 468.800 54.000 ;
        RECT 468.000 53.200 469.000 53.800 ;
        RECT 468.400 52.400 469.000 53.200 ;
        RECT 470.000 53.700 474.000 54.300 ;
        RECT 470.000 52.800 470.800 53.700 ;
        RECT 473.200 52.800 474.000 53.700 ;
        RECT 468.400 51.600 469.200 52.400 ;
        RECT 471.600 52.200 472.400 52.400 ;
        RECT 474.800 52.200 475.400 55.800 ;
        RECT 476.400 55.600 477.200 56.400 ;
        RECT 478.000 55.600 478.800 57.200 ;
        RECT 479.800 56.300 480.400 57.800 ;
        RECT 482.800 56.300 483.600 57.200 ;
        RECT 484.600 56.300 485.200 57.800 ;
        RECT 486.000 56.300 486.800 56.400 ;
        RECT 479.700 55.700 483.600 56.300 ;
        RECT 484.500 55.700 486.800 56.300 ;
        RECT 487.600 56.000 488.400 59.800 ;
        RECT 490.800 56.000 491.600 59.800 ;
        RECT 487.600 55.800 491.600 56.000 ;
        RECT 492.400 55.800 493.200 59.800 ;
        RECT 479.800 54.400 480.400 55.700 ;
        RECT 482.800 55.600 483.600 55.700 ;
        RECT 484.600 54.400 485.200 55.700 ;
        RECT 486.000 55.600 486.800 55.700 ;
        RECT 487.800 55.400 491.400 55.800 ;
        RECT 488.400 54.400 489.200 54.800 ;
        RECT 492.400 54.400 493.000 55.800 ;
        RECT 494.000 55.600 494.800 57.200 ;
        RECT 479.600 53.600 480.400 54.400 ;
        RECT 484.400 53.600 485.200 54.400 ;
        RECT 487.600 53.800 489.200 54.400 ;
        RECT 487.600 53.600 488.400 53.800 ;
        RECT 490.600 53.600 493.200 54.400 ;
        RECT 495.600 54.300 496.400 59.800 ;
        RECT 497.400 56.400 498.200 57.200 ;
        RECT 497.200 55.600 498.000 56.400 ;
        RECT 498.800 55.800 499.600 59.800 ;
        RECT 503.800 56.400 504.600 57.200 ;
        RECT 497.200 54.300 498.000 54.400 ;
        RECT 495.600 53.700 498.000 54.300 ;
        RECT 476.400 52.200 477.200 52.400 ;
        RECT 471.600 51.600 473.200 52.200 ;
        RECT 474.800 51.600 477.200 52.200 ;
        RECT 472.400 51.200 473.200 51.600 ;
        RECT 466.600 50.400 469.000 51.000 ;
        RECT 463.600 48.800 464.400 50.400 ;
        RECT 465.200 42.200 466.000 50.400 ;
        RECT 468.400 46.200 469.000 50.400 ;
        RECT 476.400 50.200 477.000 51.600 ;
        RECT 479.800 50.200 480.400 53.600 ;
        RECT 481.200 50.800 482.000 52.400 ;
        RECT 484.600 50.200 485.200 53.600 ;
        RECT 486.000 50.800 486.800 52.400 ;
        RECT 489.200 51.600 490.000 53.200 ;
        RECT 490.600 50.200 491.200 53.600 ;
        RECT 492.400 50.200 493.200 50.400 ;
        RECT 471.600 49.600 475.600 50.200 ;
        RECT 468.400 42.200 469.200 46.200 ;
        RECT 471.600 42.200 472.400 49.600 ;
        RECT 474.800 42.200 475.600 49.600 ;
        RECT 476.400 42.200 477.200 50.200 ;
        RECT 479.600 49.400 481.400 50.200 ;
        RECT 484.400 49.400 486.200 50.200 ;
        RECT 480.600 42.200 481.400 49.400 ;
        RECT 485.400 42.200 486.200 49.400 ;
        RECT 490.200 49.600 491.200 50.200 ;
        RECT 491.800 49.600 493.200 50.200 ;
        RECT 490.200 42.200 491.000 49.600 ;
        RECT 491.800 48.400 492.400 49.600 ;
        RECT 491.600 47.600 492.400 48.400 ;
        RECT 495.600 42.200 496.400 53.700 ;
        RECT 497.200 53.600 498.000 53.700 ;
        RECT 497.200 52.200 498.000 52.400 ;
        RECT 499.000 52.200 499.600 55.800 ;
        RECT 503.600 55.600 504.400 56.400 ;
        RECT 505.200 55.800 506.000 59.800 ;
        RECT 500.400 52.800 501.200 54.400 ;
        RECT 502.000 52.200 502.800 52.400 ;
        RECT 497.200 51.600 499.600 52.200 ;
        RECT 501.200 51.600 502.800 52.200 ;
        RECT 503.600 52.200 504.400 52.400 ;
        RECT 505.400 52.200 506.000 55.800 ;
        RECT 506.800 54.300 507.600 54.400 ;
        RECT 510.000 54.300 510.800 59.800 ;
        RECT 511.600 55.600 512.400 57.200 ;
        RECT 513.200 55.800 514.000 59.800 ;
        RECT 517.600 58.400 519.200 59.800 ;
        RECT 517.600 57.600 520.400 58.400 ;
        RECT 517.600 56.200 519.200 57.600 ;
        RECT 506.800 53.700 510.800 54.300 ;
        RECT 511.700 54.300 512.300 55.600 ;
        RECT 513.200 55.200 515.600 55.800 ;
        RECT 514.800 55.000 515.600 55.200 ;
        RECT 516.200 54.800 517.000 55.600 ;
        RECT 516.200 54.400 516.800 54.800 ;
        RECT 513.200 54.300 514.800 54.400 ;
        RECT 511.700 53.700 514.800 54.300 ;
        RECT 506.800 52.800 507.600 53.700 ;
        RECT 508.400 52.200 509.200 52.400 ;
        RECT 503.600 51.600 506.000 52.200 ;
        RECT 507.600 51.600 509.200 52.200 ;
        RECT 497.400 50.200 498.000 51.600 ;
        RECT 501.200 51.200 502.000 51.600 ;
        RECT 503.800 50.200 504.400 51.600 ;
        RECT 507.600 51.200 508.400 51.600 ;
        RECT 497.200 42.200 498.000 50.200 ;
        RECT 498.800 49.600 502.800 50.200 ;
        RECT 498.800 42.200 499.600 49.600 ;
        RECT 502.000 42.200 502.800 49.600 ;
        RECT 503.600 42.200 504.400 50.200 ;
        RECT 505.200 49.600 509.200 50.200 ;
        RECT 505.200 42.200 506.000 49.600 ;
        RECT 508.400 42.200 509.200 49.600 ;
        RECT 510.000 42.200 510.800 53.700 ;
        RECT 513.200 53.600 514.800 53.700 ;
        RECT 516.000 53.600 516.800 54.400 ;
        RECT 517.600 52.800 518.200 56.200 ;
        RECT 522.800 55.800 523.600 59.800 ;
        RECT 518.800 55.400 520.400 55.600 ;
        RECT 518.800 54.800 520.800 55.400 ;
        RECT 521.400 55.200 523.600 55.800 ;
        RECT 521.400 55.000 522.200 55.200 ;
        RECT 524.400 55.000 525.200 59.800 ;
        RECT 528.800 58.400 529.600 59.800 ;
        RECT 527.600 57.800 529.600 58.400 ;
        RECT 533.200 57.800 534.000 59.800 ;
        RECT 537.400 58.400 538.600 59.800 ;
        RECT 537.200 57.800 538.600 58.400 ;
        RECT 527.600 57.000 528.400 57.800 ;
        RECT 533.200 57.200 533.800 57.800 ;
        RECT 529.200 56.400 530.000 57.200 ;
        RECT 531.000 56.600 533.800 57.200 ;
        RECT 537.200 57.000 538.000 57.800 ;
        RECT 531.000 56.400 531.800 56.600 ;
        RECT 520.200 54.400 520.800 54.800 ;
        RECT 518.800 53.400 519.600 54.200 ;
        RECT 520.200 53.800 523.600 54.400 ;
        RECT 522.000 53.600 523.600 53.800 ;
        RECT 525.200 54.200 526.800 54.400 ;
        RECT 529.400 54.200 530.000 56.400 ;
        RECT 539.000 55.400 539.800 55.600 ;
        RECT 542.000 55.400 542.800 59.800 ;
        RECT 539.000 54.800 542.800 55.400 ;
        RECT 535.000 54.200 535.800 54.400 ;
        RECT 525.200 53.600 536.200 54.200 ;
        RECT 528.200 53.400 529.000 53.600 ;
        RECT 517.200 52.400 518.200 52.800 ;
        RECT 516.400 52.200 518.200 52.400 ;
        RECT 519.000 52.800 519.600 53.400 ;
        RECT 519.000 52.200 521.600 52.800 ;
        RECT 516.400 51.600 517.800 52.200 ;
        RECT 520.800 52.000 521.600 52.200 ;
        RECT 526.600 52.400 527.400 52.600 ;
        RECT 535.600 52.400 536.200 53.600 ;
        RECT 537.200 52.800 538.000 53.000 ;
        RECT 526.600 52.300 531.600 52.400 ;
        RECT 532.400 52.300 533.200 52.400 ;
        RECT 526.600 51.800 533.200 52.300 ;
        RECT 530.800 51.700 533.200 51.800 ;
        RECT 530.800 51.600 531.600 51.700 ;
        RECT 532.400 51.600 533.200 51.700 ;
        RECT 535.600 51.600 536.400 52.400 ;
        RECT 537.200 52.200 541.000 52.800 ;
        RECT 540.200 52.000 541.000 52.200 ;
        RECT 517.200 50.200 517.800 51.600 ;
        RECT 518.600 51.400 519.400 51.600 ;
        RECT 518.600 50.800 522.000 51.400 ;
        RECT 521.400 50.200 522.000 50.800 ;
        RECT 524.400 51.000 530.000 51.200 ;
        RECT 524.400 50.800 530.200 51.000 ;
        RECT 524.400 50.600 534.200 50.800 ;
        RECT 513.200 49.600 515.600 50.200 ;
        RECT 517.200 49.600 519.200 50.200 ;
        RECT 513.200 42.200 514.000 49.600 ;
        RECT 514.800 49.400 515.600 49.600 ;
        RECT 517.600 42.200 519.200 49.600 ;
        RECT 521.400 49.600 523.600 50.200 ;
        RECT 521.400 49.400 522.200 49.600 ;
        RECT 522.800 42.200 523.600 49.600 ;
        RECT 524.400 42.200 525.200 50.600 ;
        RECT 529.400 50.200 534.200 50.600 ;
        RECT 527.600 49.000 533.000 49.600 ;
        RECT 527.600 48.800 528.400 49.000 ;
        RECT 532.200 48.800 533.000 49.000 ;
        RECT 533.600 49.000 534.200 50.200 ;
        RECT 535.600 50.400 536.200 51.600 ;
        RECT 538.600 51.400 539.400 51.600 ;
        RECT 542.000 51.400 542.800 54.800 ;
        RECT 538.600 50.800 542.800 51.400 ;
        RECT 535.600 49.800 538.000 50.400 ;
        RECT 535.000 49.000 535.800 49.200 ;
        RECT 533.600 48.400 535.800 49.000 ;
        RECT 537.400 48.800 538.000 49.800 ;
        RECT 537.400 48.000 538.800 48.800 ;
        RECT 531.000 47.400 531.800 47.600 ;
        RECT 533.800 47.400 534.600 47.600 ;
        RECT 527.600 46.200 528.400 47.000 ;
        RECT 531.000 46.800 534.600 47.400 ;
        RECT 533.200 46.200 533.800 46.800 ;
        RECT 537.200 46.200 538.000 47.000 ;
        RECT 527.600 45.600 529.600 46.200 ;
        RECT 528.800 42.200 529.600 45.600 ;
        RECT 533.200 42.200 534.000 46.200 ;
        RECT 537.400 42.200 538.600 46.200 ;
        RECT 542.000 42.200 542.800 50.800 ;
        RECT 543.600 55.400 544.400 59.800 ;
        RECT 547.800 58.400 549.000 59.800 ;
        RECT 547.800 57.800 549.200 58.400 ;
        RECT 552.400 57.800 553.200 59.800 ;
        RECT 556.800 58.400 557.600 59.800 ;
        RECT 556.800 57.800 558.800 58.400 ;
        RECT 548.400 57.000 549.200 57.800 ;
        RECT 552.600 57.200 553.200 57.800 ;
        RECT 552.600 56.600 555.400 57.200 ;
        RECT 554.600 56.400 555.400 56.600 ;
        RECT 556.400 56.400 557.200 57.200 ;
        RECT 558.000 57.000 558.800 57.800 ;
        RECT 546.600 55.400 547.400 55.600 ;
        RECT 543.600 54.800 547.400 55.400 ;
        RECT 543.600 51.400 544.400 54.800 ;
        RECT 550.000 54.200 551.400 54.400 ;
        RECT 556.400 54.200 557.000 56.400 ;
        RECT 561.200 55.000 562.000 59.800 ;
        RECT 562.800 55.400 563.600 59.800 ;
        RECT 567.000 58.400 568.200 59.800 ;
        RECT 567.000 57.800 568.400 58.400 ;
        RECT 571.600 57.800 572.400 59.800 ;
        RECT 576.000 58.400 576.800 59.800 ;
        RECT 576.000 57.800 578.000 58.400 ;
        RECT 567.600 57.000 568.400 57.800 ;
        RECT 571.800 57.200 572.400 57.800 ;
        RECT 571.800 56.600 574.600 57.200 ;
        RECT 573.800 56.400 574.600 56.600 ;
        RECT 575.600 56.400 576.400 57.200 ;
        RECT 577.200 57.000 578.000 57.800 ;
        RECT 565.800 55.400 566.600 55.600 ;
        RECT 562.800 54.800 566.600 55.400 ;
        RECT 559.600 54.200 561.200 54.400 ;
        RECT 550.000 53.600 561.200 54.200 ;
        RECT 548.400 52.800 549.200 53.000 ;
        RECT 545.400 52.200 549.200 52.800 ;
        RECT 545.400 52.000 546.200 52.200 ;
        RECT 547.000 51.400 547.800 51.600 ;
        RECT 543.600 50.800 547.800 51.400 ;
        RECT 543.600 42.200 544.400 50.800 ;
        RECT 550.200 50.400 550.800 53.600 ;
        RECT 557.400 53.400 558.200 53.600 ;
        RECT 556.400 52.400 557.200 52.600 ;
        RECT 559.000 52.400 559.800 52.600 ;
        RECT 554.800 51.800 559.800 52.400 ;
        RECT 554.800 51.600 555.600 51.800 ;
        RECT 562.800 51.400 563.600 54.800 ;
        RECT 569.800 54.200 570.600 54.400 ;
        RECT 572.400 54.200 573.200 54.400 ;
        RECT 575.600 54.200 576.200 56.400 ;
        RECT 580.400 55.000 581.200 59.800 ;
        RECT 578.800 54.200 580.400 54.400 ;
        RECT 569.400 53.600 580.400 54.200 ;
        RECT 567.600 52.800 568.400 53.000 ;
        RECT 564.600 52.200 568.400 52.800 ;
        RECT 564.600 52.000 565.400 52.200 ;
        RECT 566.200 51.400 567.000 51.600 ;
        RECT 556.400 51.000 562.000 51.200 ;
        RECT 556.200 50.800 562.000 51.000 ;
        RECT 548.400 49.800 550.800 50.400 ;
        RECT 552.200 50.600 562.000 50.800 ;
        RECT 552.200 50.200 557.000 50.600 ;
        RECT 548.400 48.800 549.000 49.800 ;
        RECT 547.600 48.000 549.000 48.800 ;
        RECT 550.600 49.000 551.400 49.200 ;
        RECT 552.200 49.000 552.800 50.200 ;
        RECT 550.600 48.400 552.800 49.000 ;
        RECT 553.400 49.000 558.800 49.600 ;
        RECT 553.400 48.800 554.200 49.000 ;
        RECT 558.000 48.800 558.800 49.000 ;
        RECT 551.800 47.400 552.600 47.600 ;
        RECT 554.600 47.400 555.400 47.600 ;
        RECT 548.400 46.200 549.200 47.000 ;
        RECT 551.800 46.800 555.400 47.400 ;
        RECT 552.600 46.200 553.200 46.800 ;
        RECT 558.000 46.200 558.800 47.000 ;
        RECT 547.800 42.200 549.000 46.200 ;
        RECT 552.400 42.200 553.200 46.200 ;
        RECT 556.800 45.600 558.800 46.200 ;
        RECT 556.800 42.200 557.600 45.600 ;
        RECT 561.200 42.200 562.000 50.600 ;
        RECT 562.800 50.800 567.000 51.400 ;
        RECT 562.800 42.200 563.600 50.800 ;
        RECT 569.400 50.400 570.000 53.600 ;
        RECT 576.600 53.400 577.400 53.600 ;
        RECT 575.600 52.400 576.400 52.600 ;
        RECT 578.200 52.400 579.000 52.600 ;
        RECT 574.000 51.800 579.000 52.400 ;
        RECT 574.000 51.600 574.800 51.800 ;
        RECT 575.600 51.000 581.200 51.200 ;
        RECT 575.400 50.800 581.200 51.000 ;
        RECT 567.600 49.800 570.000 50.400 ;
        RECT 571.400 50.600 581.200 50.800 ;
        RECT 571.400 50.200 576.200 50.600 ;
        RECT 567.600 48.800 568.200 49.800 ;
        RECT 566.800 48.000 568.200 48.800 ;
        RECT 569.800 49.000 570.600 49.200 ;
        RECT 571.400 49.000 572.000 50.200 ;
        RECT 569.800 48.400 572.000 49.000 ;
        RECT 572.600 49.000 578.000 49.600 ;
        RECT 572.600 48.800 573.400 49.000 ;
        RECT 577.200 48.800 578.000 49.000 ;
        RECT 571.000 47.400 571.800 47.600 ;
        RECT 573.800 47.400 574.600 47.600 ;
        RECT 567.600 46.200 568.400 47.000 ;
        RECT 571.000 46.800 574.600 47.400 ;
        RECT 571.800 46.200 572.400 46.800 ;
        RECT 577.200 46.200 578.000 47.000 ;
        RECT 567.000 42.200 568.200 46.200 ;
        RECT 571.600 42.200 572.400 46.200 ;
        RECT 576.000 45.600 578.000 46.200 ;
        RECT 576.000 42.200 576.800 45.600 ;
        RECT 580.400 42.200 581.200 50.600 ;
        RECT 2.800 28.300 3.600 39.800 ;
        RECT 4.400 28.300 5.200 28.400 ;
        RECT 2.800 27.700 5.200 28.300 ;
        RECT 1.200 24.800 2.000 26.400 ;
        RECT 2.800 22.200 3.600 27.700 ;
        RECT 4.400 26.800 5.200 27.700 ;
        RECT 6.000 26.200 6.800 39.800 ;
        RECT 7.600 31.600 8.400 33.200 ;
        RECT 9.200 26.800 10.000 28.400 ;
        RECT 10.800 26.200 11.600 39.800 ;
        RECT 12.400 31.600 13.200 33.200 ;
        RECT 14.000 31.800 14.800 39.800 ;
        RECT 15.600 32.400 16.400 39.800 ;
        RECT 18.800 32.400 19.600 39.800 ;
        RECT 21.200 33.600 22.000 34.400 ;
        RECT 21.200 32.400 21.800 33.600 ;
        RECT 22.600 32.400 23.400 39.800 ;
        RECT 15.600 31.800 19.600 32.400 ;
        RECT 20.400 31.800 21.800 32.400 ;
        RECT 22.400 31.800 23.400 32.400 ;
        RECT 26.800 31.800 27.600 39.800 ;
        RECT 30.000 32.400 30.800 39.800 ;
        RECT 28.600 31.800 30.800 32.400 ;
        RECT 14.200 30.400 14.800 31.800 ;
        RECT 20.400 31.600 21.200 31.800 ;
        RECT 18.000 30.400 18.800 30.800 ;
        RECT 14.000 29.800 16.400 30.400 ;
        RECT 18.000 29.800 19.600 30.400 ;
        RECT 14.000 29.600 14.800 29.800 ;
        RECT 6.000 25.600 7.800 26.200 ;
        RECT 10.800 25.600 12.600 26.200 ;
        RECT 14.000 25.600 14.800 26.400 ;
        RECT 15.800 26.200 16.400 29.800 ;
        RECT 18.800 29.600 19.600 29.800 ;
        RECT 17.200 27.600 18.000 29.200 ;
        RECT 22.400 28.400 23.000 31.800 ;
        RECT 23.600 28.800 24.400 30.400 ;
        RECT 26.800 29.600 27.400 31.800 ;
        RECT 28.600 31.200 29.200 31.800 ;
        RECT 28.000 30.400 29.200 31.200 ;
        RECT 20.400 27.600 23.000 28.400 ;
        RECT 25.200 28.300 26.000 28.400 ;
        RECT 26.800 28.300 27.600 29.600 ;
        RECT 25.200 28.200 27.600 28.300 ;
        RECT 24.400 27.700 27.600 28.200 ;
        RECT 24.400 27.600 26.000 27.700 ;
        RECT 20.600 26.200 21.200 27.600 ;
        RECT 24.400 27.200 25.200 27.600 ;
        RECT 22.200 26.200 25.800 26.600 ;
        RECT 7.000 24.400 7.800 25.600 ;
        RECT 6.000 23.600 7.800 24.400 ;
        RECT 7.000 22.200 7.800 23.600 ;
        RECT 11.800 22.200 12.600 25.600 ;
        RECT 14.200 24.800 15.000 25.600 ;
        RECT 15.600 22.200 16.400 26.200 ;
        RECT 20.400 22.200 21.200 26.200 ;
        RECT 22.000 26.000 26.000 26.200 ;
        RECT 22.000 22.200 22.800 26.000 ;
        RECT 25.200 22.200 26.000 26.000 ;
        RECT 26.800 22.200 27.600 27.700 ;
        RECT 28.600 27.400 29.200 30.400 ;
        RECT 30.000 28.800 30.800 30.400 ;
        RECT 28.600 26.800 30.800 27.400 ;
        RECT 31.600 26.800 32.400 28.400 ;
        RECT 30.000 22.200 30.800 26.800 ;
        RECT 33.200 26.200 34.000 39.800 ;
        RECT 37.200 33.600 38.000 34.400 ;
        RECT 34.800 31.600 35.600 33.200 ;
        RECT 37.200 32.400 37.800 33.600 ;
        RECT 38.600 32.400 39.400 39.800 ;
        RECT 36.400 31.800 37.800 32.400 ;
        RECT 38.400 31.800 39.400 32.400 ;
        RECT 42.800 32.400 43.600 39.800 ;
        RECT 46.000 32.400 46.800 39.800 ;
        RECT 42.800 31.800 46.800 32.400 ;
        RECT 47.600 31.800 48.400 39.800 ;
        RECT 36.400 31.600 37.200 31.800 ;
        RECT 34.900 30.300 35.500 31.600 ;
        RECT 38.400 30.300 39.000 31.800 ;
        RECT 43.600 30.400 44.400 30.800 ;
        RECT 47.600 30.400 48.200 31.800 ;
        RECT 34.900 29.700 39.000 30.300 ;
        RECT 38.400 28.400 39.000 29.700 ;
        RECT 39.600 28.800 40.400 30.400 ;
        RECT 42.800 29.800 44.400 30.400 ;
        RECT 46.000 29.800 48.400 30.400 ;
        RECT 42.800 29.600 43.600 29.800 ;
        RECT 36.400 27.600 39.000 28.400 ;
        RECT 41.200 28.200 42.000 28.400 ;
        RECT 40.400 27.600 42.000 28.200 ;
        RECT 44.400 27.600 45.200 29.200 ;
        RECT 36.600 26.200 37.200 27.600 ;
        RECT 40.400 27.200 41.200 27.600 ;
        RECT 38.200 26.200 41.800 26.600 ;
        RECT 46.000 26.400 46.600 29.800 ;
        RECT 47.600 29.600 48.400 29.800 ;
        RECT 33.200 25.600 35.000 26.200 ;
        RECT 34.200 24.400 35.000 25.600 ;
        RECT 34.200 23.600 35.600 24.400 ;
        RECT 34.200 22.200 35.000 23.600 ;
        RECT 36.400 22.200 37.200 26.200 ;
        RECT 38.000 26.000 42.000 26.200 ;
        RECT 38.000 22.200 38.800 26.000 ;
        RECT 41.200 22.200 42.000 26.000 ;
        RECT 46.000 22.200 46.800 26.400 ;
        RECT 47.600 26.300 48.400 26.400 ;
        RECT 49.200 26.300 50.000 26.400 ;
        RECT 47.600 25.700 50.000 26.300 ;
        RECT 47.600 25.600 48.400 25.700 ;
        RECT 47.400 24.800 48.200 25.600 ;
        RECT 49.200 24.800 50.000 25.700 ;
        RECT 50.800 22.200 51.600 39.800 ;
        RECT 52.400 32.400 53.200 39.800 ;
        RECT 55.600 32.800 56.400 39.800 ;
        RECT 52.400 31.800 55.000 32.400 ;
        RECT 55.600 31.800 56.600 32.800 ;
        RECT 58.800 32.400 59.600 39.800 ;
        RECT 60.400 32.400 61.200 32.600 ;
        RECT 63.200 32.400 64.800 39.800 ;
        RECT 58.800 31.800 61.200 32.400 ;
        RECT 62.800 31.800 64.800 32.400 ;
        RECT 67.000 32.400 67.800 32.600 ;
        RECT 68.400 32.400 69.200 39.800 ;
        RECT 67.000 31.800 69.200 32.400 ;
        RECT 52.400 29.600 53.400 30.400 ;
        RECT 52.600 28.800 53.400 29.600 ;
        RECT 54.400 29.800 55.000 31.800 ;
        RECT 54.400 29.000 55.400 29.800 ;
        RECT 54.400 27.400 55.000 29.000 ;
        RECT 56.000 28.400 56.600 31.800 ;
        RECT 62.800 30.400 63.400 31.800 ;
        RECT 67.000 31.200 67.600 31.800 ;
        RECT 64.200 30.600 67.600 31.200 ;
        RECT 70.000 31.400 70.800 39.800 ;
        RECT 74.400 36.400 75.200 39.800 ;
        RECT 73.200 35.800 75.200 36.400 ;
        RECT 78.800 35.800 79.600 39.800 ;
        RECT 83.000 35.800 84.200 39.800 ;
        RECT 73.200 35.000 74.000 35.800 ;
        RECT 78.800 35.200 79.400 35.800 ;
        RECT 76.600 34.600 80.200 35.200 ;
        RECT 82.800 35.000 83.600 35.800 ;
        RECT 76.600 34.400 77.400 34.600 ;
        RECT 79.400 34.400 80.200 34.600 ;
        RECT 73.200 33.000 74.000 33.200 ;
        RECT 77.800 33.000 78.600 33.200 ;
        RECT 73.200 32.400 78.600 33.000 ;
        RECT 79.200 33.000 81.400 33.600 ;
        RECT 79.200 31.800 79.800 33.000 ;
        RECT 80.600 32.800 81.400 33.000 ;
        RECT 83.000 33.200 84.400 34.000 ;
        RECT 83.000 32.200 83.600 33.200 ;
        RECT 75.000 31.400 79.800 31.800 ;
        RECT 70.000 31.200 79.800 31.400 ;
        RECT 81.200 31.600 83.600 32.200 ;
        RECT 70.000 31.000 75.800 31.200 ;
        RECT 70.000 30.800 75.600 31.000 ;
        RECT 64.200 30.400 65.000 30.600 ;
        RECT 62.000 29.800 63.400 30.400 ;
        RECT 76.400 30.200 77.200 30.400 ;
        RECT 66.400 29.800 67.200 30.000 ;
        RECT 62.000 29.600 63.800 29.800 ;
        RECT 62.800 29.200 63.800 29.600 ;
        RECT 55.600 27.600 56.600 28.400 ;
        RECT 58.800 27.600 60.400 28.400 ;
        RECT 61.600 27.600 62.400 28.400 ;
        RECT 52.400 26.800 55.000 27.400 ;
        RECT 52.400 22.200 53.200 26.800 ;
        RECT 56.000 26.200 56.600 27.600 ;
        RECT 61.800 27.200 62.400 27.600 ;
        RECT 60.400 26.800 61.200 27.000 ;
        RECT 55.600 25.600 56.600 26.200 ;
        RECT 58.800 26.200 61.200 26.800 ;
        RECT 61.800 26.400 62.600 27.200 ;
        RECT 55.600 22.200 56.400 25.600 ;
        RECT 58.800 22.200 59.600 26.200 ;
        RECT 63.200 25.800 63.800 29.200 ;
        RECT 64.600 29.200 67.200 29.800 ;
        RECT 72.200 29.600 77.200 30.200 ;
        RECT 79.600 30.300 80.400 30.400 ;
        RECT 81.200 30.300 81.800 31.600 ;
        RECT 87.600 31.200 88.400 39.800 ;
        RECT 89.200 32.400 90.000 39.800 ;
        RECT 90.600 32.400 91.400 32.600 ;
        RECT 89.200 31.800 91.400 32.400 ;
        RECT 93.600 32.400 95.200 39.800 ;
        RECT 97.200 32.400 98.000 32.600 ;
        RECT 98.800 32.400 99.600 39.800 ;
        RECT 101.200 33.600 102.000 34.400 ;
        RECT 101.200 32.400 101.800 33.600 ;
        RECT 102.600 32.400 103.400 39.800 ;
        RECT 93.600 31.800 95.600 32.400 ;
        RECT 97.200 31.800 99.600 32.400 ;
        RECT 100.400 31.800 101.800 32.400 ;
        RECT 102.400 31.800 103.400 32.400 ;
        RECT 84.200 30.600 88.400 31.200 ;
        RECT 90.800 31.200 91.400 31.800 ;
        RECT 90.800 30.600 94.200 31.200 ;
        RECT 84.200 30.400 85.000 30.600 ;
        RECT 79.600 29.700 81.900 30.300 ;
        RECT 85.800 29.800 86.600 30.000 ;
        RECT 79.600 29.600 80.400 29.700 ;
        RECT 72.200 29.400 73.000 29.600 ;
        RECT 64.600 28.600 65.200 29.200 ;
        RECT 64.400 27.800 65.200 28.600 ;
        RECT 73.800 28.400 74.600 28.600 ;
        RECT 81.200 28.400 81.800 29.700 ;
        RECT 82.800 29.200 86.600 29.800 ;
        RECT 82.800 29.000 83.600 29.200 ;
        RECT 67.600 28.200 69.200 28.400 ;
        RECT 65.800 27.600 69.200 28.200 ;
        RECT 70.800 27.800 81.800 28.400 ;
        RECT 70.800 27.600 72.400 27.800 ;
        RECT 65.800 27.200 66.400 27.600 ;
        RECT 64.400 26.600 66.400 27.200 ;
        RECT 67.000 26.800 67.800 27.000 ;
        RECT 64.400 26.400 66.000 26.600 ;
        RECT 67.000 26.200 69.200 26.800 ;
        RECT 63.200 24.400 64.800 25.800 ;
        RECT 63.200 23.600 66.000 24.400 ;
        RECT 63.200 22.200 64.800 23.600 ;
        RECT 68.400 22.200 69.200 26.200 ;
        RECT 70.000 22.200 70.800 27.000 ;
        RECT 75.000 25.600 75.600 27.800 ;
        RECT 80.600 27.600 81.400 27.800 ;
        RECT 87.600 27.200 88.400 30.600 ;
        RECT 93.400 30.400 94.200 30.600 ;
        RECT 95.000 30.400 95.600 31.800 ;
        RECT 100.400 31.600 101.200 31.800 ;
        RECT 95.000 30.300 96.400 30.400 ;
        RECT 100.400 30.300 101.200 30.400 ;
        RECT 91.200 29.800 92.000 30.000 ;
        RECT 95.000 29.800 101.200 30.300 ;
        RECT 91.200 29.200 93.800 29.800 ;
        RECT 93.200 28.600 93.800 29.200 ;
        RECT 94.600 29.700 101.200 29.800 ;
        RECT 94.600 29.600 96.400 29.700 ;
        RECT 100.400 29.600 101.200 29.700 ;
        RECT 94.600 29.200 95.600 29.600 ;
        RECT 89.200 28.200 90.800 28.400 ;
        RECT 89.200 27.600 92.600 28.200 ;
        RECT 93.200 27.800 94.000 28.600 ;
        RECT 84.600 26.600 88.400 27.200 ;
        RECT 92.000 27.200 92.600 27.600 ;
        RECT 90.600 26.800 91.400 27.000 ;
        RECT 84.600 26.400 85.400 26.600 ;
        RECT 73.200 24.200 74.000 25.000 ;
        RECT 74.800 24.800 75.600 25.600 ;
        RECT 76.600 25.400 77.400 25.600 ;
        RECT 76.600 24.800 79.400 25.400 ;
        RECT 78.800 24.200 79.400 24.800 ;
        RECT 82.800 24.200 83.600 25.000 ;
        RECT 73.200 23.600 75.200 24.200 ;
        RECT 74.400 22.200 75.200 23.600 ;
        RECT 78.800 22.200 79.600 24.200 ;
        RECT 82.800 23.600 84.200 24.200 ;
        RECT 83.000 22.200 84.200 23.600 ;
        RECT 87.600 22.200 88.400 26.600 ;
        RECT 89.200 26.200 91.400 26.800 ;
        RECT 92.000 26.600 94.000 27.200 ;
        RECT 92.400 26.400 94.000 26.600 ;
        RECT 89.200 22.200 90.000 26.200 ;
        RECT 94.600 25.800 95.200 29.200 ;
        RECT 102.400 28.400 103.000 31.800 ;
        RECT 106.800 31.400 107.600 39.800 ;
        RECT 111.200 36.400 112.000 39.800 ;
        RECT 110.000 35.800 112.000 36.400 ;
        RECT 115.600 35.800 116.400 39.800 ;
        RECT 119.800 35.800 121.000 39.800 ;
        RECT 110.000 35.000 110.800 35.800 ;
        RECT 115.600 35.200 116.200 35.800 ;
        RECT 113.400 34.600 117.000 35.200 ;
        RECT 119.600 35.000 120.400 35.800 ;
        RECT 113.400 34.400 114.200 34.600 ;
        RECT 116.200 34.400 117.000 34.600 ;
        RECT 110.000 33.000 110.800 33.200 ;
        RECT 114.600 33.000 115.400 33.200 ;
        RECT 110.000 32.400 115.400 33.000 ;
        RECT 116.000 33.000 118.200 33.600 ;
        RECT 116.000 31.800 116.600 33.000 ;
        RECT 117.400 32.800 118.200 33.000 ;
        RECT 119.800 33.200 121.200 34.000 ;
        RECT 119.800 32.200 120.400 33.200 ;
        RECT 111.800 31.400 116.600 31.800 ;
        RECT 106.800 31.200 116.600 31.400 ;
        RECT 118.000 31.600 120.400 32.200 ;
        RECT 106.800 31.000 112.600 31.200 ;
        RECT 106.800 30.800 112.400 31.000 ;
        RECT 118.000 30.400 118.600 31.600 ;
        RECT 124.400 31.200 125.200 39.800 ;
        RECT 126.000 32.400 126.800 39.800 ;
        RECT 127.600 32.400 128.400 32.600 ;
        RECT 130.400 32.400 132.000 39.800 ;
        RECT 126.000 31.800 128.400 32.400 ;
        RECT 130.000 31.800 132.000 32.400 ;
        RECT 134.200 32.400 135.000 32.600 ;
        RECT 135.600 32.400 136.400 39.800 ;
        RECT 134.200 31.800 136.400 32.400 ;
        RECT 142.000 32.400 142.800 39.800 ;
        RECT 143.600 32.400 144.400 32.600 ;
        RECT 142.000 31.800 144.400 32.400 ;
        RECT 146.400 31.800 148.000 39.800 ;
        RECT 149.800 32.400 150.600 32.600 ;
        RECT 151.600 32.400 152.400 39.800 ;
        RECT 149.800 31.800 152.400 32.400 ;
        RECT 121.000 30.600 125.200 31.200 ;
        RECT 121.000 30.400 121.800 30.600 ;
        RECT 103.600 28.800 104.400 30.400 ;
        RECT 113.200 30.200 114.000 30.400 ;
        RECT 109.000 29.600 114.000 30.200 ;
        RECT 118.000 29.600 118.800 30.400 ;
        RECT 122.600 29.800 123.400 30.000 ;
        RECT 109.000 29.400 109.800 29.600 ;
        RECT 111.600 29.400 112.400 29.600 ;
        RECT 110.600 28.400 111.400 28.600 ;
        RECT 118.000 28.400 118.600 29.600 ;
        RECT 119.600 29.200 123.400 29.800 ;
        RECT 119.600 29.000 120.400 29.200 ;
        RECT 96.000 27.600 96.800 28.400 ;
        RECT 98.000 27.600 99.600 28.400 ;
        RECT 100.400 27.600 103.000 28.400 ;
        RECT 105.200 28.200 106.000 28.400 ;
        RECT 104.400 27.600 106.000 28.200 ;
        RECT 107.600 27.800 118.600 28.400 ;
        RECT 107.600 27.600 109.200 27.800 ;
        RECT 96.000 27.200 96.600 27.600 ;
        RECT 95.800 26.400 96.600 27.200 ;
        RECT 97.200 26.800 98.000 27.000 ;
        RECT 97.200 26.200 99.600 26.800 ;
        RECT 100.600 26.200 101.200 27.600 ;
        RECT 104.400 27.200 105.200 27.600 ;
        RECT 102.200 26.200 105.800 26.600 ;
        RECT 93.600 22.200 95.200 25.800 ;
        RECT 98.800 22.200 99.600 26.200 ;
        RECT 100.400 22.200 101.200 26.200 ;
        RECT 102.000 26.000 106.000 26.200 ;
        RECT 102.000 22.200 102.800 26.000 ;
        RECT 105.200 22.200 106.000 26.000 ;
        RECT 106.800 22.200 107.600 27.000 ;
        RECT 111.800 25.600 112.400 27.800 ;
        RECT 117.400 27.600 118.200 27.800 ;
        RECT 124.400 27.200 125.200 30.600 ;
        RECT 130.000 30.400 130.600 31.800 ;
        RECT 134.200 31.200 134.800 31.800 ;
        RECT 131.400 30.600 134.800 31.200 ;
        RECT 131.400 30.400 132.200 30.600 ;
        RECT 146.800 30.400 147.400 31.800 ;
        RECT 148.600 30.400 149.400 30.600 ;
        RECT 129.200 29.800 130.600 30.400 ;
        RECT 133.600 29.800 134.400 30.000 ;
        RECT 129.200 29.600 131.000 29.800 ;
        RECT 130.000 29.200 131.000 29.600 ;
        RECT 126.000 27.600 127.600 28.400 ;
        RECT 128.800 27.600 129.600 28.400 ;
        RECT 121.400 26.600 125.200 27.200 ;
        RECT 129.000 27.200 129.600 27.600 ;
        RECT 127.600 26.800 128.400 27.000 ;
        RECT 121.400 26.400 122.200 26.600 ;
        RECT 110.000 24.200 110.800 25.000 ;
        RECT 111.600 24.800 112.400 25.600 ;
        RECT 113.400 25.400 114.200 25.600 ;
        RECT 113.400 24.800 116.200 25.400 ;
        RECT 115.600 24.200 116.200 24.800 ;
        RECT 119.600 24.200 120.400 25.000 ;
        RECT 110.000 23.600 112.000 24.200 ;
        RECT 111.200 22.200 112.000 23.600 ;
        RECT 115.600 22.200 116.400 24.200 ;
        RECT 119.600 23.600 121.000 24.200 ;
        RECT 119.800 22.200 121.000 23.600 ;
        RECT 124.400 22.200 125.200 26.600 ;
        RECT 126.000 26.200 128.400 26.800 ;
        RECT 129.000 26.400 129.800 27.200 ;
        RECT 126.000 22.200 126.800 26.200 ;
        RECT 130.400 25.800 131.000 29.200 ;
        RECT 131.800 29.200 134.400 29.800 ;
        RECT 146.800 29.600 147.600 30.400 ;
        RECT 148.600 29.800 150.200 30.400 ;
        RECT 149.400 29.600 150.200 29.800 ;
        RECT 131.800 28.600 132.400 29.200 ;
        RECT 131.600 27.800 132.400 28.600 ;
        RECT 146.800 28.400 147.400 29.600 ;
        RECT 134.800 28.200 136.400 28.400 ;
        RECT 133.000 27.600 136.400 28.200 ;
        RECT 142.000 27.600 143.600 28.400 ;
        RECT 144.800 27.600 145.600 28.400 ;
        RECT 133.000 27.200 133.600 27.600 ;
        RECT 131.600 26.600 133.600 27.200 ;
        RECT 145.000 27.200 145.600 27.600 ;
        RECT 146.400 27.800 147.400 28.400 ;
        RECT 148.000 28.600 148.800 28.800 ;
        RECT 148.000 28.400 150.800 28.600 ;
        RECT 148.000 28.000 152.400 28.400 ;
        RECT 150.200 27.800 152.400 28.000 ;
        RECT 134.200 26.800 135.000 27.000 ;
        RECT 143.600 26.800 144.400 27.000 ;
        RECT 131.600 26.400 133.200 26.600 ;
        RECT 134.200 26.200 136.400 26.800 ;
        RECT 130.400 24.400 132.000 25.800 ;
        RECT 129.200 23.600 132.000 24.400 ;
        RECT 130.400 22.200 132.000 23.600 ;
        RECT 135.600 22.200 136.400 26.200 ;
        RECT 142.000 26.200 144.400 26.800 ;
        RECT 145.000 26.400 145.800 27.200 ;
        RECT 142.000 22.200 142.800 26.200 ;
        RECT 146.400 25.800 147.000 27.800 ;
        RECT 150.800 27.600 152.400 27.800 ;
        RECT 147.600 26.400 149.200 27.200 ;
        RECT 149.800 26.800 150.600 27.000 ;
        RECT 153.200 26.800 154.000 28.400 ;
        RECT 149.800 26.200 152.400 26.800 ;
        RECT 146.400 24.400 148.000 25.800 ;
        RECT 146.400 23.600 149.200 24.400 ;
        RECT 146.400 22.200 148.000 23.600 ;
        RECT 151.600 22.200 152.400 26.200 ;
        RECT 154.800 26.300 155.600 39.800 ;
        RECT 156.400 31.600 157.200 33.200 ;
        RECT 158.000 26.300 158.800 26.400 ;
        RECT 154.800 25.700 158.800 26.300 ;
        RECT 154.800 25.600 156.600 25.700 ;
        RECT 155.800 24.400 156.600 25.600 ;
        RECT 158.000 24.800 158.800 25.700 ;
        RECT 154.800 23.600 156.600 24.400 ;
        RECT 155.800 22.200 156.600 23.600 ;
        RECT 159.600 22.200 160.400 39.800 ;
        RECT 161.200 26.800 162.000 28.400 ;
        RECT 162.800 26.200 163.600 39.800 ;
        RECT 164.400 31.600 165.200 33.200 ;
        RECT 168.600 32.400 170.600 39.800 ;
        RECT 176.600 32.400 177.400 39.800 ;
        RECT 178.000 33.600 178.800 34.400 ;
        RECT 178.200 32.400 178.800 33.600 ;
        RECT 181.200 33.600 182.000 34.400 ;
        RECT 181.200 32.400 181.800 33.600 ;
        RECT 182.600 32.400 183.400 39.800 ;
        RECT 168.600 31.800 171.600 32.400 ;
        RECT 176.600 31.800 177.600 32.400 ;
        RECT 178.200 31.800 179.600 32.400 ;
        RECT 169.400 31.600 171.600 31.800 ;
        RECT 166.000 27.600 166.800 29.200 ;
        RECT 167.600 28.800 168.400 30.400 ;
        RECT 169.400 28.400 170.000 31.600 ;
        RECT 170.800 30.300 171.600 30.400 ;
        RECT 175.600 30.300 176.400 30.400 ;
        RECT 170.800 29.700 176.400 30.300 ;
        RECT 170.800 28.800 171.600 29.700 ;
        RECT 175.600 28.800 176.400 29.700 ;
        RECT 177.000 30.300 177.600 31.800 ;
        RECT 178.800 31.600 179.600 31.800 ;
        RECT 180.400 31.800 181.800 32.400 ;
        RECT 182.400 31.800 183.400 32.400 ;
        RECT 186.800 32.400 187.600 39.800 ;
        RECT 191.200 38.400 192.800 39.800 ;
        RECT 191.200 37.600 194.000 38.400 ;
        RECT 188.400 32.400 189.200 32.600 ;
        RECT 191.200 32.400 192.800 37.600 ;
        RECT 186.800 31.800 189.200 32.400 ;
        RECT 190.800 31.800 192.800 32.400 ;
        RECT 195.000 32.400 195.800 32.600 ;
        RECT 196.400 32.400 197.200 39.800 ;
        RECT 195.000 31.800 197.200 32.400 ;
        RECT 198.000 32.400 198.800 39.800 ;
        RECT 201.200 32.400 202.000 39.800 ;
        RECT 198.000 31.800 202.000 32.400 ;
        RECT 202.800 31.800 203.600 39.800 ;
        RECT 206.000 35.800 206.800 39.800 ;
        RECT 180.400 31.600 181.200 31.800 ;
        RECT 180.500 30.300 181.100 31.600 ;
        RECT 177.000 29.700 181.100 30.300 ;
        RECT 177.000 28.400 177.600 29.700 ;
        RECT 182.400 28.400 183.000 31.800 ;
        RECT 190.800 30.400 191.400 31.800 ;
        RECT 195.000 31.200 195.600 31.800 ;
        RECT 192.200 30.600 195.600 31.200 ;
        RECT 192.200 30.400 193.000 30.600 ;
        RECT 198.800 30.400 199.600 30.800 ;
        RECT 202.800 30.400 203.400 31.800 ;
        RECT 206.200 31.600 206.800 35.800 ;
        RECT 209.200 31.800 210.000 39.800 ;
        RECT 206.200 31.000 208.600 31.600 ;
        RECT 183.600 28.800 184.400 30.400 ;
        RECT 190.000 29.800 191.400 30.400 ;
        RECT 194.400 29.800 195.200 30.000 ;
        RECT 190.000 29.600 191.800 29.800 ;
        RECT 190.800 29.200 191.800 29.600 ;
        RECT 169.200 28.200 170.000 28.400 ;
        RECT 172.400 28.300 173.200 28.400 ;
        RECT 174.000 28.300 174.800 28.400 ;
        RECT 172.400 28.200 174.800 28.300 ;
        RECT 167.600 27.600 170.000 28.200 ;
        RECT 171.600 27.700 175.600 28.200 ;
        RECT 171.600 27.600 173.200 27.700 ;
        RECT 174.000 27.600 175.600 27.700 ;
        RECT 177.000 27.600 179.600 28.400 ;
        RECT 180.400 27.600 183.000 28.400 ;
        RECT 185.200 28.200 186.000 28.400 ;
        RECT 184.400 27.600 186.000 28.200 ;
        RECT 186.800 27.600 188.400 28.400 ;
        RECT 189.600 27.600 190.400 28.400 ;
        RECT 167.600 26.200 168.200 27.600 ;
        RECT 171.600 27.200 172.400 27.600 ;
        RECT 174.800 27.200 175.600 27.600 ;
        RECT 169.400 26.200 173.000 26.600 ;
        RECT 174.200 26.200 177.800 26.600 ;
        RECT 178.800 26.200 179.400 27.600 ;
        RECT 180.600 26.200 181.200 27.600 ;
        RECT 184.400 27.200 185.200 27.600 ;
        RECT 189.800 27.200 190.400 27.600 ;
        RECT 188.400 26.800 189.200 27.000 ;
        RECT 182.200 26.200 185.800 26.600 ;
        RECT 186.800 26.200 189.200 26.800 ;
        RECT 189.800 26.400 190.600 27.200 ;
        RECT 162.800 25.600 164.600 26.200 ;
        RECT 163.800 22.200 164.600 25.600 ;
        RECT 166.000 22.800 166.800 26.200 ;
        RECT 167.600 23.400 168.400 26.200 ;
        RECT 169.200 26.000 173.200 26.200 ;
        RECT 169.200 22.800 170.000 26.000 ;
        RECT 166.000 22.200 170.000 22.800 ;
        RECT 172.400 22.200 173.200 26.000 ;
        RECT 174.000 26.000 178.000 26.200 ;
        RECT 174.000 22.200 174.800 26.000 ;
        RECT 177.200 22.200 178.000 26.000 ;
        RECT 178.800 22.200 179.600 26.200 ;
        RECT 180.400 22.200 181.200 26.200 ;
        RECT 182.000 26.000 186.000 26.200 ;
        RECT 182.000 22.200 182.800 26.000 ;
        RECT 185.200 22.200 186.000 26.000 ;
        RECT 186.800 22.200 187.600 26.200 ;
        RECT 191.200 25.800 191.800 29.200 ;
        RECT 192.600 29.200 195.200 29.800 ;
        RECT 198.000 29.800 199.600 30.400 ;
        RECT 201.200 29.800 203.600 30.400 ;
        RECT 198.000 29.600 198.800 29.800 ;
        RECT 192.600 28.600 193.200 29.200 ;
        RECT 192.400 27.800 193.200 28.600 ;
        RECT 195.600 28.200 197.200 28.400 ;
        RECT 193.800 27.600 197.200 28.200 ;
        RECT 199.600 27.600 200.400 29.200 ;
        RECT 193.800 27.200 194.400 27.600 ;
        RECT 192.400 26.600 194.400 27.200 ;
        RECT 195.000 26.800 195.800 27.000 ;
        RECT 192.400 26.400 194.000 26.600 ;
        RECT 195.000 26.200 197.200 26.800 ;
        RECT 191.200 22.200 192.800 25.800 ;
        RECT 196.400 22.200 197.200 26.200 ;
        RECT 201.200 26.200 201.800 29.800 ;
        RECT 202.800 29.600 203.600 29.800 ;
        RECT 206.000 29.600 206.800 30.400 ;
        RECT 204.400 27.600 205.200 29.200 ;
        RECT 206.200 28.800 206.800 29.600 ;
        RECT 206.200 28.200 207.200 28.800 ;
        RECT 206.400 28.000 207.200 28.200 ;
        RECT 208.000 27.600 208.600 31.000 ;
        RECT 209.400 30.400 210.000 31.800 ;
        RECT 210.800 31.600 211.600 33.200 ;
        RECT 209.200 29.600 210.000 30.400 ;
        RECT 208.000 27.400 208.800 27.600 ;
        RECT 205.800 27.000 208.800 27.400 ;
        RECT 204.600 26.800 208.800 27.000 ;
        RECT 204.600 26.400 206.400 26.800 ;
        RECT 201.200 22.200 202.000 26.200 ;
        RECT 202.800 25.600 203.600 26.400 ;
        RECT 204.600 26.200 205.200 26.400 ;
        RECT 209.400 26.200 210.000 29.600 ;
        RECT 212.400 30.300 213.200 39.800 ;
        RECT 212.400 29.700 216.300 30.300 ;
        RECT 212.400 26.200 213.200 29.700 ;
        RECT 215.700 28.400 216.300 29.700 ;
        RECT 214.000 26.800 214.800 28.400 ;
        RECT 215.600 26.800 216.400 28.400 ;
        RECT 202.600 24.800 203.400 25.600 ;
        RECT 204.400 22.200 205.200 26.200 ;
        RECT 208.600 25.200 210.000 26.200 ;
        RECT 211.400 25.600 213.200 26.200 ;
        RECT 217.200 26.200 218.000 39.800 ;
        RECT 218.800 31.600 219.600 33.200 ;
        RECT 220.400 32.400 221.200 39.800 ;
        RECT 221.800 32.400 222.600 32.600 ;
        RECT 220.400 31.800 222.600 32.400 ;
        RECT 224.800 32.400 226.400 39.800 ;
        RECT 228.400 32.400 229.200 32.600 ;
        RECT 230.000 32.400 230.800 39.800 ;
        RECT 224.800 31.800 227.600 32.400 ;
        RECT 228.400 31.800 230.800 32.400 ;
        RECT 222.000 31.200 222.600 31.800 ;
        RECT 226.200 31.600 227.600 31.800 ;
        RECT 231.600 31.600 232.400 33.200 ;
        RECT 222.000 30.600 225.400 31.200 ;
        RECT 224.600 30.400 225.400 30.600 ;
        RECT 226.200 30.400 226.800 31.600 ;
        RECT 222.400 29.800 223.200 30.000 ;
        RECT 226.200 29.800 227.600 30.400 ;
        RECT 222.400 29.200 225.000 29.800 ;
        RECT 224.400 28.600 225.000 29.200 ;
        RECT 225.800 29.600 227.600 29.800 ;
        RECT 225.800 29.200 226.800 29.600 ;
        RECT 220.400 28.200 222.000 28.400 ;
        RECT 220.400 27.600 223.800 28.200 ;
        RECT 224.400 27.800 225.200 28.600 ;
        RECT 223.200 27.200 223.800 27.600 ;
        RECT 221.800 26.800 222.600 27.000 ;
        RECT 220.400 26.200 222.600 26.800 ;
        RECT 223.200 26.600 225.200 27.200 ;
        RECT 223.600 26.400 225.200 26.600 ;
        RECT 217.200 25.600 219.000 26.200 ;
        RECT 208.600 24.400 209.400 25.200 ;
        RECT 211.400 24.400 212.200 25.600 ;
        RECT 218.200 24.400 219.000 25.600 ;
        RECT 208.600 23.600 210.000 24.400 ;
        RECT 210.800 23.600 212.200 24.400 ;
        RECT 217.200 23.600 219.000 24.400 ;
        RECT 208.600 22.200 209.400 23.600 ;
        RECT 211.400 22.200 212.200 23.600 ;
        RECT 218.200 22.200 219.000 23.600 ;
        RECT 220.400 22.200 221.200 26.200 ;
        RECT 225.800 25.800 226.400 29.200 ;
        RECT 227.200 27.600 228.000 28.400 ;
        RECT 229.200 27.600 230.800 28.400 ;
        RECT 227.200 27.200 227.800 27.600 ;
        RECT 227.000 26.400 227.800 27.200 ;
        RECT 228.400 26.800 229.200 27.000 ;
        RECT 228.400 26.200 230.800 26.800 ;
        RECT 233.200 26.200 234.000 39.800 ;
        RECT 239.000 32.600 239.800 39.800 ;
        RECT 238.000 31.800 239.800 32.600 ;
        RECT 241.200 39.200 245.200 39.800 ;
        RECT 241.200 31.800 242.000 39.200 ;
        RECT 242.800 31.800 243.600 38.600 ;
        RECT 244.400 32.400 245.200 39.200 ;
        RECT 247.600 32.400 248.400 39.800 ;
        RECT 244.400 31.800 248.400 32.400 ;
        RECT 249.200 32.400 250.000 39.800 ;
        RECT 252.400 39.200 256.400 39.800 ;
        RECT 252.400 32.400 253.200 39.200 ;
        RECT 249.200 31.800 253.200 32.400 ;
        RECT 254.000 31.800 254.800 38.600 ;
        RECT 255.600 31.800 256.400 39.200 ;
        RECT 238.200 28.400 238.800 31.800 ;
        RECT 243.000 31.200 243.600 31.800 ;
        RECT 254.000 31.200 254.600 31.800 ;
        RECT 257.200 31.600 258.000 33.200 ;
        RECT 239.600 29.600 240.400 31.200 ;
        RECT 241.200 29.600 242.000 31.200 ;
        RECT 243.000 30.600 245.000 31.200 ;
        RECT 244.400 30.400 245.000 30.600 ;
        RECT 246.800 30.400 247.600 30.800 ;
        RECT 250.000 30.400 250.800 30.800 ;
        RECT 252.600 30.600 254.600 31.200 ;
        RECT 252.600 30.400 253.200 30.600 ;
        RECT 244.400 29.600 245.200 30.400 ;
        RECT 246.800 29.800 248.400 30.400 ;
        RECT 247.600 29.600 248.400 29.800 ;
        RECT 249.200 29.800 250.800 30.400 ;
        RECT 249.200 29.600 250.000 29.800 ;
        RECT 252.400 29.600 253.200 30.400 ;
        RECT 255.600 30.300 256.400 31.200 ;
        RECT 257.300 30.300 257.900 31.600 ;
        RECT 255.600 29.700 257.900 30.300 ;
        RECT 255.600 29.600 256.400 29.700 ;
        RECT 234.800 28.300 235.600 28.400 ;
        RECT 238.000 28.300 238.800 28.400 ;
        RECT 241.300 28.300 241.900 29.600 ;
        RECT 243.000 28.800 243.800 29.600 ;
        RECT 243.000 28.400 243.600 28.800 ;
        RECT 234.800 27.700 237.100 28.300 ;
        RECT 234.800 26.800 235.600 27.700 ;
        RECT 236.500 26.400 237.100 27.700 ;
        RECT 238.000 27.700 241.900 28.300 ;
        RECT 238.000 27.600 238.800 27.700 ;
        RECT 242.800 27.600 243.600 28.400 ;
        RECT 224.800 22.200 226.400 25.800 ;
        RECT 230.000 22.200 230.800 26.200 ;
        RECT 232.200 25.600 234.000 26.200 ;
        RECT 232.200 22.200 233.000 25.600 ;
        RECT 236.400 24.800 237.200 26.400 ;
        RECT 238.200 24.200 238.800 27.600 ;
        RECT 244.400 26.200 245.000 29.600 ;
        RECT 246.000 28.300 246.800 29.200 ;
        RECT 250.800 28.300 251.600 29.200 ;
        RECT 246.000 27.700 251.600 28.300 ;
        RECT 246.000 27.600 246.800 27.700 ;
        RECT 250.800 27.600 251.600 27.700 ;
        RECT 252.600 26.200 253.200 29.600 ;
        RECT 253.800 28.800 254.600 29.600 ;
        RECT 254.000 28.400 254.600 28.800 ;
        RECT 254.000 27.600 254.800 28.400 ;
        RECT 258.800 26.200 259.600 39.800 ;
        RECT 262.000 31.600 262.800 33.200 ;
        RECT 260.400 28.300 261.200 28.400 ;
        RECT 263.600 28.300 264.400 39.800 ;
        RECT 269.400 38.400 270.200 39.800 ;
        RECT 268.400 37.600 270.200 38.400 ;
        RECT 269.400 32.400 270.200 37.600 ;
        RECT 270.800 33.600 271.600 34.400 ;
        RECT 271.000 32.400 271.600 33.600 ;
        RECT 274.000 33.600 274.800 34.400 ;
        RECT 274.000 32.400 274.600 33.600 ;
        RECT 275.400 32.400 276.200 39.800 ;
        RECT 269.400 31.800 270.400 32.400 ;
        RECT 271.000 31.800 272.400 32.400 ;
        RECT 268.400 28.800 269.200 30.400 ;
        RECT 269.800 28.400 270.400 31.800 ;
        RECT 271.600 31.600 272.400 31.800 ;
        RECT 273.200 31.800 274.600 32.400 ;
        RECT 275.200 31.800 276.200 32.400 ;
        RECT 282.200 32.400 283.000 39.800 ;
        RECT 288.600 38.400 289.400 39.800 ;
        RECT 287.600 37.600 289.400 38.400 ;
        RECT 283.600 33.600 284.400 34.400 ;
        RECT 283.800 32.400 284.400 33.600 ;
        RECT 288.600 32.400 289.400 37.600 ;
        RECT 299.400 38.400 300.200 39.800 ;
        RECT 299.400 37.600 301.200 38.400 ;
        RECT 290.000 33.600 290.800 34.400 ;
        RECT 290.200 32.400 290.800 33.600 ;
        RECT 298.000 33.600 298.800 34.400 ;
        RECT 298.000 32.400 298.600 33.600 ;
        RECT 299.400 32.400 300.200 37.600 ;
        RECT 306.200 32.600 307.000 39.800 ;
        RECT 282.200 31.800 283.200 32.400 ;
        RECT 283.800 31.800 285.200 32.400 ;
        RECT 288.600 31.800 289.600 32.400 ;
        RECT 290.200 31.800 291.600 32.400 ;
        RECT 273.200 31.600 274.000 31.800 ;
        RECT 271.700 30.300 272.300 31.600 ;
        RECT 275.200 30.300 275.800 31.800 ;
        RECT 271.700 29.700 275.800 30.300 ;
        RECT 275.200 28.400 275.800 29.700 ;
        RECT 276.400 30.300 277.200 30.400 ;
        RECT 281.200 30.300 282.000 30.400 ;
        RECT 276.400 29.700 282.000 30.300 ;
        RECT 276.400 28.800 277.200 29.700 ;
        RECT 281.200 28.800 282.000 29.700 ;
        RECT 282.600 30.300 283.200 31.800 ;
        RECT 284.400 31.600 285.200 31.800 ;
        RECT 286.000 30.300 286.800 30.400 ;
        RECT 282.600 29.700 286.800 30.300 ;
        RECT 282.600 28.400 283.200 29.700 ;
        RECT 286.000 29.600 286.800 29.700 ;
        RECT 287.600 28.800 288.400 30.400 ;
        RECT 289.000 28.400 289.600 31.800 ;
        RECT 290.800 31.600 291.600 31.800 ;
        RECT 295.600 32.300 296.400 32.400 ;
        RECT 297.200 32.300 298.600 32.400 ;
        RECT 295.600 31.800 298.600 32.300 ;
        RECT 299.200 31.800 300.200 32.400 ;
        RECT 305.200 31.800 307.000 32.600 ;
        RECT 311.000 32.400 311.800 39.800 ;
        RECT 317.000 38.400 317.800 39.800 ;
        RECT 317.000 37.600 318.800 38.400 ;
        RECT 312.400 33.600 313.200 34.400 ;
        RECT 312.600 32.400 313.200 33.600 ;
        RECT 315.600 33.600 316.400 34.400 ;
        RECT 315.600 32.400 316.200 33.600 ;
        RECT 317.000 32.400 317.800 37.600 ;
        RECT 311.000 31.800 312.000 32.400 ;
        RECT 312.600 31.800 314.000 32.400 ;
        RECT 295.600 31.700 298.000 31.800 ;
        RECT 295.600 31.600 296.400 31.700 ;
        RECT 297.200 31.600 298.000 31.700 ;
        RECT 299.200 28.400 299.800 31.800 ;
        RECT 300.400 28.800 301.200 30.400 ;
        RECT 305.400 28.400 306.000 31.800 ;
        RECT 306.800 30.300 307.600 31.200 ;
        RECT 308.400 30.300 309.200 30.400 ;
        RECT 306.800 29.700 309.200 30.300 ;
        RECT 306.800 29.600 307.600 29.700 ;
        RECT 308.400 29.600 309.200 29.700 ;
        RECT 310.000 28.800 310.800 30.400 ;
        RECT 311.400 30.300 312.000 31.800 ;
        RECT 313.200 31.600 314.000 31.800 ;
        RECT 314.800 31.800 316.200 32.400 ;
        RECT 316.800 31.800 317.800 32.400 ;
        RECT 314.800 31.600 315.600 31.800 ;
        RECT 314.900 30.300 315.500 31.600 ;
        RECT 311.400 29.700 315.500 30.300 ;
        RECT 311.400 28.400 312.000 29.700 ;
        RECT 316.800 28.400 317.400 31.800 ;
        RECT 318.000 28.800 318.800 30.400 ;
        RECT 260.400 27.700 264.400 28.300 ;
        RECT 260.400 26.800 261.200 27.700 ;
        RECT 263.600 26.200 264.400 27.700 ;
        RECT 265.200 26.800 266.000 28.400 ;
        RECT 266.800 28.200 267.600 28.400 ;
        RECT 266.800 27.600 268.400 28.200 ;
        RECT 269.800 27.600 272.400 28.400 ;
        RECT 273.200 27.600 275.800 28.400 ;
        RECT 278.000 28.300 278.800 28.400 ;
        RECT 279.600 28.300 280.400 28.400 ;
        RECT 278.000 28.200 280.400 28.300 ;
        RECT 277.200 27.700 281.200 28.200 ;
        RECT 277.200 27.600 278.800 27.700 ;
        RECT 279.600 27.600 281.200 27.700 ;
        RECT 282.600 27.600 285.200 28.400 ;
        RECT 286.000 28.200 286.800 28.400 ;
        RECT 286.000 27.600 287.600 28.200 ;
        RECT 289.000 27.600 291.600 28.400 ;
        RECT 297.200 27.600 299.800 28.400 ;
        RECT 302.000 28.200 302.800 28.400 ;
        RECT 301.200 27.600 302.800 28.200 ;
        RECT 305.200 27.600 306.000 28.400 ;
        RECT 308.400 28.200 309.200 28.400 ;
        RECT 308.400 27.600 310.000 28.200 ;
        RECT 311.400 27.600 314.000 28.400 ;
        RECT 314.800 27.600 317.400 28.400 ;
        RECT 319.600 28.200 320.400 28.400 ;
        RECT 318.800 27.600 320.400 28.200 ;
        RECT 267.600 27.200 268.400 27.600 ;
        RECT 267.000 26.200 270.600 26.600 ;
        RECT 271.600 26.200 272.200 27.600 ;
        RECT 273.400 26.200 274.000 27.600 ;
        RECT 277.200 27.200 278.000 27.600 ;
        RECT 280.400 27.200 281.200 27.600 ;
        RECT 275.000 26.200 278.600 26.600 ;
        RECT 279.800 26.200 283.400 26.600 ;
        RECT 284.400 26.200 285.000 27.600 ;
        RECT 286.800 27.200 287.600 27.600 ;
        RECT 286.200 26.200 289.800 26.600 ;
        RECT 290.800 26.200 291.400 27.600 ;
        RECT 297.400 26.200 298.000 27.600 ;
        RECT 301.200 27.200 302.000 27.600 ;
        RECT 299.000 26.200 302.600 26.600 ;
        RECT 238.000 22.200 238.800 24.200 ;
        RECT 243.800 22.200 245.400 26.200 ;
        RECT 252.200 22.200 253.800 26.200 ;
        RECT 257.800 25.600 259.600 26.200 ;
        RECT 262.600 25.600 264.400 26.200 ;
        RECT 266.800 26.000 270.800 26.200 ;
        RECT 257.800 24.400 258.600 25.600 ;
        RECT 257.200 23.600 258.600 24.400 ;
        RECT 257.800 22.200 258.600 23.600 ;
        RECT 262.600 22.200 263.400 25.600 ;
        RECT 266.800 22.200 267.600 26.000 ;
        RECT 270.000 22.200 270.800 26.000 ;
        RECT 271.600 22.200 272.400 26.200 ;
        RECT 273.200 22.200 274.000 26.200 ;
        RECT 274.800 26.000 278.800 26.200 ;
        RECT 274.800 22.200 275.600 26.000 ;
        RECT 278.000 22.200 278.800 26.000 ;
        RECT 279.600 26.000 283.600 26.200 ;
        RECT 279.600 22.200 280.400 26.000 ;
        RECT 282.800 22.200 283.600 26.000 ;
        RECT 284.400 22.200 285.200 26.200 ;
        RECT 286.000 26.000 290.000 26.200 ;
        RECT 286.000 22.200 286.800 26.000 ;
        RECT 289.200 22.200 290.000 26.000 ;
        RECT 290.800 22.200 291.600 26.200 ;
        RECT 297.200 22.200 298.000 26.200 ;
        RECT 298.800 26.000 302.800 26.200 ;
        RECT 298.800 22.200 299.600 26.000 ;
        RECT 302.000 22.200 302.800 26.000 ;
        RECT 303.600 24.800 304.400 26.400 ;
        RECT 305.400 24.400 306.000 27.600 ;
        RECT 309.200 27.200 310.000 27.600 ;
        RECT 308.600 26.200 312.200 26.600 ;
        RECT 313.200 26.200 313.800 27.600 ;
        RECT 315.000 26.200 315.600 27.600 ;
        RECT 318.800 27.200 319.600 27.600 ;
        RECT 316.600 26.200 320.200 26.600 ;
        RECT 305.200 22.200 306.000 24.400 ;
        RECT 308.400 26.000 312.400 26.200 ;
        RECT 308.400 22.200 309.200 26.000 ;
        RECT 311.600 22.200 312.400 26.000 ;
        RECT 313.200 22.200 314.000 26.200 ;
        RECT 314.800 22.200 315.600 26.200 ;
        RECT 316.400 26.000 320.400 26.200 ;
        RECT 316.400 22.200 317.200 26.000 ;
        RECT 319.600 22.200 320.400 26.000 ;
        RECT 321.200 22.200 322.000 39.800 ;
        RECT 322.800 24.800 323.600 26.400 ;
        RECT 324.400 24.800 325.200 26.400 ;
        RECT 326.000 22.200 326.800 39.800 ;
        RECT 330.200 32.600 331.000 39.800 ;
        RECT 329.200 31.800 331.000 32.600 ;
        RECT 333.200 33.600 334.000 34.400 ;
        RECT 333.200 32.400 333.800 33.600 ;
        RECT 334.600 32.400 335.400 39.800 ;
        RECT 332.400 31.800 333.800 32.400 ;
        RECT 334.400 31.800 335.400 32.400 ;
        RECT 339.400 32.600 340.200 39.800 ;
        RECT 339.400 31.800 341.200 32.600 ;
        RECT 343.600 31.800 344.400 39.800 ;
        RECT 345.200 32.400 346.000 39.800 ;
        RECT 348.400 32.400 349.200 39.800 ;
        RECT 345.200 31.800 349.200 32.400 ;
        RECT 329.400 30.400 330.000 31.800 ;
        RECT 332.400 31.600 333.200 31.800 ;
        RECT 329.200 29.600 330.000 30.400 ;
        RECT 330.800 29.600 331.600 31.200 ;
        RECT 334.400 30.400 335.000 31.800 ;
        RECT 334.000 29.600 335.000 30.400 ;
        RECT 329.400 28.400 330.000 29.600 ;
        RECT 334.400 28.400 335.000 29.600 ;
        RECT 335.600 30.300 336.400 30.400 ;
        RECT 338.800 30.300 339.600 31.200 ;
        RECT 335.600 29.700 339.600 30.300 ;
        RECT 335.600 28.800 336.400 29.700 ;
        RECT 338.800 29.600 339.600 29.700 ;
        RECT 340.400 28.400 341.000 31.800 ;
        RECT 343.800 30.400 344.400 31.800 ;
        RECT 350.000 31.600 350.800 33.200 ;
        RECT 351.600 32.300 352.400 39.800 ;
        RECT 357.400 32.400 358.200 39.800 ;
        RECT 358.800 33.600 359.600 34.400 ;
        RECT 359.000 32.400 359.600 33.600 ;
        RECT 353.200 32.300 354.000 32.400 ;
        RECT 351.600 31.700 354.000 32.300 ;
        RECT 357.400 31.800 358.400 32.400 ;
        RECT 359.000 31.800 360.400 32.400 ;
        RECT 347.600 30.400 348.400 30.800 ;
        RECT 343.600 29.800 346.000 30.400 ;
        RECT 347.600 30.300 349.200 30.400 ;
        RECT 350.100 30.300 350.700 31.600 ;
        RECT 347.600 29.800 350.700 30.300 ;
        RECT 343.600 29.600 344.400 29.800 ;
        RECT 329.200 27.600 330.000 28.400 ;
        RECT 332.400 27.600 335.000 28.400 ;
        RECT 337.200 28.200 338.000 28.400 ;
        RECT 336.400 27.600 338.000 28.200 ;
        RECT 340.400 28.300 341.200 28.400 ;
        RECT 343.600 28.300 344.400 28.400 ;
        RECT 340.400 27.700 344.400 28.300 ;
        RECT 340.400 27.600 341.200 27.700 ;
        RECT 343.600 27.600 344.400 27.700 ;
        RECT 327.600 24.800 328.400 26.400 ;
        RECT 329.400 24.200 330.000 27.600 ;
        RECT 332.600 26.200 333.200 27.600 ;
        RECT 336.400 27.200 337.200 27.600 ;
        RECT 334.200 26.200 337.800 26.600 ;
        RECT 329.200 22.200 330.000 24.200 ;
        RECT 332.400 22.200 333.200 26.200 ;
        RECT 334.000 26.000 338.000 26.200 ;
        RECT 334.000 22.200 334.800 26.000 ;
        RECT 337.200 22.200 338.000 26.000 ;
        RECT 340.400 24.200 341.000 27.600 ;
        RECT 342.000 26.300 342.800 26.400 ;
        RECT 343.600 26.300 344.400 26.400 ;
        RECT 342.000 25.700 344.400 26.300 ;
        RECT 345.400 26.200 346.000 29.800 ;
        RECT 348.400 29.700 350.700 29.800 ;
        RECT 348.400 29.600 349.200 29.700 ;
        RECT 346.800 27.600 347.600 29.200 ;
        RECT 351.600 26.200 352.400 31.700 ;
        RECT 353.200 31.600 354.000 31.700 ;
        RECT 356.400 28.800 357.200 30.400 ;
        RECT 357.800 28.400 358.400 31.800 ;
        RECT 359.600 31.600 360.400 31.800 ;
        RECT 353.200 28.300 354.000 28.400 ;
        RECT 354.800 28.300 355.600 28.400 ;
        RECT 353.200 28.200 355.600 28.300 ;
        RECT 357.800 28.300 360.400 28.400 ;
        RECT 361.200 28.300 362.000 28.400 ;
        RECT 353.200 27.700 356.400 28.200 ;
        RECT 353.200 26.800 354.000 27.700 ;
        RECT 354.800 27.600 356.400 27.700 ;
        RECT 357.800 27.700 362.000 28.300 ;
        RECT 357.800 27.600 360.400 27.700 ;
        RECT 361.200 27.600 362.000 27.700 ;
        RECT 362.800 28.300 363.600 39.800 ;
        RECT 364.400 32.400 365.200 39.800 ;
        RECT 366.000 32.400 366.800 32.600 ;
        RECT 368.800 32.400 370.400 39.800 ;
        RECT 364.400 31.800 366.800 32.400 ;
        RECT 368.400 31.800 370.400 32.400 ;
        RECT 372.600 32.400 373.400 32.600 ;
        RECT 374.000 32.400 374.800 39.800 ;
        RECT 372.600 31.800 374.800 32.400 ;
        RECT 368.400 30.400 369.000 31.800 ;
        RECT 372.600 31.200 373.200 31.800 ;
        RECT 369.800 30.600 373.200 31.200 ;
        RECT 375.600 31.400 376.400 39.800 ;
        RECT 380.000 36.400 380.800 39.800 ;
        RECT 378.800 35.800 380.800 36.400 ;
        RECT 384.400 35.800 385.200 39.800 ;
        RECT 388.600 35.800 389.800 39.800 ;
        RECT 378.800 35.000 379.600 35.800 ;
        RECT 384.400 35.200 385.000 35.800 ;
        RECT 382.200 34.600 385.800 35.200 ;
        RECT 388.400 35.000 389.200 35.800 ;
        RECT 382.200 34.400 383.000 34.600 ;
        RECT 385.000 34.400 385.800 34.600 ;
        RECT 378.800 33.000 379.600 33.200 ;
        RECT 383.400 33.000 384.200 33.200 ;
        RECT 378.800 32.400 384.200 33.000 ;
        RECT 384.800 33.000 387.000 33.600 ;
        RECT 384.800 31.800 385.400 33.000 ;
        RECT 386.200 32.800 387.000 33.000 ;
        RECT 388.600 33.200 390.000 34.000 ;
        RECT 388.600 32.200 389.200 33.200 ;
        RECT 380.600 31.400 385.400 31.800 ;
        RECT 375.600 31.200 385.400 31.400 ;
        RECT 386.800 31.600 389.200 32.200 ;
        RECT 375.600 31.000 381.400 31.200 ;
        RECT 375.600 30.800 381.200 31.000 ;
        RECT 369.800 30.400 370.600 30.600 ;
        RECT 367.600 29.800 369.000 30.400 ;
        RECT 382.000 30.200 382.800 30.400 ;
        RECT 372.000 29.800 372.800 30.000 ;
        RECT 367.600 29.600 369.400 29.800 ;
        RECT 368.400 29.200 369.400 29.600 ;
        RECT 364.400 28.300 366.000 28.400 ;
        RECT 362.800 27.700 366.000 28.300 ;
        RECT 355.600 27.200 356.400 27.600 ;
        RECT 355.000 26.200 358.600 26.600 ;
        RECT 359.600 26.200 360.200 27.600 ;
        RECT 342.000 24.800 342.800 25.700 ;
        RECT 343.600 25.600 344.400 25.700 ;
        RECT 343.800 24.800 344.600 25.600 ;
        RECT 340.400 22.200 341.200 24.200 ;
        RECT 345.200 22.200 346.000 26.200 ;
        RECT 350.600 25.600 352.400 26.200 ;
        RECT 354.800 26.000 358.800 26.200 ;
        RECT 350.600 22.200 351.400 25.600 ;
        RECT 354.800 22.200 355.600 26.000 ;
        RECT 358.000 22.200 358.800 26.000 ;
        RECT 359.600 22.200 360.400 26.200 ;
        RECT 361.200 24.800 362.000 26.400 ;
        RECT 362.800 22.200 363.600 27.700 ;
        RECT 364.400 27.600 366.000 27.700 ;
        RECT 367.200 27.600 368.000 28.400 ;
        RECT 367.400 27.200 368.000 27.600 ;
        RECT 366.000 26.800 366.800 27.000 ;
        RECT 364.400 26.200 366.800 26.800 ;
        RECT 367.400 26.400 368.200 27.200 ;
        RECT 364.400 22.200 365.200 26.200 ;
        RECT 368.800 25.800 369.400 29.200 ;
        RECT 370.200 29.200 372.800 29.800 ;
        RECT 377.800 29.600 382.800 30.200 ;
        RECT 385.200 30.300 386.000 30.400 ;
        RECT 386.800 30.300 387.400 31.600 ;
        RECT 393.200 31.200 394.000 39.800 ;
        RECT 394.800 32.400 395.600 39.800 ;
        RECT 398.000 32.800 398.800 39.800 ;
        RECT 394.800 31.800 397.400 32.400 ;
        RECT 398.000 31.800 399.000 32.800 ;
        RECT 401.200 32.400 402.000 39.800 ;
        RECT 402.600 32.400 403.400 32.600 ;
        RECT 401.200 31.800 403.400 32.400 ;
        RECT 405.600 32.400 407.200 39.800 ;
        RECT 409.200 32.400 410.000 32.600 ;
        RECT 410.800 32.400 411.600 39.800 ;
        RECT 405.600 31.800 407.600 32.400 ;
        RECT 409.200 31.800 411.600 32.400 ;
        RECT 389.800 30.600 394.000 31.200 ;
        RECT 389.800 30.400 390.600 30.600 ;
        RECT 385.200 29.700 387.500 30.300 ;
        RECT 391.400 29.800 392.200 30.000 ;
        RECT 385.200 29.600 386.000 29.700 ;
        RECT 377.800 29.400 378.600 29.600 ;
        RECT 380.400 29.400 381.200 29.600 ;
        RECT 370.200 28.600 370.800 29.200 ;
        RECT 370.000 27.800 370.800 28.600 ;
        RECT 379.400 28.400 380.200 28.600 ;
        RECT 386.800 28.400 387.400 29.700 ;
        RECT 388.400 29.200 392.200 29.800 ;
        RECT 388.400 29.000 389.200 29.200 ;
        RECT 373.200 28.200 374.800 28.400 ;
        RECT 371.400 27.600 374.800 28.200 ;
        RECT 376.400 27.800 387.400 28.400 ;
        RECT 376.400 27.600 378.000 27.800 ;
        RECT 371.400 27.200 372.000 27.600 ;
        RECT 370.000 26.600 372.000 27.200 ;
        RECT 372.600 26.800 373.400 27.000 ;
        RECT 370.000 26.400 371.600 26.600 ;
        RECT 372.600 26.200 374.800 26.800 ;
        RECT 368.800 22.200 370.400 25.800 ;
        RECT 374.000 22.200 374.800 26.200 ;
        RECT 375.600 22.200 376.400 27.000 ;
        RECT 380.600 25.600 381.200 27.800 ;
        RECT 386.200 27.600 387.000 27.800 ;
        RECT 393.200 27.200 394.000 30.600 ;
        RECT 394.800 29.600 395.800 30.400 ;
        RECT 395.000 28.800 395.800 29.600 ;
        RECT 396.800 29.800 397.400 31.800 ;
        RECT 396.800 29.000 397.800 29.800 ;
        RECT 396.800 27.400 397.400 29.000 ;
        RECT 398.400 28.400 399.000 31.800 ;
        RECT 402.800 31.200 403.400 31.800 ;
        RECT 402.800 30.600 406.200 31.200 ;
        RECT 405.400 30.400 406.200 30.600 ;
        RECT 407.000 30.400 407.600 31.800 ;
        RECT 407.000 30.300 408.400 30.400 ;
        RECT 412.400 30.300 413.200 30.400 ;
        RECT 403.200 29.800 404.000 30.000 ;
        RECT 407.000 29.800 413.200 30.300 ;
        RECT 403.200 29.200 405.800 29.800 ;
        RECT 405.200 28.600 405.800 29.200 ;
        RECT 406.600 29.700 413.200 29.800 ;
        RECT 406.600 29.600 408.400 29.700 ;
        RECT 412.400 29.600 413.200 29.700 ;
        RECT 406.600 29.200 407.600 29.600 ;
        RECT 398.000 28.300 399.000 28.400 ;
        RECT 401.200 28.300 402.800 28.400 ;
        RECT 398.000 28.200 402.800 28.300 ;
        RECT 398.000 27.700 404.600 28.200 ;
        RECT 405.200 27.800 406.000 28.600 ;
        RECT 398.000 27.600 399.000 27.700 ;
        RECT 401.200 27.600 404.600 27.700 ;
        RECT 390.200 26.600 394.000 27.200 ;
        RECT 390.200 26.400 391.000 26.600 ;
        RECT 378.800 24.200 379.600 25.000 ;
        RECT 380.400 24.800 381.200 25.600 ;
        RECT 382.200 25.400 383.000 25.600 ;
        RECT 382.200 24.800 385.000 25.400 ;
        RECT 384.400 24.200 385.000 24.800 ;
        RECT 388.400 24.200 389.200 25.000 ;
        RECT 378.800 23.600 380.800 24.200 ;
        RECT 380.000 22.200 380.800 23.600 ;
        RECT 384.400 22.200 385.200 24.200 ;
        RECT 388.400 23.600 389.800 24.200 ;
        RECT 388.600 22.200 389.800 23.600 ;
        RECT 393.200 22.200 394.000 26.600 ;
        RECT 394.800 26.800 397.400 27.400 ;
        RECT 394.800 22.200 395.600 26.800 ;
        RECT 398.400 26.200 399.000 27.600 ;
        RECT 404.000 27.200 404.600 27.600 ;
        RECT 402.600 26.800 403.400 27.000 ;
        RECT 398.000 25.600 399.000 26.200 ;
        RECT 401.200 26.200 403.400 26.800 ;
        RECT 404.000 26.600 406.000 27.200 ;
        RECT 404.400 26.400 406.000 26.600 ;
        RECT 398.000 22.200 398.800 25.600 ;
        RECT 401.200 22.200 402.000 26.200 ;
        RECT 406.600 25.800 407.200 29.200 ;
        RECT 408.000 27.600 408.800 28.400 ;
        RECT 410.000 27.600 411.600 28.400 ;
        RECT 408.000 27.200 408.600 27.600 ;
        RECT 407.800 26.400 408.600 27.200 ;
        RECT 409.200 26.800 410.000 27.000 ;
        RECT 412.400 26.800 413.200 28.400 ;
        RECT 409.200 26.200 411.600 26.800 ;
        RECT 405.600 22.200 407.200 25.800 ;
        RECT 410.800 22.200 411.600 26.200 ;
        RECT 414.000 26.200 414.800 39.800 ;
        RECT 419.800 38.400 420.600 39.800 ;
        RECT 418.800 37.600 420.600 38.400 ;
        RECT 415.600 31.600 416.400 33.200 ;
        RECT 419.800 32.400 420.600 37.600 ;
        RECT 421.200 33.600 422.000 34.400 ;
        RECT 421.400 32.400 422.000 33.600 ;
        RECT 419.800 31.800 420.800 32.400 ;
        RECT 421.400 31.800 422.800 32.400 ;
        RECT 418.800 28.800 419.600 30.400 ;
        RECT 420.200 28.400 420.800 31.800 ;
        RECT 422.000 31.600 422.800 31.800 ;
        RECT 422.000 30.300 422.800 30.400 ;
        RECT 422.000 29.700 424.300 30.300 ;
        RECT 422.000 29.600 422.800 29.700 ;
        RECT 423.700 28.400 424.300 29.700 ;
        RECT 417.200 28.200 418.000 28.400 ;
        RECT 417.200 27.600 418.800 28.200 ;
        RECT 420.200 27.600 422.800 28.400 ;
        RECT 418.000 27.200 418.800 27.600 ;
        RECT 417.400 26.200 421.000 26.600 ;
        RECT 422.000 26.200 422.600 27.600 ;
        RECT 423.600 26.800 424.400 28.400 ;
        RECT 425.200 26.200 426.000 39.800 ;
        RECT 426.800 32.300 427.600 33.200 ;
        RECT 430.000 32.300 430.800 39.800 ;
        RECT 435.800 36.400 436.600 39.800 ;
        RECT 435.800 35.600 437.200 36.400 ;
        RECT 426.800 31.700 430.800 32.300 ;
        RECT 426.800 31.600 427.600 31.700 ;
        RECT 428.400 26.800 429.200 28.400 ;
        RECT 430.000 28.300 430.800 31.700 ;
        RECT 431.600 31.600 432.400 33.200 ;
        RECT 435.800 32.600 436.600 35.600 ;
        RECT 434.800 31.800 436.600 32.600 ;
        RECT 440.600 32.400 441.400 39.800 ;
        RECT 442.000 33.600 442.800 34.400 ;
        RECT 442.200 32.400 442.800 33.600 ;
        RECT 440.600 31.800 441.600 32.400 ;
        RECT 442.200 31.800 443.600 32.400 ;
        RECT 435.000 28.400 435.600 31.800 ;
        RECT 436.400 30.300 437.200 31.200 ;
        RECT 436.400 29.700 438.700 30.300 ;
        RECT 436.400 29.600 437.200 29.700 ;
        RECT 438.100 28.400 438.700 29.700 ;
        RECT 439.600 28.800 440.400 30.400 ;
        RECT 441.000 30.300 441.600 31.800 ;
        RECT 442.800 31.600 443.600 31.800 ;
        RECT 449.200 30.300 450.000 30.400 ;
        RECT 441.000 29.700 450.000 30.300 ;
        RECT 441.000 28.400 441.600 29.700 ;
        RECT 449.200 29.600 450.000 29.700 ;
        RECT 433.200 28.300 434.000 28.400 ;
        RECT 430.000 27.700 434.000 28.300 ;
        RECT 430.000 26.200 430.800 27.700 ;
        RECT 433.200 27.600 434.000 27.700 ;
        RECT 434.800 27.600 435.600 28.400 ;
        RECT 438.000 28.200 438.800 28.400 ;
        RECT 438.000 27.600 439.600 28.200 ;
        RECT 441.000 27.600 443.600 28.400 ;
        RECT 444.400 28.300 445.200 28.400 ;
        RECT 449.200 28.300 450.000 28.400 ;
        RECT 444.400 27.700 450.000 28.300 ;
        RECT 444.400 27.600 445.200 27.700 ;
        RECT 414.000 25.600 415.800 26.200 ;
        RECT 415.000 22.200 415.800 25.600 ;
        RECT 417.200 26.000 421.200 26.200 ;
        RECT 417.200 22.200 418.000 26.000 ;
        RECT 420.400 22.200 421.200 26.000 ;
        RECT 422.000 22.200 422.800 26.200 ;
        RECT 425.200 25.600 427.000 26.200 ;
        RECT 430.000 25.600 431.800 26.200 ;
        RECT 426.200 24.400 427.000 25.600 ;
        RECT 425.200 23.600 427.000 24.400 ;
        RECT 426.200 22.200 427.000 23.600 ;
        RECT 431.000 22.200 431.800 25.600 ;
        RECT 433.200 24.800 434.000 26.400 ;
        RECT 435.000 24.200 435.600 27.600 ;
        RECT 438.800 27.200 439.600 27.600 ;
        RECT 438.200 26.200 441.800 26.600 ;
        RECT 442.800 26.200 443.400 27.600 ;
        RECT 449.200 26.800 450.000 27.700 ;
        RECT 450.800 28.300 451.600 39.800 ;
        RECT 452.400 31.600 453.200 33.200 ;
        RECT 454.000 28.300 454.800 28.400 ;
        RECT 450.800 27.700 454.800 28.300 ;
        RECT 450.800 26.200 451.600 27.700 ;
        RECT 454.000 26.800 454.800 27.700 ;
        RECT 455.600 26.200 456.400 39.800 ;
        RECT 459.600 33.600 460.400 34.400 ;
        RECT 457.200 31.600 458.000 33.200 ;
        RECT 459.600 32.400 460.200 33.600 ;
        RECT 461.000 32.400 461.800 39.800 ;
        RECT 458.800 31.800 460.200 32.400 ;
        RECT 458.800 31.600 459.600 31.800 ;
        RECT 460.800 31.600 462.800 32.400 ;
        RECT 465.200 31.600 466.000 33.200 ;
        RECT 460.800 28.400 461.400 31.600 ;
        RECT 462.000 28.800 462.800 30.400 ;
        RECT 458.800 27.600 461.400 28.400 ;
        RECT 463.600 28.300 464.400 28.400 ;
        RECT 466.800 28.300 467.600 39.800 ;
        RECT 470.000 39.200 474.000 39.800 ;
        RECT 470.000 31.800 470.800 39.200 ;
        RECT 471.600 31.800 472.400 38.600 ;
        RECT 473.200 32.400 474.000 39.200 ;
        RECT 476.400 32.400 477.200 39.800 ;
        RECT 473.200 31.800 477.200 32.400 ;
        RECT 478.000 39.200 482.000 39.800 ;
        RECT 478.000 31.800 478.800 39.200 ;
        RECT 479.600 31.800 480.400 38.600 ;
        RECT 481.200 32.400 482.000 39.200 ;
        RECT 484.400 32.400 485.200 39.800 ;
        RECT 488.600 38.400 489.400 39.800 ;
        RECT 487.600 37.600 489.400 38.400 ;
        RECT 481.200 31.800 485.200 32.400 ;
        RECT 488.600 32.400 489.400 37.600 ;
        RECT 494.600 38.400 495.400 39.800 ;
        RECT 494.600 37.600 496.400 38.400 ;
        RECT 490.000 33.600 490.800 34.400 ;
        RECT 490.200 32.400 490.800 33.600 ;
        RECT 493.200 33.600 494.000 34.400 ;
        RECT 493.200 32.400 493.800 33.600 ;
        RECT 494.600 32.400 495.400 37.600 ;
        RECT 499.600 33.600 500.400 34.400 ;
        RECT 499.600 32.400 500.200 33.600 ;
        RECT 501.000 32.400 501.800 39.800 ;
        RECT 488.600 31.800 489.600 32.400 ;
        RECT 490.200 31.800 491.600 32.400 ;
        RECT 471.800 31.200 472.400 31.800 ;
        RECT 479.800 31.200 480.400 31.800 ;
        RECT 470.000 29.600 470.800 31.200 ;
        RECT 471.800 30.600 473.800 31.200 ;
        RECT 473.200 30.400 473.800 30.600 ;
        RECT 475.600 30.400 476.400 30.800 ;
        RECT 473.200 29.600 474.000 30.400 ;
        RECT 475.600 29.800 477.200 30.400 ;
        RECT 476.400 29.600 477.200 29.800 ;
        RECT 478.000 29.600 478.800 31.200 ;
        RECT 479.800 30.600 481.800 31.200 ;
        RECT 481.200 30.400 481.800 30.600 ;
        RECT 483.600 30.400 484.400 30.800 ;
        RECT 481.200 29.600 482.000 30.400 ;
        RECT 483.600 29.800 485.200 30.400 ;
        RECT 484.400 29.600 485.200 29.800 ;
        RECT 486.000 30.300 486.800 30.400 ;
        RECT 487.600 30.300 488.400 30.400 ;
        RECT 486.000 29.700 488.400 30.300 ;
        RECT 486.000 29.600 486.800 29.700 ;
        RECT 471.800 28.800 472.600 29.600 ;
        RECT 471.800 28.400 472.400 28.800 ;
        RECT 463.600 28.200 467.600 28.300 ;
        RECT 462.800 27.700 467.600 28.200 ;
        RECT 462.800 27.600 464.400 27.700 ;
        RECT 459.000 26.200 459.600 27.600 ;
        RECT 462.800 27.200 463.600 27.600 ;
        RECT 460.600 26.200 464.200 26.600 ;
        RECT 466.800 26.200 467.600 27.700 ;
        RECT 468.400 26.800 469.200 28.400 ;
        RECT 471.600 27.600 472.400 28.400 ;
        RECT 473.200 26.200 473.800 29.600 ;
        RECT 474.800 27.600 475.600 29.200 ;
        RECT 479.800 28.800 480.600 29.600 ;
        RECT 479.800 28.400 480.400 28.800 ;
        RECT 479.600 27.600 480.400 28.400 ;
        RECT 481.200 26.200 481.800 29.600 ;
        RECT 482.800 27.600 483.600 29.200 ;
        RECT 487.600 28.800 488.400 29.700 ;
        RECT 489.000 28.400 489.600 31.800 ;
        RECT 490.800 31.600 491.600 31.800 ;
        RECT 492.400 31.800 493.800 32.400 ;
        RECT 494.400 31.800 495.400 32.400 ;
        RECT 498.800 31.800 500.200 32.400 ;
        RECT 500.800 31.800 501.800 32.400 ;
        RECT 505.200 32.400 506.000 39.800 ;
        RECT 508.400 39.200 512.400 39.800 ;
        RECT 508.400 32.400 509.200 39.200 ;
        RECT 505.200 31.800 509.200 32.400 ;
        RECT 510.000 31.800 510.800 38.600 ;
        RECT 511.600 31.800 512.400 39.200 ;
        RECT 492.400 31.600 493.200 31.800 ;
        RECT 494.400 28.400 495.000 31.800 ;
        RECT 498.800 31.600 499.600 31.800 ;
        RECT 495.600 28.800 496.400 30.400 ;
        RECT 500.800 28.400 501.400 31.800 ;
        RECT 510.000 31.200 510.600 31.800 ;
        RECT 506.000 30.400 506.800 30.800 ;
        RECT 508.600 30.600 510.600 31.200 ;
        RECT 508.600 30.400 509.200 30.600 ;
        RECT 502.000 28.800 502.800 30.400 ;
        RECT 505.200 29.800 506.800 30.400 ;
        RECT 505.200 29.600 506.000 29.800 ;
        RECT 508.400 29.600 509.200 30.400 ;
        RECT 511.600 30.300 512.400 31.200 ;
        RECT 513.200 30.300 514.000 39.800 ;
        RECT 516.400 32.400 517.200 39.800 ;
        RECT 519.600 39.200 523.600 39.800 ;
        RECT 519.600 32.400 520.400 39.200 ;
        RECT 516.400 31.800 520.400 32.400 ;
        RECT 521.200 31.800 522.000 38.600 ;
        RECT 522.800 31.800 523.600 39.200 ;
        RECT 527.000 32.600 527.800 39.800 ;
        RECT 526.000 31.800 527.800 32.600 ;
        RECT 529.200 32.400 530.000 39.800 ;
        RECT 533.600 38.400 535.200 39.800 ;
        RECT 532.400 37.600 535.200 38.400 ;
        RECT 530.800 32.400 531.600 32.600 ;
        RECT 533.600 32.400 535.200 37.600 ;
        RECT 529.200 31.800 531.600 32.400 ;
        RECT 533.200 31.800 535.200 32.400 ;
        RECT 537.400 32.400 538.200 32.600 ;
        RECT 538.800 32.400 539.600 39.800 ;
        RECT 537.400 31.800 539.600 32.400 ;
        RECT 541.000 32.600 541.800 39.800 ;
        RECT 541.000 31.800 542.800 32.600 ;
        RECT 545.200 31.800 546.000 39.800 ;
        RECT 546.800 32.400 547.600 39.800 ;
        RECT 550.000 32.400 550.800 39.800 ;
        RECT 546.800 31.800 550.800 32.400 ;
        RECT 521.200 31.200 521.800 31.800 ;
        RECT 517.200 30.400 518.000 30.800 ;
        RECT 519.800 30.600 521.800 31.200 ;
        RECT 519.800 30.400 520.400 30.600 ;
        RECT 511.600 29.700 514.000 30.300 ;
        RECT 511.600 29.600 512.400 29.700 ;
        RECT 486.000 28.200 486.800 28.400 ;
        RECT 486.000 27.600 487.600 28.200 ;
        RECT 489.000 27.600 491.600 28.400 ;
        RECT 492.400 27.600 495.000 28.400 ;
        RECT 497.200 28.200 498.000 28.400 ;
        RECT 496.400 27.600 498.000 28.200 ;
        RECT 498.800 27.600 501.400 28.400 ;
        RECT 503.600 28.200 504.400 28.400 ;
        RECT 502.800 27.600 504.400 28.200 ;
        RECT 506.800 27.600 507.600 29.200 ;
        RECT 486.800 27.200 487.600 27.600 ;
        RECT 486.200 26.200 489.800 26.600 ;
        RECT 490.800 26.200 491.400 27.600 ;
        RECT 492.600 26.200 493.200 27.600 ;
        RECT 496.400 27.200 497.200 27.600 ;
        RECT 494.200 26.200 497.800 26.600 ;
        RECT 499.000 26.200 499.600 27.600 ;
        RECT 502.800 27.200 503.600 27.600 ;
        RECT 500.600 26.200 504.200 26.600 ;
        RECT 508.600 26.200 509.200 29.600 ;
        RECT 509.800 28.800 510.600 29.600 ;
        RECT 510.000 28.400 510.600 28.800 ;
        RECT 510.000 27.600 510.800 28.400 ;
        RECT 434.800 22.200 435.600 24.200 ;
        RECT 438.000 26.000 442.000 26.200 ;
        RECT 438.000 22.200 438.800 26.000 ;
        RECT 441.200 22.200 442.000 26.000 ;
        RECT 442.800 22.200 443.600 26.200 ;
        RECT 450.800 25.600 452.600 26.200 ;
        RECT 455.600 25.600 457.400 26.200 ;
        RECT 451.800 22.200 452.600 25.600 ;
        RECT 456.600 22.200 457.400 25.600 ;
        RECT 458.800 22.200 459.600 26.200 ;
        RECT 460.400 26.000 464.400 26.200 ;
        RECT 460.400 22.200 461.200 26.000 ;
        RECT 463.600 22.200 464.400 26.000 ;
        RECT 465.800 25.600 467.600 26.200 ;
        RECT 465.800 22.200 466.600 25.600 ;
        RECT 472.600 22.200 474.200 26.200 ;
        RECT 480.600 22.200 482.200 26.200 ;
        RECT 486.000 26.000 490.000 26.200 ;
        RECT 486.000 22.200 486.800 26.000 ;
        RECT 489.200 22.200 490.000 26.000 ;
        RECT 490.800 22.200 491.600 26.200 ;
        RECT 492.400 22.200 493.200 26.200 ;
        RECT 494.000 26.000 498.000 26.200 ;
        RECT 494.000 22.200 494.800 26.000 ;
        RECT 497.200 22.200 498.000 26.000 ;
        RECT 498.800 22.200 499.600 26.200 ;
        RECT 500.400 26.000 504.400 26.200 ;
        RECT 500.400 22.200 501.200 26.000 ;
        RECT 503.600 22.200 504.400 26.000 ;
        RECT 508.200 22.200 509.800 26.200 ;
        RECT 513.200 22.200 514.000 29.700 ;
        RECT 514.800 30.300 515.600 30.400 ;
        RECT 516.400 30.300 518.000 30.400 ;
        RECT 514.800 29.800 518.000 30.300 ;
        RECT 514.800 29.700 517.200 29.800 ;
        RECT 514.800 29.600 515.600 29.700 ;
        RECT 516.400 29.600 517.200 29.700 ;
        RECT 519.600 29.600 520.400 30.400 ;
        RECT 522.800 29.600 523.600 31.200 ;
        RECT 518.000 27.600 518.800 29.200 ;
        RECT 514.800 24.800 515.600 26.400 ;
        RECT 519.800 26.200 520.400 29.600 ;
        RECT 521.000 28.800 521.800 29.600 ;
        RECT 521.200 28.400 521.800 28.800 ;
        RECT 526.200 28.400 526.800 31.800 ;
        RECT 527.600 29.600 528.400 31.200 ;
        RECT 533.200 30.400 533.800 31.800 ;
        RECT 537.400 31.200 538.000 31.800 ;
        RECT 534.600 30.600 538.000 31.200 ;
        RECT 534.600 30.400 535.400 30.600 ;
        RECT 532.400 29.800 533.800 30.400 ;
        RECT 538.800 30.300 539.600 30.400 ;
        RECT 540.400 30.300 541.200 31.200 ;
        RECT 536.800 29.800 537.600 30.000 ;
        RECT 532.400 29.600 534.200 29.800 ;
        RECT 533.200 29.200 534.200 29.600 ;
        RECT 521.200 28.300 522.000 28.400 ;
        RECT 526.000 28.300 526.800 28.400 ;
        RECT 521.200 27.700 526.800 28.300 ;
        RECT 521.200 27.600 522.000 27.700 ;
        RECT 526.000 27.600 526.800 27.700 ;
        RECT 529.200 27.600 530.800 28.400 ;
        RECT 532.000 27.600 532.800 28.400 ;
        RECT 519.400 22.200 521.000 26.200 ;
        RECT 524.400 24.800 525.200 26.400 ;
        RECT 526.200 24.200 526.800 27.600 ;
        RECT 532.200 27.200 532.800 27.600 ;
        RECT 530.800 26.800 531.600 27.000 ;
        RECT 526.000 22.200 526.800 24.200 ;
        RECT 529.200 26.200 531.600 26.800 ;
        RECT 532.200 26.400 533.000 27.200 ;
        RECT 529.200 22.200 530.000 26.200 ;
        RECT 533.600 25.800 534.200 29.200 ;
        RECT 535.000 29.200 537.600 29.800 ;
        RECT 538.800 29.700 541.200 30.300 ;
        RECT 538.800 29.600 539.600 29.700 ;
        RECT 540.400 29.600 541.200 29.700 ;
        RECT 535.000 28.600 535.600 29.200 ;
        RECT 534.800 27.800 535.600 28.600 ;
        RECT 542.000 28.400 542.600 31.800 ;
        RECT 545.400 30.400 546.000 31.800 ;
        RECT 551.600 31.600 552.400 33.200 ;
        RECT 553.200 32.300 554.000 39.800 ;
        RECT 554.800 32.300 555.600 32.400 ;
        RECT 553.200 31.700 555.600 32.300 ;
        RECT 549.200 30.400 550.000 30.800 ;
        RECT 545.200 29.800 547.600 30.400 ;
        RECT 549.200 29.800 550.800 30.400 ;
        RECT 545.200 29.600 546.000 29.800 ;
        RECT 538.000 28.300 539.600 28.400 ;
        RECT 540.400 28.300 541.200 28.400 ;
        RECT 538.000 28.200 541.200 28.300 ;
        RECT 536.200 27.700 541.200 28.200 ;
        RECT 536.200 27.600 539.600 27.700 ;
        RECT 540.400 27.600 541.200 27.700 ;
        RECT 542.000 28.300 542.800 28.400 ;
        RECT 542.000 27.700 545.900 28.300 ;
        RECT 542.000 27.600 542.800 27.700 ;
        RECT 536.200 27.200 536.800 27.600 ;
        RECT 534.800 26.600 536.800 27.200 ;
        RECT 537.400 26.800 538.200 27.000 ;
        RECT 534.800 26.400 536.400 26.600 ;
        RECT 537.400 26.200 539.600 26.800 ;
        RECT 533.600 22.200 535.200 25.800 ;
        RECT 538.800 22.200 539.600 26.200 ;
        RECT 542.000 24.200 542.600 27.600 ;
        RECT 545.300 26.400 545.900 27.700 ;
        RECT 543.600 24.800 544.400 26.400 ;
        RECT 545.200 25.600 546.000 26.400 ;
        RECT 547.000 26.200 547.600 29.800 ;
        RECT 550.000 29.600 550.800 29.800 ;
        RECT 548.400 27.600 549.200 29.200 ;
        RECT 553.200 26.200 554.000 31.700 ;
        RECT 554.800 31.600 555.600 31.700 ;
        RECT 554.800 26.800 555.600 28.400 ;
        RECT 545.400 24.800 546.200 25.600 ;
        RECT 542.000 22.200 542.800 24.200 ;
        RECT 546.800 22.200 547.600 26.200 ;
        RECT 552.200 25.600 554.000 26.200 ;
        RECT 552.200 22.200 553.000 25.600 ;
        RECT 556.400 22.200 557.200 39.800 ;
        RECT 560.400 33.600 561.200 34.400 ;
        RECT 560.400 32.400 561.000 33.600 ;
        RECT 561.800 32.400 562.600 39.800 ;
        RECT 559.600 31.800 561.000 32.400 ;
        RECT 561.600 31.800 562.600 32.400 ;
        RECT 566.000 32.400 566.800 39.800 ;
        RECT 570.400 38.400 572.000 39.800 ;
        RECT 569.200 37.600 572.000 38.400 ;
        RECT 567.600 32.400 568.400 32.600 ;
        RECT 570.400 32.400 572.000 37.600 ;
        RECT 566.000 31.800 568.400 32.400 ;
        RECT 570.000 31.800 572.000 32.400 ;
        RECT 574.200 32.400 575.000 32.600 ;
        RECT 575.600 32.400 576.400 39.800 ;
        RECT 574.200 31.800 576.400 32.400 ;
        RECT 579.800 32.400 580.600 39.800 ;
        RECT 581.200 33.600 582.000 34.400 ;
        RECT 581.400 32.400 582.000 33.600 ;
        RECT 579.800 31.800 580.800 32.400 ;
        RECT 581.400 31.800 582.800 32.400 ;
        RECT 559.600 31.600 560.400 31.800 ;
        RECT 561.600 28.400 562.200 31.800 ;
        RECT 570.000 30.400 570.600 31.800 ;
        RECT 574.200 31.200 574.800 31.800 ;
        RECT 571.400 30.600 574.800 31.200 ;
        RECT 571.400 30.400 572.200 30.600 ;
        RECT 562.800 28.800 563.600 30.400 ;
        RECT 569.200 29.800 570.600 30.400 ;
        RECT 573.600 29.800 574.400 30.000 ;
        RECT 569.200 29.600 571.000 29.800 ;
        RECT 570.000 29.200 571.000 29.600 ;
        RECT 559.600 27.600 562.200 28.400 ;
        RECT 564.400 28.200 565.200 28.400 ;
        RECT 563.600 27.600 565.200 28.200 ;
        RECT 566.000 27.600 567.600 28.400 ;
        RECT 568.800 27.600 569.600 28.400 ;
        RECT 558.000 24.800 558.800 26.400 ;
        RECT 559.800 26.200 560.400 27.600 ;
        RECT 563.600 27.200 564.400 27.600 ;
        RECT 569.000 27.200 569.600 27.600 ;
        RECT 567.600 26.800 568.400 27.000 ;
        RECT 561.400 26.200 565.000 26.600 ;
        RECT 566.000 26.200 568.400 26.800 ;
        RECT 569.000 26.400 569.800 27.200 ;
        RECT 559.600 22.200 560.400 26.200 ;
        RECT 561.200 26.000 565.200 26.200 ;
        RECT 561.200 22.200 562.000 26.000 ;
        RECT 564.400 22.200 565.200 26.000 ;
        RECT 566.000 22.200 566.800 26.200 ;
        RECT 570.400 25.800 571.000 29.200 ;
        RECT 571.800 29.200 574.400 29.800 ;
        RECT 571.800 28.600 572.400 29.200 ;
        RECT 578.800 28.800 579.600 30.400 ;
        RECT 571.600 27.800 572.400 28.600 ;
        RECT 580.200 28.400 580.800 31.800 ;
        RECT 582.000 31.600 582.800 31.800 ;
        RECT 574.800 28.200 576.400 28.400 ;
        RECT 573.000 27.600 576.400 28.200 ;
        RECT 577.200 28.200 578.000 28.400 ;
        RECT 577.200 27.600 578.800 28.200 ;
        RECT 580.200 27.600 582.800 28.400 ;
        RECT 573.000 27.200 573.600 27.600 ;
        RECT 578.000 27.200 578.800 27.600 ;
        RECT 571.600 26.600 573.600 27.200 ;
        RECT 574.200 26.800 575.000 27.000 ;
        RECT 571.600 26.400 573.200 26.600 ;
        RECT 574.200 26.200 576.400 26.800 ;
        RECT 577.400 26.200 581.000 26.600 ;
        RECT 582.000 26.200 582.600 27.600 ;
        RECT 570.400 22.200 572.000 25.800 ;
        RECT 575.600 22.200 576.400 26.200 ;
        RECT 577.200 26.000 581.200 26.200 ;
        RECT 577.200 22.200 578.000 26.000 ;
        RECT 580.400 22.200 581.200 26.000 ;
        RECT 582.000 22.200 582.800 26.200 ;
        RECT 1.200 15.600 2.000 17.200 ;
        RECT 2.800 2.200 3.600 19.800 ;
        RECT 5.600 14.200 6.400 19.800 ;
        RECT 10.800 15.800 11.600 19.800 ;
        RECT 12.400 16.000 13.200 19.800 ;
        RECT 15.600 16.000 16.400 19.800 ;
        RECT 12.400 15.800 16.400 16.000 ;
        RECT 17.200 15.800 18.000 19.800 ;
        RECT 21.600 16.200 23.200 19.800 ;
        RECT 11.000 14.400 11.600 15.800 ;
        RECT 12.600 15.400 16.200 15.800 ;
        RECT 17.200 15.200 19.600 15.800 ;
        RECT 18.800 15.000 19.600 15.200 ;
        RECT 20.200 14.800 21.000 15.600 ;
        RECT 14.800 14.400 15.600 14.800 ;
        RECT 20.200 14.400 20.800 14.800 ;
        RECT 4.600 13.800 6.400 14.200 ;
        RECT 4.600 13.600 6.200 13.800 ;
        RECT 10.800 13.600 13.400 14.400 ;
        RECT 14.800 13.800 16.400 14.400 ;
        RECT 15.600 13.600 16.400 13.800 ;
        RECT 17.200 13.600 18.800 14.400 ;
        RECT 20.000 13.600 20.800 14.400 ;
        RECT 4.600 10.400 5.200 13.600 ;
        RECT 12.800 12.400 13.400 13.600 ;
        RECT 6.800 11.600 8.400 12.400 ;
        RECT 12.400 11.600 13.400 12.400 ;
        RECT 14.000 11.600 14.800 13.200 ;
        RECT 21.600 12.800 22.200 16.200 ;
        RECT 26.800 15.800 27.600 19.800 ;
        RECT 22.800 15.400 24.400 15.600 ;
        RECT 22.800 14.800 24.800 15.400 ;
        RECT 25.400 15.200 27.600 15.800 ;
        RECT 28.400 15.800 29.200 19.800 ;
        RECT 32.800 16.200 34.400 19.800 ;
        RECT 28.400 15.200 30.800 15.800 ;
        RECT 25.400 15.000 26.200 15.200 ;
        RECT 30.000 15.000 30.800 15.200 ;
        RECT 24.200 14.400 24.800 14.800 ;
        RECT 31.400 14.800 32.200 15.600 ;
        RECT 31.400 14.400 32.000 14.800 ;
        RECT 22.800 13.400 23.600 14.200 ;
        RECT 24.200 13.800 27.600 14.400 ;
        RECT 26.000 13.600 27.600 13.800 ;
        RECT 28.400 13.600 30.000 14.400 ;
        RECT 31.200 13.600 32.000 14.400 ;
        RECT 21.200 12.400 22.200 12.800 ;
        RECT 20.400 12.200 22.200 12.400 ;
        RECT 23.000 12.800 23.600 13.400 ;
        RECT 32.800 12.800 33.400 16.200 ;
        RECT 38.000 15.800 38.800 19.800 ;
        RECT 34.000 15.400 35.600 15.600 ;
        RECT 34.000 14.800 36.000 15.400 ;
        RECT 36.600 15.200 38.800 15.800 ;
        RECT 36.600 15.000 37.400 15.200 ;
        RECT 39.600 15.000 40.400 19.800 ;
        RECT 44.000 18.400 44.800 19.800 ;
        RECT 42.800 17.800 44.800 18.400 ;
        RECT 48.400 17.800 49.200 19.800 ;
        RECT 52.600 18.400 53.800 19.800 ;
        RECT 52.400 17.800 53.800 18.400 ;
        RECT 42.800 17.000 43.600 17.800 ;
        RECT 48.400 17.200 49.000 17.800 ;
        RECT 44.400 16.400 45.200 17.200 ;
        RECT 46.200 16.600 49.000 17.200 ;
        RECT 52.400 17.000 53.200 17.800 ;
        RECT 46.200 16.400 47.000 16.600 ;
        RECT 35.400 14.400 36.000 14.800 ;
        RECT 34.000 13.400 34.800 14.200 ;
        RECT 35.400 13.800 38.800 14.400 ;
        RECT 37.200 13.600 38.800 13.800 ;
        RECT 40.400 14.200 42.000 14.400 ;
        RECT 44.600 14.200 45.200 16.400 ;
        RECT 54.200 15.400 55.000 15.600 ;
        RECT 57.200 15.400 58.000 19.800 ;
        RECT 54.200 14.800 58.000 15.400 ;
        RECT 58.800 15.000 59.600 19.800 ;
        RECT 63.200 18.400 64.000 19.800 ;
        RECT 62.000 17.800 64.000 18.400 ;
        RECT 67.600 17.800 68.400 19.800 ;
        RECT 71.800 18.400 73.000 19.800 ;
        RECT 71.600 17.800 73.000 18.400 ;
        RECT 62.000 17.000 62.800 17.800 ;
        RECT 67.600 17.200 68.200 17.800 ;
        RECT 63.600 16.400 64.400 17.200 ;
        RECT 65.400 16.600 68.200 17.200 ;
        RECT 71.600 17.000 72.400 17.800 ;
        RECT 65.400 16.400 66.200 16.600 ;
        RECT 50.200 14.200 51.000 14.400 ;
        RECT 40.400 13.600 51.400 14.200 ;
        RECT 43.400 13.400 44.200 13.600 ;
        RECT 23.000 12.200 25.600 12.800 ;
        RECT 32.400 12.400 33.400 12.800 ;
        RECT 20.400 11.600 21.800 12.200 ;
        RECT 24.800 12.000 25.600 12.200 ;
        RECT 31.600 12.200 33.400 12.400 ;
        RECT 34.200 12.800 34.800 13.400 ;
        RECT 34.200 12.200 36.800 12.800 ;
        RECT 31.600 11.600 33.000 12.200 ;
        RECT 36.000 12.000 36.800 12.200 ;
        RECT 41.800 12.400 42.600 12.600 ;
        RECT 44.400 12.400 45.200 12.600 ;
        RECT 50.800 12.400 51.400 13.600 ;
        RECT 52.400 12.800 53.200 13.000 ;
        RECT 41.800 11.800 46.800 12.400 ;
        RECT 46.000 11.600 46.800 11.800 ;
        RECT 50.800 11.600 51.600 12.400 ;
        RECT 52.400 12.200 56.200 12.800 ;
        RECT 55.400 12.000 56.200 12.200 ;
        RECT 4.400 9.600 5.200 10.400 ;
        RECT 9.200 9.600 10.000 11.200 ;
        RECT 10.800 10.200 11.600 10.400 ;
        RECT 12.800 10.200 13.400 11.600 ;
        RECT 21.200 10.200 21.800 11.600 ;
        RECT 22.600 11.400 23.400 11.600 ;
        RECT 22.600 10.800 26.000 11.400 ;
        RECT 25.400 10.200 26.000 10.800 ;
        RECT 32.400 10.200 33.000 11.600 ;
        RECT 33.800 11.400 34.600 11.600 ;
        RECT 33.800 10.800 37.200 11.400 ;
        RECT 36.600 10.200 37.200 10.800 ;
        RECT 39.600 11.000 45.200 11.200 ;
        RECT 39.600 10.800 45.400 11.000 ;
        RECT 39.600 10.600 49.400 10.800 ;
        RECT 10.800 9.600 12.200 10.200 ;
        RECT 12.800 9.600 13.800 10.200 ;
        RECT 4.600 7.000 5.200 9.600 ;
        RECT 6.000 7.600 6.800 9.200 ;
        RECT 11.600 8.400 12.200 9.600 ;
        RECT 11.600 7.600 12.400 8.400 ;
        RECT 4.600 6.400 8.200 7.000 ;
        RECT 4.600 6.200 5.200 6.400 ;
        RECT 4.400 2.200 5.200 6.200 ;
        RECT 7.600 2.200 8.400 6.400 ;
        RECT 13.000 2.200 13.800 9.600 ;
        RECT 17.200 9.600 19.600 10.200 ;
        RECT 21.200 9.600 23.200 10.200 ;
        RECT 17.200 2.200 18.000 9.600 ;
        RECT 18.800 9.400 19.600 9.600 ;
        RECT 21.600 8.400 23.200 9.600 ;
        RECT 25.400 9.600 27.600 10.200 ;
        RECT 25.400 9.400 26.200 9.600 ;
        RECT 21.600 7.600 24.400 8.400 ;
        RECT 21.600 2.200 23.200 7.600 ;
        RECT 26.800 2.200 27.600 9.600 ;
        RECT 28.400 9.600 30.800 10.200 ;
        RECT 32.400 9.600 34.400 10.200 ;
        RECT 28.400 2.200 29.200 9.600 ;
        RECT 30.000 9.400 30.800 9.600 ;
        RECT 32.800 8.400 34.400 9.600 ;
        RECT 36.600 9.600 38.800 10.200 ;
        RECT 36.600 9.400 37.400 9.600 ;
        RECT 32.800 7.600 35.600 8.400 ;
        RECT 32.800 2.200 34.400 7.600 ;
        RECT 38.000 2.200 38.800 9.600 ;
        RECT 39.600 2.200 40.400 10.600 ;
        RECT 44.600 10.200 49.400 10.600 ;
        RECT 42.800 9.000 48.200 9.600 ;
        RECT 42.800 8.800 43.600 9.000 ;
        RECT 47.400 8.800 48.200 9.000 ;
        RECT 48.800 9.000 49.400 10.200 ;
        RECT 50.800 10.400 51.400 11.600 ;
        RECT 53.800 11.400 54.600 11.600 ;
        RECT 57.200 11.400 58.000 14.800 ;
        RECT 59.600 14.200 61.200 14.400 ;
        RECT 63.800 14.200 64.400 16.400 ;
        RECT 73.400 15.400 74.200 15.600 ;
        RECT 76.400 15.400 77.200 19.800 ;
        RECT 73.400 14.800 77.200 15.400 ;
        RECT 78.000 15.000 78.800 19.800 ;
        RECT 82.400 18.400 83.200 19.800 ;
        RECT 81.200 17.800 83.200 18.400 ;
        RECT 86.800 17.800 87.600 19.800 ;
        RECT 91.000 18.400 92.200 19.800 ;
        RECT 90.800 17.800 92.200 18.400 ;
        RECT 81.200 17.000 82.000 17.800 ;
        RECT 86.800 17.200 87.400 17.800 ;
        RECT 82.800 16.400 83.600 17.200 ;
        RECT 84.600 16.600 87.400 17.200 ;
        RECT 90.800 17.000 91.600 17.800 ;
        RECT 84.600 16.400 85.400 16.600 ;
        RECT 69.400 14.200 70.200 14.400 ;
        RECT 59.600 13.600 70.600 14.200 ;
        RECT 62.600 13.400 63.400 13.600 ;
        RECT 61.000 12.400 61.800 12.600 ;
        RECT 63.600 12.400 64.400 12.600 ;
        RECT 70.000 12.400 70.600 13.600 ;
        RECT 71.600 12.800 72.400 13.000 ;
        RECT 61.000 11.800 66.000 12.400 ;
        RECT 65.200 11.600 66.000 11.800 ;
        RECT 70.000 11.600 70.800 12.400 ;
        RECT 71.600 12.200 75.400 12.800 ;
        RECT 74.600 12.000 75.400 12.200 ;
        RECT 53.800 10.800 58.000 11.400 ;
        RECT 50.800 9.800 53.200 10.400 ;
        RECT 50.200 9.000 51.000 9.200 ;
        RECT 48.800 8.400 51.000 9.000 ;
        RECT 52.600 8.800 53.200 9.800 ;
        RECT 52.600 8.000 54.000 8.800 ;
        RECT 46.200 7.400 47.000 7.600 ;
        RECT 49.000 7.400 49.800 7.600 ;
        RECT 42.800 6.200 43.600 7.000 ;
        RECT 46.200 6.800 49.800 7.400 ;
        RECT 48.400 6.200 49.000 6.800 ;
        RECT 52.400 6.200 53.200 7.000 ;
        RECT 42.800 5.600 44.800 6.200 ;
        RECT 44.000 2.200 44.800 5.600 ;
        RECT 48.400 2.200 49.200 6.200 ;
        RECT 52.600 2.200 53.800 6.200 ;
        RECT 57.200 2.200 58.000 10.800 ;
        RECT 58.800 11.000 64.400 11.200 ;
        RECT 58.800 10.800 64.600 11.000 ;
        RECT 58.800 10.600 68.600 10.800 ;
        RECT 58.800 2.200 59.600 10.600 ;
        RECT 63.800 10.200 68.600 10.600 ;
        RECT 62.000 9.000 67.400 9.600 ;
        RECT 62.000 8.800 62.800 9.000 ;
        RECT 66.600 8.800 67.400 9.000 ;
        RECT 68.000 9.000 68.600 10.200 ;
        RECT 70.000 10.400 70.600 11.600 ;
        RECT 73.000 11.400 73.800 11.600 ;
        RECT 76.400 11.400 77.200 14.800 ;
        RECT 78.800 14.200 80.400 14.400 ;
        RECT 83.000 14.200 83.600 16.400 ;
        RECT 92.600 15.400 93.400 15.600 ;
        RECT 95.600 15.400 96.400 19.800 ;
        RECT 92.600 14.800 96.400 15.400 ;
        RECT 97.200 15.000 98.000 19.800 ;
        RECT 101.600 18.400 102.400 19.800 ;
        RECT 100.400 17.800 102.400 18.400 ;
        RECT 106.000 17.800 106.800 19.800 ;
        RECT 110.200 18.400 111.400 19.800 ;
        RECT 110.000 17.800 111.400 18.400 ;
        RECT 100.400 17.000 101.200 17.800 ;
        RECT 106.000 17.200 106.600 17.800 ;
        RECT 102.000 16.400 102.800 17.200 ;
        RECT 103.800 16.600 106.600 17.200 ;
        RECT 110.000 17.000 110.800 17.800 ;
        RECT 103.800 16.400 104.600 16.600 ;
        RECT 88.600 14.200 89.400 14.400 ;
        RECT 78.800 13.600 89.800 14.200 ;
        RECT 81.800 13.400 82.600 13.600 ;
        RECT 80.200 12.400 81.000 12.600 ;
        RECT 82.800 12.400 83.600 12.600 ;
        RECT 89.200 12.400 89.800 13.600 ;
        RECT 90.800 12.800 91.600 13.000 ;
        RECT 80.200 11.800 85.200 12.400 ;
        RECT 84.400 11.600 85.200 11.800 ;
        RECT 89.200 11.600 90.000 12.400 ;
        RECT 90.800 12.200 94.600 12.800 ;
        RECT 93.800 12.000 94.600 12.200 ;
        RECT 73.000 10.800 77.200 11.400 ;
        RECT 70.000 9.800 72.400 10.400 ;
        RECT 69.400 9.000 70.200 9.200 ;
        RECT 68.000 8.400 70.200 9.000 ;
        RECT 71.800 8.800 72.400 9.800 ;
        RECT 71.800 8.000 73.200 8.800 ;
        RECT 65.400 7.400 66.200 7.600 ;
        RECT 68.200 7.400 69.000 7.600 ;
        RECT 62.000 6.200 62.800 7.000 ;
        RECT 65.400 6.800 69.000 7.400 ;
        RECT 67.600 6.200 68.200 6.800 ;
        RECT 71.600 6.200 72.400 7.000 ;
        RECT 62.000 5.600 64.000 6.200 ;
        RECT 63.200 2.200 64.000 5.600 ;
        RECT 67.600 2.200 68.400 6.200 ;
        RECT 71.800 2.200 73.000 6.200 ;
        RECT 76.400 2.200 77.200 10.800 ;
        RECT 78.000 11.000 83.600 11.200 ;
        RECT 78.000 10.800 83.800 11.000 ;
        RECT 78.000 10.600 87.800 10.800 ;
        RECT 78.000 2.200 78.800 10.600 ;
        RECT 83.000 10.200 87.800 10.600 ;
        RECT 81.200 9.000 86.600 9.600 ;
        RECT 81.200 8.800 82.000 9.000 ;
        RECT 85.800 8.800 86.600 9.000 ;
        RECT 87.200 9.000 87.800 10.200 ;
        RECT 89.200 10.400 89.800 11.600 ;
        RECT 92.200 11.400 93.000 11.600 ;
        RECT 95.600 11.400 96.400 14.800 ;
        RECT 98.000 14.200 99.600 14.400 ;
        RECT 102.200 14.200 102.800 16.400 ;
        RECT 111.800 15.400 112.600 15.600 ;
        RECT 114.800 15.400 115.600 19.800 ;
        RECT 111.800 14.800 115.600 15.400 ;
        RECT 116.400 15.000 117.200 19.800 ;
        RECT 120.800 18.400 121.600 19.800 ;
        RECT 119.600 17.800 121.600 18.400 ;
        RECT 125.200 17.800 126.000 19.800 ;
        RECT 129.400 18.400 130.600 19.800 ;
        RECT 129.200 17.800 130.600 18.400 ;
        RECT 119.600 17.000 120.400 17.800 ;
        RECT 125.200 17.200 125.800 17.800 ;
        RECT 121.200 16.400 122.000 17.200 ;
        RECT 123.000 16.600 125.800 17.200 ;
        RECT 129.200 17.000 130.000 17.800 ;
        RECT 123.000 16.400 123.800 16.600 ;
        RECT 107.800 14.200 108.600 14.400 ;
        RECT 98.000 13.600 109.000 14.200 ;
        RECT 101.000 13.400 101.800 13.600 ;
        RECT 99.400 12.400 100.200 12.600 ;
        RECT 102.000 12.400 102.800 12.600 ;
        RECT 108.400 12.400 109.000 13.600 ;
        RECT 110.000 12.800 110.800 13.000 ;
        RECT 99.400 11.800 104.400 12.400 ;
        RECT 103.600 11.600 104.400 11.800 ;
        RECT 108.400 11.600 109.200 12.400 ;
        RECT 110.000 12.200 113.800 12.800 ;
        RECT 113.000 12.000 113.800 12.200 ;
        RECT 92.200 10.800 96.400 11.400 ;
        RECT 89.200 9.800 91.600 10.400 ;
        RECT 88.600 9.000 89.400 9.200 ;
        RECT 87.200 8.400 89.400 9.000 ;
        RECT 91.000 8.800 91.600 9.800 ;
        RECT 91.000 8.000 92.400 8.800 ;
        RECT 84.600 7.400 85.400 7.600 ;
        RECT 87.400 7.400 88.200 7.600 ;
        RECT 81.200 6.200 82.000 7.000 ;
        RECT 84.600 6.800 88.200 7.400 ;
        RECT 86.800 6.200 87.400 6.800 ;
        RECT 90.800 6.200 91.600 7.000 ;
        RECT 81.200 5.600 83.200 6.200 ;
        RECT 82.400 2.200 83.200 5.600 ;
        RECT 86.800 2.200 87.600 6.200 ;
        RECT 91.000 2.200 92.200 6.200 ;
        RECT 95.600 2.200 96.400 10.800 ;
        RECT 97.200 11.000 102.800 11.200 ;
        RECT 97.200 10.800 103.000 11.000 ;
        RECT 97.200 10.600 107.000 10.800 ;
        RECT 97.200 2.200 98.000 10.600 ;
        RECT 102.200 10.200 107.000 10.600 ;
        RECT 100.400 9.000 105.800 9.600 ;
        RECT 100.400 8.800 101.200 9.000 ;
        RECT 105.000 8.800 105.800 9.000 ;
        RECT 106.400 9.000 107.000 10.200 ;
        RECT 108.400 10.400 109.000 11.600 ;
        RECT 111.400 11.400 112.200 11.600 ;
        RECT 114.800 11.400 115.600 14.800 ;
        RECT 117.200 14.200 118.800 14.400 ;
        RECT 121.400 14.200 122.000 16.400 ;
        RECT 131.000 15.400 131.800 15.600 ;
        RECT 134.000 15.400 134.800 19.800 ;
        RECT 131.000 14.800 134.800 15.400 ;
        RECT 140.400 15.800 141.200 19.800 ;
        RECT 144.800 16.200 146.400 19.800 ;
        RECT 140.400 15.200 142.600 15.800 ;
        RECT 143.600 15.400 145.200 15.600 ;
        RECT 141.800 15.000 142.600 15.200 ;
        RECT 127.000 14.200 127.800 14.400 ;
        RECT 117.200 13.600 128.200 14.200 ;
        RECT 120.200 13.400 121.000 13.600 ;
        RECT 118.600 12.400 119.400 12.600 ;
        RECT 118.600 11.800 123.600 12.400 ;
        RECT 122.800 11.600 123.600 11.800 ;
        RECT 111.400 10.800 115.600 11.400 ;
        RECT 108.400 9.800 110.800 10.400 ;
        RECT 107.800 9.000 108.600 9.200 ;
        RECT 106.400 8.400 108.600 9.000 ;
        RECT 110.200 8.800 110.800 9.800 ;
        RECT 110.200 8.000 111.600 8.800 ;
        RECT 103.800 7.400 104.600 7.600 ;
        RECT 106.600 7.400 107.400 7.600 ;
        RECT 100.400 6.200 101.200 7.000 ;
        RECT 103.800 6.800 107.400 7.400 ;
        RECT 106.000 6.200 106.600 6.800 ;
        RECT 110.000 6.200 110.800 7.000 ;
        RECT 100.400 5.600 102.400 6.200 ;
        RECT 101.600 2.200 102.400 5.600 ;
        RECT 106.000 2.200 106.800 6.200 ;
        RECT 110.200 2.200 111.400 6.200 ;
        RECT 114.800 2.200 115.600 10.800 ;
        RECT 116.400 11.000 122.000 11.200 ;
        RECT 116.400 10.800 122.200 11.000 ;
        RECT 116.400 10.600 126.200 10.800 ;
        RECT 116.400 2.200 117.200 10.600 ;
        RECT 121.400 10.200 126.200 10.600 ;
        RECT 119.600 9.000 125.000 9.600 ;
        RECT 119.600 8.800 120.400 9.000 ;
        RECT 124.200 8.800 125.000 9.000 ;
        RECT 125.600 9.000 126.200 10.200 ;
        RECT 127.600 10.400 128.200 13.600 ;
        RECT 129.200 12.800 130.000 13.000 ;
        RECT 129.200 12.200 133.000 12.800 ;
        RECT 132.200 12.000 133.000 12.200 ;
        RECT 130.600 11.400 131.400 11.600 ;
        RECT 134.000 11.400 134.800 14.800 ;
        RECT 143.200 14.800 145.200 15.400 ;
        RECT 143.200 14.400 143.800 14.800 ;
        RECT 140.400 13.800 143.800 14.400 ;
        RECT 140.400 13.600 142.000 13.800 ;
        RECT 144.400 13.400 145.200 14.200 ;
        RECT 144.400 12.800 145.000 13.400 ;
        RECT 142.400 12.200 145.000 12.800 ;
        RECT 145.800 12.800 146.400 16.200 ;
        RECT 150.000 15.800 150.800 19.800 ;
        RECT 151.600 16.000 152.400 19.800 ;
        RECT 154.800 16.000 155.600 19.800 ;
        RECT 151.600 15.800 155.600 16.000 ;
        RECT 156.400 15.800 157.200 19.800 ;
        RECT 147.000 14.800 147.800 15.600 ;
        RECT 148.400 15.200 150.800 15.800 ;
        RECT 151.800 15.400 155.400 15.800 ;
        RECT 148.400 15.000 149.200 15.200 ;
        RECT 147.200 14.400 147.800 14.800 ;
        RECT 152.400 14.400 153.200 14.800 ;
        RECT 156.400 14.400 157.000 15.800 ;
        RECT 147.200 13.600 148.000 14.400 ;
        RECT 149.200 13.600 150.800 14.400 ;
        RECT 151.600 13.800 153.200 14.400 ;
        RECT 151.600 13.600 152.400 13.800 ;
        RECT 154.600 13.600 157.200 14.400 ;
        RECT 145.800 12.400 146.800 12.800 ;
        RECT 145.800 12.300 147.600 12.400 ;
        RECT 153.200 12.300 154.000 13.200 ;
        RECT 145.800 12.200 154.000 12.300 ;
        RECT 142.400 12.000 143.200 12.200 ;
        RECT 146.200 11.700 154.000 12.200 ;
        RECT 146.200 11.600 147.600 11.700 ;
        RECT 153.200 11.600 154.000 11.700 ;
        RECT 144.600 11.400 145.400 11.600 ;
        RECT 130.600 10.800 134.800 11.400 ;
        RECT 127.600 9.800 130.000 10.400 ;
        RECT 127.000 9.000 127.800 9.200 ;
        RECT 125.600 8.400 127.800 9.000 ;
        RECT 129.400 8.800 130.000 9.800 ;
        RECT 129.400 8.000 130.800 8.800 ;
        RECT 123.000 7.400 123.800 7.600 ;
        RECT 125.800 7.400 126.600 7.600 ;
        RECT 119.600 6.200 120.400 7.000 ;
        RECT 123.000 6.800 126.600 7.400 ;
        RECT 125.200 6.200 125.800 6.800 ;
        RECT 129.200 6.200 130.000 7.000 ;
        RECT 119.600 5.600 121.600 6.200 ;
        RECT 120.800 2.200 121.600 5.600 ;
        RECT 125.200 2.200 126.000 6.200 ;
        RECT 129.400 2.200 130.600 6.200 ;
        RECT 134.000 2.200 134.800 10.800 ;
        RECT 142.000 10.800 145.400 11.400 ;
        RECT 142.000 10.200 142.600 10.800 ;
        RECT 146.200 10.200 146.800 11.600 ;
        RECT 154.600 10.200 155.200 13.600 ;
        RECT 156.400 10.300 157.200 10.400 ;
        RECT 158.000 10.300 158.800 19.800 ;
        RECT 159.600 15.600 160.400 17.200 ;
        RECT 161.200 15.600 162.000 17.200 ;
        RECT 156.400 10.200 158.800 10.300 ;
        RECT 140.400 9.600 142.600 10.200 ;
        RECT 140.400 2.200 141.200 9.600 ;
        RECT 141.800 9.400 142.600 9.600 ;
        RECT 144.800 9.600 146.800 10.200 ;
        RECT 148.400 9.600 150.800 10.200 ;
        RECT 144.800 2.200 146.400 9.600 ;
        RECT 148.400 9.400 149.200 9.600 ;
        RECT 150.000 2.200 150.800 9.600 ;
        RECT 154.200 9.600 155.200 10.200 ;
        RECT 155.800 9.700 158.800 10.200 ;
        RECT 155.800 9.600 157.200 9.700 ;
        RECT 154.200 2.200 155.000 9.600 ;
        RECT 155.800 8.400 156.400 9.600 ;
        RECT 155.600 7.600 156.400 8.400 ;
        RECT 158.000 2.200 158.800 9.700 ;
        RECT 162.800 12.300 163.600 19.800 ;
        RECT 166.000 17.800 166.800 19.800 ;
        RECT 164.400 16.300 165.200 16.400 ;
        RECT 166.000 16.300 166.600 17.800 ;
        RECT 164.400 15.700 166.700 16.300 ;
        RECT 164.400 15.600 165.200 15.700 ;
        RECT 166.000 14.400 166.600 15.700 ;
        RECT 167.600 15.600 168.400 17.200 ;
        RECT 169.400 16.400 170.200 17.200 ;
        RECT 169.200 15.600 170.000 16.400 ;
        RECT 170.800 15.600 171.600 19.800 ;
        RECT 166.000 14.300 166.800 14.400 ;
        RECT 169.300 14.300 169.900 15.600 ;
        RECT 166.000 13.700 169.900 14.300 ;
        RECT 166.000 13.600 166.800 13.700 ;
        RECT 164.400 12.300 165.200 12.400 ;
        RECT 162.800 11.700 165.200 12.300 ;
        RECT 162.800 2.200 163.600 11.700 ;
        RECT 164.400 10.800 165.200 11.700 ;
        RECT 166.000 10.200 166.600 13.600 ;
        RECT 169.200 12.200 170.000 12.400 ;
        RECT 171.000 12.200 171.600 15.600 ;
        RECT 175.600 15.200 176.400 19.800 ;
        RECT 178.800 16.400 179.600 19.800 ;
        RECT 178.800 15.800 179.800 16.400 ;
        RECT 175.600 14.600 178.200 15.200 ;
        RECT 172.400 12.800 173.200 14.400 ;
        RECT 175.800 12.400 176.600 13.200 ;
        RECT 174.000 12.200 174.800 12.400 ;
        RECT 169.200 11.600 171.600 12.200 ;
        RECT 173.200 11.600 174.800 12.200 ;
        RECT 175.600 11.600 176.600 12.400 ;
        RECT 177.600 13.000 178.200 14.600 ;
        RECT 179.200 14.400 179.800 15.800 ;
        RECT 182.000 15.800 182.800 19.800 ;
        RECT 186.400 18.400 188.000 19.800 ;
        RECT 186.400 17.600 189.200 18.400 ;
        RECT 186.400 16.200 188.000 17.600 ;
        RECT 182.000 15.200 184.600 15.800 ;
        RECT 183.800 15.000 184.600 15.200 ;
        RECT 185.200 14.800 186.800 15.600 ;
        RECT 178.800 14.300 179.800 14.400 ;
        RECT 182.000 14.300 183.600 14.400 ;
        RECT 178.800 14.200 183.600 14.300 ;
        RECT 187.400 14.200 188.000 16.200 ;
        RECT 191.600 15.800 192.400 19.800 ;
        RECT 193.200 16.000 194.000 19.800 ;
        RECT 196.400 16.000 197.200 19.800 ;
        RECT 193.200 15.800 197.200 16.000 ;
        RECT 198.000 15.800 198.800 19.800 ;
        RECT 199.600 16.000 200.400 19.800 ;
        RECT 202.800 16.000 203.600 19.800 ;
        RECT 199.600 15.800 203.600 16.000 ;
        RECT 204.400 15.800 205.200 19.800 ;
        RECT 206.000 15.800 206.800 19.800 ;
        RECT 207.600 16.000 208.400 19.800 ;
        RECT 210.800 16.000 211.600 19.800 ;
        RECT 214.000 17.800 214.800 19.800 ;
        RECT 207.600 15.800 211.600 16.000 ;
        RECT 188.600 14.800 189.400 15.600 ;
        RECT 190.000 15.200 192.400 15.800 ;
        RECT 193.400 15.400 197.000 15.800 ;
        RECT 190.000 15.000 190.800 15.200 ;
        RECT 178.800 14.000 184.200 14.200 ;
        RECT 178.800 13.700 186.400 14.000 ;
        RECT 178.800 13.600 179.800 13.700 ;
        RECT 182.000 13.600 186.400 13.700 ;
        RECT 177.600 12.200 178.600 13.000 ;
        RECT 169.400 10.200 170.000 11.600 ;
        RECT 173.200 11.200 174.000 11.600 ;
        RECT 177.600 10.200 178.200 12.200 ;
        RECT 179.200 10.200 179.800 13.600 ;
        RECT 183.600 13.400 186.400 13.600 ;
        RECT 185.600 13.200 186.400 13.400 ;
        RECT 187.000 13.600 188.000 14.200 ;
        RECT 188.800 14.400 189.400 14.800 ;
        RECT 194.000 14.400 194.800 14.800 ;
        RECT 198.000 14.400 198.600 15.800 ;
        RECT 199.800 15.400 203.400 15.800 ;
        RECT 200.400 14.400 201.200 14.800 ;
        RECT 204.400 14.400 205.000 15.800 ;
        RECT 206.200 14.400 206.800 15.800 ;
        RECT 207.800 15.400 211.400 15.800 ;
        RECT 212.400 15.600 213.200 17.200 ;
        RECT 210.000 14.400 210.800 14.800 ;
        RECT 214.200 14.400 214.800 17.800 ;
        RECT 188.800 13.600 189.600 14.400 ;
        RECT 190.800 13.600 192.400 14.400 ;
        RECT 193.200 13.800 194.800 14.400 ;
        RECT 193.200 13.600 194.000 13.800 ;
        RECT 196.200 13.600 198.800 14.400 ;
        RECT 199.600 13.800 201.200 14.400 ;
        RECT 199.600 13.600 200.400 13.800 ;
        RECT 202.600 13.600 205.200 14.400 ;
        RECT 206.000 13.600 208.600 14.400 ;
        RECT 210.000 14.300 211.600 14.400 ;
        RECT 214.000 14.300 214.800 14.400 ;
        RECT 210.000 13.800 214.800 14.300 ;
        RECT 210.800 13.700 214.800 13.800 ;
        RECT 210.800 13.600 211.600 13.700 ;
        RECT 214.000 13.600 214.800 13.700 ;
        RECT 187.000 12.400 187.600 13.600 ;
        RECT 184.200 12.200 185.000 12.400 ;
        RECT 184.200 11.600 185.800 12.200 ;
        RECT 186.800 11.600 187.600 12.400 ;
        RECT 194.800 11.600 195.600 13.200 ;
        RECT 196.200 12.300 196.800 13.600 ;
        RECT 201.200 12.300 202.000 13.200 ;
        RECT 196.200 11.700 202.000 12.300 ;
        RECT 185.000 11.400 185.800 11.600 ;
        RECT 187.000 10.200 187.600 11.600 ;
        RECT 196.200 10.200 196.800 11.700 ;
        RECT 201.200 11.600 202.000 11.700 ;
        RECT 198.000 10.200 198.800 10.400 ;
        RECT 202.600 10.200 203.200 13.600 ;
        RECT 208.000 12.300 208.600 13.600 ;
        RECT 204.500 11.700 208.600 12.300 ;
        RECT 204.500 10.400 205.100 11.700 ;
        RECT 204.400 10.200 205.200 10.400 ;
        RECT 165.000 9.400 166.800 10.200 ;
        RECT 165.000 2.200 165.800 9.400 ;
        RECT 169.200 2.200 170.000 10.200 ;
        RECT 170.800 9.600 174.800 10.200 ;
        RECT 170.800 2.200 171.600 9.600 ;
        RECT 174.000 2.200 174.800 9.600 ;
        RECT 175.600 9.600 178.200 10.200 ;
        RECT 175.600 2.200 176.400 9.600 ;
        RECT 178.800 9.200 179.800 10.200 ;
        RECT 182.000 9.600 184.600 10.200 ;
        RECT 178.800 2.200 179.600 9.200 ;
        RECT 182.000 2.200 182.800 9.600 ;
        RECT 183.800 9.400 184.600 9.600 ;
        RECT 186.400 2.200 188.000 10.200 ;
        RECT 190.000 9.600 192.400 10.200 ;
        RECT 190.000 9.400 190.800 9.600 ;
        RECT 191.600 2.200 192.400 9.600 ;
        RECT 195.800 9.600 196.800 10.200 ;
        RECT 197.400 9.600 198.800 10.200 ;
        RECT 202.200 9.600 203.200 10.200 ;
        RECT 203.800 9.600 205.200 10.200 ;
        RECT 206.000 10.200 206.800 10.400 ;
        RECT 208.000 10.200 208.600 11.700 ;
        RECT 209.200 11.600 210.000 13.200 ;
        RECT 214.200 10.200 214.800 13.600 ;
        RECT 215.600 12.300 216.400 12.400 ;
        RECT 217.200 12.300 218.000 19.800 ;
        RECT 221.000 18.400 221.800 19.800 ;
        RECT 220.400 17.600 221.800 18.400 ;
        RECT 218.800 15.600 219.600 17.200 ;
        RECT 221.000 16.400 221.800 17.600 ;
        RECT 227.800 16.400 228.600 19.800 ;
        RECT 221.000 15.800 222.800 16.400 ;
        RECT 215.600 11.700 218.000 12.300 ;
        RECT 215.600 10.800 216.400 11.700 ;
        RECT 217.200 10.300 218.000 11.700 ;
        RECT 220.400 10.300 221.200 10.400 ;
        RECT 206.000 9.600 207.400 10.200 ;
        RECT 208.000 9.600 209.000 10.200 ;
        RECT 195.800 2.200 196.600 9.600 ;
        RECT 197.400 8.400 198.000 9.600 ;
        RECT 197.200 7.600 198.000 8.400 ;
        RECT 202.200 6.400 203.000 9.600 ;
        RECT 203.800 8.400 204.400 9.600 ;
        RECT 203.600 7.600 204.400 8.400 ;
        RECT 206.800 8.400 207.400 9.600 ;
        RECT 206.800 7.600 207.600 8.400 ;
        RECT 201.200 5.600 203.000 6.400 ;
        RECT 202.200 2.200 203.000 5.600 ;
        RECT 208.200 2.200 209.000 9.600 ;
        RECT 214.000 9.400 215.800 10.200 ;
        RECT 215.000 2.200 215.800 9.400 ;
        RECT 217.200 9.700 221.200 10.300 ;
        RECT 217.200 2.200 218.000 9.700 ;
        RECT 220.400 8.800 221.200 9.700 ;
        RECT 222.000 2.200 222.800 15.800 ;
        RECT 226.800 15.800 228.600 16.400 ;
        RECT 223.600 13.600 224.400 15.200 ;
        RECT 225.200 13.600 226.000 15.200 ;
        RECT 223.600 12.300 224.400 12.400 ;
        RECT 225.300 12.300 225.900 13.600 ;
        RECT 223.600 11.700 225.900 12.300 ;
        RECT 223.600 11.600 224.400 11.700 ;
        RECT 226.800 2.200 227.600 15.800 ;
        RECT 230.000 14.300 230.800 19.800 ;
        RECT 231.600 15.600 232.400 17.200 ;
        RECT 233.200 15.800 234.000 19.800 ;
        RECT 237.600 16.200 239.200 19.800 ;
        RECT 233.200 15.200 235.400 15.800 ;
        RECT 236.400 15.400 238.000 15.600 ;
        RECT 234.600 15.000 235.400 15.200 ;
        RECT 236.000 14.800 238.000 15.400 ;
        RECT 236.000 14.400 236.600 14.800 ;
        RECT 231.600 14.300 232.400 14.400 ;
        RECT 230.000 13.700 232.400 14.300 ;
        RECT 228.400 10.300 229.200 10.400 ;
        RECT 230.000 10.300 230.800 13.700 ;
        RECT 231.600 13.600 232.400 13.700 ;
        RECT 233.200 13.800 236.600 14.400 ;
        RECT 233.200 13.600 234.800 13.800 ;
        RECT 237.200 13.400 238.000 14.200 ;
        RECT 237.200 12.800 237.800 13.400 ;
        RECT 235.200 12.200 237.800 12.800 ;
        RECT 238.600 12.800 239.200 16.200 ;
        RECT 242.800 15.800 243.600 19.800 ;
        RECT 245.000 18.400 245.800 19.800 ;
        RECT 245.000 17.600 246.800 18.400 ;
        RECT 245.000 16.400 245.800 17.600 ;
        RECT 251.800 16.400 252.600 19.800 ;
        RECT 245.000 15.800 246.800 16.400 ;
        RECT 239.800 14.800 240.600 15.600 ;
        RECT 241.200 15.200 243.600 15.800 ;
        RECT 241.200 15.000 242.000 15.200 ;
        RECT 240.000 14.400 240.600 14.800 ;
        RECT 240.000 13.600 240.800 14.400 ;
        RECT 242.000 13.600 243.600 14.400 ;
        RECT 238.600 12.400 239.600 12.800 ;
        RECT 238.600 12.200 240.400 12.400 ;
        RECT 235.200 12.000 236.000 12.200 ;
        RECT 239.000 11.600 240.400 12.200 ;
        RECT 237.400 11.400 238.200 11.600 ;
        RECT 228.400 9.700 230.800 10.300 ;
        RECT 234.800 10.800 238.200 11.400 ;
        RECT 234.800 10.200 235.400 10.800 ;
        RECT 239.000 10.200 239.600 11.600 ;
        RECT 228.400 8.800 229.200 9.700 ;
        RECT 230.000 2.200 230.800 9.700 ;
        RECT 233.200 9.600 235.400 10.200 ;
        RECT 233.200 2.200 234.000 9.600 ;
        RECT 234.600 9.400 235.400 9.600 ;
        RECT 237.600 9.600 239.600 10.200 ;
        RECT 241.200 9.600 243.600 10.200 ;
        RECT 237.600 6.400 239.200 9.600 ;
        RECT 241.200 9.400 242.000 9.600 ;
        RECT 237.600 5.600 240.400 6.400 ;
        RECT 237.600 2.200 239.200 5.600 ;
        RECT 242.800 2.200 243.600 9.600 ;
        RECT 244.400 8.800 245.200 10.400 ;
        RECT 246.000 2.200 246.800 15.800 ;
        RECT 250.800 15.800 252.600 16.400 ;
        RECT 254.000 16.000 254.800 19.800 ;
        RECT 257.200 16.000 258.000 19.800 ;
        RECT 254.000 15.800 258.000 16.000 ;
        RECT 258.800 15.800 259.600 19.800 ;
        RECT 263.000 16.400 263.800 19.800 ;
        RECT 262.000 15.800 263.800 16.400 ;
        RECT 265.200 15.800 266.000 19.800 ;
        RECT 269.600 16.200 271.200 19.800 ;
        RECT 247.600 13.600 248.400 15.200 ;
        RECT 249.200 13.600 250.000 15.200 ;
        RECT 247.600 12.300 248.400 12.400 ;
        RECT 250.800 12.300 251.600 15.800 ;
        RECT 254.200 15.400 257.800 15.800 ;
        RECT 254.800 14.400 255.600 14.800 ;
        RECT 258.800 14.400 259.400 15.800 ;
        RECT 254.000 13.800 255.600 14.400 ;
        RECT 254.000 13.600 254.800 13.800 ;
        RECT 257.000 13.600 259.600 14.400 ;
        RECT 260.400 13.600 261.200 15.200 ;
        RECT 247.600 11.700 251.600 12.300 ;
        RECT 247.600 11.600 248.400 11.700 ;
        RECT 250.800 2.200 251.600 11.700 ;
        RECT 255.600 11.600 256.400 13.200 ;
        RECT 252.400 8.800 253.200 10.400 ;
        RECT 257.000 10.200 257.600 13.600 ;
        RECT 258.800 10.300 259.600 10.400 ;
        RECT 262.000 10.300 262.800 15.800 ;
        RECT 265.200 15.200 267.600 15.800 ;
        RECT 266.800 15.000 267.600 15.200 ;
        RECT 268.200 14.800 269.000 15.600 ;
        RECT 268.200 14.400 268.800 14.800 ;
        RECT 265.200 13.600 266.800 14.400 ;
        RECT 268.000 13.600 268.800 14.400 ;
        RECT 269.600 12.800 270.200 16.200 ;
        RECT 274.800 15.800 275.600 19.800 ;
        RECT 276.400 16.000 277.200 19.800 ;
        RECT 279.600 16.000 280.400 19.800 ;
        RECT 276.400 15.800 280.400 16.000 ;
        RECT 281.200 15.800 282.000 19.800 ;
        RECT 282.800 15.800 283.600 19.800 ;
        RECT 287.200 18.400 288.800 19.800 ;
        RECT 287.200 17.600 290.000 18.400 ;
        RECT 287.200 16.200 288.800 17.600 ;
        RECT 270.800 15.400 272.400 15.600 ;
        RECT 270.800 14.800 272.800 15.400 ;
        RECT 273.400 15.200 275.600 15.800 ;
        RECT 276.600 15.400 280.200 15.800 ;
        RECT 273.400 15.000 274.200 15.200 ;
        RECT 272.200 14.400 272.800 14.800 ;
        RECT 277.200 14.400 278.000 14.800 ;
        RECT 281.200 14.400 281.800 15.800 ;
        RECT 282.800 15.200 285.200 15.800 ;
        RECT 284.400 15.000 285.200 15.200 ;
        RECT 285.800 14.800 286.600 15.600 ;
        RECT 285.800 14.400 286.400 14.800 ;
        RECT 270.800 13.400 271.600 14.200 ;
        RECT 272.200 13.800 275.600 14.400 ;
        RECT 274.000 13.600 275.600 13.800 ;
        RECT 276.400 13.800 278.000 14.400 ;
        RECT 276.400 13.600 277.200 13.800 ;
        RECT 279.400 13.600 282.000 14.400 ;
        RECT 282.800 13.600 284.400 14.400 ;
        RECT 285.600 13.600 286.400 14.400 ;
        RECT 287.200 14.200 287.800 16.200 ;
        RECT 292.400 15.800 293.200 19.800 ;
        RECT 301.400 16.400 302.200 19.800 ;
        RECT 288.400 14.800 290.000 15.600 ;
        RECT 290.600 15.200 293.200 15.800 ;
        RECT 300.400 15.800 302.200 16.400 ;
        RECT 303.600 15.800 304.400 19.800 ;
        RECT 305.200 16.000 306.000 19.800 ;
        RECT 308.400 16.000 309.200 19.800 ;
        RECT 305.200 15.800 309.200 16.000 ;
        RECT 290.600 15.000 291.400 15.200 ;
        RECT 291.600 14.300 293.200 14.400 ;
        RECT 297.200 14.300 298.000 14.400 ;
        RECT 291.600 14.200 298.000 14.300 ;
        RECT 287.200 13.600 288.200 14.200 ;
        RECT 291.000 14.000 298.000 14.200 ;
        RECT 269.200 12.400 270.200 12.800 ;
        RECT 268.400 12.200 270.200 12.400 ;
        RECT 271.000 12.800 271.600 13.400 ;
        RECT 271.000 12.200 273.600 12.800 ;
        RECT 268.400 11.600 269.800 12.200 ;
        RECT 272.800 12.000 273.600 12.200 ;
        RECT 278.000 11.600 278.800 13.200 ;
        RECT 258.800 10.200 262.800 10.300 ;
        RECT 256.600 9.600 257.600 10.200 ;
        RECT 258.200 9.700 262.800 10.200 ;
        RECT 258.200 9.600 259.600 9.700 ;
        RECT 256.600 8.400 257.400 9.600 ;
        RECT 258.200 8.400 258.800 9.600 ;
        RECT 255.600 7.600 257.400 8.400 ;
        RECT 258.000 7.600 258.800 8.400 ;
        RECT 256.600 2.200 257.400 7.600 ;
        RECT 262.000 2.200 262.800 9.700 ;
        RECT 263.600 8.800 264.400 10.400 ;
        RECT 269.200 10.200 269.800 11.600 ;
        RECT 270.600 11.400 271.400 11.600 ;
        RECT 270.600 10.800 274.000 11.400 ;
        RECT 273.400 10.200 274.000 10.800 ;
        RECT 279.400 10.200 280.000 13.600 ;
        RECT 287.600 12.400 288.200 13.600 ;
        RECT 288.800 13.700 298.000 14.000 ;
        RECT 288.800 13.600 293.200 13.700 ;
        RECT 297.200 13.600 298.000 13.700 ;
        RECT 298.800 13.600 299.600 15.200 ;
        RECT 288.800 13.400 291.600 13.600 ;
        RECT 288.800 13.200 289.600 13.400 ;
        RECT 287.600 11.600 288.400 12.400 ;
        RECT 290.200 12.200 291.000 12.400 ;
        RECT 289.400 11.600 291.000 12.200 ;
        RECT 300.400 12.300 301.200 15.800 ;
        RECT 303.800 14.400 304.400 15.800 ;
        RECT 305.400 15.400 309.000 15.800 ;
        RECT 310.000 15.600 310.800 17.200 ;
        RECT 307.600 14.400 308.400 14.800 ;
        RECT 303.600 13.600 306.200 14.400 ;
        RECT 307.600 13.800 309.200 14.400 ;
        RECT 308.400 13.600 309.200 13.800 ;
        RECT 305.600 12.400 306.200 13.600 ;
        RECT 300.400 11.700 304.300 12.300 ;
        RECT 281.200 10.200 282.000 10.400 ;
        RECT 287.600 10.200 288.200 11.600 ;
        RECT 289.400 11.400 290.200 11.600 ;
        RECT 265.200 9.600 267.600 10.200 ;
        RECT 269.200 9.600 271.200 10.200 ;
        RECT 265.200 2.200 266.000 9.600 ;
        RECT 266.800 9.400 267.600 9.600 ;
        RECT 269.600 8.400 271.200 9.600 ;
        RECT 273.400 9.600 275.600 10.200 ;
        RECT 273.400 9.400 274.200 9.600 ;
        RECT 269.600 7.600 272.400 8.400 ;
        RECT 269.600 2.200 271.200 7.600 ;
        RECT 274.800 2.200 275.600 9.600 ;
        RECT 279.000 9.600 280.000 10.200 ;
        RECT 280.600 9.600 282.000 10.200 ;
        RECT 282.800 9.600 285.200 10.200 ;
        RECT 279.000 2.200 279.800 9.600 ;
        RECT 280.600 8.400 281.200 9.600 ;
        RECT 280.400 7.600 281.200 8.400 ;
        RECT 282.800 2.200 283.600 9.600 ;
        RECT 284.400 9.400 285.200 9.600 ;
        RECT 287.200 2.200 288.800 10.200 ;
        RECT 290.600 9.600 293.200 10.200 ;
        RECT 290.600 9.400 291.400 9.600 ;
        RECT 292.400 2.200 293.200 9.600 ;
        RECT 300.400 2.200 301.200 11.700 ;
        RECT 303.700 10.400 304.300 11.700 ;
        RECT 305.200 11.600 306.200 12.400 ;
        RECT 306.800 11.600 307.600 13.200 ;
        RECT 302.000 8.800 302.800 10.400 ;
        RECT 303.600 10.200 304.400 10.400 ;
        RECT 305.600 10.200 306.200 11.600 ;
        RECT 311.600 10.300 312.400 19.800 ;
        RECT 313.800 18.400 314.600 19.800 ;
        RECT 313.800 17.600 315.600 18.400 ;
        RECT 313.800 16.400 314.600 17.600 ;
        RECT 321.800 16.400 322.600 19.000 ;
        RECT 326.000 17.000 326.800 19.000 ;
        RECT 313.800 15.800 315.600 16.400 ;
        RECT 321.800 16.000 323.600 16.400 ;
        RECT 313.200 10.300 314.000 10.400 ;
        RECT 303.600 9.600 305.000 10.200 ;
        RECT 305.600 9.600 306.600 10.200 ;
        RECT 304.400 8.400 305.000 9.600 ;
        RECT 304.400 7.600 305.200 8.400 ;
        RECT 305.800 2.200 306.600 9.600 ;
        RECT 311.600 9.700 314.000 10.300 ;
        RECT 311.600 2.200 312.400 9.700 ;
        RECT 313.200 8.800 314.000 9.700 ;
        RECT 314.800 2.200 315.600 15.800 ;
        RECT 321.000 15.600 323.600 16.000 ;
        RECT 321.000 15.400 322.600 15.600 ;
        RECT 316.400 13.600 317.200 15.200 ;
        RECT 321.000 15.000 321.800 15.400 ;
        RECT 321.000 14.400 321.600 15.000 ;
        RECT 326.200 14.800 326.800 17.000 ;
        RECT 327.600 15.800 328.400 19.800 ;
        RECT 332.000 16.200 333.600 19.800 ;
        RECT 327.600 15.200 329.800 15.800 ;
        RECT 330.800 15.400 332.400 15.600 ;
        RECT 329.000 15.000 329.800 15.200 ;
        RECT 319.600 13.600 321.600 14.400 ;
        RECT 322.600 14.200 326.800 14.800 ;
        RECT 330.400 14.800 332.400 15.400 ;
        RECT 330.400 14.400 331.000 14.800 ;
        RECT 322.600 13.800 323.600 14.200 ;
        RECT 319.600 10.800 320.400 12.400 ;
        RECT 321.000 9.800 321.600 13.600 ;
        RECT 322.200 13.000 323.600 13.800 ;
        RECT 327.600 13.800 331.000 14.400 ;
        RECT 327.600 13.600 329.200 13.800 ;
        RECT 331.600 13.400 332.400 14.200 ;
        RECT 323.000 11.000 323.600 13.000 ;
        RECT 324.400 11.600 325.200 13.200 ;
        RECT 326.000 11.600 326.800 13.200 ;
        RECT 331.600 12.800 332.200 13.400 ;
        RECT 329.600 12.200 332.200 12.800 ;
        RECT 333.000 12.800 333.600 16.200 ;
        RECT 337.200 15.800 338.000 19.800 ;
        RECT 334.200 14.800 335.000 15.600 ;
        RECT 335.600 15.200 338.000 15.800 ;
        RECT 335.600 15.000 336.400 15.200 ;
        RECT 338.800 15.000 339.600 19.800 ;
        RECT 343.200 18.400 344.000 19.800 ;
        RECT 342.000 17.800 344.000 18.400 ;
        RECT 347.600 17.800 348.400 19.800 ;
        RECT 351.800 18.400 353.000 19.800 ;
        RECT 351.600 17.800 353.000 18.400 ;
        RECT 342.000 17.000 342.800 17.800 ;
        RECT 347.600 17.200 348.200 17.800 ;
        RECT 343.600 16.400 344.400 17.200 ;
        RECT 345.400 16.600 348.200 17.200 ;
        RECT 351.600 17.000 352.400 17.800 ;
        RECT 345.400 16.400 346.200 16.600 ;
        RECT 334.400 14.400 335.000 14.800 ;
        RECT 334.400 13.600 335.200 14.400 ;
        RECT 336.400 13.600 338.000 14.400 ;
        RECT 339.600 14.200 341.200 14.400 ;
        RECT 343.800 14.200 344.400 16.400 ;
        RECT 353.400 15.400 354.200 15.600 ;
        RECT 356.400 15.400 357.200 19.800 ;
        RECT 353.400 14.800 357.200 15.400 ;
        RECT 358.000 15.000 358.800 19.800 ;
        RECT 362.400 18.400 363.200 19.800 ;
        RECT 361.200 17.800 363.200 18.400 ;
        RECT 366.800 17.800 367.600 19.800 ;
        RECT 371.000 18.400 372.200 19.800 ;
        RECT 370.800 17.800 372.200 18.400 ;
        RECT 361.200 17.000 362.000 17.800 ;
        RECT 366.800 17.200 367.400 17.800 ;
        RECT 362.800 16.400 363.600 17.200 ;
        RECT 364.600 16.600 367.400 17.200 ;
        RECT 370.800 17.000 371.600 17.800 ;
        RECT 364.600 16.400 365.400 16.600 ;
        RECT 349.400 14.200 350.200 14.400 ;
        RECT 339.600 13.600 350.600 14.200 ;
        RECT 342.600 13.400 343.400 13.600 ;
        RECT 333.000 12.400 334.000 12.800 ;
        RECT 341.000 12.400 341.800 12.600 ;
        RECT 343.600 12.400 344.400 12.600 ;
        RECT 350.000 12.400 350.600 13.600 ;
        RECT 351.600 12.800 352.400 13.000 ;
        RECT 333.000 12.300 334.800 12.400 ;
        RECT 337.200 12.300 338.000 12.400 ;
        RECT 333.000 12.200 338.000 12.300 ;
        RECT 329.600 12.000 330.400 12.200 ;
        RECT 333.400 11.700 338.000 12.200 ;
        RECT 341.000 11.800 346.000 12.400 ;
        RECT 333.400 11.600 334.800 11.700 ;
        RECT 337.200 11.600 338.000 11.700 ;
        RECT 345.200 11.600 346.000 11.800 ;
        RECT 350.000 11.600 350.800 12.400 ;
        RECT 351.600 12.200 355.400 12.800 ;
        RECT 354.600 12.000 355.400 12.200 ;
        RECT 331.800 11.400 332.600 11.600 ;
        RECT 323.000 10.400 326.800 11.000 ;
        RECT 321.000 9.200 322.600 9.800 ;
        RECT 321.800 2.200 322.600 9.200 ;
        RECT 326.200 7.000 326.800 10.400 ;
        RECT 329.200 10.800 332.600 11.400 ;
        RECT 329.200 10.200 329.800 10.800 ;
        RECT 333.400 10.200 334.000 11.600 ;
        RECT 338.800 11.000 344.400 11.200 ;
        RECT 338.800 10.800 344.600 11.000 ;
        RECT 338.800 10.600 348.600 10.800 ;
        RECT 326.000 3.000 326.800 7.000 ;
        RECT 327.600 9.600 329.800 10.200 ;
        RECT 327.600 2.200 328.400 9.600 ;
        RECT 329.000 9.400 329.800 9.600 ;
        RECT 332.000 9.600 334.000 10.200 ;
        RECT 335.600 9.600 338.000 10.200 ;
        RECT 332.000 2.200 333.600 9.600 ;
        RECT 335.600 9.400 336.400 9.600 ;
        RECT 337.200 2.200 338.000 9.600 ;
        RECT 338.800 2.200 339.600 10.600 ;
        RECT 343.800 10.200 348.600 10.600 ;
        RECT 342.000 9.000 347.400 9.600 ;
        RECT 342.000 8.800 342.800 9.000 ;
        RECT 346.600 8.800 347.400 9.000 ;
        RECT 348.000 9.000 348.600 10.200 ;
        RECT 350.000 10.400 350.600 11.600 ;
        RECT 353.000 11.400 353.800 11.600 ;
        RECT 356.400 11.400 357.200 14.800 ;
        RECT 358.800 14.200 360.400 14.400 ;
        RECT 363.000 14.200 363.600 16.400 ;
        RECT 372.600 15.400 373.400 15.600 ;
        RECT 375.600 15.400 376.400 19.800 ;
        RECT 372.600 14.800 376.400 15.400 ;
        RECT 377.200 15.000 378.000 19.800 ;
        RECT 381.600 18.400 382.400 19.800 ;
        RECT 380.400 17.800 382.400 18.400 ;
        RECT 386.000 17.800 386.800 19.800 ;
        RECT 390.200 18.400 391.400 19.800 ;
        RECT 390.000 17.800 391.400 18.400 ;
        RECT 380.400 17.000 381.200 17.800 ;
        RECT 386.000 17.200 386.600 17.800 ;
        RECT 382.000 16.400 382.800 17.200 ;
        RECT 383.800 16.600 386.600 17.200 ;
        RECT 390.000 17.000 390.800 17.800 ;
        RECT 383.800 16.400 384.600 16.600 ;
        RECT 368.600 14.200 369.400 14.400 ;
        RECT 358.800 13.600 369.800 14.200 ;
        RECT 361.800 13.400 362.600 13.600 ;
        RECT 360.200 12.400 361.000 12.600 ;
        RECT 362.800 12.400 363.600 12.600 ;
        RECT 369.200 12.400 369.800 13.600 ;
        RECT 370.800 12.800 371.600 13.000 ;
        RECT 360.200 11.800 365.200 12.400 ;
        RECT 364.400 11.600 365.200 11.800 ;
        RECT 369.200 11.600 370.000 12.400 ;
        RECT 370.800 12.200 374.600 12.800 ;
        RECT 373.800 12.000 374.600 12.200 ;
        RECT 353.000 10.800 357.200 11.400 ;
        RECT 350.000 9.800 352.400 10.400 ;
        RECT 349.400 9.000 350.200 9.200 ;
        RECT 348.000 8.400 350.200 9.000 ;
        RECT 351.800 8.800 352.400 9.800 ;
        RECT 351.800 8.000 353.200 8.800 ;
        RECT 345.400 7.400 346.200 7.600 ;
        RECT 348.200 7.400 349.000 7.600 ;
        RECT 342.000 6.200 342.800 7.000 ;
        RECT 345.400 6.800 349.000 7.400 ;
        RECT 347.600 6.200 348.200 6.800 ;
        RECT 351.600 6.200 352.400 7.000 ;
        RECT 342.000 5.600 344.000 6.200 ;
        RECT 343.200 2.200 344.000 5.600 ;
        RECT 347.600 2.200 348.400 6.200 ;
        RECT 351.800 2.200 353.000 6.200 ;
        RECT 356.400 2.200 357.200 10.800 ;
        RECT 358.000 11.000 363.600 11.200 ;
        RECT 358.000 10.800 363.800 11.000 ;
        RECT 358.000 10.600 367.800 10.800 ;
        RECT 358.000 2.200 358.800 10.600 ;
        RECT 363.000 10.200 367.800 10.600 ;
        RECT 361.200 9.000 366.600 9.600 ;
        RECT 361.200 8.800 362.000 9.000 ;
        RECT 365.800 8.800 366.600 9.000 ;
        RECT 367.200 9.000 367.800 10.200 ;
        RECT 369.200 10.400 369.800 11.600 ;
        RECT 372.200 11.400 373.000 11.600 ;
        RECT 375.600 11.400 376.400 14.800 ;
        RECT 378.000 14.200 379.600 14.400 ;
        RECT 382.200 14.200 382.800 16.400 ;
        RECT 391.800 15.400 392.600 15.600 ;
        RECT 394.800 15.400 395.600 19.800 ;
        RECT 391.800 14.800 395.600 15.400 ;
        RECT 385.200 14.200 386.000 14.400 ;
        RECT 387.800 14.200 388.600 14.400 ;
        RECT 378.000 13.600 389.000 14.200 ;
        RECT 381.000 13.400 381.800 13.600 ;
        RECT 379.400 12.400 380.200 12.600 ;
        RECT 382.000 12.400 382.800 12.600 ;
        RECT 379.400 11.800 384.400 12.400 ;
        RECT 383.600 11.600 384.400 11.800 ;
        RECT 372.200 10.800 376.400 11.400 ;
        RECT 369.200 9.800 371.600 10.400 ;
        RECT 368.600 9.000 369.400 9.200 ;
        RECT 367.200 8.400 369.400 9.000 ;
        RECT 371.000 8.800 371.600 9.800 ;
        RECT 371.000 8.000 372.400 8.800 ;
        RECT 364.600 7.400 365.400 7.600 ;
        RECT 367.400 7.400 368.200 7.600 ;
        RECT 361.200 6.200 362.000 7.000 ;
        RECT 364.600 6.800 368.200 7.400 ;
        RECT 366.800 6.200 367.400 6.800 ;
        RECT 370.800 6.200 371.600 7.000 ;
        RECT 361.200 5.600 363.200 6.200 ;
        RECT 362.400 2.200 363.200 5.600 ;
        RECT 366.800 2.200 367.600 6.200 ;
        RECT 371.000 2.200 372.200 6.200 ;
        RECT 375.600 2.200 376.400 10.800 ;
        RECT 377.200 11.000 382.800 11.200 ;
        RECT 377.200 10.800 383.000 11.000 ;
        RECT 377.200 10.600 387.000 10.800 ;
        RECT 377.200 2.200 378.000 10.600 ;
        RECT 382.200 10.200 387.000 10.600 ;
        RECT 380.400 9.000 385.800 9.600 ;
        RECT 380.400 8.800 381.200 9.000 ;
        RECT 385.000 8.800 385.800 9.000 ;
        RECT 386.400 9.000 387.000 10.200 ;
        RECT 388.400 10.400 389.000 13.600 ;
        RECT 390.000 12.800 390.800 13.000 ;
        RECT 390.000 12.200 393.800 12.800 ;
        RECT 393.000 12.000 393.800 12.200 ;
        RECT 391.400 11.400 392.200 11.600 ;
        RECT 394.800 11.400 395.600 14.800 ;
        RECT 396.400 15.200 397.200 19.800 ;
        RECT 399.600 16.400 400.400 19.800 ;
        RECT 399.600 15.800 400.600 16.400 ;
        RECT 396.400 14.600 399.000 15.200 ;
        RECT 396.600 12.400 397.400 13.200 ;
        RECT 396.400 11.600 397.400 12.400 ;
        RECT 398.400 13.000 399.000 14.600 ;
        RECT 400.000 14.400 400.600 15.800 ;
        RECT 402.800 15.800 403.600 19.800 ;
        RECT 407.200 18.400 408.800 19.800 ;
        RECT 407.200 17.600 410.000 18.400 ;
        RECT 407.200 16.200 408.800 17.600 ;
        RECT 402.800 15.200 405.200 15.800 ;
        RECT 404.400 15.000 405.200 15.200 ;
        RECT 405.800 14.800 406.600 15.600 ;
        RECT 405.800 14.400 406.400 14.800 ;
        RECT 399.600 14.300 400.600 14.400 ;
        RECT 401.200 14.300 402.000 14.400 ;
        RECT 399.600 13.700 402.000 14.300 ;
        RECT 399.600 13.600 400.600 13.700 ;
        RECT 401.200 13.600 402.000 13.700 ;
        RECT 402.800 13.600 404.400 14.400 ;
        RECT 405.600 13.600 406.400 14.400 ;
        RECT 407.200 14.200 407.800 16.200 ;
        RECT 412.400 15.800 413.200 19.800 ;
        RECT 408.400 14.800 410.000 15.600 ;
        RECT 410.600 15.200 413.200 15.800 ;
        RECT 414.000 15.600 414.800 17.200 ;
        RECT 410.600 15.000 411.400 15.200 ;
        RECT 411.600 14.200 413.200 14.400 ;
        RECT 407.200 13.600 408.200 14.200 ;
        RECT 411.000 14.000 413.200 14.200 ;
        RECT 398.400 12.200 399.400 13.000 ;
        RECT 391.400 10.800 395.600 11.400 ;
        RECT 388.400 9.800 390.800 10.400 ;
        RECT 387.800 9.000 388.600 9.200 ;
        RECT 386.400 8.400 388.600 9.000 ;
        RECT 390.200 8.800 390.800 9.800 ;
        RECT 390.200 8.000 391.600 8.800 ;
        RECT 383.800 7.400 384.600 7.600 ;
        RECT 386.600 7.400 387.400 7.600 ;
        RECT 380.400 6.200 381.200 7.000 ;
        RECT 383.800 6.800 387.400 7.400 ;
        RECT 386.000 6.200 386.600 6.800 ;
        RECT 390.000 6.200 390.800 7.000 ;
        RECT 380.400 5.600 382.400 6.200 ;
        RECT 381.600 2.200 382.400 5.600 ;
        RECT 386.000 2.200 386.800 6.200 ;
        RECT 390.200 2.200 391.400 6.200 ;
        RECT 394.800 2.200 395.600 10.800 ;
        RECT 398.400 10.200 399.000 12.200 ;
        RECT 400.000 10.200 400.600 13.600 ;
        RECT 407.600 12.400 408.200 13.600 ;
        RECT 408.800 13.600 413.200 14.000 ;
        RECT 408.800 13.400 411.600 13.600 ;
        RECT 408.800 13.200 409.600 13.400 ;
        RECT 407.600 11.600 408.400 12.400 ;
        RECT 410.200 12.200 411.000 12.400 ;
        RECT 409.400 11.600 411.000 12.200 ;
        RECT 407.600 10.200 408.200 11.600 ;
        RECT 409.400 11.400 410.200 11.600 ;
        RECT 396.400 9.600 399.000 10.200 ;
        RECT 396.400 2.200 397.200 9.600 ;
        RECT 399.600 9.200 400.600 10.200 ;
        RECT 402.800 9.600 405.200 10.200 ;
        RECT 399.600 2.200 400.400 9.200 ;
        RECT 402.800 2.200 403.600 9.600 ;
        RECT 404.400 9.400 405.200 9.600 ;
        RECT 407.200 2.200 408.800 10.200 ;
        RECT 410.600 9.600 413.200 10.200 ;
        RECT 410.600 9.400 411.400 9.600 ;
        RECT 412.400 2.200 413.200 9.600 ;
        RECT 415.600 2.200 416.400 19.800 ;
        RECT 417.200 16.000 418.000 19.800 ;
        RECT 420.400 16.000 421.200 19.800 ;
        RECT 417.200 15.800 421.200 16.000 ;
        RECT 422.000 15.800 422.800 19.800 ;
        RECT 423.600 15.800 424.400 19.800 ;
        RECT 425.200 16.000 426.000 19.800 ;
        RECT 428.400 16.000 429.200 19.800 ;
        RECT 432.600 16.400 433.400 19.800 ;
        RECT 425.200 15.800 429.200 16.000 ;
        RECT 431.600 15.800 433.400 16.400 ;
        RECT 417.400 15.400 421.000 15.800 ;
        RECT 418.000 14.400 418.800 14.800 ;
        RECT 422.000 14.400 422.600 15.800 ;
        RECT 423.800 14.400 424.400 15.800 ;
        RECT 425.400 15.400 429.000 15.800 ;
        RECT 427.600 14.400 428.400 14.800 ;
        RECT 417.200 13.800 418.800 14.400 ;
        RECT 417.200 13.600 418.000 13.800 ;
        RECT 420.200 13.600 422.800 14.400 ;
        RECT 423.600 13.600 426.200 14.400 ;
        RECT 427.600 13.800 429.200 14.400 ;
        RECT 428.400 13.600 429.200 13.800 ;
        RECT 430.000 13.600 430.800 15.200 ;
        RECT 418.800 11.600 419.600 13.200 ;
        RECT 420.200 12.300 420.800 13.600 ;
        RECT 420.200 11.700 424.300 12.300 ;
        RECT 420.200 10.200 420.800 11.700 ;
        RECT 423.700 10.400 424.300 11.700 ;
        RECT 422.000 10.200 422.800 10.400 ;
        RECT 419.800 9.600 420.800 10.200 ;
        RECT 421.400 9.600 422.800 10.200 ;
        RECT 423.600 10.200 424.400 10.400 ;
        RECT 425.600 10.200 426.200 13.600 ;
        RECT 426.800 11.600 427.600 13.200 ;
        RECT 423.600 9.600 425.000 10.200 ;
        RECT 425.600 9.600 426.600 10.200 ;
        RECT 419.800 2.200 420.600 9.600 ;
        RECT 421.400 8.400 422.000 9.600 ;
        RECT 421.200 7.600 422.000 8.400 ;
        RECT 424.400 8.400 425.000 9.600 ;
        RECT 424.400 7.600 425.200 8.400 ;
        RECT 425.800 2.200 426.600 9.600 ;
        RECT 430.000 8.300 430.800 8.400 ;
        RECT 431.600 8.300 432.400 15.800 ;
        RECT 434.800 15.200 435.600 19.800 ;
        RECT 438.000 16.400 438.800 19.800 ;
        RECT 438.000 15.800 439.000 16.400 ;
        RECT 434.800 14.600 437.400 15.200 ;
        RECT 435.000 12.400 435.800 13.200 ;
        RECT 434.800 11.600 435.800 12.400 ;
        RECT 436.800 13.000 437.400 14.600 ;
        RECT 438.400 14.400 439.000 15.800 ;
        RECT 441.200 15.600 442.000 17.200 ;
        RECT 438.000 13.600 439.000 14.400 ;
        RECT 436.800 12.200 437.800 13.000 ;
        RECT 433.200 8.800 434.000 10.400 ;
        RECT 436.800 10.200 437.400 12.200 ;
        RECT 438.400 10.200 439.000 13.600 ;
        RECT 434.800 9.600 437.400 10.200 ;
        RECT 430.000 7.700 432.400 8.300 ;
        RECT 430.000 7.600 430.800 7.700 ;
        RECT 431.600 2.200 432.400 7.700 ;
        RECT 434.800 2.200 435.600 9.600 ;
        RECT 438.000 9.200 439.000 10.200 ;
        RECT 442.800 14.300 443.600 19.800 ;
        RECT 451.800 18.400 452.600 19.800 ;
        RECT 454.600 18.400 455.400 19.800 ;
        RECT 451.800 17.600 453.200 18.400 ;
        RECT 454.600 17.600 456.400 18.400 ;
        RECT 460.400 17.600 461.200 19.800 ;
        RECT 451.800 16.400 452.600 17.600 ;
        RECT 450.800 15.800 452.600 16.400 ;
        RECT 454.600 16.400 455.400 17.600 ;
        RECT 454.600 15.800 456.400 16.400 ;
        RECT 446.000 14.300 446.800 14.400 ;
        RECT 442.800 13.700 446.800 14.300 ;
        RECT 438.000 2.200 438.800 9.200 ;
        RECT 442.800 2.200 443.600 13.700 ;
        RECT 446.000 13.600 446.800 13.700 ;
        RECT 447.600 14.300 448.400 14.400 ;
        RECT 449.200 14.300 450.000 15.200 ;
        RECT 447.600 13.700 450.000 14.300 ;
        RECT 447.600 13.600 448.400 13.700 ;
        RECT 449.200 13.600 450.000 13.700 ;
        RECT 450.800 2.200 451.600 15.800 ;
        RECT 452.400 10.300 453.200 10.400 ;
        RECT 454.000 10.300 454.800 10.400 ;
        RECT 452.400 9.700 454.800 10.300 ;
        RECT 452.400 8.800 453.200 9.700 ;
        RECT 454.000 8.800 454.800 9.700 ;
        RECT 455.600 2.200 456.400 15.800 ;
        RECT 457.200 13.600 458.000 15.200 ;
        RECT 460.400 14.400 461.000 17.600 ;
        RECT 462.000 15.600 462.800 17.200 ;
        RECT 463.600 16.000 464.400 19.800 ;
        RECT 466.800 16.000 467.600 19.800 ;
        RECT 463.600 15.800 467.600 16.000 ;
        RECT 463.800 15.400 467.400 15.800 ;
        RECT 468.400 15.600 469.200 19.800 ;
        RECT 470.000 15.800 470.800 19.800 ;
        RECT 474.400 16.200 476.000 19.800 ;
        RECT 464.400 14.400 465.200 14.800 ;
        RECT 468.400 14.400 469.000 15.600 ;
        RECT 470.000 15.200 472.200 15.800 ;
        RECT 473.200 15.400 474.800 15.600 ;
        RECT 471.400 15.000 472.200 15.200 ;
        RECT 472.800 14.800 474.800 15.400 ;
        RECT 472.800 14.400 473.400 14.800 ;
        RECT 460.400 13.600 461.200 14.400 ;
        RECT 463.600 13.800 465.200 14.400 ;
        RECT 463.600 13.600 464.400 13.800 ;
        RECT 466.600 13.600 469.200 14.400 ;
        RECT 470.000 13.800 473.400 14.400 ;
        RECT 470.000 13.600 471.600 13.800 ;
        RECT 457.300 12.300 457.900 13.600 ;
        RECT 458.800 12.300 459.600 12.400 ;
        RECT 457.300 11.700 459.600 12.300 ;
        RECT 458.800 10.800 459.600 11.700 ;
        RECT 460.400 10.200 461.000 13.600 ;
        RECT 465.200 11.600 466.000 13.200 ;
        RECT 466.600 10.200 467.200 13.600 ;
        RECT 474.000 13.400 474.800 14.200 ;
        RECT 474.000 12.800 474.600 13.400 ;
        RECT 472.000 12.200 474.600 12.800 ;
        RECT 475.400 12.800 476.000 16.200 ;
        RECT 479.600 15.800 480.400 19.800 ;
        RECT 481.200 16.000 482.000 19.800 ;
        RECT 484.400 16.000 485.200 19.800 ;
        RECT 481.200 15.800 485.200 16.000 ;
        RECT 486.000 15.800 486.800 19.800 ;
        RECT 487.600 15.800 488.400 19.800 ;
        RECT 489.200 16.000 490.000 19.800 ;
        RECT 492.400 16.000 493.200 19.800 ;
        RECT 489.200 15.800 493.200 16.000 ;
        RECT 494.000 16.000 494.800 19.800 ;
        RECT 497.200 16.000 498.000 19.800 ;
        RECT 494.000 15.800 498.000 16.000 ;
        RECT 498.800 15.800 499.600 19.800 ;
        RECT 502.000 17.800 502.800 19.800 ;
        RECT 476.600 14.800 477.400 15.600 ;
        RECT 478.000 15.200 480.400 15.800 ;
        RECT 481.400 15.400 485.000 15.800 ;
        RECT 478.000 15.000 478.800 15.200 ;
        RECT 476.800 14.400 477.400 14.800 ;
        RECT 482.000 14.400 482.800 14.800 ;
        RECT 486.000 14.400 486.600 15.800 ;
        RECT 487.800 14.400 488.400 15.800 ;
        RECT 489.400 15.400 493.000 15.800 ;
        RECT 494.200 15.400 497.800 15.800 ;
        RECT 491.600 14.400 492.400 14.800 ;
        RECT 494.800 14.400 495.600 14.800 ;
        RECT 498.800 14.400 499.400 15.800 ;
        RECT 500.400 15.600 501.200 17.200 ;
        RECT 502.200 15.600 502.800 17.800 ;
        RECT 505.200 15.800 506.000 19.800 ;
        RECT 508.400 17.800 509.200 19.800 ;
        RECT 502.200 15.000 504.600 15.600 ;
        RECT 476.800 13.600 477.600 14.400 ;
        RECT 478.800 13.600 480.400 14.400 ;
        RECT 481.200 13.800 482.800 14.400 ;
        RECT 481.200 13.600 482.000 13.800 ;
        RECT 484.200 13.600 486.800 14.400 ;
        RECT 487.600 13.600 490.200 14.400 ;
        RECT 491.600 13.800 493.200 14.400 ;
        RECT 492.400 13.600 493.200 13.800 ;
        RECT 494.000 13.800 495.600 14.400 ;
        RECT 494.000 13.600 494.800 13.800 ;
        RECT 497.000 13.600 499.600 14.400 ;
        RECT 502.000 13.600 503.000 14.400 ;
        RECT 475.400 12.400 476.400 12.800 ;
        RECT 479.700 12.400 480.300 13.600 ;
        RECT 475.400 12.200 477.200 12.400 ;
        RECT 472.000 12.000 472.800 12.200 ;
        RECT 475.800 11.600 477.200 12.200 ;
        RECT 479.600 12.300 480.400 12.400 ;
        RECT 482.800 12.300 483.600 13.200 ;
        RECT 479.600 11.700 483.600 12.300 ;
        RECT 479.600 11.600 480.400 11.700 ;
        RECT 482.800 11.600 483.600 11.700 ;
        RECT 484.200 12.300 484.800 13.600 ;
        RECT 484.200 11.700 488.300 12.300 ;
        RECT 474.200 11.400 475.000 11.600 ;
        RECT 471.600 10.800 475.000 11.400 ;
        RECT 468.400 10.200 469.200 10.400 ;
        RECT 471.600 10.200 472.200 10.800 ;
        RECT 475.800 10.400 476.400 11.600 ;
        RECT 475.800 10.200 477.200 10.400 ;
        RECT 484.200 10.200 484.800 11.700 ;
        RECT 487.700 10.400 488.300 11.700 ;
        RECT 486.000 10.200 486.800 10.400 ;
        RECT 459.400 9.400 461.200 10.200 ;
        RECT 466.200 9.600 467.200 10.200 ;
        RECT 467.800 9.600 469.200 10.200 ;
        RECT 470.000 9.600 472.200 10.200 ;
        RECT 459.400 2.200 460.200 9.400 ;
        RECT 466.200 2.200 467.000 9.600 ;
        RECT 467.800 8.400 468.400 9.600 ;
        RECT 467.600 7.600 468.400 8.400 ;
        RECT 470.000 2.200 470.800 9.600 ;
        RECT 471.400 9.400 472.200 9.600 ;
        RECT 474.400 9.600 477.200 10.200 ;
        RECT 478.000 9.600 480.400 10.200 ;
        RECT 474.400 2.200 476.000 9.600 ;
        RECT 478.000 9.400 478.800 9.600 ;
        RECT 479.600 2.200 480.400 9.600 ;
        RECT 483.800 9.600 484.800 10.200 ;
        RECT 485.400 9.600 486.800 10.200 ;
        RECT 487.600 10.200 488.400 10.400 ;
        RECT 489.600 10.200 490.200 13.600 ;
        RECT 490.800 11.600 491.600 13.200 ;
        RECT 495.600 11.600 496.400 13.200 ;
        RECT 497.000 10.400 497.600 13.600 ;
        RECT 502.400 12.800 503.200 13.600 ;
        RECT 504.000 12.000 504.600 15.000 ;
        RECT 505.400 12.400 506.000 15.800 ;
        RECT 506.800 15.600 507.600 17.200 ;
        RECT 508.600 14.400 509.200 17.800 ;
        RECT 510.000 16.300 510.800 16.400 ;
        RECT 511.600 16.300 512.400 17.200 ;
        RECT 510.000 15.700 512.400 16.300 ;
        RECT 510.000 15.600 510.800 15.700 ;
        RECT 511.600 15.600 512.400 15.700 ;
        RECT 508.400 14.300 509.200 14.400 ;
        RECT 511.600 14.300 512.400 14.400 ;
        RECT 508.400 13.700 512.400 14.300 ;
        RECT 508.400 13.600 509.200 13.700 ;
        RECT 511.600 13.600 512.400 13.700 ;
        RECT 503.800 11.400 504.600 12.000 ;
        RECT 505.200 11.600 506.000 12.400 ;
        RECT 500.400 11.200 504.600 11.400 ;
        RECT 500.400 10.800 504.400 11.200 ;
        RECT 487.600 9.600 489.000 10.200 ;
        RECT 489.600 9.600 490.600 10.200 ;
        RECT 495.600 9.600 497.600 10.400 ;
        RECT 498.800 10.200 499.600 10.400 ;
        RECT 498.200 9.600 499.600 10.200 ;
        RECT 483.800 2.200 484.600 9.600 ;
        RECT 485.400 8.400 486.000 9.600 ;
        RECT 485.200 7.600 486.000 8.400 ;
        RECT 488.400 8.400 489.000 9.600 ;
        RECT 488.400 7.600 489.200 8.400 ;
        RECT 489.800 2.200 490.600 9.600 ;
        RECT 496.600 2.200 497.400 9.600 ;
        RECT 498.200 8.400 498.800 9.600 ;
        RECT 498.000 7.600 498.800 8.400 ;
        RECT 500.400 2.200 501.200 10.800 ;
        RECT 505.400 10.200 506.000 11.600 ;
        RECT 508.600 10.200 509.200 13.600 ;
        RECT 510.000 10.800 510.800 12.400 ;
        RECT 504.600 9.600 506.000 10.200 ;
        RECT 504.600 2.200 505.400 9.600 ;
        RECT 508.400 9.400 510.200 10.200 ;
        RECT 509.400 2.200 510.200 9.400 ;
        RECT 513.200 2.200 514.000 19.800 ;
        RECT 516.400 16.400 517.200 19.800 ;
        RECT 516.200 15.800 517.200 16.400 ;
        RECT 516.200 14.400 516.800 15.800 ;
        RECT 519.600 15.200 520.400 19.800 ;
        RECT 521.200 15.600 522.000 17.200 ;
        RECT 517.800 14.600 520.400 15.200 ;
        RECT 516.200 13.600 517.200 14.400 ;
        RECT 516.200 10.200 516.800 13.600 ;
        RECT 517.800 13.000 518.400 14.600 ;
        RECT 517.400 12.200 518.400 13.000 ;
        RECT 517.800 10.200 518.400 12.200 ;
        RECT 519.400 12.400 520.200 13.200 ;
        RECT 519.400 11.600 520.400 12.400 ;
        RECT 522.800 12.300 523.600 19.800 ;
        RECT 524.400 15.800 525.200 19.800 ;
        RECT 526.000 16.000 526.800 19.800 ;
        RECT 529.200 16.000 530.000 19.800 ;
        RECT 526.000 15.800 530.000 16.000 ;
        RECT 532.400 17.800 533.200 19.800 ;
        RECT 537.200 17.800 538.000 19.800 ;
        RECT 524.600 14.400 525.200 15.800 ;
        RECT 526.200 15.400 529.800 15.800 ;
        RECT 528.400 14.400 529.200 14.800 ;
        RECT 532.400 14.400 533.000 17.800 ;
        RECT 534.000 15.600 534.800 17.200 ;
        RECT 535.600 15.600 536.400 17.200 ;
        RECT 534.100 14.400 534.700 15.600 ;
        RECT 537.400 14.400 538.000 17.800 ;
        RECT 524.400 13.600 527.000 14.400 ;
        RECT 528.400 13.800 530.000 14.400 ;
        RECT 529.200 13.600 530.000 13.800 ;
        RECT 532.400 13.600 533.200 14.400 ;
        RECT 534.000 14.300 534.800 14.400 ;
        RECT 537.200 14.300 538.000 14.400 ;
        RECT 534.000 13.700 538.000 14.300 ;
        RECT 534.000 13.600 534.800 13.700 ;
        RECT 537.200 13.600 538.000 13.700 ;
        RECT 540.400 13.600 541.200 15.200 ;
        RECT 524.400 12.300 525.200 12.400 ;
        RECT 522.800 11.700 525.200 12.300 ;
        RECT 522.800 10.300 523.600 11.700 ;
        RECT 524.400 11.600 525.200 11.700 ;
        RECT 524.400 10.300 525.200 10.400 ;
        RECT 522.800 10.200 525.200 10.300 ;
        RECT 526.400 10.200 527.000 13.600 ;
        RECT 527.600 12.300 528.400 13.200 ;
        RECT 530.800 12.300 531.600 12.400 ;
        RECT 527.600 11.700 531.600 12.300 ;
        RECT 527.600 11.600 528.400 11.700 ;
        RECT 530.800 10.800 531.600 11.700 ;
        RECT 532.400 12.300 533.000 13.600 ;
        RECT 535.600 12.300 536.400 12.400 ;
        RECT 532.400 11.700 536.400 12.300 ;
        RECT 532.400 10.200 533.000 11.700 ;
        RECT 535.600 11.600 536.400 11.700 ;
        RECT 537.400 10.200 538.000 13.600 ;
        RECT 538.800 10.800 539.600 12.400 ;
        RECT 516.200 9.200 517.200 10.200 ;
        RECT 517.800 9.600 520.400 10.200 ;
        RECT 516.400 2.200 517.200 9.200 ;
        RECT 519.600 2.200 520.400 9.600 ;
        RECT 522.800 9.700 525.800 10.200 ;
        RECT 522.800 2.200 523.600 9.700 ;
        RECT 524.400 9.600 525.800 9.700 ;
        RECT 526.400 9.600 527.400 10.200 ;
        RECT 525.200 8.400 525.800 9.600 ;
        RECT 525.200 7.600 526.000 8.400 ;
        RECT 526.600 2.200 527.400 9.600 ;
        RECT 531.400 9.400 533.200 10.200 ;
        RECT 537.200 9.400 539.000 10.200 ;
        RECT 531.400 2.200 532.200 9.400 ;
        RECT 538.200 2.200 539.000 9.400 ;
        RECT 542.000 2.200 542.800 19.800 ;
        RECT 543.800 16.400 544.600 17.200 ;
        RECT 543.600 15.600 544.400 16.400 ;
        RECT 545.200 15.800 546.000 19.800 ;
        RECT 545.400 14.400 546.000 15.800 ;
        RECT 551.600 17.600 552.400 19.800 ;
        RECT 551.600 14.400 552.200 17.600 ;
        RECT 553.200 15.600 554.000 17.200 ;
        RECT 554.800 15.800 555.600 19.800 ;
        RECT 559.000 18.400 559.800 19.800 ;
        RECT 559.000 17.600 560.400 18.400 ;
        RECT 559.000 16.800 559.800 17.600 ;
        RECT 559.000 15.800 560.400 16.800 ;
        RECT 555.000 15.600 555.600 15.800 ;
        RECT 555.000 15.200 556.800 15.600 ;
        RECT 555.000 15.000 559.200 15.200 ;
        RECT 556.200 14.600 559.200 15.000 ;
        RECT 558.400 14.400 559.200 14.600 ;
        RECT 545.200 13.600 546.000 14.400 ;
        RECT 543.600 12.200 544.400 12.400 ;
        RECT 545.400 12.200 546.000 13.600 ;
        RECT 546.800 12.800 547.600 14.400 ;
        RECT 551.600 13.600 552.400 14.400 ;
        RECT 548.400 12.200 549.200 12.400 ;
        RECT 543.600 11.600 546.000 12.200 ;
        RECT 547.600 11.600 549.200 12.200 ;
        RECT 543.800 10.200 544.400 11.600 ;
        RECT 547.600 11.200 548.400 11.600 ;
        RECT 550.000 10.800 550.800 12.400 ;
        RECT 551.600 10.200 552.200 13.600 ;
        RECT 554.800 12.800 555.600 14.400 ;
        RECT 556.800 13.800 557.600 14.000 ;
        RECT 556.600 13.200 557.600 13.800 ;
        RECT 556.600 12.400 557.200 13.200 ;
        RECT 556.400 11.600 557.200 12.400 ;
        RECT 558.400 11.000 559.000 14.400 ;
        RECT 559.800 12.400 560.400 15.800 ;
        RECT 561.200 15.800 562.000 19.800 ;
        RECT 565.600 16.200 567.200 19.800 ;
        RECT 561.200 15.200 563.600 15.800 ;
        RECT 562.800 15.000 563.600 15.200 ;
        RECT 564.200 14.800 565.000 15.600 ;
        RECT 564.200 14.400 564.800 14.800 ;
        RECT 561.200 13.600 562.800 14.400 ;
        RECT 564.000 13.600 564.800 14.400 ;
        RECT 565.600 12.800 566.200 16.200 ;
        RECT 570.800 15.800 571.600 19.800 ;
        RECT 572.400 16.000 573.200 19.800 ;
        RECT 575.600 16.000 576.400 19.800 ;
        RECT 572.400 15.800 576.400 16.000 ;
        RECT 577.200 15.800 578.000 19.800 ;
        RECT 566.800 15.400 568.400 15.600 ;
        RECT 566.800 14.800 568.800 15.400 ;
        RECT 569.400 15.200 571.600 15.800 ;
        RECT 572.600 15.400 576.200 15.800 ;
        RECT 569.400 15.000 570.200 15.200 ;
        RECT 568.200 14.400 568.800 14.800 ;
        RECT 573.200 14.400 574.000 14.800 ;
        RECT 577.200 14.400 577.800 15.800 ;
        RECT 578.800 15.200 579.600 19.800 ;
        RECT 578.800 14.600 581.000 15.200 ;
        RECT 566.800 13.400 567.600 14.200 ;
        RECT 568.200 13.800 571.600 14.400 ;
        RECT 570.000 13.600 571.600 13.800 ;
        RECT 572.400 13.800 574.000 14.400 ;
        RECT 572.400 13.600 573.200 13.800 ;
        RECT 575.400 13.600 578.000 14.400 ;
        RECT 565.200 12.400 566.200 12.800 ;
        RECT 559.600 11.600 560.400 12.400 ;
        RECT 564.400 12.200 566.200 12.400 ;
        RECT 567.000 12.800 567.600 13.400 ;
        RECT 567.000 12.200 569.600 12.800 ;
        RECT 564.400 11.600 565.800 12.200 ;
        RECT 568.800 12.000 569.600 12.200 ;
        RECT 574.000 11.600 574.800 13.200 ;
        RECT 556.600 10.400 559.000 11.000 ;
        RECT 543.600 2.200 544.400 10.200 ;
        RECT 545.200 9.600 549.200 10.200 ;
        RECT 545.200 2.200 546.000 9.600 ;
        RECT 548.400 2.200 549.200 9.600 ;
        RECT 550.600 9.400 552.400 10.200 ;
        RECT 550.600 2.200 551.400 9.400 ;
        RECT 556.600 6.200 557.200 10.400 ;
        RECT 559.800 10.200 560.400 11.600 ;
        RECT 565.200 10.200 565.800 11.600 ;
        RECT 566.600 11.400 567.400 11.600 ;
        RECT 566.600 10.800 570.000 11.400 ;
        RECT 569.400 10.200 570.000 10.800 ;
        RECT 575.400 10.200 576.000 13.600 ;
        RECT 578.800 11.600 579.600 13.200 ;
        RECT 580.400 11.600 581.000 14.600 ;
        RECT 580.400 10.800 581.600 11.600 ;
        RECT 577.200 10.200 578.000 10.400 ;
        RECT 580.400 10.200 581.000 10.800 ;
        RECT 556.400 2.200 557.200 6.200 ;
        RECT 559.600 2.200 560.400 10.200 ;
        RECT 561.200 9.600 563.600 10.200 ;
        RECT 565.200 9.600 567.200 10.200 ;
        RECT 561.200 2.200 562.000 9.600 ;
        RECT 562.800 9.400 563.600 9.600 ;
        RECT 565.600 2.200 567.200 9.600 ;
        RECT 569.400 9.600 571.600 10.200 ;
        RECT 569.400 9.400 570.200 9.600 ;
        RECT 570.800 2.200 571.600 9.600 ;
        RECT 575.000 9.600 576.000 10.200 ;
        RECT 576.600 9.600 578.000 10.200 ;
        RECT 578.800 9.600 581.000 10.200 ;
        RECT 575.000 2.200 575.800 9.600 ;
        RECT 576.600 8.400 577.200 9.600 ;
        RECT 576.400 7.600 577.200 8.400 ;
        RECT 578.800 2.200 579.600 9.600 ;
      LAYER via1 ;
        RECT 7.600 403.600 8.400 404.400 ;
        RECT 46.000 417.600 46.800 418.400 ;
        RECT 15.600 403.600 16.400 404.400 ;
        RECT 20.400 409.600 21.200 410.400 ;
        RECT 31.600 411.600 32.400 412.400 ;
        RECT 38.000 409.600 38.800 410.400 ;
        RECT 44.400 413.600 45.200 414.400 ;
        RECT 62.000 413.600 62.800 414.400 ;
        RECT 50.800 412.200 51.600 413.000 ;
        RECT 58.800 411.800 59.600 412.600 ;
        RECT 81.200 413.600 82.000 414.400 ;
        RECT 84.400 413.600 85.200 414.400 ;
        RECT 70.000 412.200 70.800 413.000 ;
        RECT 63.600 410.200 64.400 411.000 ;
        RECT 78.000 411.800 78.800 412.600 ;
        RECT 82.800 410.200 83.600 411.000 ;
        RECT 65.200 407.600 66.000 408.400 ;
        RECT 126.000 414.800 126.800 415.600 ;
        RECT 119.600 413.600 120.400 414.400 ;
        RECT 108.400 412.200 109.200 413.000 ;
        RECT 116.400 411.800 117.200 412.600 ;
        RECT 132.400 413.600 133.200 414.400 ;
        RECT 100.400 403.600 101.200 404.400 ;
        RECT 121.200 410.200 122.000 411.000 ;
        RECT 103.600 403.600 104.400 404.400 ;
        RECT 145.200 409.600 146.000 410.400 ;
        RECT 153.200 414.800 154.000 415.600 ;
        RECT 159.600 413.600 160.400 414.400 ;
        RECT 174.000 413.600 174.800 414.400 ;
        RECT 167.600 411.600 168.400 412.400 ;
        RECT 164.400 409.600 165.200 410.400 ;
        RECT 166.000 409.600 166.800 410.400 ;
        RECT 162.800 403.600 163.600 404.400 ;
        RECT 175.600 409.600 176.400 410.400 ;
        RECT 186.800 411.600 187.600 412.400 ;
        RECT 191.600 413.600 192.400 414.400 ;
        RECT 193.200 411.600 194.000 412.400 ;
        RECT 194.800 411.600 195.600 412.400 ;
        RECT 209.200 415.600 210.000 416.400 ;
        RECT 199.600 411.600 200.400 412.400 ;
        RECT 188.400 403.600 189.200 404.400 ;
        RECT 209.200 403.600 210.000 404.400 ;
        RECT 218.800 403.600 219.600 404.400 ;
        RECT 220.400 417.600 221.200 418.400 ;
        RECT 225.200 412.200 226.000 413.000 ;
        RECT 233.200 411.800 234.000 412.600 ;
        RECT 239.600 411.600 240.400 412.400 ;
        RECT 238.000 410.200 238.800 411.000 ;
        RECT 220.400 403.600 221.200 404.400 ;
        RECT 247.600 412.200 248.400 413.000 ;
        RECT 255.600 411.800 256.400 412.600 ;
        RECT 260.400 410.200 261.200 411.000 ;
        RECT 242.800 403.600 243.600 404.400 ;
        RECT 274.800 411.600 275.600 412.400 ;
        RECT 294.000 413.600 294.800 414.400 ;
        RECT 302.000 413.600 302.800 414.400 ;
        RECT 282.800 412.200 283.600 413.000 ;
        RECT 276.400 409.600 277.200 410.400 ;
        RECT 295.600 410.200 296.400 411.000 ;
        RECT 278.000 405.600 278.800 406.400 ;
        RECT 321.200 412.200 322.000 413.000 ;
        RECT 329.200 411.800 330.000 412.600 ;
        RECT 334.000 410.200 334.800 411.000 ;
        RECT 316.400 403.600 317.200 404.400 ;
        RECT 340.400 413.600 341.200 414.400 ;
        RECT 372.400 415.600 373.200 416.400 ;
        RECT 374.000 414.200 374.800 415.000 ;
        RECT 385.200 411.600 386.000 412.400 ;
        RECT 356.400 403.600 357.200 404.400 ;
        RECT 367.600 406.800 368.400 407.600 ;
        RECT 370.800 406.200 371.600 407.000 ;
        RECT 366.000 404.200 366.800 405.000 ;
        RECT 367.600 404.200 368.400 405.000 ;
        RECT 369.200 404.200 370.000 405.000 ;
        RECT 374.000 406.200 374.800 407.000 ;
        RECT 377.200 406.200 378.000 407.000 ;
        RECT 378.800 404.200 379.600 405.000 ;
        RECT 380.400 404.200 381.200 405.000 ;
        RECT 418.800 415.600 419.600 416.400 ;
        RECT 420.400 414.200 421.200 415.000 ;
        RECT 431.600 411.600 432.400 412.400 ;
        RECT 402.800 403.600 403.600 404.400 ;
        RECT 414.000 406.800 414.800 407.600 ;
        RECT 417.200 406.200 418.000 407.000 ;
        RECT 412.400 404.200 413.200 405.000 ;
        RECT 414.000 404.200 414.800 405.000 ;
        RECT 415.600 404.200 416.400 405.000 ;
        RECT 420.400 406.200 421.200 407.000 ;
        RECT 423.600 406.200 424.400 407.000 ;
        RECT 425.200 404.200 426.000 405.000 ;
        RECT 426.800 404.200 427.600 405.000 ;
        RECT 479.600 415.600 480.400 416.400 ;
        RECT 481.200 414.200 482.000 415.000 ;
        RECT 492.400 411.600 493.200 412.400 ;
        RECT 463.600 403.600 464.400 404.400 ;
        RECT 474.800 406.800 475.600 407.600 ;
        RECT 478.000 406.200 478.800 407.000 ;
        RECT 473.200 404.200 474.000 405.000 ;
        RECT 474.800 404.200 475.600 405.000 ;
        RECT 476.400 404.200 477.200 405.000 ;
        RECT 481.200 406.200 482.000 407.000 ;
        RECT 484.400 406.200 485.200 407.000 ;
        RECT 486.000 404.200 486.800 405.000 ;
        RECT 487.600 404.200 488.400 405.000 ;
        RECT 521.200 413.000 522.000 413.800 ;
        RECT 530.800 412.600 531.600 413.400 ;
        RECT 514.800 411.600 515.600 412.400 ;
        RECT 537.200 411.600 538.000 412.400 ;
        RECT 522.800 408.800 523.600 409.600 ;
        RECT 527.600 407.600 528.400 408.400 ;
        RECT 524.400 406.200 525.200 407.000 ;
        RECT 521.200 404.200 522.000 405.000 ;
        RECT 522.800 404.200 523.600 405.000 ;
        RECT 527.600 406.200 528.400 407.000 ;
        RECT 530.800 406.200 531.600 407.000 ;
        RECT 532.400 404.200 533.200 405.000 ;
        RECT 534.000 404.200 534.800 405.000 ;
        RECT 535.600 404.200 536.400 405.000 ;
        RECT 566.000 415.600 566.800 416.400 ;
        RECT 567.600 414.200 568.400 415.000 ;
        RECT 558.000 411.600 558.800 412.400 ;
        RECT 545.200 403.600 546.000 404.400 ;
        RECT 550.000 403.600 550.800 404.400 ;
        RECT 561.200 406.800 562.000 407.600 ;
        RECT 564.400 406.200 565.200 407.000 ;
        RECT 559.600 404.200 560.400 405.000 ;
        RECT 561.200 404.200 562.000 405.000 ;
        RECT 562.800 404.200 563.600 405.000 ;
        RECT 567.600 406.200 568.400 407.000 ;
        RECT 570.800 406.200 571.600 407.000 ;
        RECT 572.400 404.200 573.200 405.000 ;
        RECT 574.000 404.200 574.800 405.000 ;
        RECT 2.800 389.600 3.600 390.400 ;
        RECT 7.600 387.600 8.400 388.400 ;
        RECT 15.600 387.600 16.400 388.400 ;
        RECT 20.400 387.600 21.200 388.400 ;
        RECT 22.000 387.600 22.800 388.400 ;
        RECT 6.000 383.600 6.800 384.400 ;
        RECT 41.200 391.600 42.000 392.400 ;
        RECT 30.000 385.600 30.800 386.400 ;
        RECT 41.200 389.600 42.000 390.400 ;
        RECT 42.800 387.600 43.600 388.400 ;
        RECT 47.600 387.600 48.400 388.400 ;
        RECT 49.200 387.600 50.000 388.400 ;
        RECT 66.800 391.800 67.600 392.600 ;
        RECT 34.800 383.600 35.600 384.400 ;
        RECT 57.200 385.600 58.000 386.400 ;
        RECT 60.400 383.600 61.200 384.400 ;
        RECT 66.800 386.200 67.600 387.000 ;
        RECT 74.800 387.600 75.600 388.400 ;
        RECT 71.600 386.400 72.400 387.200 ;
        RECT 70.000 383.600 70.800 384.400 ;
        RECT 76.400 385.600 77.200 386.400 ;
        RECT 89.200 389.600 90.000 390.400 ;
        RECT 82.800 387.600 83.600 388.400 ;
        RECT 100.400 387.600 101.200 388.400 ;
        RECT 94.000 383.600 94.800 384.400 ;
        RECT 108.400 387.600 109.200 388.400 ;
        RECT 127.600 392.400 128.400 393.200 ;
        RECT 138.600 391.800 139.400 392.600 ;
        RECT 149.800 391.800 150.600 392.600 ;
        RECT 130.800 391.000 131.600 391.800 ;
        RECT 111.600 385.600 112.400 386.400 ;
        RECT 130.800 386.200 131.600 387.000 ;
        RECT 113.200 383.600 114.000 384.400 ;
        RECT 138.600 386.200 139.400 387.000 ;
        RECT 161.200 389.600 162.000 390.400 ;
        RECT 146.800 387.600 147.600 388.400 ;
        RECT 149.800 386.200 150.600 387.000 ;
        RECT 169.200 389.600 170.000 390.400 ;
        RECT 158.000 387.600 158.800 388.400 ;
        RECT 162.800 387.600 163.600 388.400 ;
        RECT 170.800 387.600 171.600 388.400 ;
        RECT 178.800 389.600 179.600 390.400 ;
        RECT 186.800 389.600 187.600 390.400 ;
        RECT 175.600 387.600 176.400 388.400 ;
        RECT 188.400 387.600 189.200 388.400 ;
        RECT 190.000 387.600 190.800 388.400 ;
        RECT 194.800 391.600 195.600 392.400 ;
        RECT 199.600 389.600 200.400 390.400 ;
        RECT 196.400 387.600 197.200 388.400 ;
        RECT 201.200 387.600 202.000 388.400 ;
        RECT 226.800 397.600 227.600 398.400 ;
        RECT 204.400 385.600 205.200 386.400 ;
        RECT 218.800 385.600 219.600 386.400 ;
        RECT 223.600 387.600 224.400 388.400 ;
        RECT 228.400 387.600 229.200 388.400 ;
        RECT 257.000 391.800 257.800 392.600 ;
        RECT 230.000 385.600 230.800 386.400 ;
        RECT 242.800 387.600 243.600 388.400 ;
        RECT 246.000 383.600 246.800 384.400 ;
        RECT 252.400 383.600 253.200 384.400 ;
        RECT 257.000 386.200 257.800 387.000 ;
        RECT 270.000 387.600 270.800 388.400 ;
        RECT 284.200 391.800 285.000 392.600 ;
        RECT 305.200 397.600 306.000 398.400 ;
        RECT 274.800 387.600 275.600 388.400 ;
        RECT 284.200 386.200 285.000 387.000 ;
        RECT 273.200 383.600 274.000 384.400 ;
        RECT 281.200 383.600 282.000 384.400 ;
        RECT 292.400 387.600 293.200 388.400 ;
        RECT 287.600 383.600 288.400 384.400 ;
        RECT 298.800 385.600 299.600 386.400 ;
        RECT 303.600 387.600 304.400 388.400 ;
        RECT 316.400 389.600 317.200 390.400 ;
        RECT 321.200 389.600 322.000 390.400 ;
        RECT 326.000 391.600 326.800 392.400 ;
        RECT 311.600 387.600 312.400 388.400 ;
        RECT 318.000 387.600 318.800 388.400 ;
        RECT 322.800 387.600 323.600 388.400 ;
        RECT 310.000 383.600 310.800 384.400 ;
        RECT 343.600 392.400 344.400 393.200 ;
        RECT 346.800 391.000 347.600 391.800 ;
        RECT 353.200 389.600 354.000 390.400 ;
        RECT 327.600 385.600 328.400 386.400 ;
        RECT 346.800 386.200 347.600 387.000 ;
        RECT 351.600 385.600 352.400 386.400 ;
        RECT 358.000 387.600 358.800 388.400 ;
        RECT 364.400 385.600 365.200 386.400 ;
        RECT 362.800 383.600 363.600 384.400 ;
        RECT 369.200 389.600 370.000 390.400 ;
        RECT 374.000 389.600 374.800 390.400 ;
        RECT 404.400 392.400 405.200 393.200 ;
        RECT 407.600 391.000 408.400 391.800 ;
        RECT 402.800 385.600 403.600 386.400 ;
        RECT 390.000 383.600 390.800 384.400 ;
        RECT 407.600 386.200 408.400 387.000 ;
        RECT 414.000 389.600 414.800 390.400 ;
        RECT 418.800 389.600 419.600 390.400 ;
        RECT 423.600 389.600 424.400 390.400 ;
        RECT 422.000 387.600 422.800 388.400 ;
        RECT 428.400 389.600 429.200 390.400 ;
        RECT 455.600 394.400 456.400 395.200 ;
        RECT 458.800 395.000 459.600 395.800 ;
        RECT 454.000 392.400 454.800 393.200 ;
        RECT 444.400 383.600 445.200 384.400 ;
        RECT 460.400 385.600 461.200 386.400 ;
        RECT 454.000 384.200 454.800 385.000 ;
        RECT 455.600 384.200 456.400 385.000 ;
        RECT 457.200 384.200 458.000 385.000 ;
        RECT 458.800 384.200 459.600 385.000 ;
        RECT 462.000 384.200 462.800 385.000 ;
        RECT 465.200 384.200 466.000 385.000 ;
        RECT 466.800 384.200 467.600 385.000 ;
        RECT 468.400 384.200 469.200 385.000 ;
        RECT 487.600 385.600 488.400 386.400 ;
        RECT 498.800 389.600 499.600 390.400 ;
        RECT 495.600 385.600 496.400 386.400 ;
        RECT 490.800 383.600 491.600 384.400 ;
        RECT 505.200 389.600 506.000 390.400 ;
        RECT 510.000 389.600 510.800 390.400 ;
        RECT 529.200 395.000 530.000 395.800 ;
        RECT 526.000 393.600 526.800 394.400 ;
        RECT 543.600 397.600 544.400 398.400 ;
        RECT 530.800 392.400 531.600 393.200 ;
        RECT 519.600 388.200 520.400 389.000 ;
        RECT 529.200 388.600 530.000 389.400 ;
        RECT 502.000 383.600 502.800 384.400 ;
        RECT 524.400 387.600 525.200 388.400 ;
        RECT 519.600 384.200 520.400 385.000 ;
        RECT 521.200 384.200 522.000 385.000 ;
        RECT 522.800 384.200 523.600 385.000 ;
        RECT 526.000 384.200 526.800 385.000 ;
        RECT 529.200 384.200 530.000 385.000 ;
        RECT 530.800 384.200 531.600 385.000 ;
        RECT 532.400 384.200 533.200 385.000 ;
        RECT 534.000 384.200 534.800 385.000 ;
        RECT 564.400 395.000 565.200 395.800 ;
        RECT 561.200 393.600 562.000 394.400 ;
        RECT 566.000 392.400 566.800 393.200 ;
        RECT 554.800 388.200 555.600 389.000 ;
        RECT 564.400 388.600 565.200 389.400 ;
        RECT 559.600 387.600 560.400 388.400 ;
        RECT 554.800 384.200 555.600 385.000 ;
        RECT 556.400 384.200 557.200 385.000 ;
        RECT 558.000 384.200 558.800 385.000 ;
        RECT 561.200 384.200 562.000 385.000 ;
        RECT 564.400 384.200 565.200 385.000 ;
        RECT 566.000 384.200 566.800 385.000 ;
        RECT 567.600 384.200 568.400 385.000 ;
        RECT 569.200 384.200 570.000 385.000 ;
        RECT 578.800 383.600 579.600 384.400 ;
        RECT 17.200 373.600 18.000 374.400 ;
        RECT 14.000 367.600 14.800 368.400 ;
        RECT 41.200 377.600 42.000 378.400 ;
        RECT 26.800 369.600 27.600 370.400 ;
        RECT 28.400 369.600 29.200 370.400 ;
        RECT 34.800 371.600 35.600 372.400 ;
        RECT 65.200 373.600 66.000 374.400 ;
        RECT 54.000 372.200 54.800 373.000 ;
        RECT 62.000 371.800 62.800 372.600 ;
        RECT 66.800 370.200 67.600 371.000 ;
        RECT 49.200 363.600 50.000 364.400 ;
        RECT 73.200 373.600 74.000 374.400 ;
        RECT 68.400 369.600 69.200 370.400 ;
        RECT 74.800 363.600 75.600 364.400 ;
        RECT 82.800 372.200 83.600 373.000 ;
        RECT 90.800 371.800 91.600 372.600 ;
        RECT 102.000 372.200 102.800 373.000 ;
        RECT 95.600 370.200 96.400 371.000 ;
        RECT 78.000 363.600 78.800 364.400 ;
        RECT 110.000 371.800 110.800 372.600 ;
        RECT 121.200 372.200 122.000 373.000 ;
        RECT 114.800 370.200 115.600 371.000 ;
        RECT 97.200 367.600 98.000 368.400 ;
        RECT 150.000 373.600 150.800 374.400 ;
        RECT 145.200 372.200 146.000 373.000 ;
        RECT 134.000 370.200 134.800 371.000 ;
        RECT 116.400 365.600 117.200 366.400 ;
        RECT 166.000 374.800 166.800 375.600 ;
        RECT 153.200 371.800 154.000 372.600 ;
        RECT 172.400 371.600 173.200 372.400 ;
        RECT 158.000 370.200 158.800 371.000 ;
        RECT 140.400 363.600 141.200 364.400 ;
        RECT 183.600 371.600 184.400 372.400 ;
        RECT 191.600 369.600 192.400 370.400 ;
        RECT 190.000 363.600 190.800 364.400 ;
        RECT 202.800 375.600 203.600 376.400 ;
        RECT 199.600 369.600 200.400 370.400 ;
        RECT 204.400 369.600 205.200 370.400 ;
        RECT 217.200 369.600 218.000 370.400 ;
        RECT 222.000 369.600 222.800 370.400 ;
        RECT 225.200 369.600 226.000 370.400 ;
        RECT 239.600 373.600 240.400 374.400 ;
        RECT 246.000 377.600 246.800 378.400 ;
        RECT 262.000 377.600 262.800 378.400 ;
        RECT 271.600 377.600 272.400 378.400 ;
        RECT 250.800 373.600 251.600 374.400 ;
        RECT 249.200 371.600 250.000 372.400 ;
        RECT 255.600 367.600 256.400 368.400 ;
        RECT 262.000 369.600 262.800 370.400 ;
        RECT 273.200 373.600 274.000 374.400 ;
        RECT 287.600 375.600 288.400 376.400 ;
        RECT 282.800 373.600 283.600 374.400 ;
        RECT 274.800 371.600 275.600 372.400 ;
        RECT 276.400 371.600 277.200 372.400 ;
        RECT 266.800 363.600 267.600 364.400 ;
        RECT 286.000 369.600 286.800 370.400 ;
        RECT 311.600 377.600 312.400 378.400 ;
        RECT 330.800 377.600 331.600 378.400 ;
        RECT 316.400 372.200 317.200 373.000 ;
        RECT 310.000 369.600 310.800 370.400 ;
        RECT 324.400 371.800 325.200 372.600 ;
        RECT 335.600 372.200 336.400 373.000 ;
        RECT 329.200 370.200 330.000 371.000 ;
        RECT 343.600 371.800 344.400 372.600 ;
        RECT 353.200 371.600 354.000 372.400 ;
        RECT 348.400 370.200 349.200 371.000 ;
        RECT 354.800 369.600 355.600 370.400 ;
        RECT 364.400 371.600 365.200 372.400 ;
        RECT 367.600 371.600 368.400 372.400 ;
        RECT 366.000 369.600 366.800 370.400 ;
        RECT 375.600 371.600 376.400 372.400 ;
        RECT 386.800 377.600 387.600 378.400 ;
        RECT 369.200 363.600 370.000 364.400 ;
        RECT 380.400 367.600 381.200 368.400 ;
        RECT 391.600 372.200 392.400 373.000 ;
        RECT 399.600 371.800 400.400 372.600 ;
        RECT 404.400 370.200 405.200 371.000 ;
        RECT 428.400 375.600 429.200 376.400 ;
        RECT 430.000 374.200 430.800 375.000 ;
        RECT 441.200 371.600 442.000 372.400 ;
        RECT 438.000 370.000 438.800 370.800 ;
        RECT 412.400 363.600 413.200 364.400 ;
        RECT 423.600 366.800 424.400 367.600 ;
        RECT 426.800 366.200 427.600 367.000 ;
        RECT 422.000 364.200 422.800 365.000 ;
        RECT 423.600 364.200 424.400 365.000 ;
        RECT 425.200 364.200 426.000 365.000 ;
        RECT 430.000 366.200 430.800 367.000 ;
        RECT 433.200 366.200 434.000 367.000 ;
        RECT 434.800 364.200 435.600 365.000 ;
        RECT 436.400 364.200 437.200 365.000 ;
        RECT 474.800 375.600 475.600 376.400 ;
        RECT 476.400 374.200 477.200 375.000 ;
        RECT 487.600 371.600 488.400 372.400 ;
        RECT 458.800 363.600 459.600 364.400 ;
        RECT 470.000 366.800 470.800 367.600 ;
        RECT 473.200 366.200 474.000 367.000 ;
        RECT 468.400 364.200 469.200 365.000 ;
        RECT 470.000 364.200 470.800 365.000 ;
        RECT 471.600 364.200 472.400 365.000 ;
        RECT 476.400 366.200 477.200 367.000 ;
        RECT 479.600 366.200 480.400 367.000 ;
        RECT 506.800 373.000 507.600 373.800 ;
        RECT 481.200 364.200 482.000 365.000 ;
        RECT 482.800 364.200 483.600 365.000 ;
        RECT 516.400 372.600 517.200 373.400 ;
        RECT 530.800 377.600 531.600 378.400 ;
        RECT 502.000 371.600 502.800 372.400 ;
        RECT 508.400 368.800 509.200 369.600 ;
        RECT 513.200 367.600 514.000 368.400 ;
        RECT 510.000 366.200 510.800 367.000 ;
        RECT 506.800 364.200 507.600 365.000 ;
        RECT 508.400 364.200 509.200 365.000 ;
        RECT 513.200 366.200 514.000 367.000 ;
        RECT 516.400 366.200 517.200 367.000 ;
        RECT 518.000 364.200 518.800 365.000 ;
        RECT 519.600 364.200 520.400 365.000 ;
        RECT 521.200 364.200 522.000 365.000 ;
        RECT 535.600 363.600 536.400 364.400 ;
        RECT 556.400 373.000 557.200 373.800 ;
        RECT 566.000 372.600 566.800 373.400 ;
        RECT 580.400 377.600 581.200 378.400 ;
        RECT 551.600 371.600 552.400 372.400 ;
        RECT 558.000 368.800 558.800 369.600 ;
        RECT 562.800 367.600 563.600 368.400 ;
        RECT 545.200 363.600 546.000 364.400 ;
        RECT 559.600 366.200 560.400 367.000 ;
        RECT 556.400 364.200 557.200 365.000 ;
        RECT 558.000 364.200 558.800 365.000 ;
        RECT 562.800 366.200 563.600 367.000 ;
        RECT 566.000 366.200 566.800 367.000 ;
        RECT 567.600 364.200 568.400 365.000 ;
        RECT 569.200 364.200 570.000 365.000 ;
        RECT 570.800 364.200 571.600 365.000 ;
        RECT 4.400 351.600 5.200 352.400 ;
        RECT 9.000 351.800 9.800 352.600 ;
        RECT 20.400 357.600 21.200 358.400 ;
        RECT 4.400 349.600 5.200 350.400 ;
        RECT 6.000 347.600 6.800 348.400 ;
        RECT 9.000 346.200 9.800 347.000 ;
        RECT 17.200 347.600 18.000 348.400 ;
        RECT 12.400 343.600 13.200 344.400 ;
        RECT 18.800 345.600 19.600 346.400 ;
        RECT 23.400 351.800 24.200 352.600 ;
        RECT 28.400 351.600 29.200 352.400 ;
        RECT 34.800 357.600 35.600 358.400 ;
        RECT 20.400 343.600 21.200 344.400 ;
        RECT 23.400 346.200 24.200 347.000 ;
        RECT 33.200 345.600 34.000 346.400 ;
        RECT 36.400 345.600 37.200 346.400 ;
        RECT 34.800 343.600 35.600 344.400 ;
        RECT 52.400 349.600 53.200 350.400 ;
        RECT 57.200 349.600 58.000 350.400 ;
        RECT 50.800 347.600 51.600 348.400 ;
        RECT 54.000 347.600 54.800 348.400 ;
        RECT 44.400 343.600 45.200 344.400 ;
        RECT 73.200 345.600 74.000 346.400 ;
        RECT 74.800 343.600 75.600 344.400 ;
        RECT 84.400 345.600 85.200 346.400 ;
        RECT 81.200 343.600 82.000 344.400 ;
        RECT 108.400 352.400 109.200 353.200 ;
        RECT 111.600 351.000 112.400 351.800 ;
        RECT 111.600 346.200 112.400 347.000 ;
        RECT 116.400 347.600 117.200 348.400 ;
        RECT 94.000 343.600 94.800 344.400 ;
        RECT 123.000 351.800 123.800 352.600 ;
        RECT 124.200 349.800 125.000 350.600 ;
        RECT 119.600 347.600 120.400 348.400 ;
        RECT 118.000 343.600 118.800 344.400 ;
        RECT 123.000 346.200 123.800 347.000 ;
        RECT 130.800 347.600 131.600 348.400 ;
        RECT 132.400 347.600 133.200 348.400 ;
        RECT 127.600 343.600 128.400 344.400 ;
        RECT 143.800 351.800 144.600 352.600 ;
        RECT 145.000 349.800 145.800 350.600 ;
        RECT 143.800 346.200 144.600 347.000 ;
        RECT 151.600 347.600 152.400 348.400 ;
        RECT 167.600 352.400 168.400 353.200 ;
        RECT 170.800 351.000 171.600 351.800 ;
        RECT 148.400 343.600 149.200 344.400 ;
        RECT 186.800 352.400 187.600 353.200 ;
        RECT 198.200 351.800 199.000 352.600 ;
        RECT 190.000 351.000 190.800 351.800 ;
        RECT 223.800 351.800 224.600 352.600 ;
        RECT 199.400 349.800 200.200 350.600 ;
        RECT 170.800 346.200 171.600 347.000 ;
        RECT 153.200 343.600 154.000 344.400 ;
        RECT 209.200 349.600 210.000 350.400 ;
        RECT 190.000 346.200 190.800 347.000 ;
        RECT 172.400 343.600 173.200 344.400 ;
        RECT 194.800 345.600 195.600 346.400 ;
        RECT 198.200 346.200 199.000 347.000 ;
        RECT 206.000 347.600 206.800 348.400 ;
        RECT 214.000 347.600 214.800 348.400 ;
        RECT 209.200 345.600 210.000 346.400 ;
        RECT 225.000 349.800 225.800 350.600 ;
        RECT 236.400 349.600 237.200 350.400 ;
        RECT 223.800 346.200 224.600 347.000 ;
        RECT 231.600 347.600 232.400 348.400 ;
        RECT 238.000 347.600 238.800 348.400 ;
        RECT 242.800 347.600 243.600 348.400 ;
        RECT 244.400 347.600 245.200 348.400 ;
        RECT 250.800 357.600 251.600 358.400 ;
        RECT 249.200 347.600 250.000 348.400 ;
        RECT 241.200 343.600 242.000 344.400 ;
        RECT 247.600 343.600 248.400 344.400 ;
        RECT 255.600 351.600 256.400 352.400 ;
        RECT 254.000 347.600 254.800 348.400 ;
        RECT 262.000 357.600 262.800 358.400 ;
        RECT 266.600 351.800 267.400 352.600 ;
        RECT 263.600 347.600 264.400 348.400 ;
        RECT 262.000 343.600 262.800 344.400 ;
        RECT 266.600 346.200 267.400 347.000 ;
        RECT 274.800 347.600 275.600 348.400 ;
        RECT 286.000 347.600 286.800 348.400 ;
        RECT 295.600 345.600 296.400 346.400 ;
        RECT 302.000 345.600 302.800 346.400 ;
        RECT 326.000 355.600 326.800 356.400 ;
        RECT 308.400 345.600 309.200 346.400 ;
        RECT 310.000 345.600 310.800 346.400 ;
        RECT 311.600 343.600 312.400 344.400 ;
        RECT 326.000 349.600 326.800 350.400 ;
        RECT 321.200 345.600 322.000 346.400 ;
        RECT 327.600 347.600 328.400 348.400 ;
        RECT 319.600 343.600 320.400 344.400 ;
        RECT 346.800 352.400 347.600 353.200 ;
        RECT 350.000 351.000 350.800 351.800 ;
        RECT 351.600 349.600 352.400 350.400 ;
        RECT 330.800 345.600 331.600 346.400 ;
        RECT 345.200 345.600 346.000 346.400 ;
        RECT 350.000 346.200 350.800 347.000 ;
        RECT 369.200 352.400 370.000 353.200 ;
        RECT 380.200 351.800 381.000 352.600 ;
        RECT 372.400 351.000 373.200 351.800 ;
        RECT 374.000 349.600 374.800 350.400 ;
        RECT 353.200 345.600 354.000 346.400 ;
        RECT 367.600 345.600 368.400 346.400 ;
        RECT 354.800 343.600 355.600 344.400 ;
        RECT 372.400 346.200 373.200 347.000 ;
        RECT 380.200 346.200 381.000 347.000 ;
        RECT 383.600 343.600 384.400 344.400 ;
        RECT 391.600 347.600 392.400 348.400 ;
        RECT 407.600 352.400 408.400 353.200 ;
        RECT 410.800 351.000 411.600 351.800 ;
        RECT 415.600 349.600 416.400 350.400 ;
        RECT 426.800 349.600 427.600 350.400 ;
        RECT 434.800 349.600 435.600 350.400 ;
        RECT 390.000 343.600 390.800 344.400 ;
        RECT 410.800 346.200 411.600 347.000 ;
        RECT 417.200 347.600 418.000 348.400 ;
        RECT 423.600 347.600 424.400 348.400 ;
        RECT 438.000 347.600 438.800 348.400 ;
        RECT 393.200 343.600 394.000 344.400 ;
        RECT 430.000 343.600 430.800 344.400 ;
        RECT 441.200 351.600 442.000 352.400 ;
        RECT 439.600 345.600 440.400 346.400 ;
        RECT 442.800 345.600 443.600 346.400 ;
        RECT 449.200 345.600 450.000 346.400 ;
        RECT 454.000 347.600 454.800 348.400 ;
        RECT 471.600 351.800 472.400 352.600 ;
        RECT 481.200 357.600 482.000 358.400 ;
        RECT 471.600 346.200 472.400 347.000 ;
        RECT 460.400 343.600 461.200 344.400 ;
        RECT 468.400 343.600 469.200 344.400 ;
        RECT 476.400 346.400 477.200 347.200 ;
        RECT 495.600 352.400 496.400 353.200 ;
        RECT 498.800 351.000 499.600 351.800 ;
        RECT 511.600 357.600 512.400 358.400 ;
        RECT 498.800 346.200 499.600 347.000 ;
        RECT 532.400 355.000 533.200 355.800 ;
        RECT 529.200 353.600 530.000 354.400 ;
        RECT 534.000 352.400 534.800 353.200 ;
        RECT 522.800 348.200 523.600 349.000 ;
        RECT 532.400 348.600 533.200 349.400 ;
        RECT 511.600 343.600 512.400 344.400 ;
        RECT 527.600 347.600 528.400 348.400 ;
        RECT 547.000 347.600 547.800 348.400 ;
        RECT 522.800 344.200 523.600 345.000 ;
        RECT 524.400 344.200 525.200 345.000 ;
        RECT 526.000 344.200 526.800 345.000 ;
        RECT 529.200 344.200 530.000 345.000 ;
        RECT 532.400 344.200 533.200 345.000 ;
        RECT 534.000 344.200 534.800 345.000 ;
        RECT 535.600 344.200 536.400 345.000 ;
        RECT 537.200 344.200 538.000 345.000 ;
        RECT 567.600 355.000 568.400 355.800 ;
        RECT 564.400 353.600 565.200 354.400 ;
        RECT 569.200 352.400 570.000 353.200 ;
        RECT 558.000 348.200 558.800 349.000 ;
        RECT 567.600 348.600 568.400 349.400 ;
        RECT 562.800 347.600 563.600 348.400 ;
        RECT 558.000 344.200 558.800 345.000 ;
        RECT 559.600 344.200 560.400 345.000 ;
        RECT 561.200 344.200 562.000 345.000 ;
        RECT 564.400 344.200 565.200 345.000 ;
        RECT 567.600 344.200 568.400 345.000 ;
        RECT 569.200 344.200 570.000 345.000 ;
        RECT 570.800 344.200 571.600 345.000 ;
        RECT 572.400 344.200 573.200 345.000 ;
        RECT 582.000 343.600 582.800 344.400 ;
        RECT 4.400 334.800 5.200 335.600 ;
        RECT 22.000 337.600 22.800 338.400 ;
        RECT 10.800 333.600 11.600 334.400 ;
        RECT 6.000 323.600 6.800 324.400 ;
        RECT 25.200 331.600 26.000 332.400 ;
        RECT 22.000 323.600 22.800 324.400 ;
        RECT 38.000 333.600 38.800 334.400 ;
        RECT 28.400 323.600 29.200 324.400 ;
        RECT 33.200 323.600 34.000 324.400 ;
        RECT 41.200 323.600 42.000 324.400 ;
        RECT 54.000 331.600 54.800 332.400 ;
        RECT 47.600 327.600 48.400 328.400 ;
        RECT 54.000 323.600 54.800 324.400 ;
        RECT 71.600 331.600 72.400 332.400 ;
        RECT 66.800 329.600 67.600 330.400 ;
        RECT 65.200 327.600 66.000 328.400 ;
        RECT 71.600 325.600 72.400 326.400 ;
        RECT 78.000 323.600 78.800 324.400 ;
        RECT 113.200 337.600 114.000 338.400 ;
        RECT 86.000 329.600 86.800 330.400 ;
        RECT 118.000 333.600 118.800 334.400 ;
        RECT 146.800 334.800 147.600 335.600 ;
        RECT 134.000 333.600 134.800 334.400 ;
        RECT 100.400 323.600 101.200 324.400 ;
        RECT 113.200 329.600 114.000 330.400 ;
        RECT 130.800 329.600 131.600 330.400 ;
        RECT 156.400 333.600 157.200 334.400 ;
        RECT 180.400 334.800 181.200 335.600 ;
        RECT 183.600 333.600 184.400 334.400 ;
        RECT 186.800 323.600 187.600 324.400 ;
        RECT 210.800 333.600 211.600 334.400 ;
        RECT 204.400 332.200 205.200 333.000 ;
        RECT 225.200 334.800 226.000 335.600 ;
        RECT 228.400 333.600 229.200 334.400 ;
        RECT 236.400 334.800 237.200 335.600 ;
        RECT 212.400 331.800 213.200 332.600 ;
        RECT 239.600 333.600 240.400 334.400 ;
        RECT 217.200 330.200 218.000 331.000 ;
        RECT 199.600 323.600 200.400 324.400 ;
        RECT 247.600 329.600 248.400 330.400 ;
        RECT 266.800 337.600 267.600 338.400 ;
        RECT 244.400 323.600 245.200 324.400 ;
        RECT 265.200 333.600 266.000 334.400 ;
        RECT 273.200 331.600 274.000 332.400 ;
        RECT 260.400 323.600 261.200 324.400 ;
        RECT 279.600 329.600 280.400 330.400 ;
        RECT 295.600 331.600 296.400 332.400 ;
        RECT 326.000 334.800 326.800 335.600 ;
        RECT 314.800 333.600 315.600 334.400 ;
        RECT 289.200 323.600 290.000 324.400 ;
        RECT 310.000 329.600 310.800 330.400 ;
        RECT 321.200 331.600 322.000 332.400 ;
        RECT 334.000 337.600 334.800 338.400 ;
        RECT 332.400 333.600 333.200 334.400 ;
        RECT 345.200 333.600 346.000 334.400 ;
        RECT 338.800 332.200 339.600 333.000 ;
        RECT 346.800 331.800 347.600 332.600 ;
        RECT 356.400 337.600 357.200 338.400 ;
        RECT 353.200 331.600 354.000 332.400 ;
        RECT 351.600 330.200 352.400 331.000 ;
        RECT 367.600 333.600 368.400 334.400 ;
        RECT 382.000 333.600 382.800 334.400 ;
        RECT 361.200 332.200 362.000 333.000 ;
        RECT 369.200 331.800 370.000 332.600 ;
        RECT 374.000 330.200 374.800 331.000 ;
        RECT 410.800 333.600 411.600 334.400 ;
        RECT 399.600 332.200 400.400 333.000 ;
        RECT 393.200 329.600 394.000 330.400 ;
        RECT 407.600 331.800 408.400 332.600 ;
        RECT 423.600 333.600 424.400 334.400 ;
        RECT 436.400 334.800 437.200 335.600 ;
        RECT 418.800 332.200 419.600 333.000 ;
        RECT 412.400 330.200 413.200 331.000 ;
        RECT 394.800 323.600 395.600 324.400 ;
        RECT 426.800 331.800 427.600 332.600 ;
        RECT 474.800 337.600 475.600 338.400 ;
        RECT 494.000 337.600 494.800 338.400 ;
        RECT 431.600 330.200 432.400 331.000 ;
        RECT 460.400 331.600 461.200 332.400 ;
        RECT 414.000 323.600 414.800 324.400 ;
        RECT 458.800 329.600 459.600 330.400 ;
        RECT 513.200 337.600 514.000 338.400 ;
        RECT 474.800 329.600 475.600 330.400 ;
        RECT 476.400 330.200 477.200 331.000 ;
        RECT 497.200 333.600 498.000 334.400 ;
        RECT 500.400 331.800 501.200 332.600 ;
        RECT 495.600 330.200 496.400 331.000 ;
        RECT 521.200 337.600 522.000 338.400 ;
        RECT 537.200 335.600 538.000 336.400 ;
        RECT 538.800 334.200 539.600 335.000 ;
        RECT 546.800 331.600 547.600 332.400 ;
        RECT 532.400 326.800 533.200 327.600 ;
        RECT 535.600 326.200 536.400 327.000 ;
        RECT 530.800 324.200 531.600 325.000 ;
        RECT 532.400 324.200 533.200 325.000 ;
        RECT 534.000 324.200 534.800 325.000 ;
        RECT 538.800 326.200 539.600 327.000 ;
        RECT 542.000 326.200 542.800 327.000 ;
        RECT 559.600 332.200 560.400 333.000 ;
        RECT 543.600 324.200 544.400 325.000 ;
        RECT 545.200 324.200 546.000 325.000 ;
        RECT 572.400 330.200 573.200 331.000 ;
        RECT 554.800 323.600 555.600 324.400 ;
        RECT 4.400 309.600 5.200 310.400 ;
        RECT 1.200 303.600 2.000 304.400 ;
        RECT 17.200 307.600 18.000 308.400 ;
        RECT 14.000 303.600 14.800 304.400 ;
        RECT 28.400 309.600 29.200 310.400 ;
        RECT 26.800 307.600 27.600 308.400 ;
        RECT 23.600 305.600 24.400 306.400 ;
        RECT 30.000 307.600 30.800 308.400 ;
        RECT 49.200 311.600 50.000 312.400 ;
        RECT 53.800 311.800 54.600 312.600 ;
        RECT 34.800 307.600 35.600 308.400 ;
        RECT 41.200 307.600 42.000 308.400 ;
        RECT 39.600 305.600 40.400 306.400 ;
        RECT 49.200 309.600 50.000 310.400 ;
        RECT 50.800 307.600 51.600 308.400 ;
        RECT 53.800 306.200 54.600 307.000 ;
        RECT 33.200 303.600 34.000 304.400 ;
        RECT 38.000 303.600 38.800 304.400 ;
        RECT 62.000 307.600 62.800 308.400 ;
        RECT 74.800 317.600 75.600 318.400 ;
        RECT 70.000 307.600 70.800 308.400 ;
        RECT 68.400 305.600 69.200 306.400 ;
        RECT 65.200 303.600 66.000 304.400 ;
        RECT 86.000 307.600 86.800 308.400 ;
        RECT 81.200 303.600 82.000 304.400 ;
        RECT 95.600 309.600 96.400 310.400 ;
        RECT 106.800 309.600 107.600 310.400 ;
        RECT 92.400 305.600 93.200 306.400 ;
        RECT 100.400 305.600 101.200 306.400 ;
        RECT 108.400 307.600 109.200 308.400 ;
        RECT 98.800 303.600 99.600 304.400 ;
        RECT 102.000 303.600 102.800 304.400 ;
        RECT 114.800 303.600 115.600 304.400 ;
        RECT 124.400 305.600 125.200 306.400 ;
        RECT 132.400 309.600 133.200 310.400 ;
        RECT 130.800 307.600 131.600 308.400 ;
        RECT 126.000 303.600 126.800 304.400 ;
        RECT 129.200 303.600 130.000 304.400 ;
        RECT 143.600 309.600 144.400 310.400 ;
        RECT 142.000 307.600 142.800 308.400 ;
        RECT 134.000 305.600 134.800 306.400 ;
        RECT 145.200 307.600 146.000 308.400 ;
        RECT 146.800 307.600 147.600 308.400 ;
        RECT 150.000 303.600 150.800 304.400 ;
        RECT 161.200 305.600 162.000 306.400 ;
        RECT 159.600 303.600 160.400 304.400 ;
        RECT 172.400 305.600 173.200 306.400 ;
        RECT 170.800 303.600 171.600 304.400 ;
        RECT 194.800 312.400 195.600 313.200 ;
        RECT 198.000 311.000 198.800 311.800 ;
        RECT 199.600 313.600 200.400 314.400 ;
        RECT 214.000 312.400 214.800 313.200 ;
        RECT 217.200 311.000 218.000 311.800 ;
        RECT 198.000 306.200 198.800 307.000 ;
        RECT 178.800 303.600 179.600 304.400 ;
        RECT 180.400 303.600 181.200 304.400 ;
        RECT 217.200 306.200 218.000 307.000 ;
        RECT 231.600 311.600 232.400 312.400 ;
        RECT 231.600 309.600 232.400 310.400 ;
        RECT 239.600 307.600 240.400 308.400 ;
        RECT 252.400 309.600 253.200 310.400 ;
        RECT 273.200 317.600 274.000 318.400 ;
        RECT 263.600 309.600 264.400 310.400 ;
        RECT 249.200 305.600 250.000 306.400 ;
        RECT 271.600 309.600 272.400 310.400 ;
        RECT 287.600 312.400 288.400 313.200 ;
        RECT 290.800 311.000 291.600 311.800 ;
        RECT 311.600 312.400 312.400 313.200 ;
        RECT 314.800 311.000 315.600 311.800 ;
        RECT 290.800 306.200 291.600 307.000 ;
        RECT 314.800 306.200 315.600 307.000 ;
        RECT 297.200 303.600 298.000 304.400 ;
        RECT 335.600 309.600 336.400 310.400 ;
        RECT 351.600 317.600 352.400 318.400 ;
        RECT 342.000 309.600 342.800 310.400 ;
        RECT 348.400 309.600 349.200 310.400 ;
        RECT 330.800 307.600 331.600 308.400 ;
        RECT 337.200 307.600 338.000 308.400 ;
        RECT 343.600 307.600 344.400 308.400 ;
        RECT 356.400 311.800 357.200 312.600 ;
        RECT 367.800 311.800 368.600 312.600 ;
        RECT 378.800 317.600 379.600 318.400 ;
        RECT 356.400 306.200 357.200 307.000 ;
        RECT 369.000 309.800 369.800 310.600 ;
        RECT 364.400 307.600 365.200 308.400 ;
        RECT 361.200 306.400 362.000 307.200 ;
        RECT 367.800 306.200 368.600 307.000 ;
        RECT 375.600 307.600 376.400 308.400 ;
        RECT 377.200 307.600 378.000 308.400 ;
        RECT 388.400 309.600 389.200 310.400 ;
        RECT 391.600 309.600 392.400 310.400 ;
        RECT 404.400 313.600 405.200 314.400 ;
        RECT 382.000 305.600 382.800 306.400 ;
        RECT 388.400 305.600 389.200 306.400 ;
        RECT 396.400 305.600 397.200 306.400 ;
        RECT 401.200 307.600 402.000 308.400 ;
        RECT 418.800 312.400 419.600 313.200 ;
        RECT 422.000 311.000 422.800 311.800 ;
        RECT 394.800 303.600 395.600 304.400 ;
        RECT 402.800 305.600 403.600 306.400 ;
        RECT 422.000 306.200 422.800 307.000 ;
        RECT 438.000 309.600 438.800 310.400 ;
        RECT 441.200 307.600 442.000 308.400 ;
        RECT 450.800 307.600 451.600 308.400 ;
        RECT 458.800 309.600 459.600 310.400 ;
        RECT 460.400 307.600 461.200 308.400 ;
        RECT 433.200 303.600 434.000 304.400 ;
        RECT 466.800 311.800 467.600 312.600 ;
        RECT 476.400 317.600 477.200 318.400 ;
        RECT 466.800 306.200 467.600 307.000 ;
        RECT 462.000 303.600 462.800 304.400 ;
        RECT 474.800 307.600 475.600 308.400 ;
        RECT 471.600 306.400 472.400 307.200 ;
        RECT 497.200 317.600 498.000 318.400 ;
        RECT 478.000 305.600 478.800 306.400 ;
        RECT 479.600 306.200 480.400 307.000 ;
        RECT 511.600 314.400 512.400 315.200 ;
        RECT 514.800 315.000 515.600 315.800 ;
        RECT 510.000 312.400 510.800 313.200 ;
        RECT 529.200 311.600 530.000 312.400 ;
        RECT 500.400 305.600 501.200 306.400 ;
        RECT 516.400 305.600 517.200 306.400 ;
        RECT 510.000 304.200 510.800 305.000 ;
        RECT 511.600 304.200 512.400 305.000 ;
        RECT 513.200 304.200 514.000 305.000 ;
        RECT 514.800 304.200 515.600 305.000 ;
        RECT 518.000 304.200 518.800 305.000 ;
        RECT 521.200 304.200 522.000 305.000 ;
        RECT 522.800 304.200 523.600 305.000 ;
        RECT 524.400 304.200 525.200 305.000 ;
        RECT 535.600 311.600 536.400 312.400 ;
        RECT 562.800 313.600 563.600 314.400 ;
        RECT 543.600 305.600 544.400 306.400 ;
        RECT 545.200 306.200 546.000 307.000 ;
        RECT 566.000 307.600 566.800 308.400 ;
        RECT 564.400 306.200 565.200 307.000 ;
        RECT 582.000 303.600 582.800 304.400 ;
        RECT 2.800 289.600 3.600 290.400 ;
        RECT 17.200 291.600 18.000 292.400 ;
        RECT 23.600 291.600 24.400 292.400 ;
        RECT 46.000 297.600 46.800 298.400 ;
        RECT 4.400 283.600 5.200 284.400 ;
        RECT 10.800 283.600 11.600 284.400 ;
        RECT 17.200 283.600 18.000 284.400 ;
        RECT 39.600 293.600 40.400 294.400 ;
        RECT 44.400 293.600 45.200 294.400 ;
        RECT 41.200 291.600 42.000 292.400 ;
        RECT 49.200 291.600 50.000 292.400 ;
        RECT 36.400 283.600 37.200 284.400 ;
        RECT 55.600 289.600 56.400 290.400 ;
        RECT 90.800 297.600 91.600 298.400 ;
        RECT 70.000 289.600 70.800 290.400 ;
        RECT 60.400 285.600 61.200 286.400 ;
        RECT 74.800 291.600 75.600 292.400 ;
        RECT 84.400 293.600 85.200 294.400 ;
        RECT 86.000 291.600 86.800 292.400 ;
        RECT 81.200 283.600 82.000 284.400 ;
        RECT 98.800 294.800 99.600 295.600 ;
        RECT 103.600 297.600 104.400 298.400 ;
        RECT 102.000 293.600 102.800 294.400 ;
        RECT 90.800 289.600 91.600 290.400 ;
        RECT 130.800 295.600 131.600 296.400 ;
        RECT 156.400 297.600 157.200 298.400 ;
        RECT 119.600 293.600 120.400 294.400 ;
        RECT 121.200 291.600 122.000 292.400 ;
        RECT 116.400 283.600 117.200 284.400 ;
        RECT 132.400 289.600 133.200 290.400 ;
        RECT 143.600 289.600 144.400 290.400 ;
        RECT 135.600 283.600 136.400 284.400 ;
        RECT 148.400 291.600 149.200 292.400 ;
        RECT 190.000 294.800 190.800 295.600 ;
        RECT 183.600 293.600 184.400 294.400 ;
        RECT 174.000 291.600 174.800 292.400 ;
        RECT 175.600 291.600 176.400 292.400 ;
        RECT 169.200 283.600 170.000 284.400 ;
        RECT 185.200 289.600 186.000 290.400 ;
        RECT 202.800 292.200 203.600 293.000 ;
        RECT 210.800 291.800 211.600 292.600 ;
        RECT 215.600 290.200 216.400 291.000 ;
        RECT 198.000 285.600 198.800 286.400 ;
        RECT 244.400 297.600 245.200 298.400 ;
        RECT 231.600 293.600 232.400 294.400 ;
        RECT 226.800 290.200 227.600 291.000 ;
        RECT 252.400 294.800 253.200 295.600 ;
        RECT 255.600 293.600 256.400 294.400 ;
        RECT 262.000 292.200 262.800 293.000 ;
        RECT 270.000 291.800 270.800 292.600 ;
        RECT 281.200 292.200 282.000 293.000 ;
        RECT 289.200 291.800 290.000 292.600 ;
        RECT 274.800 290.200 275.600 291.000 ;
        RECT 257.200 283.600 258.000 284.400 ;
        RECT 294.000 290.200 294.800 291.000 ;
        RECT 276.400 283.600 277.200 284.400 ;
        RECT 311.600 294.800 312.400 295.600 ;
        RECT 302.000 289.600 302.800 290.400 ;
        RECT 303.600 289.600 304.400 290.400 ;
        RECT 340.400 293.600 341.200 294.400 ;
        RECT 334.000 292.200 334.800 293.000 ;
        RECT 342.000 291.800 342.800 292.600 ;
        RECT 367.600 297.600 368.400 298.400 ;
        RECT 353.200 292.200 354.000 293.000 ;
        RECT 361.200 291.800 362.000 292.600 ;
        RECT 346.800 290.200 347.600 291.000 ;
        RECT 329.200 283.600 330.000 284.400 ;
        RECT 372.400 292.200 373.200 293.000 ;
        RECT 393.200 294.800 394.000 295.600 ;
        RECT 380.400 291.800 381.200 292.600 ;
        RECT 366.000 290.200 366.800 291.000 ;
        RECT 348.400 283.600 349.200 284.400 ;
        RECT 385.200 290.200 386.000 291.000 ;
        RECT 414.000 297.600 414.800 298.400 ;
        RECT 418.800 292.200 419.600 293.000 ;
        RECT 439.600 294.800 440.400 295.600 ;
        RECT 442.800 293.600 443.600 294.400 ;
        RECT 457.200 293.600 458.000 294.400 ;
        RECT 466.800 293.600 467.600 294.400 ;
        RECT 431.600 290.200 432.400 291.000 ;
        RECT 457.200 289.600 458.000 290.400 ;
        RECT 470.000 291.800 470.800 292.600 ;
        RECT 463.600 289.600 464.400 290.400 ;
        RECT 465.200 290.200 466.000 291.000 ;
        RECT 490.800 294.800 491.600 295.600 ;
        RECT 494.000 293.600 494.800 294.400 ;
        RECT 508.400 293.600 509.200 294.400 ;
        RECT 511.600 293.600 512.400 294.400 ;
        RECT 516.400 293.600 517.200 294.400 ;
        RECT 514.800 291.800 515.600 292.600 ;
        RECT 482.800 287.600 483.600 288.400 ;
        RECT 510.000 290.200 510.800 291.000 ;
        RECT 524.400 287.600 525.200 288.400 ;
        RECT 527.600 287.600 528.400 288.400 ;
        RECT 551.600 295.600 552.400 296.400 ;
        RECT 553.200 294.200 554.000 295.000 ;
        RECT 564.400 291.600 565.200 292.400 ;
        RECT 529.200 283.600 530.000 284.400 ;
        RECT 546.800 286.800 547.600 287.600 ;
        RECT 550.000 286.200 550.800 287.000 ;
        RECT 545.200 284.200 546.000 285.000 ;
        RECT 546.800 284.200 547.600 285.000 ;
        RECT 548.400 284.200 549.200 285.000 ;
        RECT 553.200 286.200 554.000 287.000 ;
        RECT 556.400 286.200 557.200 287.000 ;
        RECT 558.000 284.200 558.800 285.000 ;
        RECT 559.600 284.200 560.400 285.000 ;
        RECT 9.200 271.800 10.000 272.600 ;
        RECT 2.800 263.600 3.600 264.400 ;
        RECT 9.200 266.200 10.000 267.000 ;
        RECT 17.200 267.600 18.000 268.400 ;
        RECT 14.000 266.400 14.800 267.200 ;
        RECT 12.400 263.600 13.200 264.400 ;
        RECT 18.800 265.600 19.600 266.400 ;
        RECT 30.000 277.600 30.800 278.400 ;
        RECT 22.000 263.600 22.800 264.400 ;
        RECT 28.400 265.600 29.200 266.400 ;
        RECT 34.800 269.600 35.600 270.400 ;
        RECT 36.400 267.600 37.200 268.400 ;
        RECT 31.600 263.600 32.400 264.400 ;
        RECT 57.200 277.600 58.000 278.400 ;
        RECT 39.600 263.600 40.400 264.400 ;
        RECT 46.000 265.600 46.800 266.400 ;
        RECT 55.600 265.600 56.400 266.400 ;
        RECT 50.800 263.600 51.600 264.400 ;
        RECT 60.400 271.800 61.200 272.600 ;
        RECT 60.400 266.200 61.200 267.000 ;
        RECT 71.600 269.600 72.400 270.400 ;
        RECT 68.400 267.600 69.200 268.400 ;
        RECT 87.400 271.800 88.200 272.600 ;
        RECT 82.800 269.600 83.600 270.400 ;
        RECT 65.200 266.400 66.000 267.200 ;
        RECT 84.400 267.600 85.200 268.400 ;
        RECT 87.400 266.200 88.200 267.000 ;
        RECT 79.600 263.600 80.400 264.400 ;
        RECT 95.600 267.600 96.400 268.400 ;
        RECT 92.400 263.600 93.200 264.400 ;
        RECT 100.400 265.600 101.200 266.400 ;
        RECT 105.200 265.600 106.000 266.400 ;
        RECT 106.800 265.600 107.600 266.400 ;
        RECT 126.000 277.600 126.800 278.400 ;
        RECT 121.200 269.600 122.000 270.400 ;
        RECT 124.400 267.600 125.200 268.400 ;
        RECT 118.000 263.600 118.800 264.400 ;
        RECT 130.800 269.600 131.600 270.400 ;
        RECT 132.400 267.600 133.200 268.400 ;
        RECT 134.000 267.600 134.800 268.400 ;
        RECT 153.200 271.600 154.000 272.400 ;
        RECT 145.200 269.600 146.000 270.400 ;
        RECT 146.800 269.600 147.600 270.400 ;
        RECT 154.800 267.600 155.600 268.400 ;
        RECT 127.600 263.600 128.400 264.400 ;
        RECT 161.200 269.600 162.000 270.400 ;
        RECT 169.200 269.600 170.000 270.400 ;
        RECT 158.000 265.600 158.800 266.400 ;
        RECT 166.000 267.600 166.800 268.400 ;
        RECT 178.800 273.600 179.600 274.400 ;
        RECT 177.200 267.600 178.000 268.400 ;
        RECT 193.200 272.400 194.000 273.200 ;
        RECT 196.400 271.000 197.200 271.800 ;
        RECT 212.400 272.400 213.200 273.200 ;
        RECT 218.600 271.800 219.400 272.600 ;
        RECT 215.600 271.000 216.400 271.800 ;
        RECT 196.400 266.200 197.200 267.000 ;
        RECT 215.600 266.200 216.400 267.000 ;
        RECT 198.000 263.600 198.800 264.400 ;
        RECT 218.600 266.200 219.400 267.000 ;
        RECT 242.800 269.600 243.600 270.400 ;
        RECT 249.200 269.600 250.000 270.400 ;
        RECT 234.800 265.600 235.600 266.400 ;
        RECT 244.400 267.600 245.200 268.400 ;
        RECT 250.800 267.600 251.600 268.400 ;
        RECT 255.600 268.000 256.400 268.800 ;
        RECT 265.200 269.600 266.000 270.400 ;
        RECT 271.400 271.800 272.200 272.600 ;
        RECT 262.000 267.600 262.800 268.400 ;
        RECT 271.400 266.200 272.200 267.000 ;
        RECT 285.800 271.800 286.600 272.600 ;
        RECT 279.600 267.600 280.400 268.400 ;
        RECT 281.200 267.600 282.000 268.400 ;
        RECT 282.800 265.600 283.600 266.400 ;
        RECT 285.800 266.200 286.600 267.000 ;
        RECT 294.000 267.600 294.800 268.400 ;
        RECT 316.400 269.600 317.200 270.400 ;
        RECT 321.200 269.600 322.000 270.400 ;
        RECT 324.400 269.600 325.200 270.400 ;
        RECT 305.200 265.600 306.000 266.400 ;
        RECT 311.600 265.600 312.400 266.400 ;
        RECT 318.000 267.600 318.800 268.400 ;
        RECT 326.000 267.600 326.800 268.400 ;
        RECT 321.200 265.600 322.000 266.400 ;
        RECT 329.200 265.600 330.000 266.400 ;
        RECT 334.000 267.600 334.800 268.400 ;
        RECT 338.800 267.600 339.600 268.400 ;
        RECT 356.400 272.400 357.200 273.200 ;
        RECT 362.600 271.800 363.400 272.600 ;
        RECT 359.600 271.000 360.400 271.800 ;
        RECT 332.400 263.600 333.200 264.400 ;
        RECT 340.400 265.600 341.200 266.400 ;
        RECT 359.600 266.200 360.400 267.000 ;
        RECT 342.000 263.600 342.800 264.400 ;
        RECT 362.600 266.200 363.400 267.000 ;
        RECT 386.800 277.600 387.600 278.400 ;
        RECT 385.200 273.600 386.000 274.400 ;
        RECT 382.000 271.600 382.800 272.400 ;
        RECT 370.800 267.600 371.600 268.400 ;
        RECT 377.200 267.600 378.000 268.400 ;
        RECT 394.800 271.600 395.600 272.400 ;
        RECT 380.400 265.600 381.200 266.400 ;
        RECT 391.600 263.600 392.400 264.400 ;
        RECT 396.400 265.600 397.200 266.400 ;
        RECT 409.200 277.600 410.000 278.400 ;
        RECT 402.800 265.600 403.600 266.400 ;
        RECT 409.200 263.600 410.000 264.400 ;
        RECT 410.800 277.600 411.600 278.400 ;
        RECT 428.400 272.400 429.200 273.200 ;
        RECT 431.600 271.000 432.400 271.800 ;
        RECT 455.600 277.600 456.400 278.400 ;
        RECT 451.000 271.800 451.800 272.600 ;
        RECT 462.000 277.600 462.800 278.400 ;
        RECT 452.200 269.800 453.000 270.600 ;
        RECT 412.400 265.600 413.200 266.400 ;
        RECT 410.800 263.600 411.600 264.400 ;
        RECT 431.600 266.200 432.400 267.000 ;
        RECT 436.400 265.600 437.200 266.400 ;
        RECT 442.800 267.600 443.600 268.400 ;
        RECT 451.000 266.200 451.800 267.000 ;
        RECT 434.800 263.600 435.600 264.400 ;
        RECT 458.800 267.600 459.600 268.400 ;
        RECT 460.400 267.600 461.200 268.400 ;
        RECT 482.800 273.600 483.600 274.400 ;
        RECT 466.800 267.600 467.600 268.400 ;
        RECT 465.200 266.200 466.000 267.000 ;
        RECT 521.200 273.600 522.000 274.400 ;
        RECT 484.400 266.200 485.200 267.000 ;
        RECT 510.000 269.600 510.800 270.400 ;
        RECT 502.000 263.600 502.800 264.400 ;
        RECT 503.600 266.200 504.400 267.000 ;
        RECT 559.600 273.600 560.400 274.400 ;
        RECT 524.400 267.600 525.200 268.400 ;
        RECT 522.800 266.200 523.600 267.000 ;
        RECT 534.000 267.600 534.800 268.400 ;
        RECT 578.800 273.600 579.600 274.400 ;
        RECT 543.600 267.600 544.400 268.400 ;
        RECT 540.400 263.600 541.200 264.400 ;
        RECT 542.000 266.200 542.800 267.000 ;
        RECT 562.800 267.600 563.600 268.400 ;
        RECT 561.200 266.200 562.000 267.000 ;
        RECT 580.400 269.600 581.200 270.400 ;
        RECT 6.000 249.600 6.800 250.400 ;
        RECT 9.200 243.600 10.000 244.400 ;
        RECT 20.400 253.600 21.200 254.400 ;
        RECT 41.200 249.600 42.000 250.400 ;
        RECT 30.000 243.600 30.800 244.400 ;
        RECT 38.000 243.600 38.800 244.400 ;
        RECT 46.000 251.600 46.800 252.400 ;
        RECT 57.200 254.800 58.000 255.600 ;
        RECT 65.200 254.800 66.000 255.600 ;
        RECT 60.400 253.600 61.200 254.400 ;
        RECT 76.400 257.600 77.200 258.400 ;
        RECT 74.800 253.600 75.600 254.400 ;
        RECT 66.800 243.600 67.600 244.400 ;
        RECT 87.600 253.600 88.400 254.400 ;
        RECT 118.000 253.600 118.800 254.400 ;
        RECT 130.800 254.800 131.600 255.600 ;
        RECT 111.600 251.600 112.400 252.400 ;
        RECT 97.200 243.600 98.000 244.400 ;
        RECT 146.800 254.800 147.600 255.600 ;
        RECT 137.200 253.600 138.000 254.400 ;
        RECT 158.000 257.600 158.800 258.400 ;
        RECT 170.800 257.600 171.600 258.400 ;
        RECT 153.200 253.600 154.000 254.400 ;
        RECT 162.800 251.600 163.600 252.400 ;
        RECT 164.400 249.600 165.200 250.400 ;
        RECT 177.200 251.600 178.000 252.400 ;
        RECT 185.200 243.600 186.000 244.400 ;
        RECT 199.600 257.600 200.400 258.400 ;
        RECT 218.800 257.600 219.600 258.400 ;
        RECT 204.400 252.200 205.200 253.000 ;
        RECT 212.400 251.800 213.200 252.600 ;
        RECT 223.600 252.200 224.400 253.000 ;
        RECT 217.200 250.200 218.000 251.000 ;
        RECT 236.400 250.200 237.200 251.000 ;
        RECT 262.000 257.600 262.800 258.400 ;
        RECT 258.800 253.600 259.600 254.400 ;
        RECT 247.600 252.200 248.400 253.000 ;
        RECT 238.000 243.600 238.800 244.400 ;
        RECT 255.600 251.800 256.400 252.600 ;
        RECT 281.200 253.600 282.000 254.400 ;
        RECT 266.800 252.200 267.600 253.000 ;
        RECT 274.800 251.800 275.600 252.600 ;
        RECT 260.400 250.200 261.200 251.000 ;
        RECT 242.800 243.600 243.600 244.400 ;
        RECT 279.600 250.200 280.400 251.000 ;
        RECT 313.200 254.800 314.000 255.600 ;
        RECT 295.600 252.200 296.400 253.000 ;
        RECT 303.600 251.800 304.400 252.600 ;
        RECT 319.600 253.600 320.400 254.400 ;
        RECT 308.400 250.200 309.200 251.000 ;
        RECT 343.600 251.600 344.400 252.400 ;
        RECT 345.200 249.600 346.000 250.400 ;
        RECT 353.200 251.600 354.000 252.400 ;
        RECT 367.600 257.600 368.400 258.400 ;
        RECT 364.400 249.600 365.200 250.400 ;
        RECT 383.600 253.600 384.400 254.400 ;
        RECT 388.400 253.600 389.200 254.400 ;
        RECT 372.400 252.200 373.200 253.000 ;
        RECT 380.400 251.800 381.200 252.600 ;
        RECT 393.200 251.600 394.000 252.400 ;
        RECT 385.200 250.200 386.000 251.000 ;
        RECT 399.600 257.600 400.400 258.400 ;
        RECT 398.000 251.600 398.800 252.400 ;
        RECT 418.800 257.600 419.600 258.400 ;
        RECT 415.600 253.600 416.400 254.400 ;
        RECT 404.400 252.200 405.200 253.000 ;
        RECT 430.000 253.600 430.800 254.400 ;
        RECT 441.200 257.600 442.000 258.400 ;
        RECT 439.600 253.600 440.400 254.400 ;
        RECT 423.600 252.200 424.400 253.000 ;
        RECT 417.200 250.200 418.000 251.000 ;
        RECT 431.600 251.800 432.400 252.600 ;
        RECT 463.600 257.600 464.400 258.400 ;
        RECT 462.000 253.600 462.800 254.400 ;
        RECT 436.400 250.200 437.200 251.000 ;
        RECT 452.400 251.600 453.200 252.400 ;
        RECT 455.600 251.600 456.400 252.400 ;
        RECT 466.800 251.600 467.600 252.400 ;
        RECT 452.400 245.600 453.200 246.400 ;
        RECT 490.800 257.600 491.600 258.400 ;
        RECT 478.000 249.600 478.800 250.400 ;
        RECT 486.000 249.600 486.800 250.400 ;
        RECT 489.200 249.600 490.000 250.400 ;
        RECT 510.000 257.600 510.800 258.400 ;
        RECT 510.000 254.800 510.800 255.600 ;
        RECT 521.200 257.600 522.000 258.400 ;
        RECT 497.200 251.600 498.000 252.400 ;
        RECT 498.800 251.600 499.600 252.400 ;
        RECT 513.200 253.600 514.000 254.400 ;
        RECT 532.400 257.600 533.200 258.400 ;
        RECT 524.400 253.600 525.200 254.400 ;
        RECT 532.400 254.800 533.200 255.600 ;
        RECT 535.600 253.600 536.400 254.400 ;
        RECT 543.600 253.600 544.400 254.400 ;
        RECT 542.000 251.800 542.800 252.600 ;
        RECT 537.200 250.200 538.000 251.000 ;
        RECT 562.800 253.600 563.600 254.400 ;
        RECT 566.000 251.800 566.800 252.600 ;
        RECT 554.800 247.600 555.600 248.400 ;
        RECT 561.200 250.200 562.000 251.000 ;
        RECT 578.800 247.600 579.600 248.400 ;
        RECT 15.600 232.400 16.400 233.200 ;
        RECT 22.000 231.800 22.800 232.600 ;
        RECT 33.200 231.800 34.000 232.600 ;
        RECT 18.800 231.000 19.600 231.800 ;
        RECT 18.800 226.200 19.600 227.000 ;
        RECT 1.200 223.600 2.000 224.400 ;
        RECT 22.000 226.200 22.800 227.000 ;
        RECT 30.000 227.600 30.800 228.400 ;
        RECT 26.800 226.400 27.600 227.200 ;
        RECT 25.200 223.600 26.000 224.400 ;
        RECT 33.200 226.200 34.000 227.000 ;
        RECT 41.200 227.600 42.000 228.400 ;
        RECT 38.000 226.400 38.800 227.200 ;
        RECT 57.200 232.400 58.000 233.200 ;
        RECT 60.400 231.000 61.200 231.800 ;
        RECT 82.600 231.800 83.400 232.600 ;
        RECT 55.600 225.600 56.400 226.400 ;
        RECT 42.800 223.600 43.600 224.400 ;
        RECT 60.400 226.200 61.200 227.000 ;
        RECT 62.000 226.200 62.800 227.000 ;
        RECT 79.600 223.600 80.400 224.400 ;
        RECT 82.600 226.200 83.400 227.000 ;
        RECT 90.800 227.600 91.600 228.400 ;
        RECT 95.600 227.600 96.400 228.400 ;
        RECT 111.600 232.400 112.400 233.200 ;
        RECT 114.800 231.000 115.600 231.800 ;
        RECT 130.800 232.400 131.600 233.200 ;
        RECT 141.800 231.800 142.600 232.600 ;
        RECT 134.000 231.000 134.800 231.800 ;
        RECT 153.200 229.600 154.000 230.400 ;
        RECT 114.800 226.200 115.600 227.000 ;
        RECT 97.200 223.600 98.000 224.400 ;
        RECT 134.000 226.200 134.800 227.000 ;
        RECT 116.400 223.600 117.200 224.400 ;
        RECT 141.800 226.200 142.600 227.000 ;
        RECT 159.600 229.600 160.400 230.400 ;
        RECT 150.000 227.600 150.800 228.400 ;
        RECT 178.800 232.400 179.600 233.200 ;
        RECT 182.000 231.000 182.800 231.800 ;
        RECT 196.400 229.600 197.200 230.400 ;
        RECT 162.800 223.600 163.600 224.400 ;
        RECT 182.000 226.200 182.800 227.000 ;
        RECT 164.400 223.600 165.200 224.400 ;
        RECT 212.400 232.400 213.200 233.200 ;
        RECT 215.600 231.000 216.400 231.800 ;
        RECT 231.600 232.400 232.400 233.200 ;
        RECT 234.800 231.000 235.600 231.800 ;
        RECT 215.600 226.200 216.400 227.000 ;
        RECT 198.000 223.600 198.800 224.400 ;
        RECT 234.800 226.200 235.600 227.000 ;
        RECT 217.200 223.600 218.000 224.400 ;
        RECT 236.400 225.600 237.200 226.400 ;
        RECT 238.000 223.600 238.800 224.400 ;
        RECT 239.600 233.600 240.400 234.400 ;
        RECT 258.800 233.600 259.600 234.400 ;
        RECT 242.800 229.600 243.600 230.400 ;
        RECT 246.000 227.600 246.800 228.400 ;
        RECT 244.400 226.200 245.200 227.000 ;
        RECT 270.000 229.600 270.800 230.400 ;
        RECT 265.200 227.600 266.000 228.400 ;
        RECT 262.000 223.600 262.800 224.400 ;
        RECT 263.600 226.200 264.400 227.000 ;
        RECT 282.800 225.600 283.600 226.400 ;
        RECT 281.200 223.600 282.000 224.400 ;
        RECT 297.200 233.600 298.000 234.400 ;
        RECT 314.800 229.600 315.600 230.400 ;
        RECT 310.000 227.600 310.800 228.400 ;
        RECT 302.000 225.600 302.800 226.400 ;
        RECT 308.400 226.200 309.200 227.000 ;
        RECT 326.000 223.600 326.800 224.400 ;
        RECT 332.400 225.600 333.200 226.400 ;
        RECT 329.200 223.600 330.000 224.400 ;
        RECT 358.000 233.600 358.800 234.400 ;
        RECT 340.400 226.200 341.200 227.000 ;
        RECT 338.800 223.600 339.600 224.400 ;
        RECT 359.600 229.600 360.400 230.400 ;
        RECT 362.800 227.600 363.600 228.400 ;
        RECT 378.800 232.400 379.600 233.200 ;
        RECT 382.000 231.000 382.800 231.800 ;
        RECT 401.200 235.600 402.000 236.400 ;
        RECT 382.000 226.200 382.800 227.000 ;
        RECT 364.400 223.600 365.200 224.400 ;
        RECT 383.600 226.200 384.400 227.000 ;
        RECT 404.400 227.600 405.200 228.400 ;
        RECT 402.800 226.200 403.600 227.000 ;
        RECT 433.200 237.600 434.000 238.400 ;
        RECT 439.600 237.600 440.400 238.400 ;
        RECT 450.800 237.600 451.600 238.400 ;
        RECT 441.200 233.600 442.000 234.400 ;
        RECT 438.000 231.600 438.800 232.400 ;
        RECT 428.400 223.600 429.200 224.400 ;
        RECT 434.800 225.600 435.600 226.400 ;
        RECT 436.400 225.600 437.200 226.400 ;
        RECT 444.400 231.600 445.200 232.400 ;
        RECT 442.800 229.600 443.600 230.400 ;
        RECT 455.600 233.600 456.400 234.400 ;
        RECT 457.200 225.600 458.000 226.400 ;
        RECT 465.200 231.600 466.000 232.400 ;
        RECT 463.600 227.600 464.400 228.400 ;
        RECT 470.000 229.600 470.800 230.400 ;
        RECT 473.200 229.600 474.000 230.400 ;
        RECT 474.800 227.600 475.600 228.400 ;
        RECT 460.400 223.600 461.200 224.400 ;
        RECT 470.000 223.600 470.800 224.400 ;
        RECT 476.400 225.600 477.200 226.400 ;
        RECT 486.000 233.600 486.800 234.400 ;
        RECT 481.200 231.800 482.000 232.600 ;
        RECT 508.400 233.600 509.200 234.400 ;
        RECT 478.000 223.600 478.800 224.400 ;
        RECT 481.200 226.200 482.000 227.000 ;
        RECT 527.600 233.600 528.400 234.400 ;
        RECT 489.200 227.600 490.000 228.400 ;
        RECT 492.400 227.600 493.200 228.400 ;
        RECT 486.000 226.400 486.800 227.200 ;
        RECT 490.800 226.200 491.600 227.000 ;
        RECT 511.600 227.600 512.400 228.400 ;
        RECT 510.000 226.200 510.800 227.000 ;
        RECT 551.600 233.600 552.400 234.400 ;
        RECT 529.200 229.600 530.000 230.400 ;
        RECT 570.800 233.600 571.600 234.400 ;
        RECT 534.000 226.200 534.800 227.000 ;
        RECT 554.800 227.600 555.600 228.400 ;
        RECT 553.200 226.200 554.000 227.000 ;
        RECT 564.400 227.600 565.200 228.400 ;
        RECT 572.400 229.600 573.200 230.400 ;
        RECT 577.200 229.600 578.000 230.400 ;
        RECT 6.000 211.800 6.800 212.600 ;
        RECT 1.200 210.200 2.000 211.000 ;
        RECT 18.800 203.600 19.600 204.400 ;
        RECT 20.400 210.200 21.200 211.000 ;
        RECT 38.000 203.600 38.800 204.400 ;
        RECT 55.600 213.600 56.400 214.400 ;
        RECT 44.400 212.200 45.200 213.000 ;
        RECT 52.400 211.800 53.200 212.600 ;
        RECT 57.200 210.200 58.000 211.000 ;
        RECT 39.600 203.600 40.400 204.400 ;
        RECT 58.800 210.200 59.600 211.000 ;
        RECT 76.400 203.600 77.200 204.400 ;
        RECT 94.000 213.600 94.800 214.400 ;
        RECT 97.200 213.600 98.000 214.400 ;
        RECT 82.800 212.200 83.600 213.000 ;
        RECT 90.800 211.800 91.600 212.600 ;
        RECT 95.600 210.200 96.400 211.000 ;
        RECT 78.000 203.600 78.800 204.400 ;
        RECT 127.600 213.600 128.400 214.400 ;
        RECT 116.400 212.200 117.200 213.000 ;
        RECT 124.400 211.800 125.200 212.600 ;
        RECT 129.200 210.200 130.000 211.000 ;
        RECT 111.600 203.600 112.400 204.400 ;
        RECT 135.600 210.200 136.400 211.000 ;
        RECT 153.200 203.600 154.000 204.400 ;
        RECT 154.800 210.200 155.600 211.000 ;
        RECT 172.400 203.600 173.200 204.400 ;
        RECT 220.400 217.600 221.200 218.400 ;
        RECT 180.400 203.600 181.200 204.400 ;
        RECT 186.800 209.600 187.600 210.400 ;
        RECT 191.600 211.600 192.400 212.400 ;
        RECT 204.400 213.600 205.200 214.400 ;
        RECT 207.600 211.800 208.400 212.600 ;
        RECT 201.200 209.600 202.000 210.400 ;
        RECT 202.800 210.200 203.600 211.000 ;
        RECT 271.600 217.600 272.400 218.400 ;
        RECT 222.000 211.600 222.800 212.400 ;
        RECT 217.200 207.600 218.000 208.400 ;
        RECT 246.000 213.600 246.800 214.400 ;
        RECT 233.200 207.600 234.000 208.400 ;
        RECT 239.600 209.600 240.400 210.400 ;
        RECT 246.000 209.600 246.800 210.400 ;
        RECT 258.800 211.800 259.600 212.600 ;
        RECT 252.400 209.600 253.200 210.400 ;
        RECT 254.000 210.200 254.800 211.000 ;
        RECT 284.400 217.600 285.200 218.400 ;
        RECT 279.600 211.600 280.400 212.400 ;
        RECT 284.400 209.600 285.200 210.400 ;
        RECT 298.800 217.600 299.600 218.400 ;
        RECT 310.000 213.600 310.800 214.400 ;
        RECT 318.000 213.600 318.800 214.400 ;
        RECT 303.600 212.200 304.400 213.000 ;
        RECT 311.600 211.800 312.400 212.600 ;
        RECT 316.400 210.200 317.200 211.000 ;
        RECT 342.000 215.600 342.800 216.400 ;
        RECT 327.600 212.200 328.400 213.000 ;
        RECT 335.600 211.800 336.400 212.600 ;
        RECT 364.400 217.600 365.200 218.400 ;
        RECT 340.400 210.200 341.200 211.000 ;
        RECT 322.800 207.600 323.600 208.400 ;
        RECT 348.400 213.600 349.200 214.400 ;
        RECT 351.600 211.800 352.400 212.600 ;
        RECT 346.800 210.200 347.600 211.000 ;
        RECT 388.400 217.600 389.200 218.400 ;
        RECT 374.000 209.600 374.800 210.400 ;
        RECT 380.400 209.600 381.200 210.400 ;
        RECT 407.600 217.600 408.400 218.400 ;
        RECT 409.200 214.800 410.000 215.600 ;
        RECT 412.400 213.600 413.200 214.400 ;
        RECT 415.600 213.600 416.400 214.400 ;
        RECT 418.800 211.800 419.600 212.600 ;
        RECT 399.600 209.600 400.400 210.400 ;
        RECT 414.000 210.200 414.800 211.000 ;
        RECT 436.400 213.600 437.200 214.400 ;
        RECT 439.600 211.600 440.400 212.400 ;
        RECT 431.600 207.600 432.400 208.400 ;
        RECT 486.000 217.600 486.800 218.400 ;
        RECT 452.400 209.600 453.200 210.400 ;
        RECT 463.600 209.600 464.400 210.400 ;
        RECT 465.200 209.600 466.000 210.400 ;
        RECT 474.800 209.600 475.600 210.400 ;
        RECT 481.200 209.600 482.000 210.400 ;
        RECT 495.600 217.600 496.400 218.400 ;
        RECT 510.000 217.600 510.800 218.400 ;
        RECT 489.200 213.600 490.000 214.400 ;
        RECT 497.200 213.600 498.000 214.400 ;
        RECT 506.800 214.800 507.600 215.600 ;
        RECT 500.400 213.600 501.200 214.400 ;
        RECT 486.000 209.600 486.800 210.400 ;
        RECT 521.200 217.600 522.000 218.400 ;
        RECT 513.200 213.600 514.000 214.400 ;
        RECT 521.200 214.800 522.000 215.600 ;
        RECT 542.000 217.600 542.800 218.400 ;
        RECT 524.400 213.600 525.200 214.400 ;
        RECT 527.600 213.600 528.400 214.400 ;
        RECT 502.000 209.600 502.800 210.400 ;
        RECT 534.000 209.600 534.800 210.400 ;
        RECT 548.400 211.800 549.200 212.600 ;
        RECT 542.000 209.600 542.800 210.400 ;
        RECT 543.600 210.200 544.400 211.000 ;
        RECT 564.400 213.600 565.200 214.400 ;
        RECT 567.600 213.600 568.400 214.400 ;
        RECT 561.200 207.600 562.000 208.400 ;
        RECT 562.800 210.200 563.600 211.000 ;
        RECT 580.400 207.600 581.200 208.400 ;
        RECT 1.200 186.200 2.000 187.000 ;
        RECT 18.800 183.600 19.600 184.400 ;
        RECT 20.400 186.200 21.200 187.000 ;
        RECT 42.800 187.600 43.600 188.400 ;
        RECT 44.400 185.600 45.200 186.400 ;
        RECT 38.000 183.600 38.800 184.400 ;
        RECT 50.800 185.600 51.600 186.400 ;
        RECT 68.400 189.600 69.200 190.400 ;
        RECT 63.600 187.600 64.400 188.400 ;
        RECT 70.000 187.600 70.800 188.400 ;
        RECT 52.400 183.600 53.200 184.400 ;
        RECT 57.200 183.600 58.000 184.400 ;
        RECT 62.000 183.600 62.800 184.400 ;
        RECT 78.000 185.600 78.800 186.400 ;
        RECT 76.400 183.600 77.200 184.400 ;
        RECT 86.000 191.600 86.800 192.400 ;
        RECT 87.600 185.600 88.400 186.400 ;
        RECT 92.400 187.600 93.200 188.400 ;
        RECT 94.000 185.600 94.800 186.400 ;
        RECT 108.400 187.600 109.200 188.400 ;
        RECT 113.200 187.600 114.000 188.400 ;
        RECT 102.000 183.600 102.800 184.400 ;
        RECT 111.600 183.600 112.400 184.400 ;
        RECT 129.200 189.600 130.000 190.400 ;
        RECT 121.200 187.600 122.000 188.400 ;
        RECT 122.800 186.200 123.600 187.000 ;
        RECT 119.600 183.600 120.400 184.400 ;
        RECT 146.800 186.200 147.600 187.000 ;
        RECT 164.400 183.600 165.200 184.400 ;
        RECT 166.000 186.200 166.800 187.000 ;
        RECT 185.200 185.600 186.000 186.400 ;
        RECT 183.600 183.600 184.400 184.400 ;
        RECT 191.600 191.600 192.400 192.400 ;
        RECT 191.600 189.600 192.400 190.400 ;
        RECT 193.200 187.600 194.000 188.400 ;
        RECT 202.800 193.600 203.600 194.400 ;
        RECT 202.800 189.600 203.600 190.400 ;
        RECT 198.000 187.600 198.800 188.400 ;
        RECT 204.400 187.600 205.200 188.400 ;
        RECT 215.600 191.800 216.400 192.600 ;
        RECT 186.800 183.600 187.600 184.400 ;
        RECT 196.400 183.600 197.200 184.400 ;
        RECT 207.600 183.600 208.400 184.400 ;
        RECT 212.400 185.600 213.200 186.400 ;
        RECT 215.600 186.200 216.400 187.000 ;
        RECT 223.600 187.600 224.400 188.400 ;
        RECT 226.800 187.600 227.600 188.400 ;
        RECT 220.400 186.400 221.200 187.200 ;
        RECT 225.200 186.200 226.000 187.000 ;
        RECT 247.600 189.600 248.400 190.400 ;
        RECT 265.200 197.600 266.000 198.400 ;
        RECT 260.200 191.800 261.000 192.600 ;
        RECT 246.000 187.600 246.800 188.400 ;
        RECT 249.200 187.600 250.000 188.400 ;
        RECT 242.800 183.600 243.600 184.400 ;
        RECT 250.800 185.600 251.600 186.400 ;
        RECT 257.200 185.600 258.000 186.400 ;
        RECT 260.200 186.200 261.000 187.000 ;
        RECT 268.400 187.600 269.200 188.400 ;
        RECT 276.400 187.600 277.200 188.400 ;
        RECT 274.800 186.200 275.600 187.000 ;
        RECT 273.200 183.600 274.000 184.400 ;
        RECT 298.800 187.600 299.600 188.400 ;
        RECT 314.800 189.600 315.600 190.400 ;
        RECT 308.400 187.600 309.200 188.400 ;
        RECT 292.400 183.600 293.200 184.400 ;
        RECT 310.000 187.600 310.800 188.400 ;
        RECT 313.200 187.600 314.000 188.400 ;
        RECT 318.000 187.600 318.800 188.400 ;
        RECT 324.200 191.800 325.000 192.600 ;
        RECT 335.600 189.600 336.400 190.400 ;
        RECT 324.200 186.200 325.000 187.000 ;
        RECT 321.200 183.600 322.000 184.400 ;
        RECT 351.600 197.600 352.400 198.400 ;
        RECT 346.800 191.800 347.600 192.600 ;
        RECT 374.000 197.600 374.800 198.400 ;
        RECT 332.400 187.600 333.200 188.400 ;
        RECT 342.000 187.600 342.800 188.400 ;
        RECT 346.800 186.200 347.600 187.000 ;
        RECT 380.400 197.600 381.200 198.400 ;
        RECT 354.800 187.600 355.600 188.400 ;
        RECT 358.000 187.600 358.800 188.400 ;
        RECT 351.600 186.400 352.400 187.200 ;
        RECT 356.400 186.200 357.200 187.000 ;
        RECT 377.200 189.600 378.000 190.400 ;
        RECT 402.800 197.600 403.600 198.400 ;
        RECT 388.400 189.600 389.200 190.400 ;
        RECT 374.000 183.600 374.800 184.400 ;
        RECT 390.000 187.600 390.800 188.400 ;
        RECT 391.600 185.600 392.400 186.400 ;
        RECT 399.600 185.600 400.400 186.400 ;
        RECT 401.200 185.600 402.000 186.400 ;
        RECT 409.200 197.600 410.000 198.400 ;
        RECT 404.400 185.600 405.200 186.400 ;
        RECT 423.600 192.400 424.400 193.200 ;
        RECT 426.800 191.000 427.600 191.800 ;
        RECT 471.600 197.600 472.400 198.400 ;
        RECT 466.600 191.800 467.400 192.600 ;
        RECT 426.800 186.200 427.600 187.000 ;
        RECT 428.400 186.200 429.200 187.000 ;
        RECT 433.200 185.600 434.000 186.400 ;
        RECT 462.000 189.600 462.800 190.400 ;
        RECT 478.000 189.600 478.800 190.400 ;
        RECT 460.400 187.600 461.200 188.400 ;
        RECT 463.600 187.600 464.400 188.400 ;
        RECT 466.600 186.200 467.400 187.000 ;
        RECT 474.800 187.600 475.600 188.400 ;
        RECT 481.200 187.600 482.000 188.400 ;
        RECT 487.600 189.600 488.400 190.400 ;
        RECT 497.200 197.600 498.000 198.400 ;
        RECT 505.200 197.600 506.000 198.400 ;
        RECT 500.400 191.800 501.200 192.600 ;
        RECT 511.600 191.600 512.400 192.400 ;
        RECT 484.400 185.600 485.200 186.400 ;
        RECT 500.400 186.200 501.200 187.000 ;
        RECT 508.400 187.600 509.200 188.400 ;
        RECT 505.200 186.400 506.000 187.200 ;
        RECT 510.000 185.600 510.800 186.400 ;
        RECT 513.200 185.600 514.000 186.400 ;
        RECT 524.400 197.600 525.200 198.400 ;
        RECT 534.000 197.600 534.800 198.400 ;
        RECT 521.200 187.600 522.000 188.400 ;
        RECT 524.400 185.600 525.200 186.400 ;
        RECT 530.800 187.600 531.600 188.400 ;
        RECT 514.800 183.600 515.600 184.400 ;
        RECT 532.400 185.600 533.200 186.400 ;
        RECT 537.200 197.600 538.000 198.400 ;
        RECT 535.600 187.600 536.400 188.400 ;
        RECT 545.200 189.600 546.000 190.400 ;
        RECT 556.400 191.800 557.200 192.600 ;
        RECT 542.000 187.600 542.800 188.400 ;
        RECT 548.400 187.600 549.200 188.400 ;
        RECT 540.400 183.600 541.200 184.400 ;
        RECT 553.200 185.600 554.000 186.400 ;
        RECT 556.400 186.200 557.200 187.000 ;
        RECT 564.400 187.600 565.200 188.400 ;
        RECT 567.600 187.600 568.400 188.400 ;
        RECT 561.200 186.400 562.000 187.200 ;
        RECT 566.000 186.200 566.800 187.000 ;
        RECT 583.600 183.600 584.400 184.400 ;
        RECT 12.400 173.600 13.200 174.400 ;
        RECT 6.000 172.200 6.800 173.000 ;
        RECT 14.000 171.800 14.800 172.600 ;
        RECT 33.200 174.800 34.000 175.600 ;
        RECT 44.400 174.800 45.200 175.600 ;
        RECT 47.600 173.600 48.400 174.400 ;
        RECT 18.800 170.200 19.600 171.000 ;
        RECT 1.200 163.600 2.000 164.400 ;
        RECT 33.200 167.600 34.000 168.400 ;
        RECT 58.800 173.600 59.600 174.400 ;
        RECT 60.400 171.600 61.200 172.400 ;
        RECT 44.400 165.600 45.200 166.400 ;
        RECT 55.600 163.600 56.400 164.400 ;
        RECT 89.200 174.800 90.000 175.600 ;
        RECT 74.800 171.600 75.600 172.400 ;
        RECT 92.400 173.600 93.200 174.400 ;
        RECT 103.600 173.600 104.400 174.400 ;
        RECT 106.800 173.600 107.600 174.400 ;
        RECT 81.200 169.600 82.000 170.400 ;
        RECT 110.000 171.800 110.800 172.600 ;
        RECT 105.200 170.200 106.000 171.000 ;
        RECT 100.400 163.600 101.200 164.400 ;
        RECT 122.800 163.600 123.600 164.400 ;
        RECT 138.800 171.800 139.600 172.600 ;
        RECT 127.600 169.600 128.400 170.400 ;
        RECT 134.000 170.200 134.800 171.000 ;
        RECT 154.800 173.600 155.600 174.400 ;
        RECT 158.000 171.800 158.800 172.600 ;
        RECT 151.600 163.600 152.400 164.400 ;
        RECT 153.200 170.200 154.000 171.000 ;
        RECT 178.800 174.800 179.600 175.600 ;
        RECT 182.000 173.600 182.800 174.400 ;
        RECT 186.800 171.600 187.600 172.400 ;
        RECT 207.600 175.600 208.400 176.400 ;
        RECT 204.400 173.600 205.200 174.400 ;
        RECT 198.000 171.600 198.800 172.400 ;
        RECT 202.800 171.600 203.600 172.400 ;
        RECT 170.800 163.600 171.600 164.400 ;
        RECT 178.800 165.600 179.600 166.400 ;
        RECT 199.600 169.600 200.400 170.400 ;
        RECT 215.600 169.600 216.400 170.400 ;
        RECT 220.400 167.600 221.200 168.400 ;
        RECT 234.800 173.600 235.600 174.400 ;
        RECT 238.000 171.800 238.800 172.600 ;
        RECT 226.800 169.600 227.600 170.400 ;
        RECT 230.000 169.600 230.800 170.400 ;
        RECT 231.600 169.600 232.400 170.400 ;
        RECT 233.200 170.200 234.000 171.000 ;
        RECT 265.200 173.600 266.000 174.400 ;
        RECT 268.400 173.600 269.200 174.400 ;
        RECT 308.400 177.600 309.200 178.400 ;
        RECT 276.400 173.600 277.200 174.400 ;
        RECT 271.600 171.800 272.400 172.600 ;
        RECT 250.800 163.600 251.600 164.400 ;
        RECT 266.800 170.200 267.600 171.000 ;
        RECT 292.400 173.600 293.200 174.400 ;
        RECT 326.000 177.600 326.800 178.400 ;
        RECT 295.600 171.800 296.400 172.600 ;
        RECT 284.400 167.600 285.200 168.400 ;
        RECT 290.800 170.200 291.600 171.000 ;
        RECT 305.200 167.600 306.000 168.400 ;
        RECT 310.000 169.600 310.800 170.400 ;
        RECT 319.600 169.600 320.400 170.400 ;
        RECT 351.600 177.600 352.400 178.400 ;
        RECT 335.600 169.600 336.400 170.400 ;
        RECT 346.800 169.600 347.600 170.400 ;
        RECT 353.200 171.600 354.000 172.400 ;
        RECT 351.600 169.600 352.400 170.400 ;
        RECT 362.800 175.600 363.600 176.400 ;
        RECT 361.200 171.600 362.000 172.400 ;
        RECT 372.400 177.600 373.200 178.400 ;
        RECT 361.200 167.600 362.000 168.400 ;
        RECT 394.800 177.600 395.600 178.400 ;
        RECT 374.000 173.600 374.800 174.400 ;
        RECT 375.600 171.600 376.400 172.400 ;
        RECT 380.400 171.600 381.200 172.400 ;
        RECT 390.000 171.600 390.800 172.400 ;
        RECT 385.200 169.600 386.000 170.400 ;
        RECT 391.600 169.600 392.400 170.400 ;
        RECT 399.600 169.600 400.400 170.400 ;
        RECT 415.600 177.600 416.400 178.400 ;
        RECT 398.000 163.600 398.800 164.400 ;
        RECT 404.400 163.600 405.200 164.400 ;
        RECT 439.600 177.600 440.400 178.400 ;
        RECT 433.200 173.600 434.000 174.400 ;
        RECT 426.800 171.800 427.600 172.600 ;
        RECT 417.200 169.600 418.000 170.400 ;
        RECT 422.000 170.200 422.800 171.000 ;
        RECT 449.200 174.800 450.000 175.600 ;
        RECT 474.800 177.600 475.600 178.400 ;
        RECT 455.600 173.600 456.400 174.400 ;
        RECT 458.800 173.600 459.600 174.400 ;
        RECT 452.400 171.600 453.200 172.400 ;
        RECT 462.000 171.800 462.800 172.600 ;
        RECT 457.200 170.200 458.000 171.000 ;
        RECT 476.400 177.600 477.200 178.400 ;
        RECT 486.000 177.600 486.800 178.400 ;
        RECT 482.800 174.800 483.600 175.600 ;
        RECT 492.400 177.600 493.200 178.400 ;
        RECT 489.200 173.600 490.000 174.400 ;
        RECT 500.400 177.600 501.200 178.400 ;
        RECT 519.600 177.600 520.400 178.400 ;
        RECT 498.800 169.600 499.600 170.400 ;
        RECT 516.400 173.600 517.200 174.400 ;
        RECT 511.600 171.600 512.400 172.400 ;
        RECT 518.000 171.600 518.800 172.400 ;
        RECT 510.000 169.600 510.800 170.400 ;
        RECT 513.200 167.600 514.000 168.400 ;
        RECT 530.800 169.600 531.600 170.400 ;
        RECT 527.600 165.600 528.400 166.400 ;
        RECT 538.800 171.600 539.600 172.400 ;
        RECT 545.200 171.600 546.000 172.400 ;
        RECT 550.000 171.600 550.800 172.400 ;
        RECT 553.200 171.600 554.000 172.400 ;
        RECT 558.000 170.200 558.800 171.000 ;
        RECT 535.600 163.600 536.400 164.400 ;
        RECT 551.600 163.600 552.400 164.400 ;
        RECT 575.600 167.600 576.400 168.400 ;
        RECT 20.400 157.600 21.200 158.400 ;
        RECT 7.600 145.600 8.400 146.400 ;
        RECT 6.000 143.600 6.800 144.400 ;
        RECT 15.600 149.600 16.400 150.400 ;
        RECT 18.800 145.600 19.600 146.400 ;
        RECT 36.400 149.600 37.200 150.400 ;
        RECT 41.200 149.600 42.000 150.400 ;
        RECT 38.000 147.600 38.800 148.400 ;
        RECT 46.000 147.600 46.800 148.400 ;
        RECT 50.800 147.600 51.600 148.400 ;
        RECT 74.800 153.600 75.600 154.400 ;
        RECT 70.000 151.800 70.800 152.600 ;
        RECT 22.000 143.600 22.800 144.400 ;
        RECT 33.200 143.600 34.000 144.400 ;
        RECT 54.000 143.600 54.800 144.400 ;
        RECT 66.800 145.600 67.600 146.400 ;
        RECT 70.000 146.200 70.800 147.000 ;
        RECT 78.000 147.600 78.800 148.400 ;
        RECT 74.800 146.400 75.600 147.200 ;
        RECT 82.800 143.600 83.600 144.400 ;
        RECT 90.800 143.600 91.600 144.400 ;
        RECT 97.200 145.600 98.000 146.400 ;
        RECT 98.800 145.600 99.600 146.400 ;
        RECT 106.800 147.600 107.600 148.400 ;
        RECT 113.200 151.800 114.000 152.600 ;
        RECT 143.600 151.800 144.400 152.600 ;
        RECT 110.000 145.600 110.800 146.400 ;
        RECT 113.200 146.200 114.000 147.000 ;
        RECT 121.200 147.600 122.000 148.400 ;
        RECT 188.200 151.800 189.000 152.600 ;
        RECT 199.800 151.800 200.600 152.600 ;
        RECT 118.000 146.400 118.800 147.200 ;
        RECT 134.000 145.600 134.800 146.400 ;
        RECT 143.600 146.200 144.400 147.000 ;
        RECT 148.400 146.400 149.200 147.200 ;
        RECT 148.400 143.600 149.200 144.400 ;
        RECT 153.200 146.200 154.000 147.000 ;
        RECT 172.400 149.600 173.200 150.400 ;
        RECT 201.000 149.800 201.800 150.600 ;
        RECT 170.800 143.600 171.600 144.400 ;
        RECT 188.200 146.200 189.000 147.000 ;
        RECT 196.400 147.600 197.200 148.400 ;
        RECT 193.200 143.600 194.000 144.400 ;
        RECT 199.800 146.200 200.600 147.000 ;
        RECT 207.600 147.600 208.400 148.400 ;
        RECT 215.600 151.800 216.400 152.600 ;
        RECT 212.400 147.600 213.200 148.400 ;
        RECT 215.600 146.200 216.400 147.000 ;
        RECT 223.600 147.600 224.400 148.400 ;
        RECT 220.400 146.400 221.200 147.200 ;
        RECT 220.400 143.600 221.200 144.400 ;
        RECT 228.400 145.600 229.200 146.400 ;
        RECT 239.600 153.600 240.400 154.400 ;
        RECT 234.800 151.800 235.600 152.600 ;
        RECT 231.600 145.600 232.400 146.400 ;
        RECT 234.800 146.200 235.600 147.000 ;
        RECT 226.800 143.600 227.600 144.400 ;
        RECT 230.000 143.600 230.800 144.400 ;
        RECT 242.800 147.600 243.600 148.400 ;
        RECT 239.600 146.400 240.400 147.200 ;
        RECT 244.400 145.600 245.200 146.400 ;
        RECT 257.200 147.600 258.000 148.400 ;
        RECT 258.800 147.600 259.600 148.400 ;
        RECT 279.600 151.800 280.400 152.600 ;
        RECT 308.400 153.600 309.200 154.400 ;
        RECT 274.800 149.600 275.600 150.400 ;
        RECT 273.200 147.600 274.000 148.400 ;
        RECT 276.400 147.600 277.200 148.400 ;
        RECT 279.600 146.200 280.400 147.000 ;
        RECT 287.600 147.600 288.400 148.400 ;
        RECT 284.400 146.400 285.200 147.200 ;
        RECT 294.000 146.200 294.800 147.000 ;
        RECT 314.800 147.600 315.600 148.400 ;
        RECT 311.600 143.600 312.400 144.400 ;
        RECT 313.200 146.200 314.000 147.000 ;
        RECT 356.400 157.600 357.200 158.400 ;
        RECT 348.400 149.600 349.200 150.400 ;
        RECT 356.400 149.600 357.200 150.400 ;
        RECT 330.800 143.600 331.600 144.400 ;
        RECT 364.400 149.600 365.200 150.400 ;
        RECT 370.800 149.600 371.600 150.400 ;
        RECT 385.200 151.600 386.000 152.400 ;
        RECT 385.200 149.600 386.000 150.400 ;
        RECT 391.600 149.600 392.400 150.400 ;
        RECT 343.600 143.600 344.400 144.400 ;
        RECT 361.200 145.600 362.000 146.400 ;
        RECT 380.400 147.600 381.200 148.400 ;
        RECT 374.000 145.600 374.800 146.400 ;
        RECT 386.800 147.600 387.600 148.400 ;
        RECT 390.000 147.600 390.800 148.400 ;
        RECT 393.200 147.600 394.000 148.400 ;
        RECT 418.800 157.600 419.600 158.400 ;
        RECT 414.000 149.600 414.800 150.400 ;
        RECT 394.800 145.600 395.600 146.400 ;
        RECT 415.600 149.600 416.400 150.400 ;
        RECT 410.800 145.600 411.600 146.400 ;
        RECT 447.600 157.600 448.400 158.400 ;
        RECT 431.600 145.600 432.400 146.400 ;
        RECT 433.200 145.600 434.000 146.400 ;
        RECT 439.600 149.600 440.400 150.400 ;
        RECT 436.400 143.600 437.200 144.400 ;
        RECT 458.800 149.600 459.600 150.400 ;
        RECT 486.000 157.600 486.800 158.400 ;
        RECT 449.200 145.600 450.000 146.400 ;
        RECT 466.800 147.600 467.600 148.400 ;
        RECT 470.000 147.600 470.800 148.400 ;
        RECT 468.400 146.200 469.200 147.000 ;
        RECT 487.600 149.600 488.400 150.400 ;
        RECT 516.400 149.600 517.200 150.400 ;
        RECT 505.200 147.600 506.000 148.400 ;
        RECT 538.800 153.600 539.600 154.400 ;
        RECT 527.600 149.600 528.400 150.400 ;
        RECT 529.200 149.600 530.000 150.400 ;
        RECT 542.000 151.600 542.800 152.400 ;
        RECT 540.400 149.600 541.200 150.400 ;
        RECT 510.000 143.600 510.800 144.400 ;
        RECT 524.400 143.600 525.200 144.400 ;
        RECT 532.400 145.600 533.200 146.400 ;
        RECT 543.600 147.600 544.400 148.400 ;
        RECT 559.600 157.600 560.400 158.400 ;
        RECT 554.600 151.800 555.400 152.600 ;
        RECT 570.800 149.600 571.600 150.400 ;
        RECT 551.600 145.600 552.400 146.400 ;
        RECT 554.600 146.200 555.400 147.000 ;
        RECT 562.800 147.600 563.600 148.400 ;
        RECT 564.400 146.200 565.200 147.000 ;
        RECT 4.400 131.600 5.200 132.400 ;
        RECT 14.000 129.600 14.800 130.400 ;
        RECT 23.600 131.600 24.400 132.400 ;
        RECT 25.200 131.600 26.000 132.400 ;
        RECT 30.000 131.600 30.800 132.400 ;
        RECT 44.400 137.600 45.200 138.400 ;
        RECT 41.200 129.600 42.000 130.400 ;
        RECT 57.200 133.600 58.000 134.400 ;
        RECT 50.800 129.600 51.600 130.400 ;
        RECT 57.200 129.600 58.000 130.400 ;
        RECT 62.000 129.600 62.800 130.400 ;
        RECT 68.400 131.600 69.200 132.400 ;
        RECT 63.600 123.600 64.400 124.400 ;
        RECT 71.600 123.600 72.400 124.400 ;
        RECT 81.200 129.600 82.000 130.400 ;
        RECT 97.200 129.600 98.000 130.400 ;
        RECT 105.200 129.600 106.000 130.400 ;
        RECT 121.200 137.600 122.000 138.400 ;
        RECT 129.200 137.600 130.000 138.400 ;
        RECT 102.000 123.600 102.800 124.400 ;
        RECT 119.600 129.600 120.400 130.400 ;
        RECT 127.600 129.600 128.400 130.400 ;
        RECT 143.600 134.800 144.400 135.600 ;
        RECT 151.600 134.800 152.400 135.600 ;
        RECT 146.800 133.600 147.600 134.400 ;
        RECT 158.000 133.600 158.800 134.400 ;
        RECT 164.400 131.800 165.200 132.600 ;
        RECT 159.600 130.200 160.400 131.000 ;
        RECT 142.000 123.600 142.800 124.400 ;
        RECT 174.000 127.600 174.800 128.400 ;
        RECT 177.200 123.600 178.000 124.400 ;
        RECT 201.200 137.600 202.000 138.400 ;
        RECT 182.000 129.600 182.800 130.400 ;
        RECT 185.200 129.600 186.000 130.400 ;
        RECT 196.400 129.600 197.200 130.400 ;
        RECT 231.600 133.600 232.400 134.400 ;
        RECT 201.200 129.600 202.000 130.400 ;
        RECT 210.800 127.600 211.600 128.400 ;
        RECT 204.400 123.600 205.200 124.400 ;
        RECT 218.800 129.600 219.600 130.400 ;
        RECT 223.600 123.600 224.400 124.400 ;
        RECT 231.600 129.600 232.400 130.400 ;
        RECT 238.000 129.600 238.800 130.400 ;
        RECT 250.800 133.600 251.600 134.400 ;
        RECT 268.400 129.600 269.200 130.400 ;
        RECT 274.800 129.600 275.600 130.400 ;
        RECT 276.400 129.600 277.200 130.400 ;
        RECT 302.000 134.800 302.800 135.600 ;
        RECT 324.400 137.600 325.200 138.400 ;
        RECT 305.200 133.600 306.000 134.400 ;
        RECT 308.400 133.600 309.200 134.400 ;
        RECT 314.800 133.600 315.600 134.400 ;
        RECT 289.200 129.600 290.000 130.400 ;
        RECT 311.600 131.800 312.400 132.600 ;
        RECT 306.800 130.200 307.600 131.000 ;
        RECT 302.000 123.600 302.800 124.400 ;
        RECT 332.400 134.800 333.200 135.600 ;
        RECT 335.600 133.600 336.400 134.400 ;
        RECT 343.600 134.800 344.400 135.600 ;
        RECT 351.600 134.800 352.400 135.600 ;
        RECT 370.800 137.600 371.600 138.400 ;
        RECT 358.000 133.600 358.800 134.400 ;
        RECT 332.400 125.600 333.200 126.400 ;
        RECT 343.600 129.600 344.400 130.400 ;
        RECT 354.800 131.600 355.600 132.400 ;
        RECT 367.600 129.600 368.400 130.400 ;
        RECT 378.800 135.600 379.600 136.400 ;
        RECT 386.800 137.600 387.600 138.400 ;
        RECT 393.200 137.600 394.000 138.400 ;
        RECT 366.000 127.600 366.800 128.400 ;
        RECT 380.400 129.600 381.200 130.400 ;
        RECT 382.000 123.600 382.800 124.400 ;
        RECT 410.800 137.600 411.600 138.400 ;
        RECT 393.200 129.600 394.000 130.400 ;
        RECT 404.400 133.600 405.200 134.400 ;
        RECT 426.800 137.600 427.600 138.400 ;
        RECT 399.600 131.600 400.400 132.400 ;
        RECT 406.000 131.600 406.800 132.400 ;
        RECT 414.000 131.600 414.800 132.400 ;
        RECT 415.600 131.600 416.400 132.400 ;
        RECT 426.800 134.800 427.600 135.600 ;
        RECT 462.000 137.600 462.800 138.400 ;
        RECT 430.000 133.600 430.800 134.400 ;
        RECT 433.200 133.600 434.000 134.400 ;
        RECT 441.200 131.600 442.000 132.400 ;
        RECT 479.600 137.600 480.400 138.400 ;
        RECT 465.200 129.600 466.000 130.400 ;
        RECT 471.600 129.600 472.400 130.400 ;
        RECT 521.200 137.600 522.000 138.400 ;
        RECT 495.600 133.600 496.400 134.400 ;
        RECT 484.400 132.200 485.200 133.000 ;
        RECT 497.200 130.200 498.000 131.000 ;
        RECT 510.000 123.600 510.800 124.400 ;
        RECT 516.400 129.600 517.200 130.400 ;
        RECT 526.000 129.600 526.800 130.400 ;
        RECT 529.200 123.600 530.000 124.400 ;
        RECT 535.600 129.600 536.400 130.400 ;
        RECT 540.400 129.600 541.200 130.400 ;
        RECT 548.400 133.600 549.200 134.400 ;
        RECT 562.800 134.800 563.600 135.600 ;
        RECT 566.000 133.600 566.800 134.400 ;
        RECT 574.000 134.800 574.800 135.600 ;
        RECT 577.200 133.600 578.000 134.400 ;
        RECT 2.800 109.600 3.600 110.400 ;
        RECT 23.400 111.800 24.200 112.600 ;
        RECT 6.000 105.600 6.800 106.400 ;
        RECT 12.400 103.600 13.200 104.400 ;
        RECT 17.200 103.600 18.000 104.400 ;
        RECT 23.400 106.200 24.200 107.000 ;
        RECT 38.000 107.600 38.800 108.400 ;
        RECT 33.200 105.600 34.000 106.400 ;
        RECT 42.800 109.600 43.600 110.400 ;
        RECT 44.400 109.600 45.200 110.400 ;
        RECT 47.600 105.600 48.400 106.400 ;
        RECT 49.200 103.600 50.000 104.400 ;
        RECT 54.000 105.600 54.800 106.400 ;
        RECT 60.400 107.600 61.200 108.400 ;
        RECT 78.000 113.600 78.800 114.400 ;
        RECT 73.200 111.800 74.000 112.600 ;
        RECT 55.600 103.600 56.400 104.400 ;
        RECT 66.800 103.600 67.600 104.400 ;
        RECT 73.200 106.200 74.000 107.000 ;
        RECT 81.200 107.600 82.000 108.400 ;
        RECT 78.000 106.400 78.800 107.200 ;
        RECT 89.200 107.600 90.000 108.400 ;
        RECT 94.000 105.600 94.800 106.400 ;
        RECT 105.200 109.600 106.000 110.400 ;
        RECT 111.600 109.600 112.400 110.400 ;
        RECT 106.800 107.600 107.600 108.400 ;
        RECT 102.000 105.600 102.800 106.400 ;
        RECT 100.400 103.600 101.200 104.400 ;
        RECT 122.800 105.600 123.600 106.400 ;
        RECT 127.600 105.600 128.400 106.400 ;
        RECT 124.400 103.600 125.200 104.400 ;
        RECT 151.800 111.800 152.600 112.600 ;
        RECT 153.000 109.800 153.800 110.600 ;
        RECT 182.000 113.600 182.800 114.400 ;
        RECT 143.600 105.600 144.400 106.400 ;
        RECT 145.200 105.600 146.000 106.400 ;
        RECT 151.800 106.200 152.600 107.000 ;
        RECT 159.600 107.600 160.400 108.400 ;
        RECT 162.800 105.600 163.600 106.400 ;
        RECT 164.400 106.200 165.200 107.000 ;
        RECT 183.600 107.600 184.400 108.400 ;
        RECT 169.200 105.600 170.000 106.400 ;
        RECT 188.400 107.600 189.200 108.400 ;
        RECT 194.800 107.600 195.600 108.400 ;
        RECT 201.200 107.600 202.000 108.400 ;
        RECT 233.200 111.600 234.000 112.400 ;
        RECT 214.000 107.600 214.800 108.400 ;
        RECT 196.400 103.600 197.200 104.400 ;
        RECT 206.000 103.600 206.800 104.400 ;
        RECT 233.200 109.600 234.000 110.400 ;
        RECT 252.400 117.600 253.200 118.400 ;
        RECT 247.600 111.800 248.400 112.600 ;
        RECT 234.800 107.600 235.600 108.400 ;
        RECT 242.800 109.600 243.600 110.400 ;
        RECT 244.400 109.600 245.200 110.400 ;
        RECT 247.600 106.200 248.400 107.000 ;
        RECT 255.600 107.600 256.400 108.400 ;
        RECT 252.400 106.400 253.200 107.200 ;
        RECT 257.200 105.600 258.000 106.400 ;
        RECT 268.400 109.600 269.200 110.400 ;
        RECT 263.600 107.600 264.400 108.400 ;
        RECT 271.600 107.600 272.400 108.400 ;
        RECT 289.200 113.600 290.000 114.400 ;
        RECT 284.400 111.800 285.200 112.600 ;
        RECT 278.000 109.600 278.800 110.400 ;
        RECT 279.600 109.600 280.400 110.400 ;
        RECT 306.800 117.600 307.600 118.400 ;
        RECT 258.800 103.600 259.600 104.400 ;
        RECT 265.200 103.600 266.000 104.400 ;
        RECT 284.400 106.200 285.200 107.000 ;
        RECT 292.400 107.600 293.200 108.400 ;
        RECT 298.800 107.600 299.600 108.400 ;
        RECT 289.200 106.400 290.000 107.200 ;
        RECT 300.400 103.600 301.200 104.400 ;
        RECT 345.200 117.600 346.000 118.400 ;
        RECT 308.400 106.200 309.200 107.000 ;
        RECT 348.400 117.600 349.200 118.400 ;
        RECT 329.200 107.600 330.000 108.400 ;
        RECT 326.000 103.600 326.800 104.400 ;
        RECT 327.600 106.200 328.400 107.000 ;
        RECT 356.400 117.600 357.200 118.400 ;
        RECT 362.800 113.600 363.600 114.400 ;
        RECT 351.600 109.600 352.400 110.400 ;
        RECT 367.600 109.600 368.400 110.400 ;
        RECT 375.600 109.600 376.400 110.400 ;
        RECT 356.400 103.600 357.200 104.400 ;
        RECT 378.800 109.600 379.600 110.400 ;
        RECT 380.400 109.600 381.200 110.400 ;
        RECT 386.800 107.600 387.600 108.400 ;
        RECT 382.000 105.600 382.800 106.400 ;
        RECT 417.200 117.600 418.000 118.400 ;
        RECT 398.000 107.600 398.800 108.400 ;
        RECT 399.600 105.600 400.400 106.400 ;
        RECT 401.200 103.600 402.000 104.400 ;
        RECT 422.000 111.800 422.800 112.600 ;
        RECT 449.200 117.600 450.000 118.400 ;
        RECT 417.200 109.600 418.000 110.400 ;
        RECT 406.000 105.600 406.800 106.400 ;
        RECT 418.800 107.600 419.600 108.400 ;
        RECT 422.000 106.200 422.800 107.000 ;
        RECT 430.000 107.600 430.800 108.400 ;
        RECT 433.200 107.600 434.000 108.400 ;
        RECT 426.800 106.400 427.600 107.200 ;
        RECT 431.600 106.200 432.400 107.000 ;
        RECT 457.200 117.600 458.000 118.400 ;
        RECT 458.800 107.600 459.600 108.400 ;
        RECT 463.600 117.600 464.400 118.400 ;
        RECT 470.000 111.800 470.800 112.600 ;
        RECT 462.000 107.600 462.800 108.400 ;
        RECT 466.800 109.600 467.600 110.400 ;
        RECT 470.000 106.200 470.800 107.000 ;
        RECT 478.000 107.600 478.800 108.400 ;
        RECT 479.600 107.600 480.400 108.400 ;
        RECT 474.800 106.400 475.600 107.200 ;
        RECT 502.000 117.600 502.800 118.400 ;
        RECT 521.200 117.600 522.000 118.400 ;
        RECT 518.000 113.600 518.800 114.400 ;
        RECT 481.200 103.600 482.000 104.400 ;
        RECT 484.400 106.200 485.200 107.000 ;
        RECT 524.200 111.800 525.000 112.600 ;
        RECT 535.400 111.800 536.200 112.600 ;
        RECT 562.800 113.600 563.600 114.400 ;
        RECT 503.600 106.200 504.400 107.000 ;
        RECT 524.200 106.200 525.000 107.000 ;
        RECT 551.600 109.600 552.400 110.400 ;
        RECT 582.000 117.600 582.800 118.400 ;
        RECT 532.400 107.600 533.200 108.400 ;
        RECT 529.200 103.600 530.000 104.400 ;
        RECT 535.400 106.200 536.200 107.000 ;
        RECT 543.600 107.600 544.400 108.400 ;
        RECT 540.400 103.600 541.200 104.400 ;
        RECT 545.200 106.200 546.000 107.000 ;
        RECT 566.000 107.600 566.800 108.400 ;
        RECT 564.400 106.200 565.200 107.000 ;
        RECT 2.800 97.600 3.600 98.400 ;
        RECT 22.000 97.600 22.800 98.400 ;
        RECT 9.200 83.600 10.000 84.400 ;
        RECT 18.800 89.600 19.600 90.400 ;
        RECT 25.200 91.600 26.000 92.400 ;
        RECT 30.000 91.600 30.800 92.400 ;
        RECT 33.200 87.600 34.000 88.400 ;
        RECT 39.600 89.600 40.400 90.400 ;
        RECT 52.400 95.600 53.200 96.400 ;
        RECT 47.600 85.600 48.400 86.400 ;
        RECT 58.800 95.600 59.600 96.400 ;
        RECT 63.600 93.600 64.400 94.400 ;
        RECT 62.000 91.600 62.800 92.400 ;
        RECT 65.200 91.600 66.000 92.400 ;
        RECT 71.600 89.600 72.400 90.400 ;
        RECT 76.400 89.600 77.200 90.400 ;
        RECT 74.800 87.600 75.600 88.400 ;
        RECT 87.600 97.600 88.400 98.400 ;
        RECT 94.000 95.600 94.800 96.400 ;
        RECT 105.200 97.600 106.000 98.400 ;
        RECT 97.200 93.600 98.000 94.400 ;
        RECT 110.000 93.600 110.800 94.400 ;
        RECT 126.000 97.600 126.800 98.400 ;
        RECT 119.600 93.600 120.400 94.400 ;
        RECT 146.800 97.600 147.600 98.400 ;
        RECT 175.600 97.600 176.400 98.400 ;
        RECT 129.200 91.600 130.000 92.400 ;
        RECT 134.000 91.600 134.800 92.400 ;
        RECT 143.600 83.600 144.400 84.400 ;
        RECT 153.200 89.600 154.000 90.400 ;
        RECT 166.000 93.600 166.800 94.400 ;
        RECT 162.800 91.800 163.600 92.600 ;
        RECT 158.000 90.200 158.800 91.000 ;
        RECT 177.200 91.600 178.000 92.400 ;
        RECT 223.600 97.600 224.400 98.400 ;
        RECT 185.200 91.600 186.000 92.400 ;
        RECT 186.800 91.600 187.600 92.400 ;
        RECT 194.800 91.600 195.600 92.400 ;
        RECT 201.200 89.600 202.000 90.400 ;
        RECT 206.000 83.600 206.800 84.400 ;
        RECT 217.200 93.600 218.000 94.400 ;
        RECT 212.400 91.600 213.200 92.400 ;
        RECT 218.800 91.600 219.600 92.400 ;
        RECT 214.000 83.600 214.800 84.400 ;
        RECT 236.400 93.600 237.200 94.400 ;
        RECT 223.600 89.600 224.400 90.400 ;
        RECT 241.200 91.600 242.000 92.400 ;
        RECT 246.000 91.600 246.800 92.400 ;
        RECT 239.600 83.600 240.400 84.400 ;
        RECT 263.600 94.800 264.400 95.600 ;
        RECT 266.800 93.600 267.600 94.400 ;
        RECT 254.000 91.600 254.800 92.400 ;
        RECT 282.800 89.600 283.600 90.400 ;
        RECT 302.000 89.600 302.800 90.400 ;
        RECT 316.400 91.800 317.200 92.600 ;
        RECT 310.000 89.600 310.800 90.400 ;
        RECT 311.600 90.200 312.400 91.000 ;
        RECT 308.400 83.600 309.200 84.400 ;
        RECT 335.600 91.800 336.400 92.600 ;
        RECT 329.200 83.600 330.000 84.400 ;
        RECT 330.800 90.200 331.600 91.000 ;
        RECT 345.200 87.600 346.000 88.400 ;
        RECT 348.400 87.600 349.200 88.400 ;
        RECT 374.000 97.600 374.800 98.400 ;
        RECT 374.000 94.800 374.800 95.600 ;
        RECT 393.200 97.600 394.000 98.400 ;
        RECT 377.200 93.600 378.000 94.400 ;
        RECT 391.600 93.600 392.400 94.400 ;
        RECT 382.000 91.600 382.800 92.400 ;
        RECT 407.600 97.600 408.400 98.400 ;
        RECT 410.800 97.600 411.600 98.400 ;
        RECT 396.400 93.600 397.200 94.400 ;
        RECT 382.000 87.600 382.800 88.400 ;
        RECT 388.400 89.600 389.200 90.400 ;
        RECT 407.600 89.600 408.400 90.400 ;
        RECT 409.200 89.600 410.000 90.400 ;
        RECT 414.000 93.600 414.800 94.400 ;
        RECT 426.800 93.600 427.600 94.400 ;
        RECT 433.200 93.600 434.000 94.400 ;
        RECT 462.000 97.600 462.800 98.400 ;
        RECT 422.000 89.600 422.800 90.400 ;
        RECT 436.400 91.800 437.200 92.600 ;
        RECT 431.600 90.200 432.400 91.000 ;
        RECT 462.000 94.800 462.800 95.600 ;
        RECT 470.000 94.800 470.800 95.600 ;
        RECT 465.200 93.600 466.000 94.400 ;
        RECT 479.600 95.600 480.400 96.400 ;
        RECT 476.400 93.600 477.200 94.400 ;
        RECT 490.800 97.600 491.600 98.400 ;
        RECT 510.000 97.600 510.800 98.400 ;
        RECT 494.000 93.600 494.800 94.400 ;
        RECT 497.200 91.800 498.000 92.600 ;
        RECT 490.800 89.600 491.600 90.400 ;
        RECT 492.400 90.200 493.200 91.000 ;
        RECT 511.600 97.600 512.400 98.400 ;
        RECT 542.000 93.600 542.800 94.400 ;
        RECT 516.400 92.200 517.200 93.000 ;
        RECT 524.400 91.800 525.200 92.600 ;
        RECT 529.200 90.200 530.000 91.000 ;
        RECT 530.800 90.200 531.600 91.000 ;
        RECT 548.400 87.600 549.200 88.400 ;
        RECT 550.000 97.600 550.800 98.400 ;
        RECT 554.800 93.600 555.600 94.400 ;
        RECT 558.000 91.800 558.800 92.600 ;
        RECT 553.200 90.200 554.000 91.000 ;
        RECT 567.600 87.600 568.400 88.400 ;
        RECT 570.800 87.600 571.600 88.400 ;
        RECT 2.600 71.800 3.400 72.600 ;
        RECT 2.600 66.200 3.400 67.000 ;
        RECT 18.800 69.600 19.600 70.400 ;
        RECT 15.600 67.600 16.400 68.400 ;
        RECT 31.600 71.600 32.400 72.400 ;
        RECT 31.600 69.600 32.400 70.400 ;
        RECT 33.200 67.600 34.000 68.400 ;
        RECT 26.800 63.600 27.600 64.400 ;
        RECT 44.400 69.600 45.200 70.400 ;
        RECT 36.400 67.600 37.200 68.400 ;
        RECT 38.000 65.600 38.800 66.400 ;
        RECT 34.800 63.600 35.600 64.400 ;
        RECT 46.000 67.600 46.800 68.400 ;
        RECT 73.200 73.600 74.000 74.400 ;
        RECT 78.000 77.600 78.800 78.400 ;
        RECT 50.800 65.600 51.600 66.400 ;
        RECT 74.800 67.600 75.600 68.400 ;
        RECT 70.000 63.600 70.800 64.400 ;
        RECT 76.400 65.600 77.200 66.400 ;
        RECT 82.800 73.600 83.600 74.400 ;
        RECT 78.000 63.600 78.800 64.400 ;
        RECT 86.000 67.600 86.800 68.400 ;
        RECT 89.200 63.600 90.000 64.400 ;
        RECT 94.000 67.600 94.800 68.400 ;
        RECT 92.400 65.600 93.200 66.400 ;
        RECT 98.800 67.600 99.600 68.400 ;
        RECT 105.200 69.600 106.000 70.400 ;
        RECT 122.800 69.600 123.600 70.400 ;
        RECT 97.200 63.600 98.000 64.400 ;
        RECT 113.200 65.600 114.000 66.400 ;
        RECT 145.200 71.800 146.000 72.600 ;
        RECT 130.800 67.600 131.600 68.400 ;
        RECT 134.000 67.600 134.800 68.400 ;
        RECT 137.200 67.600 138.000 68.400 ;
        RECT 145.200 66.200 146.000 67.000 ;
        RECT 153.200 67.600 154.000 68.400 ;
        RECT 150.000 66.400 150.800 67.200 ;
        RECT 154.800 66.200 155.600 67.000 ;
        RECT 175.600 69.600 176.400 70.400 ;
        RECT 185.200 77.600 186.000 78.400 ;
        RECT 190.000 77.600 190.800 78.400 ;
        RECT 182.000 69.600 182.800 70.400 ;
        RECT 172.400 63.600 173.200 64.400 ;
        RECT 180.400 65.600 181.200 66.400 ;
        RECT 188.400 67.600 189.200 68.400 ;
        RECT 186.800 65.600 187.600 66.400 ;
        RECT 194.800 77.600 195.600 78.400 ;
        RECT 199.600 69.600 200.400 70.400 ;
        RECT 196.400 65.600 197.200 66.400 ;
        RECT 210.800 71.600 211.600 72.400 ;
        RECT 222.000 77.600 222.800 78.400 ;
        RECT 206.000 65.600 206.800 66.400 ;
        RECT 212.400 67.600 213.200 68.400 ;
        RECT 215.600 65.600 216.400 66.400 ;
        RECT 220.400 65.600 221.200 66.400 ;
        RECT 244.400 73.600 245.200 74.400 ;
        RECT 223.600 65.600 224.400 66.400 ;
        RECT 225.200 65.600 226.000 66.400 ;
        RECT 247.600 71.600 248.400 72.400 ;
        RECT 246.000 69.600 246.800 70.400 ;
        RECT 250.800 69.600 251.600 70.400 ;
        RECT 238.000 63.600 238.800 64.400 ;
        RECT 254.000 67.600 254.800 68.400 ;
        RECT 255.600 67.600 256.400 68.400 ;
        RECT 260.400 71.600 261.200 72.400 ;
        RECT 258.800 63.600 259.600 64.400 ;
        RECT 276.400 77.600 277.200 78.400 ;
        RECT 286.000 77.600 286.800 78.400 ;
        RECT 287.600 73.600 288.400 74.400 ;
        RECT 262.000 65.600 262.800 66.400 ;
        RECT 263.600 65.600 264.400 66.400 ;
        RECT 268.400 69.600 269.200 70.400 ;
        RECT 270.000 69.600 270.800 70.400 ;
        RECT 276.400 69.600 277.200 70.400 ;
        RECT 284.400 71.600 285.200 72.400 ;
        RECT 279.600 65.600 280.400 66.400 ;
        RECT 295.600 65.600 296.400 66.400 ;
        RECT 302.000 69.600 302.800 70.400 ;
        RECT 303.600 67.600 304.400 68.400 ;
        RECT 310.000 69.600 310.800 70.400 ;
        RECT 311.600 69.600 312.400 70.400 ;
        RECT 306.800 65.600 307.600 66.400 ;
        RECT 305.200 63.600 306.000 64.400 ;
        RECT 316.400 65.600 317.200 66.400 ;
        RECT 319.600 65.600 320.400 66.400 ;
        RECT 327.600 65.600 328.400 66.400 ;
        RECT 334.000 71.800 334.800 72.600 ;
        RECT 361.200 77.600 362.000 78.400 ;
        RECT 326.000 63.600 326.800 64.400 ;
        RECT 334.000 66.200 334.800 67.000 ;
        RECT 342.000 67.600 342.800 68.400 ;
        RECT 345.200 67.600 346.000 68.400 ;
        RECT 338.800 66.400 339.600 67.200 ;
        RECT 338.800 63.600 339.600 64.400 ;
        RECT 343.600 66.200 344.400 67.000 ;
        RECT 364.400 67.600 365.200 68.400 ;
        RECT 362.800 66.200 363.600 67.000 ;
        RECT 383.600 77.600 384.400 78.400 ;
        RECT 380.400 63.600 381.200 64.400 ;
        RECT 399.600 69.600 400.400 70.400 ;
        RECT 401.200 67.600 402.000 68.400 ;
        RECT 414.000 71.600 414.800 72.400 ;
        RECT 412.400 67.600 413.200 68.400 ;
        RECT 415.600 65.600 416.400 66.400 ;
        RECT 423.600 67.600 424.400 68.400 ;
        RECT 428.400 77.600 429.200 78.400 ;
        RECT 439.600 71.800 440.400 72.600 ;
        RECT 468.400 77.600 469.200 78.400 ;
        RECT 463.400 71.800 464.200 72.600 ;
        RECT 422.000 65.600 422.800 66.400 ;
        RECT 426.800 65.600 427.600 66.400 ;
        RECT 420.400 63.600 421.200 64.400 ;
        RECT 430.000 65.600 430.800 66.400 ;
        RECT 455.600 69.600 456.400 70.400 ;
        RECT 439.600 66.200 440.400 67.000 ;
        RECT 434.800 63.600 435.600 64.400 ;
        RECT 447.600 67.600 448.400 68.400 ;
        RECT 458.800 69.600 459.600 70.400 ;
        RECT 474.800 69.600 475.600 70.400 ;
        RECT 457.200 67.600 458.000 68.400 ;
        RECT 444.400 66.400 445.200 67.200 ;
        RECT 460.400 67.600 461.200 68.400 ;
        RECT 463.400 66.200 464.200 67.000 ;
        RECT 471.600 67.600 472.400 68.400 ;
        RECT 478.000 65.600 478.800 66.400 ;
        RECT 479.600 65.600 480.400 66.400 ;
        RECT 484.400 65.600 485.200 66.400 ;
        RECT 518.000 73.600 518.800 74.400 ;
        RECT 529.200 77.600 530.000 78.400 ;
        RECT 490.800 69.600 491.600 70.400 ;
        RECT 497.200 69.600 498.000 70.400 ;
        RECT 492.400 67.600 493.200 68.400 ;
        RECT 498.800 67.600 499.600 68.400 ;
        RECT 500.400 65.600 501.200 66.400 ;
        RECT 506.800 69.600 507.600 70.400 ;
        RECT 532.400 73.600 533.200 74.400 ;
        RECT 529.200 69.600 530.000 70.400 ;
        RECT 508.400 67.600 509.200 68.400 ;
        RECT 513.200 65.600 514.000 66.400 ;
        RECT 514.800 65.600 515.600 66.400 ;
        RECT 530.800 67.600 531.600 68.400 ;
        RECT 535.600 69.600 536.400 70.400 ;
        RECT 559.600 73.600 560.400 74.400 ;
        RECT 578.800 73.600 579.600 74.400 ;
        RECT 540.400 67.600 541.200 68.400 ;
        RECT 542.000 66.200 542.800 67.000 ;
        RECT 561.200 66.200 562.000 67.000 ;
        RECT 572.400 67.600 573.200 68.400 ;
        RECT 580.400 69.600 581.200 70.400 ;
        RECT 9.200 57.600 10.000 58.400 ;
        RECT 1.200 51.600 2.000 52.400 ;
        RECT 9.200 49.600 10.000 50.400 ;
        RECT 14.000 49.600 14.800 50.400 ;
        RECT 18.800 51.600 19.600 52.400 ;
        RECT 30.000 53.600 30.800 54.400 ;
        RECT 25.200 51.600 26.000 52.400 ;
        RECT 31.600 51.600 32.400 52.400 ;
        RECT 41.200 53.600 42.000 54.400 ;
        RECT 23.600 49.600 24.400 50.400 ;
        RECT 42.800 51.600 43.600 52.400 ;
        RECT 47.600 51.600 48.400 52.400 ;
        RECT 44.400 43.600 45.200 44.400 ;
        RECT 62.000 55.600 62.800 56.400 ;
        RECT 58.800 43.600 59.600 44.400 ;
        RECT 66.800 53.600 67.600 54.400 ;
        RECT 68.400 51.600 69.200 52.400 ;
        RECT 63.600 43.600 64.400 44.400 ;
        RECT 84.400 49.600 85.200 50.400 ;
        RECT 86.000 49.600 86.800 50.400 ;
        RECT 90.800 49.600 91.600 50.400 ;
        RECT 95.600 49.600 96.400 50.400 ;
        RECT 92.400 43.600 93.200 44.400 ;
        RECT 105.200 49.600 106.000 50.400 ;
        RECT 113.200 53.600 114.000 54.400 ;
        RECT 121.200 57.600 122.000 58.400 ;
        RECT 114.800 49.600 115.600 50.400 ;
        RECT 130.800 55.600 131.600 56.400 ;
        RECT 143.600 57.600 144.400 58.400 ;
        RECT 126.000 53.600 126.800 54.400 ;
        RECT 150.000 57.600 150.800 58.400 ;
        RECT 151.600 53.600 152.400 54.400 ;
        RECT 161.200 54.800 162.000 55.600 ;
        RECT 164.400 53.600 165.200 54.400 ;
        RECT 172.400 54.800 173.200 55.600 ;
        RECT 175.600 53.600 176.400 54.400 ;
        RECT 178.800 53.600 179.600 54.400 ;
        RECT 182.000 51.800 182.800 52.600 ;
        RECT 177.200 50.200 178.000 51.000 ;
        RECT 130.800 43.600 131.600 44.400 ;
        RECT 172.400 47.600 173.200 48.400 ;
        RECT 194.800 43.600 195.600 44.400 ;
        RECT 196.400 57.600 197.200 58.400 ;
        RECT 206.000 57.600 206.800 58.400 ;
        RECT 206.000 54.800 206.800 55.600 ;
        RECT 209.200 53.600 210.000 54.400 ;
        RECT 212.400 53.600 213.200 54.400 ;
        RECT 247.600 57.600 248.400 58.400 ;
        RECT 244.400 54.800 245.200 55.600 ;
        RECT 233.200 51.600 234.000 52.400 ;
        RECT 250.800 53.600 251.600 54.400 ;
        RECT 218.800 43.600 219.600 44.400 ;
        RECT 239.600 49.600 240.400 50.400 ;
        RECT 266.800 57.600 267.600 58.400 ;
        RECT 262.000 43.600 262.800 44.400 ;
        RECT 297.200 57.600 298.000 58.400 ;
        RECT 266.800 43.600 267.600 44.400 ;
        RECT 270.000 45.600 270.800 46.400 ;
        RECT 278.000 51.600 278.800 52.400 ;
        RECT 282.800 51.600 283.600 52.400 ;
        RECT 274.800 43.600 275.600 44.400 ;
        RECT 297.200 49.600 298.000 50.400 ;
        RECT 324.400 57.600 325.200 58.400 ;
        RECT 314.800 53.600 315.600 54.400 ;
        RECT 322.800 53.600 323.600 54.400 ;
        RECT 319.600 51.600 320.400 52.400 ;
        RECT 327.600 51.600 328.400 52.400 ;
        RECT 329.200 51.600 330.000 52.400 ;
        RECT 369.200 57.600 370.000 58.400 ;
        RECT 353.200 53.600 354.000 54.400 ;
        RECT 356.400 51.800 357.200 52.600 ;
        RECT 337.200 47.600 338.000 48.400 ;
        RECT 343.600 49.600 344.400 50.400 ;
        RECT 351.600 50.200 352.400 51.000 ;
        RECT 372.400 53.600 373.200 54.400 ;
        RECT 375.600 51.800 376.400 52.600 ;
        RECT 370.800 50.200 371.600 51.000 ;
        RECT 385.200 47.600 386.000 48.400 ;
        RECT 388.400 47.600 389.200 48.400 ;
        RECT 394.800 57.600 395.600 58.400 ;
        RECT 415.600 57.600 416.400 58.400 ;
        RECT 399.600 53.600 400.400 54.400 ;
        RECT 409.200 53.600 410.000 54.400 ;
        RECT 402.800 51.800 403.600 52.600 ;
        RECT 398.000 50.200 398.800 51.000 ;
        RECT 426.800 54.800 427.600 55.600 ;
        RECT 433.200 53.600 434.000 54.400 ;
        RECT 454.000 57.600 454.800 58.400 ;
        RECT 452.400 49.600 453.200 50.400 ;
        RECT 470.000 53.600 470.800 54.400 ;
        RECT 492.400 57.600 493.200 58.400 ;
        RECT 498.800 57.600 499.600 58.400 ;
        RECT 505.200 57.600 506.000 58.400 ;
        RECT 463.600 49.600 464.400 50.400 ;
        RECT 465.200 49.600 466.000 50.400 ;
        RECT 481.200 51.600 482.000 52.400 ;
        RECT 486.000 51.600 486.800 52.400 ;
        RECT 476.400 43.600 477.200 44.400 ;
        RECT 492.400 49.600 493.200 50.400 ;
        RECT 500.400 53.600 501.200 54.400 ;
        RECT 502.000 51.600 502.800 52.400 ;
        RECT 510.000 57.600 510.800 58.400 ;
        RECT 519.600 57.600 520.400 58.400 ;
        RECT 508.400 51.600 509.200 52.400 ;
        RECT 519.600 54.800 520.400 55.600 ;
        RECT 542.000 57.600 542.800 58.400 ;
        RECT 522.800 53.600 523.600 54.400 ;
        RECT 524.400 50.200 525.200 51.000 ;
        RECT 562.800 57.600 563.600 58.400 ;
        RECT 559.600 53.600 560.400 54.400 ;
        RECT 548.400 52.200 549.200 53.000 ;
        RECT 556.400 51.800 557.200 52.600 ;
        RECT 572.400 53.600 573.200 54.400 ;
        RECT 567.600 52.200 568.400 53.000 ;
        RECT 561.200 50.200 562.000 51.000 ;
        RECT 543.600 43.600 544.400 44.400 ;
        RECT 575.600 51.800 576.400 52.600 ;
        RECT 580.400 50.200 581.200 51.000 ;
        RECT 1.200 25.600 2.000 26.400 ;
        RECT 10.800 33.600 11.600 34.400 ;
        RECT 9.200 27.600 10.000 28.400 ;
        RECT 23.600 29.600 24.400 30.400 ;
        RECT 25.200 27.600 26.000 28.400 ;
        RECT 15.600 23.600 16.400 24.400 ;
        RECT 20.400 23.600 21.200 24.400 ;
        RECT 30.000 29.600 30.800 30.400 ;
        RECT 31.600 27.600 32.400 28.400 ;
        RECT 50.800 37.600 51.600 38.400 ;
        RECT 39.600 29.600 40.400 30.400 ;
        RECT 41.200 27.600 42.000 28.400 ;
        RECT 34.800 23.600 35.600 24.400 ;
        RECT 46.000 25.600 46.800 26.400 ;
        RECT 49.200 25.600 50.000 26.400 ;
        RECT 55.600 37.600 56.400 38.400 ;
        RECT 60.400 31.800 61.200 32.600 ;
        RECT 87.600 37.600 88.400 38.400 ;
        RECT 60.400 26.200 61.200 27.000 ;
        RECT 76.400 29.600 77.200 30.400 ;
        RECT 90.600 31.800 91.400 32.600 ;
        RECT 68.400 27.600 69.200 28.400 ;
        RECT 65.200 26.400 66.000 27.200 ;
        RECT 65.200 23.600 66.000 24.400 ;
        RECT 70.000 26.200 70.800 27.000 ;
        RECT 90.600 26.200 91.400 27.000 ;
        RECT 127.600 31.800 128.400 32.600 ;
        RECT 143.600 31.800 144.400 32.600 ;
        RECT 103.600 29.600 104.400 30.400 ;
        RECT 98.800 27.600 99.600 28.400 ;
        RECT 105.200 27.600 106.000 28.400 ;
        RECT 108.400 27.600 109.200 28.400 ;
        RECT 106.800 26.200 107.600 27.000 ;
        RECT 124.400 23.600 125.200 24.400 ;
        RECT 127.600 26.200 128.400 27.000 ;
        RECT 135.600 27.600 136.400 28.400 ;
        RECT 132.400 26.400 133.200 27.200 ;
        RECT 143.600 26.200 144.400 27.000 ;
        RECT 151.600 27.600 152.400 28.400 ;
        RECT 153.200 27.600 154.000 28.400 ;
        RECT 148.400 26.400 149.200 27.200 ;
        RECT 148.400 23.600 149.200 24.400 ;
        RECT 170.800 31.600 171.600 32.400 ;
        RECT 167.600 29.600 168.400 30.400 ;
        RECT 161.200 27.600 162.000 28.400 ;
        RECT 162.800 27.600 163.600 28.400 ;
        RECT 175.600 29.600 176.400 30.400 ;
        RECT 193.200 37.600 194.000 38.400 ;
        RECT 188.400 31.800 189.200 32.600 ;
        RECT 183.600 29.600 184.400 30.400 ;
        RECT 182.000 27.600 182.800 28.400 ;
        RECT 185.200 27.600 186.000 28.400 ;
        RECT 188.400 26.200 189.200 27.000 ;
        RECT 159.600 23.600 160.400 24.400 ;
        RECT 196.400 27.600 197.200 28.400 ;
        RECT 193.200 26.400 194.000 27.200 ;
        RECT 214.000 27.600 214.800 28.400 ;
        RECT 201.200 23.600 202.000 24.400 ;
        RECT 221.800 31.800 222.600 32.600 ;
        RECT 226.800 31.600 227.600 32.400 ;
        RECT 233.200 35.600 234.000 36.400 ;
        RECT 221.800 26.200 222.600 27.000 ;
        RECT 209.200 23.600 210.000 24.400 ;
        RECT 230.000 27.600 230.800 28.400 ;
        RECT 254.000 37.600 254.800 38.400 ;
        RECT 234.800 27.600 235.600 28.400 ;
        RECT 268.400 29.600 269.200 30.400 ;
        RECT 300.400 37.600 301.200 38.400 ;
        RECT 276.400 29.600 277.200 30.400 ;
        RECT 287.600 29.600 288.400 30.400 ;
        RECT 318.000 37.600 318.800 38.400 ;
        RECT 321.200 37.600 322.000 38.400 ;
        RECT 300.400 29.600 301.200 30.400 ;
        RECT 310.000 29.600 310.800 30.400 ;
        RECT 318.000 29.600 318.800 30.400 ;
        RECT 265.200 27.600 266.000 28.400 ;
        RECT 278.000 27.600 278.800 28.400 ;
        RECT 302.000 27.600 302.800 28.400 ;
        RECT 244.400 23.600 245.200 24.400 ;
        RECT 303.600 25.600 304.400 26.400 ;
        RECT 319.600 27.600 320.400 28.400 ;
        RECT 305.200 23.600 306.000 24.400 ;
        RECT 326.000 37.600 326.800 38.400 ;
        RECT 322.800 25.600 323.600 26.400 ;
        RECT 324.400 25.600 325.200 26.400 ;
        RECT 335.600 29.600 336.400 30.400 ;
        RECT 327.600 25.600 328.400 26.400 ;
        RECT 337.200 27.600 338.000 28.400 ;
        RECT 342.000 25.600 342.800 26.400 ;
        RECT 356.400 29.600 357.200 30.400 ;
        RECT 366.000 31.800 366.800 32.600 ;
        RECT 345.200 23.600 346.000 24.400 ;
        RECT 361.200 25.600 362.000 26.400 ;
        RECT 366.000 26.200 366.800 27.000 ;
        RECT 402.600 31.800 403.400 32.600 ;
        RECT 374.000 27.600 374.800 28.400 ;
        RECT 370.800 26.400 371.600 27.200 ;
        RECT 375.600 26.200 376.400 27.000 ;
        RECT 393.200 23.600 394.000 24.400 ;
        RECT 402.600 26.200 403.400 27.000 ;
        RECT 418.800 29.600 419.600 30.400 ;
        RECT 410.800 27.600 411.600 28.400 ;
        RECT 412.400 27.600 413.200 28.400 ;
        RECT 414.000 27.600 414.800 28.400 ;
        RECT 436.400 35.600 437.200 36.400 ;
        RECT 428.400 27.600 429.200 28.400 ;
        RECT 439.600 29.600 440.400 30.400 ;
        RECT 433.200 25.600 434.000 26.400 ;
        RECT 455.600 33.600 456.400 34.400 ;
        RECT 462.000 31.600 462.800 32.400 ;
        RECT 462.000 29.600 462.800 30.400 ;
        RECT 471.600 37.600 472.400 38.400 ;
        RECT 495.600 37.600 496.400 38.400 ;
        RECT 468.400 27.600 469.200 28.400 ;
        RECT 510.000 37.600 510.800 38.400 ;
        RECT 495.600 29.600 496.400 30.400 ;
        RECT 502.000 29.600 502.800 30.400 ;
        RECT 530.800 31.800 531.600 32.600 ;
        RECT 497.200 27.600 498.000 28.400 ;
        RECT 500.400 27.600 501.200 28.400 ;
        RECT 503.600 27.600 504.400 28.400 ;
        RECT 481.200 23.600 482.000 24.400 ;
        RECT 514.800 25.600 515.600 26.400 ;
        RECT 524.400 25.600 525.200 26.400 ;
        RECT 530.800 26.200 531.600 27.000 ;
        RECT 556.400 37.600 557.200 38.400 ;
        RECT 535.600 26.400 536.400 27.200 ;
        RECT 543.600 25.600 544.400 26.400 ;
        RECT 554.800 27.600 555.600 28.400 ;
        RECT 546.800 23.600 547.600 24.400 ;
        RECT 567.600 31.800 568.400 32.600 ;
        RECT 562.800 29.600 563.600 30.400 ;
        RECT 561.200 27.600 562.000 28.400 ;
        RECT 558.000 25.600 558.800 26.400 ;
        RECT 564.400 27.600 565.200 28.400 ;
        RECT 567.600 26.200 568.400 27.000 ;
        RECT 578.800 29.600 579.600 30.400 ;
        RECT 575.600 27.600 576.400 28.400 ;
        RECT 580.400 27.600 581.200 28.400 ;
        RECT 572.400 26.400 573.200 27.200 ;
        RECT 2.800 13.600 3.600 14.400 ;
        RECT 7.600 11.600 8.400 12.400 ;
        RECT 23.600 14.800 24.400 15.600 ;
        RECT 26.800 13.600 27.600 14.400 ;
        RECT 34.800 14.800 35.600 15.600 ;
        RECT 57.200 17.600 58.000 18.400 ;
        RECT 38.000 13.600 38.800 14.400 ;
        RECT 76.400 17.600 77.200 18.400 ;
        RECT 44.400 11.800 45.200 12.600 ;
        RECT 39.600 10.200 40.400 11.000 ;
        RECT 7.600 5.600 8.400 6.400 ;
        RECT 23.600 7.600 24.400 8.400 ;
        RECT 34.800 7.600 35.600 8.400 ;
        RECT 60.400 13.600 61.200 14.400 ;
        RECT 95.600 17.600 96.400 18.400 ;
        RECT 63.600 11.800 64.400 12.600 ;
        RECT 58.800 10.200 59.600 11.000 ;
        RECT 79.600 13.600 80.400 14.400 ;
        RECT 114.800 17.600 115.600 18.400 ;
        RECT 82.800 11.800 83.600 12.600 ;
        RECT 78.000 10.200 78.800 11.000 ;
        RECT 98.800 13.600 99.600 14.400 ;
        RECT 134.000 17.600 134.800 18.400 ;
        RECT 102.000 11.800 102.800 12.600 ;
        RECT 97.200 10.200 98.000 11.000 ;
        RECT 118.000 13.600 118.800 14.400 ;
        RECT 116.400 10.200 117.200 11.000 ;
        RECT 143.600 14.800 144.400 15.600 ;
        RECT 156.400 17.600 157.200 18.400 ;
        RECT 150.000 13.600 150.800 14.400 ;
        RECT 172.400 13.600 173.200 14.400 ;
        RECT 174.000 11.600 174.800 12.400 ;
        RECT 188.400 17.600 189.200 18.400 ;
        RECT 191.600 13.600 192.400 14.400 ;
        RECT 198.000 9.600 198.800 10.400 ;
        RECT 220.400 9.600 221.200 10.400 ;
        RECT 236.400 14.800 237.200 15.600 ;
        RECT 246.000 17.600 246.800 18.400 ;
        RECT 242.800 13.600 243.600 14.400 ;
        RECT 226.800 7.600 227.600 8.400 ;
        RECT 239.600 5.600 240.400 6.400 ;
        RECT 244.400 9.600 245.200 10.400 ;
        RECT 252.400 9.600 253.200 10.400 ;
        RECT 281.200 17.600 282.000 18.400 ;
        RECT 289.200 17.600 290.000 18.400 ;
        RECT 271.600 14.800 272.400 15.600 ;
        RECT 274.800 13.600 275.600 14.400 ;
        RECT 289.200 14.800 290.000 15.600 ;
        RECT 263.600 9.600 264.400 10.400 ;
        RECT 271.600 7.600 272.400 8.400 ;
        RECT 281.200 9.600 282.000 10.400 ;
        RECT 302.000 9.600 302.800 10.400 ;
        RECT 314.800 17.600 315.600 18.400 ;
        RECT 322.800 15.600 323.600 16.400 ;
        RECT 330.800 14.800 331.600 15.600 ;
        RECT 319.600 11.600 320.400 12.400 ;
        RECT 356.400 17.600 357.200 18.400 ;
        RECT 337.200 13.600 338.000 14.400 ;
        RECT 375.600 17.600 376.400 18.400 ;
        RECT 343.600 11.800 344.400 12.600 ;
        RECT 338.800 10.200 339.600 11.000 ;
        RECT 362.800 11.800 363.600 12.600 ;
        RECT 358.000 10.200 358.800 11.000 ;
        RECT 385.200 13.600 386.000 14.400 ;
        RECT 382.000 11.800 382.800 12.600 ;
        RECT 377.200 10.200 378.000 11.000 ;
        RECT 409.200 17.600 410.000 18.400 ;
        RECT 409.200 14.800 410.000 15.600 ;
        RECT 415.600 15.600 416.400 16.400 ;
        RECT 423.600 17.600 424.400 18.400 ;
        RECT 412.400 13.600 413.200 14.400 ;
        RECT 394.800 7.600 395.600 8.400 ;
        RECT 422.000 9.600 422.800 10.400 ;
        RECT 438.000 17.600 438.800 18.400 ;
        RECT 433.200 9.600 434.000 10.400 ;
        RECT 452.400 17.600 453.200 18.400 ;
        RECT 455.600 17.600 456.400 18.400 ;
        RECT 452.400 9.600 453.200 10.400 ;
        RECT 473.200 14.800 474.000 15.600 ;
        RECT 489.200 13.600 490.000 14.400 ;
        RECT 505.200 17.600 506.000 18.400 ;
        RECT 468.400 9.600 469.200 10.400 ;
        RECT 476.400 9.600 477.200 10.400 ;
        RECT 486.000 9.600 486.800 10.400 ;
        RECT 513.200 17.600 514.000 18.400 ;
        RECT 498.800 9.600 499.600 10.400 ;
        RECT 510.000 11.600 510.800 12.400 ;
        RECT 516.400 17.600 517.200 18.400 ;
        RECT 519.600 11.600 520.400 12.400 ;
        RECT 526.000 13.600 526.800 14.400 ;
        RECT 542.000 17.600 542.800 18.400 ;
        RECT 538.800 11.600 539.600 12.400 ;
        RECT 559.600 17.600 560.400 18.400 ;
        RECT 546.800 13.600 547.600 14.400 ;
        RECT 554.800 13.600 555.600 14.400 ;
        RECT 548.400 11.600 549.200 12.400 ;
        RECT 550.000 11.600 550.800 12.400 ;
        RECT 577.200 17.600 578.000 18.400 ;
        RECT 567.600 14.800 568.400 15.600 ;
        RECT 570.800 13.600 571.600 14.400 ;
        RECT 577.200 9.600 578.000 10.400 ;
      LAYER metal2 ;
        RECT 39.600 417.600 40.400 418.400 ;
        RECT 46.000 417.600 46.800 418.400 ;
        RECT 39.700 416.400 40.300 417.600 ;
        RECT 10.800 415.600 11.600 416.400 ;
        RECT 28.400 415.600 29.200 416.400 ;
        RECT 34.800 415.600 35.600 416.400 ;
        RECT 39.600 415.600 40.400 416.400 ;
        RECT 10.900 414.400 11.500 415.600 ;
        RECT 28.500 414.400 29.100 415.600 ;
        RECT 9.200 413.600 10.000 414.400 ;
        RECT 10.800 413.600 11.600 414.400 ;
        RECT 17.200 413.600 18.000 414.400 ;
        RECT 26.800 413.600 27.600 414.400 ;
        RECT 28.400 413.600 29.200 414.400 ;
        RECT 9.300 412.400 9.900 413.600 ;
        RECT 2.800 411.600 3.600 412.400 ;
        RECT 4.400 411.600 5.200 412.400 ;
        RECT 9.200 411.600 10.000 412.400 ;
        RECT 20.400 411.600 21.200 412.400 ;
        RECT 23.600 411.600 24.400 412.400 ;
        RECT 1.200 409.600 2.000 410.400 ;
        RECT 2.900 394.400 3.500 411.600 ;
        RECT 20.500 410.400 21.100 411.600 ;
        RECT 20.400 409.600 21.200 410.400 ;
        RECT 22.000 407.600 22.800 408.400 ;
        RECT 7.600 403.600 8.400 404.400 ;
        RECT 15.600 403.600 16.400 404.400 ;
        RECT 7.700 396.400 8.300 403.600 ;
        RECT 7.600 395.600 8.400 396.400 ;
        RECT 2.800 393.600 3.600 394.400 ;
        RECT 2.900 390.400 3.500 393.600 ;
        RECT 10.800 391.600 11.600 392.400 ;
        RECT 12.400 391.600 13.200 392.400 ;
        RECT 2.800 389.600 3.600 390.400 ;
        RECT 10.900 388.400 11.500 391.600 ;
        RECT 1.200 387.600 2.000 388.400 ;
        RECT 7.600 387.600 8.400 388.400 ;
        RECT 10.800 387.600 11.600 388.400 ;
        RECT 1.300 374.400 1.900 387.600 ;
        RECT 6.000 383.600 6.800 384.400 ;
        RECT 6.100 374.400 6.700 383.600 ;
        RECT 1.200 373.600 2.000 374.400 ;
        RECT 2.800 373.600 3.600 374.400 ;
        RECT 6.000 373.600 6.800 374.400 ;
        RECT 1.200 367.600 2.000 368.400 ;
        RECT 1.300 352.400 1.900 367.600 ;
        RECT 1.200 351.600 2.000 352.400 ;
        RECT 2.900 338.300 3.500 373.600 ;
        RECT 6.000 371.600 6.800 372.400 ;
        RECT 6.100 370.400 6.700 371.600 ;
        RECT 6.000 369.600 6.800 370.400 ;
        RECT 4.400 352.300 5.200 352.400 ;
        RECT 4.400 351.700 6.700 352.300 ;
        RECT 4.400 351.600 5.200 351.700 ;
        RECT 6.100 350.400 6.700 351.700 ;
        RECT 4.400 349.600 5.200 350.400 ;
        RECT 6.000 349.600 6.800 350.400 ;
        RECT 6.000 347.600 6.800 348.400 ;
        RECT 6.100 346.400 6.700 347.600 ;
        RECT 7.700 346.400 8.300 387.600 ;
        RECT 12.500 374.400 13.100 391.600 ;
        RECT 15.700 390.400 16.300 403.600 ;
        RECT 22.100 398.400 22.700 407.600 ;
        RECT 22.000 397.600 22.800 398.400 ;
        RECT 22.000 391.600 22.800 392.400 ;
        RECT 15.600 389.600 16.400 390.400 ;
        RECT 15.600 387.600 16.400 388.400 ;
        RECT 20.400 387.600 21.200 388.400 ;
        RECT 22.000 388.300 22.800 388.400 ;
        RECT 23.700 388.300 24.300 411.600 ;
        RECT 26.900 404.400 27.500 413.600 ;
        RECT 34.900 412.400 35.500 415.600 ;
        RECT 44.400 414.300 45.200 414.400 ;
        RECT 46.100 414.300 46.700 417.600 ;
        RECT 44.400 413.700 46.700 414.300 ;
        RECT 44.400 413.600 45.200 413.700 ;
        RECT 31.600 411.600 32.400 412.400 ;
        RECT 34.800 411.600 35.600 412.400 ;
        RECT 42.800 411.600 43.600 412.400 ;
        RECT 34.800 409.600 35.600 410.400 ;
        RECT 38.000 409.600 38.800 410.400 ;
        RECT 38.100 406.400 38.700 409.600 ;
        RECT 42.900 408.400 43.500 411.600 ;
        RECT 42.800 407.600 43.600 408.400 ;
        RECT 38.000 405.600 38.800 406.400 ;
        RECT 50.800 406.200 51.600 417.800 ;
        RECT 58.800 411.600 59.600 412.600 ;
        RECT 57.200 407.600 58.000 408.400 ;
        RECT 26.800 403.600 27.600 404.400 ;
        RECT 38.000 403.600 38.800 404.400 ;
        RECT 38.100 394.400 38.700 403.600 ;
        RECT 49.200 397.600 50.000 398.400 ;
        RECT 42.800 395.600 43.600 396.400 ;
        RECT 33.200 393.600 34.000 394.400 ;
        RECT 38.000 393.600 38.800 394.400 ;
        RECT 25.200 391.600 26.000 392.400 ;
        RECT 22.000 387.700 24.300 388.300 ;
        RECT 22.000 387.600 22.800 387.700 ;
        RECT 15.700 384.400 16.300 387.600 ;
        RECT 15.600 383.600 16.400 384.400 ;
        RECT 15.700 376.400 16.300 383.600 ;
        RECT 15.600 375.600 16.400 376.400 ;
        RECT 18.800 375.600 19.600 376.400 ;
        RECT 10.800 373.600 11.600 374.400 ;
        RECT 12.400 373.600 13.200 374.400 ;
        RECT 9.200 371.600 10.000 372.400 ;
        RECT 9.300 362.400 9.900 371.600 ;
        RECT 14.000 367.600 14.800 368.400 ;
        RECT 9.200 361.600 10.000 362.400 ;
        RECT 15.700 354.400 16.300 375.600 ;
        RECT 17.200 373.600 18.000 374.400 ;
        RECT 18.900 364.400 19.500 375.600 ;
        RECT 20.500 370.400 21.100 387.600 ;
        RECT 23.600 383.600 24.400 384.400 ;
        RECT 23.700 372.400 24.300 383.600 ;
        RECT 25.300 374.400 25.900 391.600 ;
        RECT 33.300 388.400 33.900 393.600 ;
        RECT 38.100 392.400 38.700 393.600 ;
        RECT 38.000 391.600 38.800 392.400 ;
        RECT 41.200 391.600 42.000 392.400 ;
        RECT 41.200 390.300 42.000 390.400 ;
        RECT 39.700 389.700 42.000 390.300 ;
        RECT 33.200 387.600 34.000 388.400 ;
        RECT 30.000 385.600 30.800 386.400 ;
        RECT 33.200 385.600 34.000 386.400 ;
        RECT 36.400 385.600 37.200 386.400 ;
        RECT 33.300 378.400 33.900 385.600 ;
        RECT 34.800 383.600 35.600 384.400 ;
        RECT 34.900 378.400 35.500 383.600 ;
        RECT 33.200 377.600 34.000 378.400 ;
        RECT 34.800 377.600 35.600 378.400 ;
        RECT 31.600 375.600 32.400 376.400 ;
        RECT 36.400 375.600 37.200 376.400 ;
        RECT 31.700 374.400 32.300 375.600 ;
        RECT 36.500 374.400 37.100 375.600 ;
        RECT 25.200 373.600 26.000 374.400 ;
        RECT 30.000 373.600 30.800 374.400 ;
        RECT 31.600 373.600 32.400 374.400 ;
        RECT 36.400 373.600 37.200 374.400 ;
        RECT 22.000 371.600 22.800 372.400 ;
        RECT 23.600 371.600 24.400 372.400 ;
        RECT 25.200 371.600 26.000 372.400 ;
        RECT 20.400 369.600 21.200 370.400 ;
        RECT 22.100 366.400 22.700 371.600 ;
        RECT 22.000 365.600 22.800 366.400 ;
        RECT 18.800 363.600 19.600 364.400 ;
        RECT 22.000 363.600 22.800 364.400 ;
        RECT 20.400 361.600 21.200 362.400 ;
        RECT 20.500 358.400 21.100 361.600 ;
        RECT 20.400 357.600 21.200 358.400 ;
        RECT 15.600 353.600 16.400 354.400 ;
        RECT 18.800 353.600 19.600 354.400 ;
        RECT 9.000 351.800 9.800 352.600 ;
        RECT 15.600 351.800 16.400 352.600 ;
        RECT 9.000 347.000 9.600 351.800 ;
        RECT 11.600 348.400 12.400 348.600 ;
        RECT 15.800 348.400 16.400 351.800 ;
        RECT 17.200 349.600 18.000 350.400 ;
        RECT 17.300 348.400 17.900 349.600 ;
        RECT 18.900 348.400 19.500 353.600 ;
        RECT 22.100 348.400 22.700 363.600 ;
        RECT 25.300 360.400 25.900 371.600 ;
        RECT 26.800 369.600 27.600 370.400 ;
        RECT 28.400 369.600 29.200 370.400 ;
        RECT 26.900 362.400 27.500 369.600 ;
        RECT 30.100 364.400 30.700 373.600 ;
        RECT 31.600 371.600 32.400 372.400 ;
        RECT 34.800 371.600 35.600 372.400 ;
        RECT 38.000 371.600 38.800 372.400 ;
        RECT 30.000 363.600 30.800 364.400 ;
        RECT 26.800 361.600 27.600 362.400 ;
        RECT 25.200 359.600 26.000 360.400 ;
        RECT 23.400 351.800 24.200 352.600 ;
        RECT 11.600 347.800 16.400 348.400 ;
        RECT 10.800 347.000 11.600 347.200 ;
        RECT 14.200 347.000 15.000 347.200 ;
        RECT 15.800 347.000 16.400 347.800 ;
        RECT 17.200 347.600 18.000 348.400 ;
        RECT 18.800 347.600 19.600 348.400 ;
        RECT 22.000 347.600 22.800 348.400 ;
        RECT 6.000 345.600 6.800 346.400 ;
        RECT 7.600 345.600 8.400 346.400 ;
        RECT 9.000 346.200 9.800 347.000 ;
        RECT 10.800 346.400 15.000 347.000 ;
        RECT 15.600 346.200 16.400 347.000 ;
        RECT 18.900 346.400 19.500 347.600 ;
        RECT 23.400 347.000 24.000 351.800 ;
        RECT 28.400 351.600 29.200 352.400 ;
        RECT 30.000 351.800 30.800 352.600 ;
        RECT 26.000 348.400 26.800 348.600 ;
        RECT 30.200 348.400 30.800 351.800 ;
        RECT 26.000 347.800 30.800 348.400 ;
        RECT 25.200 347.000 26.000 347.200 ;
        RECT 28.600 347.000 29.400 347.200 ;
        RECT 30.200 347.000 30.800 347.800 ;
        RECT 18.800 345.600 19.600 346.400 ;
        RECT 22.000 345.600 22.800 346.400 ;
        RECT 23.400 346.200 24.200 347.000 ;
        RECT 25.200 346.400 29.400 347.000 ;
        RECT 30.000 346.200 30.800 347.000 ;
        RECT 12.400 343.600 13.200 344.400 ;
        RECT 20.400 343.600 21.200 344.400 ;
        RECT 1.300 337.700 3.500 338.300 ;
        RECT 1.300 334.400 1.900 337.700 ;
        RECT 2.600 335.000 3.400 335.800 ;
        RECT 4.400 335.000 8.600 335.600 ;
        RECT 9.200 335.000 10.000 335.800 ;
        RECT 10.800 335.600 11.600 336.400 ;
        RECT 1.200 333.600 2.000 334.400 ;
        RECT 2.600 330.200 3.200 335.000 ;
        RECT 4.400 334.800 5.200 335.000 ;
        RECT 7.800 334.800 8.600 335.000 ;
        RECT 9.400 334.200 10.000 335.000 ;
        RECT 10.900 334.400 11.500 335.600 ;
        RECT 5.200 333.600 10.000 334.200 ;
        RECT 10.800 333.600 11.600 334.400 ;
        RECT 5.200 333.400 6.000 333.600 ;
        RECT 9.400 330.200 10.000 333.600 ;
        RECT 2.600 329.400 3.400 330.200 ;
        RECT 9.200 329.400 10.000 330.200 ;
        RECT 6.000 323.600 6.800 324.400 ;
        RECT 7.600 323.600 8.400 324.400 ;
        RECT 1.200 313.600 2.000 314.400 ;
        RECT 1.300 312.400 1.900 313.600 ;
        RECT 1.200 311.600 2.000 312.400 ;
        RECT 4.400 309.600 5.200 310.400 ;
        RECT 4.500 308.400 5.100 309.600 ;
        RECT 4.400 307.600 5.200 308.400 ;
        RECT 1.200 303.600 2.000 304.400 ;
        RECT 1.300 296.400 1.900 303.600 ;
        RECT 6.100 298.400 6.700 323.600 ;
        RECT 7.700 308.400 8.300 323.600 ;
        RECT 12.500 310.400 13.100 343.600 ;
        RECT 18.800 341.600 19.600 342.400 ;
        RECT 18.900 334.400 19.500 341.600 ;
        RECT 18.800 333.600 19.600 334.400 ;
        RECT 14.000 331.600 14.800 332.400 ;
        RECT 18.900 314.400 19.500 333.600 ;
        RECT 20.500 314.400 21.100 343.600 ;
        RECT 22.100 338.400 22.700 345.600 ;
        RECT 25.200 343.600 26.000 344.400 ;
        RECT 22.000 337.600 22.800 338.400 ;
        RECT 25.300 336.400 25.900 343.600 ;
        RECT 25.200 335.600 26.000 336.400 ;
        RECT 26.800 335.600 27.600 336.400 ;
        RECT 25.200 331.600 26.000 332.400 ;
        RECT 26.900 324.400 27.500 335.600 ;
        RECT 31.700 334.400 32.300 371.600 ;
        RECT 34.900 370.400 35.500 371.600 ;
        RECT 34.800 369.600 35.600 370.400 ;
        RECT 36.400 369.600 37.200 370.400 ;
        RECT 34.800 361.600 35.600 362.400 ;
        RECT 34.900 358.400 35.500 361.600 ;
        RECT 34.800 357.600 35.600 358.400 ;
        RECT 33.200 347.600 34.000 348.400 ;
        RECT 36.500 346.400 37.100 369.600 ;
        RECT 38.100 366.400 38.700 371.600 ;
        RECT 38.000 365.600 38.800 366.400 ;
        RECT 38.100 350.300 38.700 365.600 ;
        RECT 39.700 362.400 40.300 389.700 ;
        RECT 41.200 389.600 42.000 389.700 ;
        RECT 42.900 388.400 43.500 395.600 ;
        RECT 44.400 391.600 45.200 392.400 ;
        RECT 47.600 389.600 48.400 390.400 ;
        RECT 47.700 388.400 48.300 389.600 ;
        RECT 49.300 388.400 49.900 397.600 ;
        RECT 54.000 395.600 54.800 396.400 ;
        RECT 52.400 391.600 53.200 392.400 ;
        RECT 52.500 390.400 53.100 391.600 ;
        RECT 54.100 390.400 54.700 395.600 ;
        RECT 52.400 389.600 53.200 390.400 ;
        RECT 54.000 389.600 54.800 390.400 ;
        RECT 42.800 387.600 43.600 388.400 ;
        RECT 47.600 387.600 48.400 388.400 ;
        RECT 49.200 387.600 50.000 388.400 ;
        RECT 54.000 387.600 54.800 388.400 ;
        RECT 57.300 386.400 57.900 407.600 ;
        RECT 60.400 406.200 61.200 417.800 ;
        RECT 62.000 413.600 62.800 414.400 ;
        RECT 63.600 410.200 64.400 415.800 ;
        RECT 65.200 407.600 66.000 408.400 ;
        RECT 62.000 405.600 62.800 406.400 ;
        RECT 70.000 406.200 70.800 417.800 ;
        RECT 78.000 411.800 78.800 412.600 ;
        RECT 78.100 410.400 78.700 411.800 ;
        RECT 78.000 409.600 78.800 410.400 ;
        RECT 79.600 406.200 80.400 417.800 ;
        RECT 81.200 413.600 82.000 414.400 ;
        RECT 82.800 410.200 83.600 415.800 ;
        RECT 84.400 413.600 85.200 414.400 ;
        RECT 98.800 413.600 99.600 414.400 ;
        RECT 62.100 390.400 62.700 405.600 ;
        RECT 76.400 393.600 77.200 394.400 ;
        RECT 66.800 391.800 67.600 392.600 ;
        RECT 73.000 391.800 73.800 392.600 ;
        RECT 62.000 389.600 62.800 390.400 ;
        RECT 63.600 389.600 64.400 390.400 ;
        RECT 62.100 388.400 62.700 389.600 ;
        RECT 63.700 388.400 64.300 389.600 ;
        RECT 66.800 388.400 67.400 391.800 ;
        RECT 71.800 389.800 72.600 390.600 ;
        RECT 71.800 388.400 72.400 389.800 ;
        RECT 62.000 387.600 62.800 388.400 ;
        RECT 63.600 387.600 64.400 388.400 ;
        RECT 66.800 387.800 72.400 388.400 ;
        RECT 66.800 387.000 67.400 387.800 ;
        RECT 68.200 387.000 69.000 387.200 ;
        RECT 71.600 387.000 72.400 387.200 ;
        RECT 73.200 387.000 73.800 391.800 ;
        RECT 74.800 387.600 75.600 388.400 ;
        RECT 41.200 385.600 42.000 386.400 ;
        RECT 57.200 385.600 58.000 386.400 ;
        RECT 66.800 386.200 67.600 387.000 ;
        RECT 68.200 386.400 73.800 387.000 ;
        RECT 76.500 386.400 77.100 393.600 ;
        RECT 79.600 391.600 80.400 392.400 ;
        RECT 79.700 388.400 80.300 391.600 ;
        RECT 79.600 387.600 80.400 388.400 ;
        RECT 82.800 387.600 83.600 388.400 ;
        RECT 73.000 386.200 73.800 386.400 ;
        RECT 76.400 385.600 77.200 386.400 ;
        RECT 41.300 378.400 41.900 385.600 ;
        RECT 44.400 383.600 45.200 384.400 ;
        RECT 60.400 383.600 61.200 384.400 ;
        RECT 70.000 383.600 70.800 384.400 ;
        RECT 41.200 377.600 42.000 378.400 ;
        RECT 42.800 369.600 43.600 370.400 ;
        RECT 42.900 368.400 43.500 369.600 ;
        RECT 42.800 367.600 43.600 368.400 ;
        RECT 39.600 361.600 40.400 362.400 ;
        RECT 42.900 354.400 43.500 367.600 ;
        RECT 42.800 353.600 43.600 354.400 ;
        RECT 38.100 349.700 40.300 350.300 ;
        RECT 38.000 347.600 38.800 348.400 ;
        RECT 33.200 345.600 34.000 346.400 ;
        RECT 36.400 345.600 37.200 346.400 ;
        RECT 36.500 344.400 37.100 345.600 ;
        RECT 34.800 343.600 35.600 344.400 ;
        RECT 36.400 343.600 37.200 344.400 ;
        RECT 31.600 333.600 32.400 334.400 ;
        RECT 30.000 331.600 30.800 332.400 ;
        RECT 28.400 329.600 29.200 330.400 ;
        RECT 28.500 324.400 29.100 329.600 ;
        RECT 22.000 323.600 22.800 324.400 ;
        RECT 26.800 323.600 27.600 324.400 ;
        RECT 28.400 323.600 29.200 324.400 ;
        RECT 18.800 313.600 19.600 314.400 ;
        RECT 20.400 313.600 21.200 314.400 ;
        RECT 22.100 312.400 22.700 323.600 ;
        RECT 22.000 311.600 22.800 312.400 ;
        RECT 25.200 311.600 26.000 312.400 ;
        RECT 28.500 310.400 29.100 323.600 ;
        RECT 30.100 312.400 30.700 331.600 ;
        RECT 33.200 323.600 34.000 324.400 ;
        RECT 31.600 313.600 32.400 314.400 ;
        RECT 31.700 312.400 32.300 313.600 ;
        RECT 30.000 311.600 30.800 312.400 ;
        RECT 31.600 311.600 32.400 312.400 ;
        RECT 10.800 309.600 11.600 310.400 ;
        RECT 12.400 309.600 13.200 310.400 ;
        RECT 15.600 309.600 16.400 310.400 ;
        RECT 20.400 309.600 21.200 310.400 ;
        RECT 28.400 309.600 29.200 310.400 ;
        RECT 10.900 308.400 11.500 309.600 ;
        RECT 7.600 307.600 8.400 308.400 ;
        RECT 10.800 307.600 11.600 308.400 ;
        RECT 6.000 297.600 6.800 298.400 ;
        RECT 1.200 295.600 2.000 296.400 ;
        RECT 6.000 295.600 6.800 296.400 ;
        RECT 1.300 266.400 1.900 295.600 ;
        RECT 2.800 289.600 3.600 290.400 ;
        RECT 7.600 289.600 8.400 290.400 ;
        RECT 10.900 286.400 11.500 307.600 ;
        RECT 15.700 306.400 16.300 309.600 ;
        RECT 17.200 307.600 18.000 308.400 ;
        RECT 26.800 307.600 27.600 308.400 ;
        RECT 12.400 305.600 13.200 306.400 ;
        RECT 15.600 305.600 16.400 306.400 ;
        RECT 20.400 305.600 21.200 306.400 ;
        RECT 23.600 305.600 24.400 306.400 ;
        RECT 12.500 296.400 13.100 305.600 ;
        RECT 14.000 303.600 14.800 304.400 ;
        RECT 14.100 296.400 14.700 303.600 ;
        RECT 22.000 299.600 22.800 300.400 ;
        RECT 12.400 295.600 13.200 296.400 ;
        RECT 14.000 295.600 14.800 296.400 ;
        RECT 20.400 295.600 21.200 296.400 ;
        RECT 12.500 294.400 13.100 295.600 ;
        RECT 12.400 293.600 13.200 294.400 ;
        RECT 12.400 291.600 13.200 292.400 ;
        RECT 12.500 286.400 13.100 291.600 ;
        RECT 7.600 285.600 8.400 286.400 ;
        RECT 10.800 285.600 11.600 286.400 ;
        RECT 12.400 285.600 13.200 286.400 ;
        RECT 4.400 283.600 5.200 284.400 ;
        RECT 4.500 268.400 5.100 283.600 ;
        RECT 6.000 269.600 6.800 270.400 ;
        RECT 4.400 267.600 5.200 268.400 ;
        RECT 1.200 265.600 2.000 266.400 ;
        RECT 6.100 264.400 6.700 269.600 ;
        RECT 7.700 268.400 8.300 285.600 ;
        RECT 10.800 283.600 11.600 284.400 ;
        RECT 9.200 271.800 10.000 272.600 ;
        RECT 14.100 272.400 14.700 295.600 ;
        RECT 20.500 294.400 21.100 295.600 ;
        RECT 20.400 293.600 21.200 294.400 ;
        RECT 22.100 292.400 22.700 299.600 ;
        RECT 26.900 296.300 27.500 307.600 ;
        RECT 28.500 306.400 29.100 309.600 ;
        RECT 33.300 308.400 33.900 323.600 ;
        RECT 34.900 308.400 35.500 343.600 ;
        RECT 38.100 340.400 38.700 347.600 ;
        RECT 38.000 339.600 38.800 340.400 ;
        RECT 38.000 334.300 38.800 334.400 ;
        RECT 39.700 334.300 40.300 349.700 ;
        RECT 41.200 349.600 42.000 350.400 ;
        RECT 44.500 346.400 45.100 383.600 ;
        RECT 47.600 373.600 48.400 374.400 ;
        RECT 46.000 371.600 46.800 372.400 ;
        RECT 46.100 370.400 46.700 371.600 ;
        RECT 46.000 369.600 46.800 370.400 ;
        RECT 47.700 362.400 48.300 373.600 ;
        RECT 54.000 366.200 54.800 377.800 ;
        RECT 49.200 363.600 50.000 364.400 ;
        RECT 47.600 361.600 48.400 362.400 ;
        RECT 49.300 354.300 49.900 363.600 ;
        RECT 54.000 361.600 54.800 362.400 ;
        RECT 47.700 353.700 49.900 354.300 ;
        RECT 47.700 350.400 48.300 353.700 ;
        RECT 49.200 351.600 50.000 352.400 ;
        RECT 47.600 349.600 48.400 350.400 ;
        RECT 46.000 347.600 46.800 348.400 ;
        RECT 42.800 345.600 43.600 346.400 ;
        RECT 44.400 345.600 45.200 346.400 ;
        RECT 47.600 345.600 48.400 346.400 ;
        RECT 42.900 344.400 43.500 345.600 ;
        RECT 42.800 343.600 43.600 344.400 ;
        RECT 44.400 343.600 45.200 344.400 ;
        RECT 38.000 333.700 40.300 334.300 ;
        RECT 38.000 333.600 38.800 333.700 ;
        RECT 41.200 333.600 42.000 334.400 ;
        RECT 44.500 332.400 45.100 343.600 ;
        RECT 47.700 332.400 48.300 345.600 ;
        RECT 49.300 334.400 49.900 351.600 ;
        RECT 52.400 349.600 53.200 350.400 ;
        RECT 50.800 347.600 51.600 348.400 ;
        RECT 52.500 344.400 53.100 349.600 ;
        RECT 54.100 348.400 54.700 361.600 ;
        RECT 60.500 360.400 61.100 383.600 ;
        RECT 62.000 371.600 62.800 372.600 ;
        RECT 63.600 366.200 64.400 377.800 ;
        RECT 65.200 373.600 66.000 374.400 ;
        RECT 66.800 370.200 67.600 375.800 ;
        RECT 68.400 369.600 69.200 370.400 ;
        RECT 57.200 359.600 58.000 360.400 ;
        RECT 60.400 359.600 61.200 360.400 ;
        RECT 57.300 350.400 57.900 359.600 ;
        RECT 63.600 353.600 64.400 354.400 ;
        RECT 60.400 351.600 61.200 352.400 ;
        RECT 57.200 349.600 58.000 350.400 ;
        RECT 62.000 349.600 62.800 350.400 ;
        RECT 63.700 348.400 64.300 353.600 ;
        RECT 65.200 351.600 66.000 352.400 ;
        RECT 65.300 350.400 65.900 351.600 ;
        RECT 65.200 349.600 66.000 350.400 ;
        RECT 68.400 349.600 69.200 350.400 ;
        RECT 54.000 347.600 54.800 348.400 ;
        RECT 55.600 347.600 56.400 348.400 ;
        RECT 62.000 347.600 62.800 348.400 ;
        RECT 63.600 347.600 64.400 348.400 ;
        RECT 52.400 343.600 53.200 344.400 ;
        RECT 54.100 340.400 54.700 347.600 ;
        RECT 60.400 345.600 61.200 346.400 ;
        RECT 54.000 339.600 54.800 340.400 ;
        RECT 58.800 339.600 59.600 340.400 ;
        RECT 58.900 336.400 59.500 339.600 ;
        RECT 60.500 336.400 61.100 345.600 ;
        RECT 68.500 344.400 69.100 349.600 ;
        RECT 68.400 343.600 69.200 344.400 ;
        RECT 58.800 335.600 59.600 336.400 ;
        RECT 60.400 335.600 61.200 336.400 ;
        RECT 49.200 333.600 50.000 334.400 ;
        RECT 36.400 331.600 37.200 332.400 ;
        RECT 44.400 331.600 45.200 332.400 ;
        RECT 47.600 331.600 48.400 332.400 ;
        RECT 54.000 331.600 54.800 332.400 ;
        RECT 36.500 330.400 37.100 331.600 ;
        RECT 44.500 330.400 45.100 331.600 ;
        RECT 54.100 330.400 54.700 331.600 ;
        RECT 36.400 329.600 37.200 330.400 ;
        RECT 44.400 329.600 45.200 330.400 ;
        RECT 54.000 329.600 54.800 330.400 ;
        RECT 47.600 327.600 48.400 328.400 ;
        RECT 52.400 327.600 53.200 328.400 ;
        RECT 41.200 325.600 42.000 326.400 ;
        RECT 41.300 324.400 41.900 325.600 ;
        RECT 41.200 323.600 42.000 324.400 ;
        RECT 54.000 323.600 54.800 324.400 ;
        RECT 41.300 314.400 41.900 323.600 ;
        RECT 52.400 317.600 53.200 318.400 ;
        RECT 41.200 313.600 42.000 314.400 ;
        RECT 44.400 313.600 45.200 314.400 ;
        RECT 44.500 312.400 45.100 313.600 ;
        RECT 44.400 311.600 45.200 312.400 ;
        RECT 49.200 312.300 50.000 312.400 ;
        RECT 49.200 311.700 51.500 312.300 ;
        RECT 49.200 311.600 50.000 311.700 ;
        RECT 50.900 310.400 51.500 311.700 ;
        RECT 36.400 309.600 37.200 310.400 ;
        RECT 49.200 309.600 50.000 310.400 ;
        RECT 50.800 309.600 51.600 310.400 ;
        RECT 30.000 307.600 30.800 308.400 ;
        RECT 33.200 307.600 34.000 308.400 ;
        RECT 34.800 307.600 35.600 308.400 ;
        RECT 28.400 305.600 29.200 306.400 ;
        RECT 28.400 296.300 29.200 296.400 ;
        RECT 26.900 295.700 29.200 296.300 ;
        RECT 25.200 293.600 26.000 294.400 ;
        RECT 17.200 291.600 18.000 292.400 ;
        RECT 22.000 291.600 22.800 292.400 ;
        RECT 23.600 291.600 24.400 292.400 ;
        RECT 18.800 289.600 19.600 290.400 ;
        RECT 15.600 287.600 16.400 288.400 ;
        RECT 15.700 284.400 16.300 287.600 ;
        RECT 15.600 283.600 16.400 284.400 ;
        RECT 17.200 283.600 18.000 284.400 ;
        RECT 9.200 268.400 9.800 271.800 ;
        RECT 14.000 271.600 14.800 272.400 ;
        RECT 15.400 271.800 16.200 272.600 ;
        RECT 14.200 269.800 15.000 270.600 ;
        RECT 14.200 268.400 14.800 269.800 ;
        RECT 7.600 267.600 8.400 268.400 ;
        RECT 9.200 267.800 14.800 268.400 ;
        RECT 9.200 267.000 9.800 267.800 ;
        RECT 10.600 267.000 11.400 267.200 ;
        RECT 14.000 267.000 14.800 267.200 ;
        RECT 15.600 267.000 16.200 271.800 ;
        RECT 17.300 270.400 17.900 283.600 ;
        RECT 18.900 278.400 19.500 289.600 ;
        RECT 18.800 277.600 19.600 278.400 ;
        RECT 18.900 274.400 19.500 277.600 ;
        RECT 18.800 273.600 19.600 274.400 ;
        RECT 22.000 273.600 22.800 274.400 ;
        RECT 22.100 272.400 22.700 273.600 ;
        RECT 22.000 271.600 22.800 272.400 ;
        RECT 23.600 271.600 24.400 272.400 ;
        RECT 17.200 269.600 18.000 270.400 ;
        RECT 20.400 269.600 21.200 270.400 ;
        RECT 17.200 267.600 18.000 268.400 ;
        RECT 9.200 266.200 10.000 267.000 ;
        RECT 10.600 266.400 16.200 267.000 ;
        RECT 15.400 266.200 16.200 266.400 ;
        RECT 18.800 265.600 19.600 266.400 ;
        RECT 2.800 263.600 3.600 264.400 ;
        RECT 6.000 263.600 6.800 264.400 ;
        RECT 12.400 263.600 13.200 264.400 ;
        RECT 1.200 253.600 2.000 254.400 ;
        RECT 2.900 252.400 3.500 263.600 ;
        RECT 6.000 261.600 6.800 262.400 ;
        RECT 2.800 251.600 3.600 252.400 ;
        RECT 6.100 250.400 6.700 261.600 ;
        RECT 10.800 257.600 11.600 258.400 ;
        RECT 10.900 254.400 11.500 257.600 ;
        RECT 12.500 254.400 13.100 263.600 ;
        RECT 18.900 262.400 19.500 265.600 ;
        RECT 18.800 261.600 19.600 262.400 ;
        RECT 14.000 259.600 14.800 260.400 ;
        RECT 10.800 253.600 11.600 254.400 ;
        RECT 12.400 253.600 13.200 254.400 ;
        RECT 6.000 249.600 6.800 250.400 ;
        RECT 9.200 243.600 10.000 244.400 ;
        RECT 1.200 223.600 2.000 224.400 ;
        RECT 6.000 224.200 6.800 235.800 ;
        RECT 1.200 210.200 2.000 215.800 ;
        RECT 4.400 206.200 5.200 217.800 ;
        RECT 6.000 211.600 6.800 212.600 ;
        RECT 1.200 186.200 2.000 191.800 ;
        RECT 2.800 183.600 3.600 184.400 ;
        RECT 4.400 184.200 5.200 195.800 ;
        RECT 9.300 190.400 9.900 243.600 ;
        RECT 14.100 230.200 14.700 259.600 ;
        RECT 20.500 258.400 21.100 269.600 ;
        RECT 22.000 263.600 22.800 264.400 ;
        RECT 20.400 257.600 21.200 258.400 ;
        RECT 22.100 256.400 22.700 263.600 ;
        RECT 23.700 256.400 24.300 271.600 ;
        RECT 15.600 255.600 16.400 256.400 ;
        RECT 18.800 255.600 19.600 256.400 ;
        RECT 22.000 255.600 22.800 256.400 ;
        RECT 23.600 255.600 24.400 256.400 ;
        RECT 18.900 252.400 19.500 255.600 ;
        RECT 20.400 253.600 21.200 254.400 ;
        RECT 22.000 253.600 22.800 254.400 ;
        RECT 18.800 251.600 19.600 252.400 ;
        RECT 15.600 249.600 16.400 250.400 ;
        RECT 14.000 229.400 14.800 230.200 ;
        RECT 12.400 227.600 13.200 228.400 ;
        RECT 12.500 214.400 13.100 227.600 ;
        RECT 15.600 224.200 16.400 235.800 ;
        RECT 18.800 226.200 19.600 231.800 ;
        RECT 20.500 228.400 21.100 253.600 ;
        RECT 25.300 252.400 25.900 293.600 ;
        RECT 26.900 272.400 27.500 295.700 ;
        RECT 28.400 295.600 29.200 295.700 ;
        RECT 30.100 292.400 30.700 307.600 ;
        RECT 34.900 306.400 35.500 307.600 ;
        RECT 34.800 305.600 35.600 306.400 ;
        RECT 33.200 303.600 34.000 304.400 ;
        RECT 33.300 302.400 33.900 303.600 ;
        RECT 33.200 301.600 34.000 302.400 ;
        RECT 36.500 298.400 37.100 309.600 ;
        RECT 41.200 307.600 42.000 308.400 ;
        RECT 50.800 307.600 51.600 308.400 ;
        RECT 39.600 305.600 40.400 306.400 ;
        RECT 38.000 303.600 38.800 304.400 ;
        RECT 31.600 297.600 32.400 298.400 ;
        RECT 36.400 297.600 37.200 298.400 ;
        RECT 28.400 291.600 29.200 292.400 ;
        RECT 30.000 291.600 30.800 292.400 ;
        RECT 28.500 274.400 29.100 291.600 ;
        RECT 30.000 290.300 30.800 290.400 ;
        RECT 31.700 290.300 32.300 297.600 ;
        RECT 34.800 295.600 35.600 296.400 ;
        RECT 36.400 295.600 37.200 296.400 ;
        RECT 34.900 294.400 35.500 295.600 ;
        RECT 36.500 294.400 37.100 295.600 ;
        RECT 34.800 293.600 35.600 294.400 ;
        RECT 36.400 293.600 37.200 294.400 ;
        RECT 33.200 291.600 34.000 292.400 ;
        RECT 33.300 290.400 33.900 291.600 ;
        RECT 30.000 289.700 32.300 290.300 ;
        RECT 30.000 289.600 30.800 289.700 ;
        RECT 33.200 289.600 34.000 290.400 ;
        RECT 30.000 287.600 30.800 288.400 ;
        RECT 30.100 278.400 30.700 287.600 ;
        RECT 30.000 277.600 30.800 278.400 ;
        RECT 28.400 273.600 29.200 274.400 ;
        RECT 26.800 271.600 27.600 272.400 ;
        RECT 31.600 271.600 32.400 272.400 ;
        RECT 26.800 269.600 27.600 270.400 ;
        RECT 33.300 268.400 33.900 289.600 ;
        RECT 36.400 283.600 37.200 284.400 ;
        RECT 34.800 279.600 35.600 280.400 ;
        RECT 34.900 270.400 35.500 279.600 ;
        RECT 36.500 272.400 37.100 283.600 ;
        RECT 36.400 271.600 37.200 272.400 ;
        RECT 34.800 269.600 35.600 270.400 ;
        RECT 33.200 267.600 34.000 268.400 ;
        RECT 36.400 267.600 37.200 268.400 ;
        RECT 38.100 266.400 38.700 303.600 ;
        RECT 44.400 301.600 45.200 302.400 ;
        RECT 41.200 297.600 42.000 298.400 ;
        RECT 39.600 295.600 40.400 296.400 ;
        RECT 39.700 294.400 40.300 295.600 ;
        RECT 39.600 293.600 40.400 294.400 ;
        RECT 41.300 292.400 41.900 297.600 ;
        RECT 44.500 294.400 45.100 301.600 ;
        RECT 46.000 299.600 46.800 300.400 ;
        RECT 47.600 299.600 48.400 300.400 ;
        RECT 46.100 298.400 46.700 299.600 ;
        RECT 46.000 297.600 46.800 298.400 ;
        RECT 47.700 294.400 48.300 299.600 ;
        RECT 50.900 298.400 51.500 307.600 ;
        RECT 50.800 297.600 51.600 298.400 ;
        RECT 50.800 295.600 51.600 296.400 ;
        RECT 50.900 294.400 51.500 295.600 ;
        RECT 44.400 293.600 45.200 294.400 ;
        RECT 47.600 293.600 48.400 294.400 ;
        RECT 50.800 293.600 51.600 294.400 ;
        RECT 41.200 291.600 42.000 292.400 ;
        RECT 42.800 273.600 43.600 274.400 ;
        RECT 42.900 270.400 43.500 273.600 ;
        RECT 42.800 269.600 43.600 270.400 ;
        RECT 41.200 267.600 42.000 268.400 ;
        RECT 44.500 268.300 45.100 293.600 ;
        RECT 52.500 292.400 53.100 317.600 ;
        RECT 54.100 314.400 54.700 323.600 ;
        RECT 54.000 313.600 54.800 314.400 ;
        RECT 60.500 314.300 61.100 335.600 ;
        RECT 70.100 332.400 70.700 383.600 ;
        RECT 73.200 375.600 74.000 376.400 ;
        RECT 73.300 374.400 73.900 375.600 ;
        RECT 73.200 373.600 74.000 374.400 ;
        RECT 76.400 373.600 77.200 374.400 ;
        RECT 71.600 371.600 72.400 372.400 ;
        RECT 73.300 368.400 73.900 373.600 ;
        RECT 76.500 372.400 77.100 373.600 ;
        RECT 76.400 371.600 77.200 372.400 ;
        RECT 73.200 367.600 74.000 368.400 ;
        RECT 73.300 346.400 73.900 367.600 ;
        RECT 76.500 366.400 77.100 371.600 ;
        RECT 74.800 365.600 75.600 366.400 ;
        RECT 76.400 365.600 77.200 366.400 ;
        RECT 74.900 364.400 75.500 365.600 ;
        RECT 74.800 363.600 75.600 364.400 ;
        RECT 74.900 350.400 75.500 363.600 ;
        RECT 76.500 350.400 77.100 365.600 ;
        RECT 78.000 363.600 78.800 364.400 ;
        RECT 74.800 349.600 75.600 350.400 ;
        RECT 76.400 349.600 77.200 350.400 ;
        RECT 78.000 349.600 78.800 350.400 ;
        RECT 78.100 348.400 78.700 349.600 ;
        RECT 76.400 347.600 77.200 348.400 ;
        RECT 78.000 347.600 78.800 348.400 ;
        RECT 76.500 346.400 77.100 347.600 ;
        RECT 73.200 345.600 74.000 346.400 ;
        RECT 76.400 345.600 77.200 346.400 ;
        RECT 74.800 343.600 75.600 344.400 ;
        RECT 74.900 340.400 75.500 343.600 ;
        RECT 79.700 342.400 80.300 387.600 ;
        RECT 82.800 366.200 83.600 377.800 ;
        RECT 84.500 374.400 85.100 413.600 ;
        RECT 98.900 406.400 99.500 413.600 ;
        RECT 98.800 405.600 99.600 406.400 ;
        RECT 108.400 406.200 109.200 417.800 ;
        RECT 110.000 413.600 110.800 414.400 ;
        RECT 110.100 412.400 110.700 413.600 ;
        RECT 110.000 411.600 110.800 412.400 ;
        RECT 116.400 411.800 117.200 412.600 ;
        RECT 86.000 391.600 86.800 392.400 ;
        RECT 89.200 391.600 90.000 392.400 ;
        RECT 92.400 391.600 93.200 392.400 ;
        RECT 97.200 391.600 98.000 392.400 ;
        RECT 89.300 390.400 89.900 391.600 ;
        RECT 92.500 390.400 93.100 391.600 ;
        RECT 89.200 389.600 90.000 390.400 ;
        RECT 92.400 389.600 93.200 390.400 ;
        RECT 98.900 388.400 99.500 405.600 ;
        RECT 100.400 403.600 101.200 404.400 ;
        RECT 103.600 403.600 104.400 404.400 ;
        RECT 100.500 394.400 101.100 403.600 ;
        RECT 100.400 393.600 101.200 394.400 ;
        RECT 103.700 388.400 104.300 403.600 ;
        RECT 108.400 391.600 109.200 392.400 ;
        RECT 105.200 389.600 106.000 390.400 ;
        RECT 92.400 387.600 93.200 388.400 ;
        RECT 98.800 387.600 99.600 388.400 ;
        RECT 100.400 387.600 101.200 388.400 ;
        RECT 103.600 387.600 104.400 388.400 ;
        RECT 108.400 387.600 109.200 388.400 ;
        RECT 94.000 383.600 94.800 384.400 ;
        RECT 84.400 373.600 85.200 374.400 ;
        RECT 84.500 372.400 85.100 373.600 ;
        RECT 84.400 371.600 85.200 372.400 ;
        RECT 90.800 371.600 91.600 372.600 ;
        RECT 92.400 366.200 93.200 377.800 ;
        RECT 94.100 372.400 94.700 383.600 ;
        RECT 94.000 371.600 94.800 372.400 ;
        RECT 95.600 370.200 96.400 375.800 ;
        RECT 97.200 367.600 98.000 368.400 ;
        RECT 100.400 367.600 101.200 368.400 ;
        RECT 87.600 352.300 88.400 352.400 ;
        RECT 86.100 351.700 88.400 352.300 ;
        RECT 82.800 345.600 83.600 346.400 ;
        RECT 84.400 345.600 85.200 346.400 ;
        RECT 81.200 343.600 82.000 344.400 ;
        RECT 79.600 341.600 80.400 342.400 ;
        RECT 74.800 339.600 75.600 340.400 ;
        RECT 81.300 338.400 81.900 343.600 ;
        RECT 82.900 338.400 83.500 345.600 ;
        RECT 78.000 337.600 78.800 338.400 ;
        RECT 81.200 337.600 82.000 338.400 ;
        RECT 82.800 337.600 83.600 338.400 ;
        RECT 71.600 335.600 72.400 336.400 ;
        RECT 71.700 332.400 72.300 335.600 ;
        RECT 78.100 332.400 78.700 337.600 ;
        RECT 81.200 335.600 82.000 336.400 ;
        RECT 81.300 334.400 81.900 335.600 ;
        RECT 79.600 333.600 80.400 334.400 ;
        RECT 81.200 333.600 82.000 334.400 ;
        RECT 70.000 331.600 70.800 332.400 ;
        RECT 71.600 331.600 72.400 332.400 ;
        RECT 78.000 331.600 78.800 332.400 ;
        RECT 66.800 329.600 67.600 330.400 ;
        RECT 71.600 329.600 72.400 330.400 ;
        RECT 73.200 329.600 74.000 330.400 ;
        RECT 74.800 329.600 75.600 330.400 ;
        RECT 65.200 327.600 66.000 328.400 ;
        RECT 66.900 326.400 67.500 329.600 ;
        RECT 70.000 327.600 70.800 328.400 ;
        RECT 71.700 326.400 72.300 329.600 ;
        RECT 66.800 325.600 67.600 326.400 ;
        RECT 71.600 325.600 72.400 326.400 ;
        RECT 68.400 315.600 69.200 316.400 ;
        RECT 60.500 313.700 62.700 314.300 ;
        RECT 53.800 311.800 54.600 312.600 ;
        RECT 60.400 311.800 61.200 312.600 ;
        RECT 53.800 307.000 54.400 311.800 ;
        RECT 56.400 308.400 57.200 308.600 ;
        RECT 60.600 308.400 61.200 311.800 ;
        RECT 62.100 308.400 62.700 313.700 ;
        RECT 63.600 313.600 64.400 314.400 ;
        RECT 66.800 313.600 67.600 314.400 ;
        RECT 63.700 312.400 64.300 313.600 ;
        RECT 63.600 311.600 64.400 312.400 ;
        RECT 56.400 307.800 61.200 308.400 ;
        RECT 55.600 307.000 56.400 307.200 ;
        RECT 59.000 307.000 59.800 307.200 ;
        RECT 60.600 307.000 61.200 307.800 ;
        RECT 62.000 307.600 62.800 308.400 ;
        RECT 53.800 306.200 54.600 307.000 ;
        RECT 55.600 306.400 59.800 307.000 ;
        RECT 60.400 306.200 61.200 307.000 ;
        RECT 55.600 303.600 56.400 304.400 ;
        RECT 55.700 294.300 56.300 303.600 ;
        RECT 62.100 296.400 62.700 307.600 ;
        RECT 65.200 303.600 66.000 304.400 ;
        RECT 66.900 298.400 67.500 313.600 ;
        RECT 68.500 308.400 69.100 315.600 ;
        RECT 73.300 314.400 73.900 329.600 ;
        RECT 78.000 323.600 78.800 324.400 ;
        RECT 74.800 319.600 75.600 320.400 ;
        RECT 74.900 318.400 75.500 319.600 ;
        RECT 74.800 317.600 75.600 318.400 ;
        RECT 73.200 313.600 74.000 314.400 ;
        RECT 71.600 311.600 72.400 312.400 ;
        RECT 71.700 310.400 72.300 311.600 ;
        RECT 71.600 309.600 72.400 310.400 ;
        RECT 76.400 310.300 77.200 310.400 ;
        RECT 73.300 309.700 77.200 310.300 ;
        RECT 68.400 307.600 69.200 308.400 ;
        RECT 70.000 308.300 70.800 308.400 ;
        RECT 73.300 308.300 73.900 309.700 ;
        RECT 76.400 309.600 77.200 309.700 ;
        RECT 70.000 307.700 73.900 308.300 ;
        RECT 70.000 307.600 70.800 307.700 ;
        RECT 76.400 307.600 77.200 308.400 ;
        RECT 68.400 305.600 69.200 306.400 ;
        RECT 68.500 302.400 69.100 305.600 ;
        RECT 71.600 303.600 72.400 304.400 ;
        RECT 68.400 301.600 69.200 302.400 ;
        RECT 63.600 297.600 64.400 298.400 ;
        RECT 66.800 297.600 67.600 298.400 ;
        RECT 62.000 295.600 62.800 296.400 ;
        RECT 63.700 294.400 64.300 297.600 ;
        RECT 54.100 293.700 56.300 294.300 ;
        RECT 49.200 291.600 50.000 292.400 ;
        RECT 52.400 291.600 53.200 292.400 ;
        RECT 49.300 288.400 49.900 291.600 ;
        RECT 52.500 290.400 53.100 291.600 ;
        RECT 52.400 289.600 53.200 290.400 ;
        RECT 49.200 287.600 50.000 288.400 ;
        RECT 47.600 275.600 48.400 276.400 ;
        RECT 47.700 270.400 48.300 275.600 ;
        RECT 52.400 273.600 53.200 274.400 ;
        RECT 47.600 269.600 48.400 270.400 ;
        RECT 52.500 268.400 53.100 273.600 ;
        RECT 46.000 268.300 46.800 268.400 ;
        RECT 44.500 267.700 46.800 268.300 ;
        RECT 46.000 267.600 46.800 267.700 ;
        RECT 52.400 267.600 53.200 268.400 ;
        RECT 28.400 265.600 29.200 266.400 ;
        RECT 38.000 265.600 38.800 266.400 ;
        RECT 41.200 265.600 42.000 266.400 ;
        RECT 46.000 265.600 46.800 266.400 ;
        RECT 47.600 265.600 48.400 266.400 ;
        RECT 31.600 263.600 32.400 264.400 ;
        RECT 33.200 263.600 34.000 264.400 ;
        RECT 39.600 263.600 40.400 264.400 ;
        RECT 26.800 255.600 27.600 256.400 ;
        RECT 26.900 252.400 27.500 255.600 ;
        RECT 31.700 252.400 32.300 263.600 ;
        RECT 33.300 256.400 33.900 263.600 ;
        RECT 33.200 255.600 34.000 256.400 ;
        RECT 39.700 256.300 40.300 263.600 ;
        RECT 41.300 258.400 41.900 265.600 ;
        RECT 46.100 264.400 46.700 265.600 ;
        RECT 46.000 263.600 46.800 264.400 ;
        RECT 41.200 257.600 42.000 258.400 ;
        RECT 38.100 255.700 40.300 256.300 ;
        RECT 33.300 252.400 33.900 255.600 ;
        RECT 38.100 252.400 38.700 255.700 ;
        RECT 46.100 254.400 46.700 263.600 ;
        RECT 47.700 258.400 48.300 265.600 ;
        RECT 49.200 263.600 50.000 264.400 ;
        RECT 50.800 263.600 51.600 264.400 ;
        RECT 47.600 257.600 48.400 258.400 ;
        RECT 49.300 256.400 49.900 263.600 ;
        RECT 50.900 256.400 51.500 263.600 ;
        RECT 54.100 260.400 54.700 293.700 ;
        RECT 62.000 293.600 62.800 294.400 ;
        RECT 63.600 293.600 64.400 294.400 ;
        RECT 68.400 293.600 69.200 294.400 ;
        RECT 62.100 292.400 62.700 293.600 ;
        RECT 55.600 291.600 56.400 292.400 ;
        RECT 57.200 291.600 58.000 292.400 ;
        RECT 62.000 291.600 62.800 292.400 ;
        RECT 65.200 291.600 66.000 292.400 ;
        RECT 55.700 290.400 56.300 291.600 ;
        RECT 55.600 289.600 56.400 290.400 ;
        RECT 55.700 276.400 56.300 289.600 ;
        RECT 57.300 278.400 57.900 291.600 ;
        RECT 60.400 285.600 61.200 286.400 ;
        RECT 65.200 283.600 66.000 284.400 ;
        RECT 57.200 277.600 58.000 278.400 ;
        RECT 55.600 275.600 56.400 276.400 ;
        RECT 58.800 275.600 59.600 276.400 ;
        RECT 55.600 269.600 56.400 270.400 ;
        RECT 55.700 266.400 56.300 269.600 ;
        RECT 58.900 268.400 59.500 275.600 ;
        RECT 60.400 271.800 61.200 272.600 ;
        RECT 60.400 268.400 61.000 271.800 ;
        RECT 65.300 270.400 65.900 283.600 ;
        RECT 67.000 271.800 67.800 272.600 ;
        RECT 68.500 272.400 69.100 293.600 ;
        RECT 70.000 289.600 70.800 290.400 ;
        RECT 70.100 286.400 70.700 289.600 ;
        RECT 70.000 285.600 70.800 286.400 ;
        RECT 70.100 280.400 70.700 285.600 ;
        RECT 70.000 279.600 70.800 280.400 ;
        RECT 65.200 269.600 66.000 270.400 ;
        RECT 64.400 268.400 65.200 268.600 ;
        RECT 58.800 267.600 59.600 268.400 ;
        RECT 60.400 267.800 65.200 268.400 ;
        RECT 60.400 267.000 61.000 267.800 ;
        RECT 61.800 267.000 62.600 267.200 ;
        RECT 65.200 267.000 66.000 267.200 ;
        RECT 67.200 267.000 67.800 271.800 ;
        RECT 68.400 271.600 69.200 272.400 ;
        RECT 68.500 270.400 69.100 271.600 ;
        RECT 71.700 270.400 72.300 303.600 ;
        RECT 76.500 298.400 77.100 307.600 ;
        RECT 78.100 298.400 78.700 323.600 ;
        RECT 79.700 320.400 80.300 333.600 ;
        RECT 84.500 332.400 85.100 345.600 ;
        RECT 84.400 331.600 85.200 332.400 ;
        RECT 86.100 330.400 86.700 351.700 ;
        RECT 87.600 351.600 88.400 351.700 ;
        RECT 89.200 351.600 90.000 352.400 ;
        RECT 87.700 350.400 88.300 351.600 ;
        RECT 87.600 349.600 88.400 350.400 ;
        RECT 89.300 348.400 89.900 351.600 ;
        RECT 89.200 347.600 90.000 348.400 ;
        RECT 89.200 343.600 90.000 344.400 ;
        RECT 94.000 343.600 94.800 344.400 ;
        RECT 98.800 344.200 99.600 355.800 ;
        RECT 100.500 350.400 101.100 367.600 ;
        RECT 102.000 366.200 102.800 377.800 ;
        RECT 110.100 376.400 110.700 411.600 ;
        RECT 116.500 408.400 117.100 411.800 ;
        RECT 116.400 407.600 117.200 408.400 ;
        RECT 118.000 406.200 118.800 417.800 ;
        RECT 220.400 417.600 221.200 418.400 ;
        RECT 220.500 416.400 221.100 417.600 ;
        RECT 119.600 413.600 120.400 414.400 ;
        RECT 111.600 387.600 112.400 388.400 ;
        RECT 111.700 386.400 112.300 387.600 ;
        RECT 111.600 385.600 112.400 386.400 ;
        RECT 113.200 383.600 114.000 384.400 ;
        RECT 118.000 384.200 118.800 395.800 ;
        RECT 119.700 390.400 120.300 413.600 ;
        RECT 121.200 410.200 122.000 415.800 ;
        RECT 124.200 415.000 125.000 415.800 ;
        RECT 126.000 415.000 130.200 415.600 ;
        RECT 130.800 415.000 131.600 415.800 ;
        RECT 138.800 415.600 139.600 416.400 ;
        RECT 145.200 415.600 146.000 416.400 ;
        RECT 150.000 415.600 150.800 416.400 ;
        RECT 122.800 413.600 123.600 414.400 ;
        RECT 124.200 410.200 124.800 415.000 ;
        RECT 126.000 414.800 126.800 415.000 ;
        RECT 129.400 414.800 130.200 415.000 ;
        RECT 131.000 414.200 131.600 415.000 ;
        RECT 126.800 413.600 131.600 414.200 ;
        RECT 132.400 413.600 133.200 414.400 ;
        RECT 134.000 413.600 134.800 414.400 ;
        RECT 126.800 413.400 127.600 413.600 ;
        RECT 124.200 409.400 125.000 410.200 ;
        RECT 126.000 409.600 126.800 410.400 ;
        RECT 131.000 410.200 131.600 413.600 ;
        RECT 126.100 408.400 126.700 409.600 ;
        RECT 130.800 409.400 131.600 410.200 ;
        RECT 126.000 407.600 126.800 408.400 ;
        RECT 132.500 398.400 133.100 413.600 ;
        RECT 138.900 410.400 139.500 415.600 ;
        RECT 150.100 414.400 150.700 415.600 ;
        RECT 151.400 415.000 152.200 415.800 ;
        RECT 153.200 415.000 157.400 415.600 ;
        RECT 158.000 415.000 158.800 415.800 ;
        RECT 174.000 415.600 174.800 416.400 ;
        RECT 198.000 415.600 198.800 416.400 ;
        RECT 202.800 415.600 203.600 416.400 ;
        RECT 209.200 415.600 210.000 416.400 ;
        RECT 210.800 415.600 211.600 416.400 ;
        RECT 217.200 415.600 218.000 416.400 ;
        RECT 220.400 415.600 221.200 416.400 ;
        RECT 143.600 413.600 144.400 414.400 ;
        RECT 148.400 413.600 149.200 414.400 ;
        RECT 150.000 413.600 150.800 414.400 ;
        RECT 142.000 411.600 142.800 412.400 ;
        RECT 142.100 410.400 142.700 411.600 ;
        RECT 138.800 409.600 139.600 410.400 ;
        RECT 142.000 409.600 142.800 410.400 ;
        RECT 145.200 409.600 146.000 410.400 ;
        RECT 132.400 397.600 133.200 398.400 ;
        RECT 145.300 396.400 145.900 409.600 ;
        RECT 119.600 389.600 120.400 390.400 ;
        RECT 126.000 389.400 126.800 390.400 ;
        RECT 127.600 384.200 128.400 395.800 ;
        RECT 145.200 395.600 146.000 396.400 ;
        RECT 148.500 394.400 149.100 413.600 ;
        RECT 151.400 410.200 152.000 415.000 ;
        RECT 153.200 414.800 154.000 415.000 ;
        RECT 156.600 414.800 157.400 415.000 ;
        RECT 158.200 414.200 158.800 415.000 ;
        RECT 174.100 414.400 174.700 415.600 ;
        RECT 198.100 414.400 198.700 415.600 ;
        RECT 154.000 413.600 158.800 414.200 ;
        RECT 159.600 413.600 160.400 414.400 ;
        RECT 161.200 413.600 162.000 414.400 ;
        RECT 170.800 413.600 171.600 414.400 ;
        RECT 174.000 413.600 174.800 414.400 ;
        RECT 182.000 413.600 182.800 414.400 ;
        RECT 191.600 413.600 192.400 414.400 ;
        RECT 193.200 413.600 194.000 414.400 ;
        RECT 198.000 413.600 198.800 414.400 ;
        RECT 154.000 413.400 154.800 413.600 ;
        RECT 158.200 410.200 158.800 413.600 ;
        RECT 151.400 409.400 152.200 410.200 ;
        RECT 158.000 409.400 158.800 410.200 ;
        RECT 153.200 407.600 154.000 408.400 ;
        RECT 159.700 404.400 160.300 413.600 ;
        RECT 159.600 403.600 160.400 404.400 ;
        RECT 161.300 398.400 161.900 413.600 ;
        RECT 167.600 411.600 168.400 412.400 ;
        RECT 164.400 409.600 165.200 410.400 ;
        RECT 166.000 409.600 166.800 410.400 ;
        RECT 166.100 404.400 166.700 409.600 ;
        RECT 162.800 403.600 163.600 404.400 ;
        RECT 166.000 403.600 166.800 404.400 ;
        RECT 161.200 397.600 162.000 398.400 ;
        RECT 140.400 393.600 141.200 394.400 ;
        RECT 148.400 393.600 149.200 394.400 ;
        RECT 159.600 393.600 160.400 394.400 ;
        RECT 138.600 391.800 139.400 392.600 ;
        RECT 129.200 387.600 130.000 388.400 ;
        RECT 127.600 381.600 128.400 382.400 ;
        RECT 110.000 375.600 110.800 376.400 ;
        RECT 110.000 371.800 110.800 372.600 ;
        RECT 110.100 370.400 110.700 371.800 ;
        RECT 110.000 369.600 110.800 370.400 ;
        RECT 111.600 366.200 112.400 377.800 ;
        RECT 114.800 370.200 115.600 375.800 ;
        RECT 116.400 365.600 117.200 366.400 ;
        RECT 121.200 366.200 122.000 377.800 ;
        RECT 127.700 372.400 128.300 381.600 ;
        RECT 129.300 376.400 129.900 387.600 ;
        RECT 130.800 386.200 131.600 391.800 ;
        RECT 137.200 387.600 138.000 388.400 ;
        RECT 137.300 386.400 137.900 387.600 ;
        RECT 138.600 387.000 139.200 391.800 ;
        RECT 140.500 390.400 141.100 393.600 ;
        RECT 145.200 391.800 146.000 392.600 ;
        RECT 140.400 389.600 141.200 390.400 ;
        RECT 141.200 388.400 142.000 388.600 ;
        RECT 145.400 388.400 146.000 391.800 ;
        RECT 149.800 391.800 150.600 392.600 ;
        RECT 156.400 391.800 157.200 392.600 ;
        RECT 141.200 387.800 146.000 388.400 ;
        RECT 140.400 387.000 141.200 387.200 ;
        RECT 143.800 387.000 144.600 387.200 ;
        RECT 145.400 387.000 146.000 387.800 ;
        RECT 146.800 387.600 147.600 388.400 ;
        RECT 148.400 387.600 149.200 388.400 ;
        RECT 137.200 385.600 138.000 386.400 ;
        RECT 138.600 386.200 139.400 387.000 ;
        RECT 140.400 386.400 144.600 387.000 ;
        RECT 145.200 386.200 146.000 387.000 ;
        RECT 129.200 375.600 130.000 376.400 ;
        RECT 129.300 374.400 129.900 375.600 ;
        RECT 129.200 373.600 130.000 374.400 ;
        RECT 127.600 371.600 128.400 372.400 ;
        RECT 130.800 366.200 131.600 377.800 ;
        RECT 134.000 370.200 134.800 375.800 ;
        RECT 145.200 366.200 146.000 377.800 ;
        RECT 146.900 372.400 147.500 387.600 ;
        RECT 148.500 384.400 149.100 387.600 ;
        RECT 149.800 387.000 150.400 391.800 ;
        RECT 152.400 388.400 153.200 388.600 ;
        RECT 156.600 388.400 157.200 391.800 ;
        RECT 158.000 391.600 158.800 392.400 ;
        RECT 158.100 388.400 158.700 391.600 ;
        RECT 159.700 388.400 160.300 393.600 ;
        RECT 162.900 390.400 163.500 403.600 ;
        RECT 170.900 394.400 171.500 413.600 ;
        RECT 172.400 411.600 173.200 412.400 ;
        RECT 177.200 411.600 178.000 412.400 ;
        RECT 178.800 411.600 179.600 412.400 ;
        RECT 180.400 411.600 181.200 412.400 ;
        RECT 172.500 408.400 173.100 411.600 ;
        RECT 177.300 410.400 177.900 411.600 ;
        RECT 178.900 410.400 179.500 411.600 ;
        RECT 182.100 410.400 182.700 413.600 ;
        RECT 186.800 411.600 187.600 412.400 ;
        RECT 175.600 409.600 176.400 410.400 ;
        RECT 177.200 409.600 178.000 410.400 ;
        RECT 178.800 409.600 179.600 410.400 ;
        RECT 182.000 409.600 182.800 410.400 ;
        RECT 172.400 407.600 173.200 408.400 ;
        RECT 175.700 400.400 176.300 409.600 ;
        RECT 186.900 402.400 187.500 411.600 ;
        RECT 191.700 408.400 192.300 413.600 ;
        RECT 210.900 412.400 211.500 415.600 ;
        RECT 217.300 414.400 217.900 415.600 ;
        RECT 212.400 413.600 213.200 414.400 ;
        RECT 217.200 413.600 218.000 414.400 ;
        RECT 193.200 411.600 194.000 412.400 ;
        RECT 194.800 411.600 195.600 412.400 ;
        RECT 199.600 411.600 200.400 412.400 ;
        RECT 201.200 411.600 202.000 412.400 ;
        RECT 207.600 411.600 208.400 412.400 ;
        RECT 210.800 411.600 211.600 412.400 ;
        RECT 191.600 407.600 192.400 408.400 ;
        RECT 193.300 404.400 193.900 411.600 ;
        RECT 199.700 410.400 200.300 411.600 ;
        RECT 199.600 409.600 200.400 410.400 ;
        RECT 188.400 403.600 189.200 404.400 ;
        RECT 193.200 403.600 194.000 404.400 ;
        RECT 209.200 403.600 210.000 404.400 ;
        RECT 186.800 401.600 187.600 402.400 ;
        RECT 175.600 399.600 176.400 400.400 ;
        RECT 188.500 398.400 189.100 403.600 ;
        RECT 209.300 402.400 209.900 403.600 ;
        RECT 209.200 401.600 210.000 402.400 ;
        RECT 180.400 397.600 181.200 398.400 ;
        RECT 188.400 397.600 189.200 398.400 ;
        RECT 199.600 397.600 200.400 398.400 ;
        RECT 178.800 396.300 179.600 396.400 ;
        RECT 174.100 395.700 179.600 396.300 ;
        RECT 164.500 393.700 168.300 394.300 ;
        RECT 164.500 392.400 165.100 393.700 ;
        RECT 164.400 391.600 165.200 392.400 ;
        RECT 166.000 391.600 166.800 392.400 ;
        RECT 166.100 390.400 166.700 391.600 ;
        RECT 167.700 390.400 168.300 393.700 ;
        RECT 170.800 393.600 171.600 394.400 ;
        RECT 170.800 391.600 171.600 392.400 ;
        RECT 172.400 392.300 173.200 392.400 ;
        RECT 174.100 392.300 174.700 395.700 ;
        RECT 178.800 395.600 179.600 395.700 ;
        RECT 175.600 393.600 176.400 394.400 ;
        RECT 172.400 391.700 174.700 392.300 ;
        RECT 172.400 391.600 173.200 391.700 ;
        RECT 161.200 389.600 162.000 390.400 ;
        RECT 162.800 389.600 163.600 390.400 ;
        RECT 166.000 389.600 166.800 390.400 ;
        RECT 167.600 389.600 168.400 390.400 ;
        RECT 169.200 389.600 170.000 390.400 ;
        RECT 161.300 388.400 161.900 389.600 ;
        RECT 152.400 387.800 157.200 388.400 ;
        RECT 151.600 387.000 152.400 387.200 ;
        RECT 155.000 387.000 155.800 387.200 ;
        RECT 156.600 387.000 157.200 387.800 ;
        RECT 158.000 387.600 158.800 388.400 ;
        RECT 159.600 387.600 160.400 388.400 ;
        RECT 161.200 387.600 162.000 388.400 ;
        RECT 162.800 387.600 163.600 388.400 ;
        RECT 166.000 387.600 166.800 388.400 ;
        RECT 149.800 386.200 150.600 387.000 ;
        RECT 151.600 386.400 155.800 387.000 ;
        RECT 156.400 386.200 157.200 387.000 ;
        RECT 162.900 386.400 163.500 387.600 ;
        RECT 169.300 386.400 169.900 389.600 ;
        RECT 170.900 388.400 171.500 391.600 ;
        RECT 172.400 389.600 173.200 390.400 ;
        RECT 175.700 388.400 176.300 393.600 ;
        RECT 177.200 391.600 178.000 392.400 ;
        RECT 177.300 388.400 177.900 391.600 ;
        RECT 178.800 389.600 179.600 390.400 ;
        RECT 178.900 388.400 179.500 389.600 ;
        RECT 170.800 387.600 171.600 388.400 ;
        RECT 175.600 387.600 176.400 388.400 ;
        RECT 177.200 387.600 178.000 388.400 ;
        RECT 178.800 387.600 179.600 388.400 ;
        RECT 162.800 385.600 163.600 386.400 ;
        RECT 169.200 385.600 170.000 386.400 ;
        RECT 148.400 383.600 149.200 384.400 ;
        RECT 151.600 383.600 152.400 384.400 ;
        RECT 151.700 380.400 152.300 383.600 ;
        RECT 151.600 379.600 152.400 380.400 ;
        RECT 153.200 377.600 154.000 378.400 ;
        RECT 150.000 373.600 150.800 374.400 ;
        RECT 146.800 371.600 147.600 372.400 ;
        RECT 100.400 349.600 101.200 350.400 ;
        RECT 106.800 349.400 107.600 350.200 ;
        RECT 102.000 347.600 102.800 348.400 ;
        RECT 89.300 336.400 89.900 343.600 ;
        RECT 89.200 335.600 90.000 336.400 ;
        RECT 89.200 333.600 90.000 334.400 ;
        RECT 94.100 332.400 94.700 343.600 ;
        RECT 102.100 338.400 102.700 347.600 ;
        RECT 106.900 346.400 107.500 349.400 ;
        RECT 106.800 345.600 107.600 346.400 ;
        RECT 108.400 344.200 109.200 355.800 ;
        RECT 111.600 346.200 112.400 351.800 ;
        RECT 113.200 351.600 114.000 352.400 ;
        RECT 116.500 350.400 117.100 365.600 ;
        RECT 130.800 363.600 131.600 364.400 ;
        RECT 140.400 363.600 141.200 364.400 ;
        RECT 118.000 351.600 118.800 352.400 ;
        RECT 123.000 351.800 123.800 352.600 ;
        RECT 129.200 351.800 130.000 352.600 ;
        RECT 130.900 352.400 131.500 363.600 ;
        RECT 150.100 354.400 150.700 373.600 ;
        RECT 153.300 372.600 153.900 377.600 ;
        RECT 153.200 371.800 154.000 372.600 ;
        RECT 154.800 366.200 155.600 377.800 ;
        RECT 175.700 376.400 176.300 387.600 ;
        RECT 180.500 376.400 181.100 397.600 ;
        RECT 183.600 395.600 184.400 396.400 ;
        RECT 185.200 395.600 186.000 396.400 ;
        RECT 183.700 392.400 184.300 395.600 ;
        RECT 183.600 391.600 184.400 392.400 ;
        RECT 158.000 370.200 158.800 375.800 ;
        RECT 161.200 375.000 162.000 375.800 ;
        RECT 162.600 375.000 166.800 375.600 ;
        RECT 167.800 375.000 168.600 375.800 ;
        RECT 175.600 375.600 176.400 376.400 ;
        RECT 178.800 375.600 179.600 376.400 ;
        RECT 180.400 375.600 181.200 376.400 ;
        RECT 159.600 373.600 160.400 374.400 ;
        RECT 161.200 374.200 161.800 375.000 ;
        RECT 162.600 374.800 163.400 375.000 ;
        RECT 166.000 374.800 166.800 375.000 ;
        RECT 161.200 373.600 166.000 374.200 ;
        RECT 159.700 360.400 160.300 373.600 ;
        RECT 161.200 370.200 161.800 373.600 ;
        RECT 165.200 373.400 166.000 373.600 ;
        RECT 161.200 369.400 162.000 370.200 ;
        RECT 162.800 369.600 163.600 370.400 ;
        RECT 168.000 370.200 168.600 375.000 ;
        RECT 178.900 372.400 179.500 375.600 ;
        RECT 185.300 372.400 185.900 395.600 ;
        RECT 194.800 391.600 195.600 392.400 ;
        RECT 199.700 390.400 200.300 397.600 ;
        RECT 202.800 391.600 203.600 392.400 ;
        RECT 204.400 391.600 205.200 392.400 ;
        RECT 186.800 389.600 187.600 390.400 ;
        RECT 188.400 389.600 189.200 390.400 ;
        RECT 196.400 389.600 197.200 390.400 ;
        RECT 199.600 389.600 200.400 390.400 ;
        RECT 186.900 386.400 187.500 389.600 ;
        RECT 188.500 388.400 189.100 389.600 ;
        RECT 196.500 388.400 197.100 389.600 ;
        RECT 202.900 388.400 203.500 391.600 ;
        RECT 188.400 387.600 189.200 388.400 ;
        RECT 190.000 387.600 190.800 388.400 ;
        RECT 196.400 387.600 197.200 388.400 ;
        RECT 198.000 387.600 198.800 388.400 ;
        RECT 201.200 387.600 202.000 388.400 ;
        RECT 202.800 387.600 203.600 388.400 ;
        RECT 190.100 386.400 190.700 387.600 ;
        RECT 196.500 386.400 197.100 387.600 ;
        RECT 186.800 385.600 187.600 386.400 ;
        RECT 190.000 385.600 190.800 386.400 ;
        RECT 196.400 385.600 197.200 386.400 ;
        RECT 172.400 371.600 173.200 372.400 ;
        RECT 177.200 371.600 178.000 372.400 ;
        RECT 178.800 371.600 179.600 372.400 ;
        RECT 183.600 371.600 184.400 372.400 ;
        RECT 185.200 371.600 186.000 372.400 ;
        RECT 167.800 369.400 168.600 370.200 ;
        RECT 172.500 368.400 173.100 371.600 ;
        RECT 172.400 367.600 173.200 368.400 ;
        RECT 177.300 364.400 177.900 371.600 ;
        RECT 186.900 370.400 187.500 385.600 ;
        RECT 191.600 383.600 192.400 384.400 ;
        RECT 191.700 378.300 192.300 383.600 ;
        RECT 190.100 377.700 192.300 378.300 ;
        RECT 186.800 369.600 187.600 370.400 ;
        RECT 190.100 370.300 190.700 377.700 ;
        RECT 191.600 375.600 192.400 376.400 ;
        RECT 194.800 375.600 195.600 376.400 ;
        RECT 194.900 374.400 195.500 375.600 ;
        RECT 196.500 374.400 197.100 385.600 ;
        RECT 198.100 378.400 198.700 387.600 ;
        RECT 198.000 377.600 198.800 378.400 ;
        RECT 191.600 374.300 192.400 374.400 ;
        RECT 191.600 373.700 193.900 374.300 ;
        RECT 191.600 373.600 192.400 373.700 ;
        RECT 191.600 370.300 192.400 370.400 ;
        RECT 190.100 369.700 192.400 370.300 ;
        RECT 191.600 369.600 192.400 369.700 ;
        RECT 193.300 368.400 193.900 373.700 ;
        RECT 194.800 373.600 195.600 374.400 ;
        RECT 196.400 373.600 197.200 374.400 ;
        RECT 199.600 373.600 200.400 374.400 ;
        RECT 199.600 371.600 200.400 372.400 ;
        RECT 199.700 370.400 200.300 371.600 ;
        RECT 199.600 369.600 200.400 370.400 ;
        RECT 190.000 367.600 190.800 368.400 ;
        RECT 193.200 367.600 194.000 368.400 ;
        RECT 190.100 364.400 190.700 367.600 ;
        RECT 201.300 364.400 201.900 387.600 ;
        RECT 204.500 386.400 205.100 391.600 ;
        RECT 207.600 389.600 208.400 390.400 ;
        RECT 209.200 389.600 210.000 390.400 ;
        RECT 204.400 385.600 205.200 386.400 ;
        RECT 207.700 376.400 208.300 389.600 ;
        RECT 202.800 375.600 203.600 376.400 ;
        RECT 204.400 375.600 205.200 376.400 ;
        RECT 207.600 375.600 208.400 376.400 ;
        RECT 204.500 370.400 205.100 375.600 ;
        RECT 209.300 372.400 209.900 389.600 ;
        RECT 210.900 376.400 211.500 411.600 ;
        RECT 218.800 409.600 219.600 410.400 ;
        RECT 218.900 404.400 219.500 409.600 ;
        RECT 225.200 406.200 226.000 417.800 ;
        RECT 228.400 411.600 229.200 412.400 ;
        RECT 233.200 411.600 234.000 412.600 ;
        RECT 228.500 410.400 229.100 411.600 ;
        RECT 228.400 409.600 229.200 410.400 ;
        RECT 218.800 403.600 219.600 404.400 ;
        RECT 220.400 403.600 221.200 404.400 ;
        RECT 226.800 403.600 227.600 404.400 ;
        RECT 215.600 397.600 216.400 398.400 ;
        RECT 214.000 393.600 214.800 394.400 ;
        RECT 212.400 387.600 213.200 388.400 ;
        RECT 214.100 382.400 214.700 393.600 ;
        RECT 215.700 390.400 216.300 397.600 ;
        RECT 218.900 392.300 219.500 403.600 ;
        RECT 220.500 394.400 221.100 403.600 ;
        RECT 226.900 398.400 227.500 403.600 ;
        RECT 226.800 397.600 227.600 398.400 ;
        RECT 220.400 393.600 221.200 394.400 ;
        RECT 220.400 392.300 221.200 392.400 ;
        RECT 218.900 391.700 221.200 392.300 ;
        RECT 220.400 391.600 221.200 391.700 ;
        RECT 225.200 391.600 226.000 392.400 ;
        RECT 215.600 389.600 216.400 390.400 ;
        RECT 214.000 381.600 214.800 382.400 ;
        RECT 210.800 375.600 211.600 376.400 ;
        RECT 212.400 373.600 213.200 374.400 ;
        RECT 207.600 371.600 208.400 372.400 ;
        RECT 209.200 371.600 210.000 372.400 ;
        RECT 210.800 371.600 211.600 372.400 ;
        RECT 212.500 370.400 213.100 373.600 ;
        RECT 204.400 369.600 205.200 370.400 ;
        RECT 212.400 369.600 213.200 370.400 ;
        RECT 215.700 368.400 216.300 389.600 ;
        RECT 220.400 387.600 221.200 388.400 ;
        RECT 223.600 387.600 224.400 388.400 ;
        RECT 218.800 385.600 219.600 386.400 ;
        RECT 218.900 372.400 219.500 385.600 ;
        RECT 220.500 374.400 221.100 387.600 ;
        RECT 225.300 386.300 225.900 391.600 ;
        RECT 228.500 390.400 229.100 409.600 ;
        RECT 234.800 406.200 235.600 417.800 ;
        RECT 238.000 410.200 238.800 415.800 ;
        RECT 241.200 415.600 242.000 416.400 ;
        RECT 244.400 413.600 245.200 414.400 ;
        RECT 239.600 411.600 240.400 412.400 ;
        RECT 242.800 403.600 243.600 404.400 ;
        RECT 233.200 399.600 234.000 400.400 ;
        RECT 233.300 390.400 233.900 399.600 ;
        RECT 234.800 395.600 235.600 396.400 ;
        RECT 242.800 393.600 243.600 394.400 ;
        RECT 239.600 392.300 240.400 392.400 ;
        RECT 239.600 391.700 241.900 392.300 ;
        RECT 239.600 391.600 240.400 391.700 ;
        RECT 228.400 389.600 229.200 390.400 ;
        RECT 233.200 389.600 234.000 390.400 ;
        RECT 238.000 389.600 238.800 390.400 ;
        RECT 238.100 388.400 238.700 389.600 ;
        RECT 228.400 387.600 229.200 388.400 ;
        RECT 238.000 387.600 238.800 388.400 ;
        RECT 230.000 386.300 230.800 386.400 ;
        RECT 225.300 385.700 230.800 386.300 ;
        RECT 230.000 385.600 230.800 385.700 ;
        RECT 233.200 377.600 234.000 378.400 ;
        RECT 230.000 375.600 230.800 376.400 ;
        RECT 231.800 375.600 232.600 375.800 ;
        RECT 230.100 374.400 230.700 375.600 ;
        RECT 231.800 375.000 237.400 375.600 ;
        RECT 238.000 375.000 238.800 375.800 ;
        RECT 239.600 375.600 240.400 376.400 ;
        RECT 220.400 373.600 221.200 374.400 ;
        RECT 223.600 373.600 224.400 374.400 ;
        RECT 225.200 373.600 226.000 374.400 ;
        RECT 228.400 373.600 229.200 374.400 ;
        RECT 230.000 373.600 230.800 374.400 ;
        RECT 217.200 371.600 218.000 372.400 ;
        RECT 218.800 371.600 219.600 372.400 ;
        RECT 217.300 370.400 217.900 371.600 ;
        RECT 217.200 369.600 218.000 370.400 ;
        RECT 207.600 367.600 208.400 368.400 ;
        RECT 215.600 367.600 216.400 368.400 ;
        RECT 177.200 363.600 178.000 364.400 ;
        RECT 190.000 363.600 190.800 364.400 ;
        RECT 201.200 363.600 202.000 364.400 ;
        RECT 159.600 359.600 160.400 360.400 ;
        RECT 166.000 357.600 166.800 358.400 ;
        RECT 150.000 353.600 150.800 354.400 ;
        RECT 116.400 349.600 117.200 350.400 ;
        RECT 116.400 347.600 117.200 348.400 ;
        RECT 113.200 343.600 114.000 344.400 ;
        RECT 113.300 340.300 113.900 343.600 ;
        RECT 116.500 342.400 117.100 347.600 ;
        RECT 118.100 344.400 118.700 351.600 ;
        RECT 121.200 349.600 122.000 350.400 ;
        RECT 121.300 348.400 121.900 349.600 ;
        RECT 119.600 347.600 120.400 348.400 ;
        RECT 121.200 347.600 122.000 348.400 ;
        RECT 123.000 347.000 123.600 351.800 ;
        RECT 124.200 349.800 125.000 350.600 ;
        RECT 124.400 348.400 125.000 349.800 ;
        RECT 129.400 348.400 130.000 351.800 ;
        RECT 130.800 351.600 131.600 352.400 ;
        RECT 135.600 351.600 136.400 352.400 ;
        RECT 137.200 351.600 138.000 352.400 ;
        RECT 143.800 351.800 144.600 352.600 ;
        RECT 150.000 351.800 150.800 352.600 ;
        RECT 130.900 348.400 131.500 351.600 ;
        RECT 132.400 349.600 133.200 350.400 ;
        RECT 132.500 348.400 133.100 349.600 ;
        RECT 124.400 347.800 130.000 348.400 ;
        RECT 124.400 347.000 125.200 347.200 ;
        RECT 127.800 347.000 128.600 347.200 ;
        RECT 129.400 347.000 130.000 347.800 ;
        RECT 130.800 347.600 131.600 348.400 ;
        RECT 132.400 347.600 133.200 348.400 ;
        RECT 123.000 346.400 128.600 347.000 ;
        RECT 123.000 346.200 123.800 346.400 ;
        RECT 129.200 346.200 130.000 347.000 ;
        RECT 118.000 343.600 118.800 344.400 ;
        RECT 122.800 343.600 123.600 344.400 ;
        RECT 127.600 343.600 128.400 344.400 ;
        RECT 116.400 341.600 117.200 342.400 ;
        RECT 111.700 339.700 113.900 340.300 ;
        RECT 102.000 337.600 102.800 338.400 ;
        RECT 108.400 337.600 109.200 338.400 ;
        RECT 102.100 336.400 102.700 337.600 ;
        RECT 95.600 335.600 96.400 336.400 ;
        RECT 102.000 335.600 102.800 336.400 ;
        RECT 103.600 335.600 104.400 336.400 ;
        RECT 95.700 334.400 96.300 335.600 ;
        RECT 102.100 334.400 102.700 335.600 ;
        RECT 108.500 334.400 109.100 337.600 ;
        RECT 95.600 333.600 96.400 334.400 ;
        RECT 97.200 333.600 98.000 334.400 ;
        RECT 102.000 333.600 102.800 334.400 ;
        RECT 106.800 333.600 107.600 334.400 ;
        RECT 108.400 333.600 109.200 334.400 ;
        RECT 89.200 331.600 90.000 332.400 ;
        RECT 90.800 331.600 91.600 332.400 ;
        RECT 94.000 331.600 94.800 332.400 ;
        RECT 95.600 331.600 96.400 332.400 ;
        RECT 89.300 330.400 89.900 331.600 ;
        RECT 86.000 329.600 86.800 330.400 ;
        RECT 89.200 329.600 90.000 330.400 ;
        RECT 81.200 325.600 82.000 326.400 ;
        RECT 79.600 319.600 80.400 320.400 ;
        RECT 79.600 307.600 80.400 308.400 ;
        RECT 81.300 306.300 81.900 325.600 ;
        RECT 84.400 309.600 85.200 310.400 ;
        RECT 84.500 308.400 85.100 309.600 ;
        RECT 86.100 308.400 86.700 329.600 ;
        RECT 82.800 307.600 83.600 308.400 ;
        RECT 84.400 307.600 85.200 308.400 ;
        RECT 86.000 307.600 86.800 308.400 ;
        RECT 82.900 306.400 83.500 307.600 ;
        RECT 79.700 305.700 81.900 306.300 ;
        RECT 73.200 297.600 74.000 298.400 ;
        RECT 76.400 297.600 77.200 298.400 ;
        RECT 78.000 297.600 78.800 298.400 ;
        RECT 73.300 294.400 73.900 297.600 ;
        RECT 74.800 295.600 75.600 296.400 ;
        RECT 76.400 295.600 77.200 296.400 ;
        RECT 78.000 295.600 78.800 296.400 ;
        RECT 73.200 293.600 74.000 294.400 ;
        RECT 74.900 292.400 75.500 295.600 ;
        RECT 76.500 292.400 77.100 295.600 ;
        RECT 78.100 292.400 78.700 295.600 ;
        RECT 79.700 294.400 80.300 305.700 ;
        RECT 82.800 305.600 83.600 306.400 ;
        RECT 84.400 305.600 85.200 306.400 ;
        RECT 87.600 305.600 88.400 306.400 ;
        RECT 81.200 303.600 82.000 304.400 ;
        RECT 79.600 293.600 80.400 294.400 ;
        RECT 74.800 291.600 75.600 292.400 ;
        RECT 76.400 291.600 77.200 292.400 ;
        RECT 78.000 291.600 78.800 292.400 ;
        RECT 74.900 290.400 75.500 291.600 ;
        RECT 74.800 289.600 75.600 290.400 ;
        RECT 81.300 288.400 81.900 303.600 ;
        RECT 82.800 299.600 83.600 300.400 ;
        RECT 82.900 288.400 83.500 299.600 ;
        RECT 84.500 294.400 85.100 305.600 ;
        RECT 89.300 294.400 89.900 329.600 ;
        RECT 90.900 316.400 91.500 331.600 ;
        RECT 97.300 330.400 97.900 333.600 ;
        RECT 102.000 331.600 102.800 332.400 ;
        RECT 110.000 331.600 110.800 332.400 ;
        RECT 97.200 329.600 98.000 330.400 ;
        RECT 90.800 315.600 91.600 316.400 ;
        RECT 95.600 309.600 96.400 310.400 ;
        RECT 97.300 308.400 97.900 329.600 ;
        RECT 100.400 323.600 101.200 324.400 ;
        RECT 98.800 312.300 99.600 312.400 ;
        RECT 100.500 312.300 101.100 323.600 ;
        RECT 98.800 311.700 101.100 312.300 ;
        RECT 98.800 311.600 99.600 311.700 ;
        RECT 92.400 308.300 93.200 308.400 ;
        RECT 90.900 307.700 93.200 308.300 ;
        RECT 90.900 302.400 91.500 307.700 ;
        RECT 92.400 307.600 93.200 307.700 ;
        RECT 97.200 307.600 98.000 308.400 ;
        RECT 102.100 306.400 102.700 331.600 ;
        RECT 110.000 311.600 110.800 312.400 ;
        RECT 106.800 309.600 107.600 310.400 ;
        RECT 103.600 307.600 104.400 308.400 ;
        RECT 105.200 307.600 106.000 308.400 ;
        RECT 108.400 307.600 109.200 308.400 ;
        RECT 92.400 305.600 93.200 306.400 ;
        RECT 100.400 305.600 101.200 306.400 ;
        RECT 102.000 305.600 102.800 306.400 ;
        RECT 90.800 301.600 91.600 302.400 ;
        RECT 90.900 298.400 91.500 301.600 ;
        RECT 90.800 297.600 91.600 298.400 ;
        RECT 92.500 294.400 93.100 305.600 ;
        RECT 98.800 303.600 99.600 304.400 ;
        RECT 102.000 303.600 102.800 304.400 ;
        RECT 98.900 298.400 99.500 303.600 ;
        RECT 103.700 298.400 104.300 307.600 ;
        RECT 105.300 306.400 105.900 307.600 ;
        RECT 105.200 305.600 106.000 306.400 ;
        RECT 98.800 297.600 99.600 298.400 ;
        RECT 102.000 297.600 102.800 298.400 ;
        RECT 103.600 297.600 104.400 298.400 ;
        RECT 102.100 296.300 102.700 297.600 ;
        RECT 108.500 296.300 109.100 307.600 ;
        RECT 110.100 298.400 110.700 311.600 ;
        RECT 111.700 310.400 112.300 339.700 ;
        RECT 113.200 337.600 114.000 338.400 ;
        RECT 116.500 336.400 117.100 341.600 ;
        RECT 118.100 336.400 118.700 343.600 ;
        RECT 119.600 341.600 120.400 342.400 ;
        RECT 116.400 335.600 117.200 336.400 ;
        RECT 118.000 335.600 118.800 336.400 ;
        RECT 118.100 334.400 118.700 335.600 ;
        RECT 118.000 333.600 118.800 334.400 ;
        RECT 119.700 332.400 120.300 341.600 ;
        RECT 122.900 332.400 123.500 343.600 ;
        RECT 124.400 337.600 125.200 338.400 ;
        RECT 113.200 331.600 114.000 332.400 ;
        RECT 119.600 331.600 120.400 332.400 ;
        RECT 122.800 331.600 123.600 332.400 ;
        RECT 113.200 329.600 114.000 330.400 ;
        RECT 119.600 329.600 120.400 330.400 ;
        RECT 111.600 309.600 112.400 310.400 ;
        RECT 113.300 308.400 113.900 329.600 ;
        RECT 122.800 319.600 123.600 320.400 ;
        RECT 119.600 313.600 120.400 314.400 ;
        RECT 122.900 312.400 123.500 319.600 ;
        RECT 124.500 312.400 125.100 337.600 ;
        RECT 126.000 333.600 126.800 334.400 ;
        RECT 127.700 316.400 128.300 343.600 ;
        RECT 130.900 334.400 131.500 347.600 ;
        RECT 137.300 346.400 137.900 351.600 ;
        RECT 142.000 347.600 142.800 348.400 ;
        RECT 143.800 347.000 144.400 351.800 ;
        RECT 145.000 349.800 145.800 350.600 ;
        RECT 145.200 348.400 145.800 349.800 ;
        RECT 150.200 348.400 150.800 351.800 ;
        RECT 145.200 347.800 150.800 348.400 ;
        RECT 145.200 347.000 146.000 347.200 ;
        RECT 148.600 347.000 149.400 347.200 ;
        RECT 150.200 347.000 150.800 347.800 ;
        RECT 151.600 347.600 152.400 348.400 ;
        RECT 143.800 346.400 149.400 347.000 ;
        RECT 137.200 345.600 138.000 346.400 ;
        RECT 143.800 346.200 144.600 346.400 ;
        RECT 150.000 346.200 150.800 347.000 ;
        RECT 140.400 343.600 141.200 344.400 ;
        RECT 148.400 343.600 149.200 344.400 ;
        RECT 151.700 344.300 152.300 347.600 ;
        RECT 153.200 344.300 154.000 344.400 ;
        RECT 151.700 343.700 154.000 344.300 ;
        RECT 140.500 338.400 141.100 343.600 ;
        RECT 151.700 342.400 152.300 343.700 ;
        RECT 153.200 343.600 154.000 343.700 ;
        RECT 154.800 343.600 155.600 344.400 ;
        RECT 158.000 344.200 158.800 355.800 ;
        RECT 159.600 353.600 160.400 354.400 ;
        RECT 159.700 350.400 160.300 353.600 ;
        RECT 159.600 349.600 160.400 350.400 ;
        RECT 166.100 350.200 166.700 357.600 ;
        RECT 166.000 349.400 166.800 350.200 ;
        RECT 167.600 344.200 168.400 355.800 ;
        RECT 170.800 346.200 171.600 351.800 ;
        RECT 172.400 347.600 173.200 348.400 ;
        RECT 172.500 344.400 173.100 347.600 ;
        RECT 172.400 343.600 173.200 344.400 ;
        RECT 177.200 344.200 178.000 355.800 ;
        RECT 185.200 355.600 186.000 356.400 ;
        RECT 178.800 353.600 179.600 354.400 ;
        RECT 178.900 350.400 179.500 353.600 ;
        RECT 178.800 349.600 179.600 350.400 ;
        RECT 185.300 350.200 185.900 355.600 ;
        RECT 185.200 349.400 186.000 350.200 ;
        RECT 183.600 347.600 184.400 348.400 ;
        RECT 151.600 341.600 152.400 342.400 ;
        RECT 153.300 340.400 153.900 343.600 ;
        RECT 153.200 339.600 154.000 340.400 ;
        RECT 140.400 337.600 141.200 338.400 ;
        RECT 145.000 335.000 145.800 335.800 ;
        RECT 146.800 335.000 151.000 335.600 ;
        RECT 151.600 335.000 152.400 335.800 ;
        RECT 130.800 333.600 131.600 334.400 ;
        RECT 134.000 333.600 134.800 334.400 ;
        RECT 137.200 333.600 138.000 334.400 ;
        RECT 143.600 333.600 144.400 334.400 ;
        RECT 137.300 332.400 137.900 333.600 ;
        RECT 130.800 331.600 131.600 332.400 ;
        RECT 137.200 331.600 138.000 332.400 ;
        RECT 138.800 331.600 139.600 332.400 ;
        RECT 130.900 330.400 131.500 331.600 ;
        RECT 130.800 329.600 131.600 330.400 ;
        RECT 145.000 330.200 145.600 335.000 ;
        RECT 146.800 334.800 147.600 335.000 ;
        RECT 150.200 334.800 151.000 335.000 ;
        RECT 151.800 334.200 152.400 335.000 ;
        RECT 154.900 334.400 155.500 343.600 ;
        RECT 174.000 339.600 174.800 340.400 ;
        RECT 162.800 337.600 163.600 338.400 ;
        RECT 172.400 337.600 173.200 338.400 ;
        RECT 162.900 336.400 163.500 337.600 ;
        RECT 159.600 335.600 160.400 336.400 ;
        RECT 162.800 335.600 163.600 336.400 ;
        RECT 164.400 335.600 165.200 336.400 ;
        RECT 172.500 334.400 173.100 337.600 ;
        RECT 174.100 334.400 174.700 339.600 ;
        RECT 175.600 335.000 176.400 335.800 ;
        RECT 177.000 335.000 181.200 335.600 ;
        RECT 182.200 335.000 183.000 335.800 ;
        RECT 147.600 333.600 152.400 334.200 ;
        RECT 154.800 333.600 155.600 334.400 ;
        RECT 156.400 333.600 157.200 334.400 ;
        RECT 159.600 333.600 160.400 334.400 ;
        RECT 172.400 333.600 173.200 334.400 ;
        RECT 174.000 333.600 174.800 334.400 ;
        RECT 175.600 334.200 176.200 335.000 ;
        RECT 177.000 334.800 177.800 335.000 ;
        RECT 180.400 334.800 181.200 335.000 ;
        RECT 175.600 333.600 180.400 334.200 ;
        RECT 147.600 333.400 148.400 333.600 ;
        RECT 151.800 330.200 152.400 333.600 ;
        RECT 154.900 332.400 155.500 333.600 ;
        RECT 154.800 331.600 155.600 332.400 ;
        RECT 158.000 331.600 158.800 332.400 ;
        RECT 167.600 331.600 168.400 332.400 ;
        RECT 130.900 320.400 131.500 329.600 ;
        RECT 145.000 329.400 145.800 330.200 ;
        RECT 151.600 329.400 152.400 330.200 ;
        RECT 146.800 323.600 147.600 324.400 ;
        RECT 130.800 319.600 131.600 320.400 ;
        RECT 127.600 315.600 128.400 316.400 ;
        RECT 122.800 311.600 123.600 312.400 ;
        RECT 124.400 311.600 125.200 312.400 ;
        RECT 127.600 311.600 128.400 312.400 ;
        RECT 113.200 307.600 114.000 308.400 ;
        RECT 118.000 307.600 118.800 308.400 ;
        RECT 116.400 305.600 117.200 306.400 ;
        RECT 114.800 303.600 115.600 304.400 ;
        RECT 114.900 300.400 115.500 303.600 ;
        RECT 114.800 299.600 115.600 300.400 ;
        RECT 110.000 297.600 110.800 298.400 ;
        RECT 113.200 297.600 114.000 298.400 ;
        RECT 113.300 296.400 113.900 297.600 ;
        RECT 94.000 295.000 94.800 295.800 ;
        RECT 95.400 295.000 99.600 295.600 ;
        RECT 100.600 295.000 101.400 295.800 ;
        RECT 102.100 295.700 104.300 296.300 ;
        RECT 84.400 293.600 85.200 294.400 ;
        RECT 86.000 293.600 86.800 294.400 ;
        RECT 87.600 293.600 88.400 294.400 ;
        RECT 89.200 293.600 90.000 294.400 ;
        RECT 92.400 293.600 93.200 294.400 ;
        RECT 94.000 294.200 94.600 295.000 ;
        RECT 95.400 294.800 96.200 295.000 ;
        RECT 98.800 294.800 99.600 295.000 ;
        RECT 94.000 293.600 98.800 294.200 ;
        RECT 86.100 292.400 86.700 293.600 ;
        RECT 87.700 292.400 88.300 293.600 ;
        RECT 86.000 291.600 86.800 292.400 ;
        RECT 87.600 291.600 88.400 292.400 ;
        RECT 90.800 291.600 91.600 292.400 ;
        RECT 76.400 287.600 77.200 288.400 ;
        RECT 81.200 287.600 82.000 288.400 ;
        RECT 82.800 287.600 83.600 288.400 ;
        RECT 76.500 270.400 77.100 287.600 ;
        RECT 81.200 283.600 82.000 284.400 ;
        RECT 79.600 277.600 80.400 278.400 ;
        RECT 79.700 272.400 80.300 277.600 ;
        RECT 79.600 271.600 80.400 272.400 ;
        RECT 68.400 269.600 69.200 270.400 ;
        RECT 71.600 269.600 72.400 270.400 ;
        RECT 76.400 269.600 77.200 270.400 ;
        RECT 68.400 267.600 69.200 268.400 ;
        RECT 55.600 265.600 56.400 266.400 ;
        RECT 60.400 266.200 61.200 267.000 ;
        RECT 61.800 266.400 66.000 267.000 ;
        RECT 67.000 266.200 67.800 267.000 ;
        RECT 62.000 263.600 62.800 264.400 ;
        RECT 54.000 259.600 54.800 260.400 ;
        RECT 49.200 255.600 50.000 256.400 ;
        RECT 50.800 255.600 51.600 256.400 ;
        RECT 52.400 255.000 53.200 255.800 ;
        RECT 53.800 255.000 58.000 255.600 ;
        RECT 59.000 255.000 59.800 255.800 ;
        RECT 39.600 253.600 40.400 254.400 ;
        RECT 46.000 253.600 46.800 254.400 ;
        RECT 52.400 254.200 53.000 255.000 ;
        RECT 53.800 254.800 54.600 255.000 ;
        RECT 57.200 254.800 58.000 255.000 ;
        RECT 52.400 253.600 57.200 254.200 ;
        RECT 25.200 251.600 26.000 252.400 ;
        RECT 26.800 251.600 27.600 252.400 ;
        RECT 31.600 251.600 32.400 252.400 ;
        RECT 33.200 251.600 34.000 252.400 ;
        RECT 34.800 251.600 35.600 252.400 ;
        RECT 38.000 251.600 38.800 252.400 ;
        RECT 46.000 251.600 46.800 252.400 ;
        RECT 34.900 250.400 35.500 251.600 ;
        RECT 46.100 250.400 46.700 251.600 ;
        RECT 31.600 249.600 32.400 250.400 ;
        RECT 34.800 249.600 35.600 250.400 ;
        RECT 41.200 249.600 42.000 250.400 ;
        RECT 46.000 249.600 46.800 250.400 ;
        RECT 52.400 250.200 53.000 253.600 ;
        RECT 56.400 253.400 57.200 253.600 ;
        RECT 59.200 250.200 59.800 255.000 ;
        RECT 63.400 255.000 64.200 255.800 ;
        RECT 65.200 255.000 69.400 255.600 ;
        RECT 70.000 255.000 70.800 255.800 ;
        RECT 60.400 253.600 61.200 254.400 ;
        RECT 62.000 253.600 62.800 254.400 ;
        RECT 30.000 243.600 30.800 244.400 ;
        RECT 22.000 231.800 22.800 232.600 ;
        RECT 28.600 231.800 29.400 232.600 ;
        RECT 22.000 228.400 22.600 231.800 ;
        RECT 26.000 228.400 26.800 228.600 ;
        RECT 20.400 227.600 21.200 228.400 ;
        RECT 22.000 227.800 26.800 228.400 ;
        RECT 22.000 227.000 22.600 227.800 ;
        RECT 23.400 227.000 24.200 227.200 ;
        RECT 26.800 227.000 27.600 227.200 ;
        RECT 28.800 227.000 29.400 231.800 ;
        RECT 30.100 228.400 30.700 243.600 ;
        RECT 31.700 228.400 32.300 249.600 ;
        RECT 52.400 249.400 53.200 250.200 ;
        RECT 59.000 249.400 59.800 250.200 ;
        RECT 63.400 250.200 64.000 255.000 ;
        RECT 65.200 254.800 66.000 255.000 ;
        RECT 68.600 254.800 69.400 255.000 ;
        RECT 70.200 254.200 70.800 255.000 ;
        RECT 66.000 253.600 70.800 254.200 ;
        RECT 66.000 253.400 66.800 253.600 ;
        RECT 70.200 250.200 70.800 253.600 ;
        RECT 71.700 252.400 72.300 269.600 ;
        RECT 76.400 267.600 77.200 268.400 ;
        RECT 73.200 263.600 74.000 264.400 ;
        RECT 73.300 254.400 73.900 263.600 ;
        RECT 76.500 258.400 77.100 267.600 ;
        RECT 79.600 263.600 80.400 264.400 ;
        RECT 76.400 257.600 77.200 258.400 ;
        RECT 78.000 257.600 78.800 258.400 ;
        RECT 78.100 256.400 78.700 257.600 ;
        RECT 78.000 255.600 78.800 256.400 ;
        RECT 73.200 253.600 74.000 254.400 ;
        RECT 74.800 253.600 75.600 254.400 ;
        RECT 78.000 253.600 78.800 254.400 ;
        RECT 71.600 251.600 72.400 252.400 ;
        RECT 63.400 249.400 64.200 250.200 ;
        RECT 70.000 249.400 70.800 250.200 ;
        RECT 38.000 243.600 38.800 244.400 ;
        RECT 54.000 243.600 54.800 244.400 ;
        RECT 66.800 243.600 67.600 244.400 ;
        RECT 33.200 231.800 34.000 232.600 ;
        RECT 33.200 228.400 33.800 231.800 ;
        RECT 38.100 230.400 38.700 243.600 ;
        RECT 39.800 231.800 40.600 232.600 ;
        RECT 38.000 229.600 38.800 230.400 ;
        RECT 37.200 228.400 38.000 228.600 ;
        RECT 30.000 227.600 30.800 228.400 ;
        RECT 31.600 227.600 32.400 228.400 ;
        RECT 33.200 227.800 38.000 228.400 ;
        RECT 22.000 226.200 22.800 227.000 ;
        RECT 23.400 226.400 27.600 227.000 ;
        RECT 28.600 226.200 29.400 227.000 ;
        RECT 33.200 227.000 33.800 227.800 ;
        RECT 34.600 227.000 35.400 227.200 ;
        RECT 38.000 227.000 38.800 227.200 ;
        RECT 40.000 227.000 40.600 231.800 ;
        RECT 41.200 229.600 42.000 230.400 ;
        RECT 41.300 228.400 41.900 229.600 ;
        RECT 41.200 227.600 42.000 228.400 ;
        RECT 33.200 226.200 34.000 227.000 ;
        RECT 34.600 226.400 38.800 227.000 ;
        RECT 39.800 226.200 40.600 227.000 ;
        RECT 25.200 223.600 26.000 224.400 ;
        RECT 34.800 223.600 35.600 224.400 ;
        RECT 42.800 223.600 43.600 224.400 ;
        RECT 47.600 224.200 48.400 235.800 ;
        RECT 12.400 213.600 13.200 214.400 ;
        RECT 12.500 212.400 13.100 213.600 ;
        RECT 12.400 211.600 13.200 212.400 ;
        RECT 12.500 190.400 13.100 211.600 ;
        RECT 14.000 206.200 14.800 217.800 ;
        RECT 20.400 210.200 21.200 215.800 ;
        RECT 23.600 206.200 24.400 217.800 ;
        RECT 18.800 203.600 19.600 204.400 ;
        RECT 9.200 189.600 10.000 190.400 ;
        RECT 12.400 189.600 13.200 190.400 ;
        RECT 1.200 163.600 2.000 164.400 ;
        RECT 1.300 148.400 1.900 163.600 ;
        RECT 2.900 150.400 3.500 183.600 ;
        RECT 6.000 166.200 6.800 177.800 ;
        RECT 12.500 174.400 13.100 189.600 ;
        RECT 14.000 184.200 14.800 195.800 ;
        RECT 18.900 186.400 19.500 203.600 ;
        RECT 18.800 185.600 19.600 186.400 ;
        RECT 20.400 186.200 21.200 191.800 ;
        RECT 18.800 183.600 19.600 184.400 ;
        RECT 23.600 184.200 24.400 195.800 ;
        RECT 25.300 190.200 25.900 223.600 ;
        RECT 26.800 215.600 27.600 216.400 ;
        RECT 26.900 212.400 27.500 215.600 ;
        RECT 31.600 213.600 32.400 214.400 ;
        RECT 31.700 212.400 32.300 213.600 ;
        RECT 26.800 211.600 27.600 212.400 ;
        RECT 31.600 211.600 32.400 212.400 ;
        RECT 31.700 190.400 32.300 211.600 ;
        RECT 33.200 206.200 34.000 217.800 ;
        RECT 34.900 216.400 35.500 223.600 ;
        RECT 34.800 215.600 35.600 216.400 ;
        RECT 38.000 203.600 38.800 204.400 ;
        RECT 39.600 203.600 40.400 204.400 ;
        RECT 25.200 189.400 26.000 190.200 ;
        RECT 31.600 189.600 32.400 190.400 ;
        RECT 25.200 185.600 26.000 186.400 ;
        RECT 14.000 175.600 14.800 176.400 ;
        RECT 12.400 173.600 13.200 174.400 ;
        RECT 14.100 172.600 14.700 175.600 ;
        RECT 14.000 171.800 14.800 172.600 ;
        RECT 15.600 166.200 16.400 177.800 ;
        RECT 23.600 177.600 24.400 178.400 ;
        RECT 18.800 170.200 19.600 175.800 ;
        RECT 23.700 172.400 24.300 177.600 ;
        RECT 25.300 176.400 25.900 185.600 ;
        RECT 26.800 183.600 27.600 184.400 ;
        RECT 33.200 184.200 34.000 195.800 ;
        RECT 38.100 186.400 38.700 203.600 ;
        RECT 42.900 194.400 43.500 223.600 ;
        RECT 54.100 222.400 54.700 243.600 ;
        RECT 55.600 233.600 56.400 234.400 ;
        RECT 55.700 230.200 56.300 233.600 ;
        RECT 55.600 229.400 56.400 230.200 ;
        RECT 55.600 225.600 56.400 226.400 ;
        RECT 54.000 221.600 54.800 222.400 ;
        RECT 52.400 219.600 53.200 220.400 ;
        RECT 44.400 206.200 45.200 217.800 ;
        RECT 52.500 212.600 53.100 219.600 ;
        RECT 52.400 211.800 53.200 212.600 ;
        RECT 54.000 206.200 54.800 217.800 ;
        RECT 55.700 214.400 56.300 225.600 ;
        RECT 57.200 224.200 58.000 235.800 ;
        RECT 60.400 226.200 61.200 231.800 ;
        RECT 62.000 226.200 62.800 231.800 ;
        RECT 65.200 224.200 66.000 235.800 ;
        RECT 66.900 230.200 67.500 243.600 ;
        RECT 66.800 229.400 67.600 230.200 ;
        RECT 70.000 227.600 70.800 228.400 ;
        RECT 65.200 221.600 66.000 222.400 ;
        RECT 55.600 213.600 56.400 214.400 ;
        RECT 57.200 210.200 58.000 215.800 ;
        RECT 58.800 210.200 59.600 215.800 ;
        RECT 62.000 206.200 62.800 217.800 ;
        RECT 65.300 212.400 65.900 221.600 ;
        RECT 70.100 214.400 70.700 227.600 ;
        RECT 74.800 224.200 75.600 235.800 ;
        RECT 79.700 232.400 80.300 263.600 ;
        RECT 81.300 252.400 81.900 283.600 ;
        RECT 82.800 269.600 83.600 270.400 ;
        RECT 82.900 266.400 83.500 269.600 ;
        RECT 86.100 268.400 86.700 291.600 ;
        RECT 90.800 289.600 91.600 290.400 ;
        RECT 94.000 290.200 94.600 293.600 ;
        RECT 98.000 293.400 98.800 293.600 ;
        RECT 95.600 291.600 96.400 292.400 ;
        RECT 94.000 289.400 94.800 290.200 ;
        RECT 95.700 276.400 96.300 291.600 ;
        RECT 100.800 290.200 101.400 295.000 ;
        RECT 102.000 293.600 102.800 294.400 ;
        RECT 100.600 289.400 101.400 290.200 ;
        RECT 95.600 275.600 96.400 276.400 ;
        RECT 87.400 271.800 88.200 272.600 ;
        RECT 94.000 271.800 94.800 272.600 ;
        RECT 84.400 267.600 85.200 268.400 ;
        RECT 86.000 267.600 86.800 268.400 ;
        RECT 87.400 267.000 88.000 271.800 ;
        RECT 90.000 268.400 90.800 268.600 ;
        RECT 94.200 268.400 94.800 271.800 ;
        RECT 95.700 268.400 96.300 275.600 ;
        RECT 97.200 269.600 98.000 270.400 ;
        RECT 90.000 267.800 94.800 268.400 ;
        RECT 89.200 267.000 90.000 267.200 ;
        RECT 92.600 267.000 93.400 267.200 ;
        RECT 94.200 267.000 94.800 267.800 ;
        RECT 95.600 267.600 96.400 268.400 ;
        RECT 98.800 267.600 99.600 268.400 ;
        RECT 102.000 267.600 102.800 268.400 ;
        RECT 82.800 265.600 83.600 266.400 ;
        RECT 87.400 266.200 88.200 267.000 ;
        RECT 89.200 266.400 93.400 267.000 ;
        RECT 94.000 266.200 94.800 267.000 ;
        RECT 100.400 265.600 101.200 266.400 ;
        RECT 102.000 265.600 102.800 266.400 ;
        RECT 92.400 263.600 93.200 264.400 ;
        RECT 92.500 262.400 93.100 263.600 ;
        RECT 92.400 261.600 93.200 262.400 ;
        RECT 90.800 257.600 91.600 258.400 ;
        RECT 90.900 256.400 91.500 257.600 ;
        RECT 90.800 255.600 91.600 256.400 ;
        RECT 82.800 253.600 83.600 254.400 ;
        RECT 87.600 253.600 88.400 254.400 ;
        RECT 82.900 252.400 83.500 253.600 ;
        RECT 81.200 251.600 82.000 252.400 ;
        RECT 82.800 251.600 83.600 252.400 ;
        RECT 92.500 250.300 93.100 261.600 ;
        RECT 102.100 260.400 102.700 265.600 ;
        RECT 102.000 259.600 102.800 260.400 ;
        RECT 94.000 255.600 94.800 256.400 ;
        RECT 97.200 253.600 98.000 254.400 ;
        RECT 102.000 253.600 102.800 254.400 ;
        RECT 97.300 252.400 97.900 253.600 ;
        RECT 103.700 252.400 104.300 295.700 ;
        RECT 106.900 295.700 109.100 296.300 ;
        RECT 106.900 294.400 107.500 295.700 ;
        RECT 113.200 295.600 114.000 296.400 ;
        RECT 105.200 293.600 106.000 294.400 ;
        RECT 106.800 293.600 107.600 294.400 ;
        RECT 108.400 293.600 109.200 294.400 ;
        RECT 113.200 293.600 114.000 294.400 ;
        RECT 105.300 268.300 105.900 293.600 ;
        RECT 108.500 292.400 109.100 293.600 ;
        RECT 106.800 291.600 107.600 292.400 ;
        RECT 108.400 291.600 109.200 292.400 ;
        RECT 106.900 270.400 107.500 291.600 ;
        RECT 113.300 290.400 113.900 293.600 ;
        RECT 113.200 289.600 114.000 290.400 ;
        RECT 116.500 288.400 117.100 305.600 ;
        RECT 118.100 304.400 118.700 307.600 ;
        RECT 124.500 306.400 125.100 311.600 ;
        RECT 130.900 308.400 131.500 319.600 ;
        RECT 137.200 313.600 138.000 314.400 ;
        RECT 137.300 312.400 137.900 313.600 ;
        RECT 137.200 311.600 138.000 312.400 ;
        RECT 143.600 311.600 144.400 312.400 ;
        RECT 150.000 311.600 150.800 312.400 ;
        RECT 151.600 311.600 152.400 312.400 ;
        RECT 153.200 311.600 154.000 312.400 ;
        RECT 158.100 312.300 158.700 331.600 ;
        RECT 167.700 312.400 168.300 331.600 ;
        RECT 175.600 330.200 176.200 333.600 ;
        RECT 179.600 333.400 180.400 333.600 ;
        RECT 182.400 330.200 183.000 335.000 ;
        RECT 183.700 334.400 184.300 347.600 ;
        RECT 186.800 344.200 187.600 355.800 ;
        RECT 190.100 354.300 190.700 363.600 ;
        RECT 194.800 359.600 195.600 360.400 ;
        RECT 190.100 353.700 192.300 354.300 ;
        RECT 190.000 346.200 190.800 351.800 ;
        RECT 191.700 350.400 192.300 353.700 ;
        RECT 191.600 349.600 192.400 350.400 ;
        RECT 194.900 346.400 195.500 359.600 ;
        RECT 201.300 354.400 201.900 363.600 ;
        RECT 201.200 353.600 202.000 354.400 ;
        RECT 215.600 353.600 216.400 354.400 ;
        RECT 198.200 351.800 199.000 352.600 ;
        RECT 196.400 349.600 197.200 350.400 ;
        RECT 196.400 347.600 197.200 348.400 ;
        RECT 198.200 347.000 198.800 351.800 ;
        RECT 199.600 351.600 200.400 352.400 ;
        RECT 204.400 351.800 205.200 352.600 ;
        RECT 199.400 349.800 200.200 350.600 ;
        RECT 199.600 348.400 200.200 349.800 ;
        RECT 204.600 348.400 205.200 351.800 ;
        RECT 207.600 351.600 208.400 352.400 ;
        RECT 207.700 348.400 208.300 351.600 ;
        RECT 209.200 349.600 210.000 350.400 ;
        RECT 214.000 349.600 214.800 350.400 ;
        RECT 214.100 348.400 214.700 349.600 ;
        RECT 199.600 347.800 205.200 348.400 ;
        RECT 199.600 347.000 200.400 347.200 ;
        RECT 203.000 347.000 203.800 347.200 ;
        RECT 204.600 347.000 205.200 347.800 ;
        RECT 206.000 347.600 206.800 348.400 ;
        RECT 207.600 347.600 208.400 348.400 ;
        RECT 209.200 347.600 210.000 348.400 ;
        RECT 214.000 347.600 214.800 348.400 ;
        RECT 198.200 346.400 203.800 347.000 ;
        RECT 194.800 345.600 195.600 346.400 ;
        RECT 198.200 346.200 199.000 346.400 ;
        RECT 204.400 346.200 205.200 347.000 ;
        RECT 194.900 344.400 195.500 345.600 ;
        RECT 194.800 343.600 195.600 344.400 ;
        RECT 206.100 338.400 206.700 347.600 ;
        RECT 209.300 346.400 209.900 347.600 ;
        RECT 215.700 346.400 216.300 353.600 ;
        RECT 218.800 348.300 219.600 348.400 ;
        RECT 220.500 348.300 221.100 373.600 ;
        RECT 222.000 369.600 222.800 370.400 ;
        RECT 223.700 366.400 224.300 373.600 ;
        RECT 225.200 369.600 226.000 370.400 ;
        RECT 231.800 370.200 232.400 375.000 ;
        RECT 233.200 374.800 234.000 375.000 ;
        RECT 236.600 374.800 237.400 375.000 ;
        RECT 238.200 374.200 238.800 375.000 ;
        RECT 239.700 374.400 240.300 375.600 ;
        RECT 233.200 373.600 238.800 374.200 ;
        RECT 239.600 373.600 240.400 374.400 ;
        RECT 233.200 372.200 233.800 373.600 ;
        RECT 233.000 371.400 233.800 372.200 ;
        RECT 238.200 370.200 238.800 373.600 ;
        RECT 225.300 368.400 225.900 369.600 ;
        RECT 231.800 369.400 232.600 370.200 ;
        RECT 238.000 369.400 238.800 370.200 ;
        RECT 239.600 369.600 240.400 370.400 ;
        RECT 225.200 367.600 226.000 368.400 ;
        RECT 223.600 365.600 224.400 366.400 ;
        RECT 223.700 358.400 224.300 365.600 ;
        RECT 223.600 357.600 224.400 358.400 ;
        RECT 223.800 351.800 224.600 352.600 ;
        RECT 230.000 351.800 230.800 352.600 ;
        RECT 239.700 352.400 240.300 369.600 ;
        RECT 241.300 368.400 241.900 391.700 ;
        RECT 242.900 388.400 243.500 393.600 ;
        RECT 242.800 387.600 243.600 388.400 ;
        RECT 244.500 386.400 245.100 413.600 ;
        RECT 247.600 406.200 248.400 417.800 ;
        RECT 255.600 415.600 256.400 416.400 ;
        RECT 255.700 412.600 256.300 415.600 ;
        RECT 249.200 411.600 250.000 412.400 ;
        RECT 255.600 411.800 256.400 412.600 ;
        RECT 249.300 410.400 249.900 411.600 ;
        RECT 249.200 409.600 250.000 410.400 ;
        RECT 255.700 402.400 256.300 411.800 ;
        RECT 257.200 406.200 258.000 417.800 ;
        RECT 260.400 410.200 261.200 415.800 ;
        RECT 266.800 413.600 267.600 414.400 ;
        RECT 270.000 413.600 270.800 414.400 ;
        RECT 271.600 413.600 272.400 414.400 ;
        RECT 265.200 411.600 266.000 412.400 ;
        RECT 266.900 404.400 267.500 413.600 ;
        RECT 266.800 404.300 267.600 404.400 ;
        RECT 266.800 403.700 269.100 404.300 ;
        RECT 266.800 403.600 267.600 403.700 ;
        RECT 254.000 401.600 254.800 402.400 ;
        RECT 255.600 401.600 256.400 402.400 ;
        RECT 247.600 393.600 248.400 394.400 ;
        RECT 247.700 388.400 248.300 393.600 ;
        RECT 254.100 392.400 254.700 401.600 ;
        RECT 254.000 391.600 254.800 392.400 ;
        RECT 257.000 391.800 257.800 392.600 ;
        RECT 263.600 391.800 264.400 392.600 ;
        RECT 249.200 389.600 250.000 390.400 ;
        RECT 254.000 389.600 254.800 390.400 ;
        RECT 247.600 387.600 248.400 388.400 ;
        RECT 244.400 385.600 245.200 386.400 ;
        RECT 249.300 384.400 249.900 389.600 ;
        RECT 254.100 386.400 254.700 389.600 ;
        RECT 255.600 387.600 256.400 388.400 ;
        RECT 255.700 386.400 256.300 387.600 ;
        RECT 257.000 387.000 257.600 391.800 ;
        RECT 259.600 388.400 260.400 388.600 ;
        RECT 263.800 388.400 264.400 391.800 ;
        RECT 266.800 391.600 267.600 392.400 ;
        RECT 259.600 387.800 264.400 388.400 ;
        RECT 258.800 387.000 259.600 387.200 ;
        RECT 262.200 387.000 263.000 387.200 ;
        RECT 263.800 387.000 264.400 387.800 ;
        RECT 265.200 387.600 266.000 388.400 ;
        RECT 254.000 385.600 254.800 386.400 ;
        RECT 255.600 385.600 256.400 386.400 ;
        RECT 257.000 386.200 257.800 387.000 ;
        RECT 258.800 386.400 263.000 387.000 ;
        RECT 263.600 386.200 264.400 387.000 ;
        RECT 246.000 383.600 246.800 384.400 ;
        RECT 249.200 383.600 250.000 384.400 ;
        RECT 252.400 383.600 253.200 384.400 ;
        RECT 246.000 381.600 246.800 382.400 ;
        RECT 246.100 378.400 246.700 381.600 ;
        RECT 252.500 378.400 253.100 383.600 ;
        RECT 254.100 382.400 254.700 385.600 ;
        RECT 258.800 383.600 259.600 384.400 ;
        RECT 254.000 381.600 254.800 382.400 ;
        RECT 258.900 380.400 259.500 383.600 ;
        RECT 258.800 379.600 259.600 380.400 ;
        RECT 262.000 379.600 262.800 380.400 ;
        RECT 262.100 378.400 262.700 379.600 ;
        RECT 242.800 377.600 243.600 378.400 ;
        RECT 246.000 377.600 246.800 378.400 ;
        RECT 252.400 377.600 253.200 378.400 ;
        RECT 262.000 377.600 262.800 378.400 ;
        RECT 242.900 376.400 243.500 377.600 ;
        RECT 242.800 375.600 243.600 376.400 ;
        RECT 250.800 373.600 251.600 374.400 ;
        RECT 252.500 372.400 253.100 377.600 ;
        RECT 255.600 375.600 256.400 376.400 ;
        RECT 255.700 372.400 256.300 375.600 ;
        RECT 257.200 373.600 258.000 374.400 ;
        RECT 257.300 372.400 257.900 373.600 ;
        RECT 244.400 371.600 245.200 372.400 ;
        RECT 249.200 371.600 250.000 372.400 ;
        RECT 252.400 371.600 253.200 372.400 ;
        RECT 255.600 371.600 256.400 372.400 ;
        RECT 257.200 371.600 258.000 372.400 ;
        RECT 262.000 371.600 262.800 372.400 ;
        RECT 241.200 367.600 242.000 368.400 ;
        RECT 244.400 361.600 245.200 362.400 ;
        RECT 244.500 358.400 245.100 361.600 ;
        RECT 249.300 358.400 249.900 371.600 ;
        RECT 255.700 370.400 256.300 371.600 ;
        RECT 262.100 370.400 262.700 371.600 ;
        RECT 255.600 369.600 256.400 370.400 ;
        RECT 262.000 369.600 262.800 370.400 ;
        RECT 263.600 369.600 264.400 370.400 ;
        RECT 263.700 368.400 264.300 369.600 ;
        RECT 250.800 367.600 251.600 368.400 ;
        RECT 255.600 367.600 256.400 368.400 ;
        RECT 263.600 367.600 264.400 368.400 ;
        RECT 250.900 358.400 251.500 367.600 ;
        RECT 265.300 366.300 265.900 387.600 ;
        RECT 266.900 380.400 267.500 391.600 ;
        RECT 266.800 379.600 267.600 380.400 ;
        RECT 268.500 374.400 269.100 403.700 ;
        RECT 270.100 390.400 270.700 413.600 ;
        RECT 273.200 411.600 274.000 412.400 ;
        RECT 274.800 411.600 275.600 412.400 ;
        RECT 273.300 398.400 273.900 411.600 ;
        RECT 273.200 397.600 274.000 398.400 ;
        RECT 271.600 391.600 272.400 392.400 ;
        RECT 274.900 390.400 275.500 411.600 ;
        RECT 276.400 409.600 277.200 410.400 ;
        RECT 276.500 392.400 277.100 409.600 ;
        RECT 278.000 405.600 278.800 406.400 ;
        RECT 282.800 406.200 283.600 417.800 ;
        RECT 292.400 406.200 293.200 417.800 ;
        RECT 294.000 413.600 294.800 414.400 ;
        RECT 295.600 410.200 296.400 415.800 ;
        RECT 302.000 413.600 302.800 414.400 ;
        RECT 319.600 409.600 320.400 410.400 ;
        RECT 300.400 407.600 301.200 408.400 ;
        RECT 300.500 398.400 301.100 407.600 ;
        RECT 316.400 404.300 317.200 404.400 ;
        RECT 316.400 403.700 318.700 404.300 ;
        RECT 316.400 403.600 317.200 403.700 ;
        RECT 305.200 399.600 306.000 400.400 ;
        RECT 305.300 398.400 305.900 399.600 ;
        RECT 278.000 397.600 278.800 398.400 ;
        RECT 300.400 397.600 301.200 398.400 ;
        RECT 305.200 397.600 306.000 398.400 ;
        RECT 316.400 397.600 317.200 398.400 ;
        RECT 276.400 391.600 277.200 392.400 ;
        RECT 270.000 389.600 270.800 390.400 ;
        RECT 274.800 389.600 275.600 390.400 ;
        RECT 270.100 388.400 270.700 389.600 ;
        RECT 270.000 387.600 270.800 388.400 ;
        RECT 274.800 387.600 275.600 388.400 ;
        RECT 276.400 387.600 277.200 388.400 ;
        RECT 271.600 385.600 272.400 386.400 ;
        RECT 271.700 378.400 272.300 385.600 ;
        RECT 273.200 383.600 274.000 384.400 ;
        RECT 270.000 377.600 270.800 378.400 ;
        RECT 271.600 377.600 272.400 378.400 ;
        RECT 270.100 376.400 270.700 377.600 ;
        RECT 270.000 375.600 270.800 376.400 ;
        RECT 273.300 374.400 273.900 383.600 ;
        RECT 276.500 378.400 277.100 387.600 ;
        RECT 276.400 377.600 277.200 378.400 ;
        RECT 278.100 376.400 278.700 397.600 ;
        RECT 279.600 391.600 280.400 392.400 ;
        RECT 281.200 391.600 282.000 392.400 ;
        RECT 284.200 391.800 285.000 392.600 ;
        RECT 290.800 391.800 291.600 392.600 ;
        RECT 274.800 375.600 275.600 376.400 ;
        RECT 278.000 375.600 278.800 376.400 ;
        RECT 268.400 373.600 269.200 374.400 ;
        RECT 273.200 373.600 274.000 374.400 ;
        RECT 274.900 372.400 275.500 375.600 ;
        RECT 266.800 371.600 267.600 372.400 ;
        RECT 274.800 371.600 275.600 372.400 ;
        RECT 276.400 371.600 277.200 372.400 ;
        RECT 278.100 370.400 278.700 375.600 ;
        RECT 279.700 374.400 280.300 391.600 ;
        RECT 281.300 390.400 281.900 391.600 ;
        RECT 281.200 389.600 282.000 390.400 ;
        RECT 282.800 387.600 283.600 388.400 ;
        RECT 281.200 383.600 282.000 384.400 ;
        RECT 279.600 373.600 280.400 374.400 ;
        RECT 278.000 369.600 278.800 370.400 ;
        RECT 263.700 365.700 265.900 366.300 ;
        RECT 244.400 357.600 245.200 358.400 ;
        RECT 249.200 357.600 250.000 358.400 ;
        RECT 250.800 357.600 251.600 358.400 ;
        RECT 262.000 357.600 262.800 358.400 ;
        RECT 218.800 347.700 221.100 348.300 ;
        RECT 218.800 347.600 219.600 347.700 ;
        RECT 222.000 347.600 222.800 348.400 ;
        RECT 218.900 346.400 219.500 347.600 ;
        RECT 223.800 347.000 224.400 351.800 ;
        RECT 225.000 349.800 225.800 350.600 ;
        RECT 225.200 348.400 225.800 349.800 ;
        RECT 228.400 349.600 229.200 350.400 ;
        RECT 230.200 348.400 230.800 351.800 ;
        RECT 233.200 351.600 234.000 352.400 ;
        RECT 239.600 351.600 240.400 352.400 ;
        RECT 231.600 349.600 232.400 350.400 ;
        RECT 236.400 349.600 237.200 350.400 ;
        RECT 231.700 348.400 232.300 349.600 ;
        RECT 244.500 348.400 245.100 357.600 ;
        RECT 247.600 351.600 248.400 352.400 ;
        RECT 255.600 351.600 256.400 352.400 ;
        RECT 247.600 349.600 248.400 350.400 ;
        RECT 249.200 349.600 250.000 350.400 ;
        RECT 225.200 347.800 230.800 348.400 ;
        RECT 225.200 347.000 226.000 347.200 ;
        RECT 228.600 347.000 229.400 347.200 ;
        RECT 230.200 347.000 230.800 347.800 ;
        RECT 231.600 347.600 232.400 348.400 ;
        RECT 238.000 347.600 238.800 348.400 ;
        RECT 242.800 347.600 243.600 348.400 ;
        RECT 244.400 347.600 245.200 348.400 ;
        RECT 223.800 346.400 229.400 347.000 ;
        RECT 209.200 345.600 210.000 346.400 ;
        RECT 215.600 345.600 216.400 346.400 ;
        RECT 218.800 345.600 219.600 346.400 ;
        RECT 223.800 346.200 224.600 346.400 ;
        RECT 230.000 346.200 230.800 347.000 ;
        RECT 231.700 346.400 232.300 347.600 ;
        RECT 231.600 345.600 232.400 346.400 ;
        RECT 225.200 343.600 226.000 344.400 ;
        RECT 231.700 344.300 232.300 345.600 ;
        RECT 230.100 343.700 232.300 344.300 ;
        RECT 183.600 333.600 184.400 334.400 ;
        RECT 175.600 329.400 176.400 330.200 ;
        RECT 182.200 329.400 183.000 330.200 ;
        RECT 204.400 326.200 205.200 337.800 ;
        RECT 206.000 337.600 206.800 338.400 ;
        RECT 210.800 333.600 211.600 334.400 ;
        RECT 172.400 323.600 173.200 324.400 ;
        RECT 186.800 323.600 187.600 324.400 ;
        RECT 199.600 323.600 200.400 324.400 ;
        RECT 156.500 311.700 158.700 312.300 ;
        RECT 143.700 310.400 144.300 311.600 ;
        RECT 150.100 310.400 150.700 311.600 ;
        RECT 132.400 309.600 133.200 310.400 ;
        RECT 134.000 309.600 134.800 310.400 ;
        RECT 143.600 309.600 144.400 310.400 ;
        RECT 150.000 309.600 150.800 310.400 ;
        RECT 130.800 307.600 131.600 308.400 ;
        RECT 134.100 306.400 134.700 309.600 ;
        RECT 151.700 308.400 152.300 311.600 ;
        RECT 142.000 307.600 142.800 308.400 ;
        RECT 145.200 307.600 146.000 308.400 ;
        RECT 146.800 307.600 147.600 308.400 ;
        RECT 151.600 307.600 152.400 308.400 ;
        RECT 124.400 305.600 125.200 306.400 ;
        RECT 134.000 305.600 134.800 306.400 ;
        RECT 118.000 303.600 118.800 304.400 ;
        RECT 121.200 303.600 122.000 304.400 ;
        RECT 126.000 303.600 126.800 304.400 ;
        RECT 127.600 303.600 128.400 304.400 ;
        RECT 129.200 303.600 130.000 304.400 ;
        RECT 119.600 295.600 120.400 296.400 ;
        RECT 119.700 294.400 120.300 295.600 ;
        RECT 119.600 293.600 120.400 294.400 ;
        RECT 121.300 292.400 121.900 303.600 ;
        RECT 122.800 293.600 123.600 294.400 ;
        RECT 126.100 292.400 126.700 303.600 ;
        RECT 127.700 294.400 128.300 303.600 ;
        RECT 129.300 302.400 129.900 303.600 ;
        RECT 129.200 301.600 130.000 302.400 ;
        RECT 137.200 297.600 138.000 298.400 ;
        RECT 130.800 295.600 131.600 296.400 ;
        RECT 132.400 295.600 133.200 296.400 ;
        RECT 127.600 293.600 128.400 294.400 ;
        RECT 129.200 293.600 130.000 294.400 ;
        RECT 121.200 291.600 122.000 292.400 ;
        RECT 126.000 291.600 126.800 292.400 ;
        RECT 122.800 289.600 123.600 290.400 ;
        RECT 116.400 287.600 117.200 288.400 ;
        RECT 108.400 285.600 109.200 286.400 ;
        RECT 122.900 284.400 123.500 289.600 ;
        RECT 129.300 286.400 129.900 293.600 ;
        RECT 132.500 290.400 133.100 295.600 ;
        RECT 137.300 292.400 137.900 297.600 ;
        RECT 137.200 291.600 138.000 292.400 ;
        RECT 132.400 289.600 133.200 290.400 ;
        RECT 132.400 287.600 133.200 288.400 ;
        RECT 129.200 285.600 130.000 286.400 ;
        RECT 111.600 283.600 112.400 284.400 ;
        RECT 116.400 283.600 117.200 284.400 ;
        RECT 122.800 283.600 123.600 284.400 ;
        RECT 108.400 279.600 109.200 280.400 ;
        RECT 106.800 269.600 107.600 270.400 ;
        RECT 105.300 267.700 107.500 268.300 ;
        RECT 106.900 266.400 107.500 267.700 ;
        RECT 105.200 265.600 106.000 266.400 ;
        RECT 106.800 265.600 107.600 266.400 ;
        RECT 105.300 254.400 105.900 265.600 ;
        RECT 105.200 253.600 106.000 254.400 ;
        RECT 97.200 251.600 98.000 252.400 ;
        RECT 103.600 251.600 104.400 252.400 ;
        RECT 94.000 250.300 94.800 250.400 ;
        RECT 92.500 249.700 94.800 250.300 ;
        RECT 94.000 249.600 94.800 249.700 ;
        RECT 90.800 247.600 91.600 248.400 ;
        RECT 98.800 247.600 99.600 248.400 ;
        RECT 103.600 247.600 104.400 248.400 ;
        RECT 84.400 233.600 85.200 234.400 ;
        RECT 79.600 231.600 80.400 232.400 ;
        RECT 82.600 231.800 83.400 232.600 ;
        RECT 89.200 231.800 90.000 232.600 ;
        RECT 81.200 227.600 82.000 228.400 ;
        RECT 82.600 227.000 83.200 231.800 ;
        RECT 85.200 228.400 86.000 228.600 ;
        RECT 89.400 228.400 90.000 231.800 ;
        RECT 90.900 228.400 91.500 247.600 ;
        RECT 97.200 243.600 98.000 244.400 ;
        RECT 92.400 231.600 93.200 232.400 ;
        RECT 85.200 227.800 90.000 228.400 ;
        RECT 84.400 227.000 85.200 227.200 ;
        RECT 87.800 227.000 88.600 227.200 ;
        RECT 89.400 227.000 90.000 227.800 ;
        RECT 90.800 227.600 91.600 228.400 ;
        RECT 95.600 228.300 96.400 228.400 ;
        RECT 97.300 228.300 97.900 243.600 ;
        RECT 95.600 227.700 97.900 228.300 ;
        RECT 95.600 227.600 96.400 227.700 ;
        RECT 82.600 226.200 83.400 227.000 ;
        RECT 84.400 226.400 88.600 227.000 ;
        RECT 89.200 226.200 90.000 227.000 ;
        RECT 79.600 223.600 80.400 224.400 ;
        RECT 92.400 223.600 93.200 224.400 ;
        RECT 97.200 223.600 98.000 224.400 ;
        RECT 102.000 224.200 102.800 235.800 ;
        RECT 106.800 227.600 107.600 228.400 ;
        RECT 92.500 220.300 93.100 223.600 ;
        RECT 97.300 222.400 97.900 223.600 ;
        RECT 97.200 221.600 98.000 222.400 ;
        RECT 103.600 221.600 104.400 222.400 ;
        RECT 90.900 219.700 93.100 220.300 ;
        RECT 70.000 213.600 70.800 214.400 ;
        RECT 70.100 212.400 70.700 213.600 ;
        RECT 65.200 211.600 66.000 212.400 ;
        RECT 70.000 211.600 70.800 212.400 ;
        RECT 71.600 206.200 72.400 217.800 ;
        RECT 82.800 206.200 83.600 217.800 ;
        RECT 90.900 212.600 91.500 219.700 ;
        RECT 90.800 211.800 91.600 212.600 ;
        RECT 92.400 206.200 93.200 217.800 ;
        RECT 94.000 213.600 94.800 214.400 ;
        RECT 95.600 210.200 96.400 215.800 ;
        RECT 97.200 213.600 98.000 214.400 ;
        RECT 44.400 203.600 45.200 204.400 ;
        RECT 76.400 203.600 77.200 204.400 ;
        RECT 78.000 204.300 78.800 204.400 ;
        RECT 78.000 203.700 80.300 204.300 ;
        RECT 78.000 203.600 78.800 203.700 ;
        RECT 42.800 193.600 43.600 194.400 ;
        RECT 39.600 191.600 40.400 192.400 ;
        RECT 42.800 191.600 43.600 192.400 ;
        RECT 39.700 190.400 40.300 191.600 ;
        RECT 39.600 189.600 40.400 190.400 ;
        RECT 42.900 188.400 43.500 191.600 ;
        RECT 44.500 188.400 45.100 203.600 ;
        RECT 76.500 196.400 77.100 203.600 ;
        RECT 76.400 195.600 77.200 196.400 ;
        RECT 49.200 191.600 50.000 192.400 ;
        RECT 55.600 191.600 56.400 192.400 ;
        RECT 60.400 191.600 61.200 192.400 ;
        RECT 65.200 191.600 66.000 192.400 ;
        RECT 68.400 191.600 69.200 192.400 ;
        RECT 78.000 191.600 78.800 192.400 ;
        RECT 54.000 189.600 54.800 190.400 ;
        RECT 42.800 187.600 43.600 188.400 ;
        RECT 44.400 187.600 45.200 188.400 ;
        RECT 46.000 187.600 46.800 188.400 ;
        RECT 44.500 186.400 45.100 187.600 ;
        RECT 46.100 186.400 46.700 187.600 ;
        RECT 38.000 185.600 38.800 186.400 ;
        RECT 44.400 185.600 45.200 186.400 ;
        RECT 46.000 185.600 46.800 186.400 ;
        RECT 50.800 185.600 51.600 186.400 ;
        RECT 38.000 183.600 38.800 184.400 ;
        RECT 39.600 183.600 40.400 184.400 ;
        RECT 25.200 175.600 26.000 176.400 ;
        RECT 22.000 171.600 22.800 172.400 ;
        RECT 23.600 171.600 24.400 172.400 ;
        RECT 20.400 169.600 21.200 170.400 ;
        RECT 20.500 158.400 21.100 169.600 ;
        RECT 18.800 157.600 19.600 158.400 ;
        RECT 20.400 157.600 21.200 158.400 ;
        RECT 18.900 152.400 19.500 157.600 ;
        RECT 22.100 154.400 22.700 171.600 ;
        RECT 23.600 155.600 24.400 156.400 ;
        RECT 22.000 153.600 22.800 154.400 ;
        RECT 12.400 151.600 13.200 152.400 ;
        RECT 18.800 151.600 19.600 152.400 ;
        RECT 2.800 149.600 3.600 150.400 ;
        RECT 7.600 149.600 8.400 150.400 ;
        RECT 10.800 149.600 11.600 150.400 ;
        RECT 15.600 149.600 16.400 150.400 ;
        RECT 20.400 149.600 21.200 150.400 ;
        RECT 1.200 147.600 2.000 148.400 ;
        RECT 1.300 136.400 1.900 147.600 ;
        RECT 2.900 146.300 3.500 149.600 ;
        RECT 7.700 146.400 8.300 149.600 ;
        RECT 9.200 147.600 10.000 148.400 ;
        RECT 7.600 146.300 8.400 146.400 ;
        RECT 2.900 145.700 5.100 146.300 ;
        RECT 1.200 135.600 2.000 136.400 ;
        RECT 1.200 127.600 2.000 128.400 ;
        RECT 1.300 110.400 1.900 127.600 ;
        RECT 2.900 110.400 3.500 145.700 ;
        RECT 4.500 134.400 5.100 145.700 ;
        RECT 6.100 145.700 8.400 146.300 ;
        RECT 6.100 144.400 6.700 145.700 ;
        RECT 7.600 145.600 8.400 145.700 ;
        RECT 6.000 143.600 6.800 144.400 ;
        RECT 7.600 135.600 8.400 136.400 ;
        RECT 9.300 134.400 9.900 147.600 ;
        RECT 4.400 133.600 5.200 134.400 ;
        RECT 9.200 133.600 10.000 134.400 ;
        RECT 4.500 132.400 5.100 133.600 ;
        RECT 10.900 132.400 11.500 149.600 ;
        RECT 14.000 148.300 14.800 148.400 ;
        RECT 14.000 147.700 16.300 148.300 ;
        RECT 14.000 147.600 14.800 147.700 ;
        RECT 14.000 137.600 14.800 138.400 ;
        RECT 4.400 131.600 5.200 132.400 ;
        RECT 10.800 131.600 11.600 132.400 ;
        RECT 14.100 130.400 14.700 137.600 ;
        RECT 15.700 136.400 16.300 147.700 ;
        RECT 20.500 146.400 21.100 149.600 ;
        RECT 23.700 148.400 24.300 155.600 ;
        RECT 25.300 150.400 25.900 175.600 ;
        RECT 26.900 174.400 27.500 183.600 ;
        RECT 39.700 178.400 40.300 183.600 ;
        RECT 39.600 177.600 40.400 178.400 ;
        RECT 28.400 175.000 29.200 175.800 ;
        RECT 30.000 175.600 30.800 176.400 ;
        RECT 29.800 175.000 34.000 175.600 ;
        RECT 35.000 175.000 35.800 175.800 ;
        RECT 26.800 173.600 27.600 174.400 ;
        RECT 28.400 174.200 29.000 175.000 ;
        RECT 29.800 174.800 30.600 175.000 ;
        RECT 33.200 174.800 34.000 175.000 ;
        RECT 28.400 173.600 33.200 174.200 ;
        RECT 26.900 156.400 27.500 173.600 ;
        RECT 28.400 170.200 29.000 173.600 ;
        RECT 32.400 173.400 33.200 173.600 ;
        RECT 33.200 171.600 34.000 172.400 ;
        RECT 28.400 169.400 29.200 170.200 ;
        RECT 33.300 168.400 33.900 171.600 ;
        RECT 35.200 170.200 35.800 175.000 ;
        RECT 39.600 175.000 40.400 175.800 ;
        RECT 41.000 175.000 45.200 175.600 ;
        RECT 46.200 175.000 47.000 175.800 ;
        RECT 38.000 173.600 38.800 174.400 ;
        RECT 39.600 174.200 40.200 175.000 ;
        RECT 41.000 174.800 41.800 175.000 ;
        RECT 44.400 174.800 45.200 175.000 ;
        RECT 39.600 173.600 44.400 174.200 ;
        RECT 38.100 172.400 38.700 173.600 ;
        RECT 38.000 171.600 38.800 172.400 ;
        RECT 35.000 169.400 35.800 170.200 ;
        RECT 39.600 170.200 40.200 173.600 ;
        RECT 43.600 173.400 44.400 173.600 ;
        RECT 41.200 171.600 42.000 172.400 ;
        RECT 39.600 169.400 40.400 170.200 ;
        RECT 33.200 167.600 34.000 168.400 ;
        RECT 33.300 158.400 33.900 167.600 ;
        RECT 41.300 158.400 41.900 171.600 ;
        RECT 46.400 170.200 47.000 175.000 ;
        RECT 47.600 173.600 48.400 174.400 ;
        RECT 47.600 171.600 48.400 172.400 ;
        RECT 50.900 172.300 51.500 185.600 ;
        RECT 52.400 183.600 53.200 184.400 ;
        RECT 52.500 176.400 53.100 183.600 ;
        RECT 52.400 175.600 53.200 176.400 ;
        RECT 54.100 174.400 54.700 189.600 ;
        RECT 60.500 186.400 61.100 191.600 ;
        RECT 65.300 190.400 65.900 191.600 ;
        RECT 68.500 190.400 69.100 191.600 ;
        RECT 63.600 189.600 64.400 190.400 ;
        RECT 65.200 189.600 66.000 190.400 ;
        RECT 66.800 189.600 67.600 190.400 ;
        RECT 68.400 189.600 69.200 190.400 ;
        RECT 63.600 187.600 64.400 188.400 ;
        RECT 60.400 185.600 61.200 186.400 ;
        RECT 57.200 183.600 58.000 184.400 ;
        RECT 62.000 183.600 62.800 184.400 ;
        RECT 55.600 175.600 56.400 176.400 ;
        RECT 54.000 173.600 54.800 174.400 ;
        RECT 57.300 172.400 57.900 183.600 ;
        RECT 60.400 175.600 61.200 176.400 ;
        RECT 58.800 173.600 59.600 174.400 ;
        RECT 52.400 172.300 53.200 172.400 ;
        RECT 50.900 171.700 53.200 172.300 ;
        RECT 52.400 171.600 53.200 171.700 ;
        RECT 57.200 171.600 58.000 172.400 ;
        RECT 46.200 169.400 47.000 170.200 ;
        RECT 44.400 165.600 45.200 166.400 ;
        RECT 33.200 157.600 34.000 158.400 ;
        RECT 41.200 157.600 42.000 158.400 ;
        RECT 26.800 155.600 27.600 156.400 ;
        RECT 31.600 151.600 32.400 152.400 ;
        RECT 33.200 151.600 34.000 152.400 ;
        RECT 36.400 151.600 37.200 152.400 ;
        RECT 31.700 150.400 32.300 151.600 ;
        RECT 33.300 150.400 33.900 151.600 ;
        RECT 36.500 150.400 37.100 151.600 ;
        RECT 47.700 150.400 48.300 171.600 ;
        RECT 58.900 170.400 59.500 173.600 ;
        RECT 60.500 172.400 61.100 175.600 ;
        RECT 60.400 171.600 61.200 172.400 ;
        RECT 62.100 170.400 62.700 183.600 ;
        RECT 66.900 174.400 67.500 189.600 ;
        RECT 70.000 187.600 70.800 188.400 ;
        RECT 71.600 187.600 72.400 188.400 ;
        RECT 73.200 188.000 74.000 188.800 ;
        RECT 70.100 174.400 70.700 187.600 ;
        RECT 71.700 176.400 72.300 187.600 ;
        RECT 73.300 186.400 73.900 188.000 ;
        RECT 73.200 185.600 74.000 186.400 ;
        RECT 74.800 185.600 75.600 186.400 ;
        RECT 78.000 185.600 78.800 186.400 ;
        RECT 71.600 175.600 72.400 176.400 ;
        RECT 74.900 174.400 75.500 185.600 ;
        RECT 76.400 183.600 77.200 184.400 ;
        RECT 66.800 173.600 67.600 174.400 ;
        RECT 70.000 173.600 70.800 174.400 ;
        RECT 74.800 173.600 75.600 174.400 ;
        RECT 74.900 172.400 75.500 173.600 ;
        RECT 76.500 172.400 77.100 183.600 ;
        RECT 63.600 171.600 64.400 172.400 ;
        RECT 65.200 171.600 66.000 172.400 ;
        RECT 70.000 171.600 70.800 172.400 ;
        RECT 74.800 171.600 75.600 172.400 ;
        RECT 76.400 171.600 77.200 172.400 ;
        RECT 49.200 169.600 50.000 170.400 ;
        RECT 58.800 169.600 59.600 170.400 ;
        RECT 62.000 169.600 62.800 170.400 ;
        RECT 49.300 168.400 49.900 169.600 ;
        RECT 49.200 167.600 50.000 168.400 ;
        RECT 55.600 163.600 56.400 164.400 ;
        RECT 49.200 153.600 50.000 154.400 ;
        RECT 49.300 152.400 49.900 153.600 ;
        RECT 55.700 152.400 56.300 163.600 ;
        RECT 63.700 154.400 64.300 171.600 ;
        RECT 78.000 167.600 78.800 168.400 ;
        RECT 63.600 153.600 64.400 154.400 ;
        RECT 74.800 153.600 75.600 154.400 ;
        RECT 49.200 152.300 50.000 152.400 ;
        RECT 49.200 151.700 51.500 152.300 ;
        RECT 49.200 151.600 50.000 151.700 ;
        RECT 25.200 149.600 26.000 150.400 ;
        RECT 28.400 149.600 29.200 150.400 ;
        RECT 31.600 149.600 32.400 150.400 ;
        RECT 33.200 149.600 34.000 150.400 ;
        RECT 36.400 149.600 37.200 150.400 ;
        RECT 41.200 149.600 42.000 150.400 ;
        RECT 47.600 149.600 48.400 150.400 ;
        RECT 49.200 149.600 50.000 150.400 ;
        RECT 23.600 147.600 24.400 148.400 ;
        RECT 18.800 145.600 19.600 146.400 ;
        RECT 20.400 145.600 21.200 146.400 ;
        RECT 18.800 143.600 19.600 144.400 ;
        RECT 15.600 135.600 16.400 136.400 ;
        RECT 14.000 129.600 14.800 130.400 ;
        RECT 14.000 125.600 14.800 126.400 ;
        RECT 4.400 123.600 5.200 124.400 ;
        RECT 10.800 123.600 11.600 124.400 ;
        RECT 1.200 109.600 2.000 110.400 ;
        RECT 2.800 109.600 3.600 110.400 ;
        RECT 1.300 108.400 1.900 109.600 ;
        RECT 2.900 108.400 3.500 109.600 ;
        RECT 1.200 107.600 2.000 108.400 ;
        RECT 2.800 107.600 3.600 108.400 ;
        RECT 2.900 104.300 3.500 107.600 ;
        RECT 1.300 103.700 3.500 104.300 ;
        RECT 1.300 94.400 1.900 103.700 ;
        RECT 2.800 101.600 3.600 102.400 ;
        RECT 2.900 98.400 3.500 101.600 ;
        RECT 2.800 97.600 3.600 98.400 ;
        RECT 4.500 96.400 5.100 123.600 ;
        RECT 10.900 112.400 11.500 123.600 ;
        RECT 12.400 115.600 13.200 116.400 ;
        RECT 6.000 111.600 6.800 112.400 ;
        RECT 10.800 111.600 11.600 112.400 ;
        RECT 7.600 109.600 8.400 110.400 ;
        RECT 12.500 108.400 13.100 115.600 ;
        RECT 14.100 110.400 14.700 125.600 ;
        RECT 14.000 109.600 14.800 110.400 ;
        RECT 18.900 108.400 19.500 143.600 ;
        RECT 20.500 132.400 21.100 145.600 ;
        RECT 22.000 143.600 22.800 144.400 ;
        RECT 20.400 131.600 21.200 132.400 ;
        RECT 22.100 126.400 22.700 143.600 ;
        RECT 23.700 136.400 24.300 147.600 ;
        RECT 25.300 142.400 25.900 149.600 ;
        RECT 31.700 148.400 32.300 149.600 ;
        RECT 30.000 147.600 30.800 148.400 ;
        RECT 31.600 147.600 32.400 148.400 ;
        RECT 38.000 147.600 38.800 148.400 ;
        RECT 39.600 147.600 40.400 148.400 ;
        RECT 26.800 145.600 27.600 146.400 ;
        RECT 25.200 141.600 26.000 142.400 ;
        RECT 26.900 138.400 27.500 145.600 ;
        RECT 30.100 138.400 30.700 147.600 ;
        RECT 38.100 146.400 38.700 147.600 ;
        RECT 39.700 146.400 40.300 147.600 ;
        RECT 38.000 145.600 38.800 146.400 ;
        RECT 39.600 145.600 40.400 146.400 ;
        RECT 41.300 144.400 41.900 149.600 ;
        RECT 46.000 147.600 46.800 148.400 ;
        RECT 46.100 146.400 46.700 147.600 ;
        RECT 46.000 145.600 46.800 146.400 ;
        RECT 33.200 143.600 34.000 144.400 ;
        RECT 41.200 143.600 42.000 144.400 ;
        RECT 44.400 143.600 45.200 144.400 ;
        RECT 33.300 140.400 33.900 143.600 ;
        RECT 34.800 141.600 35.600 142.400 ;
        RECT 33.200 139.600 34.000 140.400 ;
        RECT 26.800 137.600 27.600 138.400 ;
        RECT 30.000 137.600 30.800 138.400 ;
        RECT 30.100 136.400 30.700 137.600 ;
        RECT 34.900 136.400 35.500 141.600 ;
        RECT 44.500 138.400 45.100 143.600 ;
        RECT 44.400 137.600 45.200 138.400 ;
        RECT 23.600 135.600 24.400 136.400 ;
        RECT 28.400 135.600 29.200 136.400 ;
        RECT 30.000 135.600 30.800 136.400 ;
        RECT 33.200 135.600 34.000 136.400 ;
        RECT 34.800 135.600 35.600 136.400 ;
        RECT 38.000 135.600 38.800 136.400 ;
        RECT 28.500 134.400 29.100 135.600 ;
        RECT 28.400 133.600 29.200 134.400 ;
        RECT 23.600 131.600 24.400 132.400 ;
        RECT 25.200 131.600 26.000 132.400 ;
        RECT 30.000 131.600 30.800 132.400 ;
        RECT 25.300 128.400 25.900 131.600 ;
        RECT 30.100 130.400 30.700 131.600 ;
        RECT 30.000 129.600 30.800 130.400 ;
        RECT 25.200 127.600 26.000 128.400 ;
        RECT 22.000 125.600 22.800 126.400 ;
        RECT 22.000 123.600 22.800 124.400 ;
        RECT 22.100 110.400 22.700 123.600 ;
        RECT 23.400 111.800 24.200 112.600 ;
        RECT 30.000 111.800 30.800 112.600 ;
        RECT 22.000 109.600 22.800 110.400 ;
        RECT 9.200 107.600 10.000 108.400 ;
        RECT 12.400 107.600 13.200 108.400 ;
        RECT 18.800 107.600 19.600 108.400 ;
        RECT 22.000 107.600 22.800 108.400 ;
        RECT 6.000 105.600 6.800 106.400 ;
        RECT 9.300 102.400 9.900 107.600 ;
        RECT 23.400 107.000 24.000 111.800 ;
        RECT 26.000 108.400 26.800 108.600 ;
        RECT 30.200 108.400 30.800 111.800 ;
        RECT 33.300 110.400 33.900 135.600 ;
        RECT 38.100 134.400 38.700 135.600 ;
        RECT 38.000 133.600 38.800 134.400 ;
        RECT 44.500 132.400 45.100 137.600 ;
        RECT 44.400 131.600 45.200 132.400 ;
        RECT 38.000 129.600 38.800 130.400 ;
        RECT 41.200 129.600 42.000 130.400 ;
        RECT 41.200 113.600 42.000 114.400 ;
        RECT 36.400 111.600 37.200 112.400 ;
        RECT 36.500 110.400 37.100 111.600 ;
        RECT 31.600 109.600 32.400 110.400 ;
        RECT 33.200 109.600 34.000 110.400 ;
        RECT 36.400 109.600 37.200 110.400 ;
        RECT 38.000 109.600 38.800 110.400 ;
        RECT 26.000 107.800 30.800 108.400 ;
        RECT 25.200 107.000 26.000 107.200 ;
        RECT 28.600 107.000 29.400 107.200 ;
        RECT 30.200 107.000 30.800 107.800 ;
        RECT 15.600 105.600 16.400 106.400 ;
        RECT 23.400 106.200 24.200 107.000 ;
        RECT 25.200 106.400 29.400 107.000 ;
        RECT 30.000 106.200 30.800 107.000 ;
        RECT 12.400 103.600 13.200 104.400 ;
        RECT 17.200 103.600 18.000 104.400 ;
        RECT 28.400 103.600 29.200 104.400 ;
        RECT 9.200 101.600 10.000 102.400 ;
        RECT 4.400 95.600 5.200 96.400 ;
        RECT 1.200 93.600 2.000 94.400 ;
        RECT 1.300 68.400 1.900 93.600 ;
        RECT 9.200 91.600 10.000 92.400 ;
        RECT 10.800 91.600 11.600 92.400 ;
        RECT 9.300 86.300 9.900 91.600 ;
        RECT 10.900 88.400 11.500 91.600 ;
        RECT 10.800 87.600 11.600 88.400 ;
        RECT 9.300 85.700 11.500 86.300 ;
        RECT 9.200 83.600 10.000 84.400 ;
        RECT 9.300 76.400 9.900 83.600 ;
        RECT 9.200 75.600 10.000 76.400 ;
        RECT 2.600 71.800 3.400 72.600 ;
        RECT 9.200 71.800 10.000 72.600 ;
        RECT 1.200 67.600 2.000 68.400 ;
        RECT 2.600 67.000 3.200 71.800 ;
        RECT 5.200 68.400 6.000 68.600 ;
        RECT 9.400 68.400 10.000 71.800 ;
        RECT 5.200 67.800 10.000 68.400 ;
        RECT 4.400 67.000 5.200 67.200 ;
        RECT 7.800 67.000 8.600 67.200 ;
        RECT 9.400 67.000 10.000 67.800 ;
        RECT 2.600 66.200 3.400 67.000 ;
        RECT 4.400 66.400 8.600 67.000 ;
        RECT 7.600 65.600 8.400 66.400 ;
        RECT 9.200 66.200 10.000 67.000 ;
        RECT 4.400 63.600 5.200 64.400 ;
        RECT 2.800 57.600 3.600 58.400 ;
        RECT 4.500 56.400 5.100 63.600 ;
        RECT 9.200 59.600 10.000 60.400 ;
        RECT 9.300 58.400 9.900 59.600 ;
        RECT 10.900 58.400 11.500 85.700 ;
        RECT 12.500 74.400 13.100 103.600 ;
        RECT 14.000 99.600 14.800 100.400 ;
        RECT 14.100 94.400 14.700 99.600 ;
        RECT 14.000 94.300 14.800 94.400 ;
        RECT 14.000 93.700 16.300 94.300 ;
        RECT 14.000 93.600 14.800 93.700 ;
        RECT 14.000 91.600 14.800 92.400 ;
        RECT 14.100 80.400 14.700 91.600 ;
        RECT 14.000 79.600 14.800 80.400 ;
        RECT 12.400 73.600 13.200 74.400 ;
        RECT 12.400 71.600 13.200 72.400 ;
        RECT 14.100 70.400 14.700 79.600 ;
        RECT 15.700 72.400 16.300 93.700 ;
        RECT 17.300 82.400 17.900 103.600 ;
        RECT 18.800 101.600 19.600 102.400 ;
        RECT 22.000 101.600 22.800 102.400 ;
        RECT 18.900 90.400 19.500 101.600 ;
        RECT 22.100 98.400 22.700 101.600 ;
        RECT 28.500 98.400 29.100 103.600 ;
        RECT 22.000 97.600 22.800 98.400 ;
        RECT 28.400 97.600 29.200 98.400 ;
        RECT 31.700 96.400 32.300 109.600 ;
        RECT 38.100 108.400 38.700 109.600 ;
        RECT 41.300 108.400 41.900 113.600 ;
        RECT 46.100 112.400 46.700 145.600 ;
        RECT 47.600 141.600 48.400 142.400 ;
        RECT 47.700 134.400 48.300 141.600 ;
        RECT 49.300 138.400 49.900 149.600 ;
        RECT 50.900 148.400 51.500 151.700 ;
        RECT 54.000 151.600 54.800 152.400 ;
        RECT 55.600 151.600 56.400 152.400 ;
        RECT 60.400 151.600 61.200 152.400 ;
        RECT 66.800 152.300 67.600 152.400 ;
        RECT 65.300 151.700 67.600 152.300 ;
        RECT 50.800 147.600 51.600 148.400 ;
        RECT 54.100 148.300 54.700 151.600 ;
        RECT 55.700 150.400 56.300 151.600 ;
        RECT 60.500 150.400 61.100 151.600 ;
        RECT 55.600 149.600 56.400 150.400 ;
        RECT 60.400 149.600 61.200 150.400 ;
        RECT 55.600 148.300 56.400 148.400 ;
        RECT 54.100 147.700 56.400 148.300 ;
        RECT 55.600 147.600 56.400 147.700 ;
        RECT 62.000 147.600 62.800 148.400 ;
        RECT 55.700 144.400 56.300 147.600 ;
        RECT 62.100 146.400 62.700 147.600 ;
        RECT 58.800 145.600 59.600 146.400 ;
        RECT 62.000 145.600 62.800 146.400 ;
        RECT 54.000 143.600 54.800 144.400 ;
        RECT 55.600 143.600 56.400 144.400 ;
        RECT 49.200 137.600 50.000 138.400 ;
        RECT 47.600 133.600 48.400 134.400 ;
        RECT 52.400 133.600 53.200 134.400 ;
        RECT 52.500 130.400 53.100 133.600 ;
        RECT 54.100 130.400 54.700 143.600 ;
        RECT 58.900 134.400 59.500 145.600 ;
        RECT 65.300 144.400 65.900 151.700 ;
        RECT 66.800 151.600 67.600 151.700 ;
        RECT 70.000 151.800 70.800 152.600 ;
        RECT 74.900 152.400 75.500 153.600 ;
        RECT 70.000 148.400 70.600 151.800 ;
        RECT 74.800 151.600 75.600 152.400 ;
        RECT 76.600 151.800 77.400 152.600 ;
        RECT 74.000 148.400 74.800 148.600 ;
        RECT 68.400 147.600 69.200 148.400 ;
        RECT 70.000 147.800 74.800 148.400 ;
        RECT 70.000 147.000 70.600 147.800 ;
        RECT 71.400 147.000 72.200 147.200 ;
        RECT 74.800 147.000 75.600 147.200 ;
        RECT 76.800 147.000 77.400 151.800 ;
        RECT 79.700 150.400 80.300 203.700 ;
        RECT 87.600 195.600 88.400 196.400 ;
        RECT 87.700 192.400 88.300 195.600 ;
        RECT 103.700 192.400 104.300 221.600 ;
        RECT 106.900 214.400 107.500 227.600 ;
        RECT 106.800 213.600 107.600 214.400 ;
        RECT 86.000 191.600 86.800 192.400 ;
        RECT 87.600 191.600 88.400 192.400 ;
        RECT 103.600 191.600 104.400 192.400 ;
        RECT 87.700 186.400 88.300 191.600 ;
        RECT 94.000 189.600 94.800 190.400 ;
        RECT 92.400 187.600 93.200 188.400 ;
        RECT 92.500 186.400 93.100 187.600 ;
        RECT 94.100 186.400 94.700 189.600 ;
        RECT 103.700 188.400 104.300 191.600 ;
        RECT 97.200 187.600 98.000 188.400 ;
        RECT 103.600 187.600 104.400 188.400 ;
        RECT 87.600 185.600 88.400 186.400 ;
        RECT 92.400 185.600 93.200 186.400 ;
        RECT 94.000 185.600 94.800 186.400 ;
        RECT 81.200 183.600 82.000 184.400 ;
        RECT 102.000 183.600 102.800 184.400 ;
        RECT 81.300 172.300 81.900 183.600 ;
        RECT 102.100 178.400 102.700 183.600 ;
        RECT 92.400 177.600 93.200 178.400 ;
        RECT 102.000 177.600 102.800 178.400 ;
        RECT 82.800 175.600 83.600 176.400 ;
        RECT 82.900 174.400 83.500 175.600 ;
        RECT 84.400 175.000 85.200 175.800 ;
        RECT 90.600 175.600 91.400 175.800 ;
        RECT 85.800 175.000 91.400 175.600 ;
        RECT 82.800 173.600 83.600 174.400 ;
        RECT 84.400 174.200 85.000 175.000 ;
        RECT 85.800 174.800 86.600 175.000 ;
        RECT 89.200 174.800 90.000 175.000 ;
        RECT 84.400 173.600 90.000 174.200 ;
        RECT 81.300 171.700 83.500 172.300 ;
        RECT 81.200 169.600 82.000 170.400 ;
        RECT 79.600 149.600 80.400 150.400 ;
        RECT 78.000 147.600 78.800 148.400 ;
        RECT 66.800 145.600 67.600 146.400 ;
        RECT 70.000 146.200 70.800 147.000 ;
        RECT 71.400 146.400 75.600 147.000 ;
        RECT 76.600 146.200 77.400 147.000 ;
        RECT 78.100 146.400 78.700 147.600 ;
        RECT 78.000 145.600 78.800 146.400 ;
        RECT 60.400 143.600 61.200 144.400 ;
        RECT 65.200 143.600 66.000 144.400 ;
        RECT 60.500 138.400 61.100 143.600 ;
        RECT 74.800 141.600 75.600 142.400 ;
        RECT 62.000 139.600 62.800 140.400 ;
        RECT 60.400 137.600 61.200 138.400 ;
        RECT 57.200 133.600 58.000 134.400 ;
        RECT 58.800 133.600 59.600 134.400 ;
        RECT 62.100 134.300 62.700 139.600 ;
        RECT 68.400 135.600 69.200 136.400 ;
        RECT 60.500 133.700 62.700 134.300 ;
        RECT 57.300 132.400 57.900 133.600 ;
        RECT 57.200 131.600 58.000 132.400 ;
        RECT 50.800 129.600 51.600 130.400 ;
        RECT 52.400 129.600 53.200 130.400 ;
        RECT 54.000 129.600 54.800 130.400 ;
        RECT 57.200 129.600 58.000 130.400 ;
        RECT 50.900 118.400 51.500 129.600 ;
        RECT 47.600 117.600 48.400 118.400 ;
        RECT 50.800 117.600 51.600 118.400 ;
        RECT 52.400 117.600 53.200 118.400 ;
        RECT 46.000 111.600 46.800 112.400 ;
        RECT 42.800 109.600 43.600 110.400 ;
        RECT 44.400 109.600 45.200 110.400 ;
        RECT 42.900 108.400 43.500 109.600 ;
        RECT 33.200 107.600 34.000 108.400 ;
        RECT 36.400 107.600 37.200 108.400 ;
        RECT 38.000 107.600 38.800 108.400 ;
        RECT 41.200 107.600 42.000 108.400 ;
        RECT 42.800 107.600 43.600 108.400 ;
        RECT 33.200 105.600 34.000 106.400 ;
        RECT 34.800 105.600 35.600 106.400 ;
        RECT 33.300 104.400 33.900 105.600 ;
        RECT 33.200 103.600 34.000 104.400 ;
        RECT 26.800 95.600 27.600 96.400 ;
        RECT 31.600 95.600 32.400 96.400 ;
        RECT 26.900 94.400 27.500 95.600 ;
        RECT 26.800 93.600 27.600 94.400 ;
        RECT 20.400 91.600 21.200 92.400 ;
        RECT 25.200 91.600 26.000 92.400 ;
        RECT 30.000 91.600 30.800 92.400 ;
        RECT 18.800 89.600 19.600 90.400 ;
        RECT 17.200 81.600 18.000 82.400 ;
        RECT 15.600 71.600 16.400 72.400 ;
        RECT 17.200 71.600 18.000 72.400 ;
        RECT 18.900 72.300 19.500 89.600 ;
        RECT 20.500 78.400 21.100 91.600 ;
        RECT 20.400 77.600 21.200 78.400 ;
        RECT 25.300 74.400 25.900 91.600 ;
        RECT 31.700 90.400 32.300 95.600 ;
        RECT 34.800 93.600 35.600 94.400 ;
        RECT 36.500 92.400 37.100 107.600 ;
        RECT 38.100 94.400 38.700 107.600 ;
        RECT 46.100 102.400 46.700 111.600 ;
        RECT 47.700 108.400 48.300 117.600 ;
        RECT 49.200 111.600 50.000 112.400 ;
        RECT 47.600 107.600 48.400 108.400 ;
        RECT 47.700 106.400 48.300 107.600 ;
        RECT 47.600 105.600 48.400 106.400 ;
        RECT 49.300 104.400 49.900 111.600 ;
        RECT 50.800 109.600 51.600 110.400 ;
        RECT 49.200 103.600 50.000 104.400 ;
        RECT 46.000 101.600 46.800 102.400 ;
        RECT 49.300 94.400 49.900 103.600 ;
        RECT 52.500 98.300 53.100 117.600 ;
        RECT 54.100 116.400 54.700 129.600 ;
        RECT 54.000 115.600 54.800 116.400 ;
        RECT 60.500 110.400 61.100 133.700 ;
        RECT 65.200 133.600 66.000 134.400 ;
        RECT 62.000 131.600 62.800 132.400 ;
        RECT 62.100 130.400 62.700 131.600 ;
        RECT 65.300 130.400 65.900 133.600 ;
        RECT 68.500 132.400 69.100 135.600 ;
        RECT 74.900 132.400 75.500 141.600 ;
        RECT 76.400 133.600 77.200 134.400 ;
        RECT 68.400 131.600 69.200 132.400 ;
        RECT 73.200 131.600 74.000 132.400 ;
        RECT 74.800 131.600 75.600 132.400 ;
        RECT 78.000 131.600 78.800 132.400 ;
        RECT 62.000 129.600 62.800 130.400 ;
        RECT 65.200 129.600 66.000 130.400 ;
        RECT 63.600 127.600 64.400 128.400 ;
        RECT 63.700 124.400 64.300 127.600 ;
        RECT 63.600 123.600 64.400 124.400 ;
        RECT 63.700 110.400 64.300 123.600 ;
        RECT 65.300 114.400 65.900 129.600 ;
        RECT 71.600 123.600 72.400 124.400 ;
        RECT 70.000 119.600 70.800 120.400 ;
        RECT 65.200 113.600 66.000 114.400 ;
        RECT 70.100 110.400 70.700 119.600 ;
        RECT 60.400 109.600 61.200 110.400 ;
        RECT 63.600 109.600 64.400 110.400 ;
        RECT 70.000 109.600 70.800 110.400 ;
        RECT 71.700 108.400 72.300 123.600 ;
        RECT 73.300 120.400 73.900 131.600 ;
        RECT 73.200 119.600 74.000 120.400 ;
        RECT 73.200 111.800 74.000 112.600 ;
        RECT 74.900 112.400 75.500 131.600 ;
        RECT 79.700 130.400 80.300 149.600 ;
        RECT 82.900 148.400 83.500 171.700 ;
        RECT 84.400 170.200 85.000 173.600 ;
        RECT 87.600 171.600 88.400 172.400 ;
        RECT 89.400 172.200 90.000 173.600 ;
        RECT 89.400 171.400 90.200 172.200 ;
        RECT 90.800 170.200 91.400 175.000 ;
        RECT 92.500 174.400 93.100 177.600 ;
        RECT 95.800 175.600 96.600 175.800 ;
        RECT 95.800 175.000 101.400 175.600 ;
        RECT 102.000 175.000 102.800 175.800 ;
        RECT 92.400 173.600 93.200 174.400 ;
        RECT 94.000 173.600 94.800 174.400 ;
        RECT 84.400 169.400 85.200 170.200 ;
        RECT 90.600 169.400 91.400 170.200 ;
        RECT 86.000 149.600 86.800 150.400 ;
        RECT 87.600 149.600 88.400 150.400 ;
        RECT 81.200 148.300 82.000 148.400 ;
        RECT 82.800 148.300 83.600 148.400 ;
        RECT 81.200 147.700 83.600 148.300 ;
        RECT 81.200 147.600 82.000 147.700 ;
        RECT 82.800 147.600 83.600 147.700 ;
        RECT 84.400 147.600 85.200 148.400 ;
        RECT 82.800 143.600 83.600 144.400 ;
        RECT 82.900 136.400 83.500 143.600 ;
        RECT 82.800 135.600 83.600 136.400 ;
        RECT 84.500 136.300 85.100 147.600 ;
        RECT 86.100 138.400 86.700 149.600 ;
        RECT 87.700 146.300 88.300 149.600 ;
        RECT 89.200 147.600 90.000 148.400 ;
        RECT 92.400 147.600 93.200 148.400 ;
        RECT 87.700 145.700 89.900 146.300 ;
        RECT 89.300 144.400 89.900 145.700 ;
        RECT 89.200 143.600 90.000 144.400 ;
        RECT 90.800 143.600 91.600 144.400 ;
        RECT 86.000 137.600 86.800 138.400 ;
        RECT 84.500 135.700 86.700 136.300 ;
        RECT 82.800 133.600 83.600 134.400 ;
        RECT 79.600 129.600 80.400 130.400 ;
        RECT 81.200 129.600 82.000 130.400 ;
        RECT 82.900 118.400 83.500 133.600 ;
        RECT 82.800 117.600 83.600 118.400 ;
        RECT 78.000 113.600 78.800 114.400 ;
        RECT 73.200 108.400 73.800 111.800 ;
        RECT 74.800 111.600 75.600 112.400 ;
        RECT 79.800 111.800 80.600 112.600 ;
        RECT 77.200 108.400 78.000 108.600 ;
        RECT 54.000 107.600 54.800 108.400 ;
        RECT 60.400 107.600 61.200 108.400 ;
        RECT 65.200 107.600 66.000 108.400 ;
        RECT 68.400 107.600 69.200 108.400 ;
        RECT 71.600 107.600 72.400 108.400 ;
        RECT 73.200 107.800 78.000 108.400 ;
        RECT 54.100 106.400 54.700 107.600 ;
        RECT 60.500 106.400 61.100 107.600 ;
        RECT 73.200 107.000 73.800 107.800 ;
        RECT 74.600 107.000 75.400 107.200 ;
        RECT 78.000 107.000 78.800 107.200 ;
        RECT 80.000 107.000 80.600 111.800 ;
        RECT 84.400 111.600 85.200 112.400 ;
        RECT 84.500 110.400 85.100 111.600 ;
        RECT 84.400 109.600 85.200 110.400 ;
        RECT 81.200 107.600 82.000 108.400 ;
        RECT 82.800 107.600 83.600 108.400 ;
        RECT 54.000 105.600 54.800 106.400 ;
        RECT 60.400 105.600 61.200 106.400 ;
        RECT 65.200 105.600 66.000 106.400 ;
        RECT 73.200 106.200 74.000 107.000 ;
        RECT 74.600 106.400 78.800 107.000 ;
        RECT 79.800 106.200 80.600 107.000 ;
        RECT 82.900 106.400 83.500 107.600 ;
        RECT 82.800 105.600 83.600 106.400 ;
        RECT 55.600 103.600 56.400 104.400 ;
        RECT 66.800 103.600 67.600 104.400 ;
        RECT 50.900 97.700 53.100 98.300 ;
        RECT 38.000 93.600 38.800 94.400 ;
        RECT 41.200 93.600 42.000 94.400 ;
        RECT 49.200 93.600 50.000 94.400 ;
        RECT 50.900 92.400 51.500 97.700 ;
        RECT 52.400 95.600 53.200 96.400 ;
        RECT 55.700 92.400 56.300 103.600 ;
        RECT 58.800 95.600 59.600 96.400 ;
        RECT 60.400 95.600 61.200 96.400 ;
        RECT 60.500 94.400 61.100 95.600 ;
        RECT 66.900 94.400 67.500 103.600 ;
        RECT 73.200 95.600 74.000 96.400 ;
        RECT 73.300 94.400 73.900 95.600 ;
        RECT 60.400 93.600 61.200 94.400 ;
        RECT 63.600 93.600 64.400 94.400 ;
        RECT 65.200 93.600 66.000 94.400 ;
        RECT 66.800 93.600 67.600 94.400 ;
        RECT 73.200 93.600 74.000 94.400 ;
        RECT 78.000 93.600 78.800 94.400 ;
        RECT 65.300 92.400 65.900 93.600 ;
        RECT 36.400 91.600 37.200 92.400 ;
        RECT 50.800 91.600 51.600 92.400 ;
        RECT 55.600 91.600 56.400 92.400 ;
        RECT 62.000 91.600 62.800 92.400 ;
        RECT 65.200 91.600 66.000 92.400 ;
        RECT 68.400 91.600 69.200 92.400 ;
        RECT 73.200 91.600 74.000 92.400 ;
        RECT 73.300 90.400 73.900 91.600 ;
        RECT 78.100 90.400 78.700 93.600 ;
        RECT 81.200 91.600 82.000 92.400 ;
        RECT 31.600 89.600 32.400 90.400 ;
        RECT 39.600 89.600 40.400 90.400 ;
        RECT 54.000 89.600 54.800 90.400 ;
        RECT 71.600 89.600 72.400 90.400 ;
        RECT 73.200 89.600 74.000 90.400 ;
        RECT 76.400 89.600 77.200 90.400 ;
        RECT 78.000 89.600 78.800 90.400 ;
        RECT 33.200 87.600 34.000 88.400 ;
        RECT 30.000 81.600 30.800 82.400 ;
        RECT 28.400 77.600 29.200 78.400 ;
        RECT 26.800 75.600 27.600 76.400 ;
        RECT 23.600 73.600 24.400 74.400 ;
        RECT 25.200 73.600 26.000 74.400 ;
        RECT 18.900 71.700 21.100 72.300 ;
        RECT 12.400 69.600 13.200 70.400 ;
        RECT 14.000 69.600 14.800 70.400 ;
        RECT 12.500 68.400 13.100 69.600 ;
        RECT 17.300 68.400 17.900 71.600 ;
        RECT 18.800 69.600 19.600 70.400 ;
        RECT 12.400 67.600 13.200 68.400 ;
        RECT 15.600 67.600 16.400 68.400 ;
        RECT 17.200 67.600 18.000 68.400 ;
        RECT 15.700 66.400 16.300 67.600 ;
        RECT 15.600 65.600 16.400 66.400 ;
        RECT 12.400 63.600 13.200 64.400 ;
        RECT 9.200 57.600 10.000 58.400 ;
        RECT 10.800 57.600 11.600 58.400 ;
        RECT 4.400 55.600 5.200 56.400 ;
        RECT 12.500 56.300 13.100 63.600 ;
        RECT 15.700 56.400 16.300 65.600 ;
        RECT 20.500 62.400 21.100 71.700 ;
        RECT 22.000 71.600 22.800 72.400 ;
        RECT 22.100 66.400 22.700 71.600 ;
        RECT 22.000 65.600 22.800 66.400 ;
        RECT 20.400 61.600 21.200 62.400 ;
        RECT 10.900 55.700 13.100 56.300 ;
        RECT 1.200 51.600 2.000 52.400 ;
        RECT 1.300 26.400 1.900 51.600 ;
        RECT 1.200 25.600 2.000 26.400 ;
        RECT 4.500 20.400 5.100 55.600 ;
        RECT 10.900 54.400 11.500 55.700 ;
        RECT 15.600 55.600 16.400 56.400 ;
        RECT 20.500 54.400 21.100 61.600 ;
        RECT 23.700 54.400 24.300 73.600 ;
        RECT 26.900 72.400 27.500 75.600 ;
        RECT 28.500 72.400 29.100 77.600 ;
        RECT 26.800 71.600 27.600 72.400 ;
        RECT 28.400 71.600 29.200 72.400 ;
        RECT 30.100 70.300 30.700 81.600 ;
        RECT 39.700 76.400 40.300 89.600 ;
        RECT 54.100 88.400 54.700 89.600 ;
        RECT 54.000 87.600 54.800 88.400 ;
        RECT 57.200 87.600 58.000 88.400 ;
        RECT 74.800 87.600 75.600 88.400 ;
        RECT 57.300 86.400 57.900 87.600 ;
        RECT 47.600 85.600 48.400 86.400 ;
        RECT 57.200 85.600 58.000 86.400 ;
        RECT 78.100 78.400 78.700 89.600 ;
        RECT 41.200 77.600 42.000 78.400 ;
        RECT 78.000 77.600 78.800 78.400 ;
        RECT 39.600 75.600 40.400 76.400 ;
        RECT 31.600 71.600 32.400 72.400 ;
        RECT 41.300 70.400 41.900 77.600 ;
        RECT 82.900 76.400 83.500 105.600 ;
        RECT 84.500 96.400 85.100 109.600 ;
        RECT 86.100 102.400 86.700 135.700 ;
        RECT 87.600 133.600 88.400 134.400 ;
        RECT 87.700 124.400 88.300 133.600 ;
        RECT 89.300 128.400 89.900 143.600 ;
        RECT 90.900 140.400 91.500 143.600 ;
        RECT 90.800 139.600 91.600 140.400 ;
        RECT 92.500 138.400 93.100 147.600 ;
        RECT 90.800 137.600 91.600 138.400 ;
        RECT 92.400 137.600 93.200 138.400 ;
        RECT 90.900 136.400 91.500 137.600 ;
        RECT 90.800 135.600 91.600 136.400 ;
        RECT 92.400 133.600 93.200 134.400 ;
        RECT 94.100 132.400 94.700 173.600 ;
        RECT 95.800 170.200 96.400 175.000 ;
        RECT 97.200 174.800 98.000 175.000 ;
        RECT 100.600 174.800 101.400 175.000 ;
        RECT 102.200 174.200 102.800 175.000 ;
        RECT 97.200 173.600 102.800 174.200 ;
        RECT 103.600 173.600 104.400 174.400 ;
        RECT 97.200 172.200 97.800 173.600 ;
        RECT 97.000 171.400 97.800 172.200 ;
        RECT 102.200 170.200 102.800 173.600 ;
        RECT 95.800 169.400 96.600 170.200 ;
        RECT 102.000 169.400 102.800 170.200 ;
        RECT 100.400 163.600 101.200 164.400 ;
        RECT 103.700 162.400 104.300 173.600 ;
        RECT 105.200 170.200 106.000 175.800 ;
        RECT 106.900 174.400 107.500 213.600 ;
        RECT 108.500 188.400 109.100 279.600 ;
        RECT 111.700 270.400 112.300 283.600 ;
        RECT 126.000 277.600 126.800 278.400 ;
        RECT 127.600 275.600 128.400 276.400 ;
        RECT 124.400 273.600 125.200 274.400 ;
        RECT 118.000 271.600 118.800 272.400 ;
        RECT 124.500 270.400 125.100 273.600 ;
        RECT 127.700 272.400 128.300 275.600 ;
        RECT 127.600 271.600 128.400 272.400 ;
        RECT 110.000 269.600 110.800 270.400 ;
        RECT 111.600 269.600 112.400 270.400 ;
        RECT 121.200 269.600 122.000 270.400 ;
        RECT 122.800 269.600 123.600 270.400 ;
        RECT 124.400 269.600 125.200 270.400 ;
        RECT 110.100 268.400 110.700 269.600 ;
        RECT 110.000 267.600 110.800 268.400 ;
        RECT 116.400 267.600 117.200 268.400 ;
        RECT 119.600 267.600 120.400 268.400 ;
        RECT 116.500 266.400 117.100 267.600 ;
        RECT 116.400 265.600 117.200 266.400 ;
        RECT 110.000 259.600 110.800 260.400 ;
        RECT 110.100 256.400 110.700 259.600 ;
        RECT 110.000 255.600 110.800 256.400 ;
        RECT 114.800 255.600 115.600 256.400 ;
        RECT 111.600 253.600 112.400 254.400 ;
        RECT 111.700 252.400 112.300 253.600 ;
        RECT 111.600 251.600 112.400 252.400 ;
        RECT 113.200 251.600 114.000 252.400 ;
        RECT 116.500 250.400 117.100 265.600 ;
        RECT 118.000 263.600 118.800 264.400 ;
        RECT 118.100 260.400 118.700 263.600 ;
        RECT 118.000 259.600 118.800 260.400 ;
        RECT 118.000 257.600 118.800 258.400 ;
        RECT 118.100 254.400 118.700 257.600 ;
        RECT 118.000 253.600 118.800 254.400 ;
        RECT 119.700 252.400 120.300 267.600 ;
        RECT 121.300 254.400 121.900 269.600 ;
        RECT 122.900 268.400 123.500 269.600 ;
        RECT 129.300 268.400 129.900 285.600 ;
        RECT 132.500 278.300 133.100 287.600 ;
        RECT 135.600 283.600 136.400 284.400 ;
        RECT 132.500 277.700 134.700 278.300 ;
        RECT 130.800 269.600 131.600 270.400 ;
        RECT 130.900 268.400 131.500 269.600 ;
        RECT 134.100 268.400 134.700 277.700 ;
        RECT 137.200 273.600 138.000 274.400 ;
        RECT 137.300 272.400 137.900 273.600 ;
        RECT 137.200 271.600 138.000 272.400 ;
        RECT 122.800 267.600 123.600 268.400 ;
        RECT 124.400 268.300 125.200 268.400 ;
        RECT 126.000 268.300 126.800 268.400 ;
        RECT 124.400 267.700 126.800 268.300 ;
        RECT 124.400 267.600 125.200 267.700 ;
        RECT 126.000 267.600 126.800 267.700 ;
        RECT 129.200 267.600 130.000 268.400 ;
        RECT 130.800 267.600 131.600 268.400 ;
        RECT 132.400 267.600 133.200 268.400 ;
        RECT 134.000 267.600 134.800 268.400 ;
        RECT 126.100 256.400 126.700 267.600 ;
        RECT 132.500 266.400 133.100 267.600 ;
        RECT 132.400 265.600 133.200 266.400 ;
        RECT 134.100 264.400 134.700 267.600 ;
        RECT 127.600 263.600 128.400 264.400 ;
        RECT 134.000 263.600 134.800 264.400 ;
        RECT 137.200 263.600 138.000 264.400 ;
        RECT 122.800 255.600 123.600 256.400 ;
        RECT 126.000 255.600 126.800 256.400 ;
        RECT 127.700 254.400 128.300 263.600 ;
        RECT 129.000 255.000 129.800 255.800 ;
        RECT 130.800 255.000 135.000 255.600 ;
        RECT 135.600 255.000 136.400 255.800 ;
        RECT 121.200 253.600 122.000 254.400 ;
        RECT 127.600 253.600 128.400 254.400 ;
        RECT 119.600 251.600 120.400 252.400 ;
        RECT 116.400 249.600 117.200 250.400 ;
        RECT 129.000 250.200 129.600 255.000 ;
        RECT 130.800 254.800 131.600 255.000 ;
        RECT 134.200 254.800 135.000 255.000 ;
        RECT 135.800 254.200 136.400 255.000 ;
        RECT 137.300 254.400 137.900 263.600 ;
        RECT 142.100 254.400 142.700 307.600 ;
        RECT 146.900 306.400 147.500 307.600 ;
        RECT 146.800 305.600 147.600 306.400 ;
        RECT 150.000 303.600 150.800 304.400 ;
        RECT 150.100 302.400 150.700 303.600 ;
        RECT 145.200 301.600 146.000 302.400 ;
        RECT 150.000 301.600 150.800 302.400 ;
        RECT 143.600 289.600 144.400 290.400 ;
        RECT 143.700 278.400 144.300 289.600 ;
        RECT 143.600 277.600 144.400 278.400 ;
        RECT 145.300 276.400 145.900 301.600 ;
        RECT 150.000 297.600 150.800 298.400 ;
        RECT 151.600 295.600 152.400 296.400 ;
        RECT 153.300 294.400 153.900 311.600 ;
        RECT 156.500 310.400 157.100 311.700 ;
        RECT 167.600 311.600 168.400 312.400 ;
        RECT 156.400 309.600 157.200 310.400 ;
        RECT 158.000 309.600 158.800 310.400 ;
        RECT 169.200 309.600 170.000 310.400 ;
        RECT 156.500 308.400 157.100 309.600 ;
        RECT 158.100 308.400 158.700 309.600 ;
        RECT 156.400 307.600 157.200 308.400 ;
        RECT 158.000 307.600 158.800 308.400 ;
        RECT 161.200 307.600 162.000 308.400 ;
        RECT 172.500 306.400 173.100 323.600 ;
        RECT 175.600 309.600 176.400 310.400 ;
        RECT 161.200 305.600 162.000 306.400 ;
        RECT 169.200 305.600 170.000 306.400 ;
        RECT 172.400 305.600 173.200 306.400 ;
        RECT 159.600 303.600 160.400 304.400 ;
        RECT 159.700 302.400 160.300 303.600 ;
        RECT 154.800 301.600 155.600 302.400 ;
        RECT 159.600 301.600 160.400 302.400 ;
        RECT 154.900 296.400 155.500 301.600 ;
        RECT 156.400 299.600 157.200 300.400 ;
        RECT 156.500 298.400 157.100 299.600 ;
        RECT 156.400 297.600 157.200 298.400 ;
        RECT 154.800 295.600 155.600 296.400 ;
        RECT 158.000 295.600 158.800 296.400 ;
        RECT 159.600 295.600 160.400 296.400 ;
        RECT 146.800 293.600 147.600 294.400 ;
        RECT 153.200 294.300 154.000 294.400 ;
        RECT 151.700 293.700 154.000 294.300 ;
        RECT 148.400 291.600 149.200 292.400 ;
        RECT 148.500 290.400 149.100 291.600 ;
        RECT 148.400 289.600 149.200 290.400 ;
        RECT 146.800 287.600 147.600 288.400 ;
        RECT 145.200 275.600 146.000 276.400 ;
        RECT 146.900 272.300 147.500 287.600 ;
        RECT 148.400 273.600 149.200 274.400 ;
        RECT 148.500 272.400 149.100 273.600 ;
        RECT 145.300 271.700 147.500 272.300 ;
        RECT 145.300 270.400 145.900 271.700 ;
        RECT 148.400 271.600 149.200 272.400 ;
        RECT 150.000 271.600 150.800 272.400 ;
        RECT 145.200 269.600 146.000 270.400 ;
        RECT 146.800 269.600 147.600 270.400 ;
        RECT 151.700 268.400 152.300 293.700 ;
        RECT 153.200 293.600 154.000 293.700 ;
        RECT 153.200 291.600 154.000 292.400 ;
        RECT 153.300 290.400 153.900 291.600 ;
        RECT 158.100 290.400 158.700 295.600 ;
        RECT 159.700 294.400 160.300 295.600 ;
        RECT 159.600 293.600 160.400 294.400 ;
        RECT 161.300 292.400 161.900 305.600 ;
        RECT 169.300 298.400 169.900 305.600 ;
        RECT 170.800 303.600 171.600 304.400 ;
        RECT 178.800 303.600 179.600 304.400 ;
        RECT 180.400 303.600 181.200 304.400 ;
        RECT 183.600 303.600 184.400 304.400 ;
        RECT 185.200 304.200 186.000 315.800 ;
        RECT 186.900 310.400 187.500 323.600 ;
        RECT 193.200 311.600 194.000 312.400 ;
        RECT 186.800 309.600 187.600 310.400 ;
        RECT 193.300 310.200 193.900 311.600 ;
        RECT 167.600 297.600 168.400 298.400 ;
        RECT 169.200 297.600 170.000 298.400 ;
        RECT 167.700 296.400 168.300 297.600 ;
        RECT 170.900 296.400 171.500 303.600 ;
        RECT 178.900 298.400 179.500 303.600 ;
        RECT 175.600 297.600 176.400 298.400 ;
        RECT 178.800 297.600 179.600 298.400 ;
        RECT 167.600 295.600 168.400 296.400 ;
        RECT 170.800 295.600 171.600 296.400 ;
        RECT 175.700 294.400 176.300 297.600 ;
        RECT 178.800 295.600 179.600 296.400 ;
        RECT 175.600 293.600 176.400 294.400 ;
        RECT 175.700 292.400 176.300 293.600 ;
        RECT 180.500 292.400 181.100 303.600 ;
        RECT 182.000 297.600 182.800 298.400 ;
        RECT 182.100 292.400 182.700 297.600 ;
        RECT 183.700 294.400 184.300 303.600 ;
        RECT 183.600 293.600 184.400 294.400 ;
        RECT 185.200 293.600 186.000 294.400 ;
        RECT 185.300 292.400 185.900 293.600 ;
        RECT 186.900 292.400 187.500 309.600 ;
        RECT 193.200 309.400 194.000 310.200 ;
        RECT 194.800 304.200 195.600 315.800 ;
        RECT 199.600 313.600 200.400 314.400 ;
        RECT 198.000 306.200 198.800 311.800 ;
        RECT 199.700 310.400 200.300 313.600 ;
        RECT 199.600 309.600 200.400 310.400 ;
        RECT 204.400 304.200 205.200 315.800 ;
        RECT 210.900 308.400 211.500 333.600 ;
        RECT 212.400 331.600 213.200 332.600 ;
        RECT 214.000 326.200 214.800 337.800 ;
        RECT 218.800 337.600 219.600 338.400 ;
        RECT 217.200 330.200 218.000 335.800 ;
        RECT 218.900 334.400 219.500 337.600 ;
        RECT 220.400 335.000 221.200 335.800 ;
        RECT 221.800 335.000 226.000 335.600 ;
        RECT 227.000 335.000 227.800 335.800 ;
        RECT 218.800 333.600 219.600 334.400 ;
        RECT 220.400 334.200 221.000 335.000 ;
        RECT 221.800 334.800 222.600 335.000 ;
        RECT 225.200 334.800 226.000 335.000 ;
        RECT 220.400 333.600 225.200 334.200 ;
        RECT 218.800 331.600 219.600 332.400 ;
        RECT 220.400 330.200 221.000 333.600 ;
        RECT 224.400 333.400 225.200 333.600 ;
        RECT 227.200 330.200 227.800 335.000 ;
        RECT 230.100 334.400 230.700 343.700 ;
        RECT 241.200 343.600 242.000 344.400 ;
        RECT 241.300 338.400 241.900 343.600 ;
        RECT 233.200 337.600 234.000 338.400 ;
        RECT 241.200 337.600 242.000 338.400 ;
        RECT 231.600 335.000 232.400 335.800 ;
        RECT 237.800 335.600 238.600 335.800 ;
        RECT 239.600 335.600 240.400 336.400 ;
        RECT 233.000 335.000 238.600 335.600 ;
        RECT 228.400 333.600 229.200 334.400 ;
        RECT 230.000 333.600 230.800 334.400 ;
        RECT 231.600 334.200 232.200 335.000 ;
        RECT 233.000 334.800 233.800 335.000 ;
        RECT 236.400 334.800 237.200 335.000 ;
        RECT 231.600 333.600 237.200 334.200 ;
        RECT 220.400 329.400 221.200 330.200 ;
        RECT 227.000 329.400 227.800 330.200 ;
        RECT 228.500 328.400 229.100 333.600 ;
        RECT 228.400 327.600 229.200 328.400 ;
        RECT 212.400 319.600 213.200 320.400 ;
        RECT 212.500 310.200 213.100 319.600 ;
        RECT 212.400 309.400 213.200 310.200 ;
        RECT 210.800 307.600 211.600 308.400 ;
        RECT 188.200 295.000 189.000 295.800 ;
        RECT 190.000 295.000 194.200 295.600 ;
        RECT 194.800 295.000 195.600 295.800 ;
        RECT 161.200 292.300 162.000 292.400 ;
        RECT 161.200 291.700 163.500 292.300 ;
        RECT 161.200 291.600 162.000 291.700 ;
        RECT 153.200 289.600 154.000 290.400 ;
        RECT 158.000 289.600 158.800 290.400 ;
        RECT 161.200 289.600 162.000 290.400 ;
        RECT 162.900 288.400 163.500 291.700 ;
        RECT 174.000 291.600 174.800 292.400 ;
        RECT 175.600 291.600 176.400 292.400 ;
        RECT 180.400 291.600 181.200 292.400 ;
        RECT 182.000 291.600 182.800 292.400 ;
        RECT 185.200 291.600 186.000 292.400 ;
        RECT 186.800 291.600 187.600 292.400 ;
        RECT 162.800 287.600 163.600 288.400 ;
        RECT 174.100 284.400 174.700 291.600 ;
        RECT 185.200 289.600 186.000 290.400 ;
        RECT 185.300 288.400 185.900 289.600 ;
        RECT 185.200 287.600 186.000 288.400 ;
        RECT 156.400 283.600 157.200 284.400 ;
        RECT 169.200 283.600 170.000 284.400 ;
        RECT 174.000 283.600 174.800 284.400 ;
        RECT 175.600 283.600 176.400 284.400 ;
        RECT 153.200 271.600 154.000 272.400 ;
        RECT 153.300 268.400 153.900 271.600 ;
        RECT 151.600 267.600 152.400 268.400 ;
        RECT 153.200 267.600 154.000 268.400 ;
        RECT 154.800 267.600 155.600 268.400 ;
        RECT 154.900 266.400 155.500 267.600 ;
        RECT 154.800 265.600 155.600 266.400 ;
        RECT 145.000 255.000 145.800 255.800 ;
        RECT 146.800 255.000 151.000 255.600 ;
        RECT 151.600 255.000 152.400 255.800 ;
        RECT 131.600 253.600 136.400 254.200 ;
        RECT 137.200 253.600 138.000 254.400 ;
        RECT 142.000 253.600 142.800 254.400 ;
        RECT 131.600 253.400 132.400 253.600 ;
        RECT 135.800 250.200 136.400 253.600 ;
        RECT 129.000 249.400 129.800 250.200 ;
        RECT 135.600 249.400 136.400 250.200 ;
        RECT 145.000 250.200 145.600 255.000 ;
        RECT 146.800 254.800 147.600 255.000 ;
        RECT 150.200 254.800 151.000 255.000 ;
        RECT 151.800 254.200 152.400 255.000 ;
        RECT 156.500 254.400 157.100 283.600 ;
        RECT 169.300 274.400 169.900 283.600 ;
        RECT 169.200 273.600 170.000 274.400 ;
        RECT 166.000 271.600 166.800 272.400 ;
        RECT 172.400 271.600 173.200 272.400 ;
        RECT 158.000 269.600 158.800 270.400 ;
        RECT 161.200 269.600 162.000 270.400 ;
        RECT 162.800 269.600 163.600 270.400 ;
        RECT 166.100 268.400 166.700 271.600 ;
        RECT 169.200 269.600 170.000 270.400 ;
        RECT 159.600 267.600 160.400 268.400 ;
        RECT 166.000 267.600 166.800 268.400 ;
        RECT 167.600 267.600 168.400 268.400 ;
        RECT 159.700 266.400 160.300 267.600 ;
        RECT 158.000 265.600 158.800 266.400 ;
        RECT 159.600 265.600 160.400 266.400 ;
        RECT 164.400 265.600 165.200 266.400 ;
        RECT 158.100 258.400 158.700 265.600 ;
        RECT 158.000 257.600 158.800 258.400 ;
        RECT 147.600 253.600 152.400 254.200 ;
        RECT 153.200 253.600 154.000 254.400 ;
        RECT 154.800 253.600 155.600 254.400 ;
        RECT 156.400 253.600 157.200 254.400 ;
        RECT 159.600 253.600 160.400 254.400 ;
        RECT 147.600 253.400 148.400 253.600 ;
        RECT 150.000 251.600 150.800 252.400 ;
        RECT 145.000 249.400 145.800 250.200 ;
        RECT 130.800 243.600 131.600 244.400 ;
        RECT 146.800 243.600 147.600 244.400 ;
        RECT 130.900 238.400 131.500 243.600 ;
        RECT 110.000 237.600 110.800 238.400 ;
        RECT 130.800 237.600 131.600 238.400 ;
        RECT 110.100 230.200 110.700 237.600 ;
        RECT 110.000 229.400 110.800 230.200 ;
        RECT 111.600 224.200 112.400 235.800 ;
        RECT 114.800 226.200 115.600 231.800 ;
        RECT 116.400 223.600 117.200 224.400 ;
        RECT 121.200 224.200 122.000 235.800 ;
        RECT 129.200 233.600 130.000 234.400 ;
        RECT 129.300 230.200 129.900 233.600 ;
        RECT 129.200 229.400 130.000 230.200 ;
        RECT 130.800 224.200 131.600 235.800 ;
        RECT 132.400 227.600 133.200 228.400 ;
        RECT 116.500 222.400 117.100 223.600 ;
        RECT 116.400 221.600 117.200 222.400 ;
        RECT 116.400 206.200 117.200 217.800 ;
        RECT 118.000 213.600 118.800 214.400 ;
        RECT 118.100 212.400 118.700 213.600 ;
        RECT 118.000 211.600 118.800 212.400 ;
        RECT 124.400 211.600 125.200 212.600 ;
        RECT 126.000 206.200 126.800 217.800 ;
        RECT 127.600 213.600 128.400 214.400 ;
        RECT 111.600 203.600 112.400 204.400 ;
        RECT 121.200 195.600 122.000 196.400 ;
        RECT 110.000 191.600 110.800 192.400 ;
        RECT 121.300 188.400 121.900 195.600 ;
        RECT 108.400 187.600 109.200 188.400 ;
        RECT 113.200 187.600 114.000 188.400 ;
        RECT 121.200 187.600 122.000 188.400 ;
        RECT 111.600 183.600 112.400 184.400 ;
        RECT 119.600 183.600 120.400 184.400 ;
        RECT 106.800 173.600 107.600 174.400 ;
        RECT 108.400 166.200 109.200 177.800 ;
        RECT 111.700 174.400 112.300 183.600 ;
        RECT 111.600 173.600 112.400 174.400 ;
        RECT 110.000 171.600 110.800 172.600 ;
        RECT 118.000 166.200 118.800 177.800 ;
        RECT 119.700 170.400 120.300 183.600 ;
        RECT 119.600 169.600 120.400 170.400 ;
        RECT 110.000 163.600 110.800 164.400 ;
        RECT 103.600 161.600 104.400 162.400 ;
        RECT 108.400 155.600 109.200 156.400 ;
        RECT 103.600 153.600 104.400 154.400 ;
        RECT 106.800 153.600 107.600 154.400 ;
        RECT 103.700 152.400 104.300 153.600 ;
        RECT 103.600 151.600 104.400 152.400 ;
        RECT 97.200 149.600 98.000 150.400 ;
        RECT 98.800 149.600 99.600 150.400 ;
        RECT 106.800 149.600 107.600 150.400 ;
        RECT 98.900 146.400 99.500 149.600 ;
        RECT 106.900 148.400 107.500 149.600 ;
        RECT 106.800 147.600 107.600 148.400 ;
        RECT 97.200 145.600 98.000 146.400 ;
        RECT 98.800 145.600 99.600 146.400 ;
        RECT 103.600 145.600 104.400 146.400 ;
        RECT 103.700 144.400 104.300 145.600 ;
        RECT 103.600 143.600 104.400 144.400 ;
        RECT 103.700 134.400 104.300 143.600 ;
        RECT 108.500 134.400 109.100 155.600 ;
        RECT 110.100 154.400 110.700 163.600 ;
        RECT 111.600 161.600 112.400 162.400 ;
        RECT 110.000 153.600 110.800 154.400 ;
        RECT 110.100 146.400 110.700 153.600 ;
        RECT 111.700 148.400 112.300 161.600 ;
        RECT 113.200 151.800 114.000 152.600 ;
        RECT 119.800 151.800 120.600 152.600 ;
        RECT 113.200 148.400 113.800 151.800 ;
        RECT 114.800 149.600 115.600 150.400 ;
        RECT 117.200 148.400 118.000 148.600 ;
        RECT 111.600 147.600 112.400 148.400 ;
        RECT 113.200 147.800 118.000 148.400 ;
        RECT 110.000 145.600 110.800 146.400 ;
        RECT 110.000 135.600 110.800 136.400 ;
        RECT 103.600 133.600 104.400 134.400 ;
        RECT 108.400 133.600 109.200 134.400 ;
        RECT 108.500 132.400 109.100 133.600 ;
        RECT 94.000 131.600 94.800 132.400 ;
        RECT 108.400 131.600 109.200 132.400 ;
        RECT 111.700 130.400 112.300 147.600 ;
        RECT 113.200 147.000 113.800 147.800 ;
        RECT 114.600 147.000 115.400 147.200 ;
        RECT 118.000 147.000 118.800 147.200 ;
        RECT 120.000 147.000 120.600 151.800 ;
        RECT 121.300 148.400 121.900 187.600 ;
        RECT 122.800 186.200 123.600 191.800 ;
        RECT 126.000 184.200 126.800 195.800 ;
        RECT 127.700 188.400 128.300 213.600 ;
        RECT 129.200 210.200 130.000 215.800 ;
        RECT 132.500 214.400 133.100 227.600 ;
        RECT 134.000 226.200 134.800 231.800 ;
        RECT 140.400 231.600 141.200 232.400 ;
        RECT 141.800 231.800 142.600 232.600 ;
        RECT 148.400 231.800 149.200 232.600 ;
        RECT 140.500 228.400 141.100 231.600 ;
        RECT 140.400 227.600 141.200 228.400 ;
        RECT 141.800 227.000 142.400 231.800 ;
        RECT 144.400 228.400 145.200 228.600 ;
        RECT 148.600 228.400 149.200 231.800 ;
        RECT 150.100 228.400 150.700 251.600 ;
        RECT 151.800 250.200 152.400 253.600 ;
        RECT 154.900 252.400 155.500 253.600 ;
        RECT 154.800 251.600 155.600 252.400 ;
        RECT 151.600 249.400 152.400 250.200 ;
        RECT 159.700 248.400 160.300 253.600 ;
        RECT 161.200 251.600 162.000 252.400 ;
        RECT 162.800 251.600 163.600 252.400 ;
        RECT 161.300 250.400 161.900 251.600 ;
        RECT 161.200 249.600 162.000 250.400 ;
        RECT 159.600 248.300 160.400 248.400 ;
        RECT 158.100 247.700 160.400 248.300 ;
        RECT 151.600 241.600 152.400 242.400 ;
        RECT 151.700 228.400 152.300 241.600 ;
        RECT 153.200 231.600 154.000 232.400 ;
        RECT 158.100 230.400 158.700 247.700 ;
        RECT 159.600 247.600 160.400 247.700 ;
        RECT 162.900 232.400 163.500 251.600 ;
        RECT 164.500 250.400 165.100 265.600 ;
        RECT 167.700 260.400 168.300 267.600 ;
        RECT 175.700 264.400 176.300 283.600 ;
        RECT 178.800 273.600 179.600 274.400 ;
        RECT 178.900 272.400 179.500 273.600 ;
        RECT 178.800 271.600 179.600 272.400 ;
        RECT 177.200 267.600 178.000 268.400 ;
        RECT 174.000 263.600 174.800 264.400 ;
        RECT 175.600 263.600 176.400 264.400 ;
        RECT 182.000 263.600 182.800 264.400 ;
        RECT 183.600 264.200 184.400 275.800 ;
        RECT 186.900 270.400 187.500 291.600 ;
        RECT 188.200 290.200 188.800 295.000 ;
        RECT 190.000 294.800 190.800 295.000 ;
        RECT 193.400 294.800 194.200 295.000 ;
        RECT 195.000 294.200 195.600 295.000 ;
        RECT 190.800 293.600 195.600 294.200 ;
        RECT 190.800 293.400 191.600 293.600 ;
        RECT 195.000 290.200 195.600 293.600 ;
        RECT 188.200 289.400 189.000 290.200 ;
        RECT 194.800 289.400 195.600 290.200 ;
        RECT 190.000 287.600 190.800 288.400 ;
        RECT 198.000 285.600 198.800 286.400 ;
        RECT 202.800 286.200 203.600 297.800 ;
        RECT 210.900 296.400 211.500 307.600 ;
        RECT 214.000 304.200 214.800 315.800 ;
        RECT 228.400 315.600 229.200 316.400 ;
        RECT 228.500 312.400 229.100 315.600 ;
        RECT 217.200 306.200 218.000 311.800 ;
        RECT 228.400 311.600 229.200 312.400 ;
        RECT 228.400 310.300 229.200 310.400 ;
        RECT 230.100 310.300 230.700 333.600 ;
        RECT 231.600 330.200 232.200 333.600 ;
        RECT 234.800 331.600 235.600 332.400 ;
        RECT 236.600 332.200 237.200 333.600 ;
        RECT 236.600 331.400 237.400 332.200 ;
        RECT 238.000 330.200 238.600 335.000 ;
        RECT 239.700 334.400 240.300 335.600 ;
        RECT 239.600 333.600 240.400 334.400 ;
        RECT 241.300 330.400 241.900 337.600 ;
        RECT 242.900 336.400 243.500 347.600 ;
        RECT 247.700 346.400 248.300 349.600 ;
        RECT 249.300 348.400 249.900 349.600 ;
        RECT 249.200 347.600 250.000 348.400 ;
        RECT 254.000 347.600 254.800 348.400 ;
        RECT 244.400 345.600 245.200 346.400 ;
        RECT 247.600 345.600 248.400 346.400 ;
        RECT 242.800 335.600 243.600 336.400 ;
        RECT 244.500 334.400 245.100 345.600 ;
        RECT 249.300 344.400 249.900 347.600 ;
        RECT 247.600 343.600 248.400 344.400 ;
        RECT 249.200 343.600 250.000 344.400 ;
        RECT 246.000 335.600 246.800 336.400 ;
        RECT 246.100 334.400 246.700 335.600 ;
        RECT 244.400 333.600 245.200 334.400 ;
        RECT 246.000 333.600 246.800 334.400 ;
        RECT 244.500 332.400 245.100 333.600 ;
        RECT 244.400 331.600 245.200 332.400 ;
        RECT 231.600 329.400 232.400 330.200 ;
        RECT 237.800 329.400 238.600 330.200 ;
        RECT 239.600 329.600 240.400 330.400 ;
        RECT 241.200 329.600 242.000 330.400 ;
        RECT 234.800 317.600 235.600 318.400 ;
        RECT 234.900 312.400 235.500 317.600 ;
        RECT 231.600 311.600 232.400 312.400 ;
        RECT 234.800 311.600 235.600 312.400 ;
        RECT 228.400 309.700 230.700 310.300 ;
        RECT 228.400 309.600 229.200 309.700 ;
        RECT 230.100 308.400 230.700 309.700 ;
        RECT 231.600 309.600 232.400 310.400 ;
        RECT 230.000 307.600 230.800 308.400 ;
        RECT 210.800 295.600 211.600 296.400 ;
        RECT 204.400 291.600 205.200 292.400 ;
        RECT 210.800 291.600 211.600 292.600 ;
        RECT 212.400 286.200 213.200 297.800 ;
        RECT 215.600 290.200 216.400 295.800 ;
        RECT 226.800 290.200 227.600 295.800 ;
        RECT 230.000 286.200 230.800 297.800 ;
        RECT 231.600 293.600 232.400 294.400 ;
        RECT 228.400 283.600 229.200 284.400 ;
        RECT 191.600 273.600 192.400 274.400 ;
        RECT 186.800 269.600 187.600 270.400 ;
        RECT 191.700 270.200 192.300 273.600 ;
        RECT 191.600 269.400 192.400 270.200 ;
        RECT 185.200 267.600 186.000 268.400 ;
        RECT 167.600 259.600 168.400 260.400 ;
        RECT 170.800 259.600 171.600 260.400 ;
        RECT 170.900 258.400 171.500 259.600 ;
        RECT 169.200 257.600 170.000 258.400 ;
        RECT 170.800 257.600 171.600 258.400 ;
        RECT 169.300 254.400 169.900 257.600 ;
        RECT 169.200 253.600 170.000 254.400 ;
        RECT 169.300 252.400 169.900 253.600 ;
        RECT 169.200 251.600 170.000 252.400 ;
        RECT 164.400 249.600 165.200 250.400 ;
        RECT 162.800 231.600 163.600 232.400 ;
        RECT 153.200 229.600 154.000 230.400 ;
        RECT 158.000 229.600 158.800 230.400 ;
        RECT 159.600 229.600 160.400 230.400 ;
        RECT 158.100 228.400 158.700 229.600 ;
        RECT 144.400 227.800 149.200 228.400 ;
        RECT 143.600 227.000 144.400 227.200 ;
        RECT 147.000 227.000 147.800 227.200 ;
        RECT 148.600 227.000 149.200 227.800 ;
        RECT 150.000 227.600 150.800 228.400 ;
        RECT 151.600 227.600 152.400 228.400 ;
        RECT 158.000 227.600 158.800 228.400 ;
        RECT 141.800 226.200 142.600 227.000 ;
        RECT 143.600 226.400 147.800 227.000 ;
        RECT 148.400 226.200 149.200 227.000 ;
        RECT 143.600 223.600 144.400 224.400 ;
        RECT 162.800 223.600 163.600 224.400 ;
        RECT 164.400 223.600 165.200 224.400 ;
        RECT 169.200 224.200 170.000 235.800 ;
        RECT 170.800 227.600 171.600 228.400 ;
        RECT 132.400 213.600 133.200 214.400 ;
        RECT 135.600 210.200 136.400 215.800 ;
        RECT 138.800 206.200 139.600 217.800 ;
        RECT 143.700 212.400 144.300 223.600 ;
        RECT 143.600 211.600 144.400 212.400 ;
        RECT 146.800 211.600 147.600 212.400 ;
        RECT 148.400 206.200 149.200 217.800 ;
        RECT 154.800 210.200 155.600 215.800 ;
        RECT 156.400 211.600 157.200 212.400 ;
        RECT 153.200 203.600 154.000 204.400 ;
        RECT 129.200 189.600 130.000 190.400 ;
        RECT 127.600 187.600 128.400 188.400 ;
        RECT 135.600 184.200 136.400 195.800 ;
        RECT 146.800 186.200 147.600 191.800 ;
        RECT 145.200 183.600 146.000 184.400 ;
        RECT 150.000 184.200 150.800 195.800 ;
        RECT 151.600 189.400 152.400 190.400 ;
        RECT 153.300 182.400 153.900 203.600 ;
        RECT 156.500 190.400 157.100 211.600 ;
        RECT 158.000 206.200 158.800 217.800 ;
        RECT 162.900 212.400 163.500 223.600 ;
        RECT 164.500 216.400 165.100 223.600 ;
        RECT 164.400 215.600 165.200 216.400 ;
        RECT 162.800 211.600 163.600 212.400 ;
        RECT 166.000 211.600 166.800 212.400 ;
        RECT 167.600 206.200 168.400 217.800 ;
        RECT 170.900 212.400 171.500 227.600 ;
        RECT 174.100 218.300 174.700 263.600 ;
        RECT 180.400 255.600 181.200 256.400 ;
        RECT 182.100 254.400 182.700 263.600 ;
        RECT 175.600 253.600 176.400 254.400 ;
        RECT 182.000 253.600 182.800 254.400 ;
        RECT 175.600 251.600 176.400 252.400 ;
        RECT 177.200 251.600 178.000 252.400 ;
        RECT 178.800 251.600 179.600 252.400 ;
        RECT 175.700 248.400 176.300 251.600 ;
        RECT 177.200 249.600 178.000 250.400 ;
        RECT 177.300 248.400 177.900 249.600 ;
        RECT 175.600 247.600 176.400 248.400 ;
        RECT 177.200 247.600 178.000 248.400 ;
        RECT 178.900 238.300 179.500 251.600 ;
        RECT 182.100 250.400 182.700 253.600 ;
        RECT 182.000 249.600 182.800 250.400 ;
        RECT 180.400 245.600 181.200 246.400 ;
        RECT 177.300 237.700 179.500 238.300 ;
        RECT 177.300 230.200 177.900 237.700 ;
        RECT 177.200 229.400 178.000 230.200 ;
        RECT 178.800 224.200 179.600 235.800 ;
        RECT 180.500 228.400 181.100 245.600 ;
        RECT 182.100 242.400 182.700 249.600 ;
        RECT 185.300 246.400 185.900 267.600 ;
        RECT 193.200 264.200 194.000 275.800 ;
        RECT 196.400 266.200 197.200 271.800 ;
        RECT 198.000 263.600 198.800 264.400 ;
        RECT 202.800 264.200 203.600 275.800 ;
        RECT 206.000 269.600 206.800 270.400 ;
        RECT 190.000 259.600 190.800 260.400 ;
        RECT 198.000 259.600 198.800 260.400 ;
        RECT 190.100 256.400 190.700 259.600 ;
        RECT 198.100 256.400 198.700 259.600 ;
        RECT 199.600 257.600 200.400 258.400 ;
        RECT 199.700 256.400 200.300 257.600 ;
        RECT 186.800 255.600 187.600 256.400 ;
        RECT 190.000 255.600 190.800 256.400 ;
        RECT 193.200 255.600 194.000 256.400 ;
        RECT 198.000 255.600 198.800 256.400 ;
        RECT 199.600 255.600 200.400 256.400 ;
        RECT 186.900 254.400 187.500 255.600 ;
        RECT 186.800 253.600 187.600 254.400 ;
        RECT 193.300 252.400 193.900 255.600 ;
        RECT 186.800 251.600 187.600 252.400 ;
        RECT 190.000 251.600 190.800 252.400 ;
        RECT 193.200 251.600 194.000 252.400 ;
        RECT 193.200 247.600 194.000 248.400 ;
        RECT 185.200 245.600 186.000 246.400 ;
        RECT 204.400 246.200 205.200 257.800 ;
        RECT 206.100 252.400 206.700 269.600 ;
        RECT 210.800 269.400 211.600 270.400 ;
        RECT 212.400 264.200 213.200 275.800 ;
        RECT 220.400 273.600 221.200 274.400 ;
        RECT 215.600 266.200 216.400 271.800 ;
        RECT 217.200 271.600 218.000 272.400 ;
        RECT 218.600 271.800 219.400 272.600 ;
        RECT 225.200 271.800 226.000 272.600 ;
        RECT 217.300 268.400 217.900 271.600 ;
        RECT 217.200 267.600 218.000 268.400 ;
        RECT 218.600 267.000 219.200 271.800 ;
        RECT 221.200 268.400 222.000 268.600 ;
        RECT 225.400 268.400 226.000 271.800 ;
        RECT 228.500 270.400 229.100 283.600 ;
        RECT 228.400 269.600 229.200 270.400 ;
        RECT 221.200 267.800 226.000 268.400 ;
        RECT 220.400 267.000 221.200 267.200 ;
        RECT 223.800 267.000 224.600 267.200 ;
        RECT 225.400 267.000 226.000 267.800 ;
        RECT 230.000 267.600 230.800 268.400 ;
        RECT 218.600 266.200 219.400 267.000 ;
        RECT 220.400 266.400 224.600 267.000 ;
        RECT 225.200 266.200 226.000 267.000 ;
        RECT 215.600 263.600 216.400 264.400 ;
        RECT 206.000 251.600 206.800 252.400 ;
        RECT 212.400 251.600 213.200 252.600 ;
        RECT 185.200 243.600 186.000 244.400 ;
        RECT 182.000 241.600 182.800 242.400 ;
        RECT 180.400 227.600 181.200 228.400 ;
        RECT 180.500 218.400 181.100 227.600 ;
        RECT 182.000 226.200 182.800 231.800 ;
        RECT 185.300 230.400 185.900 243.600 ;
        RECT 185.200 229.600 186.000 230.400 ;
        RECT 196.400 229.600 197.200 230.400 ;
        RECT 191.600 223.600 192.400 224.400 ;
        RECT 198.000 223.600 198.800 224.400 ;
        RECT 202.800 224.200 203.600 235.800 ;
        RECT 204.400 230.300 205.200 230.400 ;
        RECT 206.100 230.300 206.700 251.600 ;
        RECT 214.000 246.200 214.800 257.800 ;
        RECT 215.700 252.400 216.300 263.600 ;
        RECT 218.800 257.600 219.600 258.400 ;
        RECT 215.600 251.600 216.400 252.400 ;
        RECT 217.200 250.200 218.000 255.800 ;
        RECT 223.600 246.200 224.400 257.800 ;
        RECT 231.700 256.400 232.300 293.600 ;
        RECT 233.200 269.600 234.000 270.400 ;
        RECT 234.900 266.400 235.500 311.600 ;
        RECT 239.700 310.400 240.300 329.600 ;
        RECT 244.400 323.600 245.200 324.400 ;
        RECT 244.500 314.400 245.100 323.600 ;
        RECT 241.200 313.600 242.000 314.400 ;
        RECT 244.400 313.600 245.200 314.400 ;
        RECT 239.600 309.600 240.400 310.400 ;
        RECT 239.600 307.600 240.400 308.400 ;
        RECT 241.300 306.400 241.900 313.600 ;
        RECT 244.400 311.600 245.200 312.400 ;
        RECT 242.800 309.600 243.600 310.400 ;
        RECT 244.500 308.400 245.100 311.600 ;
        RECT 246.100 310.400 246.700 333.600 ;
        RECT 247.700 330.400 248.300 343.600 ;
        RECT 254.100 338.400 254.700 347.600 ;
        RECT 255.700 346.400 256.300 351.600 ;
        RECT 263.700 348.400 264.300 365.700 ;
        RECT 266.800 363.600 267.600 364.400 ;
        RECT 266.900 354.400 267.500 363.600 ;
        RECT 268.400 355.600 269.200 356.400 ;
        RECT 266.800 353.600 267.600 354.400 ;
        RECT 276.400 353.600 277.200 354.400 ;
        RECT 266.600 351.800 267.400 352.600 ;
        RECT 273.200 351.800 274.000 352.600 ;
        RECT 265.200 349.600 266.000 350.400 ;
        RECT 265.300 348.400 265.900 349.600 ;
        RECT 263.600 347.600 264.400 348.400 ;
        RECT 265.200 347.600 266.000 348.400 ;
        RECT 255.600 345.600 256.400 346.400 ;
        RECT 250.800 338.300 251.600 338.400 ;
        RECT 250.800 337.700 253.100 338.300 ;
        RECT 250.800 337.600 251.600 337.700 ;
        RECT 250.900 334.400 251.500 337.600 ;
        RECT 250.800 333.600 251.600 334.400 ;
        RECT 252.500 332.400 253.100 337.700 ;
        RECT 254.000 337.600 254.800 338.400 ;
        RECT 254.100 336.400 254.700 337.600 ;
        RECT 254.000 335.600 254.800 336.400 ;
        RECT 250.800 331.600 251.600 332.400 ;
        RECT 252.400 331.600 253.200 332.400 ;
        RECT 254.000 331.600 254.800 332.400 ;
        RECT 250.900 330.400 251.500 331.600 ;
        RECT 247.600 329.600 248.400 330.400 ;
        RECT 250.800 329.600 251.600 330.400 ;
        RECT 247.700 312.400 248.300 329.600 ;
        RECT 254.100 328.400 254.700 331.600 ;
        RECT 255.700 330.400 256.300 345.600 ;
        RECT 262.000 343.600 262.800 344.400 ;
        RECT 262.100 342.400 262.700 343.600 ;
        RECT 262.000 341.600 262.800 342.400 ;
        RECT 262.000 339.600 262.800 340.400 ;
        RECT 262.100 334.400 262.700 339.600 ;
        RECT 263.700 336.400 264.300 347.600 ;
        RECT 266.600 347.000 267.200 351.800 ;
        RECT 269.200 348.400 270.000 348.600 ;
        RECT 273.400 348.400 274.000 351.800 ;
        RECT 276.500 350.400 277.100 353.600 ;
        RECT 278.000 351.600 278.800 352.400 ;
        RECT 281.300 352.300 281.900 383.600 ;
        RECT 282.900 374.400 283.500 387.600 ;
        RECT 284.200 387.000 284.800 391.800 ;
        RECT 286.800 388.400 287.600 388.600 ;
        RECT 291.000 388.400 291.600 391.800 ;
        RECT 308.400 391.600 309.200 392.400 ;
        RECT 311.600 391.600 312.400 392.400 ;
        RECT 313.200 391.600 314.000 392.400 ;
        RECT 311.700 390.400 312.300 391.600 ;
        RECT 316.500 390.400 317.100 397.600 ;
        RECT 292.400 389.600 293.200 390.400 ;
        RECT 302.000 389.600 302.800 390.400 ;
        RECT 311.600 389.600 312.400 390.400 ;
        RECT 316.400 389.600 317.200 390.400 ;
        RECT 292.500 388.400 293.100 389.600 ;
        RECT 286.800 387.800 291.600 388.400 ;
        RECT 286.000 387.000 286.800 387.200 ;
        RECT 289.400 387.000 290.200 387.200 ;
        RECT 291.000 387.000 291.600 387.800 ;
        RECT 292.400 387.600 293.200 388.400 ;
        RECT 298.800 387.600 299.600 388.400 ;
        RECT 284.200 386.200 285.000 387.000 ;
        RECT 286.000 386.400 290.200 387.000 ;
        RECT 290.800 386.200 291.600 387.000 ;
        RECT 298.900 386.400 299.500 387.600 ;
        RECT 302.100 386.400 302.700 389.600 ;
        RECT 318.100 388.400 318.700 403.700 ;
        RECT 303.600 387.600 304.400 388.400 ;
        RECT 311.600 387.600 312.400 388.400 ;
        RECT 318.000 387.600 318.800 388.400 ;
        RECT 298.800 385.600 299.600 386.400 ;
        RECT 302.000 385.600 302.800 386.400 ;
        RECT 286.000 383.600 286.800 384.400 ;
        RECT 287.600 383.600 288.400 384.400 ;
        RECT 282.800 373.600 283.600 374.400 ;
        RECT 286.100 370.400 286.700 383.600 ;
        RECT 287.600 381.600 288.400 382.400 ;
        RECT 287.700 378.400 288.300 381.600 ;
        RECT 287.600 377.600 288.400 378.400 ;
        RECT 287.600 375.600 288.400 376.400 ;
        RECT 289.200 373.600 290.000 374.400 ;
        RECT 289.200 371.600 290.000 372.400 ;
        RECT 286.000 369.600 286.800 370.400 ;
        RECT 282.800 352.300 283.600 352.400 ;
        RECT 281.300 351.700 283.600 352.300 ;
        RECT 282.800 351.600 283.600 351.700 ;
        RECT 274.800 349.600 275.600 350.400 ;
        RECT 276.400 349.600 277.200 350.400 ;
        RECT 274.900 348.400 275.500 349.600 ;
        RECT 269.200 347.800 274.000 348.400 ;
        RECT 268.400 347.000 269.200 347.200 ;
        RECT 271.800 347.000 272.600 347.200 ;
        RECT 273.400 347.000 274.000 347.800 ;
        RECT 274.800 347.600 275.600 348.400 ;
        RECT 276.400 347.600 277.200 348.400 ;
        RECT 266.600 346.200 267.400 347.000 ;
        RECT 268.400 346.400 272.600 347.000 ;
        RECT 273.200 346.200 274.000 347.000 ;
        RECT 274.800 345.600 275.600 346.400 ;
        RECT 271.600 341.600 272.400 342.400 ;
        RECT 266.800 339.600 267.600 340.400 ;
        RECT 266.900 338.400 267.500 339.600 ;
        RECT 266.800 337.600 267.600 338.400 ;
        RECT 270.000 337.600 270.800 338.400 ;
        RECT 270.100 336.400 270.700 337.600 ;
        RECT 263.600 335.600 264.400 336.400 ;
        RECT 268.400 335.600 269.200 336.400 ;
        RECT 270.000 335.600 270.800 336.400 ;
        RECT 262.000 333.600 262.800 334.400 ;
        RECT 265.200 333.600 266.000 334.400 ;
        RECT 263.600 331.600 264.400 332.400 ;
        RECT 255.600 329.600 256.400 330.400 ;
        RECT 266.800 329.600 267.600 330.400 ;
        RECT 254.000 327.600 254.800 328.400 ;
        RECT 255.600 327.600 256.400 328.400 ;
        RECT 249.200 313.600 250.000 314.400 ;
        RECT 247.600 311.600 248.400 312.400 ;
        RECT 246.000 309.600 246.800 310.400 ;
        RECT 244.400 307.600 245.200 308.400 ;
        RECT 241.200 305.600 242.000 306.400 ;
        RECT 244.400 298.300 245.200 298.400 ;
        RECT 246.100 298.300 246.700 309.600 ;
        RECT 249.300 306.400 249.900 313.600 ;
        RECT 250.800 309.600 251.600 310.400 ;
        RECT 252.400 309.600 253.200 310.400 ;
        RECT 250.900 308.400 251.500 309.600 ;
        RECT 252.500 308.400 253.100 309.600 ;
        RECT 250.800 307.600 251.600 308.400 ;
        RECT 252.400 307.600 253.200 308.400 ;
        RECT 249.200 305.600 250.000 306.400 ;
        RECT 254.100 298.400 254.700 327.600 ;
        RECT 255.700 326.400 256.300 327.600 ;
        RECT 255.600 325.600 256.400 326.400 ;
        RECT 255.700 312.400 256.300 325.600 ;
        RECT 260.400 323.600 261.200 324.400 ;
        RECT 260.500 316.400 261.100 323.600 ;
        RECT 260.400 315.600 261.200 316.400 ;
        RECT 263.600 313.600 264.400 314.400 ;
        RECT 255.600 311.600 256.400 312.400 ;
        RECT 263.700 310.400 264.300 313.600 ;
        RECT 266.900 310.400 267.500 329.600 ;
        RECT 268.500 318.400 269.100 335.600 ;
        RECT 268.400 317.600 269.200 318.400 ;
        RECT 271.700 312.400 272.300 341.600 ;
        RECT 273.200 335.600 274.000 336.400 ;
        RECT 274.900 334.400 275.500 345.600 ;
        RECT 276.500 334.400 277.100 347.600 ;
        RECT 282.900 338.400 283.500 351.600 ;
        RECT 286.100 348.400 286.700 369.600 ;
        RECT 289.300 358.400 289.900 371.600 ;
        RECT 289.200 357.600 290.000 358.400 ;
        RECT 292.400 353.600 293.200 354.400 ;
        RECT 292.500 350.400 293.100 353.600 ;
        RECT 294.000 351.600 294.800 352.400 ;
        RECT 294.100 350.400 294.700 351.600 ;
        RECT 298.900 350.400 299.500 385.600 ;
        RECT 302.100 376.400 302.700 385.600 ;
        RECT 310.000 383.600 310.800 384.400 ;
        RECT 305.200 379.600 306.000 380.400 ;
        RECT 302.000 375.600 302.800 376.400 ;
        RECT 305.300 374.400 305.900 379.600 ;
        RECT 302.000 373.600 302.800 374.400 ;
        RECT 305.200 373.600 306.000 374.400 ;
        RECT 302.100 370.400 302.700 373.600 ;
        RECT 310.100 370.400 310.700 383.600 ;
        RECT 311.700 380.400 312.300 387.600 ;
        RECT 311.600 379.600 312.400 380.400 ;
        RECT 311.600 377.600 312.400 378.400 ;
        RECT 302.000 369.600 302.800 370.400 ;
        RECT 310.000 369.600 310.800 370.400 ;
        RECT 316.400 366.200 317.200 377.800 ;
        RECT 318.100 376.400 318.700 387.600 ;
        RECT 318.000 375.600 318.800 376.400 ;
        RECT 319.700 372.400 320.300 409.600 ;
        RECT 321.200 406.200 322.000 417.800 ;
        RECT 322.800 413.600 323.600 414.400 ;
        RECT 322.900 412.400 323.500 413.600 ;
        RECT 322.800 411.600 323.600 412.400 ;
        RECT 329.200 411.600 330.000 412.600 ;
        RECT 330.800 406.200 331.600 417.800 ;
        RECT 334.000 410.200 334.800 415.800 ;
        RECT 340.400 413.600 341.200 414.400 ;
        RECT 338.800 412.300 339.600 412.400 ;
        RECT 340.500 412.300 341.100 413.600 ;
        RECT 338.800 411.700 341.100 412.300 ;
        RECT 338.800 411.600 339.600 411.700 ;
        RECT 345.200 411.600 346.000 412.400 ;
        RECT 354.800 411.600 355.600 412.400 ;
        RECT 324.400 397.600 325.200 398.400 ;
        RECT 330.800 397.600 331.600 398.400 ;
        RECT 324.500 392.400 325.100 397.600 ;
        RECT 327.600 393.600 328.400 394.400 ;
        RECT 324.400 391.600 325.200 392.400 ;
        RECT 326.000 391.600 326.800 392.400 ;
        RECT 327.700 390.400 328.300 393.600 ;
        RECT 321.200 389.600 322.000 390.400 ;
        RECT 327.600 389.600 328.400 390.400 ;
        RECT 322.800 387.600 323.600 388.400 ;
        RECT 322.900 386.400 323.500 387.600 ;
        RECT 327.700 386.400 328.300 389.600 ;
        RECT 322.800 385.600 323.600 386.400 ;
        RECT 327.600 385.600 328.400 386.400 ;
        RECT 322.800 379.600 323.600 380.400 ;
        RECT 319.600 371.600 320.400 372.400 ;
        RECT 306.800 363.600 307.600 364.400 ;
        RECT 303.600 351.600 304.400 352.400 ;
        RECT 292.400 349.600 293.200 350.400 ;
        RECT 294.000 349.600 294.800 350.400 ;
        RECT 298.800 349.600 299.600 350.400 ;
        RECT 294.100 348.400 294.700 349.600 ;
        RECT 286.000 347.600 286.800 348.400 ;
        RECT 294.000 347.600 294.800 348.400 ;
        RECT 284.400 345.600 285.200 346.400 ;
        RECT 295.600 345.600 296.400 346.400 ;
        RECT 302.000 345.600 302.800 346.400 ;
        RECT 282.800 337.600 283.600 338.400 ;
        RECT 284.500 336.400 285.100 345.600 ;
        RECT 298.800 343.600 299.600 344.400 ;
        RECT 298.900 336.400 299.500 343.600 ;
        RECT 306.900 336.400 307.500 363.600 ;
        RECT 322.900 352.400 323.500 379.600 ;
        RECT 330.900 378.400 331.500 397.600 ;
        RECT 334.000 384.200 334.800 395.800 ;
        RECT 342.000 389.400 342.800 390.200 ;
        RECT 342.100 388.400 342.700 389.400 ;
        RECT 338.800 387.600 339.600 388.400 ;
        RECT 342.000 387.600 342.800 388.400 ;
        RECT 324.400 371.800 325.200 372.600 ;
        RECT 324.500 370.400 325.100 371.800 ;
        RECT 324.400 369.600 325.200 370.400 ;
        RECT 326.000 366.200 326.800 377.800 ;
        RECT 330.800 377.600 331.600 378.400 ;
        RECT 329.200 370.200 330.000 375.800 ;
        RECT 335.600 366.200 336.400 377.800 ;
        RECT 338.900 372.400 339.500 387.600 ;
        RECT 343.600 384.200 344.400 395.800 ;
        RECT 346.800 386.200 347.600 391.800 ;
        RECT 348.400 389.600 349.200 390.400 ;
        RECT 353.200 389.600 354.000 390.400 ;
        RECT 354.900 388.400 355.500 411.600 ;
        RECT 356.400 403.600 357.200 404.400 ;
        RECT 366.000 404.200 366.800 417.800 ;
        RECT 367.600 404.200 368.400 417.800 ;
        RECT 369.200 404.200 370.000 417.800 ;
        RECT 370.800 406.200 371.600 417.800 ;
        RECT 372.400 415.600 373.200 416.400 ;
        RECT 372.500 414.400 373.100 415.600 ;
        RECT 372.400 413.600 373.200 414.400 ;
        RECT 367.600 401.600 368.400 402.400 ;
        RECT 361.200 389.600 362.000 390.400 ;
        RECT 348.400 387.600 349.200 388.400 ;
        RECT 354.800 387.600 355.600 388.400 ;
        RECT 358.000 387.600 358.800 388.400 ;
        RECT 361.300 386.400 361.900 389.600 ;
        RECT 351.600 386.300 352.400 386.400 ;
        RECT 350.100 385.700 352.400 386.300 ;
        RECT 343.600 373.600 344.400 374.400 ;
        RECT 343.700 372.600 344.300 373.600 ;
        RECT 338.800 371.600 339.600 372.400 ;
        RECT 343.600 371.800 344.400 372.600 ;
        RECT 334.000 361.600 334.800 362.400 ;
        RECT 326.000 355.600 326.800 356.400 ;
        RECT 330.800 353.600 331.600 354.400 ;
        RECT 322.800 351.600 323.600 352.400 ;
        RECT 313.200 349.600 314.000 350.400 ;
        RECT 314.800 349.600 315.600 350.400 ;
        RECT 326.000 349.600 326.800 350.400 ;
        RECT 313.300 346.400 313.900 349.600 ;
        RECT 326.100 348.400 326.700 349.600 ;
        RECT 321.200 347.600 322.000 348.400 ;
        RECT 326.000 347.600 326.800 348.400 ;
        RECT 327.600 347.600 328.400 348.400 ;
        RECT 321.300 346.400 321.900 347.600 ;
        RECT 308.400 345.600 309.200 346.400 ;
        RECT 310.000 345.600 310.800 346.400 ;
        RECT 313.200 345.600 314.000 346.400 ;
        RECT 321.200 345.600 322.000 346.400 ;
        RECT 308.500 340.400 309.100 345.600 ;
        RECT 311.600 343.600 312.400 344.400 ;
        RECT 311.700 342.400 312.300 343.600 ;
        RECT 311.600 341.600 312.400 342.400 ;
        RECT 313.300 340.400 313.900 345.600 ;
        RECT 327.700 344.400 328.300 347.600 ;
        RECT 330.900 346.400 331.500 353.600 ;
        RECT 330.800 345.600 331.600 346.400 ;
        RECT 319.600 343.600 320.400 344.400 ;
        RECT 327.600 343.600 328.400 344.400 ;
        RECT 318.000 341.600 318.800 342.400 ;
        RECT 308.400 339.600 309.200 340.400 ;
        RECT 311.600 339.600 312.400 340.400 ;
        RECT 313.200 339.600 314.000 340.400 ;
        RECT 311.700 336.400 312.300 339.600 ;
        RECT 314.800 337.600 315.600 338.400 ;
        RECT 281.200 335.600 282.000 336.400 ;
        RECT 284.400 335.600 285.200 336.400 ;
        RECT 298.800 335.600 299.600 336.400 ;
        RECT 302.000 335.600 302.800 336.400 ;
        RECT 306.800 335.600 307.600 336.400 ;
        RECT 311.600 335.600 312.400 336.400 ;
        RECT 273.200 333.600 274.000 334.400 ;
        RECT 274.800 333.600 275.600 334.400 ;
        RECT 276.400 333.600 277.200 334.400 ;
        RECT 273.300 332.400 273.900 333.600 ;
        RECT 274.900 332.400 275.500 333.600 ;
        RECT 273.200 331.600 274.000 332.400 ;
        RECT 274.800 331.600 275.600 332.400 ;
        RECT 276.500 330.400 277.100 333.600 ;
        RECT 284.500 332.400 285.100 335.600 ;
        RECT 300.400 333.600 301.200 334.400 ;
        RECT 284.400 331.600 285.200 332.400 ;
        RECT 295.600 331.600 296.400 332.400 ;
        RECT 276.400 329.600 277.200 330.400 ;
        RECT 279.600 329.600 280.400 330.400 ;
        RECT 276.400 325.600 277.200 326.400 ;
        RECT 289.200 323.600 290.000 324.400 ;
        RECT 273.200 317.600 274.000 318.400 ;
        RECT 271.600 311.600 272.400 312.400 ;
        RECT 271.700 310.400 272.300 311.600 ;
        RECT 263.600 309.600 264.400 310.400 ;
        RECT 266.800 309.600 267.600 310.400 ;
        RECT 271.600 309.600 272.400 310.400 ;
        RECT 257.200 307.600 258.000 308.400 ;
        RECT 239.600 286.200 240.400 297.800 ;
        RECT 244.400 297.700 246.700 298.300 ;
        RECT 244.400 297.600 245.200 297.700 ;
        RECT 254.000 297.600 254.800 298.400 ;
        RECT 246.000 295.600 246.800 296.400 ;
        RECT 246.100 294.400 246.700 295.600 ;
        RECT 247.600 295.000 248.400 295.800 ;
        RECT 253.800 295.600 254.600 295.800 ;
        RECT 249.000 295.000 254.600 295.600 ;
        RECT 246.000 293.600 246.800 294.400 ;
        RECT 247.600 294.200 248.200 295.000 ;
        RECT 249.000 294.800 249.800 295.000 ;
        RECT 252.400 294.800 253.200 295.000 ;
        RECT 247.600 293.600 253.200 294.200 ;
        RECT 246.000 291.600 246.800 292.400 ;
        RECT 247.600 290.200 248.200 293.600 ;
        RECT 252.600 292.200 253.200 293.600 ;
        RECT 252.600 291.400 253.400 292.200 ;
        RECT 254.000 290.200 254.600 295.000 ;
        RECT 255.600 294.300 256.400 294.400 ;
        RECT 257.300 294.300 257.900 307.600 ;
        RECT 278.000 304.200 278.800 315.800 ;
        RECT 286.000 309.400 286.800 310.400 ;
        RECT 282.800 307.600 283.600 308.400 ;
        RECT 255.600 293.700 257.900 294.300 ;
        RECT 255.600 293.600 256.400 293.700 ;
        RECT 247.600 289.400 248.400 290.200 ;
        RECT 253.800 289.400 254.600 290.200 ;
        RECT 262.000 286.200 262.800 297.800 ;
        RECT 270.000 293.600 270.800 294.400 ;
        RECT 270.100 292.600 270.700 293.600 ;
        RECT 263.600 291.600 264.400 292.400 ;
        RECT 270.000 291.800 270.800 292.600 ;
        RECT 257.200 283.600 258.000 284.400 ;
        RECT 260.400 283.600 261.200 284.400 ;
        RECT 239.600 271.600 240.400 272.400 ;
        RECT 241.200 271.600 242.000 272.400 ;
        RECT 249.200 271.600 250.000 272.400 ;
        RECT 258.800 271.600 259.600 272.400 ;
        RECT 238.000 269.600 238.800 270.400 ;
        RECT 239.700 268.400 240.300 271.600 ;
        RECT 241.300 270.400 241.900 271.600 ;
        RECT 249.300 270.400 249.900 271.600 ;
        RECT 241.200 269.600 242.000 270.400 ;
        RECT 242.800 269.600 243.600 270.400 ;
        RECT 249.200 269.600 250.000 270.400 ;
        RECT 250.800 269.600 251.600 270.400 ;
        RECT 257.200 269.600 258.000 270.400 ;
        RECT 239.600 267.600 240.400 268.400 ;
        RECT 244.400 267.600 245.200 268.400 ;
        RECT 246.000 267.600 246.800 268.400 ;
        RECT 250.800 267.600 251.600 268.400 ;
        RECT 255.600 267.600 256.400 268.800 ;
        RECT 257.300 268.400 257.900 269.600 ;
        RECT 257.200 267.600 258.000 268.400 ;
        RECT 244.500 266.400 245.100 267.600 ;
        RECT 234.800 265.600 235.600 266.400 ;
        RECT 244.400 265.600 245.200 266.400 ;
        RECT 260.500 260.400 261.100 283.600 ;
        RECT 262.000 273.600 262.800 274.400 ;
        RECT 262.000 267.600 262.800 268.400 ;
        RECT 262.100 266.400 262.700 267.600 ;
        RECT 262.000 265.600 262.800 266.400 ;
        RECT 260.400 259.600 261.200 260.400 ;
        RECT 230.000 255.600 230.800 256.400 ;
        RECT 231.600 255.600 232.400 256.400 ;
        RECT 230.100 252.400 230.700 255.600 ;
        RECT 225.200 251.600 226.000 252.400 ;
        RECT 230.000 251.600 230.800 252.400 ;
        RECT 210.800 233.600 211.600 234.400 ;
        RECT 204.400 229.700 206.700 230.300 ;
        RECT 210.900 230.200 211.500 233.600 ;
        RECT 204.400 229.600 205.200 229.700 ;
        RECT 210.800 229.400 211.600 230.200 ;
        RECT 212.400 224.200 213.200 235.800 ;
        RECT 215.600 226.200 216.400 231.800 ;
        RECT 217.200 223.600 218.000 224.400 ;
        RECT 222.000 224.200 222.800 235.800 ;
        RECT 223.600 230.300 224.400 230.400 ;
        RECT 225.300 230.300 225.900 251.600 ;
        RECT 233.200 246.200 234.000 257.800 ;
        RECT 241.200 257.600 242.000 258.400 ;
        RECT 236.400 250.200 237.200 255.800 ;
        RECT 241.300 252.400 241.900 257.600 ;
        RECT 241.200 251.600 242.000 252.400 ;
        RECT 247.600 246.200 248.400 257.800 ;
        RECT 255.600 253.600 256.400 254.400 ;
        RECT 255.700 252.600 256.300 253.600 ;
        RECT 255.600 251.800 256.400 252.600 ;
        RECT 257.200 246.200 258.000 257.800 ;
        RECT 262.000 257.600 262.800 258.400 ;
        RECT 258.800 253.600 259.600 254.400 ;
        RECT 258.900 252.400 259.500 253.600 ;
        RECT 258.800 251.600 259.600 252.400 ;
        RECT 238.000 243.600 238.800 244.400 ;
        RECT 242.800 243.600 243.600 244.400 ;
        RECT 230.000 231.600 230.800 232.400 ;
        RECT 223.600 229.700 225.900 230.300 ;
        RECT 230.100 230.200 230.700 231.600 ;
        RECT 223.600 229.600 224.400 229.700 ;
        RECT 230.000 229.400 230.800 230.200 ;
        RECT 231.600 224.200 232.400 235.800 ;
        RECT 238.100 234.400 238.700 243.600 ;
        RECT 238.000 233.600 238.800 234.400 ;
        RECT 239.600 233.600 240.400 234.400 ;
        RECT 239.700 232.400 240.300 233.600 ;
        RECT 234.800 226.200 235.600 231.800 ;
        RECT 239.600 231.600 240.400 232.400 ;
        RECT 242.900 230.400 243.500 243.600 ;
        RECT 242.800 229.600 243.600 230.400 ;
        RECT 238.000 227.600 238.800 228.400 ;
        RECT 236.400 225.600 237.200 226.400 ;
        RECT 236.500 224.400 237.100 225.600 ;
        RECT 238.100 224.400 238.700 227.600 ;
        RECT 244.400 226.200 245.200 231.800 ;
        RECT 246.000 229.600 246.800 230.400 ;
        RECT 246.100 228.400 246.700 229.600 ;
        RECT 246.000 227.600 246.800 228.400 ;
        RECT 236.400 223.600 237.200 224.400 ;
        RECT 238.000 223.600 238.800 224.400 ;
        RECT 247.600 224.200 248.400 235.800 ;
        RECT 249.200 229.400 250.000 230.200 ;
        RECT 249.300 228.400 249.900 229.400 ;
        RECT 249.200 227.600 250.000 228.400 ;
        RECT 257.200 224.200 258.000 235.800 ;
        RECT 258.900 234.400 259.500 251.600 ;
        RECT 260.400 250.200 261.200 255.800 ;
        RECT 263.700 252.400 264.300 291.600 ;
        RECT 271.600 286.200 272.400 297.800 ;
        RECT 274.800 290.200 275.600 295.800 ;
        RECT 281.200 286.200 282.000 297.800 ;
        RECT 282.900 292.400 283.500 307.600 ;
        RECT 287.600 304.200 288.400 315.800 ;
        RECT 289.300 314.400 289.900 323.600 ;
        RECT 289.200 313.600 290.000 314.400 ;
        RECT 290.800 306.200 291.600 311.800 ;
        RECT 292.400 307.600 293.200 308.400 ;
        RECT 297.200 303.600 298.000 304.400 ;
        RECT 282.800 291.600 283.600 292.400 ;
        RECT 289.200 291.600 290.000 292.600 ;
        RECT 282.800 289.600 283.600 290.400 ;
        RECT 276.400 283.600 277.200 284.400 ;
        RECT 268.400 273.600 269.200 274.400 ;
        RECT 268.500 272.400 269.100 273.600 ;
        RECT 268.400 271.600 269.200 272.400 ;
        RECT 271.400 271.800 272.200 272.600 ;
        RECT 278.000 271.800 278.800 272.600 ;
        RECT 265.200 269.600 266.000 270.400 ;
        RECT 271.400 267.000 272.000 271.800 ;
        RECT 274.000 268.400 274.800 268.600 ;
        RECT 278.200 268.400 278.800 271.800 ;
        RECT 274.000 267.800 278.800 268.400 ;
        RECT 273.200 267.000 274.000 267.200 ;
        RECT 276.600 267.000 277.400 267.200 ;
        RECT 278.200 267.000 278.800 267.800 ;
        RECT 279.600 267.600 280.400 268.400 ;
        RECT 281.200 267.600 282.000 268.400 ;
        RECT 271.400 266.200 272.200 267.000 ;
        RECT 273.200 266.400 277.400 267.000 ;
        RECT 278.000 266.200 278.800 267.000 ;
        RECT 279.700 266.400 280.300 267.600 ;
        RECT 282.900 266.400 283.500 289.600 ;
        RECT 290.800 286.200 291.600 297.800 ;
        RECT 294.000 290.200 294.800 295.800 ;
        RECT 297.300 290.400 297.900 303.600 ;
        RECT 300.500 294.400 301.100 333.600 ;
        RECT 302.100 332.400 302.700 335.600 ;
        RECT 314.900 334.400 315.500 337.600 ;
        RECT 318.100 336.400 318.700 341.600 ;
        RECT 319.700 336.400 320.300 343.600 ;
        RECT 332.400 339.600 333.200 340.400 ;
        RECT 318.000 335.600 318.800 336.400 ;
        RECT 319.600 335.600 320.400 336.400 ;
        RECT 306.800 333.600 307.600 334.400 ;
        RECT 314.800 333.600 315.600 334.400 ;
        RECT 302.000 331.600 302.800 332.400 ;
        RECT 319.700 332.300 320.300 335.600 ;
        RECT 324.200 335.000 325.000 335.800 ;
        RECT 326.000 335.000 330.200 335.600 ;
        RECT 330.800 335.000 331.600 335.800 ;
        RECT 322.800 333.600 323.600 334.400 ;
        RECT 321.200 332.300 322.000 332.400 ;
        RECT 319.700 331.700 322.000 332.300 ;
        RECT 321.200 331.600 322.000 331.700 ;
        RECT 310.000 329.600 310.800 330.400 ;
        RECT 324.200 330.200 324.800 335.000 ;
        RECT 326.000 334.800 326.800 335.000 ;
        RECT 329.400 334.800 330.200 335.000 ;
        RECT 331.000 334.200 331.600 335.000 ;
        RECT 332.500 334.400 333.100 339.600 ;
        RECT 334.100 338.400 334.700 361.600 ;
        RECT 337.200 344.200 338.000 355.800 ;
        RECT 338.900 350.400 339.500 371.600 ;
        RECT 345.200 366.200 346.000 377.800 ;
        RECT 348.400 370.200 349.200 375.800 ;
        RECT 350.100 374.400 350.700 385.700 ;
        RECT 351.600 385.600 352.400 385.700 ;
        RECT 361.200 385.600 362.000 386.400 ;
        RECT 364.400 385.600 365.200 386.400 ;
        RECT 367.700 386.300 368.300 401.600 ;
        RECT 369.200 389.600 370.000 390.400 ;
        RECT 369.300 388.400 369.900 389.600 ;
        RECT 369.200 387.600 370.000 388.400 ;
        RECT 367.700 385.700 369.900 386.300 ;
        RECT 351.600 375.600 352.400 376.400 ;
        RECT 350.000 373.600 350.800 374.400 ;
        RECT 350.100 372.400 350.700 373.600 ;
        RECT 351.700 372.400 352.300 375.600 ;
        RECT 361.300 374.400 361.900 385.600 ;
        RECT 362.800 383.600 363.600 384.400 ;
        RECT 362.900 376.400 363.500 383.600 ;
        RECT 362.800 375.600 363.600 376.400 ;
        RECT 364.500 374.400 365.100 385.600 ;
        RECT 369.300 378.400 369.900 385.700 ;
        RECT 372.500 378.400 373.100 413.600 ;
        RECT 374.000 406.200 374.800 417.800 ;
        RECT 377.200 406.200 378.000 417.800 ;
        RECT 378.800 404.200 379.600 417.800 ;
        RECT 380.400 404.200 381.200 417.800 ;
        RECT 401.200 415.600 402.000 416.400 ;
        RECT 386.800 413.600 387.600 414.400 ;
        RECT 390.000 413.600 390.800 414.400 ;
        RECT 385.200 411.600 386.000 412.400 ;
        RECT 386.900 410.400 387.500 413.600 ;
        RECT 393.200 411.600 394.000 412.400 ;
        RECT 386.800 409.600 387.600 410.400 ;
        RECT 401.300 408.400 401.900 415.600 ;
        RECT 401.200 407.600 402.000 408.400 ;
        RECT 402.800 403.600 403.600 404.400 ;
        RECT 410.800 403.600 411.600 404.400 ;
        RECT 412.400 404.200 413.200 417.800 ;
        RECT 414.000 404.200 414.800 417.800 ;
        RECT 415.600 404.200 416.400 417.800 ;
        RECT 417.200 406.200 418.000 417.800 ;
        RECT 418.800 415.600 419.600 416.400 ;
        RECT 420.400 406.200 421.200 417.800 ;
        RECT 423.600 406.200 424.400 417.800 ;
        RECT 425.200 404.200 426.000 417.800 ;
        RECT 426.800 404.200 427.600 417.800 ;
        RECT 450.800 415.600 451.600 416.400 ;
        RECT 433.200 413.600 434.000 414.400 ;
        RECT 436.400 413.600 437.200 414.400 ;
        RECT 431.600 411.600 432.400 412.400 ;
        RECT 433.300 410.400 433.900 413.600 ;
        RECT 441.200 411.600 442.000 412.400 ;
        RECT 433.200 409.600 434.000 410.400 ;
        RECT 450.900 408.400 451.500 415.600 ;
        RECT 457.200 411.600 458.000 412.400 ;
        RECT 450.800 407.600 451.600 408.400 ;
        RECT 402.900 400.400 403.500 403.600 ;
        RECT 402.800 399.600 403.600 400.400 ;
        RECT 374.000 389.600 374.800 390.400 ;
        RECT 377.200 389.600 378.000 390.400 ;
        RECT 374.100 388.400 374.700 389.600 ;
        RECT 374.000 387.600 374.800 388.400 ;
        RECT 369.200 377.600 370.000 378.400 ;
        RECT 372.400 377.600 373.200 378.400 ;
        RECT 374.100 376.400 374.700 387.600 ;
        RECT 390.000 383.600 390.800 384.400 ;
        RECT 394.800 384.200 395.600 395.800 ;
        RECT 396.400 389.600 397.200 390.400 ;
        RECT 402.800 389.400 403.600 390.400 ;
        RECT 402.800 385.600 403.600 386.400 ;
        RECT 386.800 378.300 387.600 378.400 ;
        RECT 385.300 377.700 387.600 378.300 ;
        RECT 385.300 376.400 385.900 377.700 ;
        RECT 386.800 377.600 387.600 377.700 ;
        RECT 390.100 376.400 390.700 383.600 ;
        RECT 367.600 375.600 368.400 376.400 ;
        RECT 372.400 376.300 373.200 376.400 ;
        RECT 374.000 376.300 374.800 376.400 ;
        RECT 372.400 375.700 374.800 376.300 ;
        RECT 372.400 375.600 373.200 375.700 ;
        RECT 374.000 375.600 374.800 375.700 ;
        RECT 382.000 375.600 382.800 376.400 ;
        RECT 385.200 375.600 386.000 376.400 ;
        RECT 390.000 375.600 390.800 376.400 ;
        RECT 361.200 373.600 362.000 374.400 ;
        RECT 362.800 373.600 363.600 374.400 ;
        RECT 364.400 373.600 365.200 374.400 ;
        RECT 362.900 372.400 363.500 373.600 ;
        RECT 367.700 372.400 368.300 375.600 ;
        RECT 382.100 374.400 382.700 375.600 ;
        RECT 385.300 374.400 385.900 375.600 ;
        RECT 382.000 373.600 382.800 374.400 ;
        RECT 385.200 373.600 386.000 374.400 ;
        RECT 350.000 371.600 350.800 372.400 ;
        RECT 351.600 371.600 352.400 372.400 ;
        RECT 353.200 371.600 354.000 372.400 ;
        RECT 362.800 371.600 363.600 372.400 ;
        RECT 364.400 371.600 365.200 372.400 ;
        RECT 367.600 371.600 368.400 372.400 ;
        RECT 375.600 371.600 376.400 372.400 ;
        RECT 377.200 371.600 378.000 372.400 ;
        RECT 380.400 371.600 381.200 372.400 ;
        RECT 353.300 370.400 353.900 371.600 ;
        RECT 353.200 369.600 354.000 370.400 ;
        RECT 354.800 369.600 355.600 370.400 ;
        RECT 338.800 349.600 339.600 350.400 ;
        RECT 345.200 349.400 346.000 350.400 ;
        RECT 345.200 345.600 346.000 346.400 ;
        RECT 334.000 337.600 334.800 338.400 ;
        RECT 326.800 333.600 331.600 334.200 ;
        RECT 332.400 333.600 333.200 334.400 ;
        RECT 326.800 333.400 327.600 333.600 ;
        RECT 331.000 330.200 331.600 333.600 ;
        RECT 324.200 329.400 325.000 330.200 ;
        RECT 330.800 329.400 331.600 330.200 ;
        RECT 302.000 327.600 302.800 328.400 ;
        RECT 338.800 326.200 339.600 337.800 ;
        RECT 345.300 334.400 345.900 345.600 ;
        RECT 346.800 344.200 347.600 355.800 ;
        RECT 348.400 347.600 349.200 348.400 ;
        RECT 350.000 346.200 350.800 351.800 ;
        RECT 351.600 349.600 352.400 350.400 ;
        RECT 353.300 346.400 353.900 369.600 ;
        RECT 354.900 368.400 355.500 369.600 ;
        RECT 354.800 367.600 355.600 368.400 ;
        RECT 353.200 345.600 354.000 346.400 ;
        RECT 354.800 343.600 355.600 344.400 ;
        RECT 359.600 344.200 360.400 355.800 ;
        RECT 364.500 350.400 365.100 371.600 ;
        RECT 375.700 370.400 376.300 371.600 ;
        RECT 377.300 370.400 377.900 371.600 ;
        RECT 380.500 370.400 381.100 371.600 ;
        RECT 366.000 369.600 366.800 370.400 ;
        RECT 375.600 369.600 376.400 370.400 ;
        RECT 377.200 369.600 378.000 370.400 ;
        RECT 380.400 369.600 381.200 370.400 ;
        RECT 366.100 368.400 366.700 369.600 ;
        RECT 366.000 367.600 366.800 368.400 ;
        RECT 377.300 368.300 377.900 369.600 ;
        RECT 375.700 367.700 377.900 368.300 ;
        RECT 369.200 363.600 370.000 364.400 ;
        RECT 369.300 358.400 369.900 363.600 ;
        RECT 369.200 357.600 370.000 358.400 ;
        RECT 364.400 349.600 365.200 350.400 ;
        RECT 367.600 345.600 368.400 346.400 ;
        RECT 356.400 339.600 357.200 340.400 ;
        RECT 356.500 338.400 357.100 339.600 ;
        RECT 345.200 333.600 346.000 334.400 ;
        RECT 340.400 331.600 341.200 332.400 ;
        RECT 346.800 331.600 347.600 332.600 ;
        RECT 326.000 323.600 326.800 324.400 ;
        RECT 326.100 320.400 326.700 323.600 ;
        RECT 326.000 319.600 326.800 320.400 ;
        RECT 302.000 304.200 302.800 315.800 ;
        RECT 310.000 313.600 310.800 314.400 ;
        RECT 303.600 309.600 304.400 310.400 ;
        RECT 310.100 310.200 310.700 313.600 ;
        RECT 303.700 308.400 304.300 309.600 ;
        RECT 310.000 309.400 310.800 310.200 ;
        RECT 303.600 307.600 304.400 308.400 ;
        RECT 311.600 304.200 312.400 315.800 ;
        RECT 337.200 315.600 338.000 316.400 ;
        RECT 314.800 306.200 315.600 311.800 ;
        RECT 316.400 311.600 317.200 312.400 ;
        RECT 322.800 311.600 323.600 312.400 ;
        RECT 327.600 311.600 328.400 312.400 ;
        RECT 330.800 311.600 331.600 312.400 ;
        RECT 332.400 311.600 333.200 312.400 ;
        RECT 316.500 310.400 317.100 311.600 ;
        RECT 327.700 310.400 328.300 311.600 ;
        RECT 330.900 310.400 331.500 311.600 ;
        RECT 316.400 309.600 317.200 310.400 ;
        RECT 327.600 309.600 328.400 310.400 ;
        RECT 330.800 309.600 331.600 310.400 ;
        RECT 321.200 307.600 322.000 308.400 ;
        RECT 330.800 307.600 331.600 308.400 ;
        RECT 306.800 295.000 307.600 295.800 ;
        RECT 308.200 295.000 312.400 295.600 ;
        RECT 313.400 295.000 314.200 295.800 ;
        RECT 300.400 293.600 301.200 294.400 ;
        RECT 305.200 293.600 306.000 294.400 ;
        RECT 306.800 294.200 307.400 295.000 ;
        RECT 308.200 294.800 309.000 295.000 ;
        RECT 311.600 294.800 312.400 295.000 ;
        RECT 306.800 293.600 311.600 294.200 ;
        RECT 303.600 291.600 304.400 292.400 ;
        RECT 297.200 289.600 298.000 290.400 ;
        RECT 302.000 289.600 302.800 290.400 ;
        RECT 303.600 289.600 304.400 290.400 ;
        RECT 285.800 271.800 286.600 272.600 ;
        RECT 292.400 271.800 293.200 272.600 ;
        RECT 284.400 267.600 285.200 268.400 ;
        RECT 284.500 266.400 285.100 267.600 ;
        RECT 285.800 267.000 286.400 271.800 ;
        RECT 288.400 268.400 289.200 268.600 ;
        RECT 292.600 268.400 293.200 271.800 ;
        RECT 303.700 270.400 304.300 289.600 ;
        RECT 305.300 274.400 305.900 293.600 ;
        RECT 306.800 290.200 307.400 293.600 ;
        RECT 310.800 293.400 311.600 293.600 ;
        RECT 313.600 290.200 314.200 295.000 ;
        RECT 321.300 294.400 321.900 307.600 ;
        RECT 332.500 306.400 333.100 311.600 ;
        RECT 335.600 309.600 336.400 310.400 ;
        RECT 337.300 308.400 337.900 315.600 ;
        RECT 338.800 311.600 339.600 312.400 ;
        RECT 338.900 308.400 339.500 311.600 ;
        RECT 337.200 307.600 338.000 308.400 ;
        RECT 338.800 307.600 339.600 308.400 ;
        RECT 332.400 305.600 333.200 306.400 ;
        RECT 322.800 303.600 323.600 304.400 ;
        RECT 322.900 294.400 323.500 303.600 ;
        RECT 327.600 295.600 328.400 296.400 ;
        RECT 321.200 293.600 322.000 294.400 ;
        RECT 322.800 293.600 323.600 294.400 ;
        RECT 306.800 289.400 307.600 290.200 ;
        RECT 313.400 289.400 314.200 290.200 ;
        RECT 316.400 289.600 317.200 290.400 ;
        RECT 318.000 283.600 318.800 284.400 ;
        RECT 305.200 273.600 306.000 274.400 ;
        RECT 313.200 273.600 314.000 274.400 ;
        RECT 295.600 269.600 296.400 270.400 ;
        RECT 300.400 269.600 301.200 270.400 ;
        RECT 303.600 269.600 304.400 270.400 ;
        RECT 295.700 268.400 296.300 269.600 ;
        RECT 305.300 268.400 305.900 273.600 ;
        RECT 313.300 272.400 313.900 273.600 ;
        RECT 311.600 271.600 312.400 272.400 ;
        RECT 313.200 271.600 314.000 272.400 ;
        RECT 311.700 270.400 312.300 271.600 ;
        RECT 308.400 270.300 309.200 270.400 ;
        RECT 308.400 269.700 310.700 270.300 ;
        RECT 308.400 269.600 309.200 269.700 ;
        RECT 288.400 267.800 293.200 268.400 ;
        RECT 287.600 267.000 288.400 267.200 ;
        RECT 291.000 267.000 291.800 267.200 ;
        RECT 292.600 267.000 293.200 267.800 ;
        RECT 294.000 267.600 294.800 268.400 ;
        RECT 295.600 267.600 296.400 268.400 ;
        RECT 305.200 267.600 306.000 268.400 ;
        RECT 308.400 267.600 309.200 268.400 ;
        RECT 279.600 265.600 280.400 266.400 ;
        RECT 282.800 265.600 283.600 266.400 ;
        RECT 284.400 265.600 285.200 266.400 ;
        RECT 285.800 266.200 286.600 267.000 ;
        RECT 287.600 266.400 291.800 267.000 ;
        RECT 292.400 266.200 293.200 267.000 ;
        RECT 305.200 265.600 306.000 266.400 ;
        RECT 310.100 264.400 310.700 269.700 ;
        RECT 311.600 269.600 312.400 270.400 ;
        RECT 316.400 269.600 317.200 270.400 ;
        RECT 318.100 268.400 318.700 283.600 ;
        RECT 321.300 272.300 321.900 293.600 ;
        RECT 319.700 271.700 321.900 272.300 ;
        RECT 319.700 268.400 320.300 271.700 ;
        RECT 327.700 270.400 328.300 295.600 ;
        RECT 334.000 286.200 334.800 297.800 ;
        RECT 340.500 294.400 341.100 331.600 ;
        RECT 348.400 326.200 349.200 337.800 ;
        RECT 356.400 337.600 357.200 338.400 ;
        RECT 351.600 330.200 352.400 335.800 ;
        RECT 354.800 335.600 355.600 336.400 ;
        RECT 354.900 332.400 355.500 335.600 ;
        RECT 353.200 331.600 354.000 332.400 ;
        RECT 354.800 331.600 355.600 332.400 ;
        RECT 351.600 327.600 352.400 328.400 ;
        RECT 351.700 318.400 352.300 327.600 ;
        RECT 361.200 326.200 362.000 337.800 ;
        RECT 367.700 334.400 368.300 345.600 ;
        RECT 369.200 344.200 370.000 355.800 ;
        RECT 370.800 347.600 371.600 348.400 ;
        RECT 372.400 346.200 373.200 351.800 ;
        RECT 374.000 349.600 374.800 350.400 ;
        RECT 375.700 340.400 376.300 367.700 ;
        RECT 380.400 367.600 381.200 368.400 ;
        RECT 391.600 366.200 392.400 377.800 ;
        RECT 393.200 377.600 394.000 378.400 ;
        RECT 393.300 372.400 393.900 377.600 ;
        RECT 393.200 371.600 394.000 372.400 ;
        RECT 399.600 371.600 400.400 372.600 ;
        RECT 401.200 366.200 402.000 377.800 ;
        RECT 378.800 357.600 379.600 358.400 ;
        RECT 378.900 348.400 379.500 357.600 ;
        RECT 380.200 351.800 381.000 352.600 ;
        RECT 386.800 351.800 387.600 352.600 ;
        RECT 378.800 347.600 379.600 348.400 ;
        RECT 380.200 347.000 380.800 351.800 ;
        RECT 382.800 348.400 383.600 348.600 ;
        RECT 387.000 348.400 387.600 351.800 ;
        RECT 382.800 347.800 387.600 348.400 ;
        RECT 382.000 347.000 382.800 347.200 ;
        RECT 385.400 347.000 386.200 347.200 ;
        RECT 387.000 347.000 387.600 347.800 ;
        RECT 391.600 347.600 392.400 348.400 ;
        RECT 380.200 346.200 381.000 347.000 ;
        RECT 382.000 346.400 386.200 347.000 ;
        RECT 386.800 346.200 387.600 347.000 ;
        RECT 383.600 343.600 384.400 344.400 ;
        RECT 390.000 343.600 390.800 344.400 ;
        RECT 375.600 339.600 376.400 340.400 ;
        RECT 367.600 333.600 368.400 334.400 ;
        RECT 369.200 331.600 370.000 332.600 ;
        RECT 370.800 326.200 371.600 337.800 ;
        RECT 374.000 330.200 374.800 335.800 ;
        RECT 375.700 334.400 376.300 339.600 ;
        RECT 375.600 333.600 376.400 334.400 ;
        RECT 382.000 333.600 382.800 334.400 ;
        RECT 351.600 317.600 352.400 318.400 ;
        RECT 364.400 317.600 365.200 318.400 ;
        RECT 342.000 315.600 342.800 316.400 ;
        RECT 342.100 310.400 342.700 315.600 ;
        RECT 353.200 313.600 354.000 314.400 ;
        RECT 354.800 313.600 355.600 314.400 ;
        RECT 343.600 311.600 344.400 312.400 ;
        RECT 345.200 311.600 346.000 312.400 ;
        RECT 343.700 310.400 344.300 311.600 ;
        RECT 353.300 310.400 353.900 313.600 ;
        RECT 342.000 309.600 342.800 310.400 ;
        RECT 343.600 309.600 344.400 310.400 ;
        RECT 348.400 309.600 349.200 310.400 ;
        RECT 353.200 309.600 354.000 310.400 ;
        RECT 354.900 308.400 355.500 313.600 ;
        RECT 356.400 311.800 357.200 312.600 ;
        RECT 363.000 311.800 363.800 312.600 ;
        RECT 356.400 308.400 357.000 311.800 ;
        RECT 360.400 308.400 361.200 308.600 ;
        RECT 343.600 307.600 344.400 308.400 ;
        RECT 354.800 307.600 355.600 308.400 ;
        RECT 356.400 307.800 361.200 308.400 ;
        RECT 343.700 306.400 344.300 307.600 ;
        RECT 356.400 307.000 357.000 307.800 ;
        RECT 357.800 307.000 358.600 307.200 ;
        RECT 361.200 307.000 362.000 307.200 ;
        RECT 363.200 307.000 363.800 311.800 ;
        RECT 364.500 308.400 365.100 317.600 ;
        RECT 367.800 311.800 368.600 312.600 ;
        RECT 374.000 311.800 374.800 312.600 ;
        RECT 375.700 312.400 376.300 333.600 ;
        RECT 383.700 332.400 384.300 343.600 ;
        RECT 390.100 336.400 390.700 343.600 ;
        RECT 391.700 340.400 392.300 347.600 ;
        RECT 393.200 343.600 394.000 344.400 ;
        RECT 398.000 344.200 398.800 355.800 ;
        RECT 402.900 348.400 403.500 385.600 ;
        RECT 404.400 384.200 405.200 395.800 ;
        RECT 407.600 386.200 408.400 391.800 ;
        RECT 410.900 388.400 411.500 403.600 ;
        RECT 414.000 389.600 414.800 390.400 ;
        RECT 418.800 389.600 419.600 390.400 ;
        RECT 423.600 390.300 424.400 390.400 ;
        RECT 422.100 389.700 424.400 390.300 ;
        RECT 418.900 388.400 419.500 389.600 ;
        RECT 422.100 388.400 422.700 389.700 ;
        RECT 423.600 389.600 424.400 389.700 ;
        RECT 428.400 389.600 429.200 390.400 ;
        RECT 410.800 387.600 411.600 388.400 ;
        RECT 418.800 387.600 419.600 388.400 ;
        RECT 422.000 387.600 422.800 388.400 ;
        RECT 404.400 370.200 405.200 375.800 ;
        RECT 410.900 374.400 411.500 387.600 ;
        RECT 434.800 383.600 435.600 384.400 ;
        RECT 444.400 383.600 445.200 384.400 ;
        RECT 434.900 380.400 435.500 383.600 ;
        RECT 444.500 380.400 445.100 383.600 ;
        RECT 434.800 379.600 435.600 380.400 ;
        RECT 439.600 379.600 440.400 380.400 ;
        RECT 444.400 379.600 445.200 380.400 ;
        RECT 420.400 377.600 421.200 378.400 ;
        RECT 410.800 373.600 411.600 374.400 ;
        RECT 406.000 371.600 406.800 372.400 ;
        RECT 406.000 349.400 406.800 350.400 ;
        RECT 402.800 347.600 403.600 348.400 ;
        RECT 393.300 340.400 393.900 343.600 ;
        RECT 391.600 339.600 392.400 340.400 ;
        RECT 393.200 339.600 394.000 340.400 ;
        RECT 390.000 335.600 390.800 336.400 ;
        RECT 386.800 333.600 387.600 334.400 ;
        RECT 388.400 333.600 389.200 334.400 ;
        RECT 390.000 333.600 390.800 334.400 ;
        RECT 386.900 332.400 387.500 333.600 ;
        RECT 377.200 331.600 378.000 332.400 ;
        RECT 380.400 331.600 381.200 332.400 ;
        RECT 383.600 331.600 384.400 332.400 ;
        RECT 385.200 331.600 386.000 332.400 ;
        RECT 386.800 331.600 387.600 332.400 ;
        RECT 377.300 328.400 377.900 331.600 ;
        RECT 378.800 329.600 379.600 330.400 ;
        RECT 377.200 327.600 378.000 328.400 ;
        RECT 377.200 323.600 378.000 324.400 ;
        RECT 377.300 316.400 377.900 323.600 ;
        RECT 378.900 318.400 379.500 329.600 ;
        RECT 380.500 324.400 381.100 331.600 ;
        RECT 383.600 329.600 384.400 330.400 ;
        RECT 380.400 323.600 381.200 324.400 ;
        RECT 382.000 321.600 382.800 322.400 ;
        RECT 378.800 317.600 379.600 318.400 ;
        RECT 377.200 315.600 378.000 316.400 ;
        RECT 364.400 307.600 365.200 308.400 ;
        RECT 366.000 307.600 366.800 308.400 ;
        RECT 343.600 305.600 344.400 306.400 ;
        RECT 356.400 306.200 357.200 307.000 ;
        RECT 357.800 306.400 362.000 307.000 ;
        RECT 363.000 306.200 363.800 307.000 ;
        RECT 367.800 307.000 368.400 311.800 ;
        RECT 369.000 309.800 369.800 310.600 ;
        RECT 369.200 308.400 369.800 309.800 ;
        RECT 374.200 308.400 374.800 311.800 ;
        RECT 375.600 311.600 376.400 312.400 ;
        RECT 375.700 310.400 376.300 311.600 ;
        RECT 375.600 309.600 376.400 310.400 ;
        RECT 380.400 309.600 381.200 310.400 ;
        RECT 369.200 307.800 374.800 308.400 ;
        RECT 369.200 307.000 370.000 307.200 ;
        RECT 372.600 307.000 373.400 307.200 ;
        RECT 374.200 307.000 374.800 307.800 ;
        RECT 375.600 307.600 376.400 308.400 ;
        RECT 377.200 307.600 378.000 308.400 ;
        RECT 367.800 306.400 373.400 307.000 ;
        RECT 367.800 306.200 368.600 306.400 ;
        RECT 374.000 306.200 374.800 307.000 ;
        RECT 375.700 306.400 376.300 307.600 ;
        RECT 375.600 305.600 376.400 306.400 ;
        RECT 343.700 300.400 344.300 305.600 ;
        RECT 369.200 303.600 370.000 304.400 ;
        RECT 343.600 299.600 344.400 300.400 ;
        RECT 367.600 299.600 368.400 300.400 ;
        RECT 367.700 298.400 368.300 299.600 ;
        RECT 340.400 293.600 341.200 294.400 ;
        RECT 340.500 292.400 341.100 293.600 ;
        RECT 340.400 291.600 341.200 292.400 ;
        RECT 342.000 291.800 342.800 292.600 ;
        RECT 342.100 288.400 342.700 291.800 ;
        RECT 342.000 287.600 342.800 288.400 ;
        RECT 343.600 286.200 344.400 297.800 ;
        RECT 346.800 290.200 347.600 295.800 ;
        RECT 353.200 286.200 354.000 297.800 ;
        RECT 361.200 293.600 362.000 294.400 ;
        RECT 361.300 292.600 361.900 293.600 ;
        RECT 354.800 291.600 355.600 292.400 ;
        RECT 361.200 291.800 362.000 292.600 ;
        RECT 362.800 286.200 363.600 297.800 ;
        RECT 367.600 297.600 368.400 298.400 ;
        RECT 366.000 290.200 366.800 295.800 ;
        RECT 369.300 294.400 369.900 303.600 ;
        RECT 377.300 302.400 377.900 307.600 ;
        RECT 382.100 306.400 382.700 321.600 ;
        RECT 385.300 318.400 385.900 331.600 ;
        RECT 388.500 324.400 389.100 333.600 ;
        RECT 388.400 323.600 389.200 324.400 ;
        RECT 390.100 322.400 390.700 333.600 ;
        RECT 393.200 329.600 394.000 330.400 ;
        RECT 391.600 323.600 392.400 324.400 ;
        RECT 390.000 321.600 390.800 322.400 ;
        RECT 385.200 317.600 386.000 318.400 ;
        RECT 391.700 310.400 392.300 323.600 ;
        RECT 385.200 309.600 386.000 310.400 ;
        RECT 388.400 309.600 389.200 310.400 ;
        RECT 391.600 309.600 392.400 310.400 ;
        RECT 386.800 307.600 387.600 308.400 ;
        RECT 382.000 305.600 382.800 306.400 ;
        RECT 388.400 305.600 389.200 306.400 ;
        RECT 391.700 304.400 392.300 309.600 ;
        RECT 393.300 308.400 393.900 329.600 ;
        RECT 399.600 326.200 400.400 337.800 ;
        RECT 402.900 332.400 403.500 347.600 ;
        RECT 407.600 344.200 408.400 355.800 ;
        RECT 410.900 354.400 411.500 373.600 ;
        RECT 418.800 371.600 419.600 372.400 ;
        RECT 412.400 363.600 413.200 364.400 ;
        RECT 410.800 353.600 411.600 354.400 ;
        RECT 418.900 352.400 419.500 371.600 ;
        RECT 410.800 346.200 411.600 351.800 ;
        RECT 412.400 351.600 413.200 352.400 ;
        RECT 417.200 351.600 418.000 352.400 ;
        RECT 418.800 351.600 419.600 352.400 ;
        RECT 417.300 350.400 417.900 351.600 ;
        RECT 412.400 349.600 413.200 350.400 ;
        RECT 415.600 349.600 416.400 350.400 ;
        RECT 417.200 349.600 418.000 350.400 ;
        RECT 417.200 347.600 418.000 348.400 ;
        RECT 418.900 340.400 419.500 351.600 ;
        RECT 418.800 339.600 419.600 340.400 ;
        RECT 407.600 337.600 408.400 338.400 ;
        RECT 407.700 332.600 408.300 337.600 ;
        RECT 402.800 331.600 403.600 332.400 ;
        RECT 407.600 331.800 408.400 332.600 ;
        RECT 409.200 326.200 410.000 337.800 ;
        RECT 410.800 333.600 411.600 334.400 ;
        RECT 394.800 323.600 395.600 324.400 ;
        RECT 394.900 322.400 395.500 323.600 ;
        RECT 394.800 321.600 395.600 322.400 ;
        RECT 404.400 313.600 405.200 314.400 ;
        RECT 396.400 309.600 397.200 310.400 ;
        RECT 393.200 307.600 394.000 308.400 ;
        RECT 396.400 307.600 397.200 308.400 ;
        RECT 401.200 307.600 402.000 308.400 ;
        RECT 396.500 306.400 397.100 307.600 ;
        RECT 396.400 305.600 397.200 306.400 ;
        RECT 402.800 306.300 403.600 306.400 ;
        RECT 401.300 305.700 403.600 306.300 ;
        RECT 391.600 303.600 392.400 304.400 ;
        RECT 394.800 303.600 395.600 304.400 ;
        RECT 398.000 303.600 398.800 304.400 ;
        RECT 377.200 301.600 378.000 302.400 ;
        RECT 369.200 293.600 370.000 294.400 ;
        RECT 372.400 286.200 373.200 297.800 ;
        RECT 374.000 291.600 374.800 292.400 ;
        RECT 329.200 283.600 330.000 284.400 ;
        RECT 348.400 283.600 349.200 284.400 ;
        RECT 330.800 271.600 331.600 272.400 ;
        RECT 321.200 269.600 322.000 270.400 ;
        RECT 324.400 269.600 325.200 270.400 ;
        RECT 327.600 269.600 328.400 270.400 ;
        RECT 311.600 267.600 312.400 268.400 ;
        RECT 318.000 267.600 318.800 268.400 ;
        RECT 319.600 267.600 320.400 268.400 ;
        RECT 311.700 266.400 312.300 267.600 ;
        RECT 311.600 265.600 312.400 266.400 ;
        RECT 273.200 263.600 274.000 264.400 ;
        RECT 287.600 263.600 288.400 264.400 ;
        RECT 310.000 263.600 310.800 264.400 ;
        RECT 263.600 251.600 264.400 252.400 ;
        RECT 266.800 246.200 267.600 257.800 ;
        RECT 273.300 256.400 273.900 263.600 ;
        RECT 319.700 258.400 320.300 267.600 ;
        RECT 321.200 265.600 322.000 266.400 ;
        RECT 324.500 262.400 325.100 269.600 ;
        RECT 326.000 267.600 326.800 268.400 ;
        RECT 329.200 267.600 330.000 268.400 ;
        RECT 324.400 261.600 325.200 262.400 ;
        RECT 273.200 255.600 274.000 256.400 ;
        RECT 268.400 251.600 269.200 252.400 ;
        RECT 274.800 251.800 275.600 252.600 ;
        RECT 274.900 250.400 275.500 251.800 ;
        RECT 274.800 249.600 275.600 250.400 ;
        RECT 276.400 246.200 277.200 257.800 ;
        RECT 289.200 257.600 290.000 258.400 ;
        RECT 279.600 250.200 280.400 255.800 ;
        RECT 281.200 253.600 282.000 254.400 ;
        RECT 289.300 252.400 289.900 257.600 ;
        RECT 289.200 251.600 290.000 252.400 ;
        RECT 295.600 246.200 296.400 257.800 ;
        RECT 297.200 251.600 298.000 252.400 ;
        RECT 303.600 251.600 304.400 252.600 ;
        RECT 305.200 246.200 306.000 257.800 ;
        RECT 319.600 257.600 320.400 258.400 ;
        RECT 308.400 250.200 309.200 255.800 ;
        RECT 311.400 255.000 312.200 255.800 ;
        RECT 313.200 255.000 317.400 255.600 ;
        RECT 318.000 255.000 318.800 255.800 ;
        RECT 319.600 255.600 320.400 256.400 ;
        RECT 310.000 253.600 310.800 254.400 ;
        RECT 311.400 250.200 312.000 255.000 ;
        RECT 313.200 254.800 314.000 255.000 ;
        RECT 316.600 254.800 317.400 255.000 ;
        RECT 318.200 254.200 318.800 255.000 ;
        RECT 319.700 254.400 320.300 255.600 ;
        RECT 324.500 254.400 325.100 261.600 ;
        RECT 326.100 256.400 326.700 267.600 ;
        RECT 329.300 266.400 329.900 267.600 ;
        RECT 329.200 265.600 330.000 266.400 ;
        RECT 329.200 261.600 330.000 262.400 ;
        RECT 330.900 262.300 331.500 271.600 ;
        RECT 334.000 269.600 334.800 270.400 ;
        RECT 334.000 267.600 334.800 268.400 ;
        RECT 338.800 267.600 339.600 268.400 ;
        RECT 342.000 267.600 342.800 268.400 ;
        RECT 334.000 265.600 334.800 266.400 ;
        RECT 340.400 265.600 341.200 266.400 ;
        RECT 332.400 263.600 333.200 264.400 ;
        RECT 330.900 261.700 333.100 262.300 ;
        RECT 329.300 258.400 329.900 261.600 ;
        RECT 327.600 257.600 328.400 258.400 ;
        RECT 329.200 257.600 330.000 258.400 ;
        RECT 330.800 257.600 331.600 258.400 ;
        RECT 326.000 255.600 326.800 256.400 ;
        RECT 327.700 254.400 328.300 257.600 ;
        RECT 330.900 254.400 331.500 257.600 ;
        RECT 332.500 254.400 333.100 261.700 ;
        RECT 314.000 253.600 318.800 254.200 ;
        RECT 319.600 253.600 320.400 254.400 ;
        RECT 321.200 253.600 322.000 254.400 ;
        RECT 324.400 253.600 325.200 254.400 ;
        RECT 327.600 253.600 328.400 254.400 ;
        RECT 330.800 253.600 331.600 254.400 ;
        RECT 332.400 253.600 333.200 254.400 ;
        RECT 314.000 253.400 314.800 253.600 ;
        RECT 311.400 249.400 312.200 250.200 ;
        RECT 313.200 249.600 314.000 250.400 ;
        RECT 318.200 250.200 318.800 253.600 ;
        RECT 332.500 252.400 333.100 253.600 ;
        RECT 334.100 252.400 334.700 265.600 ;
        RECT 342.100 264.400 342.700 267.600 ;
        RECT 345.200 265.600 346.000 266.400 ;
        RECT 342.000 263.600 342.800 264.400 ;
        RECT 345.300 258.400 345.900 265.600 ;
        RECT 346.800 264.200 347.600 275.800 ;
        RECT 348.500 274.400 349.100 283.600 ;
        RECT 348.400 273.600 349.200 274.400 ;
        RECT 354.800 271.600 355.600 272.400 ;
        RECT 354.900 270.200 355.500 271.600 ;
        RECT 354.800 269.400 355.600 270.200 ;
        RECT 351.600 267.600 352.400 268.400 ;
        RECT 340.400 257.600 341.200 258.400 ;
        RECT 345.200 257.600 346.000 258.400 ;
        RECT 340.500 256.400 341.100 257.600 ;
        RECT 340.400 255.600 341.200 256.400 ;
        RECT 350.000 256.300 350.800 256.400 ;
        RECT 348.500 255.700 350.800 256.300 ;
        RECT 348.500 254.400 349.100 255.700 ;
        RECT 350.000 255.600 350.800 255.700 ;
        RECT 343.600 253.600 344.400 254.400 ;
        RECT 348.400 253.600 349.200 254.400 ;
        RECT 350.000 253.600 350.800 254.400 ;
        RECT 343.700 252.400 344.300 253.600 ;
        RECT 322.800 251.600 323.600 252.400 ;
        RECT 324.400 251.600 325.200 252.400 ;
        RECT 332.400 251.600 333.200 252.400 ;
        RECT 334.000 251.600 334.800 252.400 ;
        RECT 337.200 251.600 338.000 252.400 ;
        RECT 343.600 251.600 344.400 252.400 ;
        RECT 313.300 248.400 313.900 249.600 ;
        RECT 318.000 249.400 318.800 250.200 ;
        RECT 321.200 249.600 322.000 250.400 ;
        RECT 322.900 250.300 323.500 251.600 ;
        RECT 324.400 250.300 325.200 250.400 ;
        RECT 322.900 249.700 325.200 250.300 ;
        RECT 324.400 249.600 325.200 249.700 ;
        RECT 334.000 249.600 334.800 250.400 ;
        RECT 345.200 249.600 346.000 250.400 ;
        RECT 313.200 247.600 314.000 248.400 ;
        RECT 258.800 233.600 259.600 234.400 ;
        RECT 263.600 226.200 264.400 231.800 ;
        RECT 265.200 227.600 266.000 228.400 ;
        RECT 262.000 223.600 262.800 224.400 ;
        RECT 174.100 217.700 176.300 218.300 ;
        RECT 174.000 215.600 174.800 216.400 ;
        RECT 170.800 211.600 171.600 212.400 ;
        RECT 156.400 189.600 157.200 190.400 ;
        RECT 159.600 184.200 160.400 195.800 ;
        RECT 166.000 186.200 166.800 191.800 ;
        RECT 164.400 184.300 165.200 184.400 ;
        RECT 162.900 183.700 165.200 184.300 ;
        RECT 169.200 184.200 170.000 195.800 ;
        RECT 170.900 188.400 171.500 211.600 ;
        RECT 172.400 203.600 173.200 204.400 ;
        RECT 170.800 187.600 171.600 188.400 ;
        RECT 172.500 186.400 173.100 203.600 ;
        RECT 175.700 190.400 176.300 217.700 ;
        RECT 180.400 217.600 181.200 218.400 ;
        RECT 191.700 216.400 192.300 223.600 ;
        RECT 204.400 217.600 205.200 218.400 ;
        RECT 188.400 215.600 189.200 216.400 ;
        RECT 191.600 215.600 192.400 216.400 ;
        RECT 177.200 213.600 178.000 214.400 ;
        RECT 182.000 213.600 182.800 214.400 ;
        RECT 183.600 213.600 184.400 214.400 ;
        RECT 183.700 212.400 184.300 213.600 ;
        RECT 191.700 212.400 192.300 215.600 ;
        RECT 193.200 213.600 194.000 214.400 ;
        RECT 196.400 213.600 197.200 214.400 ;
        RECT 183.600 211.600 184.400 212.400 ;
        RECT 188.400 211.600 189.200 212.400 ;
        RECT 191.600 211.600 192.400 212.400 ;
        RECT 193.200 211.600 194.000 212.400 ;
        RECT 186.800 209.600 187.600 210.400 ;
        RECT 180.400 203.600 181.200 204.400 ;
        RECT 175.600 189.600 176.400 190.400 ;
        RECT 172.400 185.600 173.200 186.400 ;
        RECT 178.800 184.200 179.600 195.800 ;
        RECT 180.500 190.400 181.100 203.600 ;
        RECT 186.900 196.400 187.500 209.600 ;
        RECT 188.500 208.400 189.100 211.600 ;
        RECT 193.300 208.400 193.900 211.600 ;
        RECT 196.500 210.400 197.100 213.600 ;
        RECT 198.000 211.600 198.800 212.400 ;
        RECT 196.400 209.600 197.200 210.400 ;
        RECT 201.200 209.600 202.000 210.400 ;
        RECT 202.800 210.200 203.600 215.800 ;
        RECT 204.500 214.400 205.100 217.600 ;
        RECT 204.400 213.600 205.200 214.400 ;
        RECT 201.300 208.400 201.900 209.600 ;
        RECT 188.400 207.600 189.200 208.400 ;
        RECT 193.200 207.600 194.000 208.400 ;
        RECT 201.200 207.600 202.000 208.400 ;
        RECT 186.800 195.600 187.600 196.400 ;
        RECT 190.000 195.600 190.800 196.400 ;
        RECT 188.400 191.600 189.200 192.400 ;
        RECT 180.400 189.600 181.200 190.400 ;
        RECT 185.200 185.600 186.000 186.400 ;
        RECT 153.200 181.600 154.000 182.400 ;
        RECT 124.400 173.600 125.200 174.400 ;
        RECT 132.400 171.600 133.200 172.400 ;
        RECT 127.600 169.600 128.400 170.400 ;
        RECT 134.000 170.200 134.800 175.800 ;
        RECT 137.200 166.200 138.000 177.800 ;
        RECT 145.200 173.600 146.000 174.400 ;
        RECT 138.800 171.800 139.600 172.600 ;
        RECT 145.300 172.400 145.900 173.600 ;
        RECT 138.900 166.400 139.500 171.800 ;
        RECT 145.200 171.600 146.000 172.400 ;
        RECT 138.800 165.600 139.600 166.400 ;
        RECT 146.800 166.200 147.600 177.800 ;
        RECT 153.200 170.200 154.000 175.800 ;
        RECT 154.800 173.600 155.600 174.400 ;
        RECT 156.400 166.200 157.200 177.800 ;
        RECT 158.000 171.600 158.800 172.600 ;
        RECT 122.800 163.600 123.600 164.400 ;
        RECT 151.600 163.600 152.400 164.400 ;
        RECT 122.900 158.400 123.500 163.600 ;
        RECT 122.800 157.600 123.600 158.400 ;
        RECT 142.000 153.600 142.800 154.400 ;
        RECT 122.800 149.600 123.600 150.400 ;
        RECT 126.000 149.600 126.800 150.400 ;
        RECT 129.200 149.600 130.000 150.400 ;
        RECT 135.600 149.600 136.400 150.400 ;
        RECT 121.200 147.600 122.000 148.400 ;
        RECT 113.200 146.200 114.000 147.000 ;
        RECT 114.600 146.400 118.800 147.000 ;
        RECT 116.500 134.400 117.100 146.400 ;
        RECT 119.800 146.200 120.600 147.000 ;
        RECT 121.200 145.600 122.000 146.400 ;
        RECT 121.300 138.400 121.900 145.600 ;
        RECT 122.900 144.400 123.500 149.600 ;
        RECT 122.800 143.600 123.600 144.400 ;
        RECT 118.000 137.600 118.800 138.400 ;
        RECT 121.200 137.600 122.000 138.400 ;
        RECT 114.800 134.300 115.600 134.400 ;
        RECT 113.300 133.700 115.600 134.300 ;
        RECT 113.300 132.400 113.900 133.700 ;
        RECT 114.800 133.600 115.600 133.700 ;
        RECT 116.400 133.600 117.200 134.400 ;
        RECT 113.200 131.600 114.000 132.400 ;
        RECT 114.800 131.600 115.600 132.400 ;
        RECT 97.200 129.600 98.000 130.400 ;
        RECT 105.200 129.600 106.000 130.400 ;
        RECT 111.600 129.600 112.400 130.400 ;
        RECT 97.300 128.400 97.900 129.600 ;
        RECT 89.200 127.600 90.000 128.400 ;
        RECT 97.200 127.600 98.000 128.400 ;
        RECT 87.600 123.600 88.400 124.400 ;
        RECT 102.000 123.600 102.800 124.400 ;
        RECT 102.100 120.400 102.700 123.600 ;
        RECT 105.300 122.400 105.900 129.600 ;
        RECT 105.200 121.600 106.000 122.400 ;
        RECT 102.000 119.600 102.800 120.400 ;
        RECT 108.400 115.600 109.200 116.400 ;
        RECT 108.500 112.400 109.100 115.600 ;
        RECT 92.400 111.600 93.200 112.400 ;
        RECT 97.200 111.600 98.000 112.400 ;
        RECT 108.400 111.600 109.200 112.400 ;
        RECT 111.600 111.600 112.400 112.400 ;
        RECT 97.300 110.400 97.900 111.600 ;
        RECT 111.700 110.400 112.300 111.600 ;
        RECT 89.200 109.600 90.000 110.400 ;
        RECT 97.200 109.600 98.000 110.400 ;
        RECT 98.800 109.600 99.600 110.400 ;
        RECT 105.200 109.600 106.000 110.400 ;
        RECT 108.400 109.600 109.200 110.400 ;
        RECT 111.600 109.600 112.400 110.400 ;
        RECT 87.600 107.600 88.400 108.400 ;
        RECT 89.200 107.600 90.000 108.400 ;
        RECT 103.600 107.600 104.400 108.400 ;
        RECT 106.800 107.600 107.600 108.400 ;
        RECT 86.000 101.600 86.800 102.400 ;
        RECT 87.700 98.400 88.300 107.600 ;
        RECT 89.300 106.400 89.900 107.600 ;
        RECT 89.200 105.600 90.000 106.400 ;
        RECT 94.000 105.600 94.800 106.400 ;
        RECT 98.800 105.600 99.600 106.400 ;
        RECT 102.000 105.600 102.800 106.400 ;
        RECT 90.800 103.600 91.600 104.400 ;
        RECT 100.400 103.600 101.200 104.400 ;
        RECT 105.200 103.600 106.000 104.400 ;
        RECT 87.600 97.600 88.400 98.400 ;
        RECT 84.400 95.600 85.200 96.400 ;
        RECT 84.500 94.400 85.100 95.600 ;
        RECT 90.900 94.400 91.500 103.600 ;
        RECT 100.500 98.400 101.100 103.600 ;
        RECT 105.300 98.400 105.900 103.600 ;
        RECT 100.400 97.600 101.200 98.400 ;
        RECT 105.200 97.600 106.000 98.400 ;
        RECT 106.900 96.400 107.500 107.600 ;
        RECT 108.500 96.400 109.100 109.600 ;
        RECT 110.000 107.600 110.800 108.400 ;
        RECT 110.100 106.400 110.700 107.600 ;
        RECT 110.000 105.600 110.800 106.400 ;
        RECT 94.000 95.600 94.800 96.400 ;
        RECT 98.800 95.600 99.600 96.400 ;
        RECT 100.400 95.600 101.200 96.400 ;
        RECT 106.800 95.600 107.600 96.400 ;
        RECT 108.400 95.600 109.200 96.400 ;
        RECT 84.400 93.600 85.200 94.400 ;
        RECT 89.200 93.600 90.000 94.400 ;
        RECT 90.800 93.600 91.600 94.400 ;
        RECT 97.200 93.600 98.000 94.400 ;
        RECT 98.900 92.400 99.500 95.600 ;
        RECT 108.500 92.400 109.100 95.600 ;
        RECT 110.000 94.300 110.800 94.400 ;
        RECT 111.700 94.300 112.300 109.600 ;
        RECT 110.000 93.700 112.300 94.300 ;
        RECT 110.000 93.600 110.800 93.700 ;
        RECT 95.600 91.600 96.400 92.400 ;
        RECT 98.800 91.600 99.600 92.400 ;
        RECT 102.000 91.600 102.800 92.400 ;
        RECT 108.400 91.600 109.200 92.400 ;
        RECT 84.400 89.600 85.200 90.400 ;
        RECT 66.800 75.600 67.600 76.400 ;
        RECT 76.400 75.600 77.200 76.400 ;
        RECT 82.800 75.600 83.600 76.400 ;
        RECT 66.900 72.400 67.500 75.600 ;
        RECT 73.200 73.600 74.000 74.400 ;
        RECT 44.400 71.600 45.200 72.400 ;
        RECT 63.600 71.600 64.400 72.400 ;
        RECT 66.800 71.600 67.600 72.400 ;
        RECT 74.800 71.600 75.600 72.400 ;
        RECT 44.500 70.400 45.100 71.600 ;
        RECT 31.600 70.300 32.400 70.400 ;
        RECT 30.100 69.700 32.400 70.300 ;
        RECT 31.600 69.600 32.400 69.700 ;
        RECT 41.200 69.600 42.000 70.400 ;
        RECT 42.800 69.600 43.600 70.400 ;
        RECT 44.400 69.600 45.200 70.400 ;
        RECT 50.800 69.600 51.600 70.400 ;
        RECT 55.600 69.600 56.400 70.400 ;
        RECT 62.000 69.600 62.800 70.400 ;
        RECT 42.900 68.400 43.500 69.600 ;
        RECT 33.200 67.600 34.000 68.400 ;
        RECT 36.400 67.600 37.200 68.400 ;
        RECT 42.800 67.600 43.600 68.400 ;
        RECT 46.000 67.600 46.800 68.400 ;
        RECT 31.600 65.600 32.400 66.400 ;
        RECT 31.700 64.400 32.300 65.600 ;
        RECT 26.800 63.600 27.600 64.400 ;
        RECT 31.600 63.600 32.400 64.400 ;
        RECT 25.200 57.600 26.000 58.400 ;
        RECT 10.800 53.600 11.600 54.400 ;
        RECT 12.400 53.600 13.200 54.400 ;
        RECT 20.400 53.600 21.200 54.400 ;
        RECT 23.600 53.600 24.400 54.400 ;
        RECT 9.200 51.600 10.000 52.400 ;
        RECT 9.300 50.400 9.900 51.600 ;
        RECT 9.200 49.600 10.000 50.400 ;
        RECT 10.900 36.300 11.500 53.600 ;
        RECT 9.300 35.700 11.500 36.300 ;
        RECT 7.600 31.600 8.400 32.400 ;
        RECT 9.300 30.300 9.900 35.700 ;
        RECT 10.800 33.600 11.600 34.400 ;
        RECT 12.500 32.400 13.100 53.600 ;
        RECT 25.300 52.400 25.900 57.600 ;
        RECT 14.000 51.600 14.800 52.400 ;
        RECT 18.800 51.600 19.600 52.400 ;
        RECT 20.400 51.600 21.200 52.400 ;
        RECT 25.200 51.600 26.000 52.400 ;
        RECT 14.100 50.400 14.700 51.600 ;
        RECT 18.900 50.400 19.500 51.600 ;
        RECT 14.000 49.600 14.800 50.400 ;
        RECT 18.800 49.600 19.600 50.400 ;
        RECT 23.600 49.600 24.400 50.400 ;
        RECT 17.200 43.600 18.000 44.400 ;
        RECT 12.400 31.600 13.200 32.400 ;
        RECT 17.300 30.400 17.900 43.600 ;
        RECT 26.900 34.400 27.500 63.600 ;
        RECT 30.000 57.600 30.800 58.400 ;
        RECT 30.100 54.400 30.700 57.600 ;
        RECT 30.000 53.600 30.800 54.400 ;
        RECT 31.700 52.400 32.300 63.600 ;
        RECT 33.300 60.400 33.900 67.600 ;
        RECT 38.000 65.600 38.800 66.400 ;
        RECT 38.100 64.400 38.700 65.600 ;
        RECT 34.800 63.600 35.600 64.400 ;
        RECT 38.000 63.600 38.800 64.400 ;
        RECT 33.200 59.600 34.000 60.400 ;
        RECT 33.300 56.400 33.900 59.600 ;
        RECT 33.200 55.600 34.000 56.400 ;
        RECT 34.900 54.400 35.500 63.600 ;
        RECT 42.800 61.600 43.600 62.400 ;
        RECT 41.200 57.600 42.000 58.400 ;
        RECT 36.400 55.600 37.200 56.400 ;
        RECT 38.000 55.600 38.800 56.400 ;
        RECT 36.500 54.400 37.100 55.600 ;
        RECT 34.800 53.600 35.600 54.400 ;
        RECT 36.400 53.600 37.200 54.400 ;
        RECT 28.400 51.600 29.200 52.400 ;
        RECT 31.600 51.600 32.400 52.400 ;
        RECT 34.900 50.400 35.500 53.600 ;
        RECT 38.100 52.400 38.700 55.600 ;
        RECT 41.300 54.400 41.900 57.600 ;
        RECT 41.200 53.600 42.000 54.400 ;
        RECT 42.900 52.400 43.500 61.600 ;
        RECT 38.000 51.600 38.800 52.400 ;
        RECT 39.600 51.600 40.400 52.400 ;
        RECT 42.800 51.600 43.600 52.400 ;
        RECT 34.800 49.600 35.600 50.400 ;
        RECT 46.100 48.400 46.700 67.600 ;
        RECT 50.800 65.600 51.600 66.400 ;
        RECT 50.900 64.400 51.500 65.600 ;
        RECT 50.800 63.600 51.600 64.400 ;
        RECT 55.700 62.400 56.300 69.600 ;
        RECT 57.200 67.600 58.000 68.400 ;
        RECT 60.400 67.600 61.200 68.400 ;
        RECT 62.000 67.600 62.800 68.400 ;
        RECT 55.600 61.600 56.400 62.400 ;
        RECT 57.300 56.400 57.900 67.600 ;
        RECT 60.500 56.400 61.100 67.600 ;
        RECT 63.700 64.400 64.300 71.600 ;
        RECT 74.900 68.400 75.500 71.600 ;
        RECT 76.500 68.400 77.100 75.600 ;
        RECT 79.600 73.600 80.400 74.400 ;
        RECT 82.800 73.600 83.600 74.400 ;
        RECT 79.700 70.400 80.300 73.600 ;
        RECT 102.100 72.400 102.700 91.600 ;
        RECT 103.600 79.600 104.400 80.400 ;
        RECT 97.200 71.600 98.000 72.400 ;
        RECT 102.000 71.600 102.800 72.400 ;
        RECT 79.600 69.600 80.400 70.400 ;
        RECT 97.300 68.400 97.900 71.600 ;
        RECT 103.700 68.400 104.300 79.600 ;
        RECT 113.300 74.400 113.900 131.600 ;
        RECT 114.900 124.400 115.500 131.600 ;
        RECT 118.100 128.400 118.700 137.600 ;
        RECT 119.600 129.600 120.400 130.400 ;
        RECT 118.000 127.600 118.800 128.400 ;
        RECT 114.800 123.600 115.600 124.400 ;
        RECT 118.100 118.400 118.700 127.600 ;
        RECT 114.800 117.600 115.600 118.400 ;
        RECT 118.000 117.600 118.800 118.400 ;
        RECT 114.900 112.400 115.500 117.600 ;
        RECT 114.800 111.600 115.600 112.400 ;
        RECT 121.200 111.600 122.000 112.400 ;
        RECT 116.400 109.600 117.200 110.400 ;
        RECT 114.800 99.600 115.600 100.400 ;
        RECT 114.900 96.400 115.500 99.600 ;
        RECT 114.800 95.600 115.600 96.400 ;
        RECT 114.800 87.600 115.600 88.400 ;
        RECT 113.200 73.600 114.000 74.400 ;
        RECT 105.200 71.600 106.000 72.400 ;
        RECT 108.400 71.600 109.200 72.400 ;
        RECT 105.200 69.600 106.000 70.400 ;
        RECT 74.800 67.600 75.600 68.400 ;
        RECT 76.400 67.600 77.200 68.400 ;
        RECT 86.000 67.600 86.800 68.400 ;
        RECT 92.400 67.600 93.200 68.400 ;
        RECT 94.000 67.600 94.800 68.400 ;
        RECT 97.200 67.600 98.000 68.400 ;
        RECT 98.800 67.600 99.600 68.400 ;
        RECT 103.600 67.600 104.400 68.400 ;
        RECT 63.600 63.600 64.400 64.400 ;
        RECT 70.000 63.600 70.800 64.400 ;
        RECT 63.700 56.400 64.300 63.600 ;
        RECT 54.000 55.600 54.800 56.400 ;
        RECT 57.200 55.600 58.000 56.400 ;
        RECT 60.400 55.600 61.200 56.400 ;
        RECT 62.000 55.600 62.800 56.400 ;
        RECT 63.600 55.600 64.400 56.400 ;
        RECT 66.800 55.600 67.600 56.400 ;
        RECT 50.800 54.300 51.600 54.400 ;
        RECT 47.700 53.700 51.600 54.300 ;
        RECT 47.700 52.400 48.300 53.700 ;
        RECT 50.800 53.600 51.600 53.700 ;
        RECT 54.100 52.400 54.700 55.600 ;
        RECT 66.900 54.400 67.500 55.600 ;
        RECT 66.800 53.600 67.600 54.400 ;
        RECT 47.600 51.600 48.400 52.400 ;
        RECT 54.000 51.600 54.800 52.400 ;
        RECT 68.400 51.600 69.200 52.400 ;
        RECT 49.200 49.600 50.000 50.400 ;
        RECT 50.800 49.600 51.600 50.400 ;
        RECT 55.600 49.600 56.400 50.400 ;
        RECT 42.800 47.600 43.600 48.400 ;
        RECT 46.000 47.600 46.800 48.400 ;
        RECT 30.000 35.600 30.800 36.400 ;
        RECT 20.400 33.600 21.200 34.400 ;
        RECT 26.800 33.600 27.600 34.400 ;
        RECT 20.500 32.400 21.100 33.600 ;
        RECT 20.400 31.600 21.200 32.400 ;
        RECT 30.100 30.400 30.700 35.600 ;
        RECT 42.900 34.400 43.500 47.600 ;
        RECT 44.400 43.600 45.200 44.400 ;
        RECT 42.800 33.600 43.600 34.400 ;
        RECT 36.400 31.600 37.200 32.400 ;
        RECT 39.600 31.600 40.400 32.400 ;
        RECT 39.700 30.400 40.300 31.600 ;
        RECT 42.900 30.400 43.500 33.600 ;
        RECT 44.500 30.400 45.100 43.600 ;
        RECT 50.900 38.400 51.500 49.600 ;
        RECT 55.700 38.400 56.300 49.600 ;
        RECT 58.800 43.600 59.600 44.400 ;
        RECT 63.600 43.600 64.400 44.400 ;
        RECT 50.800 37.600 51.600 38.400 ;
        RECT 55.600 37.600 56.400 38.400 ;
        RECT 52.400 33.600 53.200 34.400 ;
        RECT 52.500 30.400 53.100 33.600 ;
        RECT 7.700 29.700 9.900 30.300 ;
        RECT 6.000 23.600 6.800 24.400 ;
        RECT 1.200 19.600 2.000 20.400 ;
        RECT 4.400 19.600 5.200 20.400 ;
        RECT 1.300 16.400 1.900 19.600 ;
        RECT 1.200 15.600 2.000 16.400 ;
        RECT 2.800 13.600 3.600 14.400 ;
        RECT 6.100 8.400 6.700 23.600 ;
        RECT 7.700 12.400 8.300 29.700 ;
        RECT 14.000 29.600 14.800 30.400 ;
        RECT 17.200 29.600 18.000 30.400 ;
        RECT 18.800 29.600 19.600 30.400 ;
        RECT 23.600 29.600 24.400 30.400 ;
        RECT 30.000 29.600 30.800 30.400 ;
        RECT 31.600 29.600 32.400 30.400 ;
        RECT 39.600 29.600 40.400 30.400 ;
        RECT 42.800 29.600 43.600 30.400 ;
        RECT 44.400 29.600 45.200 30.400 ;
        RECT 49.200 29.600 50.000 30.400 ;
        RECT 52.400 29.600 53.200 30.400 ;
        RECT 9.200 27.600 10.000 28.400 ;
        RECT 7.600 11.600 8.400 12.400 ;
        RECT 9.300 10.400 9.900 27.600 ;
        RECT 14.100 26.400 14.700 29.600 ;
        RECT 31.700 28.400 32.300 29.600 ;
        RECT 17.200 27.600 18.000 28.400 ;
        RECT 25.200 27.600 26.000 28.400 ;
        RECT 31.600 27.600 32.400 28.400 ;
        RECT 41.200 27.600 42.000 28.400 ;
        RECT 44.400 27.600 45.200 28.400 ;
        RECT 17.300 26.400 17.900 27.600 ;
        RECT 41.300 26.400 41.900 27.600 ;
        RECT 49.300 26.400 49.900 29.600 ;
        RECT 58.900 28.400 59.500 43.600 ;
        RECT 60.400 31.800 61.200 32.600 ;
        RECT 63.700 32.400 64.300 43.600 ;
        RECT 68.400 37.600 69.200 38.400 ;
        RECT 60.400 28.400 61.000 31.800 ;
        RECT 63.600 31.600 64.400 32.400 ;
        RECT 67.000 31.800 67.800 32.600 ;
        RECT 64.400 28.400 65.200 28.600 ;
        RECT 58.800 27.600 59.600 28.400 ;
        RECT 60.400 27.800 65.200 28.400 ;
        RECT 60.400 27.000 61.000 27.800 ;
        RECT 61.800 27.000 62.600 27.200 ;
        RECT 65.200 27.000 66.000 27.200 ;
        RECT 67.200 27.000 67.800 31.800 ;
        RECT 68.500 28.400 69.100 37.600 ;
        RECT 70.100 34.400 70.700 63.600 ;
        RECT 74.900 52.400 75.500 67.600 ;
        RECT 76.500 66.400 77.100 67.600 ;
        RECT 86.100 66.400 86.700 67.600 ;
        RECT 92.500 66.400 93.100 67.600 ;
        RECT 94.100 66.400 94.700 67.600 ;
        RECT 76.400 65.600 77.200 66.400 ;
        RECT 86.000 65.600 86.800 66.400 ;
        RECT 92.400 65.600 93.200 66.400 ;
        RECT 94.000 65.600 94.800 66.400 ;
        RECT 97.300 66.300 97.900 67.600 ;
        RECT 103.700 66.400 104.300 67.600 ;
        RECT 97.300 65.700 99.500 66.300 ;
        RECT 78.000 63.600 78.800 64.400 ;
        RECT 89.200 63.600 90.000 64.400 ;
        RECT 97.200 63.600 98.000 64.400 ;
        RECT 78.100 56.400 78.700 63.600 ;
        RECT 79.600 61.600 80.400 62.400 ;
        RECT 78.000 55.600 78.800 56.400 ;
        RECT 79.700 54.400 80.300 61.600 ;
        RECT 86.000 57.600 86.800 58.400 ;
        RECT 81.200 55.600 82.000 56.400 ;
        RECT 86.000 55.600 86.800 56.400 ;
        RECT 89.300 56.300 89.900 63.600 ;
        RECT 97.300 58.400 97.900 63.600 ;
        RECT 97.200 57.600 98.000 58.400 ;
        RECT 89.300 55.700 91.500 56.300 ;
        RECT 79.600 53.600 80.400 54.400 ;
        RECT 81.300 52.400 81.900 55.600 ;
        RECT 74.800 51.600 75.600 52.400 ;
        RECT 76.400 51.600 77.200 52.400 ;
        RECT 78.000 51.600 78.800 52.400 ;
        RECT 81.200 51.600 82.000 52.400 ;
        RECT 76.500 48.400 77.100 51.600 ;
        RECT 86.100 50.400 86.700 55.600 ;
        RECT 89.200 53.600 90.000 54.400 ;
        RECT 90.900 52.400 91.500 55.700 ;
        RECT 98.900 54.400 99.500 65.700 ;
        RECT 103.600 65.600 104.400 66.400 ;
        RECT 105.300 64.400 105.900 69.600 ;
        RECT 106.800 65.600 107.600 66.400 ;
        RECT 100.400 63.600 101.200 64.400 ;
        RECT 105.200 63.600 106.000 64.400 ;
        RECT 95.600 53.600 96.400 54.400 ;
        RECT 98.800 53.600 99.600 54.400 ;
        RECT 90.800 51.600 91.600 52.400 ;
        RECT 90.900 50.400 91.500 51.600 ;
        RECT 95.700 50.400 96.300 53.600 ;
        RECT 84.400 49.600 85.200 50.400 ;
        RECT 86.000 49.600 86.800 50.400 ;
        RECT 90.800 49.600 91.600 50.400 ;
        RECT 95.600 49.600 96.400 50.400 ;
        RECT 100.500 48.400 101.100 63.600 ;
        RECT 106.900 56.400 107.500 65.600 ;
        RECT 108.500 62.400 109.100 71.600 ;
        RECT 116.500 70.400 117.100 109.600 ;
        RECT 122.900 106.400 123.500 143.600 ;
        RECT 126.100 134.400 126.700 149.600 ;
        RECT 127.600 145.600 128.400 146.400 ;
        RECT 127.700 142.400 128.300 145.600 ;
        RECT 127.600 141.600 128.400 142.400 ;
        RECT 129.300 138.400 129.900 149.600 ;
        RECT 134.000 147.600 134.800 148.400 ;
        RECT 134.000 145.600 134.800 146.400 ;
        RECT 135.700 142.400 136.300 149.600 ;
        RECT 142.100 148.400 142.700 153.600 ;
        RECT 143.600 151.800 144.400 152.600 ;
        RECT 150.200 151.800 151.000 152.600 ;
        RECT 143.600 148.400 144.200 151.800 ;
        RECT 147.600 148.400 148.400 148.600 ;
        RECT 142.000 147.600 142.800 148.400 ;
        RECT 143.600 147.800 148.400 148.400 ;
        RECT 143.600 147.000 144.200 147.800 ;
        RECT 145.000 147.000 145.800 147.200 ;
        RECT 148.400 147.000 149.200 147.200 ;
        RECT 150.400 147.000 151.000 151.800 ;
        RECT 143.600 146.200 144.400 147.000 ;
        RECT 145.000 146.400 149.200 147.000 ;
        RECT 146.800 145.600 147.600 146.400 ;
        RECT 150.200 146.200 151.000 147.000 ;
        RECT 151.700 146.400 152.300 163.600 ;
        RECT 151.600 145.600 152.400 146.400 ;
        RECT 153.200 146.200 154.000 151.800 ;
        RECT 148.400 143.600 149.200 144.400 ;
        RECT 156.400 144.200 157.200 155.800 ;
        RECT 158.000 151.600 158.800 152.400 ;
        RECT 158.100 150.200 158.700 151.600 ;
        RECT 158.000 149.400 158.800 150.200 ;
        RECT 162.900 144.400 163.500 183.700 ;
        RECT 164.400 183.600 165.200 183.700 ;
        RECT 183.600 183.600 184.400 184.400 ;
        RECT 185.300 182.400 185.900 185.600 ;
        RECT 186.800 183.600 187.600 184.400 ;
        RECT 172.400 181.600 173.200 182.400 ;
        RECT 185.200 181.600 186.000 182.400 ;
        RECT 164.400 171.600 165.200 172.400 ;
        RECT 164.500 150.400 165.100 171.600 ;
        RECT 166.000 166.200 166.800 177.800 ;
        RECT 172.500 174.400 173.100 181.600 ;
        RECT 186.900 178.400 187.500 183.600 ;
        RECT 186.800 177.600 187.600 178.400 ;
        RECT 174.000 175.000 174.800 175.800 ;
        RECT 175.400 175.000 179.600 175.600 ;
        RECT 180.600 175.000 181.400 175.800 ;
        RECT 185.200 175.600 186.000 176.400 ;
        RECT 172.400 173.600 173.200 174.400 ;
        RECT 174.000 174.200 174.600 175.000 ;
        RECT 175.400 174.800 176.200 175.000 ;
        RECT 178.800 174.800 179.600 175.000 ;
        RECT 174.000 173.600 178.800 174.200 ;
        RECT 174.000 170.200 174.600 173.600 ;
        RECT 178.000 173.400 178.800 173.600 ;
        RECT 180.800 170.200 181.400 175.000 ;
        RECT 182.000 173.600 182.800 174.400 ;
        RECT 183.600 173.600 184.400 174.400 ;
        RECT 182.100 172.400 182.700 173.600 ;
        RECT 182.000 171.600 182.800 172.400 ;
        RECT 174.000 169.400 174.800 170.200 ;
        RECT 180.600 169.400 181.400 170.200 ;
        RECT 178.800 165.600 179.600 166.400 ;
        RECT 170.800 163.600 171.600 164.400 ;
        RECT 170.900 162.400 171.500 163.600 ;
        RECT 170.800 161.600 171.600 162.400 ;
        RECT 164.400 149.600 165.200 150.400 ;
        RECT 158.000 143.600 158.800 144.400 ;
        RECT 162.800 143.600 163.600 144.400 ;
        RECT 135.600 141.600 136.400 142.400 ;
        RECT 129.200 137.600 130.000 138.400 ;
        RECT 148.500 136.400 149.100 143.600 ;
        RECT 138.800 135.000 139.600 135.800 ;
        RECT 140.200 135.000 144.400 135.600 ;
        RECT 145.400 135.000 146.200 135.800 ;
        RECT 146.800 135.600 147.600 136.400 ;
        RECT 148.400 135.600 149.200 136.400 ;
        RECT 126.000 133.600 126.800 134.400 ;
        RECT 130.800 133.600 131.600 134.400 ;
        RECT 138.800 134.200 139.400 135.000 ;
        RECT 140.200 134.800 141.000 135.000 ;
        RECT 143.600 134.800 144.400 135.000 ;
        RECT 138.800 133.600 143.600 134.200 ;
        RECT 126.000 131.600 126.800 132.400 ;
        RECT 122.800 105.600 123.600 106.400 ;
        RECT 124.400 103.600 125.200 104.400 ;
        RECT 124.500 100.400 125.100 103.600 ;
        RECT 124.400 99.600 125.200 100.400 ;
        RECT 126.100 98.400 126.700 131.600 ;
        RECT 127.600 129.600 128.400 130.400 ;
        RECT 138.800 130.200 139.400 133.600 ;
        RECT 142.800 133.400 143.600 133.600 ;
        RECT 145.600 130.200 146.200 135.000 ;
        RECT 146.900 134.400 147.500 135.600 ;
        RECT 149.800 135.000 150.600 135.800 ;
        RECT 151.600 135.000 155.800 135.600 ;
        RECT 156.400 135.000 157.200 135.800 ;
        RECT 146.800 133.600 147.600 134.400 ;
        RECT 148.400 133.600 149.200 134.400 ;
        RECT 148.500 130.400 149.100 133.600 ;
        RECT 127.700 128.400 128.300 129.600 ;
        RECT 138.800 129.400 139.600 130.200 ;
        RECT 145.400 129.400 146.200 130.200 ;
        RECT 148.400 129.600 149.200 130.400 ;
        RECT 149.800 130.200 150.400 135.000 ;
        RECT 151.600 134.800 152.400 135.000 ;
        RECT 155.000 134.800 155.800 135.000 ;
        RECT 156.600 134.200 157.200 135.000 ;
        RECT 158.100 134.400 158.700 143.600 ;
        RECT 152.400 133.600 157.200 134.200 ;
        RECT 158.000 133.600 158.800 134.400 ;
        RECT 152.400 133.400 153.200 133.600 ;
        RECT 156.600 130.200 157.200 133.600 ;
        RECT 127.600 127.600 128.400 128.400 ;
        RECT 142.000 123.600 142.800 124.400 ;
        RECT 130.800 117.600 131.600 118.400 ;
        RECT 130.900 110.400 131.500 117.600 ;
        RECT 137.200 115.600 138.000 116.400 ;
        RECT 134.000 111.600 134.800 112.400 ;
        RECT 134.100 110.400 134.700 111.600 ;
        RECT 127.600 109.600 128.400 110.400 ;
        RECT 130.800 109.600 131.600 110.400 ;
        RECT 134.000 109.600 134.800 110.400 ;
        RECT 127.600 107.600 128.400 108.400 ;
        RECT 127.700 106.400 128.300 107.600 ;
        RECT 127.600 105.600 128.400 106.400 ;
        RECT 119.700 97.700 123.500 98.300 ;
        RECT 119.700 94.400 120.300 97.700 ;
        RECT 121.200 95.600 122.000 96.400 ;
        RECT 122.900 96.300 123.500 97.700 ;
        RECT 126.000 97.600 126.800 98.400 ;
        RECT 124.400 96.300 125.200 96.400 ;
        RECT 122.900 95.700 125.200 96.300 ;
        RECT 124.400 95.600 125.200 95.700 ;
        RECT 119.600 93.600 120.400 94.400 ;
        RECT 121.300 92.400 121.900 95.600 ;
        RECT 122.800 93.600 123.600 94.400 ;
        RECT 121.200 91.600 122.000 92.400 ;
        RECT 124.400 91.600 125.200 92.400 ;
        RECT 121.200 85.600 122.000 86.400 ;
        RECT 121.300 82.400 121.900 85.600 ;
        RECT 121.200 81.600 122.000 82.400 ;
        RECT 110.000 69.600 110.800 70.400 ;
        RECT 116.400 69.600 117.200 70.400 ;
        RECT 119.600 69.600 120.400 70.400 ;
        RECT 110.100 64.400 110.700 69.600 ;
        RECT 118.000 67.600 118.800 68.400 ;
        RECT 113.200 65.600 114.000 66.400 ;
        RECT 110.000 63.600 110.800 64.400 ;
        RECT 118.100 62.400 118.700 67.600 ;
        RECT 119.700 62.400 120.300 69.600 ;
        RECT 121.300 68.400 121.900 81.600 ;
        RECT 122.800 69.600 123.600 70.400 ;
        RECT 121.200 67.600 122.000 68.400 ;
        RECT 121.200 63.600 122.000 64.400 ;
        RECT 122.800 63.600 123.600 64.400 ;
        RECT 108.400 61.600 109.200 62.400 ;
        RECT 113.200 61.600 114.000 62.400 ;
        RECT 114.800 61.600 115.600 62.400 ;
        RECT 118.000 61.600 118.800 62.400 ;
        RECT 119.600 61.600 120.400 62.400 ;
        RECT 106.800 55.600 107.600 56.400 ;
        RECT 110.000 55.600 110.800 56.400 ;
        RECT 110.100 54.400 110.700 55.600 ;
        RECT 113.300 54.400 113.900 61.600 ;
        RECT 102.000 53.600 102.800 54.400 ;
        RECT 110.000 53.600 110.800 54.400 ;
        RECT 111.600 53.600 112.400 54.400 ;
        RECT 113.200 53.600 114.000 54.400 ;
        RECT 102.100 52.400 102.700 53.600 ;
        RECT 111.700 52.400 112.300 53.600 ;
        RECT 114.900 52.400 115.500 61.600 ;
        RECT 121.300 58.400 121.900 63.600 ;
        RECT 121.200 57.600 122.000 58.400 ;
        RECT 122.900 56.400 123.500 63.600 ;
        RECT 116.400 55.600 117.200 56.400 ;
        RECT 122.800 55.600 123.600 56.400 ;
        RECT 122.900 54.400 123.500 55.600 ;
        RECT 122.800 53.600 123.600 54.400 ;
        RECT 102.000 51.600 102.800 52.400 ;
        RECT 111.600 51.600 112.400 52.400 ;
        RECT 114.800 51.600 115.600 52.400 ;
        RECT 118.000 51.600 118.800 52.400 ;
        RECT 124.500 52.300 125.100 91.600 ;
        RECT 126.000 72.300 126.800 72.400 ;
        RECT 127.700 72.300 128.300 105.600 ;
        RECT 130.900 96.400 131.500 109.600 ;
        RECT 135.600 105.600 136.400 106.400 ;
        RECT 134.000 97.600 134.800 98.400 ;
        RECT 130.800 95.600 131.600 96.400 ;
        RECT 134.100 92.400 134.700 97.600 ;
        RECT 140.400 93.600 141.200 94.400 ;
        RECT 129.200 91.600 130.000 92.400 ;
        RECT 134.000 91.600 134.800 92.400 ;
        RECT 126.000 71.700 128.300 72.300 ;
        RECT 126.000 71.600 126.800 71.700 ;
        RECT 129.300 60.400 129.900 91.600 ;
        RECT 140.500 90.400 141.100 93.600 ;
        RECT 140.400 89.600 141.200 90.400 ;
        RECT 130.800 73.600 131.600 74.400 ;
        RECT 137.200 73.600 138.000 74.400 ;
        RECT 130.900 68.400 131.500 73.600 ;
        RECT 137.300 68.400 137.900 73.600 ;
        RECT 142.100 70.400 142.700 123.600 ;
        RECT 148.500 112.300 149.100 129.600 ;
        RECT 149.800 129.400 150.600 130.200 ;
        RECT 156.400 129.400 157.200 130.200 ;
        RECT 158.100 128.300 158.700 133.600 ;
        RECT 159.600 130.200 160.400 135.800 ;
        RECT 158.100 127.700 160.300 128.300 ;
        RECT 151.600 123.600 152.400 124.400 ;
        RECT 151.700 118.400 152.300 123.600 ;
        RECT 151.600 117.600 152.400 118.400 ;
        RECT 148.500 111.700 150.700 112.300 ;
        RECT 148.400 109.600 149.200 110.400 ;
        RECT 150.100 108.400 150.700 111.700 ;
        RECT 151.800 111.800 152.600 112.600 ;
        RECT 158.000 111.800 158.800 112.600 ;
        RECT 150.000 107.600 150.800 108.400 ;
        RECT 150.100 106.400 150.700 107.600 ;
        RECT 151.800 107.000 152.400 111.800 ;
        RECT 153.000 109.800 153.800 110.600 ;
        RECT 153.200 108.400 153.800 109.800 ;
        RECT 156.400 109.600 157.200 110.400 ;
        RECT 158.200 108.400 158.800 111.800 ;
        RECT 159.700 108.400 160.300 127.700 ;
        RECT 162.800 126.200 163.600 137.800 ;
        RECT 164.500 136.400 165.100 149.600 ;
        RECT 166.000 144.200 166.800 155.800 ;
        RECT 172.400 149.600 173.200 150.400 ;
        RECT 170.800 143.600 171.600 144.400 ;
        RECT 164.400 135.600 165.200 136.400 ;
        RECT 164.400 131.600 165.200 132.600 ;
        RECT 170.900 132.400 171.500 143.600 ;
        RECT 183.700 142.400 184.300 173.600 ;
        RECT 185.300 172.400 185.900 175.600 ;
        RECT 185.200 171.600 186.000 172.400 ;
        RECT 186.800 171.600 187.600 172.400 ;
        RECT 188.500 156.400 189.100 191.600 ;
        RECT 190.100 174.400 190.700 195.600 ;
        RECT 191.600 191.600 192.400 192.400 ;
        RECT 191.600 189.600 192.400 190.400 ;
        RECT 193.300 188.400 193.900 207.600 ;
        RECT 198.000 203.600 198.800 204.400 ;
        RECT 198.100 196.400 198.700 203.600 ;
        RECT 198.000 195.600 198.800 196.400 ;
        RECT 199.600 191.600 200.400 192.400 ;
        RECT 201.300 190.300 201.900 207.600 ;
        RECT 206.000 206.200 206.800 217.800 ;
        RECT 207.600 213.600 208.400 214.400 ;
        RECT 207.700 212.600 208.300 213.600 ;
        RECT 207.600 211.800 208.400 212.600 ;
        RECT 215.600 206.200 216.400 217.800 ;
        RECT 217.300 212.400 217.900 223.600 ;
        RECT 220.400 217.600 221.200 218.400 ;
        RECT 225.200 217.600 226.000 218.400 ;
        RECT 225.300 216.400 225.900 217.600 ;
        RECT 225.200 215.600 226.000 216.400 ;
        RECT 230.000 213.600 230.800 214.400 ;
        RECT 234.800 213.600 235.600 214.400 ;
        RECT 217.200 211.600 218.000 212.400 ;
        RECT 222.000 211.600 222.800 212.400 ;
        RECT 226.800 211.600 227.600 212.400 ;
        RECT 236.400 212.300 237.200 212.400 ;
        RECT 238.100 212.300 238.700 223.600 ;
        RECT 241.200 213.600 242.000 214.400 ;
        RECT 246.000 213.600 246.800 214.400 ;
        RECT 247.600 213.600 248.400 214.400 ;
        RECT 241.300 212.400 241.900 213.600 ;
        RECT 247.700 212.400 248.300 213.600 ;
        RECT 236.400 211.700 238.700 212.300 ;
        RECT 236.400 211.600 237.200 211.700 ;
        RECT 241.200 211.600 242.000 212.400 ;
        RECT 242.800 211.600 243.600 212.400 ;
        RECT 247.600 211.600 248.400 212.400 ;
        RECT 249.200 211.600 250.000 212.400 ;
        RECT 233.200 209.600 234.000 210.400 ;
        RECT 239.600 209.600 240.400 210.400 ;
        RECT 233.300 208.400 233.900 209.600 ;
        RECT 217.200 207.600 218.000 208.400 ;
        RECT 233.200 207.600 234.000 208.400 ;
        RECT 202.800 193.600 203.600 194.400 ;
        RECT 206.000 191.600 206.800 192.400 ;
        RECT 215.600 191.800 216.400 192.600 ;
        RECT 217.300 192.400 217.900 207.600 ;
        RECT 239.700 206.400 240.300 209.600 ;
        RECT 239.600 205.600 240.400 206.400 ;
        RECT 223.600 195.600 224.400 196.400 ;
        RECT 202.800 190.300 203.600 190.400 ;
        RECT 201.300 189.700 203.600 190.300 ;
        RECT 202.800 189.600 203.600 189.700 ;
        RECT 193.200 187.600 194.000 188.400 ;
        RECT 198.000 187.600 198.800 188.400 ;
        RECT 204.400 188.300 205.200 188.400 ;
        RECT 206.100 188.300 206.700 191.600 ;
        RECT 204.400 187.700 206.700 188.300 ;
        RECT 215.600 188.400 216.200 191.800 ;
        RECT 217.200 191.600 218.000 192.400 ;
        RECT 222.200 191.800 223.000 192.600 ;
        RECT 217.200 189.600 218.000 190.400 ;
        RECT 219.600 188.400 220.400 188.600 ;
        RECT 215.600 187.800 220.400 188.400 ;
        RECT 204.400 187.600 205.200 187.700 ;
        RECT 198.100 186.400 198.700 187.600 ;
        RECT 215.600 187.000 216.200 187.800 ;
        RECT 217.000 187.000 217.800 187.200 ;
        RECT 220.400 187.000 221.200 187.200 ;
        RECT 222.400 187.000 223.000 191.800 ;
        RECT 223.700 188.400 224.300 195.600 ;
        RECT 223.600 187.600 224.400 188.400 ;
        RECT 198.000 185.600 198.800 186.400 ;
        RECT 212.400 185.600 213.200 186.400 ;
        RECT 215.600 186.200 216.400 187.000 ;
        RECT 217.000 186.400 221.200 187.000 ;
        RECT 222.200 186.200 223.000 187.000 ;
        RECT 225.200 186.200 226.000 191.800 ;
        RECT 226.800 191.600 227.600 192.400 ;
        RECT 226.900 188.400 227.500 191.600 ;
        RECT 226.800 187.600 227.600 188.400 ;
        RECT 196.400 183.600 197.200 184.400 ;
        RECT 207.600 183.600 208.400 184.400 ;
        RECT 210.800 183.600 211.600 184.400 ;
        RECT 228.400 184.200 229.200 195.800 ;
        RECT 230.000 193.600 230.800 194.400 ;
        RECT 230.100 190.200 230.700 193.600 ;
        RECT 230.000 189.400 230.800 190.200 ;
        RECT 234.800 187.600 235.600 188.400 ;
        RECT 193.200 177.600 194.000 178.400 ;
        RECT 193.300 174.400 193.900 177.600 ;
        RECT 190.000 173.600 190.800 174.400 ;
        RECT 193.200 173.600 194.000 174.400 ;
        RECT 196.500 172.400 197.100 183.600 ;
        RECT 204.400 177.600 205.200 178.400 ;
        RECT 207.700 178.300 208.300 183.600 ;
        RECT 207.700 177.700 209.900 178.300 ;
        RECT 201.200 175.600 202.000 176.400 ;
        RECT 201.300 174.400 201.900 175.600 ;
        RECT 204.500 174.400 205.100 177.600 ;
        RECT 209.300 176.400 209.900 177.700 ;
        RECT 210.900 176.400 211.500 183.600 ;
        RECT 207.600 175.600 208.400 176.400 ;
        RECT 209.200 175.600 210.000 176.400 ;
        RECT 210.800 175.600 211.600 176.400 ;
        RECT 217.200 175.600 218.000 176.400 ;
        RECT 210.900 174.400 211.500 175.600 ;
        RECT 199.600 173.600 200.400 174.400 ;
        RECT 201.200 173.600 202.000 174.400 ;
        RECT 204.400 173.600 205.200 174.400 ;
        RECT 210.800 173.600 211.600 174.400 ;
        RECT 196.400 171.600 197.200 172.400 ;
        RECT 198.000 171.600 198.800 172.400 ;
        RECT 198.100 170.400 198.700 171.600 ;
        RECT 199.700 170.400 200.300 173.600 ;
        RECT 202.800 171.600 203.600 172.400 ;
        RECT 212.400 171.600 213.200 172.400 ;
        RECT 215.600 171.600 216.400 172.400 ;
        RECT 217.300 170.400 217.900 175.600 ;
        RECT 222.000 173.600 222.800 174.400 ;
        RECT 223.600 173.600 224.400 174.400 ;
        RECT 220.400 171.600 221.200 172.400 ;
        RECT 223.700 170.400 224.300 173.600 ;
        RECT 226.800 171.600 227.600 172.400 ;
        RECT 226.900 170.400 227.500 171.600 ;
        RECT 198.000 169.600 198.800 170.400 ;
        RECT 199.600 169.600 200.400 170.400 ;
        RECT 215.600 169.600 216.400 170.400 ;
        RECT 217.200 169.600 218.000 170.400 ;
        RECT 223.600 169.600 224.400 170.400 ;
        RECT 226.800 169.600 227.600 170.400 ;
        RECT 230.000 169.600 230.800 170.400 ;
        RECT 231.600 169.600 232.400 170.400 ;
        RECT 233.200 170.200 234.000 175.800 ;
        RECT 234.900 174.400 235.500 187.600 ;
        RECT 238.000 184.200 238.800 195.800 ;
        RECT 242.900 192.300 243.500 211.600 ;
        RECT 246.000 209.600 246.800 210.400 ;
        RECT 246.100 208.400 246.700 209.600 ;
        RECT 246.000 207.600 246.800 208.400 ;
        RECT 244.400 192.300 245.200 192.400 ;
        RECT 242.900 191.700 245.200 192.300 ;
        RECT 244.400 191.600 245.200 191.700 ;
        RECT 247.700 190.400 248.300 211.600 ;
        RECT 249.300 210.400 249.900 211.600 ;
        RECT 249.200 209.600 250.000 210.400 ;
        RECT 252.400 209.600 253.200 210.400 ;
        RECT 254.000 210.200 254.800 215.800 ;
        RECT 249.200 207.600 250.000 208.400 ;
        RECT 249.200 205.600 250.000 206.400 ;
        RECT 247.600 189.600 248.400 190.400 ;
        RECT 249.300 188.400 249.900 205.600 ;
        RECT 252.500 204.400 253.100 209.600 ;
        RECT 257.200 206.200 258.000 217.800 ;
        RECT 258.800 213.600 259.600 214.400 ;
        RECT 258.900 212.600 259.500 213.600 ;
        RECT 258.800 211.800 259.600 212.600 ;
        RECT 265.300 212.400 265.900 227.600 ;
        RECT 266.800 224.200 267.600 235.800 ;
        RECT 270.000 229.600 270.800 230.400 ;
        RECT 265.200 211.600 266.000 212.400 ;
        RECT 265.200 207.600 266.000 208.400 ;
        RECT 252.400 203.600 253.200 204.400 ;
        RECT 265.300 198.400 265.900 207.600 ;
        RECT 266.800 206.200 267.600 217.800 ;
        RECT 270.100 208.400 270.700 229.600 ;
        RECT 273.200 223.600 274.000 224.400 ;
        RECT 276.400 224.200 277.200 235.800 ;
        RECT 297.200 233.600 298.000 234.400 ;
        RECT 289.200 232.300 290.000 232.400 ;
        RECT 287.700 231.700 290.000 232.300 ;
        RECT 284.400 229.600 285.200 230.400 ;
        RECT 281.200 225.600 282.000 226.400 ;
        RECT 282.800 225.600 283.600 226.400 ;
        RECT 281.300 224.400 281.900 225.600 ;
        RECT 281.200 223.600 282.000 224.400 ;
        RECT 271.600 217.600 272.400 218.400 ;
        RECT 273.300 216.400 273.900 223.600 ;
        RECT 282.900 218.400 283.500 225.600 ;
        RECT 284.500 218.400 285.100 229.600 ;
        RECT 282.800 217.600 283.600 218.400 ;
        RECT 284.400 217.600 285.200 218.400 ;
        RECT 273.200 215.600 274.000 216.400 ;
        RECT 281.200 214.300 282.000 214.400 ;
        RECT 282.900 214.300 283.500 217.600 ;
        RECT 287.700 214.400 288.300 231.700 ;
        RECT 289.200 231.600 290.000 231.700 ;
        RECT 305.200 231.600 306.000 232.400 ;
        RECT 294.000 229.600 294.800 230.400 ;
        RECT 295.600 229.600 296.400 230.400 ;
        RECT 306.800 229.600 307.600 230.400 ;
        RECT 295.700 228.400 296.300 229.600 ;
        RECT 295.600 227.600 296.400 228.400 ;
        RECT 302.000 225.600 302.800 226.400 ;
        RECT 308.400 226.200 309.200 231.800 ;
        RECT 310.000 227.600 310.800 228.400 ;
        RECT 294.000 217.600 294.800 218.400 ;
        RECT 298.800 217.600 299.600 218.400 ;
        RECT 294.100 216.400 294.700 217.600 ;
        RECT 298.900 216.400 299.500 217.600 ;
        RECT 292.400 215.600 293.200 216.400 ;
        RECT 294.000 215.600 294.800 216.400 ;
        RECT 298.800 215.600 299.600 216.400 ;
        RECT 281.200 213.700 283.500 214.300 ;
        RECT 281.200 213.600 282.000 213.700 ;
        RECT 287.600 213.600 288.400 214.400 ;
        RECT 276.400 211.600 277.200 212.400 ;
        RECT 279.600 211.600 280.400 212.400 ;
        RECT 284.400 211.600 285.200 212.400 ;
        RECT 273.200 209.600 274.000 210.400 ;
        RECT 270.000 207.600 270.800 208.400 ;
        RECT 265.200 197.600 266.000 198.400 ;
        RECT 255.600 191.600 256.400 192.400 ;
        RECT 260.200 191.800 261.000 192.600 ;
        RECT 266.800 191.800 267.600 192.600 ;
        RECT 273.300 192.400 273.900 209.600 ;
        RECT 250.800 189.600 251.600 190.400 ;
        RECT 246.000 187.600 246.800 188.400 ;
        RECT 249.200 187.600 250.000 188.400 ;
        RECT 242.800 185.600 243.600 186.400 ;
        RECT 242.900 184.400 243.500 185.600 ;
        RECT 242.800 183.600 243.600 184.400 ;
        RECT 234.800 173.600 235.600 174.400 ;
        RECT 231.700 168.400 232.300 169.600 ;
        RECT 220.400 167.600 221.200 168.400 ;
        RECT 231.600 167.600 232.400 168.400 ;
        RECT 236.400 166.200 237.200 177.800 ;
        RECT 238.000 171.600 238.800 172.600 ;
        RECT 246.000 166.200 246.800 177.800 ;
        RECT 249.300 174.400 249.900 187.600 ;
        RECT 250.900 186.400 251.500 189.600 ;
        RECT 258.800 187.600 259.600 188.400 ;
        RECT 260.200 187.000 260.800 191.800 ;
        RECT 262.800 188.400 263.600 188.600 ;
        RECT 267.000 188.400 267.600 191.800 ;
        RECT 273.200 191.600 274.000 192.400 ;
        RECT 262.800 187.800 267.600 188.400 ;
        RECT 262.000 187.000 262.800 187.200 ;
        RECT 265.400 187.000 266.200 187.200 ;
        RECT 267.000 187.000 267.600 187.800 ;
        RECT 268.400 187.600 269.200 188.400 ;
        RECT 250.800 185.600 251.600 186.400 ;
        RECT 257.200 185.600 258.000 186.400 ;
        RECT 260.200 186.200 261.000 187.000 ;
        RECT 262.000 186.400 266.200 187.000 ;
        RECT 266.800 186.200 267.600 187.000 ;
        RECT 268.500 186.400 269.100 187.600 ;
        RECT 268.400 185.600 269.200 186.400 ;
        RECT 274.800 186.200 275.600 191.800 ;
        RECT 276.500 188.400 277.100 211.600 ;
        RECT 281.200 209.600 282.000 210.400 ;
        RECT 284.400 209.600 285.200 210.400 ;
        RECT 281.300 208.400 281.900 209.600 ;
        RECT 281.200 207.600 282.000 208.400 ;
        RECT 303.600 206.200 304.400 217.800 ;
        RECT 310.100 214.400 310.700 227.600 ;
        RECT 311.600 224.200 312.400 235.800 ;
        RECT 314.800 229.600 315.600 230.400 ;
        RECT 314.900 222.400 315.500 229.600 ;
        RECT 321.200 224.200 322.000 235.800 ;
        RECT 327.600 233.600 328.400 234.400 ;
        RECT 327.700 232.400 328.300 233.600 ;
        RECT 327.600 231.600 328.400 232.400 ;
        RECT 338.800 231.600 339.600 232.400 ;
        RECT 332.400 225.600 333.200 226.400 ;
        RECT 340.400 226.200 341.200 231.800 ;
        RECT 332.500 224.400 333.100 225.600 ;
        RECT 326.000 223.600 326.800 224.400 ;
        RECT 329.200 223.600 330.000 224.400 ;
        RECT 332.400 223.600 333.200 224.400 ;
        RECT 338.800 223.600 339.600 224.400 ;
        RECT 343.600 224.200 344.400 235.800 ;
        RECT 345.300 230.200 345.900 249.600 ;
        RECT 351.700 230.400 352.300 267.600 ;
        RECT 356.400 264.200 357.200 275.800 ;
        RECT 364.400 273.600 365.200 274.400 ;
        RECT 362.600 271.800 363.400 272.600 ;
        RECT 364.500 272.400 365.100 273.600 ;
        RECT 358.000 267.600 358.800 268.400 ;
        RECT 359.600 266.200 360.400 271.800 ;
        RECT 361.200 269.600 362.000 270.400 ;
        RECT 361.300 268.400 361.900 269.600 ;
        RECT 361.200 267.600 362.000 268.400 ;
        RECT 362.600 267.000 363.200 271.800 ;
        RECT 364.400 271.600 365.200 272.400 ;
        RECT 369.200 271.800 370.000 272.600 ;
        RECT 365.200 268.400 366.000 268.600 ;
        RECT 369.400 268.400 370.000 271.800 ;
        RECT 372.400 271.600 373.200 272.400 ;
        RECT 370.800 269.600 371.600 270.400 ;
        RECT 365.200 267.800 370.000 268.400 ;
        RECT 364.400 267.000 365.200 267.200 ;
        RECT 367.800 267.000 368.600 267.200 ;
        RECT 369.400 267.000 370.000 267.800 ;
        RECT 370.800 267.600 371.600 268.400 ;
        RECT 362.600 266.200 363.400 267.000 ;
        RECT 364.400 266.400 368.600 267.000 ;
        RECT 369.200 266.200 370.000 267.000 ;
        RECT 370.900 264.400 371.500 267.600 ;
        RECT 370.800 263.600 371.600 264.400 ;
        RECT 358.000 261.600 358.800 262.400 ;
        RECT 353.200 255.600 354.000 256.400 ;
        RECT 356.400 255.600 357.200 256.400 ;
        RECT 356.500 254.400 357.100 255.600 ;
        RECT 356.400 253.600 357.200 254.400 ;
        RECT 353.200 251.600 354.000 252.400 ;
        RECT 356.400 251.600 357.200 252.400 ;
        RECT 353.300 250.400 353.900 251.600 ;
        RECT 358.100 250.400 358.700 261.600 ;
        RECT 372.500 260.400 373.100 271.600 ;
        RECT 377.300 270.400 377.900 301.600 ;
        RECT 394.900 298.400 395.500 303.600 ;
        RECT 380.400 291.800 381.200 292.600 ;
        RECT 380.500 286.400 381.100 291.800 ;
        RECT 380.400 285.600 381.200 286.400 ;
        RECT 382.000 286.200 382.800 297.800 ;
        RECT 386.800 297.600 387.600 298.400 ;
        RECT 394.800 297.600 395.600 298.400 ;
        RECT 383.600 289.600 384.400 290.400 ;
        RECT 385.200 290.200 386.000 295.800 ;
        RECT 386.900 294.400 387.500 297.600 ;
        RECT 388.400 295.000 389.200 295.800 ;
        RECT 389.800 295.000 394.000 295.600 ;
        RECT 395.000 295.000 395.800 295.800 ;
        RECT 386.800 293.600 387.600 294.400 ;
        RECT 388.400 294.200 389.000 295.000 ;
        RECT 389.800 294.800 390.600 295.000 ;
        RECT 393.200 294.800 394.000 295.000 ;
        RECT 388.400 293.600 393.200 294.200 ;
        RECT 388.400 290.200 389.000 293.600 ;
        RECT 392.400 293.400 393.200 293.600 ;
        RECT 395.200 290.200 395.800 295.000 ;
        RECT 398.100 290.400 398.700 303.600 ;
        RECT 401.300 292.400 401.900 305.700 ;
        RECT 402.800 305.600 403.600 305.700 ;
        RECT 409.200 304.200 410.000 315.800 ;
        RECT 410.900 310.400 411.500 333.600 ;
        RECT 412.400 330.200 413.200 335.800 ;
        RECT 418.800 326.200 419.600 337.800 ;
        RECT 414.000 323.600 414.800 324.400 ;
        RECT 410.800 309.600 411.600 310.400 ;
        RECT 414.100 308.400 414.700 323.600 ;
        RECT 417.200 317.600 418.000 318.400 ;
        RECT 417.300 310.200 417.900 317.600 ;
        RECT 417.200 309.400 418.000 310.200 ;
        RECT 414.000 307.600 414.800 308.400 ;
        RECT 418.800 304.200 419.600 315.800 ;
        RECT 414.000 301.600 414.800 302.400 ;
        RECT 414.100 298.400 414.700 301.600 ;
        RECT 414.000 297.600 414.800 298.400 ;
        RECT 404.400 295.600 405.200 296.400 ;
        RECT 402.800 293.600 403.600 294.400 ;
        RECT 401.200 291.600 402.000 292.400 ;
        RECT 382.000 273.600 382.800 274.400 ;
        RECT 382.100 272.400 382.700 273.600 ;
        RECT 382.000 271.600 382.800 272.400 ;
        RECT 377.200 269.600 378.000 270.400 ;
        RECT 382.100 268.400 382.700 271.600 ;
        RECT 383.700 270.400 384.300 289.600 ;
        RECT 388.400 289.400 389.200 290.200 ;
        RECT 395.000 289.400 395.800 290.200 ;
        RECT 398.000 289.600 398.800 290.400 ;
        RECT 390.000 287.600 390.800 288.400 ;
        RECT 398.100 278.400 398.700 289.600 ;
        RECT 386.800 277.600 387.600 278.400 ;
        RECT 398.000 277.600 398.800 278.400 ;
        RECT 402.900 274.400 403.500 293.600 ;
        RECT 404.500 290.400 405.100 295.600 ;
        RECT 412.400 293.600 413.200 294.400 ;
        RECT 407.600 291.600 408.400 292.400 ;
        RECT 410.800 292.300 411.600 292.400 ;
        RECT 409.300 291.700 411.600 292.300 ;
        RECT 404.400 289.600 405.200 290.400 ;
        RECT 409.300 278.400 409.900 291.700 ;
        RECT 410.800 291.600 411.600 291.700 ;
        RECT 412.500 290.300 413.100 293.600 ;
        RECT 410.900 289.700 413.100 290.300 ;
        RECT 410.900 278.400 411.500 289.700 ;
        RECT 418.800 286.200 419.600 297.800 ;
        RECT 420.500 292.400 421.100 377.600 ;
        RECT 422.000 364.200 422.800 377.800 ;
        RECT 423.600 364.200 424.400 377.800 ;
        RECT 425.200 364.200 426.000 377.800 ;
        RECT 426.800 366.200 427.600 377.800 ;
        RECT 428.400 377.600 429.200 378.400 ;
        RECT 428.500 376.400 429.100 377.600 ;
        RECT 428.400 375.600 429.200 376.400 ;
        RECT 430.000 366.200 430.800 377.800 ;
        RECT 433.200 366.200 434.000 377.800 ;
        RECT 434.800 364.200 435.600 377.800 ;
        RECT 436.400 364.200 437.200 377.800 ;
        RECT 438.000 371.600 438.800 372.400 ;
        RECT 438.100 370.800 438.700 371.600 ;
        RECT 438.000 370.000 438.800 370.800 ;
        RECT 425.200 353.600 426.000 354.400 ;
        RECT 431.600 353.600 432.400 354.400 ;
        RECT 425.300 348.400 425.900 353.600 ;
        RECT 431.700 352.400 432.300 353.600 ;
        RECT 426.800 351.600 427.600 352.400 ;
        RECT 431.600 351.600 432.400 352.400 ;
        RECT 426.900 350.400 427.500 351.600 ;
        RECT 426.800 349.600 427.600 350.400 ;
        RECT 430.000 349.600 430.800 350.400 ;
        RECT 434.800 349.600 435.600 350.400 ;
        RECT 426.900 348.400 427.500 349.600 ;
        RECT 423.600 347.600 424.400 348.400 ;
        RECT 425.200 347.600 426.000 348.400 ;
        RECT 426.800 347.600 427.600 348.400 ;
        RECT 438.000 347.600 438.800 348.400 ;
        RECT 423.700 346.400 424.300 347.600 ;
        RECT 439.700 346.400 440.300 379.600 ;
        RECT 450.900 376.400 451.500 407.600 ;
        RECT 457.300 400.400 457.900 411.600 ;
        RECT 463.600 403.600 464.400 404.400 ;
        RECT 473.200 404.200 474.000 417.800 ;
        RECT 474.800 404.200 475.600 417.800 ;
        RECT 476.400 404.200 477.200 417.800 ;
        RECT 478.000 406.200 478.800 417.800 ;
        RECT 479.600 415.600 480.400 416.400 ;
        RECT 457.200 399.600 458.000 400.400 ;
        RECT 454.000 384.200 454.800 397.800 ;
        RECT 455.600 384.200 456.400 397.800 ;
        RECT 457.200 384.200 458.000 397.800 ;
        RECT 458.800 384.200 459.600 395.800 ;
        RECT 460.400 385.600 461.200 386.400 ;
        RECT 460.500 378.400 461.100 385.600 ;
        RECT 462.000 384.200 462.800 395.800 ;
        RECT 465.200 384.200 466.000 395.800 ;
        RECT 466.800 384.200 467.600 397.800 ;
        RECT 468.400 384.200 469.200 397.800 ;
        RECT 474.800 391.600 475.600 392.400 ;
        RECT 473.200 389.600 474.000 390.400 ;
        RECT 474.900 388.400 475.500 391.600 ;
        RECT 474.800 387.600 475.600 388.400 ;
        RECT 478.000 387.600 478.800 388.400 ;
        RECT 479.700 386.400 480.300 415.600 ;
        RECT 481.200 406.200 482.000 417.800 ;
        RECT 484.400 406.200 485.200 417.800 ;
        RECT 486.000 404.200 486.800 417.800 ;
        RECT 487.600 404.200 488.400 417.800 ;
        RECT 506.800 415.600 507.600 416.400 ;
        RECT 514.800 415.600 515.600 416.400 ;
        RECT 494.000 413.600 494.800 414.400 ;
        RECT 497.200 413.600 498.000 414.400 ;
        RECT 492.400 411.600 493.200 412.400 ;
        RECT 494.100 410.400 494.700 413.600 ;
        RECT 514.900 412.400 515.500 415.600 ;
        RECT 502.000 411.600 502.800 412.400 ;
        RECT 514.800 411.600 515.600 412.400 ;
        RECT 494.000 409.600 494.800 410.400 ;
        RECT 521.200 404.200 522.000 417.800 ;
        RECT 522.800 404.200 523.600 417.800 ;
        RECT 524.400 406.200 525.200 417.800 ;
        RECT 526.000 413.600 526.800 414.400 ;
        RECT 527.600 406.200 528.400 417.800 ;
        RECT 529.200 415.600 530.000 416.400 ;
        RECT 529.300 404.300 529.900 415.600 ;
        RECT 530.800 406.200 531.600 417.800 ;
        RECT 527.700 403.700 529.900 404.300 ;
        RECT 532.400 404.200 533.200 417.800 ;
        RECT 534.000 404.200 534.800 417.800 ;
        RECT 535.600 404.200 536.400 417.800 ;
        RECT 543.600 413.600 544.400 414.400 ;
        RECT 537.200 411.600 538.000 412.400 ;
        RECT 481.200 389.600 482.000 390.400 ;
        RECT 498.800 389.600 499.600 390.400 ;
        RECT 505.200 389.600 506.000 390.400 ;
        RECT 510.000 389.600 510.800 390.400 ;
        RECT 514.800 389.600 515.600 390.400 ;
        RECT 474.800 385.600 475.600 386.400 ;
        RECT 479.600 385.600 480.400 386.400 ;
        RECT 487.600 385.600 488.400 386.400 ;
        RECT 495.600 385.600 496.400 386.400 ;
        RECT 460.400 377.600 461.200 378.400 ;
        RECT 450.800 375.600 451.600 376.400 ;
        RECT 455.600 375.600 456.400 376.400 ;
        RECT 441.200 371.600 442.000 372.400 ;
        RECT 446.000 371.600 446.800 372.400 ;
        RECT 458.800 363.600 459.600 364.400 ;
        RECT 468.400 364.200 469.200 377.800 ;
        RECT 470.000 364.200 470.800 377.800 ;
        RECT 471.600 364.200 472.400 377.800 ;
        RECT 473.200 366.200 474.000 377.800 ;
        RECT 474.900 376.400 475.500 385.600 ;
        RECT 474.800 375.600 475.600 376.400 ;
        RECT 441.200 351.600 442.000 352.400 ;
        RECT 450.800 351.600 451.600 352.400 ;
        RECT 457.200 351.600 458.000 352.400 ;
        RECT 449.200 347.600 450.000 348.400 ;
        RECT 449.300 346.400 449.900 347.600 ;
        RECT 450.900 346.400 451.500 351.600 ;
        RECT 457.300 350.400 457.900 351.600 ;
        RECT 452.400 349.600 453.200 350.400 ;
        RECT 457.200 349.600 458.000 350.400 ;
        RECT 454.000 347.600 454.800 348.400 ;
        RECT 423.600 345.600 424.400 346.400 ;
        RECT 439.600 345.600 440.400 346.400 ;
        RECT 442.800 345.600 443.600 346.400 ;
        RECT 449.200 345.600 450.000 346.400 ;
        RECT 450.800 345.600 451.600 346.400 ;
        RECT 442.900 344.400 443.500 345.600 ;
        RECT 430.000 343.600 430.800 344.400 ;
        RECT 442.800 343.600 443.600 344.400 ;
        RECT 455.600 343.600 456.400 344.400 ;
        RECT 423.600 333.600 424.400 334.400 ;
        RECT 426.800 331.600 427.600 332.600 ;
        RECT 426.800 325.600 427.600 326.400 ;
        RECT 428.400 326.200 429.200 337.800 ;
        RECT 430.100 334.400 430.700 343.600 ;
        RECT 449.200 339.600 450.000 340.400 ;
        RECT 450.800 339.600 451.600 340.400 ;
        RECT 430.000 333.600 430.800 334.400 ;
        RECT 431.600 330.200 432.400 335.800 ;
        RECT 434.600 335.000 435.400 335.800 ;
        RECT 436.400 335.000 440.600 335.600 ;
        RECT 441.200 335.000 442.000 335.800 ;
        RECT 433.200 333.600 434.000 334.400 ;
        RECT 434.600 330.200 435.200 335.000 ;
        RECT 436.400 334.800 437.200 335.000 ;
        RECT 439.800 334.800 440.600 335.000 ;
        RECT 441.400 334.200 442.000 335.000 ;
        RECT 437.200 333.600 442.000 334.200 ;
        RECT 447.600 333.600 448.400 334.400 ;
        RECT 437.200 333.400 438.000 333.600 ;
        RECT 436.400 331.600 437.200 332.400 ;
        RECT 434.600 329.400 435.400 330.200 ;
        RECT 436.500 328.400 437.100 331.600 ;
        RECT 441.400 330.200 442.000 333.600 ;
        RECT 449.300 332.400 449.900 339.600 ;
        RECT 449.200 331.600 450.000 332.400 ;
        RECT 441.200 329.400 442.000 330.200 ;
        RECT 436.400 327.600 437.200 328.400 ;
        RECT 422.000 306.200 422.800 311.800 ;
        RECT 425.200 311.600 426.000 312.400 ;
        RECT 423.600 309.600 424.400 310.400 ;
        RECT 423.700 308.400 424.300 309.600 ;
        RECT 425.300 308.400 425.900 311.600 ;
        RECT 423.600 307.600 424.400 308.400 ;
        RECT 425.200 307.600 426.000 308.400 ;
        RECT 425.200 303.600 426.000 304.400 ;
        RECT 425.300 292.400 425.900 303.600 ;
        RECT 420.400 291.600 421.200 292.400 ;
        RECT 425.200 291.600 426.000 292.400 ;
        RECT 409.200 277.600 410.000 278.400 ;
        RECT 410.800 277.600 411.600 278.400 ;
        RECT 385.200 273.600 386.000 274.400 ;
        RECT 402.800 273.600 403.600 274.400 ;
        RECT 412.400 273.600 413.200 274.400 ;
        RECT 385.300 272.400 385.900 273.600 ;
        RECT 385.200 271.600 386.000 272.400 ;
        RECT 388.400 271.600 389.200 272.400 ;
        RECT 394.800 271.600 395.600 272.400 ;
        RECT 398.000 272.300 398.800 272.400 ;
        RECT 396.500 271.700 398.800 272.300 ;
        RECT 388.500 270.400 389.100 271.600 ;
        RECT 383.600 269.600 384.400 270.400 ;
        RECT 386.800 269.600 387.600 270.400 ;
        RECT 388.400 269.600 389.200 270.400 ;
        RECT 390.000 269.600 390.800 270.400 ;
        RECT 374.000 267.600 374.800 268.400 ;
        RECT 377.200 267.600 378.000 268.400 ;
        RECT 382.000 267.600 382.800 268.400 ;
        RECT 372.400 259.600 373.200 260.400 ;
        RECT 366.000 257.600 366.800 258.400 ;
        RECT 367.600 257.600 368.400 258.400 ;
        RECT 366.100 256.400 366.700 257.600 ;
        RECT 366.000 255.600 366.800 256.400 ;
        RECT 362.800 253.600 363.600 254.400 ;
        RECT 366.100 252.400 366.700 255.600 ;
        RECT 367.700 254.400 368.300 257.600 ;
        RECT 367.600 253.600 368.400 254.400 ;
        RECT 361.200 251.600 362.000 252.400 ;
        RECT 366.000 251.600 366.800 252.400 ;
        RECT 353.200 249.600 354.000 250.400 ;
        RECT 358.000 249.600 358.800 250.400 ;
        RECT 364.400 249.600 365.200 250.400 ;
        RECT 372.400 246.200 373.200 257.800 ;
        RECT 374.100 254.400 374.700 267.600 ;
        RECT 380.400 265.600 381.200 266.400 ;
        RECT 383.700 264.400 384.300 269.600 ;
        RECT 383.600 263.600 384.400 264.400 ;
        RECT 374.000 253.600 374.800 254.400 ;
        RECT 380.400 251.600 381.200 252.600 ;
        RECT 382.000 246.200 382.800 257.800 ;
        RECT 383.600 253.600 384.400 254.400 ;
        RECT 385.200 250.200 386.000 255.800 ;
        RECT 386.900 252.400 387.500 269.600 ;
        RECT 390.100 268.400 390.700 269.600 ;
        RECT 390.000 267.600 390.800 268.400 ;
        RECT 396.500 266.400 397.100 271.700 ;
        RECT 398.000 271.600 398.800 271.700 ;
        RECT 402.900 268.400 403.500 273.600 ;
        RECT 404.400 271.600 405.200 272.400 ;
        RECT 406.000 269.600 406.800 270.400 ;
        RECT 402.800 267.600 403.600 268.400 ;
        RECT 406.100 266.400 406.700 269.600 ;
        RECT 412.500 266.400 413.100 273.600 ;
        RECT 393.200 265.600 394.000 266.400 ;
        RECT 396.400 265.600 397.200 266.400 ;
        RECT 402.800 265.600 403.600 266.400 ;
        RECT 406.000 265.600 406.800 266.400 ;
        RECT 412.400 265.600 413.200 266.400 ;
        RECT 393.300 264.400 393.900 265.600 ;
        RECT 388.400 263.600 389.200 264.400 ;
        RECT 391.600 263.600 392.400 264.400 ;
        RECT 393.200 263.600 394.000 264.400 ;
        RECT 396.400 263.600 397.200 264.400 ;
        RECT 398.000 263.600 398.800 264.400 ;
        RECT 388.500 254.400 389.100 263.600 ;
        RECT 391.700 254.400 392.300 263.600 ;
        RECT 393.200 259.600 394.000 260.400 ;
        RECT 388.400 253.600 389.200 254.400 ;
        RECT 391.600 253.600 392.400 254.400 ;
        RECT 393.300 252.400 393.900 259.600 ;
        RECT 396.500 258.400 397.100 263.600 ;
        RECT 398.100 260.400 398.700 263.600 ;
        RECT 398.000 259.600 398.800 260.400 ;
        RECT 406.100 258.400 406.700 265.600 ;
        RECT 409.200 263.600 410.000 264.400 ;
        RECT 410.800 263.600 411.600 264.400 ;
        RECT 418.800 264.200 419.600 275.800 ;
        RECT 420.500 270.400 421.100 291.600 ;
        RECT 422.000 273.600 422.800 274.400 ;
        RECT 420.400 269.600 421.200 270.400 ;
        RECT 396.400 257.600 397.200 258.400 ;
        RECT 399.600 257.600 400.400 258.400 ;
        RECT 394.800 255.600 395.600 256.400 ;
        RECT 386.800 251.600 387.600 252.400 ;
        RECT 390.000 251.600 390.800 252.400 ;
        RECT 393.200 251.600 394.000 252.400 ;
        RECT 398.000 251.600 398.800 252.400 ;
        RECT 404.400 246.200 405.200 257.800 ;
        RECT 406.000 257.600 406.800 258.400 ;
        RECT 409.300 252.400 409.900 263.600 ;
        RECT 410.900 256.400 411.500 263.600 ;
        RECT 410.800 255.600 411.600 256.400 ;
        RECT 409.200 251.600 410.000 252.400 ;
        RECT 414.000 246.200 414.800 257.800 ;
        RECT 418.800 257.600 419.600 258.400 ;
        RECT 415.600 253.600 416.400 254.400 ;
        RECT 417.200 250.200 418.000 255.800 ;
        RECT 345.200 229.400 346.000 230.200 ;
        RECT 351.600 229.600 352.400 230.400 ;
        RECT 345.200 223.600 346.000 224.400 ;
        RECT 353.200 224.200 354.000 235.800 ;
        RECT 358.000 234.300 358.800 234.400 ;
        RECT 358.000 233.700 360.300 234.300 ;
        RECT 358.000 233.600 358.800 233.700 ;
        RECT 359.700 230.400 360.300 233.700 ;
        RECT 359.600 229.600 360.400 230.400 ;
        RECT 362.800 229.600 363.600 230.400 ;
        RECT 362.900 228.400 363.500 229.600 ;
        RECT 362.800 227.600 363.600 228.400 ;
        RECT 364.400 223.600 365.200 224.400 ;
        RECT 369.200 224.200 370.000 235.800 ;
        RECT 375.600 229.600 376.400 230.400 ;
        RECT 378.800 224.200 379.600 235.800 ;
        RECT 382.000 226.200 382.800 231.800 ;
        RECT 383.600 226.200 384.400 231.800 ;
        RECT 386.800 224.200 387.600 235.800 ;
        RECT 388.400 229.400 389.200 230.200 ;
        RECT 394.800 229.600 395.600 230.400 ;
        RECT 314.800 221.600 315.600 222.400 ;
        RECT 326.000 221.600 326.800 222.400 ;
        RECT 310.000 213.600 310.800 214.400 ;
        RECT 305.200 211.600 306.000 212.400 ;
        RECT 311.600 211.600 312.400 212.600 ;
        RECT 298.800 203.600 299.600 204.400 ;
        RECT 276.400 187.600 277.200 188.400 ;
        RECT 273.200 183.600 274.000 184.400 ;
        RECT 249.200 173.600 250.000 174.400 ;
        RECT 265.200 173.600 266.000 174.400 ;
        RECT 266.800 170.200 267.600 175.800 ;
        RECT 268.400 173.600 269.200 174.400 ;
        RECT 270.000 166.200 270.800 177.800 ;
        RECT 276.500 174.400 277.100 187.600 ;
        RECT 278.000 184.200 278.800 195.800 ;
        RECT 279.600 189.400 280.400 190.400 ;
        RECT 287.600 184.200 288.400 195.800 ;
        RECT 298.900 188.400 299.500 203.600 ;
        RECT 302.000 191.600 302.800 192.400 ;
        RECT 303.600 191.600 304.400 192.400 ;
        RECT 303.700 190.400 304.300 191.600 ;
        RECT 303.600 189.600 304.400 190.400 ;
        RECT 298.800 187.600 299.600 188.400 ;
        RECT 292.400 185.600 293.200 186.400 ;
        RECT 292.500 184.400 293.100 185.600 ;
        RECT 292.400 183.600 293.200 184.400 ;
        RECT 276.400 173.600 277.200 174.400 ;
        RECT 271.600 171.800 272.400 172.600 ;
        RECT 271.700 170.400 272.300 171.800 ;
        RECT 271.600 169.600 272.400 170.400 ;
        RECT 279.600 166.200 280.400 177.800 ;
        RECT 290.800 170.200 291.600 175.800 ;
        RECT 292.400 173.600 293.200 174.400 ;
        RECT 284.400 167.600 285.200 168.400 ;
        RECT 294.000 166.200 294.800 177.800 ;
        RECT 295.600 171.800 296.400 172.600 ;
        RECT 295.700 166.400 296.300 171.800 ;
        RECT 298.900 170.400 299.500 187.600 ;
        RECT 298.800 169.600 299.600 170.400 ;
        RECT 295.600 165.600 296.400 166.400 ;
        RECT 303.600 166.200 304.400 177.800 ;
        RECT 305.300 168.400 305.900 211.600 ;
        RECT 313.200 206.200 314.000 217.800 ;
        RECT 316.400 210.200 317.200 215.800 ;
        RECT 318.000 213.600 318.800 214.400 ;
        RECT 318.100 212.400 318.700 213.600 ;
        RECT 318.000 211.600 318.800 212.400 ;
        RECT 321.200 211.600 322.000 212.400 ;
        RECT 321.300 208.300 321.900 211.600 ;
        RECT 322.800 208.300 323.600 208.400 ;
        RECT 321.300 207.700 323.600 208.300 ;
        RECT 322.800 207.600 323.600 207.700 ;
        RECT 326.100 198.400 326.700 221.600 ;
        RECT 329.300 218.400 329.900 223.600 ;
        RECT 327.600 206.200 328.400 217.800 ;
        RECT 329.200 217.600 330.000 218.400 ;
        RECT 335.600 215.600 336.400 216.400 ;
        RECT 329.200 213.600 330.000 214.400 ;
        RECT 329.300 212.400 329.900 213.600 ;
        RECT 335.700 212.600 336.300 215.600 ;
        RECT 329.200 211.600 330.000 212.400 ;
        RECT 335.600 211.800 336.400 212.600 ;
        RECT 337.200 206.200 338.000 217.800 ;
        RECT 338.900 212.400 339.500 223.600 ;
        RECT 338.800 211.600 339.600 212.400 ;
        RECT 340.400 210.200 341.200 215.800 ;
        RECT 342.000 215.600 342.800 216.400 ;
        RECT 345.300 212.400 345.900 223.600 ;
        RECT 388.500 218.400 389.100 229.400 ;
        RECT 396.400 224.200 397.200 235.800 ;
        RECT 401.200 235.600 402.000 236.400 ;
        RECT 402.800 226.200 403.600 231.800 ;
        RECT 404.400 229.600 405.200 230.400 ;
        RECT 404.500 228.400 405.100 229.600 ;
        RECT 404.400 227.600 405.200 228.400 ;
        RECT 406.000 224.200 406.800 235.800 ;
        RECT 407.600 229.400 408.400 230.200 ;
        RECT 414.000 229.600 414.800 230.400 ;
        RECT 407.700 218.400 408.300 229.400 ;
        RECT 414.100 222.300 414.700 229.600 ;
        RECT 415.600 224.200 416.400 235.800 ;
        RECT 422.100 234.400 422.700 273.600 ;
        RECT 426.900 270.200 427.500 325.600 ;
        RECT 428.400 315.600 429.200 316.400 ;
        RECT 428.500 308.400 429.100 315.600 ;
        RECT 444.400 313.600 445.200 314.400 ;
        RECT 444.500 312.400 445.100 313.600 ;
        RECT 434.800 311.600 435.600 312.400 ;
        RECT 438.000 311.600 438.800 312.400 ;
        RECT 444.400 311.600 445.200 312.400 ;
        RECT 434.900 310.400 435.500 311.600 ;
        RECT 438.100 310.400 438.700 311.600 ;
        RECT 430.000 309.600 430.800 310.400 ;
        RECT 434.800 309.600 435.600 310.400 ;
        RECT 438.000 309.600 438.800 310.400 ;
        RECT 439.600 309.600 440.400 310.400 ;
        RECT 450.900 308.400 451.500 339.600 ;
        RECT 454.000 333.600 454.800 334.400 ;
        RECT 455.700 332.400 456.300 343.600 ;
        RECT 455.600 331.600 456.400 332.400 ;
        RECT 457.300 326.400 457.900 349.600 ;
        RECT 458.900 348.400 459.500 363.600 ;
        RECT 474.900 354.400 475.500 375.600 ;
        RECT 476.400 366.200 477.200 377.800 ;
        RECT 479.600 366.200 480.400 377.800 ;
        RECT 481.200 364.200 482.000 377.800 ;
        RECT 482.800 364.200 483.600 377.800 ;
        RECT 487.700 376.400 488.300 385.600 ;
        RECT 490.800 383.600 491.600 384.400 ;
        RECT 487.600 375.600 488.400 376.400 ;
        RECT 487.600 371.600 488.400 372.400 ;
        RECT 489.200 370.300 490.000 370.400 ;
        RECT 490.900 370.300 491.500 383.600 ;
        RECT 497.200 375.600 498.000 376.400 ;
        RECT 492.400 371.600 493.200 372.400 ;
        RECT 489.200 369.700 491.500 370.300 ;
        RECT 489.200 369.600 490.000 369.700 ;
        RECT 498.900 364.400 499.500 389.600 ;
        RECT 502.000 383.600 502.800 384.400 ;
        RECT 502.100 376.400 502.700 383.600 ;
        RECT 510.100 380.400 510.700 389.600 ;
        RECT 514.900 384.400 515.500 389.600 ;
        RECT 514.800 383.600 515.600 384.400 ;
        RECT 519.600 384.200 520.400 397.800 ;
        RECT 521.200 384.200 522.000 397.800 ;
        RECT 522.800 384.200 523.600 395.800 ;
        RECT 524.400 387.600 525.200 388.400 ;
        RECT 524.500 380.400 525.100 387.600 ;
        RECT 526.000 384.200 526.800 395.800 ;
        RECT 527.700 386.400 528.300 403.700 ;
        RECT 537.300 402.400 537.900 411.600 ;
        RECT 537.200 401.600 538.000 402.400 ;
        RECT 543.700 398.400 544.300 413.600 ;
        RECT 546.800 411.600 547.600 412.400 ;
        RECT 558.000 411.600 558.800 412.400 ;
        RECT 545.200 403.600 546.000 404.400 ;
        RECT 527.600 385.600 528.400 386.400 ;
        RECT 510.000 379.600 510.800 380.400 ;
        RECT 524.400 379.600 525.200 380.400 ;
        RECT 502.000 375.600 502.800 376.400 ;
        RECT 502.100 372.400 502.700 375.600 ;
        RECT 502.000 371.600 502.800 372.400 ;
        RECT 498.800 363.600 499.600 364.400 ;
        RECT 506.800 364.200 507.600 377.800 ;
        RECT 508.400 364.200 509.200 377.800 ;
        RECT 510.000 366.200 510.800 377.800 ;
        RECT 511.600 371.600 512.400 372.400 ;
        RECT 511.700 358.400 512.300 371.600 ;
        RECT 513.200 366.200 514.000 377.800 ;
        RECT 514.800 375.600 515.600 376.400 ;
        RECT 514.900 372.400 515.500 375.600 ;
        RECT 514.800 371.600 515.600 372.400 ;
        RECT 516.400 366.200 517.200 377.800 ;
        RECT 518.000 364.200 518.800 377.800 ;
        RECT 519.600 364.200 520.400 377.800 ;
        RECT 521.200 364.200 522.000 377.800 ;
        RECT 527.700 372.400 528.300 385.600 ;
        RECT 529.200 384.200 530.000 395.800 ;
        RECT 530.800 384.200 531.600 397.800 ;
        RECT 532.400 384.200 533.200 397.800 ;
        RECT 534.000 384.200 534.800 397.800 ;
        RECT 543.600 397.600 544.400 398.400 ;
        RECT 545.300 388.400 545.900 403.600 ;
        RECT 545.200 387.600 546.000 388.400 ;
        RECT 530.800 379.600 531.600 380.400 ;
        RECT 530.900 378.400 531.500 379.600 ;
        RECT 530.800 377.600 531.600 378.400 ;
        RECT 546.900 374.400 547.500 411.600 ;
        RECT 550.000 403.600 550.800 404.400 ;
        RECT 559.600 404.200 560.400 417.800 ;
        RECT 561.200 404.200 562.000 417.800 ;
        RECT 562.800 404.200 563.600 417.800 ;
        RECT 564.400 406.200 565.200 417.800 ;
        RECT 566.000 415.600 566.800 416.400 ;
        RECT 546.800 373.600 547.600 374.400 ;
        RECT 527.600 371.600 528.400 372.400 ;
        RECT 542.000 371.600 542.800 372.400 ;
        RECT 542.100 364.400 542.700 371.600 ;
        RECT 535.600 363.600 536.400 364.400 ;
        RECT 542.000 363.600 542.800 364.400 ;
        RECT 545.200 363.600 546.000 364.400 ;
        RECT 481.200 357.600 482.000 358.400 ;
        RECT 511.600 357.600 512.400 358.400 ;
        RECT 474.800 353.600 475.600 354.400 ;
        RECT 484.400 353.600 485.200 354.400 ;
        RECT 463.600 351.600 464.400 352.400 ;
        RECT 468.400 351.600 469.200 352.400 ;
        RECT 471.600 351.800 472.400 352.600 ;
        RECT 478.200 351.800 479.000 352.600 ;
        RECT 463.700 350.400 464.300 351.600 ;
        RECT 463.600 349.600 464.400 350.400 ;
        RECT 471.600 348.400 472.200 351.800 ;
        RECT 475.600 348.400 476.400 348.600 ;
        RECT 458.800 347.600 459.600 348.400 ;
        RECT 463.600 347.600 464.400 348.400 ;
        RECT 468.400 347.600 469.200 348.400 ;
        RECT 471.600 347.800 476.400 348.400 ;
        RECT 458.900 346.400 459.500 347.600 ;
        RECT 458.800 345.600 459.600 346.400 ;
        RECT 458.900 330.400 459.500 345.600 ;
        RECT 460.400 343.600 461.200 344.400 ;
        RECT 460.500 334.400 461.100 343.600 ;
        RECT 463.700 336.400 464.300 347.600 ;
        RECT 471.600 347.000 472.200 347.800 ;
        RECT 473.000 347.000 473.800 347.200 ;
        RECT 476.400 347.000 477.200 347.200 ;
        RECT 478.400 347.000 479.000 351.800 ;
        RECT 471.600 346.200 472.400 347.000 ;
        RECT 473.000 346.400 477.200 347.000 ;
        RECT 468.400 343.600 469.200 344.400 ;
        RECT 473.200 343.600 474.000 344.400 ;
        RECT 463.600 335.600 464.400 336.400 ;
        RECT 460.400 333.600 461.200 334.400 ;
        RECT 468.500 332.400 469.100 343.600 ;
        RECT 470.000 339.600 470.800 340.400 ;
        RECT 470.100 334.400 470.700 339.600 ;
        RECT 473.300 338.400 473.900 343.600 ;
        RECT 474.900 338.400 475.500 346.400 ;
        RECT 478.200 346.200 479.000 347.000 ;
        RECT 486.000 344.200 486.800 355.800 ;
        RECT 494.100 350.200 494.700 350.300 ;
        RECT 494.000 349.400 494.800 350.200 ;
        RECT 487.600 347.600 488.400 348.400 ;
        RECT 473.200 337.600 474.000 338.400 ;
        RECT 474.800 337.600 475.600 338.400 ;
        RECT 470.000 333.600 470.800 334.400 ;
        RECT 460.400 331.600 461.200 332.400 ;
        RECT 468.400 331.600 469.200 332.400 ;
        RECT 458.800 329.600 459.600 330.400 ;
        RECT 468.400 329.600 469.200 330.400 ;
        RECT 474.800 329.600 475.600 330.400 ;
        RECT 476.400 330.200 477.200 335.800 ;
        RECT 463.600 327.600 464.400 328.400 ;
        RECT 457.200 325.600 458.000 326.400 ;
        RECT 455.600 323.600 456.400 324.400 ;
        RECT 454.000 312.300 454.800 312.400 ;
        RECT 455.700 312.300 456.300 323.600 ;
        RECT 458.800 313.600 459.600 314.400 ;
        RECT 454.000 311.700 456.300 312.300 ;
        RECT 454.000 311.600 454.800 311.700 ;
        RECT 428.400 307.600 429.200 308.400 ;
        RECT 441.200 307.600 442.000 308.400 ;
        RECT 450.800 307.600 451.600 308.400 ;
        RECT 452.400 307.600 453.200 308.400 ;
        RECT 441.300 306.400 441.900 307.600 ;
        RECT 441.200 305.600 442.000 306.400 ;
        RECT 433.200 303.600 434.000 304.400 ;
        RECT 449.200 303.600 450.000 304.400 ;
        RECT 428.400 286.200 429.200 297.800 ;
        RECT 431.600 290.200 432.400 295.800 ;
        RECT 433.300 294.400 433.900 303.600 ;
        RECT 449.300 296.400 449.900 303.600 ;
        RECT 434.800 295.000 435.600 295.800 ;
        RECT 436.200 295.000 440.400 295.600 ;
        RECT 441.400 295.000 442.200 295.800 ;
        RECT 449.200 295.600 450.000 296.400 ;
        RECT 433.200 293.600 434.000 294.400 ;
        RECT 434.800 294.200 435.400 295.000 ;
        RECT 436.200 294.800 437.000 295.000 ;
        RECT 439.600 294.800 440.400 295.000 ;
        RECT 434.800 293.600 439.600 294.200 ;
        RECT 434.800 290.200 435.400 293.600 ;
        RECT 438.800 293.400 439.600 293.600 ;
        RECT 441.600 290.200 442.200 295.000 ;
        RECT 452.500 294.400 453.100 307.600 ;
        RECT 442.800 293.600 443.600 294.400 ;
        RECT 452.400 293.600 453.200 294.400 ;
        RECT 452.500 290.400 453.100 293.600 ;
        RECT 454.100 292.400 454.700 311.600 ;
        RECT 458.900 310.400 459.500 313.600 ;
        RECT 457.200 309.600 458.000 310.400 ;
        RECT 458.800 309.600 459.600 310.400 ;
        RECT 463.700 308.400 464.300 327.600 ;
        RECT 476.400 325.600 477.200 326.400 ;
        RECT 479.600 326.200 480.400 337.800 ;
        RECT 487.700 332.400 488.300 347.600 ;
        RECT 494.100 338.400 494.700 349.400 ;
        RECT 495.600 344.200 496.400 355.800 ;
        RECT 497.200 347.600 498.000 348.400 ;
        RECT 486.000 331.600 486.800 332.400 ;
        RECT 487.600 331.600 488.400 332.400 ;
        RECT 476.500 318.400 477.100 325.600 ;
        RECT 468.400 317.600 469.200 318.400 ;
        RECT 476.400 317.600 477.200 318.400 ;
        RECT 466.800 311.800 467.600 312.600 ;
        RECT 473.400 311.800 474.200 312.600 ;
        RECT 466.800 308.400 467.400 311.800 ;
        RECT 470.800 308.400 471.600 308.600 ;
        RECT 460.400 307.600 461.200 308.400 ;
        RECT 463.600 307.600 464.400 308.400 ;
        RECT 466.800 307.800 471.600 308.400 ;
        RECT 466.800 307.000 467.400 307.800 ;
        RECT 468.200 307.000 469.000 307.200 ;
        RECT 471.600 307.000 472.400 307.200 ;
        RECT 473.600 307.000 474.200 311.800 ;
        RECT 474.800 309.600 475.600 310.400 ;
        RECT 474.900 308.400 475.500 309.600 ;
        RECT 474.800 307.600 475.600 308.400 ;
        RECT 462.000 305.600 462.800 306.400 ;
        RECT 466.800 306.200 467.600 307.000 ;
        RECT 468.200 306.400 472.400 307.000 ;
        RECT 473.400 306.200 474.200 307.000 ;
        RECT 478.000 305.600 478.800 306.400 ;
        RECT 479.600 306.200 480.400 311.800 ;
        RECT 481.200 309.600 482.000 310.400 ;
        RECT 462.100 304.400 462.700 305.600 ;
        RECT 481.300 304.400 481.900 309.600 ;
        RECT 455.600 303.600 456.400 304.400 ;
        RECT 462.000 303.600 462.800 304.400 ;
        RECT 481.200 303.600 482.000 304.400 ;
        RECT 482.800 304.200 483.600 315.800 ;
        RECT 484.400 309.400 485.200 310.400 ;
        RECT 486.100 306.300 486.700 331.600 ;
        RECT 489.200 326.200 490.000 337.800 ;
        RECT 494.000 337.600 494.800 338.400 ;
        RECT 495.600 330.200 496.400 335.800 ;
        RECT 497.300 334.400 497.900 347.600 ;
        RECT 498.800 346.200 499.600 351.800 ;
        RECT 518.000 349.600 518.800 350.400 ;
        RECT 521.200 347.600 522.000 348.400 ;
        RECT 511.600 345.600 512.400 346.400 ;
        RECT 511.700 344.400 512.300 345.600 ;
        RECT 511.600 343.600 512.400 344.400 ;
        RECT 497.200 333.600 498.000 334.400 ;
        RECT 498.800 326.200 499.600 337.800 ;
        RECT 500.400 331.800 501.200 332.600 ;
        RECT 500.500 318.400 501.100 331.800 ;
        RECT 506.800 331.600 507.600 332.400 ;
        RECT 508.400 326.200 509.200 337.800 ;
        RECT 511.700 332.400 512.300 343.600 ;
        RECT 521.300 338.400 521.900 347.600 ;
        RECT 522.800 344.200 523.600 357.800 ;
        RECT 524.400 344.200 525.200 357.800 ;
        RECT 526.000 344.200 526.800 355.800 ;
        RECT 527.600 347.600 528.400 348.400 ;
        RECT 529.200 344.200 530.000 355.800 ;
        RECT 530.800 345.600 531.600 346.400 ;
        RECT 530.900 340.400 531.500 345.600 ;
        RECT 532.400 344.200 533.200 355.800 ;
        RECT 534.000 344.200 534.800 357.800 ;
        RECT 535.600 344.200 536.400 357.800 ;
        RECT 537.200 344.200 538.000 357.800 ;
        RECT 530.800 339.600 531.600 340.400 ;
        RECT 537.200 339.600 538.000 340.400 ;
        RECT 545.300 340.300 545.900 363.600 ;
        RECT 546.800 347.600 547.800 348.400 ;
        RECT 545.300 339.700 547.500 340.300 ;
        RECT 513.200 337.600 514.000 338.400 ;
        RECT 521.200 337.600 522.000 338.400 ;
        RECT 511.600 331.600 512.400 332.400 ;
        RECT 530.800 324.200 531.600 337.800 ;
        RECT 532.400 324.200 533.200 337.800 ;
        RECT 534.000 324.200 534.800 337.800 ;
        RECT 535.600 326.200 536.400 337.800 ;
        RECT 537.300 336.400 537.900 339.600 ;
        RECT 537.200 335.600 538.000 336.400 ;
        RECT 538.800 326.200 539.600 337.800 ;
        RECT 540.400 335.600 541.200 336.400 ;
        RECT 540.500 334.400 541.100 335.600 ;
        RECT 540.400 333.600 541.200 334.400 ;
        RECT 542.000 326.200 542.800 337.800 ;
        RECT 543.600 324.200 544.400 337.800 ;
        RECT 545.200 324.200 546.000 337.800 ;
        RECT 546.900 332.400 547.500 339.700 ;
        RECT 550.100 336.400 550.700 403.600 ;
        RECT 566.100 402.400 566.700 415.600 ;
        RECT 567.600 406.200 568.400 417.800 ;
        RECT 569.200 413.600 570.000 414.400 ;
        RECT 570.800 406.200 571.600 417.800 ;
        RECT 572.400 404.200 573.200 417.800 ;
        RECT 574.000 404.200 574.800 417.800 ;
        RECT 580.400 413.600 581.200 414.400 ;
        RECT 551.600 401.600 552.400 402.400 ;
        RECT 562.800 401.600 563.600 402.400 ;
        RECT 566.000 401.600 566.800 402.400 ;
        RECT 551.700 390.400 552.300 401.600 ;
        RECT 551.600 389.600 552.400 390.400 ;
        RECT 551.700 372.400 552.300 389.600 ;
        RECT 554.800 384.200 555.600 397.800 ;
        RECT 556.400 384.200 557.200 397.800 ;
        RECT 558.000 384.200 558.800 395.800 ;
        RECT 559.600 387.600 560.400 388.400 ;
        RECT 561.200 384.200 562.000 395.800 ;
        RECT 562.900 386.400 563.500 401.600 ;
        RECT 562.800 385.600 563.600 386.400 ;
        RECT 562.900 382.300 563.500 385.600 ;
        RECT 564.400 384.200 565.200 395.800 ;
        RECT 566.000 384.200 566.800 397.800 ;
        RECT 567.600 384.200 568.400 397.800 ;
        RECT 569.200 384.200 570.000 397.800 ;
        RECT 578.800 383.600 579.600 384.400 ;
        RECT 562.900 381.700 565.100 382.300 ;
        RECT 551.600 371.600 552.400 372.400 ;
        RECT 551.700 350.400 552.300 371.600 ;
        RECT 556.400 364.200 557.200 377.800 ;
        RECT 558.000 364.200 558.800 377.800 ;
        RECT 559.600 366.200 560.400 377.800 ;
        RECT 561.200 373.600 562.000 374.400 ;
        RECT 562.800 366.200 563.600 377.800 ;
        RECT 564.500 376.400 565.100 381.700 ;
        RECT 564.400 375.600 565.200 376.400 ;
        RECT 564.500 364.300 565.100 375.600 ;
        RECT 566.000 366.200 566.800 377.800 ;
        RECT 564.500 363.700 566.700 364.300 ;
        RECT 567.600 364.200 568.400 377.800 ;
        RECT 569.200 364.200 570.000 377.800 ;
        RECT 570.800 364.200 571.600 377.800 ;
        RECT 578.900 374.400 579.500 383.600 ;
        RECT 580.500 378.400 581.100 413.600 ;
        RECT 580.400 377.600 581.200 378.400 ;
        RECT 578.800 373.600 579.600 374.400 ;
        RECT 551.600 349.600 552.400 350.400 ;
        RECT 553.200 349.600 554.000 350.400 ;
        RECT 550.000 335.600 550.800 336.400 ;
        RECT 553.300 334.400 553.900 349.600 ;
        RECT 558.000 344.200 558.800 357.800 ;
        RECT 559.600 344.200 560.400 357.800 ;
        RECT 561.200 344.200 562.000 355.800 ;
        RECT 562.800 347.600 563.600 348.400 ;
        RECT 564.400 344.200 565.200 355.800 ;
        RECT 566.100 346.400 566.700 363.700 ;
        RECT 566.000 345.600 566.800 346.400 ;
        RECT 566.100 340.400 566.700 345.600 ;
        RECT 567.600 344.200 568.400 355.800 ;
        RECT 569.200 344.200 570.000 357.800 ;
        RECT 570.800 344.200 571.600 357.800 ;
        RECT 572.400 344.200 573.200 357.800 ;
        RECT 578.800 343.600 579.600 344.400 ;
        RECT 582.000 343.600 582.800 344.400 ;
        RECT 566.000 339.600 566.800 340.400 ;
        RECT 553.200 333.600 554.000 334.400 ;
        RECT 546.800 331.600 547.600 332.400 ;
        RECT 497.200 317.600 498.000 318.400 ;
        RECT 500.400 317.600 501.200 318.400 ;
        RECT 487.600 307.600 488.400 308.400 ;
        RECT 486.100 305.700 488.300 306.300 ;
        RECT 454.000 291.600 454.800 292.400 ;
        RECT 434.800 289.400 435.600 290.200 ;
        RECT 441.400 289.400 442.200 290.200 ;
        RECT 452.400 289.600 453.200 290.400 ;
        RECT 436.400 285.600 437.200 286.400 ;
        RECT 455.700 278.400 456.300 303.600 ;
        RECT 462.100 294.400 462.700 303.600 ;
        RECT 487.700 298.400 488.300 305.700 ;
        RECT 492.400 304.200 493.200 315.800 ;
        RECT 500.400 305.600 501.200 306.400 ;
        RECT 510.000 304.200 510.800 317.800 ;
        RECT 511.600 304.200 512.400 317.800 ;
        RECT 513.200 304.200 514.000 317.800 ;
        RECT 514.800 304.200 515.600 315.800 ;
        RECT 516.400 307.600 517.200 308.400 ;
        RECT 516.500 306.400 517.100 307.600 ;
        RECT 516.400 305.600 517.200 306.400 ;
        RECT 457.200 293.600 458.000 294.400 ;
        RECT 458.800 293.600 459.600 294.400 ;
        RECT 462.000 293.600 462.800 294.400 ;
        RECT 460.400 291.600 461.200 292.400 ;
        RECT 462.000 291.600 462.800 292.400 ;
        RECT 457.200 289.600 458.000 290.400 ;
        RECT 457.300 288.400 457.900 289.600 ;
        RECT 457.200 287.600 458.000 288.400 ;
        RECT 460.400 287.600 461.200 288.400 ;
        RECT 462.100 278.400 462.700 291.600 ;
        RECT 463.600 289.600 464.400 290.400 ;
        RECT 465.200 290.200 466.000 295.800 ;
        RECT 466.800 293.600 467.600 294.400 ;
        RECT 455.600 277.600 456.400 278.400 ;
        RECT 462.000 277.600 462.800 278.400 ;
        RECT 426.800 269.400 427.600 270.200 ;
        RECT 428.400 264.200 429.200 275.800 ;
        RECT 433.200 273.600 434.000 274.400 ;
        RECT 430.000 267.600 430.800 268.400 ;
        RECT 423.600 246.200 424.400 257.800 ;
        RECT 430.100 254.400 430.700 267.600 ;
        RECT 431.600 266.200 432.400 271.800 ;
        RECT 433.300 270.400 433.900 273.600 ;
        RECT 438.000 271.600 438.800 272.400 ;
        RECT 451.000 271.800 451.800 272.600 ;
        RECT 457.200 271.800 458.000 272.600 ;
        RECT 433.200 269.600 434.000 270.400 ;
        RECT 439.600 269.600 440.400 270.400 ;
        RECT 444.400 269.600 445.200 270.400 ;
        RECT 442.800 268.300 443.600 268.400 ;
        RECT 441.300 267.700 443.600 268.300 ;
        RECT 436.400 265.600 437.200 266.400 ;
        RECT 434.800 263.600 435.600 264.400 ;
        RECT 434.900 260.400 435.500 263.600 ;
        RECT 434.800 259.600 435.600 260.400 ;
        RECT 431.600 257.600 432.400 258.400 ;
        RECT 436.500 258.300 437.100 265.600 ;
        RECT 439.600 259.600 440.400 260.400 ;
        RECT 430.000 253.600 430.800 254.400 ;
        RECT 431.700 252.600 432.300 257.600 ;
        RECT 431.600 251.800 432.400 252.600 ;
        RECT 433.200 246.200 434.000 257.800 ;
        RECT 434.900 257.700 437.100 258.300 ;
        RECT 433.200 237.600 434.000 238.400 ;
        RECT 425.200 235.600 426.000 236.400 ;
        RECT 422.000 233.600 422.800 234.400 ;
        RECT 425.300 232.400 425.900 235.600 ;
        RECT 430.000 233.600 430.800 234.400 ;
        RECT 425.200 231.600 426.000 232.400 ;
        RECT 430.100 230.400 430.700 233.600 ;
        RECT 430.000 229.600 430.800 230.400 ;
        RECT 434.900 230.300 435.500 257.700 ;
        RECT 436.400 250.200 437.200 255.800 ;
        RECT 439.700 254.400 440.300 259.600 ;
        RECT 441.300 258.400 441.900 267.700 ;
        RECT 442.800 267.600 443.600 267.700 ;
        RECT 444.500 264.400 445.100 269.600 ;
        RECT 449.200 267.600 450.000 268.400 ;
        RECT 444.400 263.600 445.200 264.400 ;
        RECT 441.200 257.600 442.000 258.400 ;
        RECT 442.800 255.600 443.600 256.400 ;
        RECT 439.600 253.600 440.400 254.400 ;
        RECT 438.000 251.600 438.800 252.400 ;
        RECT 441.200 251.600 442.000 252.400 ;
        RECT 439.600 243.600 440.400 244.400 ;
        RECT 439.700 238.400 440.300 243.600 ;
        RECT 439.600 237.600 440.400 238.400 ;
        RECT 441.300 234.400 441.900 251.600 ;
        RECT 442.900 250.400 443.500 255.600 ;
        RECT 442.800 249.600 443.600 250.400 ;
        RECT 449.300 246.400 449.900 267.600 ;
        RECT 451.000 267.000 451.600 271.800 ;
        RECT 452.200 269.800 453.000 270.600 ;
        RECT 452.400 268.400 453.000 269.800 ;
        RECT 457.400 268.400 458.000 271.800 ;
        RECT 463.600 271.600 464.400 272.400 ;
        RECT 460.400 269.600 461.200 270.400 ;
        RECT 460.500 268.400 461.100 269.600 ;
        RECT 452.400 267.800 458.000 268.400 ;
        RECT 452.400 267.000 453.200 267.200 ;
        RECT 455.800 267.000 456.600 267.200 ;
        RECT 457.400 267.000 458.000 267.800 ;
        RECT 458.800 267.600 459.600 268.400 ;
        RECT 460.400 267.600 461.200 268.400 ;
        RECT 451.000 266.400 456.600 267.000 ;
        RECT 451.000 266.200 451.800 266.400 ;
        RECT 457.200 266.200 458.000 267.000 ;
        RECT 457.200 263.600 458.000 264.400 ;
        RECT 452.400 259.600 453.200 260.400 ;
        RECT 452.500 252.400 453.100 259.600 ;
        RECT 457.300 258.400 457.900 263.600 ;
        RECT 458.900 260.400 459.500 267.600 ;
        RECT 458.800 259.600 459.600 260.400 ;
        RECT 463.700 258.400 464.300 271.600 ;
        RECT 465.200 266.200 466.000 271.800 ;
        RECT 466.900 268.400 467.500 293.600 ;
        RECT 468.400 286.200 469.200 297.800 ;
        RECT 470.000 291.600 470.800 292.600 ;
        RECT 478.000 286.200 478.800 297.800 ;
        RECT 487.600 297.600 488.400 298.400 ;
        RECT 486.000 295.000 486.800 295.800 ;
        RECT 487.400 295.000 491.600 295.600 ;
        RECT 492.600 295.000 493.400 295.800 ;
        RECT 484.400 293.600 485.200 294.400 ;
        RECT 486.000 294.200 486.600 295.000 ;
        RECT 487.400 294.800 488.200 295.000 ;
        RECT 490.800 294.800 491.600 295.000 ;
        RECT 486.000 293.600 490.800 294.200 ;
        RECT 482.800 287.600 483.600 288.400 ;
        RECT 466.800 267.600 467.600 268.400 ;
        RECT 468.400 264.200 469.200 275.800 ;
        RECT 470.000 269.400 470.800 270.200 ;
        RECT 457.200 257.600 458.000 258.400 ;
        RECT 463.600 257.600 464.400 258.400 ;
        RECT 458.800 255.600 459.600 256.400 ;
        RECT 468.400 255.600 469.200 256.400 ;
        RECT 450.800 251.600 451.600 252.400 ;
        RECT 452.400 251.600 453.200 252.400 ;
        RECT 455.600 251.600 456.400 252.400 ;
        RECT 458.900 252.300 459.500 255.600 ;
        RECT 468.500 254.400 469.100 255.600 ;
        RECT 462.000 253.600 462.800 254.400 ;
        RECT 465.200 253.600 466.000 254.400 ;
        RECT 468.400 253.600 469.200 254.400 ;
        RECT 460.400 252.300 461.200 252.400 ;
        RECT 458.900 251.700 461.200 252.300 ;
        RECT 460.400 251.600 461.200 251.700 ;
        RECT 450.900 248.400 451.500 251.600 ;
        RECT 454.000 249.600 454.800 250.400 ;
        RECT 455.700 248.400 456.300 251.600 ;
        RECT 460.500 248.400 461.100 251.600 ;
        RECT 450.800 247.600 451.600 248.400 ;
        RECT 452.400 247.600 453.200 248.400 ;
        RECT 455.600 247.600 456.400 248.400 ;
        RECT 460.400 247.600 461.200 248.400 ;
        RECT 452.500 246.400 453.100 247.600 ;
        RECT 449.200 245.600 450.000 246.400 ;
        RECT 452.400 245.600 453.200 246.400 ;
        RECT 450.800 241.600 451.600 242.400 ;
        RECT 450.900 238.400 451.500 241.600 ;
        RECT 455.700 240.400 456.300 247.600 ;
        RECT 455.600 239.600 456.400 240.400 ;
        RECT 450.800 237.600 451.600 238.400 ;
        RECT 462.100 236.400 462.700 253.600 ;
        RECT 465.300 238.400 465.900 253.600 ;
        RECT 466.800 251.600 467.600 252.400 ;
        RECT 468.400 249.600 469.200 250.400 ;
        RECT 470.100 250.300 470.700 269.400 ;
        RECT 478.000 264.200 478.800 275.800 ;
        RECT 484.500 274.400 485.100 293.600 ;
        RECT 486.000 290.200 486.600 293.600 ;
        RECT 490.000 293.400 490.800 293.600 ;
        RECT 490.800 291.600 491.600 292.400 ;
        RECT 486.000 289.400 486.800 290.200 ;
        RECT 479.600 273.600 480.400 274.400 ;
        RECT 482.800 273.600 483.600 274.400 ;
        RECT 484.400 273.600 485.200 274.400 ;
        RECT 471.600 251.600 472.400 252.400 ;
        RECT 474.800 251.600 475.600 252.400 ;
        RECT 470.100 249.700 472.300 250.300 ;
        RECT 468.400 245.600 469.200 246.400 ;
        RECT 466.800 239.600 467.600 240.400 ;
        RECT 465.200 237.600 466.000 238.400 ;
        RECT 462.000 235.600 462.800 236.400 ;
        RECT 441.200 233.600 442.000 234.400 ;
        RECT 442.800 233.600 443.600 234.400 ;
        RECT 455.600 233.600 456.400 234.400 ;
        RECT 438.000 231.600 438.800 232.400 ;
        RECT 436.400 230.300 437.200 230.400 ;
        RECT 434.900 229.700 437.200 230.300 ;
        RECT 436.400 229.600 437.200 229.700 ;
        RECT 436.500 226.400 437.100 229.600 ;
        RECT 434.800 225.600 435.600 226.400 ;
        RECT 436.400 225.600 437.200 226.400 ;
        RECT 428.400 223.600 429.200 224.400 ;
        RECT 414.100 221.700 416.300 222.300 ;
        RECT 364.400 218.300 365.200 218.400 ;
        RECT 345.200 211.600 346.000 212.400 ;
        RECT 346.800 210.200 347.600 215.800 ;
        RECT 348.400 213.600 349.200 214.400 ;
        RECT 350.000 206.200 350.800 217.800 ;
        RECT 351.600 211.800 352.400 212.600 ;
        RECT 351.700 198.400 352.300 211.800 ;
        RECT 358.000 211.600 358.800 212.400 ;
        RECT 326.000 197.600 326.800 198.400 ;
        RECT 351.600 197.600 352.400 198.400 ;
        RECT 306.800 193.600 307.600 194.400 ;
        RECT 321.200 193.600 322.000 194.400 ;
        RECT 321.300 192.400 321.900 193.600 ;
        RECT 311.600 191.600 312.400 192.400 ;
        RECT 321.200 191.600 322.000 192.400 ;
        RECT 324.200 191.800 325.000 192.600 ;
        RECT 330.800 191.800 331.600 192.600 ;
        RECT 314.800 189.600 315.600 190.400 ;
        RECT 308.400 187.600 309.200 188.400 ;
        RECT 310.000 187.600 310.800 188.400 ;
        RECT 313.200 187.600 314.000 188.400 ;
        RECT 310.100 186.400 310.700 187.600 ;
        RECT 313.300 186.400 313.900 187.600 ;
        RECT 310.000 185.600 310.800 186.400 ;
        RECT 313.200 185.600 314.000 186.400 ;
        RECT 308.400 177.600 309.200 178.400 ;
        RECT 310.100 170.400 310.700 185.600 ;
        RECT 314.900 184.400 315.500 189.600 ;
        RECT 318.000 187.600 318.800 188.400 ;
        RECT 322.800 187.600 323.600 188.400 ;
        RECT 314.800 184.300 315.600 184.400 ;
        RECT 314.800 183.700 317.100 184.300 ;
        RECT 314.800 183.600 315.600 183.700 ;
        RECT 313.200 177.600 314.000 178.400 ;
        RECT 313.300 174.400 313.900 177.600 ;
        RECT 313.200 173.600 314.000 174.400 ;
        RECT 316.500 172.400 317.100 183.700 ;
        RECT 316.400 171.600 317.200 172.400 ;
        RECT 318.100 170.400 318.700 187.600 ;
        RECT 322.900 186.400 323.500 187.600 ;
        RECT 324.200 187.000 324.800 191.800 ;
        RECT 326.800 188.400 327.600 188.600 ;
        RECT 331.000 188.400 331.600 191.800 ;
        RECT 338.800 191.600 339.600 192.400 ;
        RECT 343.600 191.600 344.400 192.400 ;
        RECT 346.800 191.800 347.600 192.600 ;
        RECT 353.400 191.800 354.200 192.600 ;
        RECT 335.600 189.600 336.400 190.400 ;
        RECT 326.800 187.800 331.600 188.400 ;
        RECT 326.000 187.000 326.800 187.200 ;
        RECT 329.400 187.000 330.200 187.200 ;
        RECT 331.000 187.000 331.600 187.800 ;
        RECT 332.400 187.600 333.200 188.400 ;
        RECT 322.800 185.600 323.600 186.400 ;
        RECT 324.200 186.200 325.000 187.000 ;
        RECT 326.000 186.400 330.200 187.000 ;
        RECT 330.800 186.200 331.600 187.000 ;
        RECT 332.400 185.600 333.200 186.400 ;
        RECT 321.200 183.600 322.000 184.400 ;
        RECT 321.300 176.400 321.900 183.600 ;
        RECT 326.000 179.600 326.800 180.400 ;
        RECT 326.100 178.400 326.700 179.600 ;
        RECT 326.000 177.600 326.800 178.400 ;
        RECT 332.500 176.400 333.100 185.600 ;
        RECT 335.700 184.400 336.300 189.600 ;
        RECT 335.600 183.600 336.400 184.400 ;
        RECT 321.200 175.600 322.000 176.400 ;
        RECT 332.400 175.600 333.200 176.400 ;
        RECT 321.200 173.600 322.000 174.400 ;
        RECT 324.400 173.600 325.200 174.400 ;
        RECT 330.800 173.600 331.600 174.400 ;
        RECT 319.600 171.600 320.400 172.400 ;
        RECT 319.700 170.400 320.300 171.600 ;
        RECT 321.300 170.400 321.900 173.600 ;
        RECT 310.000 169.600 310.800 170.400 ;
        RECT 318.000 169.600 318.800 170.400 ;
        RECT 319.600 169.600 320.400 170.400 ;
        RECT 321.200 169.600 322.000 170.400 ;
        RECT 326.000 169.600 326.800 170.400 ;
        RECT 305.200 167.600 306.000 168.400 ;
        RECT 247.600 163.600 248.400 164.400 ;
        RECT 250.800 163.600 251.600 164.400 ;
        RECT 244.400 157.600 245.200 158.400 ;
        RECT 188.400 155.600 189.200 156.400 ;
        RECT 239.600 153.600 240.400 154.400 ;
        RECT 188.200 151.800 189.000 152.600 ;
        RECT 194.800 151.800 195.600 152.600 ;
        RECT 188.200 147.000 188.800 151.800 ;
        RECT 190.800 148.400 191.600 148.600 ;
        RECT 195.000 148.400 195.600 151.800 ;
        RECT 199.800 151.800 200.600 152.600 ;
        RECT 206.000 151.800 206.800 152.600 ;
        RECT 190.800 147.800 195.600 148.400 ;
        RECT 190.000 147.000 190.800 147.200 ;
        RECT 193.400 147.000 194.200 147.200 ;
        RECT 195.000 147.000 195.600 147.800 ;
        RECT 196.400 147.600 197.200 148.400 ;
        RECT 198.000 147.600 198.800 148.400 ;
        RECT 188.200 146.200 189.000 147.000 ;
        RECT 190.000 146.400 194.200 147.000 ;
        RECT 183.600 141.600 184.400 142.400 ;
        RECT 170.800 131.600 171.600 132.400 ;
        RECT 172.400 126.200 173.200 137.800 ;
        RECT 188.400 135.600 189.200 136.400 ;
        RECT 178.800 133.600 179.600 134.400 ;
        RECT 183.600 133.600 184.400 134.400 ;
        RECT 182.000 131.600 182.800 132.400 ;
        RECT 182.100 130.400 182.700 131.600 ;
        RECT 182.000 129.600 182.800 130.400 ;
        RECT 174.000 127.600 174.800 128.400 ;
        RECT 153.200 107.800 158.800 108.400 ;
        RECT 153.200 107.000 154.000 107.200 ;
        RECT 156.600 107.000 157.400 107.200 ;
        RECT 158.200 107.000 158.800 107.800 ;
        RECT 159.600 107.600 160.400 108.400 ;
        RECT 151.800 106.400 157.400 107.000 ;
        RECT 143.600 105.600 144.400 106.400 ;
        RECT 145.200 105.600 146.000 106.400 ;
        RECT 150.000 105.600 150.800 106.400 ;
        RECT 151.800 106.200 152.600 106.400 ;
        RECT 158.000 106.200 158.800 107.000 ;
        RECT 159.700 106.400 160.300 107.600 ;
        RECT 159.600 105.600 160.400 106.400 ;
        RECT 162.800 105.600 163.600 106.400 ;
        RECT 164.400 106.200 165.200 111.800 ;
        RECT 153.200 103.600 154.000 104.400 ;
        RECT 167.600 104.200 168.400 115.800 ;
        RECT 169.200 113.600 170.000 114.400 ;
        RECT 169.300 110.200 169.900 113.600 ;
        RECT 174.100 110.400 174.700 127.600 ;
        RECT 177.200 123.600 178.000 124.400 ;
        RECT 177.300 120.400 177.900 123.600 ;
        RECT 177.200 119.600 178.000 120.400 ;
        RECT 169.200 109.400 170.000 110.200 ;
        RECT 174.000 109.600 174.800 110.400 ;
        RECT 169.200 105.600 170.000 106.400 ;
        RECT 146.800 101.600 147.600 102.400 ;
        RECT 146.900 98.400 147.500 101.600 ;
        RECT 145.200 97.600 146.000 98.400 ;
        RECT 146.800 97.600 147.600 98.400 ;
        RECT 145.300 94.400 145.900 97.600 ;
        RECT 145.200 93.600 146.000 94.400 ;
        RECT 153.300 92.400 153.900 103.600 ;
        RECT 156.400 93.600 157.200 94.400 ;
        RECT 145.200 91.600 146.000 92.400 ;
        RECT 150.000 91.600 150.800 92.400 ;
        RECT 153.200 91.600 154.000 92.400 ;
        RECT 145.300 90.400 145.900 91.600 ;
        RECT 150.100 90.400 150.700 91.600 ;
        RECT 153.300 90.400 153.900 91.600 ;
        RECT 145.200 89.600 146.000 90.400 ;
        RECT 146.800 89.600 147.600 90.400 ;
        RECT 150.000 89.600 150.800 90.400 ;
        RECT 153.200 89.600 154.000 90.400 ;
        RECT 146.900 88.400 147.500 89.600 ;
        RECT 146.800 87.600 147.600 88.400 ;
        RECT 156.500 86.400 157.100 93.600 ;
        RECT 158.000 90.200 158.800 95.800 ;
        RECT 156.400 85.600 157.200 86.400 ;
        RECT 161.200 86.200 162.000 97.800 ;
        RECT 162.800 93.600 163.600 94.400 ;
        RECT 166.000 93.600 166.800 94.400 ;
        RECT 162.900 92.600 163.500 93.600 ;
        RECT 162.800 91.800 163.600 92.600 ;
        RECT 143.600 83.600 144.400 84.400 ;
        RECT 143.700 70.400 144.300 83.600 ;
        RECT 145.200 71.800 146.000 72.600 ;
        RECT 151.800 71.800 152.600 72.600 ;
        RECT 142.000 69.600 142.800 70.400 ;
        RECT 143.600 69.600 144.400 70.400 ;
        RECT 145.200 68.400 145.800 71.800 ;
        RECT 149.200 68.400 150.000 68.600 ;
        RECT 130.800 67.600 131.600 68.400 ;
        RECT 134.000 67.600 134.800 68.400 ;
        RECT 137.200 67.600 138.000 68.400 ;
        RECT 143.600 67.600 144.400 68.400 ;
        RECT 145.200 67.800 150.000 68.400 ;
        RECT 127.600 59.600 128.400 60.400 ;
        RECT 129.200 59.600 130.000 60.400 ;
        RECT 126.000 53.600 126.800 54.400 ;
        RECT 127.700 52.400 128.300 59.600 ;
        RECT 132.400 57.600 133.200 58.400 ;
        RECT 132.500 56.400 133.100 57.600 ;
        RECT 130.800 55.600 131.600 56.400 ;
        RECT 132.400 55.600 133.200 56.400 ;
        RECT 129.200 53.600 130.000 54.400 ;
        RECT 124.500 51.700 126.700 52.300 ;
        RECT 114.900 50.400 115.500 51.600 ;
        RECT 105.200 49.600 106.000 50.400 ;
        RECT 114.800 49.600 115.600 50.400 ;
        RECT 124.400 49.600 125.200 50.400 ;
        RECT 76.400 47.600 77.200 48.400 ;
        RECT 100.400 47.600 101.200 48.400 ;
        RECT 87.600 45.600 88.400 46.400 ;
        RECT 73.200 43.600 74.000 44.400 ;
        RECT 81.200 43.600 82.000 44.400 ;
        RECT 73.300 38.400 73.900 43.600 ;
        RECT 73.200 37.600 74.000 38.400 ;
        RECT 70.000 33.600 70.800 34.400 ;
        RECT 68.400 27.600 69.200 28.400 ;
        RECT 14.000 25.600 14.800 26.400 ;
        RECT 17.200 25.600 18.000 26.400 ;
        RECT 28.400 25.600 29.200 26.400 ;
        RECT 41.200 25.600 42.000 26.400 ;
        RECT 46.000 25.600 46.800 26.400 ;
        RECT 49.200 25.600 50.000 26.400 ;
        RECT 57.200 25.600 58.000 26.400 ;
        RECT 60.400 26.200 61.200 27.000 ;
        RECT 61.800 26.400 66.000 27.000 ;
        RECT 67.000 26.200 67.800 27.000 ;
        RECT 70.000 26.200 70.800 31.800 ;
        RECT 15.600 23.600 16.400 24.400 ;
        RECT 20.400 23.600 21.200 24.400 ;
        RECT 15.700 16.300 16.300 23.600 ;
        RECT 20.500 18.400 21.100 23.600 ;
        RECT 20.400 17.600 21.200 18.400 ;
        RECT 14.100 15.700 16.300 16.300 ;
        RECT 14.100 12.400 14.700 15.700 ;
        RECT 18.800 15.000 19.600 15.800 ;
        RECT 20.200 15.000 24.400 15.600 ;
        RECT 25.400 15.000 26.200 15.800 ;
        RECT 15.600 13.600 16.400 14.400 ;
        RECT 17.200 13.600 18.000 14.400 ;
        RECT 18.800 14.200 19.400 15.000 ;
        RECT 20.200 14.800 21.000 15.000 ;
        RECT 23.600 14.800 24.400 15.000 ;
        RECT 18.800 13.600 23.600 14.200 ;
        RECT 12.400 11.600 13.200 12.400 ;
        RECT 14.000 11.600 14.800 12.400 ;
        RECT 15.700 10.400 16.300 13.600 ;
        RECT 9.200 9.600 10.000 10.400 ;
        RECT 10.800 9.600 11.600 10.400 ;
        RECT 15.600 9.600 16.400 10.400 ;
        RECT 18.800 10.200 19.400 13.600 ;
        RECT 22.800 13.400 23.600 13.600 ;
        RECT 25.600 10.200 26.200 15.000 ;
        RECT 28.500 14.400 29.100 25.600 ;
        RECT 34.800 23.600 35.600 24.400 ;
        RECT 34.900 20.400 35.500 23.600 ;
        RECT 34.800 19.600 35.600 20.400 ;
        RECT 57.300 18.400 57.900 25.600 ;
        RECT 65.200 23.600 66.000 24.400 ;
        RECT 73.200 24.200 74.000 35.800 ;
        RECT 76.400 31.600 77.200 32.400 ;
        RECT 76.500 30.400 77.100 31.600 ;
        RECT 81.300 30.400 81.900 43.600 ;
        RECT 87.700 38.400 88.300 45.600 ;
        RECT 92.400 43.600 93.200 44.400 ;
        RECT 102.000 43.600 102.800 44.400 ;
        RECT 87.600 37.600 88.400 38.400 ;
        RECT 76.400 29.600 77.200 30.400 ;
        RECT 79.600 29.600 80.400 30.400 ;
        RECT 81.200 29.600 82.000 30.400 ;
        RECT 76.400 19.600 77.200 20.400 ;
        RECT 76.500 18.400 77.100 19.600 ;
        RECT 38.000 17.600 38.800 18.400 ;
        RECT 30.000 15.000 30.800 15.800 ;
        RECT 31.400 15.000 35.600 15.600 ;
        RECT 36.600 15.000 37.400 15.800 ;
        RECT 26.800 13.600 27.600 14.400 ;
        RECT 28.400 13.600 29.200 14.400 ;
        RECT 30.000 14.200 30.600 15.000 ;
        RECT 31.400 14.800 32.200 15.000 ;
        RECT 34.800 14.800 35.600 15.000 ;
        RECT 30.000 13.600 34.800 14.200 ;
        RECT 26.900 12.400 27.500 13.600 ;
        RECT 26.800 11.600 27.600 12.400 ;
        RECT 10.900 8.400 11.500 9.600 ;
        RECT 18.800 9.400 19.600 10.200 ;
        RECT 25.400 9.400 26.200 10.200 ;
        RECT 30.000 10.200 30.600 13.600 ;
        RECT 34.000 13.400 34.800 13.600 ;
        RECT 30.000 9.400 30.800 10.200 ;
        RECT 34.800 9.600 35.600 10.400 ;
        RECT 36.800 10.200 37.400 15.000 ;
        RECT 38.100 14.400 38.700 17.600 ;
        RECT 38.000 13.600 38.800 14.400 ;
        RECT 39.600 10.200 40.400 15.800 ;
        RECT 34.900 8.400 35.500 9.600 ;
        RECT 36.600 9.400 37.400 10.200 ;
        RECT 6.000 7.600 6.800 8.400 ;
        RECT 7.600 7.600 8.400 8.400 ;
        RECT 10.800 7.600 11.600 8.400 ;
        RECT 23.600 7.600 24.400 8.400 ;
        RECT 34.800 7.600 35.600 8.400 ;
        RECT 7.700 6.400 8.300 7.600 ;
        RECT 7.600 5.600 8.400 6.400 ;
        RECT 42.800 6.200 43.600 17.800 ;
        RECT 44.400 11.800 45.200 12.600 ;
        RECT 44.500 8.400 45.100 11.800 ;
        RECT 50.800 11.600 51.600 12.400 ;
        RECT 44.400 7.600 45.200 8.400 ;
        RECT 52.400 6.200 53.200 17.800 ;
        RECT 57.200 17.600 58.000 18.400 ;
        RECT 58.800 10.200 59.600 15.800 ;
        RECT 60.400 13.600 61.200 14.400 ;
        RECT 60.500 12.400 61.100 13.600 ;
        RECT 60.400 11.600 61.200 12.400 ;
        RECT 62.000 6.200 62.800 17.800 ;
        RECT 63.600 11.600 64.400 12.600 ;
        RECT 70.000 11.600 70.800 12.400 ;
        RECT 71.600 6.200 72.400 17.800 ;
        RECT 76.400 17.600 77.200 18.400 ;
        RECT 78.000 10.200 78.800 15.800 ;
        RECT 79.700 14.400 80.300 29.600 ;
        RECT 82.800 24.200 83.600 35.800 ;
        RECT 90.600 31.800 91.400 32.600 ;
        RECT 92.500 32.400 93.100 43.600 ;
        RECT 98.800 37.600 99.600 38.400 ;
        RECT 89.200 27.600 90.000 28.400 ;
        RECT 90.600 27.000 91.200 31.800 ;
        RECT 92.400 31.600 93.200 32.400 ;
        RECT 97.200 31.800 98.000 32.600 ;
        RECT 93.200 28.400 94.000 28.600 ;
        RECT 97.400 28.400 98.000 31.800 ;
        RECT 98.900 28.400 99.500 37.600 ;
        RECT 100.400 32.300 101.200 32.400 ;
        RECT 102.100 32.300 102.700 43.600 ;
        RECT 103.600 33.600 104.400 34.400 ;
        RECT 100.400 31.700 102.700 32.300 ;
        RECT 100.400 31.600 101.200 31.700 ;
        RECT 103.700 30.400 104.300 33.600 ;
        RECT 100.400 29.600 101.200 30.400 ;
        RECT 103.600 29.600 104.400 30.400 ;
        RECT 105.300 28.400 105.900 49.600 ;
        RECT 124.500 48.400 125.100 49.600 ;
        RECT 124.400 47.600 125.200 48.400 ;
        RECT 93.200 27.800 98.000 28.400 ;
        RECT 92.400 27.000 93.200 27.200 ;
        RECT 95.800 27.000 96.600 27.200 ;
        RECT 97.400 27.000 98.000 27.800 ;
        RECT 98.800 27.600 99.600 28.400 ;
        RECT 100.400 27.600 101.200 28.400 ;
        RECT 105.200 27.600 106.000 28.400 ;
        RECT 90.600 26.200 91.400 27.000 ;
        RECT 92.400 26.400 96.600 27.000 ;
        RECT 97.200 26.200 98.000 27.000 ;
        RECT 106.800 26.200 107.600 31.800 ;
        RECT 108.400 27.600 109.200 28.400 ;
        RECT 102.000 23.600 102.800 24.400 ;
        RECT 79.600 13.600 80.400 14.400 ;
        RECT 81.200 6.200 82.000 17.800 ;
        RECT 82.800 11.800 83.600 12.600 ;
        RECT 82.900 10.400 83.500 11.800 ;
        RECT 89.200 11.600 90.000 12.400 ;
        RECT 82.800 9.600 83.600 10.400 ;
        RECT 90.800 6.200 91.600 17.800 ;
        RECT 95.600 17.600 96.400 18.400 ;
        RECT 97.200 10.200 98.000 15.800 ;
        RECT 98.800 13.600 99.600 14.400 ;
        RECT 98.900 12.400 99.500 13.600 ;
        RECT 98.800 11.600 99.600 12.400 ;
        RECT 100.400 6.200 101.200 17.800 ;
        RECT 102.100 12.600 102.700 23.600 ;
        RECT 102.000 11.800 102.800 12.600 ;
        RECT 108.500 12.400 109.100 27.600 ;
        RECT 110.000 24.200 110.800 35.800 ;
        RECT 118.000 31.600 118.800 32.400 ;
        RECT 118.100 30.400 118.700 31.600 ;
        RECT 111.600 29.400 112.400 30.400 ;
        RECT 118.000 29.600 118.800 30.400 ;
        RECT 108.400 11.600 109.200 12.400 ;
        RECT 110.000 6.200 110.800 17.800 ;
        RECT 114.800 17.600 115.600 18.400 ;
        RECT 116.400 10.200 117.200 15.800 ;
        RECT 118.100 14.400 118.700 29.600 ;
        RECT 119.600 24.200 120.400 35.800 ;
        RECT 126.100 28.400 126.700 51.700 ;
        RECT 127.600 51.600 128.400 52.400 ;
        RECT 129.300 50.400 129.900 53.600 ;
        RECT 129.200 49.600 130.000 50.400 ;
        RECT 130.800 43.600 131.600 44.400 ;
        RECT 134.100 44.300 134.700 67.600 ;
        RECT 143.700 64.400 144.300 67.600 ;
        RECT 145.200 67.000 145.800 67.800 ;
        RECT 146.600 67.000 147.400 67.200 ;
        RECT 150.000 67.000 150.800 67.200 ;
        RECT 152.000 67.000 152.600 71.800 ;
        RECT 153.200 67.600 154.000 68.400 ;
        RECT 145.200 66.200 146.000 67.000 ;
        RECT 146.600 66.400 150.800 67.000 ;
        RECT 151.800 66.200 152.600 67.000 ;
        RECT 153.300 66.400 153.900 67.600 ;
        RECT 153.200 65.600 154.000 66.400 ;
        RECT 154.800 66.200 155.600 71.800 ;
        RECT 143.600 63.600 144.400 64.400 ;
        RECT 146.800 63.600 147.600 64.400 ;
        RECT 153.200 63.600 154.000 64.400 ;
        RECT 146.900 62.400 147.500 63.600 ;
        RECT 140.400 61.600 141.200 62.400 ;
        RECT 146.800 61.600 147.600 62.400 ;
        RECT 148.400 61.600 149.200 62.400 ;
        RECT 140.500 52.400 141.100 61.600 ;
        RECT 143.600 57.600 144.400 58.400 ;
        RECT 146.800 55.600 147.600 56.400 ;
        RECT 146.900 52.400 147.500 55.600 ;
        RECT 140.400 51.600 141.200 52.400 ;
        RECT 146.800 51.600 147.600 52.400 ;
        RECT 132.500 43.700 134.700 44.300 ;
        RECT 130.900 34.400 131.500 43.600 ;
        RECT 130.800 33.600 131.600 34.400 ;
        RECT 127.600 31.800 128.400 32.600 ;
        RECT 127.600 28.400 128.200 31.800 ;
        RECT 132.500 30.400 133.100 43.700 ;
        RECT 140.400 35.600 141.200 36.400 ;
        RECT 134.200 31.800 135.000 32.600 ;
        RECT 132.400 29.600 133.200 30.400 ;
        RECT 131.600 28.400 132.400 28.600 ;
        RECT 126.000 27.600 126.800 28.400 ;
        RECT 127.600 27.800 132.400 28.400 ;
        RECT 127.600 27.000 128.200 27.800 ;
        RECT 129.000 27.000 129.800 27.200 ;
        RECT 132.400 27.000 133.200 27.200 ;
        RECT 134.400 27.000 135.000 31.800 ;
        RECT 135.600 29.600 136.400 30.400 ;
        RECT 135.700 28.400 136.300 29.600 ;
        RECT 135.600 27.600 136.400 28.400 ;
        RECT 127.600 26.200 128.400 27.000 ;
        RECT 129.000 26.400 133.200 27.000 ;
        RECT 134.200 26.200 135.000 27.000 ;
        RECT 122.800 23.600 123.600 24.400 ;
        RECT 124.400 23.600 125.200 24.400 ;
        RECT 129.200 23.600 130.000 24.400 ;
        RECT 134.000 23.600 134.800 24.400 ;
        RECT 118.000 13.600 118.800 14.400 ;
        RECT 119.600 6.200 120.400 17.800 ;
        RECT 122.900 12.400 123.500 23.600 ;
        RECT 124.500 22.400 125.100 23.600 ;
        RECT 124.400 21.600 125.200 22.400 ;
        RECT 134.100 18.400 134.700 23.600 ;
        RECT 140.500 18.400 141.100 35.600 ;
        RECT 143.600 31.800 144.400 32.600 ;
        RECT 148.500 32.400 149.100 61.600 ;
        RECT 150.000 59.600 150.800 60.400 ;
        RECT 150.100 58.400 150.700 59.600 ;
        RECT 150.000 57.600 150.800 58.400 ;
        RECT 151.600 55.600 152.400 56.400 ;
        RECT 151.700 54.400 152.300 55.600 ;
        RECT 153.300 54.400 153.900 63.600 ;
        RECT 156.500 60.400 157.100 85.600 ;
        RECT 158.000 64.200 158.800 75.800 ;
        RECT 166.100 70.400 166.700 93.600 ;
        RECT 169.300 92.400 169.900 105.600 ;
        RECT 177.200 104.200 178.000 115.800 ;
        RECT 182.000 113.600 182.800 114.400 ;
        RECT 183.700 108.400 184.300 133.600 ;
        RECT 188.500 132.400 189.100 135.600 ;
        RECT 191.700 134.400 192.300 146.400 ;
        RECT 193.200 145.600 194.000 146.400 ;
        RECT 194.800 146.200 195.600 147.000 ;
        RECT 193.200 143.600 194.000 144.400 ;
        RECT 193.300 136.400 193.900 143.600 ;
        RECT 193.200 135.600 194.000 136.400 ;
        RECT 196.500 134.400 197.100 147.600 ;
        RECT 198.100 146.400 198.700 147.600 ;
        RECT 199.800 147.000 200.400 151.800 ;
        RECT 201.000 149.800 201.800 150.600 ;
        RECT 201.200 148.400 201.800 149.800 ;
        RECT 206.200 148.400 206.800 151.800 ;
        RECT 209.200 151.600 210.000 152.400 ;
        RECT 215.600 151.800 216.400 152.600 ;
        RECT 221.800 151.800 222.600 152.600 ;
        RECT 214.000 149.600 214.800 150.400 ;
        RECT 214.100 148.400 214.700 149.600 ;
        RECT 215.600 148.400 216.200 151.800 ;
        RECT 220.600 149.800 221.400 150.600 ;
        RECT 220.600 148.400 221.200 149.800 ;
        RECT 201.200 147.800 206.800 148.400 ;
        RECT 201.200 147.000 202.000 147.200 ;
        RECT 204.600 147.000 205.400 147.200 ;
        RECT 206.200 147.000 206.800 147.800 ;
        RECT 207.600 147.600 208.400 148.400 ;
        RECT 212.400 147.600 213.200 148.400 ;
        RECT 214.000 147.600 214.800 148.400 ;
        RECT 215.600 147.800 221.200 148.400 ;
        RECT 199.800 146.400 205.400 147.000 ;
        RECT 198.000 145.600 198.800 146.400 ;
        RECT 199.800 146.200 200.600 146.400 ;
        RECT 206.000 146.200 206.800 147.000 ;
        RECT 209.200 143.600 210.000 144.400 ;
        RECT 206.000 141.600 206.800 142.400 ;
        RECT 201.200 137.600 202.000 138.400 ;
        RECT 206.100 136.400 206.700 141.600 ;
        RECT 198.000 135.600 198.800 136.400 ;
        RECT 206.000 135.600 206.800 136.400 ;
        RECT 198.100 134.400 198.700 135.600 ;
        RECT 191.600 133.600 192.400 134.400 ;
        RECT 196.400 133.600 197.200 134.400 ;
        RECT 198.000 133.600 198.800 134.400 ;
        RECT 188.400 131.600 189.200 132.400 ;
        RECT 191.600 131.600 192.400 132.400 ;
        RECT 193.200 131.600 194.000 132.400 ;
        RECT 185.200 129.600 186.000 130.400 ;
        RECT 188.400 129.600 189.200 130.400 ;
        RECT 188.500 114.400 189.100 129.600 ;
        RECT 188.400 113.600 189.200 114.400 ;
        RECT 191.700 112.400 192.300 131.600 ;
        RECT 196.500 130.400 197.100 133.600 ;
        RECT 196.400 129.600 197.200 130.400 ;
        RECT 201.200 129.600 202.000 130.400 ;
        RECT 207.600 130.300 208.400 130.400 ;
        RECT 209.300 130.300 209.900 143.600 ;
        RECT 210.800 131.600 211.600 132.400 ;
        RECT 210.900 130.400 211.500 131.600 ;
        RECT 207.600 129.700 209.900 130.300 ;
        RECT 207.600 129.600 208.400 129.700 ;
        RECT 210.800 129.600 211.600 130.400 ;
        RECT 193.200 123.600 194.000 124.400 ;
        RECT 204.400 123.600 205.200 124.400 ;
        RECT 193.300 112.400 193.900 123.600 ;
        RECT 201.200 117.600 202.000 118.400 ;
        RECT 191.600 111.600 192.400 112.400 ;
        RECT 193.200 111.600 194.000 112.400 ;
        RECT 196.400 111.600 197.200 112.400 ;
        RECT 191.700 110.400 192.300 111.600 ;
        RECT 201.300 110.400 201.900 117.600 ;
        RECT 204.500 112.400 205.100 123.600 ;
        RECT 207.700 118.400 208.300 129.600 ;
        RECT 210.800 127.600 211.600 128.400 ;
        RECT 207.600 117.600 208.400 118.400 ;
        RECT 212.500 116.400 213.100 147.600 ;
        RECT 215.600 147.000 216.200 147.800 ;
        RECT 217.000 147.000 217.800 147.200 ;
        RECT 220.400 147.000 221.200 147.200 ;
        RECT 222.000 147.000 222.600 151.800 ;
        RECT 225.200 151.600 226.000 152.400 ;
        RECT 234.800 151.800 235.600 152.600 ;
        RECT 241.400 151.800 242.200 152.600 ;
        RECT 225.300 150.400 225.900 151.600 ;
        RECT 225.200 149.600 226.000 150.400 ;
        RECT 234.800 148.400 235.400 151.800 ;
        RECT 238.800 148.400 239.600 148.600 ;
        RECT 223.600 147.600 224.400 148.400 ;
        RECT 228.400 147.600 229.200 148.400 ;
        RECT 231.600 147.600 232.400 148.400 ;
        RECT 234.800 147.800 239.600 148.400 ;
        RECT 214.000 145.600 214.800 146.400 ;
        RECT 215.600 146.200 216.400 147.000 ;
        RECT 217.000 146.400 222.600 147.000 ;
        RECT 221.800 146.200 222.600 146.400 ;
        RECT 214.100 134.400 214.700 145.600 ;
        RECT 220.400 143.600 221.200 144.400 ;
        RECT 223.700 134.400 224.300 147.600 ;
        RECT 228.500 146.400 229.100 147.600 ;
        RECT 234.800 147.000 235.400 147.800 ;
        RECT 236.200 147.000 237.000 147.200 ;
        RECT 239.600 147.000 240.400 147.200 ;
        RECT 241.600 147.000 242.200 151.800 ;
        RECT 242.800 147.600 243.600 148.400 ;
        RECT 228.400 145.600 229.200 146.400 ;
        RECT 231.600 146.300 232.400 146.400 ;
        RECT 231.600 145.700 233.900 146.300 ;
        RECT 234.800 146.200 235.600 147.000 ;
        RECT 236.200 146.400 240.400 147.000 ;
        RECT 241.400 146.200 242.200 147.000 ;
        RECT 231.600 145.600 232.400 145.700 ;
        RECT 228.500 144.400 229.100 145.600 ;
        RECT 226.800 143.600 227.600 144.400 ;
        RECT 228.400 143.600 229.200 144.400 ;
        RECT 230.000 143.600 230.800 144.400 ;
        RECT 226.900 140.400 227.500 143.600 ;
        RECT 226.800 139.600 227.600 140.400 ;
        RECT 225.200 137.600 226.000 138.400 ;
        RECT 225.300 134.400 225.900 137.600 ;
        RECT 230.100 136.400 230.700 143.600 ;
        RECT 226.800 135.600 227.600 136.400 ;
        RECT 230.000 135.600 230.800 136.400 ;
        RECT 226.900 134.400 227.500 135.600 ;
        RECT 233.300 134.400 233.900 145.700 ;
        RECT 242.900 138.400 243.500 147.600 ;
        RECT 244.500 146.400 245.100 157.600 ;
        RECT 246.000 149.600 246.800 150.400 ;
        RECT 246.100 148.400 246.700 149.600 ;
        RECT 246.000 147.600 246.800 148.400 ;
        RECT 244.400 145.600 245.200 146.400 ;
        RECT 242.800 137.600 243.600 138.400 ;
        RECT 214.000 133.600 214.800 134.400 ;
        RECT 215.600 133.600 216.400 134.400 ;
        RECT 223.600 133.600 224.400 134.400 ;
        RECT 225.200 133.600 226.000 134.400 ;
        RECT 226.800 133.600 227.600 134.400 ;
        RECT 228.400 133.600 229.200 134.400 ;
        RECT 231.600 133.600 232.400 134.400 ;
        RECT 233.200 133.600 234.000 134.400 ;
        RECT 238.000 133.600 238.800 134.400 ;
        RECT 215.700 132.400 216.300 133.600 ;
        RECT 214.000 131.600 214.800 132.400 ;
        RECT 215.600 131.600 216.400 132.400 ;
        RECT 223.600 131.600 224.400 132.400 ;
        RECT 214.100 122.400 214.700 131.600 ;
        RECT 223.700 130.400 224.300 131.600 ;
        RECT 218.800 129.600 219.600 130.400 ;
        RECT 222.000 129.600 222.800 130.400 ;
        RECT 223.600 129.600 224.400 130.400 ;
        RECT 214.000 121.600 214.800 122.400 ;
        RECT 209.200 115.600 210.000 116.400 ;
        RECT 212.400 115.600 213.200 116.400 ;
        RECT 204.400 111.600 205.200 112.400 ;
        RECT 207.600 111.600 208.400 112.400 ;
        RECT 191.600 109.600 192.400 110.400 ;
        RECT 201.200 109.600 202.000 110.400 ;
        RECT 202.800 109.600 203.600 110.400 ;
        RECT 183.600 107.600 184.400 108.400 ;
        RECT 188.400 107.600 189.200 108.400 ;
        RECT 194.800 107.600 195.600 108.400 ;
        RECT 201.200 107.600 202.000 108.400 ;
        RECT 183.700 98.400 184.300 107.600 ;
        RECT 169.200 91.600 170.000 92.400 ;
        RECT 170.800 86.200 171.600 97.800 ;
        RECT 175.600 97.600 176.400 98.400 ;
        RECT 183.600 97.600 184.400 98.400 ;
        RECT 175.700 96.400 176.300 97.600 ;
        RECT 183.700 96.400 184.300 97.600 ;
        RECT 175.600 95.600 176.400 96.400 ;
        RECT 180.400 95.600 181.200 96.400 ;
        RECT 183.600 95.600 184.400 96.400 ;
        RECT 186.800 95.600 187.600 96.400 ;
        RECT 177.200 91.600 178.000 92.400 ;
        RECT 175.600 87.600 176.400 88.400 ;
        RECT 175.700 78.400 176.300 87.600 ;
        RECT 175.600 77.600 176.400 78.400 ;
        RECT 159.600 69.400 160.400 70.400 ;
        RECT 166.000 69.600 166.800 70.400 ;
        RECT 164.400 65.600 165.200 66.400 ;
        RECT 156.400 59.600 157.200 60.400 ;
        RECT 156.400 55.000 157.200 55.800 ;
        RECT 162.600 55.600 163.400 55.800 ;
        RECT 157.800 55.000 163.400 55.600 ;
        RECT 151.600 53.600 152.400 54.400 ;
        RECT 153.200 53.600 154.000 54.400 ;
        RECT 156.400 54.200 157.000 55.000 ;
        RECT 157.800 54.800 158.600 55.000 ;
        RECT 161.200 54.800 162.000 55.000 ;
        RECT 156.400 53.600 162.000 54.200 ;
        RECT 156.400 50.200 157.000 53.600 ;
        RECT 161.400 52.200 162.000 53.600 ;
        RECT 161.400 51.400 162.200 52.200 ;
        RECT 162.800 50.200 163.400 55.000 ;
        RECT 164.500 54.400 165.100 65.600 ;
        RECT 166.100 62.400 166.700 69.600 ;
        RECT 167.600 64.200 168.400 75.800 ;
        RECT 174.000 73.600 174.800 74.400 ;
        RECT 174.100 68.400 174.700 73.600 ;
        RECT 175.600 70.300 176.400 70.400 ;
        RECT 177.300 70.300 177.900 91.600 ;
        RECT 180.500 72.400 181.100 95.600 ;
        RECT 185.200 91.600 186.000 92.400 ;
        RECT 186.800 91.600 187.600 92.400 ;
        RECT 185.300 78.400 185.900 91.600 ;
        RECT 185.200 77.600 186.000 78.400 ;
        RECT 186.900 74.400 187.500 91.600 ;
        RECT 186.800 73.600 187.600 74.400 ;
        RECT 180.400 71.600 181.200 72.400 ;
        RECT 188.500 72.300 189.100 107.600 ;
        RECT 196.400 103.600 197.200 104.400 ;
        RECT 201.200 103.600 202.000 104.400 ;
        RECT 196.500 100.400 197.100 103.600 ;
        RECT 196.400 99.600 197.200 100.400 ;
        RECT 190.000 97.600 190.800 98.400 ;
        RECT 196.400 97.600 197.200 98.400 ;
        RECT 190.100 96.400 190.700 97.600 ;
        RECT 190.000 95.600 190.800 96.400 ;
        RECT 196.500 94.400 197.100 97.600 ;
        RECT 201.300 94.400 201.900 103.600 ;
        RECT 202.900 98.400 203.500 109.600 ;
        RECT 207.700 108.400 208.300 111.600 ;
        RECT 209.300 110.400 209.900 115.600 ;
        RECT 210.800 111.600 211.600 112.400 ;
        RECT 210.900 110.400 211.500 111.600 ;
        RECT 209.200 109.600 210.000 110.400 ;
        RECT 210.800 109.600 211.600 110.400 ;
        RECT 214.100 108.400 214.700 121.600 ;
        RECT 217.200 111.600 218.000 112.400 ;
        RECT 217.300 110.400 217.900 111.600 ;
        RECT 222.100 110.400 222.700 129.600 ;
        RECT 223.600 123.600 224.400 124.400 ;
        RECT 223.700 110.400 224.300 123.600 ;
        RECT 226.900 122.400 227.500 133.600 ;
        RECT 228.500 132.400 229.100 133.600 ;
        RECT 228.400 131.600 229.200 132.400 ;
        RECT 234.800 131.600 235.600 132.400 ;
        RECT 238.100 130.400 238.700 133.600 ;
        RECT 247.700 132.400 248.300 163.600 ;
        RECT 255.600 151.600 256.400 152.400 ;
        RECT 271.600 151.600 272.400 152.400 ;
        RECT 279.600 151.800 280.400 152.600 ;
        RECT 286.200 151.800 287.000 152.600 ;
        RECT 255.700 150.400 256.300 151.600 ;
        RECT 255.600 149.600 256.400 150.400 ;
        RECT 263.600 149.600 264.400 150.400 ;
        RECT 266.800 149.600 267.600 150.400 ;
        RECT 270.000 149.600 270.800 150.400 ;
        RECT 250.800 143.600 251.600 144.400 ;
        RECT 250.900 136.400 251.500 143.600 ;
        RECT 255.700 136.400 256.300 149.600 ;
        RECT 257.200 147.600 258.000 148.400 ;
        RECT 258.800 147.600 259.600 148.400 ;
        RECT 265.200 147.600 266.000 148.400 ;
        RECT 270.100 148.300 270.700 149.600 ;
        RECT 271.700 148.400 272.300 151.600 ;
        RECT 274.800 149.600 275.600 150.400 ;
        RECT 268.500 147.700 270.700 148.300 ;
        RECT 258.900 146.400 259.500 147.600 ;
        RECT 258.800 145.600 259.600 146.400 ;
        RECT 263.600 145.600 264.400 146.400 ;
        RECT 258.900 144.400 259.500 145.600 ;
        RECT 265.300 144.400 265.900 147.600 ;
        RECT 258.800 143.600 259.600 144.400 ;
        RECT 265.200 143.600 266.000 144.400 ;
        RECT 258.900 136.400 259.500 143.600 ;
        RECT 250.800 136.300 251.600 136.400 ;
        RECT 249.300 135.700 251.600 136.300 ;
        RECT 249.300 132.400 249.900 135.700 ;
        RECT 250.800 135.600 251.600 135.700 ;
        RECT 255.600 135.600 256.400 136.400 ;
        RECT 258.800 135.600 259.600 136.400 ;
        RECT 255.700 134.400 256.300 135.600 ;
        RECT 250.800 133.600 251.600 134.400 ;
        RECT 255.600 133.600 256.400 134.400 ;
        RECT 265.200 133.600 266.000 134.400 ;
        RECT 244.400 131.600 245.200 132.400 ;
        RECT 246.000 131.600 246.800 132.400 ;
        RECT 247.600 131.600 248.400 132.400 ;
        RECT 249.200 131.600 250.000 132.400 ;
        RECT 231.600 129.600 232.400 130.400 ;
        RECT 238.000 129.600 238.800 130.400 ;
        RECT 226.800 121.600 227.600 122.400 ;
        RECT 226.800 117.600 227.600 118.400 ;
        RECT 228.400 117.600 229.200 118.400 ;
        RECT 217.200 109.600 218.000 110.400 ;
        RECT 220.400 109.600 221.200 110.400 ;
        RECT 222.000 109.600 222.800 110.400 ;
        RECT 223.600 109.600 224.400 110.400 ;
        RECT 204.400 107.600 205.200 108.400 ;
        RECT 207.600 107.600 208.400 108.400 ;
        RECT 209.200 107.600 210.000 108.400 ;
        RECT 214.000 107.600 214.800 108.400 ;
        RECT 218.800 107.600 219.600 108.400 ;
        RECT 215.600 105.600 216.400 106.400 ;
        RECT 206.000 103.600 206.800 104.400 ;
        RECT 202.800 97.600 203.600 98.400 ;
        RECT 194.800 93.600 195.600 94.400 ;
        RECT 196.400 93.600 197.200 94.400 ;
        RECT 201.200 93.600 202.000 94.400 ;
        RECT 202.800 93.600 203.600 94.400 ;
        RECT 194.800 91.600 195.600 92.400 ;
        RECT 198.000 91.600 198.800 92.400 ;
        RECT 194.900 90.400 195.500 91.600 ;
        RECT 194.800 89.600 195.600 90.400 ;
        RECT 190.000 81.600 190.800 82.400 ;
        RECT 190.100 78.400 190.700 81.600 ;
        RECT 194.900 78.400 195.500 89.600 ;
        RECT 190.000 77.600 190.800 78.400 ;
        RECT 194.800 77.600 195.600 78.400 ;
        RECT 186.900 71.700 189.100 72.300 ;
        RECT 175.600 69.700 177.900 70.300 ;
        RECT 175.600 69.600 176.400 69.700 ;
        RECT 182.000 69.600 182.800 70.400 ;
        RECT 183.600 69.600 184.400 70.400 ;
        RECT 174.000 67.600 174.800 68.400 ;
        RECT 180.400 65.600 181.200 66.400 ;
        RECT 183.700 64.400 184.300 69.600 ;
        RECT 186.900 68.400 187.500 71.700 ;
        RECT 191.600 71.600 192.400 72.400 ;
        RECT 188.400 69.600 189.200 70.400 ;
        RECT 188.500 68.400 189.100 69.600 ;
        RECT 186.800 67.600 187.600 68.400 ;
        RECT 188.400 67.600 189.200 68.400 ;
        RECT 186.900 66.400 187.500 67.600 ;
        RECT 186.800 65.600 187.600 66.400 ;
        RECT 191.700 64.400 192.300 71.600 ;
        RECT 193.200 69.600 194.000 70.400 ;
        RECT 198.100 70.300 198.700 91.600 ;
        RECT 201.300 90.400 201.900 93.600 ;
        RECT 202.900 92.400 203.500 93.600 ;
        RECT 206.100 92.400 206.700 103.600 ;
        RECT 212.400 99.600 213.200 100.400 ;
        RECT 207.600 93.600 208.400 94.400 ;
        RECT 212.500 92.400 213.100 99.600 ;
        RECT 202.800 91.600 203.600 92.400 ;
        RECT 206.000 91.600 206.800 92.400 ;
        RECT 212.400 91.600 213.200 92.400 ;
        RECT 215.700 90.400 216.300 105.600 ;
        RECT 218.900 104.400 219.500 107.600 ;
        RECT 218.800 103.600 219.600 104.400 ;
        RECT 220.500 102.400 221.100 109.600 ;
        RECT 220.400 101.600 221.200 102.400 ;
        RECT 220.500 100.400 221.100 101.600 ;
        RECT 220.400 99.600 221.200 100.400 ;
        RECT 218.800 97.600 219.600 98.400 ;
        RECT 217.200 93.600 218.000 94.400 ;
        RECT 201.200 89.600 202.000 90.400 ;
        RECT 202.800 89.600 203.600 90.400 ;
        RECT 215.600 89.600 216.400 90.400 ;
        RECT 202.900 88.400 203.500 89.600 ;
        RECT 202.800 87.600 203.600 88.400 ;
        RECT 199.600 83.600 200.400 84.400 ;
        RECT 206.000 83.600 206.800 84.400 ;
        RECT 214.000 83.600 214.800 84.400 ;
        RECT 199.700 78.400 200.300 83.600 ;
        RECT 199.600 77.600 200.400 78.400 ;
        RECT 202.800 71.600 203.600 72.400 ;
        RECT 199.600 70.300 200.400 70.400 ;
        RECT 198.100 69.700 200.400 70.300 ;
        RECT 199.600 69.600 200.400 69.700 ;
        RECT 196.400 67.600 197.200 68.400 ;
        RECT 198.000 67.600 198.800 68.400 ;
        RECT 196.500 66.400 197.100 67.600 ;
        RECT 198.100 66.400 198.700 67.600 ;
        RECT 196.400 65.600 197.200 66.400 ;
        RECT 198.000 65.600 198.800 66.400 ;
        RECT 172.400 63.600 173.200 64.400 ;
        RECT 183.600 63.600 184.400 64.400 ;
        RECT 191.600 63.600 192.400 64.400 ;
        RECT 196.400 63.600 197.200 64.400 ;
        RECT 166.000 61.600 166.800 62.400 ;
        RECT 178.800 61.600 179.600 62.400 ;
        RECT 166.000 59.600 166.800 60.400 ;
        RECT 166.100 54.400 166.700 59.600 ;
        RECT 167.600 55.000 168.400 55.800 ;
        RECT 169.000 55.000 173.200 55.600 ;
        RECT 174.200 55.000 175.000 55.800 ;
        RECT 164.400 53.600 165.200 54.400 ;
        RECT 166.000 53.600 166.800 54.400 ;
        RECT 167.600 54.200 168.200 55.000 ;
        RECT 169.000 54.800 169.800 55.000 ;
        RECT 172.400 54.800 173.200 55.000 ;
        RECT 167.600 53.600 172.400 54.200 ;
        RECT 156.400 49.400 157.200 50.200 ;
        RECT 162.600 49.400 163.400 50.200 ;
        RECT 167.600 50.200 168.200 53.600 ;
        RECT 171.600 53.400 172.400 53.600 ;
        RECT 172.400 51.600 173.200 52.400 ;
        RECT 167.600 49.400 168.400 50.200 ;
        RECT 172.500 48.400 173.100 51.600 ;
        RECT 174.400 50.200 175.000 55.000 ;
        RECT 175.600 53.600 176.400 54.400 ;
        RECT 177.200 50.200 178.000 55.800 ;
        RECT 178.900 54.400 179.500 61.600 ;
        RECT 178.800 53.600 179.600 54.400 ;
        RECT 174.200 49.400 175.000 50.200 ;
        RECT 172.400 47.600 173.200 48.400 ;
        RECT 156.400 45.600 157.200 46.400 ;
        RECT 174.000 45.600 174.800 46.400 ;
        RECT 180.400 46.200 181.200 57.800 ;
        RECT 182.000 51.600 182.800 52.600 ;
        RECT 153.200 41.600 154.000 42.400 ;
        RECT 151.600 35.600 152.400 36.400 ;
        RECT 143.600 28.400 144.200 31.800 ;
        RECT 148.400 31.600 149.200 32.400 ;
        RECT 149.800 31.800 150.600 32.600 ;
        RECT 148.600 29.800 149.400 30.600 ;
        RECT 148.600 28.400 149.200 29.800 ;
        RECT 142.000 27.600 142.800 28.400 ;
        RECT 143.600 27.800 149.200 28.400 ;
        RECT 142.100 22.400 142.700 27.600 ;
        RECT 143.600 27.000 144.200 27.800 ;
        RECT 145.000 27.000 145.800 27.200 ;
        RECT 148.400 27.000 149.200 27.200 ;
        RECT 150.000 27.000 150.600 31.800 ;
        RECT 151.700 28.400 152.300 35.600 ;
        RECT 153.300 28.400 153.900 41.600 ;
        RECT 156.500 32.400 157.100 45.600 ;
        RECT 158.000 43.600 158.800 44.400 ;
        RECT 158.100 38.400 158.700 43.600 ;
        RECT 158.000 37.600 158.800 38.400 ;
        RECT 164.400 37.600 165.200 38.400 ;
        RECT 158.000 33.600 158.800 34.400 ;
        RECT 156.400 31.600 157.200 32.400 ;
        RECT 158.100 30.300 158.700 33.600 ;
        RECT 164.500 32.400 165.100 37.600 ;
        RECT 164.400 31.600 165.200 32.400 ;
        RECT 170.800 31.600 171.600 32.400 ;
        RECT 156.500 29.700 158.700 30.300 ;
        RECT 151.600 27.600 152.400 28.400 ;
        RECT 153.200 27.600 154.000 28.400 ;
        RECT 143.600 26.200 144.400 27.000 ;
        RECT 145.000 26.400 150.600 27.000 ;
        RECT 153.300 26.400 153.900 27.600 ;
        RECT 149.800 26.200 150.600 26.400 ;
        RECT 153.200 25.600 154.000 26.400 ;
        RECT 148.400 23.600 149.200 24.400 ;
        RECT 154.800 23.600 155.600 24.400 ;
        RECT 142.000 21.600 142.800 22.400 ;
        RECT 148.500 18.400 149.100 23.600 ;
        RECT 122.800 11.600 123.600 12.400 ;
        RECT 129.200 6.200 130.000 17.800 ;
        RECT 134.000 17.600 134.800 18.400 ;
        RECT 140.400 17.600 141.200 18.400 ;
        RECT 148.400 17.600 149.200 18.400 ;
        RECT 140.500 14.400 141.100 17.600 ;
        RECT 154.900 16.400 155.500 23.600 ;
        RECT 156.500 18.400 157.100 29.700 ;
        RECT 161.200 27.600 162.000 28.400 ;
        RECT 162.800 27.600 163.600 28.400 ;
        RECT 164.500 28.300 165.100 31.600 ;
        RECT 167.600 29.600 168.400 30.400 ;
        RECT 172.400 29.600 173.200 30.400 ;
        RECT 166.000 28.300 166.800 28.400 ;
        RECT 164.500 27.700 166.800 28.300 ;
        RECT 166.000 27.600 166.800 27.700 ;
        RECT 159.600 23.600 160.400 24.400 ;
        RECT 159.700 22.400 160.300 23.600 ;
        RECT 159.600 21.600 160.400 22.400 ;
        RECT 156.400 17.600 157.200 18.400 ;
        RECT 161.300 16.400 161.900 27.600 ;
        RECT 141.800 15.000 142.600 15.800 ;
        RECT 143.600 15.000 147.800 15.600 ;
        RECT 148.400 15.000 149.200 15.800 ;
        RECT 151.600 15.600 152.400 16.400 ;
        RECT 154.800 15.600 155.600 16.400 ;
        RECT 159.600 15.600 160.400 16.400 ;
        RECT 161.200 15.600 162.000 16.400 ;
        RECT 164.400 15.600 165.200 16.400 ;
        RECT 166.100 16.300 166.700 27.600 ;
        RECT 172.500 22.400 173.100 29.600 ;
        RECT 174.100 28.400 174.700 45.600 ;
        RECT 177.200 43.600 178.000 44.400 ;
        RECT 175.600 39.600 176.400 40.400 ;
        RECT 175.700 30.400 176.300 39.600 ;
        RECT 175.600 29.600 176.400 30.400 ;
        RECT 174.000 27.600 174.800 28.400 ;
        RECT 172.400 21.600 173.200 22.400 ;
        RECT 167.600 16.300 168.400 16.400 ;
        RECT 166.100 15.700 168.400 16.300 ;
        RECT 167.600 15.600 168.400 15.700 ;
        RECT 170.800 15.600 171.600 16.400 ;
        RECT 140.400 13.600 141.200 14.400 ;
        RECT 141.800 10.200 142.400 15.000 ;
        RECT 143.600 14.800 144.400 15.000 ;
        RECT 147.000 14.800 147.800 15.000 ;
        RECT 148.600 14.200 149.200 15.000 ;
        RECT 151.700 14.400 152.300 15.600 ;
        RECT 161.300 14.400 161.900 15.600 ;
        RECT 172.500 14.400 173.100 21.600 ;
        RECT 177.300 20.400 177.900 43.600 ;
        RECT 183.700 40.400 184.300 63.600 ;
        RECT 196.500 58.400 197.100 63.600 ;
        RECT 190.000 46.200 190.800 57.800 ;
        RECT 196.400 57.600 197.200 58.400 ;
        RECT 199.700 56.300 200.300 69.600 ;
        RECT 202.900 68.400 203.500 71.600 ;
        RECT 206.100 70.400 206.700 83.600 ;
        RECT 210.800 71.600 211.600 72.400 ;
        RECT 206.000 69.600 206.800 70.400 ;
        RECT 212.400 70.300 213.200 70.400 ;
        RECT 214.100 70.300 214.700 83.600 ;
        RECT 217.300 82.400 217.900 93.600 ;
        RECT 218.900 92.400 219.500 97.600 ;
        RECT 220.400 93.600 221.200 94.400 ;
        RECT 218.800 91.600 219.600 92.400 ;
        RECT 218.800 85.600 219.600 86.400 ;
        RECT 217.200 81.600 218.000 82.400 ;
        RECT 218.900 70.400 219.500 85.600 ;
        RECT 220.500 74.400 221.100 93.600 ;
        RECT 222.100 90.300 222.700 109.600 ;
        RECT 226.900 108.400 227.500 117.600 ;
        RECT 228.500 110.400 229.100 117.600 ;
        RECT 230.000 111.600 230.800 112.400 ;
        RECT 233.200 112.300 234.000 112.400 ;
        RECT 233.200 111.700 235.500 112.300 ;
        RECT 233.200 111.600 234.000 111.700 ;
        RECT 228.400 109.600 229.200 110.400 ;
        RECT 223.600 107.600 224.400 108.400 ;
        RECT 225.200 107.600 226.000 108.400 ;
        RECT 226.800 107.600 227.600 108.400 ;
        RECT 230.100 106.400 230.700 111.600 ;
        RECT 234.900 110.400 235.500 111.700 ;
        RECT 242.800 111.600 243.600 112.400 ;
        RECT 242.900 110.400 243.500 111.600 ;
        RECT 244.500 110.400 245.100 131.600 ;
        RECT 246.100 128.400 246.700 131.600 ;
        RECT 246.000 127.600 246.800 128.400 ;
        RECT 250.900 122.400 251.500 133.600 ;
        RECT 265.300 132.400 265.900 133.600 ;
        RECT 268.500 132.400 269.100 147.700 ;
        RECT 271.600 147.600 272.400 148.400 ;
        RECT 273.200 147.600 274.000 148.400 ;
        RECT 270.000 145.600 270.800 146.400 ;
        RECT 270.100 134.400 270.700 145.600 ;
        RECT 270.000 133.600 270.800 134.400 ;
        RECT 252.400 131.600 253.200 132.400 ;
        RECT 265.200 131.600 266.000 132.400 ;
        RECT 268.400 131.600 269.200 132.400 ;
        RECT 252.500 130.400 253.100 131.600 ;
        RECT 252.400 129.600 253.200 130.400 ;
        RECT 268.400 129.600 269.200 130.400 ;
        RECT 271.600 129.600 272.400 130.400 ;
        RECT 252.400 127.600 253.200 128.400 ;
        RECT 250.800 121.600 251.600 122.400 ;
        RECT 252.500 118.400 253.100 127.600 ;
        RECT 265.200 123.600 266.000 124.400 ;
        RECT 265.300 118.400 265.900 123.600 ;
        RECT 270.000 121.600 270.800 122.400 ;
        RECT 252.400 117.600 253.200 118.400 ;
        RECT 265.200 117.600 266.000 118.400 ;
        RECT 247.600 111.800 248.400 112.600 ;
        RECT 253.800 111.800 254.600 112.600 ;
        RECT 265.300 112.400 265.900 117.600 ;
        RECT 233.200 109.600 234.000 110.400 ;
        RECT 234.800 109.600 235.600 110.400 ;
        RECT 241.200 109.600 242.000 110.400 ;
        RECT 242.800 109.600 243.600 110.400 ;
        RECT 244.400 109.600 245.200 110.400 ;
        RECT 233.300 108.400 233.900 109.600 ;
        RECT 233.200 107.600 234.000 108.400 ;
        RECT 234.800 107.600 235.600 108.400 ;
        RECT 239.600 107.600 240.400 108.400 ;
        RECT 223.600 105.600 224.400 106.400 ;
        RECT 230.000 105.600 230.800 106.400 ;
        RECT 223.700 98.400 224.300 105.600 ;
        RECT 233.300 98.400 233.900 107.600 ;
        RECT 234.900 104.400 235.500 107.600 ;
        RECT 239.700 106.400 240.300 107.600 ;
        RECT 239.600 105.600 240.400 106.400 ;
        RECT 234.800 103.600 235.600 104.400 ;
        RECT 223.600 97.600 224.400 98.400 ;
        RECT 230.000 97.600 230.800 98.400 ;
        RECT 233.200 97.600 234.000 98.400 ;
        RECT 230.100 94.400 230.700 97.600 ;
        RECT 233.200 95.600 234.000 96.400 ;
        RECT 230.000 93.600 230.800 94.400 ;
        RECT 233.300 92.400 233.900 95.600 ;
        RECT 241.300 94.400 241.900 109.600 ;
        RECT 242.800 103.600 243.600 104.400 ;
        RECT 242.900 96.400 243.500 103.600 ;
        RECT 242.800 95.600 243.600 96.400 ;
        RECT 236.400 93.600 237.200 94.400 ;
        RECT 241.200 93.600 242.000 94.400 ;
        RECT 244.500 92.400 245.100 109.600 ;
        RECT 247.600 108.400 248.200 111.800 ;
        RECT 252.600 109.800 253.400 110.600 ;
        RECT 252.600 108.400 253.200 109.800 ;
        RECT 246.000 107.600 246.800 108.400 ;
        RECT 247.600 107.800 253.200 108.400 ;
        RECT 246.100 96.400 246.700 107.600 ;
        RECT 247.600 107.000 248.200 107.800 ;
        RECT 249.000 107.000 249.800 107.200 ;
        RECT 252.400 107.000 253.200 107.200 ;
        RECT 254.000 107.000 254.600 111.800 ;
        RECT 260.400 111.600 261.200 112.400 ;
        RECT 265.200 111.600 266.000 112.400 ;
        RECT 255.600 107.600 256.400 108.400 ;
        RECT 247.600 106.200 248.400 107.000 ;
        RECT 249.000 106.400 254.600 107.000 ;
        RECT 253.800 106.200 254.600 106.400 ;
        RECT 257.200 105.600 258.000 106.400 ;
        RECT 257.300 104.400 257.900 105.600 ;
        RECT 257.200 103.600 258.000 104.400 ;
        RECT 258.800 103.600 259.600 104.400 ;
        RECT 260.500 102.400 261.100 111.600 ;
        RECT 268.400 109.600 269.200 110.400 ;
        RECT 263.600 107.600 264.400 108.400 ;
        RECT 265.200 103.600 266.000 104.400 ;
        RECT 265.300 102.400 265.900 103.600 ;
        RECT 260.400 101.600 261.200 102.400 ;
        RECT 265.200 101.600 266.000 102.400 ;
        RECT 270.100 98.400 270.700 121.600 ;
        RECT 273.300 116.400 273.900 147.600 ;
        RECT 274.900 146.400 275.500 149.600 ;
        RECT 279.600 148.400 280.200 151.800 ;
        RECT 281.200 149.600 282.000 150.400 ;
        RECT 283.600 148.400 284.400 148.600 ;
        RECT 276.400 147.600 277.200 148.400 ;
        RECT 278.000 147.600 278.800 148.400 ;
        RECT 279.600 147.800 284.400 148.400 ;
        RECT 274.800 145.600 275.600 146.400 ;
        RECT 276.500 138.400 277.100 147.600 ;
        RECT 278.100 142.400 278.700 147.600 ;
        RECT 279.600 147.000 280.200 147.800 ;
        RECT 281.000 147.000 281.800 147.200 ;
        RECT 284.400 147.000 285.200 147.200 ;
        RECT 286.400 147.000 287.000 151.800 ;
        RECT 287.600 147.600 288.400 148.400 ;
        RECT 279.600 146.200 280.400 147.000 ;
        RECT 281.000 146.400 285.200 147.000 ;
        RECT 286.200 146.200 287.000 147.000 ;
        RECT 287.700 144.400 288.300 147.600 ;
        RECT 294.000 146.200 294.800 151.800 ;
        RECT 279.600 143.600 280.400 144.400 ;
        RECT 287.600 143.600 288.400 144.400 ;
        RECT 297.200 144.200 298.000 155.800 ;
        RECT 298.800 153.600 299.600 154.400 ;
        RECT 298.900 150.200 299.500 153.600 ;
        RECT 305.300 150.400 305.900 167.600 ;
        RECT 298.800 149.400 299.600 150.200 ;
        RECT 305.200 149.600 306.000 150.400 ;
        RECT 306.800 144.200 307.600 155.800 ;
        RECT 308.400 153.600 309.200 154.400 ;
        RECT 278.000 141.600 278.800 142.400 ;
        RECT 276.400 137.600 277.200 138.400 ;
        RECT 274.800 129.600 275.600 130.400 ;
        RECT 276.400 129.600 277.200 130.400 ;
        RECT 274.900 122.400 275.500 129.600 ;
        RECT 274.800 121.600 275.600 122.400 ;
        RECT 276.500 120.400 277.100 129.600 ;
        RECT 276.400 119.600 277.200 120.400 ;
        RECT 273.200 115.600 274.000 116.400 ;
        RECT 273.300 112.300 273.900 115.600 ;
        RECT 274.800 112.300 275.600 112.400 ;
        RECT 273.300 111.700 275.600 112.300 ;
        RECT 274.800 111.600 275.600 111.700 ;
        RECT 278.000 111.600 278.800 112.400 ;
        RECT 278.100 110.400 278.700 111.600 ;
        RECT 279.700 110.400 280.300 143.600 ;
        RECT 281.200 137.600 282.000 138.400 ;
        RECT 281.300 136.400 281.900 137.600 ;
        RECT 281.200 135.600 282.000 136.400 ;
        RECT 295.600 135.600 296.400 136.400 ;
        RECT 295.700 134.400 296.300 135.600 ;
        RECT 297.200 135.000 298.000 135.800 ;
        RECT 303.400 135.600 304.200 135.800 ;
        RECT 298.600 135.000 304.200 135.600 ;
        RECT 281.200 134.300 282.000 134.400 ;
        RECT 281.200 133.700 283.500 134.300 ;
        RECT 281.200 133.600 282.000 133.700 ;
        RECT 281.200 111.600 282.000 112.400 ;
        RECT 274.800 109.600 275.600 110.400 ;
        RECT 278.000 109.600 278.800 110.400 ;
        RECT 279.600 109.600 280.400 110.400 ;
        RECT 271.600 107.600 272.400 108.400 ;
        RECT 268.400 97.600 269.200 98.400 ;
        RECT 270.000 97.600 270.800 98.400 ;
        RECT 246.000 95.600 246.800 96.400 ;
        RECT 246.100 92.400 246.700 95.600 ;
        RECT 258.800 95.000 259.600 95.800 ;
        RECT 260.200 95.000 264.400 95.600 ;
        RECT 265.400 95.000 266.200 95.800 ;
        RECT 255.600 93.600 256.400 94.400 ;
        RECT 257.200 93.600 258.000 94.400 ;
        RECT 258.800 94.200 259.400 95.000 ;
        RECT 260.200 94.800 261.000 95.000 ;
        RECT 263.600 94.800 264.400 95.000 ;
        RECT 258.800 93.600 263.600 94.200 ;
        RECT 226.800 91.600 227.600 92.400 ;
        RECT 233.200 91.600 234.000 92.400 ;
        RECT 234.800 91.600 235.600 92.400 ;
        RECT 241.200 91.600 242.000 92.400 ;
        RECT 244.400 92.300 245.200 92.400 ;
        RECT 242.900 91.700 245.200 92.300 ;
        RECT 223.600 90.300 224.400 90.400 ;
        RECT 222.100 89.700 224.400 90.300 ;
        RECT 223.600 89.600 224.400 89.700 ;
        RECT 225.200 89.600 226.000 90.400 ;
        RECT 222.000 87.600 222.800 88.400 ;
        RECT 222.100 78.400 222.700 87.600 ;
        RECT 225.300 84.400 225.900 89.600 ;
        RECT 225.200 83.600 226.000 84.400 ;
        RECT 222.000 77.600 222.800 78.400 ;
        RECT 220.400 73.600 221.200 74.400 ;
        RECT 226.900 70.400 227.500 91.600 ;
        RECT 234.900 90.400 235.500 91.600 ;
        RECT 234.800 89.600 235.600 90.400 ;
        RECT 239.600 89.600 240.400 90.400 ;
        RECT 228.400 73.600 229.200 74.400 ;
        RECT 212.400 69.700 214.700 70.300 ;
        RECT 212.400 69.600 213.200 69.700 ;
        RECT 218.800 69.600 219.600 70.400 ;
        RECT 226.800 69.600 227.600 70.400 ;
        RECT 202.800 67.600 203.600 68.400 ;
        RECT 212.400 67.600 213.200 68.400 ;
        RECT 223.600 67.600 224.400 68.400 ;
        RECT 226.800 67.600 227.600 68.400 ;
        RECT 228.400 67.600 229.200 68.400 ;
        RECT 202.900 58.400 203.500 67.600 ;
        RECT 206.000 65.600 206.800 66.400 ;
        RECT 212.500 64.400 213.100 67.600 ;
        RECT 223.700 66.400 224.300 67.600 ;
        RECT 214.000 65.600 214.800 66.400 ;
        RECT 215.600 65.600 216.400 66.400 ;
        RECT 220.400 65.600 221.200 66.400 ;
        RECT 223.600 66.300 224.400 66.400 ;
        RECT 222.100 65.700 224.400 66.300 ;
        RECT 212.400 63.600 213.200 64.400 ;
        RECT 206.000 61.600 206.800 62.400 ;
        RECT 214.100 62.300 214.700 65.600 ;
        RECT 220.500 64.400 221.100 65.600 ;
        RECT 220.400 63.600 221.200 64.400 ;
        RECT 212.500 61.700 214.700 62.300 ;
        RECT 206.100 58.400 206.700 61.600 ;
        RECT 202.800 57.600 203.600 58.400 ;
        RECT 206.000 57.600 206.800 58.400 ;
        RECT 198.100 55.700 200.300 56.300 ;
        RECT 198.100 54.400 198.700 55.700 ;
        RECT 201.200 55.000 202.000 55.800 ;
        RECT 207.400 55.600 208.200 55.800 ;
        RECT 202.600 55.000 208.200 55.600 ;
        RECT 198.000 53.600 198.800 54.400 ;
        RECT 199.600 53.600 200.400 54.400 ;
        RECT 201.200 54.200 201.800 55.000 ;
        RECT 202.600 54.800 203.400 55.000 ;
        RECT 206.000 54.800 206.800 55.000 ;
        RECT 201.200 53.600 206.800 54.200 ;
        RECT 193.200 47.600 194.000 48.400 ;
        RECT 183.600 39.600 184.400 40.400 ;
        RECT 193.300 38.400 193.900 47.600 ;
        RECT 194.800 44.300 195.600 44.400 ;
        RECT 194.800 43.700 197.100 44.300 ;
        RECT 194.800 43.600 195.600 43.700 ;
        RECT 193.200 37.600 194.000 38.400 ;
        RECT 178.800 31.600 179.600 32.400 ;
        RECT 188.400 31.800 189.200 32.600 ;
        RECT 195.000 31.800 195.800 32.600 ;
        RECT 178.900 22.400 179.500 31.600 ;
        RECT 183.600 29.600 184.400 30.400 ;
        RECT 188.400 28.400 189.000 31.800 ;
        RECT 192.400 28.400 193.200 28.600 ;
        RECT 182.000 27.600 182.800 28.400 ;
        RECT 185.200 27.600 186.000 28.400 ;
        RECT 186.800 27.600 187.600 28.400 ;
        RECT 188.400 27.800 193.200 28.400 ;
        RECT 182.100 26.400 182.700 27.600 ;
        RECT 182.000 25.600 182.800 26.400 ;
        RECT 185.300 22.400 185.900 27.600 ;
        RECT 178.800 21.600 179.600 22.400 ;
        RECT 185.200 21.600 186.000 22.400 ;
        RECT 177.200 19.600 178.000 20.400 ;
        RECT 174.000 17.600 174.800 18.400 ;
        RECT 144.400 13.600 149.200 14.200 ;
        RECT 150.000 13.600 150.800 14.400 ;
        RECT 151.600 13.600 152.400 14.400 ;
        RECT 161.200 13.600 162.000 14.400 ;
        RECT 172.400 13.600 173.200 14.400 ;
        RECT 144.400 13.400 145.200 13.600 ;
        RECT 148.600 10.200 149.200 13.600 ;
        RECT 174.100 12.400 174.700 17.600 ;
        RECT 174.000 11.600 174.800 12.400 ;
        RECT 175.600 12.300 176.400 12.400 ;
        RECT 177.300 12.300 177.900 19.600 ;
        RECT 178.900 12.400 179.500 21.600 ;
        RECT 186.900 18.400 187.500 27.600 ;
        RECT 188.400 27.000 189.000 27.800 ;
        RECT 189.800 27.000 190.600 27.200 ;
        RECT 193.200 27.000 194.000 27.200 ;
        RECT 195.200 27.000 195.800 31.800 ;
        RECT 196.500 30.400 197.100 43.700 ;
        RECT 198.100 42.400 198.700 53.600 ;
        RECT 199.700 46.400 200.300 53.600 ;
        RECT 201.200 50.200 201.800 53.600 ;
        RECT 206.200 52.200 206.800 53.600 ;
        RECT 206.200 51.400 207.000 52.200 ;
        RECT 207.600 50.200 208.200 55.000 ;
        RECT 212.500 54.400 213.100 61.700 ;
        RECT 222.100 58.400 222.700 65.700 ;
        RECT 223.600 65.600 224.400 65.700 ;
        RECT 225.200 66.300 226.000 66.400 ;
        RECT 228.500 66.300 229.100 67.600 ;
        RECT 225.200 65.700 229.100 66.300 ;
        RECT 225.200 65.600 226.000 65.700 ;
        RECT 226.800 63.600 227.600 64.400 ;
        RECT 226.900 58.400 227.500 63.600 ;
        RECT 215.600 57.600 216.400 58.400 ;
        RECT 222.000 57.600 222.800 58.400 ;
        RECT 226.800 57.600 227.600 58.400 ;
        RECT 233.200 58.300 234.000 58.400 ;
        RECT 234.900 58.300 235.500 89.600 ;
        RECT 239.700 84.400 240.300 89.600 ;
        RECT 239.600 83.600 240.400 84.400 ;
        RECT 239.700 70.300 240.300 83.600 ;
        RECT 241.200 70.300 242.000 70.400 ;
        RECT 239.700 69.700 242.000 70.300 ;
        RECT 241.200 69.600 242.000 69.700 ;
        RECT 239.600 67.600 240.400 68.400 ;
        RECT 236.400 65.600 237.200 66.400 ;
        RECT 233.200 57.700 235.500 58.300 ;
        RECT 233.200 57.600 234.000 57.700 ;
        RECT 215.700 54.400 216.300 57.600 ;
        RECT 223.600 55.600 224.400 56.400 ;
        RECT 230.000 55.600 230.800 56.400 ;
        RECT 209.200 53.600 210.000 54.400 ;
        RECT 212.400 53.600 213.200 54.400 ;
        RECT 215.600 53.600 216.400 54.400 ;
        RECT 217.200 53.600 218.000 54.400 ;
        RECT 220.400 53.600 221.200 54.400 ;
        RECT 217.300 52.400 217.900 53.600 ;
        RECT 217.200 51.600 218.000 52.400 ;
        RECT 201.200 49.400 202.000 50.200 ;
        RECT 207.400 49.400 208.200 50.200 ;
        RECT 210.800 49.600 211.600 50.400 ;
        RECT 210.900 46.400 211.500 49.600 ;
        RECT 199.600 45.600 200.400 46.400 ;
        RECT 207.600 45.600 208.400 46.400 ;
        RECT 210.800 45.600 211.600 46.400 ;
        RECT 198.000 41.600 198.800 42.400 ;
        RECT 199.600 31.600 200.400 32.400 ;
        RECT 204.400 31.600 205.200 32.400 ;
        RECT 196.400 29.600 197.200 30.400 ;
        RECT 198.000 29.600 198.800 30.400 ;
        RECT 198.100 28.400 198.700 29.600 ;
        RECT 199.700 28.400 200.300 31.600 ;
        RECT 204.500 28.400 205.100 31.600 ;
        RECT 206.000 29.600 206.800 30.400 ;
        RECT 206.100 28.400 206.700 29.600 ;
        RECT 196.400 27.600 197.200 28.400 ;
        RECT 198.000 27.600 198.800 28.400 ;
        RECT 199.600 27.600 200.400 28.400 ;
        RECT 204.400 27.600 205.200 28.400 ;
        RECT 206.000 27.600 206.800 28.400 ;
        RECT 188.400 26.200 189.200 27.000 ;
        RECT 189.800 26.400 194.000 27.000 ;
        RECT 195.000 26.200 195.800 27.000 ;
        RECT 196.500 26.400 197.100 27.600 ;
        RECT 196.400 25.600 197.200 26.400 ;
        RECT 202.800 25.600 203.600 26.400 ;
        RECT 201.200 23.600 202.000 24.400 ;
        RECT 193.200 21.600 194.000 22.400 ;
        RECT 188.400 19.600 189.200 20.400 ;
        RECT 188.500 18.400 189.100 19.600 ;
        RECT 186.800 17.600 187.600 18.400 ;
        RECT 188.400 17.600 189.200 18.400 ;
        RECT 191.600 17.600 192.400 18.400 ;
        RECT 183.800 15.600 184.600 15.800 ;
        RECT 183.800 15.000 189.400 15.600 ;
        RECT 190.000 15.000 190.800 15.800 ;
        RECT 182.000 13.600 182.800 14.400 ;
        RECT 175.600 11.700 177.900 12.300 ;
        RECT 175.600 11.600 176.400 11.700 ;
        RECT 178.800 11.600 179.600 12.400 ;
        RECT 141.800 9.400 142.600 10.200 ;
        RECT 148.400 9.400 149.200 10.200 ;
        RECT 183.800 10.200 184.400 15.000 ;
        RECT 185.200 14.800 186.000 15.000 ;
        RECT 188.600 14.800 189.400 15.000 ;
        RECT 190.200 14.200 190.800 15.000 ;
        RECT 191.700 14.400 192.300 17.600 ;
        RECT 193.300 14.400 193.900 21.600 ;
        RECT 199.600 17.600 200.400 18.400 ;
        RECT 194.800 15.600 195.600 16.400 ;
        RECT 199.700 16.300 200.300 17.600 ;
        RECT 198.100 15.700 200.300 16.300 ;
        RECT 185.200 13.600 190.800 14.200 ;
        RECT 191.600 13.600 192.400 14.400 ;
        RECT 193.200 13.600 194.000 14.400 ;
        RECT 185.200 12.200 185.800 13.600 ;
        RECT 185.000 11.400 185.800 12.200 ;
        RECT 190.200 10.200 190.800 13.600 ;
        RECT 194.900 12.400 195.500 15.600 ;
        RECT 194.800 11.600 195.600 12.400 ;
        RECT 198.100 10.400 198.700 15.700 ;
        RECT 199.600 13.600 200.400 14.400 ;
        RECT 199.700 12.400 200.300 13.600 ;
        RECT 199.600 11.600 200.400 12.400 ;
        RECT 183.800 9.400 184.600 10.200 ;
        RECT 190.000 9.400 190.800 10.200 ;
        RECT 198.000 9.600 198.800 10.400 ;
        RECT 201.300 8.400 201.900 23.600 ;
        RECT 202.900 20.400 203.500 25.600 ;
        RECT 202.800 19.600 203.600 20.400 ;
        RECT 206.000 11.600 206.800 12.400 ;
        RECT 206.100 10.400 206.700 11.600 ;
        RECT 206.000 10.300 206.800 10.400 ;
        RECT 207.700 10.300 208.300 45.600 ;
        RECT 217.300 36.400 217.900 51.600 ;
        RECT 218.800 43.600 219.600 44.400 ;
        RECT 218.900 38.400 219.500 43.600 ;
        RECT 218.800 37.600 219.600 38.400 ;
        RECT 217.200 35.600 218.000 36.400 ;
        RECT 218.800 35.600 219.600 36.400 ;
        RECT 218.900 34.300 219.500 35.600 ;
        RECT 217.300 33.700 219.500 34.300 ;
        RECT 210.800 31.600 211.600 32.400 ;
        RECT 215.600 31.600 216.400 32.400 ;
        RECT 210.900 30.400 211.500 31.600 ;
        RECT 210.800 29.600 211.600 30.400 ;
        RECT 214.000 27.600 214.800 28.400 ;
        RECT 209.200 25.600 210.000 26.400 ;
        RECT 209.300 24.400 209.900 25.600 ;
        RECT 209.200 23.600 210.000 24.400 ;
        RECT 210.800 23.600 211.600 24.400 ;
        RECT 210.900 18.400 211.500 23.600 ;
        RECT 215.700 18.400 216.300 31.600 ;
        RECT 217.300 26.400 217.900 33.700 ;
        RECT 218.800 31.600 219.600 32.400 ;
        RECT 218.800 29.600 219.600 30.400 ;
        RECT 218.900 26.400 219.500 29.600 ;
        RECT 220.500 28.400 221.100 53.600 ;
        RECT 230.100 52.400 230.700 55.600 ;
        RECT 233.300 52.400 233.900 57.600 ;
        RECT 234.800 53.600 235.600 54.400 ;
        RECT 234.900 52.400 235.500 53.600 ;
        RECT 230.000 51.600 230.800 52.400 ;
        RECT 233.200 51.600 234.000 52.400 ;
        RECT 234.800 51.600 235.600 52.400 ;
        RECT 236.500 50.400 237.100 65.600 ;
        RECT 238.000 63.600 238.800 64.400 ;
        RECT 242.900 58.400 243.500 91.700 ;
        RECT 244.400 91.600 245.200 91.700 ;
        RECT 246.000 91.600 246.800 92.400 ;
        RECT 247.600 91.600 248.400 92.400 ;
        RECT 249.200 91.600 250.000 92.400 ;
        RECT 254.000 91.600 254.800 92.400 ;
        RECT 249.300 86.400 249.900 91.600 ;
        RECT 254.100 90.400 254.700 91.600 ;
        RECT 254.000 89.600 254.800 90.400 ;
        RECT 257.300 88.400 257.900 93.600 ;
        RECT 258.800 90.200 259.400 93.600 ;
        RECT 262.800 93.400 263.600 93.600 ;
        RECT 258.800 89.400 259.600 90.200 ;
        RECT 260.400 89.600 261.200 90.400 ;
        RECT 265.600 90.200 266.200 95.000 ;
        RECT 268.500 94.400 269.100 97.600 ;
        RECT 266.800 93.600 267.600 94.400 ;
        RECT 268.400 93.600 269.200 94.400 ;
        RECT 265.400 89.400 266.200 90.200 ;
        RECT 257.200 87.600 258.000 88.400 ;
        RECT 249.200 85.600 250.000 86.400 ;
        RECT 244.400 73.600 245.200 74.400 ;
        RECT 270.000 73.600 270.800 74.400 ;
        RECT 244.400 71.600 245.200 72.400 ;
        RECT 247.600 71.600 248.400 72.400 ;
        RECT 250.800 71.600 251.600 72.400 ;
        RECT 254.000 71.600 254.800 72.400 ;
        RECT 258.800 71.600 259.600 72.400 ;
        RECT 260.400 71.600 261.200 72.400 ;
        RECT 244.500 64.400 245.100 71.600 ;
        RECT 246.000 69.600 246.800 70.400 ;
        RECT 246.000 65.600 246.800 66.400 ;
        RECT 247.700 64.400 248.300 71.600 ;
        RECT 250.900 70.400 251.500 71.600 ;
        RECT 258.900 70.400 259.500 71.600 ;
        RECT 270.100 70.400 270.700 73.600 ;
        RECT 271.700 72.400 272.300 107.600 ;
        RECT 273.200 105.600 274.000 106.400 ;
        RECT 274.900 96.400 275.500 109.600 ;
        RECT 276.400 107.600 277.200 108.400 ;
        RECT 274.800 95.600 275.600 96.400 ;
        RECT 276.500 94.400 277.100 107.600 ;
        RECT 281.300 106.400 281.900 111.600 ;
        RECT 282.900 110.400 283.500 133.700 ;
        RECT 284.400 133.600 285.200 134.400 ;
        RECT 294.000 133.600 294.800 134.400 ;
        RECT 295.600 133.600 296.400 134.400 ;
        RECT 297.200 134.200 297.800 135.000 ;
        RECT 298.600 134.800 299.400 135.000 ;
        RECT 302.000 134.800 302.800 135.000 ;
        RECT 297.200 133.600 302.800 134.200 ;
        RECT 284.500 132.400 285.100 133.600 ;
        RECT 284.400 131.600 285.200 132.400 ;
        RECT 289.200 129.600 290.000 130.400 ;
        RECT 297.200 130.200 297.800 133.600 ;
        RECT 298.800 131.600 299.600 132.400 ;
        RECT 302.200 132.200 302.800 133.600 ;
        RECT 297.200 129.400 298.000 130.200 ;
        RECT 289.200 113.600 290.000 114.400 ;
        RECT 284.400 111.800 285.200 112.600 ;
        RECT 291.000 111.800 291.800 112.600 ;
        RECT 282.800 109.600 283.600 110.400 ;
        RECT 284.400 108.400 285.000 111.800 ;
        RECT 288.400 108.400 289.200 108.600 ;
        RECT 282.800 107.600 283.600 108.400 ;
        RECT 284.400 107.800 289.200 108.400 ;
        RECT 281.200 105.600 282.000 106.400 ;
        RECT 282.900 104.400 283.500 107.600 ;
        RECT 284.400 107.000 285.000 107.800 ;
        RECT 285.800 107.000 286.600 107.200 ;
        RECT 289.200 107.000 290.000 107.200 ;
        RECT 291.200 107.000 291.800 111.800 ;
        RECT 297.200 109.600 298.000 110.400 ;
        RECT 292.400 107.600 293.200 108.400 ;
        RECT 284.400 106.200 285.200 107.000 ;
        RECT 285.800 106.400 290.000 107.000 ;
        RECT 291.000 106.200 291.800 107.000 ;
        RECT 292.500 104.400 293.100 107.600 ;
        RECT 282.800 103.600 283.600 104.400 ;
        RECT 292.400 103.600 293.200 104.400 ;
        RECT 287.600 101.600 288.400 102.400 ;
        RECT 287.700 98.400 288.300 101.600 ;
        RECT 287.600 97.600 288.400 98.400 ;
        RECT 282.800 95.600 283.600 96.400 ;
        RECT 276.400 93.600 277.200 94.400 ;
        RECT 282.900 92.400 283.500 95.600 ;
        RECT 297.300 94.400 297.900 109.600 ;
        RECT 298.900 108.400 299.500 131.600 ;
        RECT 302.200 131.400 303.000 132.200 ;
        RECT 303.600 130.200 304.200 135.000 ;
        RECT 305.200 133.600 306.000 134.400 ;
        RECT 306.800 130.200 307.600 135.800 ;
        RECT 308.500 134.400 309.100 153.600 ;
        RECT 313.200 146.200 314.000 151.800 ;
        RECT 314.800 147.600 315.600 148.400 ;
        RECT 311.600 143.600 312.400 144.400 ;
        RECT 311.700 142.400 312.300 143.600 ;
        RECT 311.600 141.600 312.400 142.400 ;
        RECT 308.400 133.600 309.200 134.400 ;
        RECT 303.400 129.400 304.200 130.200 ;
        RECT 306.800 125.600 307.600 126.400 ;
        RECT 310.000 126.200 310.800 137.800 ;
        RECT 314.900 134.400 315.500 147.600 ;
        RECT 316.400 144.200 317.200 155.800 ;
        RECT 318.000 149.400 318.800 150.400 ;
        RECT 319.700 146.300 320.300 169.600 ;
        RECT 330.900 168.400 331.500 173.600 ;
        RECT 332.500 170.400 333.100 175.600 ;
        RECT 337.200 173.600 338.000 174.400 ;
        RECT 337.300 172.400 337.900 173.600 ;
        RECT 337.200 172.300 338.000 172.400 ;
        RECT 338.900 172.300 339.500 191.600 ;
        RECT 342.000 187.600 342.800 188.400 ;
        RECT 343.700 186.400 344.300 191.600 ;
        RECT 346.800 188.400 347.400 191.800 ;
        RECT 350.800 188.400 351.600 188.600 ;
        RECT 345.200 187.600 346.000 188.400 ;
        RECT 346.800 187.800 351.600 188.400 ;
        RECT 343.600 185.600 344.400 186.400 ;
        RECT 343.600 179.600 344.400 180.400 ;
        RECT 340.400 175.600 341.200 176.400 ;
        RECT 342.000 173.600 342.800 174.400 ;
        RECT 337.200 171.700 339.500 172.300 ;
        RECT 337.200 171.600 338.000 171.700 ;
        RECT 342.100 170.400 342.700 173.600 ;
        RECT 343.700 172.400 344.300 179.600 ;
        RECT 345.300 176.400 345.900 187.600 ;
        RECT 346.800 187.000 347.400 187.800 ;
        RECT 348.200 187.000 349.000 187.200 ;
        RECT 351.600 187.000 352.400 187.200 ;
        RECT 353.600 187.000 354.200 191.800 ;
        RECT 354.800 187.600 355.600 188.400 ;
        RECT 346.800 186.200 347.600 187.000 ;
        RECT 348.200 186.400 352.400 187.000 ;
        RECT 353.400 186.200 354.200 187.000 ;
        RECT 356.400 186.200 357.200 191.800 ;
        RECT 358.100 188.400 358.700 211.600 ;
        RECT 359.600 206.200 360.400 217.800 ;
        RECT 364.400 217.700 366.700 218.300 ;
        RECT 364.400 217.600 365.200 217.700 ;
        RECT 366.100 216.400 366.700 217.700 ;
        RECT 370.800 217.600 371.600 218.400 ;
        RECT 388.400 217.600 389.200 218.400 ;
        RECT 407.600 217.600 408.400 218.400 ;
        RECT 366.000 215.600 366.800 216.400 ;
        RECT 366.100 214.400 366.700 215.600 ;
        RECT 366.000 213.600 366.800 214.400 ;
        RECT 370.900 212.400 371.500 217.600 ;
        RECT 380.400 215.600 381.200 216.400 ;
        RECT 383.800 215.600 384.600 215.800 ;
        RECT 383.800 215.000 389.400 215.600 ;
        RECT 390.000 215.000 390.800 215.800 ;
        RECT 393.200 215.600 394.000 216.400 ;
        RECT 375.600 213.600 376.400 214.400 ;
        RECT 382.000 213.600 382.800 214.400 ;
        RECT 370.800 211.600 371.600 212.400 ;
        RECT 377.200 211.600 378.000 212.400 ;
        RECT 374.000 209.600 374.800 210.400 ;
        RECT 380.400 209.600 381.200 210.400 ;
        RECT 370.800 207.600 371.600 208.400 ;
        RECT 374.100 198.400 374.700 209.600 ;
        RECT 382.100 208.300 382.700 213.600 ;
        RECT 383.800 210.200 384.400 215.000 ;
        RECT 385.200 214.800 386.000 215.000 ;
        RECT 388.600 214.800 389.400 215.000 ;
        RECT 390.200 214.200 390.800 215.000 ;
        RECT 404.400 215.000 405.200 215.800 ;
        RECT 405.800 215.000 410.000 215.600 ;
        RECT 411.000 215.000 411.800 215.800 ;
        RECT 385.200 213.600 390.800 214.200 ;
        RECT 393.200 213.600 394.000 214.400 ;
        RECT 401.200 213.600 402.000 214.400 ;
        RECT 402.800 213.600 403.600 214.400 ;
        RECT 404.400 214.200 405.000 215.000 ;
        RECT 405.800 214.800 406.600 215.000 ;
        RECT 409.200 214.800 410.000 215.000 ;
        RECT 404.400 213.600 409.200 214.200 ;
        RECT 385.200 212.200 385.800 213.600 ;
        RECT 385.000 211.400 385.800 212.200 ;
        RECT 390.200 210.200 390.800 213.600 ;
        RECT 383.800 209.400 384.600 210.200 ;
        RECT 390.000 209.400 390.800 210.200 ;
        RECT 380.500 207.700 382.700 208.300 ;
        RECT 380.500 198.400 381.100 207.700 ;
        RECT 393.300 198.400 393.900 213.600 ;
        RECT 396.400 211.600 397.200 212.400 ;
        RECT 399.600 211.600 400.400 212.400 ;
        RECT 396.400 209.600 397.200 210.400 ;
        RECT 399.600 209.600 400.400 210.400 ;
        RECT 396.500 208.400 397.100 209.600 ;
        RECT 396.400 207.600 397.200 208.400 ;
        RECT 401.300 198.400 401.900 213.600 ;
        RECT 402.900 198.400 403.500 213.600 ;
        RECT 404.400 210.200 405.000 213.600 ;
        RECT 408.400 213.400 409.200 213.600 ;
        RECT 411.200 210.200 411.800 215.000 ;
        RECT 412.400 213.600 413.200 214.400 ;
        RECT 412.500 212.400 413.100 213.600 ;
        RECT 412.400 211.600 413.200 212.400 ;
        RECT 414.000 210.200 414.800 215.800 ;
        RECT 415.700 214.400 416.300 221.700 ;
        RECT 441.300 218.400 441.900 233.600 ;
        RECT 466.900 232.400 467.500 239.600 ;
        RECT 442.800 231.600 443.600 232.400 ;
        RECT 444.400 231.600 445.200 232.400 ;
        RECT 452.400 231.600 453.200 232.400 ;
        RECT 458.800 231.600 459.600 232.400 ;
        RECT 465.200 231.600 466.000 232.400 ;
        RECT 466.800 231.600 467.600 232.400 ;
        RECT 442.900 230.400 443.500 231.600 ;
        RECT 442.800 229.600 443.600 230.400 ;
        RECT 444.500 226.400 445.100 231.600 ;
        RECT 452.500 230.400 453.100 231.600 ;
        RECT 449.200 229.600 450.000 230.400 ;
        RECT 452.400 229.600 453.200 230.400 ;
        RECT 444.400 225.600 445.200 226.400 ;
        RECT 442.800 219.600 443.600 220.400 ;
        RECT 415.600 213.600 416.400 214.400 ;
        RECT 415.600 211.600 416.400 212.400 ;
        RECT 404.400 209.400 405.200 210.200 ;
        RECT 411.000 209.400 411.800 210.200 ;
        RECT 410.800 207.600 411.600 208.400 ;
        RECT 374.000 197.600 374.800 198.400 ;
        RECT 380.400 197.600 381.200 198.400 ;
        RECT 393.200 197.600 394.000 198.400 ;
        RECT 401.200 197.600 402.000 198.400 ;
        RECT 402.800 197.600 403.600 198.400 ;
        RECT 409.200 197.600 410.000 198.400 ;
        RECT 358.000 187.600 358.800 188.400 ;
        RECT 351.600 183.600 352.400 184.400 ;
        RECT 359.600 184.200 360.400 195.800 ;
        RECT 361.200 189.400 362.000 190.200 ;
        RECT 351.700 178.400 352.300 183.600 ;
        RECT 361.300 180.400 361.900 189.400 ;
        RECT 369.200 184.200 370.000 195.800 ;
        RECT 393.300 190.400 393.900 197.600 ;
        RECT 372.400 189.600 373.200 190.400 ;
        RECT 377.200 189.600 378.000 190.400 ;
        RECT 382.000 189.600 382.800 190.400 ;
        RECT 383.600 189.600 384.400 190.400 ;
        RECT 385.200 189.600 386.000 190.400 ;
        RECT 388.400 189.600 389.200 190.400 ;
        RECT 393.200 189.600 394.000 190.400 ;
        RECT 396.400 190.300 397.200 190.400 ;
        RECT 394.900 189.700 397.200 190.300 ;
        RECT 361.200 179.600 362.000 180.400 ;
        RECT 372.500 178.400 373.100 189.600 ;
        RECT 378.800 185.600 379.600 186.400 ;
        RECT 374.000 183.600 374.800 184.400 ;
        RECT 374.100 180.400 374.700 183.600 ;
        RECT 374.000 179.600 374.800 180.400 ;
        RECT 378.900 178.400 379.500 185.600 ;
        RECT 383.700 178.400 384.300 189.600 ;
        RECT 385.300 188.400 385.900 189.600 ;
        RECT 388.500 188.400 389.100 189.600 ;
        RECT 385.200 187.600 386.000 188.400 ;
        RECT 388.400 187.600 389.200 188.400 ;
        RECT 390.000 187.600 390.800 188.400 ;
        RECT 390.100 178.400 390.700 187.600 ;
        RECT 391.600 185.600 392.400 186.400 ;
        RECT 391.600 181.600 392.400 182.400 ;
        RECT 351.600 177.600 352.400 178.400 ;
        RECT 372.400 177.600 373.200 178.400 ;
        RECT 374.000 177.600 374.800 178.400 ;
        RECT 378.800 177.600 379.600 178.400 ;
        RECT 383.600 177.600 384.400 178.400 ;
        RECT 390.000 177.600 390.800 178.400 ;
        RECT 345.200 175.600 346.000 176.400 ;
        RECT 356.400 175.600 357.200 176.400 ;
        RECT 362.800 175.600 363.600 176.400 ;
        RECT 364.400 175.600 365.200 176.400 ;
        RECT 369.200 175.600 370.000 176.400 ;
        RECT 356.500 174.400 357.100 175.600 ;
        RECT 348.400 173.600 349.200 174.400 ;
        RECT 356.400 173.600 357.200 174.400 ;
        RECT 361.200 173.600 362.000 174.400 ;
        RECT 361.300 172.400 361.900 173.600 ;
        RECT 364.500 172.400 365.100 175.600 ;
        RECT 366.000 173.600 366.800 174.400 ;
        RECT 343.600 171.600 344.400 172.400 ;
        RECT 348.400 171.600 349.200 172.400 ;
        RECT 353.200 171.600 354.000 172.400 ;
        RECT 361.200 171.600 362.000 172.400 ;
        RECT 364.400 171.600 365.200 172.400 ;
        RECT 348.500 170.400 349.100 171.600 ;
        RECT 332.400 169.600 333.200 170.400 ;
        RECT 335.600 169.600 336.400 170.400 ;
        RECT 342.000 169.600 342.800 170.400 ;
        RECT 346.800 169.600 347.600 170.400 ;
        RECT 348.400 169.600 349.200 170.400 ;
        RECT 351.600 169.600 352.400 170.400 ;
        RECT 361.200 169.600 362.000 170.400 ;
        RECT 346.900 168.400 347.500 169.600 ;
        RECT 361.300 168.400 361.900 169.600 ;
        RECT 330.800 167.600 331.600 168.400 ;
        RECT 346.800 167.600 347.600 168.400 ;
        RECT 361.200 167.600 362.000 168.400 ;
        RECT 356.400 165.600 357.200 166.400 ;
        RECT 356.500 158.400 357.100 165.600 ;
        RECT 356.400 157.600 357.200 158.400 ;
        RECT 324.400 155.600 325.200 156.400 ;
        RECT 318.100 145.700 320.300 146.300 ;
        RECT 314.800 133.600 315.600 134.400 ;
        RECT 311.600 131.800 312.400 132.600 ;
        RECT 311.700 128.400 312.300 131.800 ;
        RECT 311.600 127.600 312.400 128.400 ;
        RECT 302.000 123.600 302.800 124.400 ;
        RECT 306.900 118.400 307.500 125.600 ;
        RECT 313.200 123.600 314.000 124.400 ;
        RECT 310.000 121.600 310.800 122.400 ;
        RECT 306.800 117.600 307.600 118.400 ;
        RECT 298.800 107.600 299.600 108.400 ;
        RECT 298.900 94.400 299.500 107.600 ;
        RECT 308.400 106.200 309.200 111.800 ;
        RECT 300.400 103.600 301.200 104.400 ;
        RECT 300.500 96.400 301.100 103.600 ;
        RECT 303.600 97.600 304.400 98.400 ;
        RECT 303.700 96.400 304.300 97.600 ;
        RECT 300.400 95.600 301.200 96.400 ;
        RECT 303.600 95.600 304.400 96.400 ;
        RECT 286.000 93.600 286.800 94.400 ;
        RECT 292.400 93.600 293.200 94.400 ;
        RECT 297.200 93.600 298.000 94.400 ;
        RECT 298.800 93.600 299.600 94.400 ;
        RECT 302.000 93.600 302.800 94.400 ;
        RECT 282.800 91.600 283.600 92.400 ;
        RECT 282.800 89.600 283.600 90.400 ;
        RECT 282.900 88.400 283.500 89.600 ;
        RECT 276.400 87.600 277.200 88.400 ;
        RECT 282.800 87.600 283.600 88.400 ;
        RECT 276.500 78.400 277.100 87.600 ;
        RECT 286.100 78.400 286.700 93.600 ;
        RECT 292.500 90.400 293.100 93.600 ;
        RECT 295.600 91.600 296.400 92.400 ;
        RECT 302.000 91.600 302.800 92.400 ;
        RECT 302.100 90.400 302.700 91.600 ;
        RECT 292.400 89.600 293.200 90.400 ;
        RECT 302.000 89.600 302.800 90.400 ;
        RECT 290.800 87.600 291.600 88.400 ;
        RECT 276.400 77.600 277.200 78.400 ;
        RECT 286.000 77.600 286.800 78.400 ;
        RECT 287.600 73.600 288.400 74.400 ;
        RECT 271.600 71.600 272.400 72.400 ;
        RECT 273.200 71.600 274.000 72.400 ;
        RECT 284.400 71.600 285.200 72.400 ;
        RECT 286.000 71.600 286.800 72.400 ;
        RECT 250.800 69.600 251.600 70.400 ;
        RECT 254.000 69.600 254.800 70.400 ;
        RECT 258.800 69.600 259.600 70.400 ;
        RECT 268.400 69.600 269.200 70.400 ;
        RECT 270.000 69.600 270.800 70.400 ;
        RECT 254.100 68.400 254.700 69.600 ;
        RECT 268.500 68.400 269.100 69.600 ;
        RECT 249.200 67.600 250.000 68.400 ;
        RECT 254.000 67.600 254.800 68.400 ;
        RECT 255.600 67.600 256.400 68.400 ;
        RECT 266.800 67.600 267.600 68.400 ;
        RECT 268.400 67.600 269.200 68.400 ;
        RECT 255.700 66.400 256.300 67.600 ;
        RECT 255.600 65.600 256.400 66.400 ;
        RECT 262.000 65.600 262.800 66.400 ;
        RECT 263.600 65.600 264.400 66.400 ;
        RECT 262.100 64.400 262.700 65.600 ;
        RECT 244.400 63.600 245.200 64.400 ;
        RECT 247.600 63.600 248.400 64.400 ;
        RECT 258.800 63.600 259.600 64.400 ;
        RECT 262.000 63.600 262.800 64.400 ;
        RECT 247.700 58.400 248.300 63.600 ;
        RECT 239.600 57.600 240.400 58.400 ;
        RECT 242.800 57.600 243.600 58.400 ;
        RECT 247.600 57.600 248.400 58.400 ;
        RECT 239.700 50.400 240.300 57.600 ;
        RECT 241.200 55.600 242.000 56.400 ;
        RECT 241.300 54.400 241.900 55.600 ;
        RECT 242.600 55.000 243.400 55.800 ;
        RECT 244.400 55.000 248.600 55.600 ;
        RECT 249.200 55.000 250.000 55.800 ;
        RECT 241.200 53.600 242.000 54.400 ;
        RECT 236.400 49.600 237.200 50.400 ;
        RECT 239.600 49.600 240.400 50.400 ;
        RECT 242.600 50.200 243.200 55.000 ;
        RECT 244.400 54.800 245.200 55.000 ;
        RECT 247.800 54.800 248.600 55.000 ;
        RECT 249.400 54.200 250.000 55.000 ;
        RECT 258.900 54.400 259.500 63.600 ;
        RECT 266.900 58.400 267.500 67.600 ;
        RECT 273.300 64.400 273.900 71.600 ;
        RECT 286.100 70.400 286.700 71.600 ;
        RECT 287.700 70.400 288.300 73.600 ;
        RECT 303.700 70.400 304.300 95.600 ;
        RECT 306.800 93.600 307.600 94.400 ;
        RECT 310.100 90.400 310.700 121.600 ;
        RECT 311.600 104.200 312.400 115.800 ;
        RECT 313.300 110.200 313.900 123.600 ;
        RECT 313.200 109.400 314.000 110.200 ;
        RECT 314.900 108.400 315.500 133.600 ;
        RECT 318.100 132.400 318.700 145.700 ;
        RECT 324.500 138.400 325.100 155.600 ;
        RECT 326.000 144.200 326.800 155.800 ;
        RECT 364.500 154.400 365.100 171.600 ;
        RECT 369.300 168.400 369.900 175.600 ;
        RECT 374.100 174.400 374.700 177.600 ;
        RECT 377.200 175.600 378.000 176.400 ;
        RECT 377.300 174.400 377.900 175.600 ;
        RECT 372.400 173.600 373.200 174.400 ;
        RECT 374.000 173.600 374.800 174.400 ;
        RECT 377.200 173.600 378.000 174.400 ;
        RECT 382.000 173.600 382.800 174.400 ;
        RECT 386.800 173.600 387.600 174.400 ;
        RECT 369.200 168.300 370.000 168.400 ;
        RECT 367.700 167.700 370.000 168.300 ;
        RECT 364.400 153.600 365.200 154.400 ;
        RECT 367.700 152.400 368.300 167.700 ;
        RECT 369.200 167.600 370.000 167.700 ;
        RECT 370.800 155.600 371.600 156.400 ;
        RECT 369.200 153.600 370.000 154.400 ;
        RECT 351.600 151.600 352.400 152.400 ;
        RECT 367.600 151.600 368.400 152.400 ;
        RECT 348.400 149.600 349.200 150.400 ;
        RECT 346.800 147.600 347.600 148.400 ;
        RECT 346.900 146.400 347.500 147.600 ;
        RECT 330.800 145.600 331.600 146.400 ;
        RECT 337.200 145.600 338.000 146.400 ;
        RECT 346.800 145.600 347.600 146.400 ;
        RECT 330.900 144.400 331.500 145.600 ;
        RECT 330.800 143.600 331.600 144.400 ;
        RECT 326.000 141.600 326.800 142.400 ;
        RECT 318.000 131.600 318.800 132.400 ;
        RECT 319.600 126.200 320.400 137.800 ;
        RECT 324.400 137.600 325.200 138.400 ;
        RECT 326.100 134.400 326.700 141.600 ;
        RECT 327.600 135.000 328.400 135.800 ;
        RECT 333.800 135.600 334.600 135.800 ;
        RECT 329.000 135.000 334.600 135.600 ;
        RECT 326.000 133.600 326.800 134.400 ;
        RECT 327.600 134.200 328.200 135.000 ;
        RECT 329.000 134.800 329.800 135.000 ;
        RECT 332.400 134.800 333.200 135.000 ;
        RECT 327.600 133.600 333.200 134.200 ;
        RECT 327.600 130.200 328.200 133.600 ;
        RECT 332.600 132.200 333.200 133.600 ;
        RECT 332.600 131.400 333.400 132.200 ;
        RECT 334.000 130.200 334.600 135.000 ;
        RECT 337.300 134.400 337.900 145.600 ;
        RECT 343.600 143.600 344.400 144.400 ;
        RECT 343.700 138.400 344.300 143.600 ;
        RECT 348.500 142.400 349.100 149.600 ;
        RECT 351.700 142.400 352.300 151.600 ;
        RECT 356.400 149.600 357.200 150.400 ;
        RECT 364.400 149.600 365.200 150.400 ;
        RECT 367.600 149.600 368.400 150.400 ;
        RECT 354.800 147.600 355.600 148.400 ;
        RECT 348.400 141.600 349.200 142.400 ;
        RECT 351.600 141.600 352.400 142.400 ;
        RECT 343.600 137.600 344.400 138.400 ;
        RECT 338.800 135.000 339.600 135.800 ;
        RECT 345.000 135.600 345.800 135.800 ;
        RECT 340.200 135.000 345.800 135.600 ;
        RECT 335.600 133.600 336.400 134.400 ;
        RECT 337.200 133.600 338.000 134.400 ;
        RECT 338.800 134.200 339.400 135.000 ;
        RECT 340.200 134.800 341.000 135.000 ;
        RECT 343.600 134.800 344.400 135.000 ;
        RECT 338.800 133.600 344.400 134.200 ;
        RECT 327.600 129.400 328.400 130.200 ;
        RECT 333.800 129.400 334.600 130.200 ;
        RECT 338.800 130.200 339.400 133.600 ;
        RECT 343.800 132.200 344.400 133.600 ;
        RECT 343.800 131.400 344.600 132.200 ;
        RECT 338.800 129.400 339.600 130.200 ;
        RECT 343.600 129.600 344.400 130.400 ;
        RECT 345.200 130.200 345.800 135.000 ;
        RECT 349.800 135.000 350.600 135.800 ;
        RECT 354.900 135.600 355.500 147.600 ;
        RECT 356.500 144.400 357.100 149.600 ;
        RECT 362.800 147.600 363.600 148.400 ;
        RECT 362.900 146.400 363.500 147.600 ;
        RECT 358.000 145.600 358.800 146.400 ;
        RECT 361.200 145.600 362.000 146.400 ;
        RECT 362.800 145.600 363.600 146.400 ;
        RECT 356.400 143.600 357.200 144.400 ;
        RECT 358.100 136.400 358.700 145.600 ;
        RECT 351.600 135.000 355.800 135.600 ;
        RECT 356.400 135.000 357.200 135.800 ;
        RECT 358.000 135.600 358.800 136.400 ;
        RECT 348.400 133.600 349.200 134.400 ;
        RECT 345.000 129.400 345.800 130.200 ;
        RECT 345.200 127.600 346.000 128.400 ;
        RECT 332.400 125.600 333.200 126.400 ;
        RECT 345.300 118.400 345.900 127.600 ;
        RECT 348.500 118.400 349.100 133.600 ;
        RECT 349.800 130.200 350.400 135.000 ;
        RECT 351.600 134.800 352.400 135.000 ;
        RECT 355.000 134.800 355.800 135.000 ;
        RECT 356.600 134.200 357.200 135.000 ;
        RECT 358.100 134.400 358.700 135.600 ;
        RECT 361.300 134.400 361.900 145.600 ;
        RECT 362.800 141.600 363.600 142.400 ;
        RECT 352.400 133.600 357.200 134.200 ;
        RECT 358.000 133.600 358.800 134.400 ;
        RECT 361.200 133.600 362.000 134.400 ;
        RECT 352.400 133.400 353.200 133.600 ;
        RECT 354.800 131.600 355.600 132.400 ;
        RECT 356.600 130.200 357.200 133.600 ;
        RECT 358.000 131.600 358.800 132.400 ;
        RECT 349.800 129.400 350.600 130.200 ;
        RECT 356.400 129.400 357.200 130.200 ;
        RECT 356.400 127.600 357.200 128.400 ;
        RECT 356.500 118.400 357.100 127.600 ;
        RECT 345.200 117.600 346.000 118.400 ;
        RECT 348.400 117.600 349.200 118.400 ;
        RECT 356.400 117.600 357.200 118.400 ;
        RECT 314.800 107.600 315.600 108.400 ;
        RECT 321.200 104.200 322.000 115.800 ;
        RECT 327.600 106.200 328.400 111.800 ;
        RECT 329.200 107.600 330.000 108.400 ;
        RECT 326.000 103.600 326.800 104.400 ;
        RECT 330.800 104.200 331.600 115.800 ;
        RECT 332.400 113.600 333.200 114.400 ;
        RECT 332.500 110.200 333.100 113.600 ;
        RECT 332.400 109.400 333.200 110.200 ;
        RECT 340.400 104.200 341.200 115.800 ;
        RECT 351.600 110.300 352.400 110.400 ;
        RECT 350.100 109.700 352.400 110.300 ;
        RECT 326.100 102.400 326.700 103.600 ;
        RECT 326.000 101.600 326.800 102.400 ;
        RECT 310.000 89.600 310.800 90.400 ;
        RECT 311.600 90.200 312.400 95.800 ;
        RECT 314.800 86.200 315.600 97.800 ;
        RECT 316.400 91.800 317.200 92.600 ;
        RECT 316.500 90.400 317.100 91.800 ;
        RECT 322.800 91.600 323.600 92.400 ;
        RECT 316.400 89.600 317.200 90.400 ;
        RECT 324.400 86.200 325.200 97.800 ;
        RECT 330.800 90.200 331.600 95.800 ;
        RECT 334.000 86.200 334.800 97.800 ;
        RECT 335.600 91.800 336.400 92.600 ;
        RECT 335.700 88.400 336.300 91.800 ;
        RECT 342.000 91.600 342.800 92.400 ;
        RECT 335.600 87.600 336.400 88.400 ;
        RECT 343.600 86.200 344.400 97.800 ;
        RECT 350.100 92.400 350.700 109.700 ;
        RECT 351.600 109.600 352.400 109.700 ;
        RECT 356.400 103.600 357.200 104.400 ;
        RECT 356.400 101.600 357.200 102.400 ;
        RECT 356.500 96.400 357.100 101.600 ;
        RECT 356.400 95.600 357.200 96.400 ;
        RECT 358.100 94.400 358.700 131.600 ;
        RECT 362.900 114.400 363.500 141.600 ;
        RECT 364.500 138.400 365.100 149.600 ;
        RECT 369.300 148.400 369.900 153.600 ;
        RECT 370.900 150.400 371.500 155.600 ;
        RECT 370.800 149.600 371.600 150.400 ;
        RECT 372.500 148.400 373.100 173.600 ;
        RECT 374.100 170.400 374.700 173.600 ;
        RECT 382.100 172.400 382.700 173.600 ;
        RECT 386.900 172.400 387.500 173.600 ;
        RECT 375.600 171.600 376.400 172.400 ;
        RECT 380.400 171.600 381.200 172.400 ;
        RECT 382.000 171.600 382.800 172.400 ;
        RECT 386.800 171.600 387.600 172.400 ;
        RECT 388.400 171.600 389.200 172.400 ;
        RECT 390.000 171.600 390.800 172.400 ;
        RECT 374.000 169.600 374.800 170.400 ;
        RECT 374.100 154.400 374.700 169.600 ;
        RECT 375.700 166.400 376.300 171.600 ;
        RECT 380.500 170.400 381.100 171.600 ;
        RECT 388.500 170.400 389.100 171.600 ;
        RECT 391.700 170.400 392.300 181.600 ;
        RECT 394.900 178.400 395.500 189.700 ;
        RECT 396.400 189.600 397.200 189.700 ;
        RECT 407.600 189.600 408.400 190.400 ;
        RECT 406.000 187.600 406.800 188.400 ;
        RECT 399.600 185.600 400.400 186.400 ;
        RECT 401.200 185.600 402.000 186.400 ;
        RECT 404.400 185.600 405.200 186.400 ;
        RECT 399.700 182.400 400.300 185.600 ;
        RECT 399.600 181.600 400.400 182.400 ;
        RECT 401.300 178.400 401.900 185.600 ;
        RECT 404.500 178.400 405.100 185.600 ;
        RECT 394.800 177.600 395.600 178.400 ;
        RECT 401.200 177.600 402.000 178.400 ;
        RECT 404.400 177.600 405.200 178.400 ;
        RECT 393.200 175.600 394.000 176.400 ;
        RECT 396.400 175.600 397.200 176.400 ;
        RECT 393.300 170.400 393.900 175.600 ;
        RECT 396.500 174.400 397.100 175.600 ;
        RECT 406.100 174.400 406.700 187.600 ;
        RECT 407.600 185.600 408.400 186.400 ;
        RECT 407.700 176.300 408.300 185.600 ;
        RECT 409.200 176.300 410.000 176.400 ;
        RECT 407.700 175.700 410.000 176.300 ;
        RECT 409.200 175.600 410.000 175.700 ;
        RECT 396.400 173.600 397.200 174.400 ;
        RECT 406.000 173.600 406.800 174.400 ;
        RECT 406.100 172.400 406.700 173.600 ;
        RECT 401.200 171.600 402.000 172.400 ;
        RECT 406.000 171.600 406.800 172.400 ;
        RECT 401.300 170.400 401.900 171.600 ;
        RECT 380.400 169.600 381.200 170.400 ;
        RECT 385.200 169.600 386.000 170.400 ;
        RECT 388.400 169.600 389.200 170.400 ;
        RECT 391.600 169.600 392.400 170.400 ;
        RECT 393.200 169.600 394.000 170.400 ;
        RECT 396.400 169.600 397.200 170.400 ;
        RECT 399.600 169.600 400.400 170.400 ;
        RECT 401.200 169.600 402.000 170.400 ;
        RECT 377.200 167.600 378.000 168.400 ;
        RECT 375.600 165.600 376.400 166.400 ;
        RECT 375.700 158.400 376.300 165.600 ;
        RECT 375.600 157.600 376.400 158.400 ;
        RECT 375.600 155.600 376.400 156.400 ;
        RECT 374.000 153.600 374.800 154.400 ;
        RECT 374.000 151.600 374.800 152.400 ;
        RECT 375.700 150.400 376.300 155.600 ;
        RECT 375.600 149.600 376.400 150.400 ;
        RECT 369.200 147.600 370.000 148.400 ;
        RECT 372.400 147.600 373.200 148.400 ;
        RECT 375.600 147.600 376.400 148.400 ;
        RECT 374.000 145.600 374.800 146.400 ;
        RECT 377.300 144.300 377.900 167.600 ;
        RECT 380.500 156.400 381.100 169.600 ;
        RECT 385.300 168.400 385.900 169.600 ;
        RECT 391.700 168.400 392.300 169.600 ;
        RECT 385.200 167.600 386.000 168.400 ;
        RECT 391.600 167.600 392.400 168.400 ;
        RECT 406.000 167.600 406.800 168.400 ;
        RECT 398.000 163.600 398.800 164.400 ;
        RECT 404.400 163.600 405.200 164.400 ;
        RECT 398.100 160.400 398.700 163.600 ;
        RECT 398.000 159.600 398.800 160.400 ;
        RECT 402.800 159.600 403.600 160.400 ;
        RECT 398.000 157.600 398.800 158.400 ;
        RECT 380.400 155.600 381.200 156.400 ;
        RECT 380.400 153.600 381.200 154.400 ;
        RECT 380.500 152.400 381.100 153.600 ;
        RECT 380.400 151.600 381.200 152.400 ;
        RECT 382.000 151.600 382.800 152.400 ;
        RECT 385.200 151.600 386.000 152.400 ;
        RECT 388.400 151.600 389.200 152.400 ;
        RECT 380.400 147.600 381.200 148.400 ;
        RECT 382.100 146.400 382.700 151.600 ;
        RECT 388.500 150.400 389.100 151.600 ;
        RECT 398.100 150.400 398.700 157.600 ;
        RECT 385.200 149.600 386.000 150.400 ;
        RECT 388.400 149.600 389.200 150.400 ;
        RECT 391.600 149.600 392.400 150.400 ;
        RECT 398.000 149.600 398.800 150.400 ;
        RECT 382.000 145.600 382.800 146.400 ;
        RECT 385.300 144.400 385.900 149.600 ;
        RECT 386.800 147.600 387.600 148.400 ;
        RECT 390.000 147.600 390.800 148.400 ;
        RECT 375.700 143.700 377.900 144.300 ;
        RECT 374.000 139.600 374.800 140.400 ;
        RECT 364.400 137.600 365.200 138.400 ;
        RECT 369.200 137.600 370.000 138.400 ;
        RECT 370.800 137.600 371.600 138.400 ;
        RECT 364.500 130.400 365.100 137.600 ;
        RECT 369.300 136.400 369.900 137.600 ;
        RECT 369.200 135.600 370.000 136.400 ;
        RECT 367.600 133.600 368.400 134.400 ;
        RECT 372.400 133.600 373.200 134.400 ;
        RECT 367.700 130.400 368.300 133.600 ;
        RECT 364.400 129.600 365.200 130.400 ;
        RECT 367.600 129.600 368.400 130.400 ;
        RECT 366.000 127.600 366.800 128.400 ;
        RECT 362.800 113.600 363.600 114.400 ;
        RECT 367.600 111.600 368.400 112.400 ;
        RECT 370.800 111.600 371.600 112.400 ;
        RECT 367.700 110.400 368.300 111.600 ;
        RECT 359.600 109.600 360.400 110.400 ;
        RECT 367.600 109.600 368.400 110.400 ;
        RECT 366.000 107.600 366.800 108.400 ;
        RECT 374.100 98.400 374.700 139.600 ;
        RECT 375.700 134.400 376.300 143.700 ;
        RECT 380.400 143.600 381.200 144.400 ;
        RECT 385.200 143.600 386.000 144.400 ;
        RECT 380.500 138.400 381.100 143.600 ;
        RECT 380.400 137.600 381.200 138.400 ;
        RECT 383.600 137.600 384.400 138.400 ;
        RECT 386.800 137.600 387.600 138.400 ;
        RECT 377.200 135.600 378.000 136.400 ;
        RECT 378.800 135.600 379.600 136.400 ;
        RECT 375.600 133.600 376.400 134.400 ;
        RECT 383.700 130.400 384.300 137.600 ;
        RECT 386.800 135.600 387.600 136.400 ;
        RECT 388.400 135.600 389.200 136.400 ;
        RECT 385.200 133.600 386.000 134.400 ;
        RECT 385.300 132.400 385.900 133.600 ;
        RECT 385.200 131.600 386.000 132.400 ;
        RECT 380.400 129.600 381.200 130.400 ;
        RECT 383.600 129.600 384.400 130.400 ;
        RECT 382.000 123.600 382.800 124.400 ;
        RECT 380.400 117.600 381.200 118.400 ;
        RECT 380.500 110.400 381.100 117.600 ;
        RECT 382.100 112.400 382.700 123.600 ;
        RECT 382.000 111.600 382.800 112.400 ;
        RECT 375.600 109.600 376.400 110.400 ;
        RECT 378.800 109.600 379.600 110.400 ;
        RECT 380.400 109.600 381.200 110.400 ;
        RECT 378.900 106.400 379.500 109.600 ;
        RECT 378.800 105.600 379.600 106.400 ;
        RECT 378.800 101.600 379.600 102.400 ;
        RECT 366.000 97.600 366.800 98.400 ;
        RECT 374.000 97.600 374.800 98.400 ;
        RECT 366.100 94.400 366.700 97.600 ;
        RECT 378.900 96.400 379.500 101.600 ;
        RECT 369.200 95.000 370.000 95.800 ;
        RECT 375.400 95.600 376.200 95.800 ;
        RECT 378.800 95.600 379.600 96.400 ;
        RECT 370.600 95.000 376.200 95.600 ;
        RECT 358.000 93.600 358.800 94.400 ;
        RECT 366.000 93.600 366.800 94.400 ;
        RECT 369.200 94.200 369.800 95.000 ;
        RECT 370.600 94.800 371.400 95.000 ;
        RECT 374.000 94.800 374.800 95.000 ;
        RECT 369.200 93.600 374.800 94.200 ;
        RECT 350.000 91.600 350.800 92.400 ;
        RECT 367.600 91.600 368.400 92.400 ;
        RECT 345.200 87.600 346.000 88.400 ;
        RECT 348.400 88.300 349.200 88.400 ;
        RECT 350.100 88.300 350.700 91.600 ;
        RECT 369.200 90.200 369.800 93.600 ;
        RECT 374.200 92.200 374.800 93.600 ;
        RECT 374.200 91.400 375.000 92.200 ;
        RECT 375.600 90.200 376.200 95.000 ;
        RECT 377.200 93.600 378.000 94.400 ;
        RECT 369.200 89.400 370.000 90.200 ;
        RECT 375.400 89.400 376.200 90.200 ;
        RECT 377.300 88.400 377.900 93.600 ;
        RECT 348.400 87.700 350.700 88.300 ;
        RECT 348.400 87.600 349.200 87.700 ;
        RECT 377.200 87.600 378.000 88.400 ;
        RECT 308.400 83.600 309.200 84.400 ;
        RECT 329.200 83.600 330.000 84.400 ;
        RECT 308.500 72.400 309.100 83.600 ;
        RECT 329.300 74.400 329.900 83.600 ;
        RECT 316.400 73.600 317.200 74.400 ;
        RECT 329.200 73.600 330.000 74.400 ;
        RECT 306.800 71.600 307.600 72.400 ;
        RECT 308.400 71.600 309.200 72.400 ;
        RECT 276.400 69.600 277.200 70.400 ;
        RECT 282.800 70.300 283.600 70.400 ;
        RECT 282.800 69.700 285.100 70.300 ;
        RECT 282.800 69.600 283.600 69.700 ;
        RECT 273.200 63.600 274.000 64.400 ;
        RECT 273.200 59.600 274.000 60.400 ;
        RECT 260.400 57.600 261.200 58.400 ;
        RECT 266.800 57.600 267.600 58.400 ;
        RECT 245.200 53.600 250.000 54.200 ;
        RECT 250.800 53.600 251.600 54.400 ;
        RECT 255.600 53.600 256.400 54.400 ;
        RECT 258.800 53.600 259.600 54.400 ;
        RECT 245.200 53.400 246.000 53.600 ;
        RECT 249.400 50.200 250.000 53.600 ;
        RECT 252.400 51.600 253.200 52.400 ;
        RECT 242.600 49.400 243.400 50.200 ;
        RECT 249.200 49.400 250.000 50.200 ;
        RECT 252.500 44.400 253.100 51.600 ;
        RECT 255.700 50.400 256.300 53.600 ;
        RECT 258.800 51.600 259.600 52.400 ;
        RECT 255.600 49.600 256.400 50.400 ;
        RECT 252.400 43.600 253.200 44.400 ;
        RECT 254.000 39.600 254.800 40.400 ;
        RECT 254.100 38.400 254.700 39.600 ;
        RECT 247.600 37.600 248.400 38.400 ;
        RECT 254.000 37.600 254.800 38.400 ;
        RECT 233.200 35.600 234.000 36.400 ;
        RECT 242.800 33.600 243.600 34.400 ;
        RECT 221.800 31.800 222.600 32.600 ;
        RECT 220.400 27.600 221.200 28.400 ;
        RECT 221.800 27.000 222.400 31.800 ;
        RECT 226.800 31.600 227.600 32.400 ;
        RECT 228.400 31.800 229.200 32.600 ;
        RECT 224.400 28.400 225.200 28.600 ;
        RECT 228.600 28.400 229.200 31.800 ;
        RECT 231.600 32.300 232.400 32.400 ;
        RECT 231.600 31.700 233.900 32.300 ;
        RECT 231.600 31.600 232.400 31.700 ;
        RECT 224.400 27.800 229.200 28.400 ;
        RECT 223.600 27.000 224.400 27.200 ;
        RECT 227.000 27.000 227.800 27.200 ;
        RECT 228.600 27.000 229.200 27.800 ;
        RECT 230.000 27.600 230.800 28.400 ;
        RECT 217.200 25.600 218.000 26.400 ;
        RECT 218.800 25.600 219.600 26.400 ;
        RECT 221.800 26.200 222.600 27.000 ;
        RECT 223.600 26.400 227.800 27.000 ;
        RECT 228.400 26.200 229.200 27.000 ;
        RECT 217.200 23.600 218.000 24.400 ;
        RECT 217.300 22.400 217.900 23.600 ;
        RECT 217.200 21.600 218.000 22.400 ;
        RECT 210.800 17.600 211.600 18.400 ;
        RECT 215.600 17.600 216.400 18.400 ;
        RECT 218.900 16.400 219.500 25.600 ;
        RECT 230.100 24.400 230.700 27.600 ;
        RECT 230.000 23.600 230.800 24.400 ;
        RECT 231.600 23.600 232.400 24.400 ;
        RECT 220.400 17.600 221.200 18.400 ;
        RECT 225.200 17.600 226.000 18.400 ;
        RECT 212.400 15.600 213.200 16.400 ;
        RECT 218.800 15.600 219.600 16.400 ;
        RECT 212.500 14.400 213.100 15.600 ;
        RECT 212.400 13.600 213.200 14.400 ;
        RECT 223.600 13.600 224.400 14.400 ;
        RECT 209.200 11.600 210.000 12.400 ;
        RECT 223.600 12.300 224.400 12.400 ;
        RECT 220.500 11.700 224.400 12.300 ;
        RECT 206.000 9.700 208.300 10.300 ;
        RECT 206.000 9.600 206.800 9.700 ;
        RECT 209.300 8.400 209.900 11.600 ;
        RECT 220.500 10.400 221.100 11.700 ;
        RECT 223.600 11.600 224.400 11.700 ;
        RECT 220.400 9.600 221.200 10.400 ;
        RECT 225.300 8.400 225.900 17.600 ;
        RECT 231.700 16.400 232.300 23.600 ;
        RECT 233.300 22.400 233.900 31.700 ;
        RECT 234.800 31.600 235.600 32.400 ;
        RECT 234.900 28.400 235.500 31.600 ;
        RECT 239.600 29.600 240.400 30.400 ;
        RECT 234.800 27.600 235.600 28.400 ;
        RECT 239.700 22.400 240.300 29.600 ;
        RECT 242.900 28.400 243.500 33.600 ;
        RECT 246.000 31.600 246.800 32.400 ;
        RECT 246.100 28.400 246.700 31.600 ;
        RECT 247.700 30.400 248.300 37.600 ;
        RECT 250.900 33.700 259.500 34.300 ;
        RECT 250.900 32.400 251.500 33.700 ;
        RECT 258.900 32.400 259.500 33.700 ;
        RECT 250.800 31.600 251.600 32.400 ;
        RECT 257.200 31.600 258.000 32.400 ;
        RECT 258.800 31.600 259.600 32.400 ;
        RECT 247.600 29.600 248.400 30.400 ;
        RECT 249.200 29.600 250.000 30.400 ;
        RECT 242.800 27.600 243.600 28.400 ;
        RECT 246.000 27.600 246.800 28.400 ;
        RECT 254.000 27.600 254.800 28.400 ;
        RECT 255.600 27.600 256.400 28.400 ;
        RECT 244.400 24.300 245.200 24.400 ;
        RECT 244.400 23.700 246.700 24.300 ;
        RECT 244.400 23.600 245.200 23.700 ;
        RECT 233.200 21.600 234.000 22.400 ;
        RECT 239.600 21.600 240.400 22.400 ;
        RECT 244.400 21.600 245.200 22.400 ;
        RECT 246.100 22.300 246.700 23.700 ;
        RECT 254.100 22.400 254.700 27.600 ;
        RECT 246.100 21.700 251.500 22.300 ;
        RECT 244.500 18.400 245.100 21.600 ;
        RECT 249.200 19.600 250.000 20.400 ;
        RECT 244.400 17.600 245.200 18.400 ;
        RECT 246.000 17.600 246.800 18.400 ;
        RECT 231.600 15.600 232.400 16.400 ;
        RECT 234.600 15.000 235.400 15.800 ;
        RECT 236.400 15.000 240.600 15.600 ;
        RECT 241.200 15.000 242.000 15.800 ;
        RECT 231.600 13.600 232.400 14.400 ;
        RECT 233.200 13.600 234.000 14.400 ;
        RECT 201.200 7.600 202.000 8.400 ;
        RECT 209.200 7.600 210.000 8.400 ;
        RECT 225.200 7.600 226.000 8.400 ;
        RECT 226.800 7.600 227.600 8.400 ;
        RECT 233.300 6.400 233.900 13.600 ;
        RECT 234.600 10.200 235.200 15.000 ;
        RECT 236.400 14.800 237.200 15.000 ;
        RECT 239.800 14.800 240.600 15.000 ;
        RECT 241.400 14.200 242.000 15.000 ;
        RECT 249.300 14.400 249.900 19.600 ;
        RECT 250.900 18.300 251.500 21.700 ;
        RECT 254.000 21.600 254.800 22.400 ;
        RECT 254.000 18.300 254.800 18.400 ;
        RECT 250.900 17.700 254.800 18.300 ;
        RECT 254.000 17.600 254.800 17.700 ;
        RECT 237.200 13.600 242.000 14.200 ;
        RECT 242.800 13.600 243.600 14.400 ;
        RECT 244.400 13.600 245.200 14.400 ;
        RECT 246.000 13.600 246.800 14.400 ;
        RECT 247.600 13.600 248.400 14.400 ;
        RECT 249.200 13.600 250.000 14.400 ;
        RECT 254.000 13.600 254.800 14.400 ;
        RECT 237.200 13.400 238.000 13.600 ;
        RECT 241.400 10.200 242.000 13.600 ;
        RECT 234.600 9.400 235.400 10.200 ;
        RECT 241.200 9.400 242.000 10.200 ;
        RECT 242.900 8.400 243.500 13.600 ;
        RECT 244.500 10.400 245.100 13.600 ;
        RECT 246.100 12.300 246.700 13.600 ;
        RECT 255.700 12.400 256.300 27.600 ;
        RECT 257.200 23.600 258.000 24.400 ;
        RECT 247.600 12.300 248.400 12.400 ;
        RECT 246.100 11.700 248.400 12.300 ;
        RECT 247.600 11.600 248.400 11.700 ;
        RECT 255.600 11.600 256.400 12.400 ;
        RECT 244.400 9.600 245.200 10.400 ;
        RECT 252.400 10.300 253.200 10.400 ;
        RECT 257.300 10.300 257.900 23.600 ;
        RECT 260.500 14.400 261.100 57.600 ;
        RECT 273.300 52.400 273.900 59.600 ;
        RECT 276.500 56.400 277.100 69.600 ;
        RECT 279.600 68.300 280.400 68.400 ;
        RECT 279.600 67.700 281.900 68.300 ;
        RECT 279.600 67.600 280.400 67.700 ;
        RECT 279.600 65.600 280.400 66.400 ;
        RECT 279.700 58.400 280.300 65.600 ;
        RECT 281.300 60.400 281.900 67.700 ;
        RECT 282.800 67.600 283.600 68.400 ;
        RECT 284.500 66.400 285.100 69.700 ;
        RECT 286.000 69.600 286.800 70.400 ;
        RECT 287.600 69.600 288.400 70.400 ;
        RECT 298.800 69.600 299.600 70.400 ;
        RECT 302.000 69.600 302.800 70.400 ;
        RECT 303.600 69.600 304.400 70.400 ;
        RECT 306.900 70.300 307.500 71.600 ;
        RECT 308.400 70.300 309.200 70.400 ;
        RECT 306.900 69.700 309.200 70.300 ;
        RECT 308.400 69.600 309.200 69.700 ;
        RECT 310.000 69.600 310.800 70.400 ;
        RECT 311.600 69.600 312.400 70.400 ;
        RECT 290.800 67.600 291.600 68.400 ;
        RECT 295.600 68.300 296.400 68.400 ;
        RECT 295.600 67.700 301.100 68.300 ;
        RECT 295.600 67.600 296.400 67.700 ;
        RECT 282.800 65.600 283.600 66.400 ;
        RECT 284.400 65.600 285.200 66.400 ;
        RECT 281.200 59.600 282.000 60.400 ;
        RECT 278.000 57.600 278.800 58.400 ;
        RECT 279.600 57.600 280.400 58.400 ;
        RECT 276.400 55.600 277.200 56.400 ;
        RECT 278.100 54.400 278.700 57.600 ;
        RECT 282.900 56.400 283.500 65.600 ;
        RECT 284.500 58.400 285.100 65.600 ;
        RECT 286.000 63.600 286.800 64.400 ;
        RECT 290.900 64.300 291.500 67.600 ;
        RECT 295.600 66.300 296.400 66.400 ;
        RECT 295.600 65.700 297.900 66.300 ;
        RECT 295.600 65.600 296.400 65.700 ;
        RECT 287.700 63.700 291.500 64.300 ;
        RECT 284.400 57.600 285.200 58.400 ;
        RECT 286.100 56.400 286.700 63.600 ;
        RECT 287.700 60.400 288.300 63.700 ;
        RECT 287.600 59.600 288.400 60.400 ;
        RECT 297.300 58.400 297.900 65.700 ;
        RECT 300.500 62.300 301.100 67.700 ;
        RECT 302.100 64.400 302.700 69.600 ;
        RECT 303.600 67.600 304.400 68.400 ;
        RECT 308.400 67.600 309.200 68.400 ;
        RECT 303.700 66.400 304.300 67.600 ;
        RECT 303.600 65.600 304.400 66.400 ;
        RECT 306.800 65.600 307.600 66.400 ;
        RECT 310.100 64.400 310.700 69.600 ;
        RECT 316.500 66.400 317.100 73.600 ;
        RECT 334.000 71.800 334.800 72.600 ;
        RECT 340.600 71.800 341.400 72.600 ;
        RECT 322.800 69.600 323.600 70.400 ;
        RECT 324.400 69.600 325.200 70.400 ;
        RECT 329.200 69.600 330.000 70.400 ;
        RECT 321.200 67.600 322.000 68.400 ;
        RECT 321.300 66.400 321.900 67.600 ;
        RECT 316.400 65.600 317.200 66.400 ;
        RECT 319.600 65.600 320.400 66.400 ;
        RECT 321.200 65.600 322.000 66.400 ;
        RECT 324.500 64.400 325.100 69.600 ;
        RECT 327.600 65.600 328.400 66.400 ;
        RECT 302.000 63.600 302.800 64.400 ;
        RECT 303.600 63.600 304.400 64.400 ;
        RECT 305.200 63.600 306.000 64.400 ;
        RECT 310.000 63.600 310.800 64.400 ;
        RECT 324.400 63.600 325.200 64.400 ;
        RECT 326.000 63.600 326.800 64.400 ;
        RECT 303.700 62.300 304.300 63.600 ;
        RECT 300.500 61.700 304.300 62.300 ;
        RECT 297.200 57.600 298.000 58.400 ;
        RECT 282.800 55.600 283.600 56.400 ;
        RECT 286.000 55.600 286.800 56.400 ;
        RECT 300.400 55.600 301.200 56.400 ;
        RECT 305.300 56.300 305.900 63.600 ;
        RECT 324.500 58.400 325.100 63.600 ;
        RECT 324.400 57.600 325.200 58.400 ;
        RECT 326.100 56.400 326.700 63.600 ;
        RECT 303.700 55.700 305.900 56.300 ;
        RECT 282.900 54.400 283.500 55.600 ;
        RECT 303.700 54.400 304.300 55.700 ;
        RECT 306.800 55.600 307.600 56.400 ;
        RECT 311.600 55.600 312.400 56.400 ;
        RECT 316.400 55.600 317.200 56.400 ;
        RECT 326.000 55.600 326.800 56.400 ;
        RECT 278.000 53.600 278.800 54.400 ;
        RECT 282.800 53.600 283.600 54.400 ;
        RECT 292.400 53.600 293.200 54.400 ;
        RECT 300.400 53.600 301.200 54.400 ;
        RECT 303.600 53.600 304.400 54.400 ;
        RECT 305.200 53.600 306.000 54.400 ;
        RECT 263.600 51.600 264.400 52.400 ;
        RECT 273.200 51.600 274.000 52.400 ;
        RECT 276.400 51.600 277.200 52.400 ;
        RECT 278.000 51.600 278.800 52.400 ;
        RECT 282.800 51.600 283.600 52.400 ;
        RECT 294.000 51.600 294.800 52.400 ;
        RECT 278.100 50.400 278.700 51.600 ;
        RECT 278.000 49.600 278.800 50.400 ;
        RECT 265.200 47.600 266.000 48.400 ;
        RECT 268.400 47.600 269.200 48.400 ;
        RECT 265.300 44.400 265.900 47.600 ;
        RECT 262.000 43.600 262.800 44.400 ;
        RECT 265.200 43.600 266.000 44.400 ;
        RECT 266.800 43.600 267.600 44.400 ;
        RECT 262.100 34.400 262.700 43.600 ;
        RECT 266.900 38.400 267.500 43.600 ;
        RECT 268.500 38.400 269.100 47.600 ;
        RECT 278.100 46.400 278.700 49.600 ;
        RECT 270.000 45.600 270.800 46.400 ;
        RECT 278.000 45.600 278.800 46.400 ;
        RECT 274.800 43.600 275.600 44.400 ;
        RECT 266.800 37.600 267.600 38.400 ;
        RECT 268.400 37.600 269.200 38.400 ;
        RECT 268.400 35.600 269.200 36.400 ;
        RECT 262.000 33.600 262.800 34.400 ;
        RECT 262.000 31.600 262.800 32.400 ;
        RECT 262.100 30.400 262.700 31.600 ;
        RECT 268.500 30.400 269.100 35.600 ;
        RECT 273.200 32.300 274.000 32.400 ;
        RECT 274.900 32.300 275.500 43.600 ;
        RECT 287.600 41.600 288.400 42.400 ;
        RECT 287.700 38.400 288.300 41.600 ;
        RECT 287.600 37.600 288.400 38.400 ;
        RECT 294.100 34.400 294.700 51.600 ;
        RECT 297.200 49.600 298.000 50.400 ;
        RECT 300.500 38.400 301.100 53.600 ;
        RECT 305.200 52.300 306.000 52.400 ;
        RECT 306.900 52.300 307.500 55.600 ;
        RECT 308.400 53.600 309.200 54.400 ;
        RECT 305.200 51.700 307.500 52.300 ;
        RECT 305.200 51.600 306.000 51.700 ;
        RECT 308.400 47.600 309.200 48.400 ;
        RECT 300.400 37.600 301.200 38.400 ;
        RECT 303.600 37.600 304.400 38.400 ;
        RECT 284.400 33.600 285.200 34.400 ;
        RECT 294.000 33.600 294.800 34.400 ;
        RECT 298.800 33.600 299.600 34.400 ;
        RECT 284.500 32.400 285.100 33.600 ;
        RECT 273.200 31.700 275.500 32.300 ;
        RECT 273.200 31.600 274.000 31.700 ;
        RECT 284.400 31.600 285.200 32.400 ;
        RECT 286.000 31.600 286.800 32.400 ;
        RECT 290.800 31.600 291.600 32.400 ;
        RECT 295.600 31.600 296.400 32.400 ;
        RECT 273.300 30.400 273.900 31.600 ;
        RECT 286.100 30.400 286.700 31.600 ;
        RECT 295.700 30.400 296.300 31.600 ;
        RECT 262.000 29.600 262.800 30.400 ;
        RECT 268.400 29.600 269.200 30.400 ;
        RECT 273.200 29.600 274.000 30.400 ;
        RECT 276.400 29.600 277.200 30.400 ;
        RECT 281.200 29.600 282.000 30.400 ;
        RECT 286.000 29.600 286.800 30.400 ;
        RECT 287.600 29.600 288.400 30.400 ;
        RECT 295.600 29.600 296.400 30.400 ;
        RECT 265.200 27.600 266.000 28.400 ;
        RECT 266.800 27.600 267.600 28.400 ;
        RECT 265.300 24.400 265.900 27.600 ;
        RECT 276.500 24.400 277.100 29.600 ;
        RECT 278.000 27.600 278.800 28.400 ;
        RECT 278.100 26.400 278.700 27.600 ;
        RECT 278.000 25.600 278.800 26.400 ;
        RECT 265.200 23.600 266.000 24.400 ;
        RECT 276.400 23.600 277.200 24.400 ;
        RECT 265.200 19.600 266.000 20.400 ;
        RECT 263.600 15.600 264.400 16.400 ;
        RECT 260.400 13.600 261.200 14.400 ;
        RECT 263.700 10.400 264.300 15.600 ;
        RECT 265.300 14.400 265.900 19.600 ;
        RECT 281.300 18.400 281.900 29.600 ;
        RECT 286.000 27.600 286.800 28.400 ;
        RECT 287.700 18.400 288.300 29.600 ;
        RECT 297.200 27.600 298.000 28.400 ;
        RECT 281.200 17.600 282.000 18.400 ;
        RECT 287.600 17.600 288.400 18.400 ;
        RECT 289.200 17.600 290.000 18.400 ;
        RECT 297.300 16.400 297.900 27.600 ;
        RECT 266.800 15.000 267.600 15.800 ;
        RECT 268.200 15.000 272.400 15.600 ;
        RECT 273.400 15.000 274.200 15.800 ;
        RECT 274.800 15.600 275.600 16.400 ;
        RECT 276.400 15.600 277.200 16.400 ;
        RECT 265.200 13.600 266.000 14.400 ;
        RECT 266.800 14.200 267.400 15.000 ;
        RECT 268.200 14.800 269.000 15.000 ;
        RECT 271.600 14.800 272.400 15.000 ;
        RECT 266.800 13.600 271.600 14.200 ;
        RECT 252.400 9.700 257.900 10.300 ;
        RECT 252.400 9.600 253.200 9.700 ;
        RECT 263.600 9.600 264.400 10.400 ;
        RECT 266.800 10.200 267.400 13.600 ;
        RECT 270.800 13.400 271.600 13.600 ;
        RECT 273.600 10.200 274.200 15.000 ;
        RECT 274.900 14.400 275.500 15.600 ;
        RECT 276.500 14.400 277.100 15.600 ;
        RECT 284.400 15.000 285.200 15.800 ;
        RECT 290.600 15.600 291.400 15.800 ;
        RECT 297.200 15.600 298.000 16.400 ;
        RECT 285.800 15.000 291.400 15.600 ;
        RECT 274.800 13.600 275.600 14.400 ;
        RECT 276.400 13.600 277.200 14.400 ;
        RECT 282.800 13.600 283.600 14.400 ;
        RECT 284.400 14.200 285.000 15.000 ;
        RECT 285.800 14.800 286.600 15.000 ;
        RECT 289.200 14.800 290.000 15.000 ;
        RECT 284.400 13.600 290.000 14.200 ;
        RECT 278.000 11.600 278.800 12.400 ;
        RECT 281.200 12.300 282.000 12.400 ;
        RECT 282.900 12.300 283.500 13.600 ;
        RECT 281.200 11.700 283.500 12.300 ;
        RECT 281.200 11.600 282.000 11.700 ;
        RECT 278.100 10.400 278.700 11.600 ;
        RECT 281.300 10.400 281.900 11.600 ;
        RECT 252.500 8.400 253.100 9.600 ;
        RECT 266.800 9.400 267.600 10.200 ;
        RECT 273.400 9.400 274.200 10.200 ;
        RECT 278.000 9.600 278.800 10.400 ;
        RECT 281.200 9.600 282.000 10.400 ;
        RECT 284.400 10.200 285.000 13.600 ;
        RECT 289.400 12.200 290.000 13.600 ;
        RECT 289.400 11.400 290.200 12.200 ;
        RECT 290.800 10.200 291.400 15.000 ;
        RECT 297.300 14.400 297.900 15.600 ;
        RECT 298.900 14.400 299.500 33.600 ;
        RECT 302.000 31.600 302.800 32.400 ;
        RECT 300.400 29.600 301.200 30.400 ;
        RECT 300.500 24.400 301.100 29.600 ;
        RECT 302.100 28.400 302.700 31.600 ;
        RECT 302.000 27.600 302.800 28.400 ;
        RECT 303.700 26.400 304.300 37.600 ;
        RECT 308.500 30.400 309.100 47.600 ;
        RECT 311.700 30.400 312.300 55.600 ;
        RECT 314.800 53.600 315.600 54.400 ;
        RECT 318.000 53.600 318.800 54.400 ;
        RECT 322.800 53.600 323.600 54.400 ;
        RECT 326.000 53.600 326.800 54.400 ;
        RECT 313.200 51.600 314.000 52.400 ;
        RECT 313.300 46.400 313.900 51.600 ;
        RECT 313.200 45.600 314.000 46.400 ;
        RECT 318.100 42.400 318.700 53.600 ;
        RECT 319.600 51.600 320.400 52.400 ;
        RECT 321.200 51.600 322.000 52.400 ;
        RECT 319.700 50.300 320.300 51.600 ;
        RECT 319.700 49.700 321.900 50.300 ;
        RECT 318.000 41.600 318.800 42.400 ;
        RECT 316.400 39.600 317.200 40.400 ;
        RECT 318.000 39.600 318.800 40.400 ;
        RECT 313.200 33.600 314.000 34.400 ;
        RECT 313.300 32.400 313.900 33.600 ;
        RECT 313.200 31.600 314.000 32.400 ;
        RECT 308.400 29.600 309.200 30.400 ;
        RECT 310.000 30.300 310.800 30.400 ;
        RECT 311.600 30.300 312.400 30.400 ;
        RECT 310.000 29.700 312.400 30.300 ;
        RECT 316.500 30.300 317.100 39.600 ;
        RECT 318.100 38.400 318.700 39.600 ;
        RECT 321.300 38.400 321.900 49.700 ;
        RECT 326.100 38.400 326.700 53.600 ;
        RECT 329.300 52.400 329.900 69.600 ;
        RECT 334.000 68.400 334.600 71.800 ;
        RECT 338.000 68.400 338.800 68.600 ;
        RECT 332.400 67.600 333.200 68.400 ;
        RECT 334.000 67.800 338.800 68.400 ;
        RECT 332.500 56.400 333.100 67.600 ;
        RECT 334.000 67.000 334.600 67.800 ;
        RECT 335.400 67.000 336.200 67.200 ;
        RECT 338.800 67.000 339.600 67.200 ;
        RECT 340.800 67.000 341.400 71.800 ;
        RECT 342.000 67.600 342.800 68.400 ;
        RECT 334.000 66.200 334.800 67.000 ;
        RECT 335.400 66.400 339.600 67.000 ;
        RECT 340.600 66.200 341.400 67.000 ;
        RECT 334.000 63.600 334.800 64.400 ;
        RECT 338.800 63.600 339.600 64.400 ;
        RECT 332.400 55.600 333.200 56.400 ;
        RECT 334.100 52.400 334.700 63.600 ;
        RECT 338.900 56.400 339.500 63.600 ;
        RECT 342.100 60.400 342.700 67.600 ;
        RECT 343.600 66.200 344.400 71.800 ;
        RECT 345.300 68.400 345.900 87.600 ;
        RECT 361.200 77.600 362.000 78.400 ;
        RECT 345.200 67.600 346.000 68.400 ;
        RECT 346.800 64.200 347.600 75.800 ;
        RECT 348.400 69.400 349.200 70.200 ;
        RECT 348.500 62.400 349.100 69.400 ;
        RECT 353.200 67.600 354.000 68.400 ;
        RECT 348.400 61.600 349.200 62.400 ;
        RECT 342.000 59.600 342.800 60.400 ;
        RECT 338.800 55.600 339.600 56.400 ;
        RECT 348.400 55.600 349.200 56.400 ;
        RECT 338.800 53.600 339.600 54.400 ;
        RECT 340.400 53.600 341.200 54.400 ;
        RECT 338.900 52.400 339.500 53.600 ;
        RECT 340.500 52.400 341.100 53.600 ;
        RECT 348.500 52.400 349.100 55.600 ;
        RECT 350.000 53.600 350.800 54.400 ;
        RECT 327.600 51.600 328.400 52.400 ;
        RECT 329.200 51.600 330.000 52.400 ;
        RECT 330.800 51.600 331.600 52.400 ;
        RECT 332.400 51.600 333.200 52.400 ;
        RECT 334.000 51.600 334.800 52.400 ;
        RECT 338.800 51.600 339.600 52.400 ;
        RECT 340.400 51.600 341.200 52.400 ;
        RECT 346.800 51.600 347.600 52.400 ;
        RECT 348.400 51.600 349.200 52.400 ;
        RECT 327.700 48.400 328.300 51.600 ;
        RECT 327.600 47.600 328.400 48.400 ;
        RECT 329.300 40.400 329.900 51.600 ;
        RECT 329.200 39.600 330.000 40.400 ;
        RECT 318.000 37.600 318.800 38.400 ;
        RECT 321.200 37.600 322.000 38.400 ;
        RECT 326.000 37.600 326.800 38.400 ;
        RECT 330.900 34.400 331.500 51.600 ;
        RECT 350.100 50.400 350.700 53.600 ;
        RECT 337.200 49.600 338.000 50.400 ;
        RECT 343.600 49.600 344.400 50.400 ;
        RECT 350.000 49.600 350.800 50.400 ;
        RECT 351.600 50.200 352.400 55.800 ;
        RECT 353.300 54.400 353.900 67.600 ;
        RECT 356.400 64.200 357.200 75.800 ;
        RECT 362.800 66.200 363.600 71.800 ;
        RECT 364.400 67.600 365.200 68.400 ;
        RECT 366.000 64.200 366.800 75.800 ;
        RECT 367.600 71.600 368.400 72.400 ;
        RECT 367.700 70.200 368.300 71.600 ;
        RECT 367.600 69.400 368.400 70.200 ;
        RECT 372.400 67.600 373.200 68.400 ;
        RECT 353.200 53.600 354.000 54.400 ;
        RECT 337.300 48.400 337.900 49.600 ;
        RECT 337.200 47.600 338.000 48.400 ;
        RECT 348.400 47.600 349.200 48.400 ;
        RECT 330.800 33.600 331.600 34.400 ;
        RECT 322.800 31.600 323.600 32.400 ;
        RECT 318.000 30.300 318.800 30.400 ;
        RECT 316.500 29.700 318.800 30.300 ;
        RECT 310.000 29.600 310.800 29.700 ;
        RECT 311.600 29.600 312.400 29.700 ;
        RECT 318.000 29.600 318.800 29.700 ;
        RECT 308.400 27.600 309.200 28.400 ;
        RECT 303.600 25.600 304.400 26.400 ;
        RECT 300.400 23.600 301.200 24.400 ;
        RECT 305.200 23.600 306.000 24.400 ;
        RECT 300.500 16.400 301.100 23.600 ;
        RECT 310.100 20.400 310.700 29.600 ;
        RECT 314.800 27.600 315.600 28.400 ;
        RECT 319.600 27.600 320.400 28.400 ;
        RECT 302.000 19.600 302.800 20.400 ;
        RECT 310.000 19.600 310.800 20.400 ;
        RECT 300.400 15.600 301.200 16.400 ;
        RECT 297.200 13.600 298.000 14.400 ;
        RECT 298.800 13.600 299.600 14.400 ;
        RECT 302.100 10.400 302.700 19.600 ;
        RECT 314.900 18.400 315.500 27.600 ;
        RECT 322.900 26.400 323.500 31.600 ;
        RECT 330.900 30.400 331.500 33.600 ;
        RECT 332.400 31.600 333.200 32.400 ;
        RECT 334.000 31.600 334.800 32.400 ;
        RECT 327.600 29.600 328.400 30.400 ;
        RECT 329.200 29.600 330.000 30.400 ;
        RECT 330.800 29.600 331.600 30.400 ;
        RECT 324.400 27.600 325.200 28.400 ;
        RECT 324.500 26.400 325.100 27.600 ;
        RECT 327.700 26.400 328.300 29.600 ;
        RECT 316.400 25.600 317.200 26.400 ;
        RECT 322.800 25.600 323.600 26.400 ;
        RECT 324.400 25.600 325.200 26.400 ;
        RECT 327.600 25.600 328.400 26.400 ;
        RECT 310.000 17.600 310.800 18.400 ;
        RECT 314.800 17.600 315.600 18.400 ;
        RECT 310.100 16.400 310.700 17.600 ;
        RECT 316.500 16.400 317.100 25.600 ;
        RECT 324.400 19.600 325.200 20.400 ;
        RECT 306.800 15.600 307.600 16.400 ;
        RECT 308.400 15.600 309.200 16.400 ;
        RECT 310.000 15.600 310.800 16.400 ;
        RECT 316.400 15.600 317.200 16.400 ;
        RECT 322.800 15.600 323.600 16.400 ;
        RECT 306.900 12.400 307.500 15.600 ;
        RECT 308.500 14.400 309.100 15.600 ;
        RECT 316.500 14.400 317.100 15.600 ;
        RECT 308.400 13.600 309.200 14.400 ;
        RECT 316.400 13.600 317.200 14.400 ;
        RECT 324.500 12.400 325.100 19.600 ;
        RECT 332.500 18.400 333.100 31.600 ;
        RECT 334.100 30.400 334.700 31.600 ;
        RECT 348.500 30.400 349.100 47.600 ;
        RECT 350.100 38.400 350.700 49.600 ;
        RECT 354.800 46.200 355.600 57.800 ;
        RECT 356.400 51.600 357.200 52.600 ;
        RECT 364.400 46.200 365.200 57.800 ;
        RECT 369.200 57.600 370.000 58.400 ;
        RECT 369.300 56.400 369.900 57.600 ;
        RECT 369.200 55.600 370.000 56.400 ;
        RECT 370.800 50.200 371.600 55.800 ;
        RECT 372.500 54.400 373.100 67.600 ;
        RECT 375.600 64.200 376.400 75.800 ;
        RECT 380.500 68.400 381.100 109.600 ;
        RECT 382.000 105.600 382.800 106.400 ;
        RECT 382.000 103.600 382.800 104.400 ;
        RECT 382.100 100.400 382.700 103.600 ;
        RECT 382.000 99.600 382.800 100.400 ;
        RECT 382.100 92.400 382.700 99.600 ;
        RECT 385.300 96.400 385.900 131.600 ;
        RECT 386.900 110.400 387.500 135.600 ;
        RECT 388.500 134.400 389.100 135.600 ;
        RECT 388.400 133.600 389.200 134.400 ;
        RECT 390.000 133.600 390.800 134.400 ;
        RECT 391.700 126.300 392.300 149.600 ;
        RECT 402.900 148.400 403.500 159.600 ;
        RECT 404.500 154.400 405.100 163.600 ;
        RECT 404.400 153.600 405.200 154.400 ;
        RECT 406.100 150.400 406.700 167.600 ;
        RECT 409.300 150.400 409.900 175.600 ;
        RECT 410.900 174.400 411.500 207.600 ;
        RECT 414.000 184.200 414.800 195.800 ;
        RECT 414.000 179.600 414.800 180.400 ;
        RECT 410.800 173.600 411.600 174.400 ;
        RECT 410.900 172.400 411.500 173.600 ;
        RECT 410.800 171.600 411.600 172.400 ;
        RECT 412.400 171.600 413.200 172.400 ;
        RECT 412.500 170.300 413.100 171.600 ;
        RECT 410.900 169.700 413.100 170.300 ;
        RECT 404.400 149.600 405.200 150.400 ;
        RECT 406.000 150.300 406.800 150.400 ;
        RECT 406.000 149.700 408.300 150.300 ;
        RECT 406.000 149.600 406.800 149.700 ;
        RECT 393.200 147.600 394.000 148.400 ;
        RECT 402.800 147.600 403.600 148.400 ;
        RECT 404.500 148.300 405.100 149.600 ;
        RECT 404.500 147.700 406.700 148.300 ;
        RECT 393.300 138.400 393.900 147.600 ;
        RECT 394.800 145.600 395.600 146.400 ;
        RECT 399.600 143.600 400.400 144.400 ;
        RECT 401.200 143.600 402.000 144.400 ;
        RECT 393.200 137.600 394.000 138.400 ;
        RECT 399.700 136.400 400.300 143.600 ;
        RECT 401.300 138.400 401.900 143.600 ;
        RECT 401.200 137.600 402.000 138.400 ;
        RECT 404.400 137.600 405.200 138.400 ;
        RECT 398.000 135.600 398.800 136.400 ;
        RECT 399.600 135.600 400.400 136.400 ;
        RECT 398.100 134.400 398.700 135.600 ;
        RECT 404.500 134.400 405.100 137.600 ;
        RECT 398.000 133.600 398.800 134.400 ;
        RECT 404.400 133.600 405.200 134.400 ;
        RECT 406.100 132.400 406.700 147.700 ;
        RECT 407.700 132.400 408.300 149.700 ;
        RECT 409.200 149.600 410.000 150.400 ;
        RECT 410.900 148.400 411.500 169.700 ;
        RECT 414.100 150.400 414.700 179.600 ;
        RECT 415.700 178.400 416.300 211.600 ;
        RECT 417.200 206.200 418.000 217.800 ;
        RECT 418.800 211.800 419.600 212.600 ;
        RECT 418.900 210.400 419.500 211.800 ;
        RECT 425.200 211.600 426.000 212.400 ;
        RECT 418.800 209.600 419.600 210.400 ;
        RECT 420.400 189.600 421.200 190.400 ;
        RECT 420.500 184.400 421.100 189.600 ;
        RECT 420.400 183.600 421.200 184.400 ;
        RECT 423.600 184.200 424.400 195.800 ;
        RECT 425.300 188.400 425.900 211.600 ;
        RECT 426.800 206.200 427.600 217.800 ;
        RECT 441.200 217.600 442.000 218.400 ;
        RECT 442.900 216.400 443.500 219.600 ;
        RECT 438.000 215.600 438.800 216.400 ;
        RECT 442.800 215.600 443.600 216.400 ;
        RECT 436.400 213.600 437.200 214.400 ;
        RECT 433.200 211.600 434.000 212.400 ;
        RECT 431.600 207.600 432.400 208.400 ;
        RECT 436.500 204.400 437.100 213.600 ;
        RECT 436.400 203.600 437.200 204.400 ;
        RECT 425.200 187.600 426.000 188.400 ;
        RECT 425.300 182.400 425.900 187.600 ;
        RECT 426.800 186.200 427.600 191.800 ;
        RECT 428.400 186.200 429.200 191.800 ;
        RECT 430.000 189.600 430.800 190.400 ;
        RECT 425.200 181.600 426.000 182.400 ;
        RECT 415.600 177.600 416.400 178.400 ;
        RECT 418.800 173.600 419.600 174.400 ;
        RECT 420.400 173.600 421.200 174.400 ;
        RECT 417.200 169.600 418.000 170.400 ;
        RECT 417.300 158.400 417.900 169.600 ;
        RECT 418.900 158.400 419.500 173.600 ;
        RECT 420.500 172.400 421.100 173.600 ;
        RECT 420.400 171.600 421.200 172.400 ;
        RECT 417.200 157.600 418.000 158.400 ;
        RECT 418.800 157.600 419.600 158.400 ;
        RECT 420.500 156.400 421.100 171.600 ;
        RECT 422.000 170.200 422.800 175.800 ;
        RECT 425.200 166.200 426.000 177.800 ;
        RECT 426.800 171.800 427.600 172.600 ;
        RECT 420.400 155.600 421.200 156.400 ;
        RECT 415.600 151.600 416.400 152.400 ;
        RECT 415.700 150.400 416.300 151.600 ;
        RECT 412.400 149.600 413.200 150.400 ;
        RECT 414.000 149.600 414.800 150.400 ;
        RECT 415.600 149.600 416.400 150.400 ;
        RECT 420.400 149.600 421.200 150.400 ;
        RECT 410.800 147.600 411.600 148.400 ;
        RECT 410.800 145.600 411.600 146.400 ;
        RECT 410.800 143.600 411.600 144.400 ;
        RECT 410.900 138.400 411.500 143.600 ;
        RECT 414.100 142.400 414.700 149.600 ;
        RECT 420.500 146.400 421.100 149.600 ;
        RECT 425.200 147.600 426.000 148.400 ;
        RECT 420.400 145.600 421.200 146.400 ;
        RECT 414.000 141.600 414.800 142.400 ;
        RECT 426.900 140.400 427.500 171.800 ;
        RECT 428.400 149.600 429.200 150.400 ;
        RECT 428.400 147.600 429.200 148.400 ;
        RECT 428.400 145.600 429.200 146.400 ;
        RECT 428.500 144.400 429.100 145.600 ;
        RECT 428.400 143.600 429.200 144.400 ;
        RECT 426.800 139.600 427.600 140.400 ;
        RECT 430.100 138.400 430.700 189.600 ;
        RECT 431.600 184.200 432.400 195.800 ;
        RECT 438.100 190.400 438.700 215.600 ;
        RECT 439.600 211.600 440.400 212.400 ;
        RECT 444.500 210.400 445.100 225.600 ;
        RECT 449.300 214.400 449.900 229.600 ;
        RECT 463.600 227.600 464.400 228.400 ;
        RECT 466.800 227.600 467.600 228.400 ;
        RECT 454.000 226.300 454.800 226.400 ;
        RECT 454.000 225.700 456.300 226.300 ;
        RECT 454.000 225.600 454.800 225.700 ;
        RECT 452.400 219.600 453.200 220.400 ;
        RECT 449.200 213.600 450.000 214.400 ;
        RECT 444.400 209.600 445.200 210.400 ;
        RECT 439.600 203.600 440.400 204.400 ;
        RECT 449.300 204.300 449.900 213.600 ;
        RECT 452.500 210.400 453.100 219.600 ;
        RECT 455.700 218.400 456.300 225.700 ;
        RECT 457.200 225.600 458.000 226.400 ;
        RECT 458.800 225.600 459.600 226.400 ;
        RECT 458.900 220.400 459.500 225.600 ;
        RECT 460.400 223.600 461.200 224.400 ;
        RECT 458.800 219.600 459.600 220.400 ;
        RECT 455.600 217.600 456.400 218.400 ;
        RECT 457.200 215.600 458.000 216.400 ;
        RECT 457.200 213.600 458.000 214.400 ;
        RECT 458.800 213.600 459.600 214.400 ;
        RECT 452.400 209.600 453.200 210.400 ;
        RECT 449.300 203.700 451.500 204.300 ;
        RECT 433.200 189.400 434.000 190.400 ;
        RECT 438.000 189.600 438.800 190.400 ;
        RECT 433.200 185.600 434.000 186.400 ;
        RECT 433.300 174.400 433.900 185.600 ;
        RECT 433.200 173.600 434.000 174.400 ;
        RECT 431.600 171.600 432.400 172.400 ;
        RECT 431.700 170.400 432.300 171.600 ;
        RECT 431.600 169.600 432.400 170.400 ;
        RECT 434.800 166.200 435.600 177.800 ;
        RECT 431.600 145.600 432.400 146.400 ;
        RECT 433.200 145.600 434.000 146.400 ;
        RECT 433.300 144.400 433.900 145.600 ;
        RECT 433.200 143.600 434.000 144.400 ;
        RECT 436.400 143.600 437.200 144.400 ;
        RECT 431.600 141.600 432.400 142.400 ;
        RECT 410.800 137.600 411.600 138.400 ;
        RECT 426.800 137.600 427.600 138.400 ;
        RECT 430.000 137.600 430.800 138.400 ;
        RECT 418.800 135.600 419.600 136.400 ;
        RECT 399.600 131.600 400.400 132.400 ;
        RECT 406.000 131.600 406.800 132.400 ;
        RECT 407.600 131.600 408.400 132.400 ;
        RECT 414.000 131.600 414.800 132.400 ;
        RECT 415.600 131.600 416.400 132.400 ;
        RECT 417.200 131.600 418.000 132.400 ;
        RECT 393.200 129.600 394.000 130.400 ;
        RECT 393.300 128.400 393.900 129.600 ;
        RECT 393.200 127.600 394.000 128.400 ;
        RECT 396.400 127.600 397.200 128.400 ;
        RECT 391.700 125.700 393.900 126.300 ;
        RECT 388.400 113.600 389.200 114.400 ;
        RECT 386.800 109.600 387.600 110.400 ;
        RECT 388.500 108.400 389.100 113.600 ;
        RECT 393.300 112.400 393.900 125.700 ;
        RECT 394.800 113.600 395.600 114.400 ;
        RECT 394.900 112.400 395.500 113.600 ;
        RECT 390.000 111.600 390.800 112.400 ;
        RECT 393.200 111.600 394.000 112.400 ;
        RECT 394.800 111.600 395.600 112.400 ;
        RECT 386.800 107.600 387.600 108.400 ;
        RECT 388.400 107.600 389.200 108.400 ;
        RECT 393.300 98.400 393.900 111.600 ;
        RECT 396.500 108.400 397.100 127.600 ;
        RECT 406.100 120.400 406.700 131.600 ;
        RECT 407.700 128.400 408.300 131.600 ;
        RECT 407.600 127.600 408.400 128.400 ;
        RECT 399.600 119.600 400.400 120.400 ;
        RECT 406.000 119.600 406.800 120.400 ;
        RECT 396.400 107.600 397.200 108.400 ;
        RECT 398.000 107.600 398.800 108.400 ;
        RECT 394.800 103.600 395.600 104.400 ;
        RECT 394.900 98.400 395.500 103.600 ;
        RECT 398.100 102.400 398.700 107.600 ;
        RECT 399.700 106.400 400.300 119.600 ;
        RECT 414.100 116.400 414.700 131.600 ;
        RECT 415.700 130.400 416.300 131.600 ;
        RECT 415.600 129.600 416.400 130.400 ;
        RECT 417.300 118.400 417.900 131.600 ;
        RECT 418.900 126.400 419.500 135.600 ;
        RECT 422.000 135.000 422.800 135.800 ;
        RECT 423.400 135.000 427.600 135.600 ;
        RECT 428.600 135.000 429.400 135.800 ;
        RECT 420.400 133.600 421.200 134.400 ;
        RECT 422.000 134.200 422.600 135.000 ;
        RECT 423.400 134.800 424.200 135.000 ;
        RECT 426.800 134.800 427.600 135.000 ;
        RECT 422.000 133.600 426.800 134.200 ;
        RECT 422.000 130.200 422.600 133.600 ;
        RECT 426.000 133.400 426.800 133.600 ;
        RECT 428.800 130.200 429.400 135.000 ;
        RECT 430.000 133.600 430.800 134.400 ;
        RECT 430.100 132.400 430.700 133.600 ;
        RECT 430.000 131.600 430.800 132.400 ;
        RECT 431.700 130.400 432.300 141.600 ;
        RECT 433.300 134.400 433.900 143.600 ;
        RECT 433.200 133.600 434.000 134.400 ;
        RECT 434.800 131.600 435.600 132.400 ;
        RECT 422.000 129.400 422.800 130.200 ;
        RECT 428.600 129.400 429.400 130.200 ;
        RECT 431.600 129.600 432.400 130.400 ;
        RECT 418.800 126.300 419.600 126.400 ;
        RECT 418.800 125.700 421.100 126.300 ;
        RECT 418.800 125.600 419.600 125.700 ;
        RECT 417.200 117.600 418.000 118.400 ;
        RECT 414.000 115.600 414.800 116.400 ;
        RECT 417.200 115.600 418.000 116.400 ;
        RECT 406.000 113.600 406.800 114.400 ;
        RECT 406.100 110.400 406.700 113.600 ;
        RECT 407.600 111.600 408.400 112.400 ;
        RECT 412.400 111.600 413.200 112.400 ;
        RECT 414.000 111.600 414.800 112.400 ;
        RECT 406.000 109.600 406.800 110.400 ;
        RECT 399.600 105.600 400.400 106.400 ;
        RECT 406.000 105.600 406.800 106.400 ;
        RECT 396.400 101.600 397.200 102.400 ;
        RECT 398.000 101.600 398.800 102.400 ;
        RECT 388.400 97.600 389.200 98.400 ;
        RECT 393.200 97.600 394.000 98.400 ;
        RECT 394.800 97.600 395.600 98.400 ;
        RECT 385.200 95.600 386.000 96.400 ;
        RECT 383.600 93.600 384.400 94.400 ;
        RECT 382.000 91.600 382.800 92.400 ;
        RECT 382.000 89.600 382.800 90.400 ;
        RECT 382.100 88.400 382.700 89.600 ;
        RECT 382.000 87.600 382.800 88.400 ;
        RECT 383.700 78.400 384.300 93.600 ;
        RECT 385.200 91.600 386.000 92.400 ;
        RECT 385.300 90.400 385.900 91.600 ;
        RECT 388.500 90.400 389.100 97.600 ;
        RECT 390.000 95.600 390.800 96.400 ;
        RECT 394.800 95.600 395.600 96.400 ;
        RECT 390.100 94.400 390.700 95.600 ;
        RECT 390.000 93.600 390.800 94.400 ;
        RECT 391.600 93.600 392.400 94.400 ;
        RECT 391.700 92.400 392.300 93.600 ;
        RECT 390.000 91.600 390.800 92.400 ;
        RECT 391.600 91.600 392.400 92.400 ;
        RECT 385.200 89.600 386.000 90.400 ;
        RECT 388.400 89.600 389.200 90.400 ;
        RECT 394.900 88.400 395.500 95.600 ;
        RECT 396.500 94.400 397.100 101.600 ;
        RECT 396.400 93.600 397.200 94.400 ;
        RECT 398.000 94.300 398.800 94.400 ;
        RECT 399.700 94.300 400.300 105.600 ;
        RECT 401.200 103.600 402.000 104.400 ;
        RECT 398.000 93.700 400.300 94.300 ;
        RECT 398.000 93.600 398.800 93.700 ;
        RECT 398.100 92.400 398.700 93.600 ;
        RECT 398.000 91.600 398.800 92.400 ;
        RECT 401.300 88.400 401.900 103.600 ;
        RECT 406.100 102.400 406.700 105.600 ;
        RECT 406.000 101.600 406.800 102.400 ;
        RECT 407.700 98.400 408.300 111.600 ;
        RECT 412.400 109.600 413.200 110.400 ;
        RECT 414.100 108.400 414.700 111.600 ;
        RECT 417.300 110.400 417.900 115.600 ;
        RECT 417.200 109.600 418.000 110.400 ;
        RECT 420.500 108.400 421.100 125.700 ;
        RECT 431.700 118.400 432.300 129.600 ;
        RECT 434.900 128.400 435.500 131.600 ;
        RECT 436.500 128.400 437.100 143.600 ;
        RECT 438.100 140.400 438.700 189.600 ;
        RECT 439.700 178.400 440.300 203.600 ;
        RECT 450.900 198.400 451.500 203.700 ;
        RECT 450.800 197.600 451.600 198.400 ;
        RECT 441.200 184.200 442.000 195.800 ;
        RECT 452.500 192.400 453.100 209.600 ;
        RECT 452.400 191.600 453.200 192.400 ;
        RECT 452.400 189.600 453.200 190.400 ;
        RECT 454.000 189.600 454.800 190.400 ;
        RECT 452.500 188.400 453.100 189.600 ;
        RECT 454.100 188.400 454.700 189.600 ;
        RECT 452.400 187.600 453.200 188.400 ;
        RECT 454.000 187.600 454.800 188.400 ;
        RECT 457.300 186.400 457.900 213.600 ;
        RECT 458.900 212.400 459.500 213.600 ;
        RECT 460.500 212.400 461.100 223.600 ;
        RECT 465.200 215.600 466.000 216.400 ;
        RECT 465.200 213.600 466.000 214.400 ;
        RECT 458.800 211.600 459.600 212.400 ;
        RECT 460.400 211.600 461.200 212.400 ;
        RECT 463.600 209.600 464.400 210.400 ;
        RECT 465.200 209.600 466.000 210.400 ;
        RECT 462.000 199.600 462.800 200.400 ;
        RECT 462.100 190.400 462.700 199.600 ;
        RECT 462.000 189.600 462.800 190.400 ;
        RECT 463.700 188.400 464.300 209.600 ;
        RECT 465.300 204.400 465.900 209.600 ;
        RECT 466.900 208.400 467.500 227.600 ;
        RECT 468.500 214.400 469.100 245.600 ;
        RECT 470.000 231.600 470.800 232.400 ;
        RECT 470.100 230.400 470.700 231.600 ;
        RECT 470.000 229.600 470.800 230.400 ;
        RECT 470.000 223.600 470.800 224.400 ;
        RECT 470.100 220.400 470.700 223.600 ;
        RECT 470.000 219.600 470.800 220.400 ;
        RECT 468.400 213.600 469.200 214.400 ;
        RECT 466.800 207.600 467.600 208.400 ;
        RECT 466.900 206.400 467.500 207.600 ;
        RECT 466.800 205.600 467.600 206.400 ;
        RECT 465.200 203.600 466.000 204.400 ;
        RECT 468.500 200.400 469.100 213.600 ;
        RECT 470.000 211.600 470.800 212.400 ;
        RECT 470.100 204.400 470.700 211.600 ;
        RECT 470.000 203.600 470.800 204.400 ;
        RECT 468.400 199.600 469.200 200.400 ;
        RECT 471.700 198.400 472.300 249.700 ;
        RECT 474.900 242.400 475.500 251.600 ;
        RECT 478.000 250.300 478.800 250.400 ;
        RECT 479.700 250.300 480.300 273.600 ;
        RECT 482.900 272.400 483.500 273.600 ;
        RECT 482.800 271.600 483.600 272.400 ;
        RECT 484.400 266.200 485.200 271.800 ;
        RECT 487.600 264.200 488.400 275.800 ;
        RECT 489.200 271.600 490.000 272.400 ;
        RECT 489.300 270.200 489.900 271.600 ;
        RECT 489.200 269.400 490.000 270.200 ;
        RECT 487.600 261.600 488.400 262.400 ;
        RECT 481.200 259.600 482.000 260.400 ;
        RECT 481.300 254.400 481.900 259.600 ;
        RECT 487.700 254.400 488.300 261.600 ;
        RECT 490.900 258.400 491.500 291.600 ;
        RECT 492.800 290.200 493.400 295.000 ;
        RECT 494.000 293.600 494.800 294.400 ;
        RECT 508.400 293.600 509.200 294.400 ;
        RECT 494.100 292.400 494.700 293.600 ;
        RECT 494.000 291.600 494.800 292.400 ;
        RECT 510.000 290.200 510.800 295.800 ;
        RECT 511.600 293.600 512.400 294.400 ;
        RECT 492.600 289.400 493.400 290.200 ;
        RECT 495.600 269.600 496.400 270.400 ;
        RECT 492.400 267.600 493.200 268.400 ;
        RECT 490.800 257.600 491.600 258.400 ;
        RECT 481.200 253.600 482.000 254.400 ;
        RECT 487.600 253.600 488.400 254.400 ;
        RECT 486.000 251.600 486.800 252.400 ;
        RECT 478.000 249.700 480.300 250.300 ;
        RECT 478.000 249.600 478.800 249.700 ;
        RECT 482.800 249.600 483.600 250.400 ;
        RECT 486.000 249.600 486.800 250.400 ;
        RECT 489.200 249.600 490.000 250.400 ;
        RECT 482.900 244.400 483.500 249.600 ;
        RECT 482.800 243.600 483.600 244.400 ;
        RECT 474.800 241.600 475.600 242.400 ;
        RECT 476.400 233.600 477.200 234.400 ;
        RECT 486.000 233.600 486.800 234.400 ;
        RECT 473.200 229.600 474.000 230.400 ;
        RECT 473.300 224.400 473.900 229.600 ;
        RECT 474.800 227.600 475.600 228.400 ;
        RECT 473.200 223.600 474.000 224.400 ;
        RECT 474.900 222.400 475.500 227.600 ;
        RECT 476.500 226.400 477.100 233.600 ;
        RECT 481.200 231.800 482.000 232.600 ;
        RECT 486.100 232.400 486.700 233.600 ;
        RECT 481.200 228.400 481.800 231.800 ;
        RECT 486.000 231.600 486.800 232.400 ;
        RECT 487.800 231.800 488.600 232.600 ;
        RECT 485.200 228.400 486.000 228.600 ;
        RECT 479.600 227.600 480.400 228.400 ;
        RECT 481.200 227.800 486.000 228.400 ;
        RECT 479.700 226.400 480.300 227.600 ;
        RECT 481.200 227.000 481.800 227.800 ;
        RECT 482.600 227.000 483.400 227.200 ;
        RECT 486.000 227.000 486.800 227.200 ;
        RECT 488.000 227.000 488.600 231.800 ;
        RECT 489.200 227.600 490.000 228.400 ;
        RECT 476.400 225.600 477.200 226.400 ;
        RECT 479.600 225.600 480.400 226.400 ;
        RECT 481.200 226.200 482.000 227.000 ;
        RECT 482.600 226.400 486.800 227.000 ;
        RECT 487.800 226.200 488.600 227.000 ;
        RECT 489.300 224.400 489.900 227.600 ;
        RECT 490.800 226.200 491.600 231.800 ;
        RECT 492.500 228.400 493.100 267.600 ;
        RECT 497.200 264.200 498.000 275.800 ;
        RECT 503.600 266.200 504.400 271.800 ;
        RECT 502.000 263.600 502.800 264.400 ;
        RECT 506.800 264.200 507.600 275.800 ;
        RECT 511.700 270.400 512.300 293.600 ;
        RECT 513.200 286.200 514.000 297.800 ;
        RECT 516.500 294.400 517.100 305.600 ;
        RECT 518.000 304.200 518.800 315.800 ;
        RECT 521.200 304.200 522.000 315.800 ;
        RECT 522.800 304.200 523.600 317.800 ;
        RECT 524.400 304.200 525.200 317.800 ;
        RECT 529.200 311.600 530.000 312.400 ;
        RECT 535.600 311.600 536.400 312.400 ;
        RECT 529.200 309.600 530.000 310.400 ;
        RECT 537.200 309.600 538.000 310.400 ;
        RECT 543.600 305.600 544.400 306.400 ;
        RECT 545.200 306.200 546.000 311.800 ;
        RECT 546.900 306.400 547.500 331.600 ;
        RECT 559.600 326.200 560.400 337.800 ;
        RECT 561.200 331.600 562.000 332.400 ;
        RECT 566.000 331.600 566.800 332.400 ;
        RECT 554.800 323.600 555.600 324.400 ;
        RECT 546.800 305.600 547.600 306.400 ;
        RECT 532.400 303.600 533.200 304.400 ;
        RECT 548.400 304.200 549.200 315.800 ;
        RECT 550.000 309.400 550.800 310.200 ;
        RECT 550.100 304.400 550.700 309.400 ;
        RECT 551.600 307.600 552.400 308.400 ;
        RECT 550.000 303.600 550.800 304.400 ;
        RECT 516.400 293.600 517.200 294.400 ;
        RECT 514.800 291.800 515.600 292.600 ;
        RECT 514.900 288.400 515.500 291.800 ;
        RECT 514.800 287.600 515.600 288.400 ;
        RECT 522.800 286.200 523.600 297.800 ;
        RECT 524.400 287.600 525.200 288.400 ;
        RECT 527.600 287.600 528.400 288.400 ;
        RECT 510.000 269.600 510.800 270.400 ;
        RECT 511.600 269.600 512.400 270.400 ;
        RECT 502.100 262.400 502.700 263.600 ;
        RECT 502.000 261.600 502.800 262.400 ;
        RECT 494.000 259.600 494.800 260.400 ;
        RECT 494.100 256.400 494.700 259.600 ;
        RECT 510.100 258.400 510.700 269.600 ;
        RECT 511.700 268.400 512.300 269.600 ;
        RECT 511.600 267.600 512.400 268.400 ;
        RECT 516.400 264.200 517.200 275.800 ;
        RECT 521.200 273.600 522.000 274.400 ;
        RECT 521.300 272.400 521.900 273.600 ;
        RECT 521.200 271.600 522.000 272.400 ;
        RECT 521.200 269.600 522.000 270.400 ;
        RECT 521.300 258.400 521.900 269.600 ;
        RECT 522.800 266.200 523.600 271.800 ;
        RECT 524.500 268.400 525.100 287.600 ;
        RECT 529.200 283.600 530.000 284.400 ;
        RECT 524.400 267.600 525.200 268.400 ;
        RECT 526.000 264.200 526.800 275.800 ;
        RECT 527.600 271.600 528.400 272.400 ;
        RECT 527.700 270.200 528.300 271.600 ;
        RECT 527.600 269.400 528.400 270.200 ;
        RECT 529.300 258.400 529.900 283.600 ;
        RECT 532.500 258.400 533.100 303.600 ;
        RECT 545.200 284.200 546.000 297.800 ;
        RECT 546.800 284.200 547.600 297.800 ;
        RECT 548.400 284.200 549.200 297.800 ;
        RECT 550.000 286.200 550.800 297.800 ;
        RECT 551.700 296.400 552.300 307.600 ;
        RECT 558.000 304.200 558.800 315.800 ;
        RECT 551.600 295.600 552.400 296.400 ;
        RECT 534.000 267.600 534.800 268.400 ;
        RECT 535.600 264.200 536.400 275.800 ;
        RECT 542.000 266.200 542.800 271.800 ;
        RECT 543.600 267.600 544.400 268.400 ;
        RECT 540.400 263.600 541.200 264.400 ;
        RECT 510.000 257.600 510.800 258.400 ;
        RECT 521.200 257.600 522.000 258.400 ;
        RECT 529.200 257.600 530.000 258.400 ;
        RECT 532.400 257.600 533.200 258.400 ;
        RECT 494.000 255.600 494.800 256.400 ;
        RECT 498.800 255.600 499.600 256.400 ;
        RECT 502.000 255.600 502.800 256.400 ;
        RECT 505.200 255.000 506.000 255.800 ;
        RECT 511.400 255.600 512.200 255.800 ;
        RECT 506.600 255.000 512.200 255.600 ;
        RECT 502.000 253.600 502.800 254.400 ;
        RECT 505.200 254.200 505.800 255.000 ;
        RECT 506.600 254.800 507.400 255.000 ;
        RECT 510.000 254.800 510.800 255.000 ;
        RECT 505.200 253.600 510.800 254.200 ;
        RECT 497.200 251.600 498.000 252.400 ;
        RECT 498.800 251.600 499.600 252.400 ;
        RECT 502.000 251.600 502.800 252.400 ;
        RECT 492.400 227.600 493.200 228.400 ;
        RECT 478.000 223.600 478.800 224.400 ;
        RECT 486.000 223.600 486.800 224.400 ;
        RECT 489.200 223.600 490.000 224.400 ;
        RECT 494.000 224.200 494.800 235.800 ;
        RECT 495.600 231.600 496.400 232.400 ;
        RECT 495.700 230.200 496.300 231.600 ;
        RECT 497.300 230.400 497.900 251.600 ;
        RECT 498.900 234.400 499.500 251.600 ;
        RECT 498.800 233.600 499.600 234.400 ;
        RECT 495.600 229.400 496.400 230.200 ;
        RECT 497.200 229.600 498.000 230.400 ;
        RECT 502.100 226.400 502.700 251.600 ;
        RECT 505.200 250.200 505.800 253.600 ;
        RECT 510.200 252.200 510.800 253.600 ;
        RECT 510.200 251.400 511.000 252.200 ;
        RECT 511.600 250.200 512.200 255.000 ;
        RECT 516.600 255.600 517.400 255.800 ;
        RECT 516.600 255.000 522.200 255.600 ;
        RECT 522.800 255.000 523.600 255.800 ;
        RECT 513.200 253.600 514.000 254.400 ;
        RECT 514.800 253.600 515.600 254.400 ;
        RECT 514.900 252.400 515.500 253.600 ;
        RECT 514.800 251.600 515.600 252.400 ;
        RECT 505.200 249.400 506.000 250.200 ;
        RECT 511.400 249.400 512.200 250.200 ;
        RECT 516.600 250.200 517.200 255.000 ;
        RECT 518.000 254.800 518.800 255.000 ;
        RECT 521.400 254.800 522.200 255.000 ;
        RECT 523.000 254.200 523.600 255.000 ;
        RECT 527.600 255.000 528.400 255.800 ;
        RECT 529.000 255.000 533.200 255.600 ;
        RECT 534.200 255.000 535.000 255.800 ;
        RECT 518.000 253.600 523.600 254.200 ;
        RECT 524.400 253.600 525.200 254.400 ;
        RECT 527.600 254.200 528.200 255.000 ;
        RECT 529.000 254.800 529.800 255.000 ;
        RECT 532.400 254.800 533.200 255.000 ;
        RECT 527.600 253.600 532.400 254.200 ;
        RECT 518.000 252.200 518.600 253.600 ;
        RECT 517.800 251.400 518.600 252.200 ;
        RECT 523.000 250.200 523.600 253.600 ;
        RECT 516.600 249.400 517.400 250.200 ;
        RECT 522.800 249.400 523.600 250.200 ;
        RECT 495.600 225.600 496.400 226.400 ;
        RECT 502.000 225.600 502.800 226.400 ;
        RECT 474.800 221.600 475.600 222.400 ;
        RECT 476.400 215.600 477.200 216.400 ;
        RECT 476.500 214.400 477.100 215.600 ;
        RECT 476.400 213.600 477.200 214.400 ;
        RECT 478.100 212.400 478.700 223.600 ;
        RECT 486.100 218.400 486.700 223.600 ;
        RECT 494.000 219.600 494.800 220.400 ;
        RECT 486.000 217.600 486.800 218.400 ;
        RECT 487.600 215.600 488.400 216.400 ;
        RECT 490.800 215.600 491.600 216.400 ;
        RECT 490.900 214.400 491.500 215.600 ;
        RECT 482.800 213.600 483.600 214.400 ;
        RECT 489.200 213.600 490.000 214.400 ;
        RECT 490.800 213.600 491.600 214.400 ;
        RECT 474.800 211.600 475.600 212.400 ;
        RECT 476.400 211.600 477.200 212.400 ;
        RECT 478.000 211.600 478.800 212.400 ;
        RECT 482.800 211.600 483.600 212.400 ;
        RECT 492.400 211.600 493.200 212.400 ;
        RECT 474.900 210.400 475.500 211.600 ;
        RECT 482.900 210.400 483.500 211.600 ;
        RECT 474.800 209.600 475.600 210.400 ;
        RECT 481.200 209.600 482.000 210.400 ;
        RECT 482.800 209.600 483.600 210.400 ;
        RECT 486.000 209.600 486.800 210.400 ;
        RECT 474.900 208.400 475.500 209.600 ;
        RECT 474.800 207.600 475.600 208.400 ;
        RECT 479.600 207.600 480.400 208.400 ;
        RECT 474.800 203.600 475.600 204.400 ;
        RECT 471.600 197.600 472.400 198.400 ;
        RECT 466.600 191.800 467.400 192.600 ;
        RECT 473.200 191.800 474.000 192.600 ;
        RECT 460.400 187.600 461.200 188.400 ;
        RECT 463.600 187.600 464.400 188.400 ;
        RECT 465.200 187.600 466.000 188.400 ;
        RECT 460.500 186.400 461.100 187.600 ;
        RECT 465.300 186.400 465.900 187.600 ;
        RECT 466.600 187.000 467.200 191.800 ;
        RECT 469.200 188.400 470.000 188.600 ;
        RECT 473.400 188.400 474.000 191.800 ;
        RECT 474.900 188.400 475.500 203.600 ;
        RECT 478.000 189.600 478.800 190.400 ;
        RECT 469.200 187.800 474.000 188.400 ;
        RECT 468.400 187.000 469.200 187.200 ;
        RECT 471.800 187.000 472.600 187.200 ;
        RECT 473.400 187.000 474.000 187.800 ;
        RECT 474.800 187.600 475.600 188.400 ;
        RECT 476.400 187.600 477.200 188.400 ;
        RECT 457.200 185.600 458.000 186.400 ;
        RECT 460.400 185.600 461.200 186.400 ;
        RECT 465.200 185.600 466.000 186.400 ;
        RECT 466.600 186.200 467.400 187.000 ;
        RECT 468.400 186.400 472.600 187.000 ;
        RECT 473.200 186.200 474.000 187.000 ;
        RECT 476.500 186.400 477.100 187.600 ;
        RECT 476.400 185.600 477.200 186.400 ;
        RECT 457.300 180.400 457.900 185.600 ;
        RECT 474.800 183.600 475.600 184.400 ;
        RECT 478.100 184.300 478.700 189.600 ;
        RECT 476.500 183.700 478.700 184.300 ;
        RECT 458.800 181.600 459.600 182.400 ;
        RECT 457.200 179.600 458.000 180.400 ;
        RECT 439.600 177.600 440.400 178.400 ;
        RECT 447.400 175.000 448.200 175.800 ;
        RECT 449.200 175.000 453.400 175.600 ;
        RECT 454.000 175.000 454.800 175.800 ;
        RECT 446.000 173.600 446.800 174.400 ;
        RECT 447.400 170.200 448.000 175.000 ;
        RECT 449.200 174.800 450.000 175.000 ;
        RECT 452.600 174.800 453.400 175.000 ;
        RECT 454.200 174.200 454.800 175.000 ;
        RECT 450.000 173.600 454.800 174.200 ;
        RECT 455.600 173.600 456.400 174.400 ;
        RECT 450.000 173.400 450.800 173.600 ;
        RECT 452.400 171.600 453.200 172.400 ;
        RECT 454.200 170.200 454.800 173.600 ;
        RECT 447.400 169.400 448.200 170.200 ;
        RECT 454.000 169.400 454.800 170.200 ;
        RECT 455.700 158.400 456.300 173.600 ;
        RECT 457.200 170.200 458.000 175.800 ;
        RECT 458.900 174.400 459.500 181.600 ;
        RECT 474.900 178.400 475.500 183.600 ;
        RECT 476.500 180.400 477.100 183.700 ;
        RECT 476.400 179.600 477.200 180.400 ;
        RECT 476.500 178.400 477.100 179.600 ;
        RECT 458.800 173.600 459.600 174.400 ;
        RECT 460.400 166.200 461.200 177.800 ;
        RECT 462.000 171.600 462.800 172.600 ;
        RECT 468.400 171.600 469.200 172.400 ;
        RECT 468.500 164.300 469.100 171.600 ;
        RECT 470.000 166.200 470.800 177.800 ;
        RECT 474.800 177.600 475.600 178.400 ;
        RECT 476.400 177.600 477.200 178.400 ;
        RECT 479.700 174.400 480.300 207.600 ;
        RECT 481.300 206.400 481.900 209.600 ;
        RECT 481.200 205.600 482.000 206.400 ;
        RECT 481.300 200.400 481.900 205.600 ;
        RECT 481.200 199.600 482.000 200.400 ;
        RECT 486.000 199.600 486.800 200.400 ;
        RECT 486.100 188.400 486.700 199.600 ;
        RECT 490.800 192.300 491.600 192.400 ;
        RECT 489.300 191.700 491.600 192.300 ;
        RECT 487.600 189.600 488.400 190.400 ;
        RECT 481.200 187.600 482.000 188.400 ;
        RECT 486.000 187.600 486.800 188.400 ;
        RECT 484.400 185.600 485.200 186.400 ;
        RECT 484.500 184.400 485.100 185.600 ;
        RECT 489.300 184.400 489.900 191.700 ;
        RECT 490.800 191.600 491.600 191.700 ;
        RECT 492.400 189.600 493.200 190.400 ;
        RECT 492.500 188.400 493.100 189.600 ;
        RECT 494.100 188.400 494.700 219.600 ;
        RECT 495.700 218.400 496.300 225.600 ;
        RECT 503.600 224.200 504.400 235.800 ;
        RECT 508.400 233.600 509.200 234.400 ;
        RECT 508.500 232.400 509.100 233.600 ;
        RECT 508.400 231.600 509.200 232.400 ;
        RECT 510.000 226.200 510.800 231.800 ;
        RECT 511.600 227.600 512.400 228.400 ;
        RECT 510.000 223.600 510.800 224.400 ;
        RECT 513.200 224.200 514.000 235.800 ;
        RECT 514.800 231.600 515.600 232.400 ;
        RECT 514.900 230.200 515.500 231.600 ;
        RECT 514.800 229.400 515.600 230.200 ;
        RECT 521.200 229.600 522.000 230.400 ;
        RECT 497.200 221.600 498.000 222.400 ;
        RECT 495.600 217.600 496.400 218.400 ;
        RECT 497.300 214.400 497.900 221.600 ;
        RECT 510.100 218.400 510.700 223.600 ;
        RECT 521.300 218.400 521.900 229.600 ;
        RECT 522.800 224.200 523.600 235.800 ;
        RECT 524.500 224.400 525.100 253.600 ;
        RECT 527.600 250.200 528.200 253.600 ;
        RECT 531.600 253.400 532.400 253.600 ;
        RECT 534.400 250.200 535.000 255.000 ;
        RECT 535.600 253.600 536.400 254.400 ;
        RECT 527.600 249.400 528.400 250.200 ;
        RECT 534.200 249.400 535.000 250.200 ;
        RECT 527.600 234.300 528.400 234.400 ;
        RECT 527.600 233.700 529.900 234.300 ;
        RECT 527.600 233.600 528.400 233.700 ;
        RECT 529.300 230.400 529.900 233.700 ;
        RECT 529.200 229.600 530.000 230.400 ;
        RECT 534.000 226.200 534.800 231.800 ;
        RECT 524.400 223.600 525.200 224.400 ;
        RECT 510.000 217.600 510.800 218.400 ;
        RECT 521.200 217.600 522.000 218.400 ;
        RECT 498.800 215.600 499.600 216.400 ;
        RECT 498.900 214.400 499.500 215.600 ;
        RECT 505.000 215.000 505.800 215.800 ;
        RECT 506.800 215.000 511.000 215.600 ;
        RECT 511.600 215.000 512.400 215.800 ;
        RECT 495.600 213.600 496.400 214.400 ;
        RECT 497.200 213.600 498.000 214.400 ;
        RECT 498.800 213.600 499.600 214.400 ;
        RECT 500.400 213.600 501.200 214.400 ;
        RECT 502.000 213.600 502.800 214.400 ;
        RECT 495.700 212.400 496.300 213.600 ;
        RECT 495.600 211.600 496.400 212.400 ;
        RECT 497.200 211.600 498.000 212.400 ;
        RECT 497.300 198.400 497.900 211.600 ;
        RECT 498.900 200.400 499.500 213.600 ;
        RECT 502.100 210.400 502.700 213.600 ;
        RECT 502.000 209.600 502.800 210.400 ;
        RECT 505.000 210.200 505.600 215.000 ;
        RECT 506.800 214.800 507.600 215.000 ;
        RECT 510.200 214.800 511.000 215.000 ;
        RECT 511.800 214.200 512.400 215.000 ;
        RECT 516.400 215.000 517.200 215.800 ;
        RECT 517.800 215.000 522.000 215.600 ;
        RECT 523.000 215.000 523.800 215.800 ;
        RECT 524.400 215.600 525.200 216.400 ;
        RECT 529.200 215.600 530.000 216.400 ;
        RECT 507.600 213.600 512.400 214.200 ;
        RECT 513.200 213.600 514.000 214.400 ;
        RECT 514.800 213.600 515.600 214.400 ;
        RECT 516.400 214.200 517.000 215.000 ;
        RECT 517.800 214.800 518.600 215.000 ;
        RECT 521.200 214.800 522.000 215.000 ;
        RECT 516.400 213.600 521.200 214.200 ;
        RECT 507.600 213.400 508.400 213.600 ;
        RECT 511.800 210.200 512.400 213.600 ;
        RECT 502.100 208.400 502.700 209.600 ;
        RECT 505.000 209.400 505.800 210.200 ;
        RECT 511.600 209.400 512.400 210.200 ;
        RECT 502.000 207.600 502.800 208.400 ;
        RECT 505.200 207.600 506.000 208.400 ;
        RECT 498.800 199.600 499.600 200.400 ;
        RECT 505.300 198.400 505.900 207.600 ;
        RECT 497.200 197.600 498.000 198.400 ;
        RECT 505.200 197.600 506.000 198.400 ;
        RECT 500.400 191.800 501.200 192.600 ;
        RECT 507.000 191.800 507.800 192.600 ;
        RECT 514.900 192.400 515.500 213.600 ;
        RECT 516.400 210.200 517.000 213.600 ;
        RECT 520.400 213.400 521.200 213.600 ;
        RECT 521.200 211.600 522.000 212.400 ;
        RECT 516.400 209.400 517.200 210.200 ;
        RECT 500.400 188.400 501.000 191.800 ;
        RECT 504.400 188.400 505.200 188.600 ;
        RECT 492.400 187.600 493.200 188.400 ;
        RECT 494.000 187.600 494.800 188.400 ;
        RECT 497.200 187.600 498.000 188.400 ;
        RECT 498.800 187.600 499.600 188.400 ;
        RECT 500.400 187.800 505.200 188.400 ;
        RECT 497.300 186.400 497.900 187.600 ;
        RECT 494.000 185.600 494.800 186.400 ;
        RECT 497.200 185.600 498.000 186.400 ;
        RECT 484.400 183.600 485.200 184.400 ;
        RECT 489.200 183.600 490.000 184.400 ;
        RECT 492.400 183.600 493.200 184.400 ;
        RECT 486.000 181.600 486.800 182.400 ;
        RECT 486.100 178.400 486.700 181.600 ;
        RECT 486.000 177.600 486.800 178.400 ;
        RECT 481.000 175.000 481.800 175.800 ;
        RECT 482.800 175.000 487.000 175.600 ;
        RECT 487.600 175.000 488.400 175.800 ;
        RECT 479.600 173.600 480.400 174.400 ;
        RECT 468.500 163.700 470.700 164.300 ;
        RECT 447.600 157.600 448.400 158.400 ;
        RECT 455.600 157.600 456.400 158.400 ;
        RECT 463.600 155.600 464.400 156.400 ;
        RECT 439.600 153.600 440.400 154.400 ;
        RECT 439.700 150.400 440.300 153.600 ;
        RECT 450.800 151.600 451.600 152.400 ;
        RECT 462.000 151.600 462.800 152.400 ;
        RECT 450.900 150.400 451.500 151.600 ;
        RECT 439.600 149.600 440.400 150.400 ;
        RECT 450.800 149.600 451.600 150.400 ;
        RECT 458.800 149.600 459.600 150.400 ;
        RECT 444.400 147.600 445.200 148.400 ;
        RECT 444.500 146.400 445.100 147.600 ;
        RECT 444.400 145.600 445.200 146.400 ;
        RECT 449.200 145.600 450.000 146.400 ;
        RECT 455.600 145.600 456.400 146.400 ;
        RECT 438.000 139.600 438.800 140.400 ;
        RECT 444.500 138.400 445.100 145.600 ;
        RECT 449.300 138.400 449.900 145.600 ;
        RECT 455.700 142.400 456.300 145.600 ;
        RECT 455.600 141.600 456.400 142.400 ;
        RECT 462.000 141.600 462.800 142.400 ;
        RECT 450.800 139.600 451.600 140.400 ;
        RECT 444.400 137.600 445.200 138.400 ;
        RECT 449.200 137.600 450.000 138.400 ;
        RECT 449.300 136.400 449.900 137.600 ;
        RECT 449.200 135.600 450.000 136.400 ;
        RECT 438.000 133.600 438.800 134.400 ;
        RECT 434.800 127.600 435.600 128.400 ;
        RECT 436.400 127.600 437.200 128.400 ;
        RECT 433.200 119.600 434.000 120.400 ;
        RECT 431.600 117.600 432.400 118.400 ;
        RECT 431.700 116.400 432.300 117.600 ;
        RECT 431.600 115.600 432.400 116.400 ;
        RECT 422.000 111.800 422.800 112.600 ;
        RECT 428.600 111.800 429.400 112.600 ;
        RECT 422.000 108.400 422.600 111.800 ;
        RECT 423.600 109.600 424.400 110.400 ;
        RECT 426.000 108.400 426.800 108.600 ;
        RECT 410.800 107.600 411.600 108.400 ;
        RECT 414.000 107.600 414.800 108.400 ;
        RECT 418.800 107.600 419.600 108.400 ;
        RECT 420.400 107.600 421.200 108.400 ;
        RECT 422.000 107.800 426.800 108.400 ;
        RECT 410.900 98.400 411.500 107.600 ;
        RECT 417.200 103.600 418.000 104.400 ;
        RECT 407.600 97.600 408.400 98.400 ;
        RECT 410.800 97.600 411.600 98.400 ;
        RECT 409.200 95.600 410.000 96.400 ;
        RECT 402.800 93.600 403.600 94.400 ;
        RECT 402.900 90.400 403.500 93.600 ;
        RECT 407.600 91.600 408.400 92.400 ;
        RECT 407.700 90.400 408.300 91.600 ;
        RECT 409.300 90.400 409.900 95.600 ;
        RECT 414.000 93.600 414.800 94.400 ;
        RECT 414.100 90.400 414.700 93.600 ;
        RECT 417.300 92.400 417.900 103.600 ;
        RECT 418.900 94.400 419.500 107.600 ;
        RECT 422.000 107.000 422.600 107.800 ;
        RECT 423.400 107.000 424.200 107.200 ;
        RECT 426.800 107.000 427.600 107.200 ;
        RECT 428.800 107.000 429.400 111.800 ;
        RECT 430.000 107.600 430.800 108.400 ;
        RECT 422.000 106.200 422.800 107.000 ;
        RECT 423.400 106.400 427.600 107.000 ;
        RECT 428.600 106.200 429.400 107.000 ;
        RECT 430.100 106.400 430.700 107.600 ;
        RECT 430.000 105.600 430.800 106.400 ;
        RECT 431.600 106.200 432.400 111.800 ;
        RECT 433.300 108.400 433.900 119.600 ;
        RECT 433.200 107.600 434.000 108.400 ;
        RECT 423.600 97.600 424.400 98.400 ;
        RECT 423.700 94.400 424.300 97.600 ;
        RECT 426.800 95.600 427.600 96.400 ;
        RECT 426.900 94.400 427.500 95.600 ;
        RECT 418.800 93.600 419.600 94.400 ;
        RECT 423.600 93.600 424.400 94.400 ;
        RECT 426.800 93.600 427.600 94.400 ;
        RECT 430.000 93.600 430.800 94.400 ;
        RECT 417.200 91.600 418.000 92.400 ;
        RECT 418.900 90.400 419.500 93.600 ;
        RECT 422.000 91.600 422.800 92.400 ;
        RECT 402.800 89.600 403.600 90.400 ;
        RECT 407.600 89.600 408.400 90.400 ;
        RECT 409.200 89.600 410.000 90.400 ;
        RECT 414.000 89.600 414.800 90.400 ;
        RECT 418.800 89.600 419.600 90.400 ;
        RECT 422.000 89.600 422.800 90.400 ;
        RECT 391.600 87.600 392.400 88.400 ;
        RECT 394.800 87.600 395.600 88.400 ;
        RECT 401.200 87.600 402.000 88.400 ;
        RECT 391.700 78.400 392.300 87.600 ;
        RECT 383.600 77.600 384.400 78.400 ;
        RECT 391.600 77.600 392.400 78.400 ;
        RECT 385.200 71.600 386.000 72.400 ;
        RECT 396.400 71.600 397.200 72.400 ;
        RECT 399.600 71.600 400.400 72.400 ;
        RECT 406.000 71.600 406.800 72.400 ;
        RECT 380.400 67.600 381.200 68.400 ;
        RECT 380.400 63.600 381.200 64.400 ;
        RECT 380.500 60.400 381.100 63.600 ;
        RECT 380.400 59.600 381.200 60.400 ;
        RECT 372.400 53.600 373.200 54.400 ;
        RECT 374.000 46.200 374.800 57.800 ;
        RECT 375.600 57.600 376.400 58.400 ;
        RECT 375.700 52.600 376.300 57.600 ;
        RECT 375.600 51.800 376.400 52.600 ;
        RECT 383.600 46.200 384.400 57.800 ;
        RECT 385.300 56.400 385.900 71.600 ;
        RECT 394.800 69.600 395.600 70.400 ;
        RECT 390.000 67.600 390.800 68.400 ;
        RECT 390.000 59.600 390.800 60.400 ;
        RECT 390.100 56.400 390.700 59.600 ;
        RECT 394.900 58.400 395.500 69.600 ;
        RECT 396.500 68.400 397.100 71.600 ;
        RECT 399.700 70.400 400.300 71.600 ;
        RECT 407.700 70.400 408.300 89.600 ;
        RECT 412.400 87.600 413.200 88.400 ;
        RECT 409.200 81.600 410.000 82.400 ;
        RECT 399.600 69.600 400.400 70.400 ;
        RECT 407.600 69.600 408.400 70.400 ;
        RECT 396.400 67.600 397.200 68.400 ;
        RECT 401.200 67.600 402.000 68.400 ;
        RECT 401.300 60.400 401.900 67.600 ;
        RECT 401.200 59.600 402.000 60.400 ;
        RECT 394.800 57.600 395.600 58.400 ;
        RECT 385.200 55.600 386.000 56.400 ;
        RECT 390.000 55.600 390.800 56.400 ;
        RECT 396.400 55.600 397.200 56.400 ;
        RECT 396.500 54.400 397.100 55.600 ;
        RECT 385.200 53.600 386.000 54.400 ;
        RECT 396.400 53.600 397.200 54.400 ;
        RECT 385.300 48.400 385.900 53.600 ;
        RECT 398.000 50.200 398.800 55.800 ;
        RECT 399.600 53.600 400.400 54.400 ;
        RECT 385.200 47.600 386.000 48.400 ;
        RECT 388.400 47.600 389.200 48.400 ;
        RECT 394.800 47.600 395.600 48.400 ;
        RECT 356.400 41.600 357.200 42.400 ;
        RECT 350.000 37.600 350.800 38.400 ;
        RECT 354.800 37.600 355.600 38.400 ;
        RECT 353.200 31.600 354.000 32.400 ;
        RECT 334.000 29.600 334.800 30.400 ;
        RECT 335.600 29.600 336.400 30.400 ;
        RECT 348.400 29.600 349.200 30.400 ;
        RECT 354.900 28.400 355.500 37.600 ;
        RECT 356.500 30.400 357.100 41.600 ;
        RECT 359.600 31.600 360.400 32.400 ;
        RECT 366.000 31.800 366.800 32.600 ;
        RECT 372.600 31.800 373.400 32.600 ;
        RECT 356.400 29.600 357.200 30.400 ;
        RECT 366.000 28.400 366.600 31.800 ;
        RECT 367.600 29.600 368.400 30.400 ;
        RECT 370.000 28.400 370.800 28.600 ;
        RECT 337.200 27.600 338.000 28.400 ;
        RECT 343.600 27.600 344.400 28.400 ;
        RECT 346.800 27.600 347.600 28.400 ;
        RECT 354.800 27.600 355.600 28.400 ;
        RECT 361.200 27.600 362.000 28.400 ;
        RECT 366.000 27.800 370.800 28.400 ;
        RECT 337.300 24.400 337.900 27.600 ;
        RECT 342.000 25.600 342.800 26.400 ;
        RECT 346.900 25.700 347.500 27.600 ;
        RECT 366.000 27.000 366.600 27.800 ;
        RECT 367.400 27.000 368.200 27.200 ;
        RECT 370.800 27.000 371.600 27.200 ;
        RECT 372.800 27.000 373.400 31.800 ;
        RECT 374.000 27.600 374.800 28.400 ;
        RECT 361.200 25.600 362.000 26.400 ;
        RECT 366.000 26.200 366.800 27.000 ;
        RECT 367.400 26.400 371.600 27.000 ;
        RECT 372.600 26.200 373.400 27.000 ;
        RECT 375.600 26.200 376.400 31.800 ;
        RECT 342.100 24.400 342.700 25.600 ;
        RECT 337.200 23.600 338.000 24.400 ;
        RECT 342.000 23.600 342.800 24.400 ;
        RECT 345.200 23.600 346.000 24.400 ;
        RECT 378.800 24.200 379.600 35.800 ;
        RECT 385.300 30.400 385.900 47.600 ;
        RECT 380.400 29.400 381.200 30.400 ;
        RECT 385.200 29.600 386.000 30.400 ;
        RECT 345.300 20.400 345.900 23.600 ;
        RECT 356.400 21.600 357.200 22.400 ;
        RECT 345.200 19.600 346.000 20.400 ;
        RECT 356.500 18.400 357.100 21.600 ;
        RECT 332.400 17.600 333.200 18.400 ;
        RECT 337.200 17.600 338.000 18.400 ;
        RECT 327.600 15.600 328.400 16.400 ;
        RECT 327.700 14.400 328.300 15.600 ;
        RECT 329.000 15.000 329.800 15.800 ;
        RECT 330.800 15.000 335.000 15.600 ;
        RECT 335.600 15.000 336.400 15.800 ;
        RECT 326.000 13.600 326.800 14.400 ;
        RECT 327.600 13.600 328.400 14.400 ;
        RECT 326.100 12.400 326.700 13.600 ;
        RECT 305.200 11.600 306.000 12.400 ;
        RECT 306.800 11.600 307.600 12.400 ;
        RECT 319.600 11.600 320.400 12.400 ;
        RECT 324.400 11.600 325.200 12.400 ;
        RECT 326.000 11.600 326.800 12.400 ;
        RECT 284.400 9.400 285.200 10.200 ;
        RECT 290.600 9.400 291.400 10.200 ;
        RECT 302.000 9.600 302.800 10.400 ;
        RECT 329.000 10.200 329.600 15.000 ;
        RECT 330.800 14.800 331.600 15.000 ;
        RECT 334.200 14.800 335.000 15.000 ;
        RECT 335.800 14.200 336.400 15.000 ;
        RECT 337.300 14.400 337.900 17.600 ;
        RECT 331.600 13.600 336.400 14.200 ;
        RECT 337.200 13.600 338.000 14.400 ;
        RECT 331.600 13.400 332.400 13.600 ;
        RECT 335.800 10.200 336.400 13.600 ;
        RECT 337.200 11.600 338.000 12.400 ;
        RECT 338.800 10.200 339.600 15.800 ;
        RECT 329.000 9.400 329.800 10.200 ;
        RECT 335.600 9.400 336.400 10.200 ;
        RECT 242.800 7.600 243.600 8.400 ;
        RECT 252.400 7.600 253.200 8.400 ;
        RECT 255.600 7.600 256.400 8.400 ;
        RECT 271.600 7.600 272.400 8.400 ;
        RECT 201.200 5.600 202.000 6.400 ;
        RECT 233.200 5.600 234.000 6.400 ;
        RECT 239.600 5.600 240.400 6.400 ;
        RECT 342.000 6.200 342.800 17.800 ;
        RECT 350.000 13.600 350.800 14.400 ;
        RECT 343.600 11.800 344.400 12.600 ;
        RECT 350.100 12.400 350.700 13.600 ;
        RECT 343.700 6.400 344.300 11.800 ;
        RECT 350.000 11.600 350.800 12.400 ;
        RECT 343.600 5.600 344.400 6.400 ;
        RECT 351.600 6.200 352.400 17.800 ;
        RECT 356.400 17.600 357.200 18.400 ;
        RECT 358.000 10.200 358.800 15.800 ;
        RECT 361.200 6.200 362.000 17.800 ;
        RECT 369.200 13.600 370.000 14.400 ;
        RECT 362.800 11.800 363.600 12.600 ;
        RECT 369.300 12.400 369.900 13.600 ;
        RECT 362.900 8.400 363.500 11.800 ;
        RECT 369.200 11.600 370.000 12.400 ;
        RECT 362.800 7.600 363.600 8.400 ;
        RECT 370.800 6.200 371.600 17.800 ;
        RECT 375.600 17.600 376.400 18.400 ;
        RECT 375.700 16.400 376.300 17.600 ;
        RECT 375.600 15.600 376.400 16.400 ;
        RECT 377.200 10.200 378.000 15.800 ;
        RECT 380.400 6.200 381.200 17.800 ;
        RECT 385.300 14.400 385.900 29.600 ;
        RECT 388.400 24.200 389.200 35.800 ;
        RECT 394.900 30.400 395.500 47.600 ;
        RECT 401.200 46.200 402.000 57.800 ;
        RECT 409.300 54.400 409.900 81.600 ;
        RECT 410.800 71.600 411.600 72.400 ;
        RECT 410.900 70.400 411.500 71.600 ;
        RECT 412.500 70.400 413.100 87.600 ;
        RECT 423.700 78.400 424.300 93.600 ;
        RECT 428.400 91.600 429.200 92.400 ;
        RECT 425.200 89.600 426.000 90.400 ;
        RECT 428.500 78.400 429.100 91.600 ;
        RECT 431.600 90.200 432.400 95.800 ;
        RECT 433.300 94.400 433.900 107.600 ;
        RECT 434.800 104.200 435.600 115.800 ;
        RECT 438.100 110.400 438.700 133.600 ;
        RECT 441.200 131.600 442.000 132.400 ;
        RECT 449.200 117.600 450.000 118.400 ;
        RECT 436.400 109.400 437.200 110.400 ;
        RECT 438.000 109.600 438.800 110.400 ;
        RECT 433.200 93.600 434.000 94.400 ;
        RECT 433.300 82.400 433.900 93.600 ;
        RECT 434.800 86.200 435.600 97.800 ;
        RECT 436.400 91.800 437.200 92.600 ;
        RECT 436.500 88.400 437.100 91.800 ;
        RECT 436.400 87.600 437.200 88.400 ;
        RECT 433.200 81.600 434.000 82.400 ;
        RECT 423.600 77.600 424.400 78.400 ;
        RECT 426.800 77.600 427.600 78.400 ;
        RECT 428.400 77.600 429.200 78.400 ;
        RECT 414.000 75.600 414.800 76.400 ;
        RECT 414.100 72.400 414.700 75.600 ;
        RECT 423.600 73.600 424.400 74.400 ;
        RECT 414.000 71.600 414.800 72.400 ;
        RECT 410.800 69.600 411.600 70.400 ;
        RECT 412.400 69.600 413.200 70.400 ;
        RECT 423.700 68.400 424.300 73.600 ;
        RECT 426.900 72.400 427.500 77.600 ;
        RECT 438.100 74.400 438.700 109.600 ;
        RECT 444.400 104.200 445.200 115.800 ;
        RECT 450.900 98.400 451.500 139.600 ;
        RECT 462.100 138.400 462.700 141.600 ;
        RECT 454.000 137.600 454.800 138.400 ;
        RECT 462.000 137.600 462.800 138.400 ;
        RECT 452.400 135.600 453.200 136.400 ;
        RECT 452.500 100.400 453.100 135.600 ;
        RECT 457.200 133.600 458.000 134.400 ;
        RECT 457.300 132.400 457.900 133.600 ;
        RECT 457.200 131.600 458.000 132.400 ;
        RECT 458.800 131.600 459.600 132.400 ;
        RECT 457.300 118.400 457.900 131.600 ;
        RECT 457.200 117.600 458.000 118.400 ;
        RECT 458.900 112.400 459.500 131.600 ;
        RECT 463.700 130.400 464.300 155.600 ;
        RECT 466.800 149.600 467.600 150.400 ;
        RECT 466.800 147.600 467.600 148.400 ;
        RECT 468.400 146.200 469.200 151.800 ;
        RECT 470.100 148.400 470.700 163.700 ;
        RECT 470.000 147.600 470.800 148.400 ;
        RECT 471.600 144.200 472.400 155.800 ;
        RECT 473.200 149.400 474.000 150.400 ;
        RECT 478.000 149.600 478.800 150.400 ;
        RECT 474.800 147.600 475.600 148.400 ;
        RECT 474.900 138.400 475.500 147.600 ;
        RECT 479.700 138.400 480.300 173.600 ;
        RECT 481.000 170.200 481.600 175.000 ;
        RECT 482.800 174.800 483.600 175.000 ;
        RECT 486.200 174.800 487.000 175.000 ;
        RECT 487.800 174.200 488.400 175.000 ;
        RECT 489.300 174.400 489.900 183.600 ;
        RECT 492.500 178.400 493.100 183.600 ;
        RECT 492.400 177.600 493.200 178.400 ;
        RECT 494.100 174.400 494.700 185.600 ;
        RECT 498.900 182.400 499.500 187.600 ;
        RECT 500.400 187.000 501.000 187.800 ;
        RECT 501.800 187.000 502.600 187.200 ;
        RECT 505.200 187.000 506.000 187.200 ;
        RECT 507.200 187.000 507.800 191.800 ;
        RECT 511.600 191.600 512.400 192.400 ;
        RECT 514.800 191.600 515.600 192.400 ;
        RECT 518.000 191.600 518.800 192.400 ;
        RECT 519.600 191.600 520.400 192.400 ;
        RECT 516.400 189.600 517.200 190.400 ;
        RECT 508.400 187.600 509.200 188.400 ;
        RECT 500.400 186.200 501.200 187.000 ;
        RECT 501.800 186.400 506.000 187.000 ;
        RECT 507.000 186.200 507.800 187.000 ;
        RECT 510.000 185.600 510.800 186.400 ;
        RECT 513.200 185.600 514.000 186.400 ;
        RECT 498.800 181.600 499.600 182.400 ;
        RECT 508.400 181.600 509.200 182.400 ;
        RECT 503.600 179.600 504.400 180.400 ;
        RECT 500.400 177.600 501.200 178.400 ;
        RECT 502.000 175.600 502.800 176.400 ;
        RECT 483.600 173.600 488.400 174.200 ;
        RECT 489.200 173.600 490.000 174.400 ;
        RECT 490.800 173.600 491.600 174.400 ;
        RECT 494.000 173.600 494.800 174.400 ;
        RECT 483.600 173.400 484.400 173.600 ;
        RECT 487.800 170.200 488.400 173.600 ;
        RECT 481.000 169.400 481.800 170.200 ;
        RECT 487.600 169.400 488.400 170.200 ;
        RECT 490.900 158.400 491.500 173.600 ;
        RECT 498.800 169.600 499.600 170.400 ;
        RECT 486.000 157.600 486.800 158.400 ;
        RECT 490.800 157.600 491.600 158.400 ;
        RECT 481.200 144.200 482.000 155.800 ;
        RECT 487.600 149.600 488.400 150.400 ;
        RECT 474.800 137.600 475.600 138.400 ;
        RECT 479.600 137.600 480.400 138.400 ;
        RECT 466.800 135.600 467.600 136.400 ;
        RECT 466.900 134.400 467.500 135.600 ;
        RECT 466.800 133.600 467.600 134.400 ;
        RECT 468.400 133.600 469.200 134.400 ;
        RECT 468.500 132.400 469.100 133.600 ;
        RECT 468.400 131.600 469.200 132.400 ;
        RECT 471.600 131.600 472.400 132.400 ;
        RECT 474.800 131.600 475.600 132.400 ;
        RECT 463.600 129.600 464.400 130.400 ;
        RECT 465.200 129.600 466.000 130.400 ;
        RECT 471.600 129.600 472.400 130.400 ;
        RECT 473.200 129.600 474.000 130.400 ;
        RECT 463.700 118.400 464.300 129.600 ;
        RECT 463.600 117.600 464.400 118.400 ;
        RECT 473.300 114.400 473.900 129.600 ;
        RECT 476.400 127.600 477.200 128.400 ;
        RECT 484.400 126.200 485.200 137.800 ;
        RECT 490.900 134.400 491.500 157.600 ;
        RECT 502.100 152.400 502.700 175.600 ;
        RECT 503.700 172.400 504.300 179.600 ;
        RECT 508.500 178.400 509.100 181.600 ;
        RECT 506.800 177.600 507.600 178.400 ;
        RECT 508.400 177.600 509.200 178.400 ;
        RECT 506.900 174.400 507.500 177.600 ;
        RECT 510.100 176.400 510.700 185.600 ;
        RECT 516.500 184.400 517.100 189.600 ;
        RECT 514.800 183.600 515.600 184.400 ;
        RECT 516.400 183.600 517.200 184.400 ;
        RECT 518.000 183.600 518.800 184.400 ;
        RECT 514.900 176.400 515.500 183.600 ;
        RECT 518.100 176.400 518.700 183.600 ;
        RECT 519.700 178.400 520.300 191.600 ;
        RECT 521.300 188.400 521.900 211.600 ;
        RECT 523.200 210.200 523.800 215.000 ;
        RECT 524.500 214.400 525.100 215.600 ;
        RECT 524.400 213.600 525.200 214.400 ;
        RECT 527.600 213.600 528.400 214.400 ;
        RECT 530.800 213.600 531.600 214.400 ;
        RECT 532.400 213.600 533.200 214.400 ;
        RECT 527.700 212.400 528.300 213.600 ;
        RECT 524.400 211.600 525.200 212.400 ;
        RECT 527.600 211.600 528.400 212.400 ;
        RECT 523.000 209.400 523.800 210.200 ;
        RECT 524.500 198.400 525.100 211.600 ;
        RECT 527.600 199.600 528.400 200.400 ;
        RECT 524.400 197.600 525.200 198.400 ;
        RECT 527.700 188.400 528.300 199.600 ;
        RECT 530.900 188.400 531.500 213.600 ;
        RECT 532.500 194.400 533.100 213.600 ;
        RECT 534.000 211.600 534.800 212.400 ;
        RECT 534.100 210.400 534.700 211.600 ;
        RECT 534.000 209.600 534.800 210.400 ;
        RECT 534.100 198.400 534.700 209.600 ;
        RECT 534.000 197.600 534.800 198.400 ;
        RECT 535.700 196.300 536.300 253.600 ;
        RECT 537.200 250.200 538.000 255.800 ;
        RECT 540.400 246.200 541.200 257.800 ;
        RECT 543.700 254.400 544.300 267.600 ;
        RECT 545.200 264.200 546.000 275.800 ;
        RECT 551.700 270.400 552.300 295.600 ;
        RECT 553.200 286.200 554.000 297.800 ;
        RECT 556.400 286.200 557.200 297.800 ;
        RECT 558.000 284.200 558.800 297.800 ;
        RECT 559.600 284.200 560.400 297.800 ;
        RECT 561.300 278.400 561.900 331.600 ;
        RECT 569.200 326.200 570.000 337.800 ;
        RECT 572.400 330.200 573.200 335.800 ;
        RECT 578.900 332.400 579.500 343.600 ;
        RECT 574.000 331.600 574.800 332.400 ;
        RECT 578.800 331.600 579.600 332.400 ;
        RECT 562.800 313.600 563.600 314.400 ;
        RECT 562.900 312.400 563.500 313.600 ;
        RECT 562.800 311.600 563.600 312.400 ;
        RECT 564.400 306.200 565.200 311.800 ;
        RECT 566.000 307.600 566.800 308.400 ;
        RECT 567.600 304.200 568.400 315.800 ;
        RECT 569.200 311.600 570.000 312.400 ;
        RECT 569.300 310.200 569.900 311.600 ;
        RECT 569.200 309.400 570.000 310.200 ;
        RECT 574.100 296.400 574.700 331.600 ;
        RECT 577.200 304.200 578.000 315.800 ;
        RECT 578.800 305.600 579.600 306.400 ;
        RECT 578.900 296.400 579.500 305.600 ;
        RECT 582.000 303.600 582.800 304.400 ;
        RECT 574.000 295.600 574.800 296.400 ;
        RECT 578.800 295.600 579.600 296.400 ;
        RECT 564.400 291.600 565.200 292.400 ;
        RECT 574.000 291.600 574.800 292.400 ;
        RECT 580.400 291.600 581.200 292.400 ;
        RECT 564.400 289.600 565.200 290.400 ;
        RECT 569.200 289.600 570.000 290.400 ;
        RECT 580.500 288.400 581.100 291.600 ;
        RECT 580.400 287.600 581.200 288.400 ;
        RECT 561.200 277.600 562.000 278.400 ;
        RECT 546.800 269.400 547.600 270.400 ;
        RECT 551.600 269.600 552.400 270.400 ;
        RECT 554.800 264.200 555.600 275.800 ;
        RECT 559.600 273.600 560.400 274.400 ;
        RECT 559.700 272.400 560.300 273.600 ;
        RECT 559.600 271.600 560.400 272.400 ;
        RECT 561.200 266.200 562.000 271.800 ;
        RECT 562.800 267.600 563.600 268.400 ;
        RECT 556.400 261.600 557.200 262.400 ;
        RECT 543.600 253.600 544.400 254.400 ;
        RECT 542.000 251.800 542.800 252.600 ;
        RECT 537.200 224.200 538.000 235.800 ;
        RECT 538.800 229.400 539.600 230.400 ;
        RECT 542.100 218.400 542.700 251.800 ;
        RECT 543.700 230.400 544.300 253.600 ;
        RECT 550.000 246.200 550.800 257.800 ;
        RECT 556.500 252.400 557.100 261.600 ;
        RECT 556.400 251.600 557.200 252.400 ;
        RECT 561.200 250.200 562.000 255.800 ;
        RECT 562.900 254.400 563.500 267.600 ;
        RECT 564.400 264.200 565.200 275.800 ;
        RECT 566.000 271.600 566.800 272.400 ;
        RECT 566.100 270.200 566.700 271.600 ;
        RECT 566.000 269.400 566.800 270.200 ;
        RECT 574.000 264.200 574.800 275.800 ;
        RECT 578.800 274.300 579.600 274.400 ;
        RECT 578.800 273.700 581.100 274.300 ;
        RECT 578.800 273.600 579.600 273.700 ;
        RECT 580.500 270.400 581.100 273.700 ;
        RECT 580.400 269.600 581.200 270.400 ;
        RECT 577.200 263.600 578.000 264.400 ;
        RECT 562.800 253.600 563.600 254.400 ;
        RECT 554.800 247.600 555.600 248.400 ;
        RECT 564.400 246.200 565.200 257.800 ;
        RECT 566.000 251.800 566.800 252.600 ;
        RECT 566.100 248.400 566.700 251.800 ;
        RECT 566.000 247.600 566.800 248.400 ;
        RECT 574.000 246.200 574.800 257.800 ;
        RECT 543.600 229.600 544.400 230.400 ;
        RECT 546.800 224.200 547.600 235.800 ;
        RECT 551.600 233.600 552.400 234.400 ;
        RECT 551.700 232.400 552.300 233.600 ;
        RECT 551.600 231.600 552.400 232.400 ;
        RECT 553.200 226.200 554.000 231.800 ;
        RECT 554.800 227.600 555.600 228.400 ;
        RECT 542.000 217.600 542.800 218.400 ;
        RECT 537.200 213.600 538.000 214.400 ;
        RECT 537.200 211.600 538.000 212.400 ;
        RECT 537.300 198.400 537.900 211.600 ;
        RECT 538.800 209.600 539.600 210.400 ;
        RECT 542.000 209.600 542.800 210.400 ;
        RECT 543.600 210.200 544.400 215.800 ;
        RECT 546.800 206.200 547.600 217.800 ;
        RECT 548.400 211.800 549.200 212.600 ;
        RECT 554.900 212.400 555.500 227.600 ;
        RECT 556.400 224.200 557.200 235.800 ;
        RECT 558.000 231.600 558.800 232.400 ;
        RECT 558.100 230.200 558.700 231.600 ;
        RECT 558.000 229.400 558.800 230.200 ;
        RECT 564.400 227.600 565.200 228.400 ;
        RECT 548.500 208.400 549.100 211.800 ;
        RECT 554.800 211.600 555.600 212.400 ;
        RECT 548.400 207.600 549.200 208.400 ;
        RECT 556.400 206.200 557.200 217.800 ;
        RECT 562.800 210.200 563.600 215.800 ;
        RECT 564.500 214.400 565.100 227.600 ;
        RECT 566.000 224.200 566.800 235.800 ;
        RECT 570.800 234.300 571.600 234.400 ;
        RECT 570.800 233.700 573.100 234.300 ;
        RECT 570.800 233.600 571.600 233.700 ;
        RECT 572.500 230.400 573.100 233.700 ;
        RECT 577.300 230.400 577.900 263.600 ;
        RECT 580.400 251.600 581.200 252.400 ;
        RECT 578.800 248.300 579.600 248.400 ;
        RECT 580.500 248.300 581.100 251.600 ;
        RECT 578.800 247.700 581.100 248.300 ;
        RECT 578.800 247.600 579.600 247.700 ;
        RECT 572.400 229.600 573.200 230.400 ;
        RECT 577.200 229.600 578.000 230.400 ;
        RECT 564.400 213.600 565.200 214.400 ;
        RECT 561.200 207.600 562.000 208.400 ;
        RECT 566.000 206.200 566.800 217.800 ;
        RECT 567.600 213.600 568.400 214.400 ;
        RECT 537.200 197.600 538.000 198.400 ;
        RECT 534.100 195.700 536.300 196.300 ;
        RECT 532.400 193.600 533.200 194.400 ;
        RECT 532.500 188.400 533.100 193.600 ;
        RECT 521.200 187.600 522.000 188.400 ;
        RECT 527.600 187.600 528.400 188.400 ;
        RECT 530.800 187.600 531.600 188.400 ;
        RECT 532.400 187.600 533.200 188.400 ;
        RECT 521.200 185.600 522.000 186.400 ;
        RECT 524.400 185.600 525.200 186.400 ;
        RECT 526.000 185.600 526.800 186.400 ;
        RECT 519.600 177.600 520.400 178.400 ;
        RECT 510.000 175.600 510.800 176.400 ;
        RECT 511.600 175.600 512.400 176.400 ;
        RECT 514.800 175.600 515.600 176.400 ;
        RECT 518.000 175.600 518.800 176.400 ;
        RECT 505.200 173.600 506.000 174.400 ;
        RECT 506.800 173.600 507.600 174.400 ;
        RECT 503.600 171.600 504.400 172.400 ;
        RECT 505.300 170.400 505.900 173.600 ;
        RECT 511.700 172.400 512.300 175.600 ;
        RECT 513.200 174.300 514.000 174.400 ;
        RECT 513.200 173.700 515.500 174.300 ;
        RECT 513.200 173.600 514.000 173.700 ;
        RECT 508.400 171.600 509.200 172.400 ;
        RECT 511.600 171.600 512.400 172.400 ;
        RECT 505.200 169.600 506.000 170.400 ;
        RECT 505.200 155.600 506.000 156.400 ;
        RECT 502.000 151.600 502.800 152.400 ;
        RECT 490.800 133.600 491.600 134.400 ;
        RECT 490.800 131.600 491.600 132.400 ;
        RECT 479.600 115.600 480.400 116.400 ;
        RECT 473.200 113.600 474.000 114.400 ;
        RECT 458.800 111.600 459.600 112.400 ;
        RECT 470.000 111.800 470.800 112.600 ;
        RECT 476.200 111.800 477.000 112.600 ;
        RECT 458.900 110.400 459.500 111.600 ;
        RECT 458.800 109.600 459.600 110.400 ;
        RECT 462.000 109.600 462.800 110.400 ;
        RECT 466.800 109.600 467.600 110.400 ;
        RECT 462.100 108.400 462.700 109.600 ;
        RECT 458.800 107.600 459.600 108.400 ;
        RECT 462.000 107.600 462.800 108.400 ;
        RECT 458.900 100.400 459.500 107.600 ;
        RECT 462.100 106.400 462.700 107.600 ;
        RECT 462.000 105.600 462.800 106.400 ;
        RECT 466.900 104.400 467.500 109.600 ;
        RECT 470.000 108.400 470.600 111.800 ;
        RECT 473.200 109.600 474.000 110.400 ;
        RECT 475.000 109.800 475.800 110.600 ;
        RECT 475.000 108.400 475.600 109.800 ;
        RECT 468.400 107.600 469.200 108.400 ;
        RECT 470.000 107.800 475.600 108.400 ;
        RECT 466.800 103.600 467.600 104.400 ;
        RECT 462.000 101.600 462.800 102.400 ;
        RECT 452.400 99.600 453.200 100.400 ;
        RECT 458.800 99.600 459.600 100.400 ;
        RECT 462.100 98.400 462.700 101.600 ;
        RECT 466.800 99.600 467.600 100.400 ;
        RECT 444.400 86.200 445.200 97.800 ;
        RECT 450.800 97.600 451.600 98.400 ;
        RECT 462.000 97.600 462.800 98.400 ;
        RECT 457.200 95.000 458.000 95.800 ;
        RECT 458.600 95.000 462.800 95.600 ;
        RECT 463.800 95.000 464.600 95.800 ;
        RECT 465.200 95.600 466.000 96.400 ;
        RECT 452.400 93.600 453.200 94.400 ;
        RECT 457.200 94.200 457.800 95.000 ;
        RECT 458.600 94.800 459.400 95.000 ;
        RECT 462.000 94.800 462.800 95.000 ;
        RECT 457.200 93.600 462.000 94.200 ;
        RECT 438.000 73.600 438.800 74.400 ;
        RECT 426.800 71.600 427.600 72.400 ;
        RECT 428.400 71.600 429.200 72.400 ;
        RECT 439.600 71.800 440.400 72.600 ;
        RECT 445.800 71.800 446.600 72.600 ;
        RECT 412.400 67.600 413.200 68.400 ;
        RECT 423.600 67.600 424.400 68.400 ;
        RECT 412.500 62.400 413.100 67.600 ;
        RECT 415.600 65.600 416.400 66.400 ;
        RECT 422.000 65.600 422.800 66.400 ;
        RECT 426.800 65.600 427.600 66.400 ;
        RECT 412.400 61.600 413.200 62.400 ;
        RECT 409.200 53.600 410.000 54.400 ;
        RECT 402.800 51.800 403.600 52.600 ;
        RECT 402.900 44.400 403.500 51.800 ;
        RECT 410.800 46.200 411.600 57.800 ;
        RECT 412.500 56.400 413.100 61.600 ;
        RECT 415.700 58.400 416.300 65.600 ;
        RECT 420.400 63.600 421.200 64.400 ;
        RECT 422.100 60.400 422.700 65.600 ;
        RECT 422.000 59.600 422.800 60.400 ;
        RECT 423.600 59.600 424.400 60.400 ;
        RECT 415.600 57.600 416.400 58.400 ;
        RECT 415.700 56.400 416.300 57.600 ;
        RECT 412.400 55.600 413.200 56.400 ;
        RECT 415.600 55.600 416.400 56.400 ;
        RECT 422.000 53.600 422.800 54.400 ;
        RECT 417.200 51.600 418.000 52.400 ;
        RECT 417.300 48.400 417.900 51.600 ;
        RECT 417.200 47.600 418.000 48.400 ;
        RECT 402.800 43.600 403.600 44.400 ;
        RECT 417.300 34.400 417.900 47.600 ;
        RECT 418.800 39.600 419.600 40.400 ;
        RECT 418.900 38.400 419.500 39.600 ;
        RECT 418.800 37.600 419.600 38.400 ;
        RECT 417.200 33.600 418.000 34.400 ;
        RECT 402.600 31.800 403.400 32.600 ;
        RECT 409.200 31.800 410.000 32.600 ;
        RECT 422.100 32.400 422.700 53.600 ;
        RECT 394.800 29.600 395.600 30.400 ;
        RECT 393.200 23.600 394.000 24.400 ;
        RECT 385.200 13.600 386.000 14.400 ;
        RECT 382.000 11.600 382.800 12.600 ;
        RECT 390.000 6.200 390.800 17.800 ;
        RECT 394.900 14.300 395.500 29.600 ;
        RECT 402.600 27.000 403.200 31.800 ;
        RECT 405.200 28.400 406.000 28.600 ;
        RECT 409.400 28.400 410.000 31.800 ;
        RECT 415.600 31.600 416.400 32.400 ;
        RECT 422.000 31.600 422.800 32.400 ;
        RECT 412.400 29.600 413.200 30.400 ;
        RECT 405.200 27.800 410.000 28.400 ;
        RECT 404.400 27.000 405.200 27.200 ;
        RECT 407.800 27.000 408.600 27.200 ;
        RECT 409.400 27.000 410.000 27.800 ;
        RECT 410.800 27.600 411.600 28.400 ;
        RECT 412.400 27.600 413.200 28.400 ;
        RECT 414.000 27.600 414.800 28.400 ;
        RECT 415.700 28.300 416.300 31.600 ;
        RECT 418.800 29.600 419.600 30.400 ;
        RECT 422.000 29.600 422.800 30.400 ;
        RECT 417.200 28.300 418.000 28.400 ;
        RECT 415.700 27.700 418.000 28.300 ;
        RECT 417.200 27.600 418.000 27.700 ;
        RECT 402.600 26.200 403.400 27.000 ;
        RECT 404.400 26.400 408.600 27.000 ;
        RECT 407.600 25.600 408.400 26.400 ;
        RECT 409.200 26.200 410.000 27.000 ;
        RECT 410.900 22.400 411.500 27.600 ;
        RECT 412.500 26.400 413.100 27.600 ;
        RECT 412.400 25.600 413.200 26.400 ;
        RECT 410.800 21.600 411.600 22.400 ;
        RECT 409.200 19.600 410.000 20.400 ;
        RECT 409.300 18.400 409.900 19.600 ;
        RECT 409.200 17.600 410.000 18.400 ;
        RECT 402.800 15.600 403.600 16.400 ;
        RECT 402.900 14.400 403.500 15.600 ;
        RECT 404.400 15.000 405.200 15.800 ;
        RECT 410.600 15.600 411.400 15.800 ;
        RECT 414.000 15.600 414.800 16.400 ;
        RECT 415.600 15.600 416.400 16.400 ;
        RECT 405.800 15.000 411.400 15.600 ;
        RECT 394.900 13.700 397.100 14.300 ;
        RECT 396.500 12.400 397.100 13.700 ;
        RECT 401.200 13.600 402.000 14.400 ;
        RECT 402.800 13.600 403.600 14.400 ;
        RECT 404.400 14.200 405.000 15.000 ;
        RECT 405.800 14.800 406.600 15.000 ;
        RECT 409.200 14.800 410.000 15.000 ;
        RECT 404.400 13.600 410.000 14.200 ;
        RECT 394.800 11.600 395.600 12.400 ;
        RECT 396.400 11.600 397.200 12.400 ;
        RECT 394.900 8.400 395.500 11.600 ;
        RECT 404.400 10.200 405.000 13.600 ;
        RECT 409.400 12.200 410.000 13.600 ;
        RECT 409.400 11.400 410.200 12.200 ;
        RECT 410.800 10.200 411.400 15.000 ;
        RECT 417.300 14.400 417.900 27.600 ;
        RECT 418.900 22.400 419.500 29.600 ;
        RECT 418.800 21.600 419.600 22.400 ;
        RECT 412.400 13.600 413.200 14.400 ;
        RECT 417.200 13.600 418.000 14.400 ;
        RECT 412.500 10.400 413.100 13.600 ;
        RECT 418.900 12.400 419.500 21.600 ;
        RECT 423.700 20.300 424.300 59.600 ;
        RECT 425.000 55.000 425.800 55.800 ;
        RECT 428.500 55.600 429.100 71.600 ;
        RECT 431.600 69.600 432.400 70.400 ;
        RECT 438.000 69.600 438.800 70.400 ;
        RECT 439.600 68.400 440.200 71.800 ;
        RECT 444.600 69.800 445.400 70.600 ;
        RECT 444.600 68.400 445.200 69.800 ;
        RECT 438.000 67.600 438.800 68.400 ;
        RECT 439.600 67.800 445.200 68.400 ;
        RECT 430.000 65.600 430.800 66.400 ;
        RECT 436.400 65.600 437.200 66.400 ;
        RECT 436.500 64.400 437.100 65.600 ;
        RECT 434.800 63.600 435.600 64.400 ;
        RECT 436.400 63.600 437.200 64.400 ;
        RECT 434.900 58.400 435.500 63.600 ;
        RECT 434.800 57.600 435.600 58.400 ;
        RECT 438.100 56.400 438.700 67.600 ;
        RECT 439.600 67.000 440.200 67.800 ;
        RECT 441.000 67.000 441.800 67.200 ;
        RECT 444.400 67.000 445.200 67.200 ;
        RECT 446.000 67.000 446.600 71.800 ;
        RECT 452.500 70.400 453.100 93.600 ;
        RECT 457.200 90.200 457.800 93.600 ;
        RECT 461.200 93.400 462.000 93.600 ;
        RECT 464.000 90.200 464.600 95.000 ;
        RECT 465.300 94.400 465.900 95.600 ;
        RECT 466.900 94.400 467.500 99.600 ;
        RECT 468.500 98.400 469.100 107.600 ;
        RECT 470.000 107.000 470.600 107.800 ;
        RECT 471.400 107.000 472.200 107.200 ;
        RECT 474.800 107.000 475.600 107.200 ;
        RECT 476.400 107.000 477.000 111.800 ;
        RECT 479.700 108.400 480.300 115.600 ;
        RECT 478.000 107.600 478.800 108.400 ;
        RECT 479.600 107.600 480.400 108.400 ;
        RECT 470.000 106.200 470.800 107.000 ;
        RECT 471.400 106.400 477.000 107.000 ;
        RECT 478.100 106.400 478.700 107.600 ;
        RECT 476.200 106.200 477.000 106.400 ;
        RECT 478.000 105.600 478.800 106.400 ;
        RECT 479.700 100.400 480.300 107.600 ;
        RECT 484.400 106.200 485.200 111.800 ;
        RECT 486.000 111.600 486.800 112.400 ;
        RECT 481.200 103.600 482.000 104.400 ;
        RECT 479.600 99.600 480.400 100.400 ;
        RECT 468.400 97.600 469.200 98.400 ;
        RECT 478.000 97.600 478.800 98.400 ;
        RECT 478.100 96.400 478.700 97.600 ;
        RECT 468.200 95.000 469.000 95.800 ;
        RECT 470.000 95.000 474.200 95.600 ;
        RECT 474.800 95.000 475.600 95.800 ;
        RECT 478.000 95.600 478.800 96.400 ;
        RECT 479.600 95.600 480.400 96.400 ;
        RECT 465.200 93.600 466.000 94.400 ;
        RECT 466.800 93.600 467.600 94.400 ;
        RECT 457.200 89.400 458.000 90.200 ;
        RECT 463.800 89.400 464.600 90.200 ;
        RECT 468.200 90.200 468.800 95.000 ;
        RECT 470.000 94.800 470.800 95.000 ;
        RECT 473.400 94.800 474.200 95.000 ;
        RECT 475.000 94.200 475.600 95.000 ;
        RECT 470.800 93.600 475.600 94.200 ;
        RECT 476.400 93.600 477.200 94.400 ;
        RECT 470.800 93.400 471.600 93.600 ;
        RECT 475.000 90.200 475.600 93.600 ;
        RECT 468.200 89.400 469.000 90.200 ;
        RECT 474.800 89.400 475.600 90.200 ;
        RECT 468.400 87.600 469.200 88.400 ;
        RECT 468.500 78.400 469.100 87.600 ;
        RECT 468.400 77.600 469.200 78.400 ;
        RECT 460.400 73.600 461.200 74.400 ;
        RECT 452.400 69.600 453.200 70.400 ;
        RECT 455.600 69.600 456.400 70.400 ;
        RECT 458.800 69.600 459.600 70.400 ;
        RECT 455.700 68.400 456.300 69.600 ;
        RECT 460.500 68.400 461.100 73.600 ;
        RECT 463.400 71.800 464.200 72.600 ;
        RECT 470.000 71.800 470.800 72.600 ;
        RECT 447.600 67.600 448.400 68.400 ;
        RECT 450.800 67.600 451.600 68.400 ;
        RECT 455.600 67.600 456.400 68.400 ;
        RECT 457.200 67.600 458.000 68.400 ;
        RECT 458.800 67.600 459.600 68.400 ;
        RECT 460.400 67.600 461.200 68.400 ;
        RECT 462.000 67.600 462.800 68.400 ;
        RECT 439.600 66.200 440.400 67.000 ;
        RECT 441.000 66.400 446.600 67.000 ;
        RECT 445.800 66.200 446.600 66.400 ;
        RECT 441.200 63.600 442.000 64.400 ;
        RECT 439.600 57.600 440.400 58.400 ;
        RECT 426.800 55.000 431.000 55.600 ;
        RECT 431.600 55.000 432.400 55.800 ;
        RECT 433.200 55.600 434.000 56.400 ;
        RECT 438.000 55.600 438.800 56.400 ;
        RECT 425.000 50.200 425.600 55.000 ;
        RECT 426.800 54.800 427.600 55.000 ;
        RECT 430.200 54.800 431.000 55.000 ;
        RECT 431.800 54.200 432.400 55.000 ;
        RECT 433.300 54.400 433.900 55.600 ;
        RECT 427.600 53.600 432.400 54.200 ;
        RECT 433.200 53.600 434.000 54.400 ;
        RECT 434.800 53.600 435.600 54.400 ;
        RECT 427.600 53.400 428.400 53.600 ;
        RECT 425.000 49.400 425.800 50.200 ;
        RECT 430.000 49.600 430.800 50.400 ;
        RECT 431.800 50.200 432.400 53.600 ;
        RECT 425.200 35.600 426.000 36.400 ;
        RECT 425.300 30.400 425.900 35.600 ;
        RECT 425.200 29.600 426.000 30.400 ;
        RECT 426.800 29.600 427.600 30.400 ;
        RECT 425.200 23.600 426.000 24.400 ;
        RECT 422.100 19.700 424.300 20.300 ;
        RECT 422.100 14.400 422.700 19.700 ;
        RECT 423.600 17.600 424.400 18.400 ;
        RECT 422.000 13.600 422.800 14.400 ;
        RECT 418.800 11.600 419.600 12.400 ;
        RECT 422.100 10.400 422.700 13.600 ;
        RECT 425.300 12.300 425.900 23.600 ;
        RECT 426.900 20.400 427.500 29.600 ;
        RECT 428.400 27.600 429.200 28.400 ;
        RECT 426.800 19.600 427.600 20.400 ;
        RECT 430.100 16.300 430.700 49.600 ;
        RECT 431.600 49.400 432.400 50.200 ;
        RECT 436.400 43.600 437.200 44.400 ;
        RECT 431.600 37.600 432.400 38.400 ;
        RECT 431.700 32.400 432.300 37.600 ;
        RECT 436.400 35.600 437.200 36.400 ;
        RECT 431.600 31.600 432.400 32.400 ;
        RECT 439.700 30.400 440.300 57.600 ;
        RECT 441.300 56.400 441.900 63.600 ;
        RECT 441.200 55.600 442.000 56.400 ;
        RECT 447.700 46.400 448.300 67.600 ;
        RECT 450.900 60.400 451.500 67.600 ;
        RECT 454.000 65.600 454.800 66.400 ;
        RECT 450.800 59.600 451.600 60.400 ;
        RECT 449.200 53.600 450.000 54.400 ;
        RECT 450.900 48.300 451.500 59.600 ;
        RECT 454.100 58.400 454.700 65.600 ;
        RECT 455.700 58.400 456.300 67.600 ;
        RECT 452.400 57.600 453.200 58.400 ;
        RECT 454.000 57.600 454.800 58.400 ;
        RECT 455.600 57.600 456.400 58.400 ;
        RECT 452.500 50.400 453.100 57.600 ;
        RECT 457.300 56.400 457.900 67.600 ;
        RECT 457.200 55.600 458.000 56.400 ;
        RECT 458.900 54.400 459.500 67.600 ;
        RECT 462.100 66.400 462.700 67.600 ;
        RECT 463.400 67.000 464.000 71.800 ;
        RECT 466.000 68.400 466.800 68.600 ;
        RECT 470.200 68.400 470.800 71.800 ;
        RECT 474.800 72.300 475.600 72.400 ;
        RECT 476.500 72.300 477.100 93.600 ;
        RECT 478.100 92.400 478.700 95.600 ;
        RECT 478.000 91.600 478.800 92.400 ;
        RECT 482.800 91.600 483.600 92.400 ;
        RECT 478.100 74.400 478.700 91.600 ;
        RECT 482.900 84.400 483.500 91.600 ;
        RECT 484.400 87.600 485.200 88.400 ;
        RECT 484.500 86.400 485.100 87.600 ;
        RECT 484.400 85.600 485.200 86.400 ;
        RECT 482.800 83.600 483.600 84.400 ;
        RECT 479.600 75.600 480.400 76.400 ;
        RECT 478.000 73.600 478.800 74.400 ;
        RECT 474.800 71.700 477.100 72.300 ;
        RECT 474.800 71.600 475.600 71.700 ;
        RECT 478.000 71.600 478.800 72.400 ;
        RECT 474.900 70.400 475.500 71.600 ;
        RECT 474.800 69.600 475.600 70.400 ;
        RECT 478.100 68.400 478.700 71.600 ;
        RECT 466.000 67.800 470.800 68.400 ;
        RECT 465.200 67.000 466.000 67.200 ;
        RECT 468.600 67.000 469.400 67.200 ;
        RECT 470.200 67.000 470.800 67.800 ;
        RECT 471.600 67.600 472.400 68.400 ;
        RECT 473.200 67.600 474.000 68.400 ;
        RECT 478.000 67.600 478.800 68.400 ;
        RECT 462.000 65.600 462.800 66.400 ;
        RECT 463.400 66.200 464.200 67.000 ;
        RECT 465.200 66.400 469.400 67.000 ;
        RECT 470.000 66.200 470.800 67.000 ;
        RECT 471.700 66.400 472.300 67.600 ;
        RECT 471.600 65.600 472.400 66.400 ;
        RECT 473.300 62.400 473.900 67.600 ;
        RECT 479.700 66.400 480.300 75.600 ;
        RECT 484.400 70.300 485.200 70.400 ;
        RECT 486.100 70.300 486.700 111.600 ;
        RECT 487.600 104.200 488.400 115.800 ;
        RECT 489.200 109.400 490.000 110.200 ;
        RECT 489.300 102.400 489.900 109.400 ;
        RECT 489.200 101.600 490.000 102.400 ;
        RECT 490.900 98.400 491.500 131.600 ;
        RECT 494.000 126.200 494.800 137.800 ;
        RECT 495.600 133.600 496.400 134.400 ;
        RECT 495.700 110.400 496.300 133.600 ;
        RECT 497.200 130.200 498.000 135.800 ;
        RECT 502.100 118.400 502.700 151.600 ;
        RECT 505.300 148.400 505.900 155.600 ;
        RECT 506.800 149.600 507.600 150.400 ;
        RECT 508.500 148.400 509.100 171.600 ;
        RECT 511.700 170.400 512.300 171.600 ;
        RECT 510.000 169.600 510.800 170.400 ;
        RECT 511.600 169.600 512.400 170.400 ;
        RECT 510.100 168.400 510.700 169.600 ;
        RECT 510.000 167.600 510.800 168.400 ;
        RECT 511.700 148.400 512.300 169.600 ;
        RECT 513.200 167.600 514.000 168.400 ;
        RECT 513.300 160.400 513.900 167.600 ;
        RECT 514.900 164.400 515.500 173.700 ;
        RECT 516.400 173.600 517.200 174.400 ;
        RECT 516.500 168.400 517.100 173.600 ;
        RECT 518.000 171.600 518.800 172.400 ;
        RECT 519.600 169.600 520.400 170.400 ;
        RECT 516.400 167.600 517.200 168.400 ;
        RECT 514.800 163.600 515.600 164.400 ;
        RECT 513.200 159.600 514.000 160.400 ;
        RECT 519.600 155.600 520.400 156.400 ;
        RECT 513.200 151.600 514.000 152.400 ;
        RECT 513.300 150.400 513.900 151.600 ;
        RECT 513.200 149.600 514.000 150.400 ;
        RECT 516.400 149.600 517.200 150.400 ;
        RECT 505.200 147.600 506.000 148.400 ;
        RECT 508.400 147.600 509.200 148.400 ;
        RECT 511.600 147.600 512.400 148.400 ;
        RECT 514.800 147.600 515.600 148.400 ;
        RECT 510.000 143.600 510.800 144.400 ;
        RECT 510.100 140.400 510.700 143.600 ;
        RECT 510.000 139.600 510.800 140.400 ;
        RECT 514.900 138.400 515.500 147.600 ;
        RECT 516.500 146.400 517.100 149.600 ;
        RECT 516.400 145.600 517.200 146.400 ;
        RECT 514.800 137.600 515.600 138.400 ;
        RECT 513.200 133.600 514.000 134.400 ;
        RECT 516.400 129.600 517.200 130.400 ;
        RECT 516.500 128.400 517.100 129.600 ;
        RECT 511.600 127.600 512.400 128.400 ;
        RECT 516.400 127.600 517.200 128.400 ;
        RECT 510.000 123.600 510.800 124.400 ;
        RECT 502.000 117.600 502.800 118.400 ;
        RECT 495.600 110.300 496.400 110.400 ;
        RECT 494.100 109.700 496.400 110.300 ;
        RECT 490.800 97.600 491.600 98.400 ;
        RECT 490.800 89.600 491.600 90.400 ;
        RECT 492.400 90.200 493.200 95.800 ;
        RECT 494.100 94.400 494.700 109.700 ;
        RECT 495.600 109.600 496.400 109.700 ;
        RECT 497.200 104.200 498.000 115.800 ;
        RECT 503.600 106.200 504.400 111.800 ;
        RECT 506.800 104.200 507.600 115.800 ;
        RECT 508.400 109.400 509.200 110.400 ;
        RECT 510.100 108.400 510.700 123.600 ;
        RECT 510.000 107.600 510.800 108.400 ;
        RECT 511.700 100.300 512.300 127.600 ;
        RECT 513.200 117.600 514.000 118.400 ;
        RECT 519.700 118.300 520.300 155.600 ;
        RECT 521.300 152.400 521.900 185.600 ;
        RECT 522.800 175.600 523.600 176.400 ;
        RECT 524.400 175.600 525.200 176.400 ;
        RECT 522.900 172.400 523.500 175.600 ;
        RECT 524.500 174.400 525.100 175.600 ;
        RECT 524.400 173.600 525.200 174.400 ;
        RECT 522.800 171.600 523.600 172.400 ;
        RECT 522.900 152.400 523.500 171.600 ;
        RECT 524.500 162.400 525.100 173.600 ;
        RECT 524.400 161.600 525.200 162.400 ;
        RECT 526.100 156.400 526.700 185.600 ;
        RECT 527.700 170.400 528.300 187.600 ;
        RECT 530.900 178.400 531.500 187.600 ;
        RECT 532.400 185.600 533.200 186.400 ;
        RECT 534.100 182.400 534.700 195.700 ;
        RECT 538.800 191.600 539.600 192.400 ;
        RECT 548.400 191.600 549.200 192.400 ;
        RECT 556.400 191.800 557.200 192.600 ;
        RECT 563.000 191.800 563.800 192.600 ;
        RECT 538.900 190.400 539.500 191.600 ;
        RECT 538.800 189.600 539.600 190.400 ;
        RECT 545.200 189.600 546.000 190.400 ;
        RECT 550.000 189.600 550.800 190.400 ;
        RECT 535.600 187.600 536.400 188.400 ;
        RECT 535.700 186.400 536.300 187.600 ;
        RECT 535.600 185.600 536.400 186.400 ;
        RECT 534.000 181.600 534.800 182.400 ;
        RECT 532.400 179.600 533.200 180.400 ;
        RECT 530.800 177.600 531.600 178.400 ;
        RECT 529.200 175.600 530.000 176.400 ;
        RECT 530.900 174.400 531.500 177.600 ;
        RECT 530.800 173.600 531.600 174.400 ;
        RECT 529.200 171.600 530.000 172.400 ;
        RECT 530.800 171.600 531.600 172.400 ;
        RECT 527.600 169.600 528.400 170.400 ;
        RECT 529.300 168.400 529.900 171.600 ;
        RECT 530.900 170.400 531.500 171.600 ;
        RECT 530.800 169.600 531.600 170.400 ;
        RECT 529.200 167.600 530.000 168.400 ;
        RECT 527.600 165.600 528.400 166.400 ;
        RECT 530.900 158.400 531.500 169.600 ;
        RECT 530.800 157.600 531.600 158.400 ;
        RECT 526.000 155.600 526.800 156.400 ;
        RECT 532.500 154.400 533.100 179.600 ;
        RECT 534.000 175.600 534.800 176.400 ;
        RECT 534.100 174.400 534.700 175.600 ;
        RECT 538.900 174.400 539.500 189.600 ;
        RECT 542.000 187.600 542.800 188.400 ;
        RECT 540.400 183.600 541.200 184.400 ;
        RECT 540.500 180.400 541.100 183.600 ;
        RECT 540.400 179.600 541.200 180.400 ;
        RECT 542.000 175.600 542.800 176.400 ;
        RECT 543.600 175.600 544.400 176.400 ;
        RECT 534.000 173.600 534.800 174.400 ;
        RECT 538.800 173.600 539.600 174.400 ;
        RECT 542.100 172.400 542.700 175.600 ;
        RECT 545.300 174.400 545.900 189.600 ;
        RECT 548.400 187.600 549.200 188.400 ;
        RECT 543.600 173.600 544.400 174.400 ;
        RECT 545.200 173.600 546.000 174.400 ;
        RECT 538.800 171.600 539.600 172.400 ;
        RECT 542.000 171.600 542.800 172.400 ;
        RECT 537.200 167.600 538.000 168.400 ;
        RECT 537.300 166.400 537.900 167.600 ;
        RECT 538.900 166.400 539.500 171.600 ;
        RECT 540.400 169.600 541.200 170.400 ;
        RECT 537.200 165.600 538.000 166.400 ;
        RECT 538.800 165.600 539.600 166.400 ;
        RECT 535.600 163.600 536.400 164.400 ;
        RECT 540.500 162.400 541.100 169.600 ;
        RECT 537.200 161.600 538.000 162.400 ;
        RECT 540.400 161.600 541.200 162.400 ;
        RECT 534.000 157.600 534.800 158.400 ;
        RECT 532.400 153.600 533.200 154.400 ;
        RECT 521.200 151.600 522.000 152.400 ;
        RECT 522.800 151.600 523.600 152.400 ;
        RECT 524.400 151.600 525.200 152.400 ;
        RECT 527.600 151.600 528.400 152.400 ;
        RECT 530.800 151.600 531.600 152.400 ;
        RECT 524.500 150.400 525.100 151.600 ;
        RECT 527.700 150.400 528.300 151.600 ;
        RECT 534.100 150.400 534.700 157.600 ;
        RECT 524.400 149.600 525.200 150.400 ;
        RECT 527.600 149.600 528.400 150.400 ;
        RECT 529.200 149.600 530.000 150.400 ;
        RECT 534.000 149.600 534.800 150.400 ;
        RECT 535.600 149.600 536.400 150.400 ;
        RECT 526.000 147.600 526.800 148.400 ;
        RECT 534.000 147.600 534.800 148.400 ;
        RECT 532.400 145.600 533.200 146.400 ;
        RECT 524.400 143.600 525.200 144.400 ;
        RECT 522.800 141.600 523.600 142.400 ;
        RECT 521.200 137.600 522.000 138.400 ;
        RECT 522.900 134.400 523.500 141.600 ;
        RECT 522.800 133.600 523.600 134.400 ;
        RECT 521.200 118.300 522.000 118.400 ;
        RECT 519.700 117.700 522.000 118.300 ;
        RECT 521.200 117.600 522.000 117.700 ;
        RECT 510.100 99.700 512.300 100.300 ;
        RECT 510.100 98.400 510.700 99.700 ;
        RECT 494.000 93.600 494.800 94.400 ;
        RECT 490.900 88.300 491.500 89.600 ;
        RECT 490.900 87.700 493.100 88.300 ;
        RECT 487.600 85.600 488.400 86.400 ;
        RECT 487.700 70.400 488.300 85.600 ;
        RECT 492.500 70.400 493.100 87.700 ;
        RECT 495.600 86.200 496.400 97.800 ;
        RECT 497.200 91.800 498.000 92.600 ;
        RECT 497.300 88.400 497.900 91.800 ;
        RECT 503.600 91.600 504.400 92.400 ;
        RECT 497.200 87.600 498.000 88.400 ;
        RECT 505.200 86.200 506.000 97.800 ;
        RECT 510.000 97.600 510.800 98.400 ;
        RECT 511.600 98.300 512.400 98.400 ;
        RECT 513.300 98.300 513.900 117.600 ;
        RECT 516.400 104.200 517.200 115.800 ;
        RECT 518.000 113.600 518.800 114.400 ;
        RECT 524.500 114.300 525.100 143.600 ;
        RECT 534.100 138.400 534.700 147.600 ;
        RECT 535.700 146.400 536.300 149.600 ;
        RECT 535.600 145.600 536.400 146.400 ;
        RECT 534.000 137.600 534.800 138.400 ;
        RECT 527.600 133.600 528.400 134.400 ;
        RECT 532.400 133.600 533.200 134.400 ;
        RECT 526.000 129.600 526.800 130.400 ;
        RECT 522.900 113.700 525.100 114.300 ;
        RECT 511.600 97.700 513.900 98.300 ;
        RECT 511.600 97.600 512.400 97.700 ;
        RECT 516.400 86.200 517.200 97.800 ;
        RECT 518.100 92.400 518.700 113.600 ;
        RECT 522.900 108.400 523.500 113.700 ;
        RECT 524.200 111.800 525.000 112.600 ;
        RECT 522.800 107.600 523.600 108.400 ;
        RECT 524.200 107.000 524.800 111.800 ;
        RECT 527.700 110.400 528.300 133.600 ;
        RECT 537.300 130.400 537.900 161.600 ;
        RECT 538.800 153.600 539.600 154.400 ;
        RECT 542.000 151.600 542.800 152.400 ;
        RECT 540.400 149.600 541.200 150.400 ;
        RECT 540.400 147.600 541.200 148.400 ;
        RECT 542.100 146.400 542.700 151.600 ;
        RECT 543.700 150.400 544.300 173.600 ;
        RECT 550.100 172.400 550.700 189.600 ;
        RECT 556.400 188.400 557.000 191.800 ;
        RECT 558.000 189.600 558.800 190.400 ;
        RECT 560.400 188.400 561.200 188.600 ;
        RECT 556.400 187.800 561.200 188.400 ;
        RECT 556.400 187.000 557.000 187.800 ;
        RECT 557.800 187.000 558.600 187.200 ;
        RECT 561.200 187.000 562.000 187.200 ;
        RECT 563.200 187.000 563.800 191.800 ;
        RECT 564.400 187.600 565.200 188.400 ;
        RECT 553.200 185.600 554.000 186.400 ;
        RECT 556.400 186.200 557.200 187.000 ;
        RECT 557.800 186.400 562.000 187.000 ;
        RECT 563.000 186.200 563.800 187.000 ;
        RECT 566.000 186.200 566.800 191.800 ;
        RECT 567.700 188.400 568.300 213.600 ;
        RECT 569.200 211.600 570.000 212.400 ;
        RECT 569.300 208.400 569.900 211.600 ;
        RECT 569.200 207.600 570.000 208.400 ;
        RECT 575.600 206.200 576.400 217.800 ;
        RECT 582.000 211.600 582.800 212.400 ;
        RECT 580.400 208.300 581.200 208.400 ;
        RECT 582.100 208.300 582.700 211.600 ;
        RECT 580.400 207.700 582.700 208.300 ;
        RECT 580.400 207.600 581.200 207.700 ;
        RECT 567.600 187.600 568.400 188.400 ;
        RECT 553.300 176.400 553.900 185.600 ;
        RECT 559.600 183.600 560.400 184.400 ;
        RECT 556.400 177.600 557.200 178.400 ;
        RECT 556.500 176.400 557.100 177.600 ;
        RECT 553.200 175.600 554.000 176.400 ;
        RECT 556.400 175.600 557.200 176.400 ;
        RECT 545.200 171.600 546.000 172.400 ;
        RECT 548.400 171.600 549.200 172.400 ;
        RECT 550.000 171.600 550.800 172.400 ;
        RECT 553.200 171.600 554.000 172.400 ;
        RECT 545.300 166.400 545.900 171.600 ;
        RECT 546.800 169.600 547.600 170.400 ;
        RECT 545.200 165.600 546.000 166.400 ;
        RECT 543.600 149.600 544.400 150.400 ;
        RECT 545.300 150.300 545.900 165.600 ;
        RECT 546.800 163.600 547.600 164.400 ;
        RECT 546.900 152.400 547.500 163.600 ;
        RECT 548.500 158.400 549.100 171.600 ;
        RECT 550.000 167.600 550.800 168.400 ;
        RECT 551.600 163.600 552.400 164.400 ;
        RECT 553.300 162.400 553.900 171.600 ;
        RECT 558.000 170.200 558.800 175.800 ;
        RECT 553.200 161.600 554.000 162.400 ;
        RECT 551.600 159.600 552.400 160.400 ;
        RECT 548.400 157.600 549.200 158.400 ;
        RECT 546.800 151.600 547.600 152.400 ;
        RECT 545.300 149.700 547.500 150.300 ;
        RECT 543.600 147.600 544.400 148.400 ;
        RECT 540.400 145.600 541.200 146.400 ;
        RECT 542.000 145.600 542.800 146.400 ;
        RECT 540.500 138.400 541.100 145.600 ;
        RECT 545.200 143.600 546.000 144.400 ;
        RECT 540.400 137.600 541.200 138.400 ;
        RECT 538.800 135.600 539.600 136.400 ;
        RECT 538.900 134.400 539.500 135.600 ;
        RECT 538.800 133.600 539.600 134.400 ;
        RECT 543.600 133.600 544.400 134.400 ;
        RECT 535.600 129.600 536.400 130.400 ;
        RECT 537.200 129.600 538.000 130.400 ;
        RECT 538.900 128.400 539.500 133.600 ;
        RECT 540.400 129.600 541.200 130.400 ;
        RECT 543.600 129.600 544.400 130.400 ;
        RECT 538.800 127.600 539.600 128.400 ;
        RECT 540.500 124.400 541.100 129.600 ;
        RECT 529.200 123.600 530.000 124.400 ;
        RECT 532.400 123.600 533.200 124.400 ;
        RECT 540.400 123.600 541.200 124.400 ;
        RECT 529.300 112.400 529.900 123.600 ;
        RECT 529.200 111.600 530.000 112.400 ;
        RECT 530.800 111.800 531.600 112.600 ;
        RECT 527.600 109.600 528.400 110.400 ;
        RECT 526.800 108.400 527.600 108.600 ;
        RECT 531.000 108.400 531.600 111.800 ;
        RECT 532.500 108.400 533.100 123.600 ;
        RECT 545.300 114.400 545.900 143.600 ;
        RECT 534.000 113.600 534.800 114.400 ;
        RECT 545.200 113.600 546.000 114.400 ;
        RECT 534.100 108.400 534.700 113.600 ;
        RECT 535.400 111.800 536.200 112.600 ;
        RECT 542.000 111.800 542.800 112.600 ;
        RECT 526.800 107.800 531.600 108.400 ;
        RECT 526.000 107.000 526.800 107.200 ;
        RECT 529.400 107.000 530.200 107.200 ;
        RECT 531.000 107.000 531.600 107.800 ;
        RECT 532.400 107.600 533.200 108.400 ;
        RECT 534.000 107.600 534.800 108.400 ;
        RECT 524.200 106.200 525.000 107.000 ;
        RECT 526.000 106.400 530.200 107.000 ;
        RECT 530.800 106.200 531.600 107.000 ;
        RECT 535.400 107.000 536.000 111.800 ;
        RECT 538.000 108.400 538.800 108.600 ;
        RECT 542.200 108.400 542.800 111.800 ;
        RECT 538.000 107.800 542.800 108.400 ;
        RECT 537.200 107.000 538.000 107.200 ;
        RECT 540.600 107.000 541.400 107.200 ;
        RECT 542.200 107.000 542.800 107.800 ;
        RECT 543.600 107.600 544.400 108.400 ;
        RECT 535.400 106.200 536.200 107.000 ;
        RECT 537.200 106.400 541.400 107.000 ;
        RECT 542.000 106.200 542.800 107.000 ;
        RECT 545.200 106.200 546.000 111.800 ;
        RECT 546.900 108.400 547.500 149.700 ;
        RECT 548.400 149.600 549.200 150.400 ;
        RECT 548.500 142.400 549.100 149.600 ;
        RECT 551.700 148.400 552.300 159.600 ;
        RECT 551.600 147.600 552.400 148.400 ;
        RECT 551.600 145.600 552.400 146.400 ;
        RECT 553.300 142.400 553.900 161.600 ;
        RECT 559.700 158.400 560.300 183.600 ;
        RECT 566.000 181.600 566.800 182.400 ;
        RECT 561.200 166.200 562.000 177.800 ;
        RECT 566.100 172.400 566.700 181.600 ;
        RECT 566.000 171.600 566.800 172.400 ;
        RECT 567.700 172.300 568.300 187.600 ;
        RECT 569.200 184.200 570.000 195.800 ;
        RECT 570.800 189.400 571.600 190.400 ;
        RECT 578.800 184.200 579.600 195.800 ;
        RECT 583.600 183.600 584.400 184.400 ;
        RECT 583.700 182.400 584.300 183.600 ;
        RECT 583.600 181.600 584.400 182.400 ;
        RECT 569.200 172.300 570.000 172.400 ;
        RECT 567.700 171.700 570.000 172.300 ;
        RECT 569.200 171.600 570.000 171.700 ;
        RECT 559.600 157.600 560.400 158.400 ;
        RECT 554.600 151.800 555.400 152.600 ;
        RECT 561.200 151.800 562.000 152.600 ;
        RECT 554.600 147.000 555.200 151.800 ;
        RECT 557.200 148.400 558.000 148.600 ;
        RECT 561.400 148.400 562.000 151.800 ;
        RECT 557.200 147.800 562.000 148.400 ;
        RECT 556.400 147.000 557.200 147.200 ;
        RECT 559.800 147.000 560.600 147.200 ;
        RECT 561.400 147.000 562.000 147.800 ;
        RECT 562.800 147.600 563.600 148.400 ;
        RECT 554.600 146.200 555.400 147.000 ;
        RECT 556.400 146.400 560.600 147.000 ;
        RECT 561.200 146.200 562.000 147.000 ;
        RECT 564.400 146.200 565.200 151.800 ;
        RECT 567.600 144.200 568.400 155.800 ;
        RECT 569.300 148.400 569.900 171.600 ;
        RECT 570.800 166.200 571.600 177.800 ;
        RECT 577.200 171.600 578.000 172.400 ;
        RECT 575.600 168.300 576.400 168.400 ;
        RECT 577.300 168.300 577.900 171.600 ;
        RECT 575.600 167.700 577.900 168.300 ;
        RECT 575.600 167.600 576.400 167.700 ;
        RECT 570.800 163.600 571.600 164.400 ;
        RECT 570.900 150.400 571.500 163.600 ;
        RECT 570.800 149.600 571.600 150.400 ;
        RECT 569.200 147.600 570.000 148.400 ;
        RECT 570.800 147.600 571.600 148.400 ;
        RECT 548.400 141.600 549.200 142.400 ;
        RECT 553.200 141.600 554.000 142.400 ;
        RECT 566.000 139.600 566.800 140.400 ;
        RECT 556.400 137.600 557.200 138.400 ;
        RECT 550.000 135.600 550.800 136.400 ;
        RECT 550.100 134.400 550.700 135.600 ;
        RECT 556.500 134.400 557.100 137.600 ;
        RECT 558.000 135.000 558.800 135.800 ;
        RECT 564.200 135.600 565.000 135.800 ;
        RECT 559.400 135.000 565.000 135.600 ;
        RECT 548.400 133.600 549.200 134.400 ;
        RECT 550.000 133.600 550.800 134.400 ;
        RECT 556.400 133.600 557.200 134.400 ;
        RECT 558.000 134.200 558.600 135.000 ;
        RECT 559.400 134.800 560.200 135.000 ;
        RECT 562.800 134.800 563.600 135.000 ;
        RECT 558.000 133.600 563.600 134.200 ;
        RECT 548.500 124.400 549.100 133.600 ;
        RECT 558.000 130.200 558.600 133.600 ;
        RECT 563.000 132.200 563.600 133.600 ;
        RECT 563.000 131.400 563.800 132.200 ;
        RECT 564.400 130.200 565.000 135.000 ;
        RECT 566.100 134.400 566.700 139.600 ;
        RECT 570.900 138.400 571.500 147.600 ;
        RECT 577.200 144.200 578.000 155.800 ;
        RECT 583.600 143.600 584.400 144.400 ;
        RECT 570.800 137.600 571.600 138.400 ;
        RECT 569.200 135.000 570.000 135.800 ;
        RECT 575.400 135.600 576.200 135.800 ;
        RECT 577.200 135.600 578.000 136.400 ;
        RECT 570.600 135.000 576.200 135.600 ;
        RECT 566.000 133.600 566.800 134.400 ;
        RECT 567.600 133.600 568.400 134.400 ;
        RECT 569.200 134.200 569.800 135.000 ;
        RECT 570.600 134.800 571.400 135.000 ;
        RECT 574.000 134.800 574.800 135.000 ;
        RECT 569.200 133.600 574.800 134.200 ;
        RECT 558.000 129.400 558.800 130.200 ;
        RECT 564.200 129.400 565.000 130.200 ;
        RECT 548.400 123.600 549.200 124.400 ;
        RECT 559.600 123.600 560.400 124.400 ;
        RECT 546.800 107.600 547.600 108.400 ;
        RECT 529.200 103.600 530.000 104.400 ;
        RECT 535.600 103.600 536.400 104.400 ;
        RECT 540.400 103.600 541.200 104.400 ;
        RECT 546.800 103.600 547.600 104.400 ;
        RECT 548.400 104.200 549.200 115.800 ;
        RECT 551.600 109.600 552.400 110.400 ;
        RECT 554.800 109.600 555.600 110.400 ;
        RECT 554.900 108.400 555.500 109.600 ;
        RECT 550.000 107.600 550.800 108.400 ;
        RECT 554.800 107.600 555.600 108.400 ;
        RECT 529.300 102.400 529.900 103.600 ;
        RECT 529.200 101.600 530.000 102.400 ;
        RECT 518.000 91.600 518.800 92.400 ;
        RECT 524.400 91.800 525.200 92.600 ;
        RECT 524.500 88.400 525.100 91.800 ;
        RECT 524.400 87.600 525.200 88.400 ;
        RECT 526.000 86.200 526.800 97.800 ;
        RECT 529.200 90.200 530.000 95.800 ;
        RECT 530.800 90.200 531.600 95.800 ;
        RECT 529.200 87.600 530.000 88.400 ;
        RECT 503.600 83.600 504.400 84.400 ;
        RECT 494.000 73.600 494.800 74.400 ;
        RECT 494.100 72.400 494.700 73.600 ;
        RECT 494.000 71.600 494.800 72.400 ;
        RECT 503.700 70.400 504.300 83.600 ;
        RECT 529.300 78.400 529.900 87.600 ;
        RECT 534.000 86.200 534.800 97.800 ;
        RECT 529.200 77.600 530.000 78.400 ;
        RECT 518.000 73.600 518.800 74.400 ;
        RECT 532.400 73.600 533.200 74.400 ;
        RECT 518.100 72.300 518.700 73.600 ;
        RECT 532.500 72.400 533.100 73.600 ;
        RECT 518.100 71.700 520.300 72.300 ;
        RECT 519.700 70.400 520.300 71.700 ;
        RECT 524.400 71.600 525.200 72.400 ;
        RECT 532.400 71.600 533.200 72.400 ;
        RECT 535.700 70.400 536.300 103.600 ;
        RECT 537.200 101.600 538.000 102.400 ;
        RECT 537.300 92.400 537.900 101.600 ;
        RECT 542.000 93.600 542.800 94.400 ;
        RECT 537.200 91.600 538.000 92.400 ;
        RECT 543.600 86.200 544.400 97.800 ;
        RECT 484.400 69.700 486.700 70.300 ;
        RECT 484.400 69.600 485.200 69.700 ;
        RECT 484.400 67.600 485.200 68.400 ;
        RECT 476.400 65.600 477.200 66.400 ;
        RECT 478.000 65.600 478.800 66.400 ;
        RECT 479.600 65.600 480.400 66.400 ;
        RECT 484.400 65.600 485.200 66.400 ;
        RECT 473.200 61.600 474.000 62.400 ;
        RECT 460.400 57.600 461.200 58.400 ;
        RECT 460.500 54.400 461.100 57.600 ;
        RECT 476.500 56.400 477.100 65.600 ;
        RECT 478.000 61.600 478.800 62.400 ;
        RECT 478.100 56.400 478.700 61.600 ;
        RECT 479.700 58.400 480.300 65.600 ;
        RECT 479.600 57.600 480.400 58.400 ;
        RECT 486.100 58.300 486.700 69.700 ;
        RECT 487.600 69.600 488.400 70.400 ;
        RECT 490.800 69.600 491.600 70.400 ;
        RECT 492.400 69.600 493.200 70.400 ;
        RECT 497.200 69.600 498.000 70.400 ;
        RECT 503.600 69.600 504.400 70.400 ;
        RECT 506.800 69.600 507.600 70.400 ;
        RECT 510.000 69.600 510.800 70.400 ;
        RECT 518.000 69.600 518.800 70.400 ;
        RECT 519.600 69.600 520.400 70.400 ;
        RECT 529.200 69.600 530.000 70.400 ;
        RECT 535.600 69.600 536.400 70.400 ;
        RECT 490.900 58.400 491.500 69.600 ;
        RECT 492.400 68.300 493.200 68.400 ;
        RECT 492.400 67.700 494.700 68.300 ;
        RECT 492.400 67.600 493.200 67.700 ;
        RECT 492.400 63.600 493.200 64.400 ;
        RECT 492.500 58.400 493.100 63.600 ;
        RECT 484.500 57.700 486.700 58.300 ;
        RECT 470.000 55.600 470.800 56.400 ;
        RECT 476.400 55.600 477.200 56.400 ;
        RECT 478.000 55.600 478.800 56.400 ;
        RECT 470.100 54.400 470.700 55.600 ;
        RECT 458.800 53.600 459.600 54.400 ;
        RECT 460.400 53.600 461.200 54.400 ;
        RECT 463.600 53.600 464.400 54.400 ;
        RECT 468.400 53.600 469.200 54.400 ;
        RECT 470.000 53.600 470.800 54.400 ;
        RECT 471.600 53.600 472.400 54.400 ;
        RECT 468.500 52.400 469.100 53.600 ;
        RECT 471.700 52.400 472.300 53.600 ;
        RECT 457.200 51.600 458.000 52.400 ;
        RECT 468.400 51.600 469.200 52.400 ;
        RECT 471.600 51.600 472.400 52.400 ;
        RECT 457.300 50.400 457.900 51.600 ;
        RECT 476.500 50.400 477.100 55.600 ;
        RECT 481.200 51.600 482.000 52.400 ;
        RECT 452.400 49.600 453.200 50.400 ;
        RECT 457.200 49.600 458.000 50.400 ;
        RECT 463.600 49.600 464.400 50.400 ;
        RECT 465.200 49.600 466.000 50.400 ;
        RECT 468.400 49.600 469.200 50.400 ;
        RECT 476.400 49.600 477.200 50.400 ;
        RECT 463.700 48.400 464.300 49.600 ;
        RECT 452.400 48.300 453.200 48.400 ;
        RECT 450.900 47.700 453.200 48.300 ;
        RECT 452.400 47.600 453.200 47.700 ;
        RECT 463.600 47.600 464.400 48.400 ;
        RECT 447.600 45.600 448.400 46.400 ;
        RECT 452.500 32.400 453.100 47.600 ;
        RECT 458.800 37.600 459.600 38.400 ;
        RECT 455.600 33.600 456.400 34.400 ;
        RECT 458.900 32.400 459.500 37.600 ;
        RECT 460.400 35.600 461.200 36.400 ;
        RECT 442.800 32.300 443.600 32.400 ;
        RECT 441.300 31.700 443.600 32.300 ;
        RECT 431.700 29.700 435.500 30.300 ;
        RECT 431.700 28.400 432.300 29.700 ;
        RECT 431.600 27.600 432.400 28.400 ;
        RECT 433.200 27.600 434.000 28.400 ;
        RECT 433.200 25.600 434.000 26.400 ;
        RECT 434.900 26.300 435.500 29.700 ;
        RECT 439.600 29.600 440.400 30.400 ;
        RECT 439.700 28.400 440.300 29.600 ;
        RECT 438.000 27.600 438.800 28.400 ;
        RECT 439.600 27.600 440.400 28.400 ;
        RECT 441.300 26.300 441.900 31.700 ;
        RECT 442.800 31.600 443.600 31.700 ;
        RECT 447.600 31.600 448.400 32.400 ;
        RECT 449.200 31.600 450.000 32.400 ;
        RECT 452.400 31.600 453.200 32.400 ;
        RECT 457.200 31.600 458.000 32.400 ;
        RECT 458.800 31.600 459.600 32.400 ;
        RECT 444.400 27.600 445.200 28.400 ;
        RECT 434.900 25.700 441.900 26.300 ;
        RECT 433.300 20.400 433.900 25.600 ;
        RECT 444.500 20.400 445.100 27.600 ;
        RECT 433.200 19.600 434.000 20.400 ;
        RECT 434.800 19.600 435.600 20.400 ;
        RECT 438.000 19.600 438.800 20.400 ;
        RECT 441.200 19.600 442.000 20.400 ;
        RECT 444.400 19.600 445.200 20.400 ;
        RECT 428.500 15.700 430.700 16.300 ;
        RECT 428.500 14.400 429.100 15.700 ;
        RECT 433.200 15.600 434.000 16.400 ;
        RECT 428.400 13.600 429.200 14.400 ;
        RECT 430.000 13.600 430.800 14.400 ;
        RECT 426.800 12.300 427.600 12.400 ;
        RECT 425.300 11.700 427.600 12.300 ;
        RECT 426.800 11.600 427.600 11.700 ;
        RECT 433.300 10.400 433.900 15.600 ;
        RECT 434.900 12.400 435.500 19.600 ;
        RECT 438.100 18.400 438.700 19.600 ;
        RECT 438.000 17.600 438.800 18.400 ;
        RECT 441.300 16.400 441.900 19.600 ;
        RECT 441.200 15.600 442.000 16.400 ;
        RECT 447.700 14.400 448.300 31.600 ;
        RECT 449.300 30.400 449.900 31.600 ;
        RECT 449.200 29.600 450.000 30.400 ;
        RECT 457.300 22.400 457.900 31.600 ;
        RECT 452.400 21.600 453.200 22.400 ;
        RECT 457.200 22.300 458.000 22.400 ;
        RECT 457.200 21.700 459.500 22.300 ;
        RECT 457.200 21.600 458.000 21.700 ;
        RECT 452.500 18.400 453.100 21.600 ;
        RECT 455.600 19.600 456.400 20.400 ;
        RECT 455.700 18.400 456.300 19.600 ;
        RECT 452.400 17.600 453.200 18.400 ;
        RECT 455.600 17.600 456.400 18.400 ;
        RECT 458.900 16.400 459.500 21.700 ;
        RECT 460.500 18.400 461.100 35.600 ;
        RECT 465.200 33.600 466.000 34.400 ;
        RECT 465.300 32.400 465.900 33.600 ;
        RECT 462.000 32.300 462.800 32.400 ;
        RECT 462.000 31.700 464.300 32.300 ;
        RECT 462.000 31.600 462.800 31.700 ;
        RECT 462.000 29.600 462.800 30.400 ;
        RECT 462.100 28.400 462.700 29.600 ;
        RECT 463.700 28.400 464.300 31.700 ;
        RECT 465.200 31.600 466.000 32.400 ;
        RECT 468.500 30.400 469.100 49.600 ;
        RECT 484.500 48.400 485.100 57.700 ;
        RECT 489.200 57.600 490.000 58.400 ;
        RECT 490.800 57.600 491.600 58.400 ;
        RECT 492.400 57.600 493.200 58.400 ;
        RECT 486.000 55.600 486.800 56.400 ;
        RECT 486.000 53.600 486.800 54.400 ;
        RECT 487.600 53.600 488.400 54.400 ;
        RECT 486.100 52.400 486.700 53.600 ;
        RECT 487.700 52.400 488.300 53.600 ;
        RECT 489.300 52.400 489.900 57.600 ;
        RECT 494.100 56.400 494.700 67.700 ;
        RECT 498.800 67.600 499.600 68.400 ;
        RECT 505.200 67.600 506.000 68.400 ;
        RECT 497.200 65.600 498.000 66.400 ;
        RECT 498.800 65.600 499.600 66.400 ;
        RECT 500.400 65.600 501.200 66.400 ;
        RECT 495.600 57.600 496.400 58.400 ;
        RECT 494.000 55.600 494.800 56.400 ;
        RECT 494.100 54.400 494.700 55.600 ;
        RECT 494.000 53.600 494.800 54.400 ;
        RECT 486.000 51.600 486.800 52.400 ;
        RECT 487.600 51.600 488.400 52.400 ;
        RECT 489.200 51.600 490.000 52.400 ;
        RECT 492.400 50.300 493.200 50.400 ;
        RECT 490.900 49.700 493.200 50.300 ;
        RECT 484.400 47.600 485.200 48.400 ;
        RECT 470.000 43.600 470.800 44.400 ;
        RECT 476.400 43.600 477.200 44.400 ;
        RECT 470.100 32.300 470.700 43.600 ;
        RECT 471.600 39.600 472.400 40.400 ;
        RECT 471.700 38.400 472.300 39.600 ;
        RECT 476.500 38.400 477.100 43.600 ;
        RECT 471.600 37.600 472.400 38.400 ;
        RECT 476.400 37.600 477.200 38.400 ;
        RECT 479.600 37.600 480.400 38.400 ;
        RECT 470.100 31.700 472.300 32.300 ;
        RECT 468.400 29.600 469.200 30.400 ;
        RECT 470.000 29.600 470.800 30.400 ;
        RECT 468.500 28.400 469.100 29.600 ;
        RECT 471.700 28.400 472.300 31.700 ;
        RECT 476.400 29.600 477.200 30.400 ;
        RECT 478.000 29.600 478.800 30.400 ;
        RECT 462.000 27.600 462.800 28.400 ;
        RECT 463.600 27.600 464.400 28.400 ;
        RECT 468.400 27.600 469.200 28.400 ;
        RECT 471.600 27.600 472.400 28.400 ;
        RECT 474.800 27.600 475.600 28.400 ;
        RECT 466.800 23.600 467.600 24.400 ;
        RECT 463.600 21.600 464.400 22.400 ;
        RECT 460.400 17.600 461.200 18.400 ;
        RECT 457.200 15.600 458.000 16.400 ;
        RECT 458.800 15.600 459.600 16.400 ;
        RECT 462.000 15.600 462.800 16.400 ;
        RECT 457.300 14.400 457.900 15.600 ;
        RECT 446.000 13.600 446.800 14.400 ;
        RECT 447.600 13.600 448.400 14.400 ;
        RECT 452.400 13.600 453.200 14.400 ;
        RECT 457.200 13.600 458.000 14.400 ;
        RECT 434.800 11.600 435.600 12.400 ;
        RECT 452.500 10.400 453.100 13.600 ;
        RECT 462.100 10.400 462.700 15.600 ;
        RECT 463.700 14.400 464.300 21.600 ;
        RECT 466.900 16.400 467.500 23.600 ;
        RECT 474.900 20.400 475.500 27.600 ;
        RECT 476.500 26.400 477.100 29.600 ;
        RECT 476.400 25.600 477.200 26.400 ;
        RECT 478.100 24.400 478.700 29.600 ;
        RECT 479.700 28.400 480.300 37.600 ;
        RECT 484.500 30.400 485.100 47.600 ;
        RECT 486.000 37.600 486.800 38.400 ;
        RECT 487.600 37.600 488.400 38.400 ;
        RECT 486.100 30.400 486.700 37.600 ;
        RECT 487.600 35.600 488.400 36.400 ;
        RECT 489.200 35.600 490.000 36.400 ;
        RECT 484.400 29.600 485.200 30.400 ;
        RECT 486.000 29.600 486.800 30.400 ;
        RECT 479.600 27.600 480.400 28.400 ;
        RECT 482.800 27.600 483.600 28.400 ;
        RECT 478.000 23.600 478.800 24.400 ;
        RECT 481.200 23.600 482.000 24.400 ;
        RECT 481.200 21.600 482.000 22.400 ;
        RECT 474.800 19.600 475.600 20.400 ;
        RECT 466.800 15.600 467.600 16.400 ;
        RECT 468.400 15.600 469.200 16.400 ;
        RECT 471.400 15.000 472.200 15.800 ;
        RECT 473.200 15.000 477.400 15.600 ;
        RECT 478.000 15.000 478.800 15.800 ;
        RECT 463.600 13.600 464.400 14.400 ;
        RECT 470.000 13.600 470.800 14.400 ;
        RECT 465.200 11.600 466.000 12.400 ;
        RECT 404.400 9.400 405.200 10.200 ;
        RECT 410.600 9.400 411.400 10.200 ;
        RECT 412.400 9.600 413.200 10.400 ;
        RECT 422.000 9.600 422.800 10.400 ;
        RECT 433.200 9.600 434.000 10.400 ;
        RECT 452.400 9.600 453.200 10.400 ;
        RECT 462.000 9.600 462.800 10.400 ;
        RECT 468.400 10.300 469.200 10.400 ;
        RECT 470.100 10.300 470.700 13.600 ;
        RECT 468.400 9.700 470.700 10.300 ;
        RECT 471.400 10.200 472.000 15.000 ;
        RECT 473.200 14.800 474.000 15.000 ;
        RECT 476.600 14.800 477.400 15.000 ;
        RECT 478.200 14.200 478.800 15.000 ;
        RECT 481.300 14.400 481.900 21.600 ;
        RECT 482.900 20.400 483.500 27.600 ;
        RECT 482.800 19.600 483.600 20.400 ;
        RECT 474.000 13.600 478.800 14.200 ;
        RECT 481.200 13.600 482.000 14.400 ;
        RECT 474.000 13.400 474.800 13.600 ;
        RECT 468.400 9.600 469.200 9.700 ;
        RECT 471.400 9.400 472.200 10.200 ;
        RECT 476.400 9.600 477.200 10.400 ;
        RECT 478.200 10.200 478.800 13.600 ;
        RECT 479.600 11.600 480.400 12.400 ;
        RECT 478.000 9.400 478.800 10.200 ;
        RECT 484.500 10.300 485.100 29.600 ;
        RECT 486.000 28.300 486.800 28.400 ;
        RECT 487.700 28.300 488.300 35.600 ;
        RECT 486.000 27.700 488.300 28.300 ;
        RECT 486.000 27.600 486.800 27.700 ;
        RECT 489.300 14.400 489.900 35.600 ;
        RECT 490.900 32.400 491.500 49.700 ;
        RECT 492.400 49.600 493.200 49.700 ;
        RECT 494.000 39.600 494.800 40.400 ;
        RECT 490.800 31.600 491.600 32.400 ;
        RECT 492.400 31.600 493.200 32.400 ;
        RECT 490.800 23.600 491.600 24.400 ;
        RECT 489.200 13.600 490.000 14.400 ;
        RECT 490.900 12.400 491.500 23.600 ;
        RECT 492.500 16.400 493.100 31.600 ;
        RECT 494.100 30.300 494.700 39.600 ;
        RECT 495.700 38.400 496.300 57.600 ;
        RECT 497.300 56.400 497.900 65.600 ;
        RECT 498.900 58.400 499.500 65.600 ;
        RECT 500.500 64.400 501.100 65.600 ;
        RECT 500.400 63.600 501.200 64.400 ;
        RECT 503.600 63.600 504.400 64.400 ;
        RECT 498.800 57.600 499.600 58.400 ;
        RECT 503.700 56.400 504.300 63.600 ;
        RECT 505.300 58.400 505.900 67.600 ;
        RECT 505.200 57.600 506.000 58.400 ;
        RECT 497.200 55.600 498.000 56.400 ;
        RECT 503.600 55.600 504.400 56.400 ;
        RECT 497.200 53.600 498.000 54.400 ;
        RECT 500.400 53.600 501.200 54.400 ;
        RECT 502.000 51.600 502.800 52.400 ;
        RECT 502.100 48.400 502.700 51.600 ;
        RECT 503.600 49.600 504.400 50.400 ;
        RECT 502.000 47.600 502.800 48.400 ;
        RECT 495.600 37.600 496.400 38.400 ;
        RECT 498.800 37.600 499.600 38.400 ;
        RECT 498.900 32.400 499.500 37.600 ;
        RECT 498.800 31.600 499.600 32.400 ;
        RECT 502.000 31.600 502.800 32.400 ;
        RECT 502.100 30.400 502.700 31.600 ;
        RECT 495.600 30.300 496.400 30.400 ;
        RECT 494.100 29.700 496.400 30.300 ;
        RECT 495.600 29.600 496.400 29.700 ;
        RECT 502.000 29.600 502.800 30.400 ;
        RECT 503.700 28.400 504.300 49.600 ;
        RECT 506.900 40.400 507.500 69.600 ;
        RECT 510.100 68.400 510.700 69.600 ;
        RECT 508.400 67.600 509.200 68.400 ;
        RECT 510.000 67.600 510.800 68.400 ;
        RECT 514.800 67.600 515.600 68.400 ;
        RECT 519.600 67.600 520.400 68.400 ;
        RECT 508.500 56.400 509.100 67.600 ;
        RECT 529.300 66.400 529.900 69.600 ;
        RECT 530.800 67.600 531.600 68.400 ;
        RECT 540.400 67.600 541.200 68.400 ;
        RECT 510.000 65.600 510.800 66.400 ;
        RECT 513.200 65.600 514.000 66.400 ;
        RECT 514.800 65.600 515.600 66.400 ;
        RECT 519.600 65.600 520.400 66.400 ;
        RECT 529.200 65.600 530.000 66.400 ;
        RECT 542.000 66.200 542.800 71.800 ;
        RECT 510.100 58.400 510.700 65.600 ;
        RECT 510.000 57.600 510.800 58.400 ;
        RECT 508.400 55.600 509.200 56.400 ;
        RECT 511.600 56.300 512.400 56.400 ;
        RECT 513.300 56.300 513.900 65.600 ;
        RECT 519.700 58.400 520.300 65.600 ;
        RECT 542.000 63.600 542.800 64.400 ;
        RECT 545.200 64.200 546.000 75.800 ;
        RECT 546.900 70.200 547.500 103.600 ;
        RECT 550.100 98.400 550.700 107.600 ;
        RECT 550.000 97.600 550.800 98.400 ;
        RECT 551.600 93.600 552.400 94.400 ;
        RECT 548.400 87.600 549.200 88.400 ;
        RECT 546.800 69.400 547.600 70.200 ;
        RECT 550.000 67.600 550.800 68.400 ;
        RECT 542.100 58.400 542.700 63.600 ;
        RECT 519.600 57.600 520.400 58.400 ;
        RECT 522.800 57.600 523.600 58.400 ;
        RECT 511.600 55.700 513.900 56.300 ;
        RECT 511.600 55.600 512.400 55.700 ;
        RECT 514.800 55.000 515.600 55.800 ;
        RECT 516.200 55.000 520.400 55.600 ;
        RECT 521.400 55.000 522.200 55.800 ;
        RECT 508.400 53.600 509.200 54.400 ;
        RECT 514.800 54.200 515.400 55.000 ;
        RECT 516.200 54.800 517.000 55.000 ;
        RECT 519.600 54.800 520.400 55.000 ;
        RECT 514.800 53.600 519.600 54.200 ;
        RECT 508.500 52.400 509.100 53.600 ;
        RECT 508.400 51.600 509.200 52.400 ;
        RECT 511.600 51.600 512.400 52.400 ;
        RECT 506.800 39.600 507.600 40.400 ;
        RECT 508.500 36.400 509.100 51.600 ;
        RECT 510.000 47.600 510.800 48.400 ;
        RECT 510.100 38.400 510.700 47.600 ;
        RECT 510.000 37.600 510.800 38.400 ;
        RECT 508.400 35.600 509.200 36.400 ;
        RECT 508.400 31.600 509.200 32.400 ;
        RECT 505.200 29.600 506.000 30.400 ;
        RECT 497.200 27.600 498.000 28.400 ;
        RECT 500.400 27.600 501.200 28.400 ;
        RECT 503.600 27.600 504.400 28.400 ;
        RECT 497.300 24.400 497.900 27.600 ;
        RECT 497.200 23.600 498.000 24.400 ;
        RECT 500.500 24.300 501.100 27.600 ;
        RECT 505.300 26.400 505.900 29.600 ;
        RECT 506.800 27.600 507.600 28.400 ;
        RECT 506.900 26.400 507.500 27.600 ;
        RECT 505.200 25.600 506.000 26.400 ;
        RECT 506.800 25.600 507.600 26.400 ;
        RECT 508.500 24.300 509.100 31.600 ;
        RECT 510.000 27.600 510.800 28.400 ;
        RECT 500.500 23.700 509.100 24.300 ;
        RECT 505.200 21.600 506.000 22.400 ;
        RECT 500.400 19.600 501.200 20.400 ;
        RECT 500.500 16.400 501.100 19.600 ;
        RECT 505.300 18.400 505.900 21.600 ;
        RECT 506.800 19.600 507.600 20.400 ;
        RECT 505.200 17.600 506.000 18.400 ;
        RECT 506.900 16.400 507.500 19.600 ;
        RECT 511.700 16.400 512.300 51.600 ;
        RECT 514.800 50.200 515.400 53.600 ;
        RECT 518.800 53.400 519.600 53.600 ;
        RECT 514.800 49.400 515.600 50.200 ;
        RECT 516.400 49.600 517.200 50.400 ;
        RECT 521.600 50.200 522.200 55.000 ;
        RECT 522.900 54.400 523.500 57.600 ;
        RECT 522.800 53.600 523.600 54.400 ;
        RECT 524.400 50.200 525.200 55.800 ;
        RECT 514.800 29.600 515.600 30.400 ;
        RECT 514.800 25.600 515.600 26.400 ;
        RECT 514.900 24.400 515.500 25.600 ;
        RECT 514.800 23.600 515.600 24.400 ;
        RECT 513.200 19.600 514.000 20.400 ;
        RECT 513.300 18.400 513.900 19.600 ;
        RECT 516.500 18.400 517.100 49.600 ;
        RECT 521.400 49.400 522.200 50.200 ;
        RECT 527.600 46.200 528.400 57.800 ;
        RECT 532.400 51.600 533.200 52.400 ;
        RECT 535.600 51.600 536.400 52.400 ;
        RECT 519.600 39.600 520.400 40.400 ;
        RECT 519.700 30.400 520.300 39.600 ;
        RECT 532.500 38.400 533.100 51.600 ;
        RECT 537.200 46.200 538.000 57.800 ;
        RECT 542.000 57.600 542.800 58.400 ;
        RECT 548.400 46.200 549.200 57.800 ;
        RECT 550.100 54.400 550.700 67.600 ;
        RECT 551.700 58.400 552.300 93.600 ;
        RECT 553.200 90.200 554.000 95.800 ;
        RECT 554.900 94.400 555.500 107.600 ;
        RECT 558.000 104.200 558.800 115.800 ;
        RECT 559.700 110.400 560.300 123.600 ;
        RECT 567.700 118.400 568.300 133.600 ;
        RECT 569.200 130.200 569.800 133.600 ;
        RECT 574.200 132.200 574.800 133.600 ;
        RECT 574.200 131.400 575.000 132.200 ;
        RECT 575.600 130.200 576.200 135.000 ;
        RECT 577.300 134.400 577.900 135.600 ;
        RECT 577.200 133.600 578.000 134.400 ;
        RECT 569.200 129.400 570.000 130.200 ;
        RECT 575.400 129.400 576.200 130.200 ;
        RECT 567.600 117.600 568.400 118.400 ;
        RECT 582.000 117.600 582.800 118.400 ;
        RECT 562.800 113.600 563.600 114.400 ;
        RECT 562.900 112.400 563.500 113.600 ;
        RECT 562.800 111.600 563.600 112.400 ;
        RECT 559.600 109.600 560.400 110.400 ;
        RECT 564.400 106.200 565.200 111.800 ;
        RECT 566.000 107.600 566.800 108.400 ;
        RECT 567.600 104.200 568.400 115.800 ;
        RECT 569.200 111.600 570.000 112.400 ;
        RECT 569.300 110.200 569.900 111.600 ;
        RECT 569.200 109.400 570.000 110.200 ;
        RECT 577.200 104.200 578.000 115.800 ;
        RECT 583.700 102.400 584.300 143.600 ;
        RECT 577.200 101.600 578.000 102.400 ;
        RECT 583.600 101.600 584.400 102.400 ;
        RECT 554.800 93.600 555.600 94.400 ;
        RECT 556.400 86.200 557.200 97.800 ;
        RECT 558.000 91.800 558.800 92.600 ;
        RECT 558.100 88.400 558.700 91.800 ;
        RECT 558.000 87.600 558.800 88.400 ;
        RECT 566.000 86.200 566.800 97.800 ;
        RECT 577.300 92.400 577.900 101.600 ;
        RECT 572.400 91.600 573.200 92.400 ;
        RECT 577.200 91.600 578.000 92.400 ;
        RECT 567.600 87.600 568.400 88.400 ;
        RECT 570.800 88.300 571.600 88.400 ;
        RECT 572.500 88.300 573.100 91.600 ;
        RECT 570.800 87.700 573.100 88.300 ;
        RECT 570.800 87.600 571.600 87.700 ;
        RECT 553.200 67.600 554.000 68.400 ;
        RECT 551.600 57.600 552.400 58.400 ;
        RECT 550.000 53.600 550.800 54.400 ;
        RECT 550.100 52.400 550.700 53.600 ;
        RECT 550.000 51.600 550.800 52.400 ;
        RECT 543.600 43.600 544.400 44.400 ;
        RECT 532.400 37.600 533.200 38.400 ;
        RECT 529.200 33.600 530.000 34.400 ;
        RECT 519.600 29.600 520.400 30.400 ;
        RECT 522.800 29.600 523.600 30.400 ;
        RECT 527.600 29.600 528.400 30.400 ;
        RECT 518.000 27.600 518.800 28.400 ;
        RECT 518.100 26.400 518.700 27.600 ;
        RECT 518.000 25.600 518.800 26.400 ;
        RECT 519.600 21.600 520.400 22.400 ;
        RECT 513.200 17.600 514.000 18.400 ;
        RECT 516.400 17.600 517.200 18.400 ;
        RECT 492.400 15.600 493.200 16.400 ;
        RECT 500.400 15.600 501.200 16.400 ;
        RECT 506.800 15.600 507.600 16.400 ;
        RECT 510.000 15.600 510.800 16.400 ;
        RECT 511.600 15.600 512.400 16.400 ;
        RECT 492.400 13.600 493.200 14.400 ;
        RECT 494.000 13.600 494.800 14.400 ;
        RECT 495.600 13.600 496.400 14.400 ;
        RECT 502.000 13.600 502.800 14.400 ;
        RECT 511.600 14.300 512.400 14.400 ;
        RECT 516.400 14.300 517.200 14.400 ;
        RECT 511.600 13.700 517.200 14.300 ;
        RECT 511.600 13.600 512.400 13.700 ;
        RECT 516.400 13.600 517.200 13.700 ;
        RECT 486.000 11.600 486.800 12.400 ;
        RECT 490.800 11.600 491.600 12.400 ;
        RECT 486.100 10.400 486.700 11.600 ;
        RECT 486.000 10.300 486.800 10.400 ;
        RECT 484.500 9.700 486.800 10.300 ;
        RECT 492.500 10.300 493.100 13.600 ;
        RECT 494.100 12.400 494.700 13.600 ;
        RECT 495.700 12.400 496.300 13.600 ;
        RECT 519.700 12.400 520.300 21.600 ;
        RECT 522.900 18.400 523.500 29.600 ;
        RECT 524.400 25.600 525.200 26.400 ;
        RECT 522.800 17.600 523.600 18.400 ;
        RECT 521.200 15.600 522.000 16.400 ;
        RECT 494.000 11.600 494.800 12.400 ;
        RECT 495.600 11.600 496.400 12.400 ;
        RECT 498.800 11.600 499.600 12.400 ;
        RECT 510.000 11.600 510.800 12.400 ;
        RECT 519.600 11.600 520.400 12.400 ;
        RECT 498.900 10.400 499.500 11.600 ;
        RECT 521.300 10.400 521.900 15.600 ;
        RECT 524.500 12.400 525.100 25.600 ;
        RECT 526.000 23.600 526.800 24.400 ;
        RECT 526.100 14.400 526.700 23.600 ;
        RECT 527.700 22.400 528.300 29.600 ;
        RECT 529.300 28.400 529.900 33.600 ;
        RECT 530.800 31.800 531.600 32.600 ;
        RECT 537.400 31.800 538.200 32.600 ;
        RECT 530.800 28.400 531.400 31.800 ;
        RECT 534.800 28.400 535.600 28.600 ;
        RECT 529.200 27.600 530.000 28.400 ;
        RECT 530.800 27.800 535.600 28.400 ;
        RECT 530.800 27.000 531.400 27.800 ;
        RECT 532.200 27.000 533.000 27.200 ;
        RECT 535.600 27.000 536.400 27.200 ;
        RECT 537.600 27.000 538.200 31.800 ;
        RECT 540.400 31.600 541.200 32.400 ;
        RECT 551.600 31.600 552.400 32.400 ;
        RECT 538.800 29.600 539.600 30.400 ;
        RECT 530.800 26.200 531.600 27.000 ;
        RECT 532.200 26.400 536.400 27.000 ;
        RECT 537.400 26.200 538.200 27.000 ;
        RECT 527.600 21.600 528.400 22.400 ;
        RECT 538.900 20.400 539.500 29.600 ;
        RECT 540.500 28.400 541.100 31.600 ;
        RECT 543.600 29.600 544.400 30.400 ;
        RECT 550.000 29.600 550.800 30.400 ;
        RECT 540.400 27.600 541.200 28.400 ;
        RECT 543.700 26.400 544.300 29.600 ;
        RECT 550.100 28.400 550.700 29.600 ;
        RECT 548.400 27.600 549.200 28.400 ;
        RECT 550.000 27.600 550.800 28.400 ;
        RECT 543.600 25.600 544.400 26.400 ;
        RECT 546.800 23.600 547.600 24.400 ;
        RECT 542.000 21.600 542.800 22.400 ;
        RECT 538.800 19.600 539.600 20.400 ;
        RECT 535.600 15.600 536.400 16.400 ;
        RECT 526.000 13.600 526.800 14.400 ;
        RECT 527.600 13.600 528.400 14.400 ;
        RECT 529.200 13.600 530.000 14.400 ;
        RECT 534.000 13.600 534.800 14.400 ;
        RECT 527.700 12.400 528.300 13.600 ;
        RECT 538.900 12.400 539.500 19.600 ;
        RECT 542.100 18.400 542.700 21.600 ;
        RECT 542.000 17.600 542.800 18.400 ;
        RECT 546.900 16.400 547.500 23.600 ;
        RECT 548.500 22.400 549.100 27.600 ;
        RECT 551.700 26.300 552.300 31.600 ;
        RECT 553.300 28.300 553.900 67.600 ;
        RECT 554.800 64.200 555.600 75.800 ;
        RECT 559.600 73.600 560.400 74.400 ;
        RECT 559.700 72.400 560.300 73.600 ;
        RECT 559.600 71.600 560.400 72.400 ;
        RECT 561.200 66.200 562.000 71.800 ;
        RECT 564.400 64.200 565.200 75.800 ;
        RECT 566.000 71.600 566.800 72.400 ;
        RECT 566.100 70.200 566.700 71.600 ;
        RECT 566.000 69.400 566.800 70.200 ;
        RECT 567.700 68.400 568.300 87.600 ;
        RECT 567.600 67.600 568.400 68.400 ;
        RECT 572.400 67.600 573.200 68.400 ;
        RECT 556.400 51.600 557.200 52.600 ;
        RECT 556.400 49.600 557.200 50.400 ;
        RECT 556.500 38.400 557.100 49.600 ;
        RECT 558.000 46.200 558.800 57.800 ;
        RECT 562.800 57.600 563.600 58.400 ;
        RECT 559.600 53.600 560.400 54.400 ;
        RECT 561.200 50.200 562.000 55.800 ;
        RECT 567.600 46.200 568.400 57.800 ;
        RECT 572.500 54.400 573.100 67.600 ;
        RECT 574.000 64.200 574.800 75.800 ;
        RECT 578.800 74.300 579.600 74.400 ;
        RECT 578.800 73.700 581.100 74.300 ;
        RECT 578.800 73.600 579.600 73.700 ;
        RECT 580.500 70.400 581.100 73.700 ;
        RECT 580.400 69.600 581.200 70.400 ;
        RECT 572.400 53.600 573.200 54.400 ;
        RECT 569.200 51.600 570.000 52.400 ;
        RECT 575.600 51.600 576.400 52.600 ;
        RECT 558.000 43.600 558.800 44.400 ;
        RECT 556.400 37.600 557.200 38.400 ;
        RECT 554.800 31.600 555.600 32.400 ;
        RECT 554.800 28.300 555.600 28.400 ;
        RECT 553.300 27.700 555.600 28.300 ;
        RECT 554.800 27.600 555.600 27.700 ;
        RECT 558.100 26.400 558.700 43.600 ;
        RECT 569.300 38.400 569.900 51.600 ;
        RECT 577.200 46.200 578.000 57.800 ;
        RECT 580.400 50.200 581.200 55.800 ;
        RECT 569.200 37.600 570.000 38.400 ;
        RECT 559.600 31.600 560.400 32.400 ;
        RECT 567.600 31.800 568.400 32.600 ;
        RECT 574.200 31.800 575.000 32.600 ;
        RECT 562.800 29.600 563.600 30.400 ;
        RECT 567.600 28.400 568.200 31.800 ;
        RECT 571.600 28.400 572.400 28.600 ;
        RECT 561.200 27.600 562.000 28.400 ;
        RECT 564.400 27.600 565.200 28.400 ;
        RECT 566.000 27.600 566.800 28.400 ;
        RECT 567.600 27.800 572.400 28.400 ;
        RECT 561.300 26.400 561.900 27.600 ;
        RECT 550.100 25.700 552.300 26.300 ;
        RECT 548.400 21.600 549.200 22.400 ;
        RECT 548.400 18.300 549.200 18.400 ;
        RECT 550.100 18.300 550.700 25.700 ;
        RECT 558.000 25.600 558.800 26.400 ;
        RECT 561.200 25.600 562.000 26.400 ;
        RECT 551.600 23.600 552.400 24.400 ;
        RECT 551.700 18.400 552.300 23.600 ;
        RECT 559.600 19.600 560.400 20.400 ;
        RECT 559.700 18.400 560.300 19.600 ;
        RECT 564.500 18.400 565.100 27.600 ;
        RECT 566.100 22.400 566.700 27.600 ;
        RECT 567.600 27.000 568.200 27.800 ;
        RECT 569.000 27.000 569.800 27.200 ;
        RECT 572.400 27.000 573.200 27.200 ;
        RECT 574.400 27.000 575.000 31.800 ;
        RECT 582.000 31.600 582.800 32.400 ;
        RECT 578.800 29.600 579.600 30.400 ;
        RECT 575.600 27.600 576.400 28.400 ;
        RECT 577.200 27.600 578.000 28.400 ;
        RECT 578.800 27.600 579.600 28.400 ;
        RECT 580.400 27.600 581.200 28.400 ;
        RECT 567.600 26.200 568.400 27.000 ;
        RECT 569.000 26.400 573.200 27.000 ;
        RECT 574.200 26.200 575.000 27.000 ;
        RECT 575.700 26.400 576.300 27.600 ;
        RECT 575.600 25.600 576.400 26.400 ;
        RECT 577.300 24.400 577.900 27.600 ;
        RECT 577.200 23.600 578.000 24.400 ;
        RECT 566.000 21.600 566.800 22.400 ;
        RECT 577.200 21.600 578.000 22.400 ;
        RECT 577.300 18.400 577.900 21.600 ;
        RECT 548.400 17.700 550.700 18.300 ;
        RECT 548.400 17.600 549.200 17.700 ;
        RECT 551.600 17.600 552.400 18.400 ;
        RECT 559.600 17.600 560.400 18.400 ;
        RECT 564.400 17.600 565.200 18.400 ;
        RECT 572.400 17.600 573.200 18.400 ;
        RECT 577.200 17.600 578.000 18.400 ;
        RECT 543.600 15.600 544.400 16.400 ;
        RECT 546.800 15.600 547.600 16.400 ;
        RECT 543.700 14.400 544.300 15.600 ;
        RECT 540.400 13.600 541.200 14.400 ;
        RECT 543.600 13.600 544.400 14.400 ;
        RECT 545.200 13.600 546.000 14.400 ;
        RECT 546.800 13.600 547.600 14.400 ;
        RECT 540.500 12.400 541.100 13.600 ;
        RECT 546.900 12.400 547.500 13.600 ;
        RECT 548.500 12.400 549.100 17.600 ;
        RECT 553.200 15.600 554.000 16.400 ;
        RECT 550.000 13.600 550.800 14.400 ;
        RECT 550.100 12.400 550.700 13.600 ;
        RECT 524.400 11.600 525.200 12.400 ;
        RECT 527.600 11.600 528.400 12.400 ;
        RECT 535.600 11.600 536.400 12.400 ;
        RECT 538.800 11.600 539.600 12.400 ;
        RECT 540.400 11.600 541.200 12.400 ;
        RECT 546.800 11.600 547.600 12.400 ;
        RECT 548.400 11.600 549.200 12.400 ;
        RECT 550.000 11.600 550.800 12.400 ;
        RECT 553.300 10.400 553.900 15.600 ;
        RECT 562.800 15.000 563.600 15.800 ;
        RECT 564.200 15.000 568.400 15.600 ;
        RECT 569.400 15.000 570.200 15.800 ;
        RECT 570.800 15.600 571.600 16.400 ;
        RECT 554.800 13.600 555.600 14.400 ;
        RECT 561.200 13.600 562.000 14.400 ;
        RECT 562.800 14.200 563.400 15.000 ;
        RECT 564.200 14.800 565.000 15.000 ;
        RECT 567.600 14.800 568.400 15.000 ;
        RECT 562.800 13.600 567.600 14.200 ;
        RECT 556.400 11.600 557.200 12.400 ;
        RECT 556.500 10.400 557.100 11.600 ;
        RECT 561.300 10.400 561.900 13.600 ;
        RECT 495.600 10.300 496.400 10.400 ;
        RECT 492.500 9.700 496.400 10.300 ;
        RECT 486.000 9.600 486.800 9.700 ;
        RECT 495.600 9.600 496.400 9.700 ;
        RECT 498.800 9.600 499.600 10.400 ;
        RECT 521.200 9.600 522.000 10.400 ;
        RECT 553.200 9.600 554.000 10.400 ;
        RECT 556.400 9.600 557.200 10.400 ;
        RECT 561.200 9.600 562.000 10.400 ;
        RECT 562.800 10.200 563.400 13.600 ;
        RECT 566.800 13.400 567.600 13.600 ;
        RECT 564.400 11.600 565.200 12.400 ;
        RECT 569.600 10.200 570.200 15.000 ;
        RECT 570.900 14.400 571.500 15.600 ;
        RECT 572.500 14.400 573.100 17.600 ;
        RECT 570.800 13.600 571.600 14.400 ;
        RECT 572.400 13.600 573.200 14.400 ;
        RECT 578.900 12.400 579.500 27.600 ;
        RECT 574.000 11.600 574.800 12.400 ;
        RECT 578.800 11.600 579.600 12.400 ;
        RECT 580.500 10.400 581.100 27.600 ;
        RECT 582.100 18.400 582.700 31.600 ;
        RECT 582.000 17.600 582.800 18.400 ;
        RECT 562.800 9.400 563.600 10.200 ;
        RECT 569.400 9.400 570.200 10.200 ;
        RECT 577.200 9.600 578.000 10.400 ;
        RECT 580.400 9.600 581.200 10.400 ;
        RECT 394.800 7.600 395.600 8.400 ;
        RECT 430.000 7.600 430.800 8.400 ;
      LAYER via2 ;
        RECT 126.000 389.600 126.800 390.400 ;
        RECT 151.600 189.600 152.400 190.400 ;
        RECT 210.800 269.600 211.600 270.400 ;
        RECT 286.000 309.600 286.800 310.400 ;
        RECT 402.800 389.600 403.600 390.400 ;
        RECT 345.200 349.600 346.000 350.400 ;
        RECT 406.000 349.600 406.800 350.400 ;
        RECT 279.600 189.600 280.400 190.400 ;
        RECT 484.400 309.600 485.200 310.400 ;
        RECT 546.800 347.600 547.600 348.400 ;
        RECT 111.600 29.600 112.400 30.400 ;
        RECT 159.600 69.600 160.400 70.400 ;
        RECT 318.000 149.600 318.800 150.400 ;
        RECT 433.200 189.600 434.000 190.400 ;
        RECT 380.400 29.600 381.200 30.400 ;
        RECT 436.400 109.600 437.200 110.400 ;
        RECT 473.200 149.600 474.000 150.400 ;
        RECT 546.800 269.600 547.600 270.400 ;
        RECT 538.800 229.600 539.600 230.400 ;
        RECT 508.400 109.600 509.200 110.400 ;
        RECT 570.800 189.600 571.600 190.400 ;
      LAYER metal3 ;
        RECT 34.800 416.300 35.600 416.400 ;
        RECT 39.600 416.300 40.400 416.400 ;
        RECT 34.800 415.700 40.400 416.300 ;
        RECT 34.800 415.600 35.600 415.700 ;
        RECT 39.600 415.600 40.400 415.700 ;
        RECT 138.800 416.300 139.600 416.400 ;
        RECT 145.200 416.300 146.000 416.400 ;
        RECT 138.800 415.700 146.000 416.300 ;
        RECT 138.800 415.600 139.600 415.700 ;
        RECT 145.200 415.600 146.000 415.700 ;
        RECT 150.000 416.300 150.800 416.400 ;
        RECT 174.000 416.300 174.800 416.400 ;
        RECT 150.000 415.700 174.800 416.300 ;
        RECT 150.000 415.600 150.800 415.700 ;
        RECT 174.000 415.600 174.800 415.700 ;
        RECT 202.800 416.300 203.600 416.400 ;
        RECT 209.200 416.300 210.000 416.400 ;
        RECT 202.800 415.700 210.000 416.300 ;
        RECT 202.800 415.600 203.600 415.700 ;
        RECT 209.200 415.600 210.000 415.700 ;
        RECT 217.200 416.300 218.000 416.400 ;
        RECT 220.400 416.300 221.200 416.400 ;
        RECT 217.200 415.700 221.200 416.300 ;
        RECT 217.200 415.600 218.000 415.700 ;
        RECT 220.400 415.600 221.200 415.700 ;
        RECT 241.200 416.300 242.000 416.400 ;
        RECT 255.600 416.300 256.400 416.400 ;
        RECT 241.200 415.700 256.400 416.300 ;
        RECT 241.200 415.600 242.000 415.700 ;
        RECT 255.600 415.600 256.400 415.700 ;
        RECT 418.800 416.300 419.600 416.400 ;
        RECT 479.600 416.300 480.400 416.400 ;
        RECT 418.800 415.700 480.400 416.300 ;
        RECT 418.800 415.600 419.600 415.700 ;
        RECT 479.600 415.600 480.400 415.700 ;
        RECT 506.800 416.300 507.600 416.400 ;
        RECT 514.800 416.300 515.600 416.400 ;
        RECT 506.800 415.700 515.600 416.300 ;
        RECT 506.800 415.600 507.600 415.700 ;
        RECT 514.800 415.600 515.600 415.700 ;
        RECT 10.800 414.300 11.600 414.400 ;
        RECT 17.200 414.300 18.000 414.400 ;
        RECT 28.400 414.300 29.200 414.400 ;
        RECT 44.400 414.300 45.200 414.400 ;
        RECT 10.800 413.700 45.200 414.300 ;
        RECT 10.800 413.600 11.600 413.700 ;
        RECT 17.200 413.600 18.000 413.700 ;
        RECT 28.400 413.600 29.200 413.700 ;
        RECT 44.400 413.600 45.200 413.700 ;
        RECT 62.000 414.300 62.800 414.400 ;
        RECT 81.200 414.300 82.000 414.400 ;
        RECT 84.400 414.300 85.200 414.400 ;
        RECT 110.000 414.300 110.800 414.400 ;
        RECT 62.000 413.700 110.800 414.300 ;
        RECT 62.000 413.600 62.800 413.700 ;
        RECT 81.200 413.600 82.000 413.700 ;
        RECT 84.400 413.600 85.200 413.700 ;
        RECT 110.000 413.600 110.800 413.700 ;
        RECT 122.800 414.300 123.600 414.400 ;
        RECT 134.000 414.300 134.800 414.400 ;
        RECT 122.800 413.700 134.800 414.300 ;
        RECT 122.800 413.600 123.600 413.700 ;
        RECT 134.000 413.600 134.800 413.700 ;
        RECT 143.600 414.300 144.400 414.400 ;
        RECT 148.400 414.300 149.200 414.400 ;
        RECT 193.200 414.300 194.000 414.400 ;
        RECT 143.600 413.700 149.200 414.300 ;
        RECT 143.600 413.600 144.400 413.700 ;
        RECT 148.400 413.600 149.200 413.700 ;
        RECT 150.100 413.700 194.000 414.300 ;
        RECT 4.400 412.300 5.200 412.400 ;
        RECT 9.200 412.300 10.000 412.400 ;
        RECT 20.400 412.300 21.200 412.400 ;
        RECT 31.600 412.300 32.400 412.400 ;
        RECT 38.000 412.300 38.800 412.400 ;
        RECT 42.800 412.300 43.600 412.400 ;
        RECT 4.400 411.700 43.600 412.300 ;
        RECT 4.400 411.600 5.200 411.700 ;
        RECT 9.200 411.600 10.000 411.700 ;
        RECT 20.400 411.600 21.200 411.700 ;
        RECT 31.600 411.600 32.400 411.700 ;
        RECT 38.000 411.600 38.800 411.700 ;
        RECT 42.800 411.600 43.600 411.700 ;
        RECT 58.800 412.300 59.600 412.400 ;
        RECT 150.100 412.300 150.700 413.700 ;
        RECT 193.200 413.600 194.000 413.700 ;
        RECT 198.000 414.300 198.800 414.400 ;
        RECT 212.400 414.300 213.200 414.400 ;
        RECT 244.400 414.300 245.200 414.400 ;
        RECT 198.000 413.700 245.200 414.300 ;
        RECT 198.000 413.600 198.800 413.700 ;
        RECT 212.400 413.600 213.200 413.700 ;
        RECT 244.400 413.600 245.200 413.700 ;
        RECT 266.800 414.300 267.600 414.400 ;
        RECT 271.600 414.300 272.400 414.400 ;
        RECT 266.800 413.700 272.400 414.300 ;
        RECT 266.800 413.600 267.600 413.700 ;
        RECT 271.600 413.600 272.400 413.700 ;
        RECT 294.000 414.300 294.800 414.400 ;
        RECT 302.000 414.300 302.800 414.400 ;
        RECT 322.800 414.300 323.600 414.400 ;
        RECT 372.400 414.300 373.200 414.400 ;
        RECT 294.000 413.700 373.200 414.300 ;
        RECT 294.000 413.600 294.800 413.700 ;
        RECT 302.000 413.600 302.800 413.700 ;
        RECT 322.800 413.600 323.600 413.700 ;
        RECT 372.400 413.600 373.200 413.700 ;
        RECT 386.800 414.300 387.600 414.400 ;
        RECT 390.000 414.300 390.800 414.400 ;
        RECT 386.800 413.700 390.800 414.300 ;
        RECT 386.800 413.600 387.600 413.700 ;
        RECT 390.000 413.600 390.800 413.700 ;
        RECT 433.200 414.300 434.000 414.400 ;
        RECT 436.400 414.300 437.200 414.400 ;
        RECT 433.200 413.700 437.200 414.300 ;
        RECT 433.200 413.600 434.000 413.700 ;
        RECT 436.400 413.600 437.200 413.700 ;
        RECT 494.000 414.300 494.800 414.400 ;
        RECT 497.200 414.300 498.000 414.400 ;
        RECT 494.000 413.700 498.000 414.300 ;
        RECT 494.000 413.600 494.800 413.700 ;
        RECT 497.200 413.600 498.000 413.700 ;
        RECT 526.000 414.300 526.800 414.400 ;
        RECT 543.600 414.300 544.400 414.400 ;
        RECT 526.000 413.700 544.400 414.300 ;
        RECT 526.000 413.600 526.800 413.700 ;
        RECT 543.600 413.600 544.400 413.700 ;
        RECT 569.200 414.300 570.000 414.400 ;
        RECT 580.400 414.300 581.200 414.400 ;
        RECT 569.200 413.700 581.200 414.300 ;
        RECT 569.200 413.600 570.000 413.700 ;
        RECT 580.400 413.600 581.200 413.700 ;
        RECT 58.800 411.700 150.700 412.300 ;
        RECT 167.600 412.300 168.400 412.400 ;
        RECT 177.200 412.300 178.000 412.400 ;
        RECT 167.600 411.700 178.000 412.300 ;
        RECT 58.800 411.600 59.600 411.700 ;
        RECT 167.600 411.600 168.400 411.700 ;
        RECT 177.200 411.600 178.000 411.700 ;
        RECT 180.400 412.300 181.200 412.400 ;
        RECT 186.800 412.300 187.600 412.400 ;
        RECT 180.400 411.700 187.600 412.300 ;
        RECT 180.400 411.600 181.200 411.700 ;
        RECT 186.800 411.600 187.600 411.700 ;
        RECT 194.800 412.300 195.600 412.400 ;
        RECT 201.200 412.300 202.000 412.400 ;
        RECT 194.800 411.700 202.000 412.300 ;
        RECT 194.800 411.600 195.600 411.700 ;
        RECT 201.200 411.600 202.000 411.700 ;
        RECT 207.600 412.300 208.400 412.400 ;
        RECT 210.800 412.300 211.600 412.400 ;
        RECT 207.600 411.700 211.600 412.300 ;
        RECT 207.600 411.600 208.400 411.700 ;
        RECT 210.800 411.600 211.600 411.700 ;
        RECT 233.200 412.300 234.000 412.400 ;
        RECT 239.600 412.300 240.400 412.400 ;
        RECT 233.200 411.700 240.400 412.300 ;
        RECT 233.200 411.600 234.000 411.700 ;
        RECT 239.600 411.600 240.400 411.700 ;
        RECT 265.200 412.300 266.000 412.400 ;
        RECT 273.200 412.300 274.000 412.400 ;
        RECT 265.200 411.700 274.000 412.300 ;
        RECT 265.200 411.600 266.000 411.700 ;
        RECT 273.200 411.600 274.000 411.700 ;
        RECT 329.200 412.300 330.000 412.400 ;
        RECT 338.800 412.300 339.600 412.400 ;
        RECT 329.200 411.700 339.600 412.300 ;
        RECT 329.200 411.600 330.000 411.700 ;
        RECT 338.800 411.600 339.600 411.700 ;
        RECT 345.200 412.300 346.000 412.400 ;
        RECT 354.800 412.300 355.600 412.400 ;
        RECT 345.200 411.700 355.600 412.300 ;
        RECT 345.200 411.600 346.000 411.700 ;
        RECT 354.800 411.600 355.600 411.700 ;
        RECT 385.200 412.300 386.000 412.400 ;
        RECT 393.200 412.300 394.000 412.400 ;
        RECT 385.200 411.700 394.000 412.300 ;
        RECT 385.200 411.600 386.000 411.700 ;
        RECT 393.200 411.600 394.000 411.700 ;
        RECT 431.600 412.300 432.400 412.400 ;
        RECT 441.200 412.300 442.000 412.400 ;
        RECT 431.600 411.700 442.000 412.300 ;
        RECT 431.600 411.600 432.400 411.700 ;
        RECT 441.200 411.600 442.000 411.700 ;
        RECT 492.400 412.300 493.200 412.400 ;
        RECT 502.000 412.300 502.800 412.400 ;
        RECT 492.400 411.700 502.800 412.300 ;
        RECT 492.400 411.600 493.200 411.700 ;
        RECT 502.000 411.600 502.800 411.700 ;
        RECT 546.800 412.300 547.600 412.400 ;
        RECT 558.000 412.300 558.800 412.400 ;
        RECT 546.800 411.700 558.800 412.300 ;
        RECT 546.800 411.600 547.600 411.700 ;
        RECT 558.000 411.600 558.800 411.700 ;
        RECT 1.200 410.300 2.000 410.400 ;
        RECT 34.800 410.300 35.600 410.400 ;
        RECT 1.200 409.700 35.600 410.300 ;
        RECT 1.200 409.600 2.000 409.700 ;
        RECT 34.800 409.600 35.600 409.700 ;
        RECT 78.000 410.300 78.800 410.400 ;
        RECT 126.000 410.300 126.800 410.400 ;
        RECT 78.000 409.700 126.800 410.300 ;
        RECT 78.000 409.600 78.800 409.700 ;
        RECT 126.000 409.600 126.800 409.700 ;
        RECT 142.000 410.300 142.800 410.400 ;
        RECT 164.400 410.300 165.200 410.400 ;
        RECT 178.800 410.300 179.600 410.400 ;
        RECT 142.000 409.700 179.600 410.300 ;
        RECT 142.000 409.600 142.800 409.700 ;
        RECT 164.400 409.600 165.200 409.700 ;
        RECT 178.800 409.600 179.600 409.700 ;
        RECT 182.000 410.300 182.800 410.400 ;
        RECT 199.600 410.300 200.400 410.400 ;
        RECT 218.800 410.300 219.600 410.400 ;
        RECT 182.000 409.700 219.600 410.300 ;
        RECT 182.000 409.600 182.800 409.700 ;
        RECT 199.600 409.600 200.400 409.700 ;
        RECT 218.800 409.600 219.600 409.700 ;
        RECT 228.400 410.300 229.200 410.400 ;
        RECT 249.200 410.300 250.000 410.400 ;
        RECT 319.600 410.300 320.400 410.400 ;
        RECT 228.400 409.700 320.400 410.300 ;
        RECT 228.400 409.600 229.200 409.700 ;
        RECT 249.200 409.600 250.000 409.700 ;
        RECT 319.600 409.600 320.400 409.700 ;
        RECT 42.800 408.300 43.600 408.400 ;
        RECT 57.200 408.300 58.000 408.400 ;
        RECT 65.200 408.300 66.000 408.400 ;
        RECT 42.800 407.700 66.000 408.300 ;
        RECT 42.800 407.600 43.600 407.700 ;
        RECT 57.200 407.600 58.000 407.700 ;
        RECT 65.200 407.600 66.000 407.700 ;
        RECT 116.400 408.300 117.200 408.400 ;
        RECT 153.200 408.300 154.000 408.400 ;
        RECT 116.400 407.700 154.000 408.300 ;
        RECT 116.400 407.600 117.200 407.700 ;
        RECT 153.200 407.600 154.000 407.700 ;
        RECT 172.400 408.300 173.200 408.400 ;
        RECT 191.600 408.300 192.400 408.400 ;
        RECT 300.400 408.300 301.200 408.400 ;
        RECT 172.400 407.700 301.200 408.300 ;
        RECT 172.400 407.600 173.200 407.700 ;
        RECT 191.600 407.600 192.400 407.700 ;
        RECT 300.400 407.600 301.200 407.700 ;
        RECT 401.200 408.300 402.000 408.400 ;
        RECT 450.800 408.300 451.600 408.400 ;
        RECT 401.200 407.700 451.600 408.300 ;
        RECT 401.200 407.600 402.000 407.700 ;
        RECT 450.800 407.600 451.600 407.700 ;
        RECT 38.000 406.300 38.800 406.400 ;
        RECT 62.000 406.300 62.800 406.400 ;
        RECT 38.000 405.700 62.800 406.300 ;
        RECT 38.000 405.600 38.800 405.700 ;
        RECT 62.000 405.600 62.800 405.700 ;
        RECT 98.800 406.300 99.600 406.400 ;
        RECT 278.000 406.300 278.800 406.400 ;
        RECT 98.800 405.700 278.800 406.300 ;
        RECT 98.800 405.600 99.600 405.700 ;
        RECT 278.000 405.600 278.800 405.700 ;
        RECT 26.800 404.300 27.600 404.400 ;
        RECT 38.000 404.300 38.800 404.400 ;
        RECT 26.800 403.700 38.800 404.300 ;
        RECT 26.800 403.600 27.600 403.700 ;
        RECT 38.000 403.600 38.800 403.700 ;
        RECT 159.600 404.300 160.400 404.400 ;
        RECT 166.000 404.300 166.800 404.400 ;
        RECT 193.200 404.300 194.000 404.400 ;
        RECT 226.800 404.300 227.600 404.400 ;
        RECT 159.600 403.700 227.600 404.300 ;
        RECT 159.600 403.600 160.400 403.700 ;
        RECT 166.000 403.600 166.800 403.700 ;
        RECT 193.200 403.600 194.000 403.700 ;
        RECT 226.800 403.600 227.600 403.700 ;
        RECT 242.800 404.300 243.600 404.400 ;
        RECT 266.800 404.300 267.600 404.400 ;
        RECT 242.800 403.700 267.600 404.300 ;
        RECT 242.800 403.600 243.600 403.700 ;
        RECT 266.800 403.600 267.600 403.700 ;
        RECT 356.400 404.300 357.200 404.400 ;
        RECT 410.800 404.300 411.600 404.400 ;
        RECT 356.400 403.700 411.600 404.300 ;
        RECT 356.400 403.600 357.200 403.700 ;
        RECT 410.800 403.600 411.600 403.700 ;
        RECT 463.600 403.600 464.400 404.400 ;
        RECT 186.800 402.300 187.600 402.400 ;
        RECT 201.200 402.300 202.000 402.400 ;
        RECT 186.800 401.700 202.000 402.300 ;
        RECT 186.800 401.600 187.600 401.700 ;
        RECT 201.200 401.600 202.000 401.700 ;
        RECT 209.200 402.300 210.000 402.400 ;
        RECT 254.000 402.300 254.800 402.400 ;
        RECT 209.200 401.700 254.800 402.300 ;
        RECT 209.200 401.600 210.000 401.700 ;
        RECT 254.000 401.600 254.800 401.700 ;
        RECT 255.600 402.300 256.400 402.400 ;
        RECT 367.600 402.300 368.400 402.400 ;
        RECT 255.600 401.700 368.400 402.300 ;
        RECT 255.600 401.600 256.400 401.700 ;
        RECT 367.600 401.600 368.400 401.700 ;
        RECT 537.200 402.300 538.000 402.400 ;
        RECT 551.600 402.300 552.400 402.400 ;
        RECT 537.200 401.700 552.400 402.300 ;
        RECT 537.200 401.600 538.000 401.700 ;
        RECT 551.600 401.600 552.400 401.700 ;
        RECT 562.800 402.300 563.600 402.400 ;
        RECT 566.000 402.300 566.800 402.400 ;
        RECT 562.800 401.700 566.800 402.300 ;
        RECT 562.800 401.600 563.600 401.700 ;
        RECT 566.000 401.600 566.800 401.700 ;
        RECT 175.600 400.300 176.400 400.400 ;
        RECT 233.200 400.300 234.000 400.400 ;
        RECT 305.200 400.300 306.000 400.400 ;
        RECT 175.600 399.700 306.000 400.300 ;
        RECT 175.600 399.600 176.400 399.700 ;
        RECT 233.200 399.600 234.000 399.700 ;
        RECT 305.200 399.600 306.000 399.700 ;
        RECT 402.800 400.300 403.600 400.400 ;
        RECT 438.000 400.300 438.800 400.400 ;
        RECT 402.800 399.700 438.800 400.300 ;
        RECT 402.800 399.600 403.600 399.700 ;
        RECT 438.000 399.600 438.800 399.700 ;
        RECT 457.200 400.300 458.000 400.400 ;
        RECT 473.200 400.300 474.000 400.400 ;
        RECT 457.200 399.700 474.000 400.300 ;
        RECT 457.200 399.600 458.000 399.700 ;
        RECT 473.200 399.600 474.000 399.700 ;
        RECT 22.000 398.300 22.800 398.400 ;
        RECT 49.200 398.300 50.000 398.400 ;
        RECT 22.000 397.700 50.000 398.300 ;
        RECT 22.000 397.600 22.800 397.700 ;
        RECT 49.200 397.600 50.000 397.700 ;
        RECT 132.400 398.300 133.200 398.400 ;
        RECT 161.200 398.300 162.000 398.400 ;
        RECT 180.400 398.300 181.200 398.400 ;
        RECT 132.400 397.700 181.200 398.300 ;
        RECT 132.400 397.600 133.200 397.700 ;
        RECT 161.200 397.600 162.000 397.700 ;
        RECT 180.400 397.600 181.200 397.700 ;
        RECT 188.400 398.300 189.200 398.400 ;
        RECT 199.600 398.300 200.400 398.400 ;
        RECT 188.400 397.700 200.400 398.300 ;
        RECT 188.400 397.600 189.200 397.700 ;
        RECT 199.600 397.600 200.400 397.700 ;
        RECT 201.200 398.300 202.000 398.400 ;
        RECT 215.600 398.300 216.400 398.400 ;
        RECT 201.200 397.700 216.400 398.300 ;
        RECT 201.200 397.600 202.000 397.700 ;
        RECT 215.600 397.600 216.400 397.700 ;
        RECT 273.200 398.300 274.000 398.400 ;
        RECT 278.000 398.300 278.800 398.400 ;
        RECT 316.400 398.300 317.200 398.400 ;
        RECT 324.400 398.300 325.200 398.400 ;
        RECT 330.800 398.300 331.600 398.400 ;
        RECT 273.200 397.700 331.600 398.300 ;
        RECT 273.200 397.600 274.000 397.700 ;
        RECT 278.000 397.600 278.800 397.700 ;
        RECT 316.400 397.600 317.200 397.700 ;
        RECT 324.400 397.600 325.200 397.700 ;
        RECT 330.800 397.600 331.600 397.700 ;
        RECT 7.600 396.300 8.400 396.400 ;
        RECT 42.800 396.300 43.600 396.400 ;
        RECT 54.000 396.300 54.800 396.400 ;
        RECT 7.600 395.700 54.800 396.300 ;
        RECT 7.600 395.600 8.400 395.700 ;
        RECT 42.800 395.600 43.600 395.700 ;
        RECT 54.000 395.600 54.800 395.700 ;
        RECT 145.200 396.300 146.000 396.400 ;
        RECT 183.600 396.300 184.400 396.400 ;
        RECT 185.200 396.300 186.000 396.400 ;
        RECT 234.800 396.300 235.600 396.400 ;
        RECT 145.200 395.700 235.600 396.300 ;
        RECT 145.200 395.600 146.000 395.700 ;
        RECT 183.600 395.600 184.400 395.700 ;
        RECT 185.200 395.600 186.000 395.700 ;
        RECT 234.800 395.600 235.600 395.700 ;
        RECT 2.800 394.300 3.600 394.400 ;
        RECT 33.200 394.300 34.000 394.400 ;
        RECT 2.800 393.700 34.000 394.300 ;
        RECT 2.800 393.600 3.600 393.700 ;
        RECT 33.200 393.600 34.000 393.700 ;
        RECT 38.000 394.300 38.800 394.400 ;
        RECT 76.400 394.300 77.200 394.400 ;
        RECT 100.400 394.300 101.200 394.400 ;
        RECT 38.000 393.700 101.200 394.300 ;
        RECT 38.000 393.600 38.800 393.700 ;
        RECT 76.400 393.600 77.200 393.700 ;
        RECT 100.400 393.600 101.200 393.700 ;
        RECT 148.400 394.300 149.200 394.400 ;
        RECT 159.600 394.300 160.400 394.400 ;
        RECT 170.800 394.300 171.600 394.400 ;
        RECT 175.600 394.300 176.400 394.400 ;
        RECT 214.000 394.300 214.800 394.400 ;
        RECT 148.400 393.700 214.800 394.300 ;
        RECT 148.400 393.600 149.200 393.700 ;
        RECT 159.600 393.600 160.400 393.700 ;
        RECT 170.800 393.600 171.600 393.700 ;
        RECT 175.600 393.600 176.400 393.700 ;
        RECT 214.000 393.600 214.800 393.700 ;
        RECT 220.400 394.300 221.200 394.400 ;
        RECT 242.800 394.300 243.600 394.400 ;
        RECT 247.600 394.300 248.400 394.400 ;
        RECT 220.400 393.700 248.400 394.300 ;
        RECT 220.400 393.600 221.200 393.700 ;
        RECT 242.800 393.600 243.600 393.700 ;
        RECT 247.600 393.600 248.400 393.700 ;
        RECT 22.000 392.300 22.800 392.400 ;
        RECT 25.200 392.300 26.000 392.400 ;
        RECT 22.000 391.700 26.000 392.300 ;
        RECT 22.000 391.600 22.800 391.700 ;
        RECT 25.200 391.600 26.000 391.700 ;
        RECT 41.200 392.300 42.000 392.400 ;
        RECT 44.400 392.300 45.200 392.400 ;
        RECT 41.200 391.700 45.200 392.300 ;
        RECT 41.200 391.600 42.000 391.700 ;
        RECT 44.400 391.600 45.200 391.700 ;
        RECT 79.600 392.300 80.400 392.400 ;
        RECT 86.000 392.300 86.800 392.400 ;
        RECT 79.600 391.700 86.800 392.300 ;
        RECT 79.600 391.600 80.400 391.700 ;
        RECT 86.000 391.600 86.800 391.700 ;
        RECT 89.200 392.300 90.000 392.400 ;
        RECT 97.200 392.300 98.000 392.400 ;
        RECT 108.400 392.300 109.200 392.400 ;
        RECT 114.800 392.300 115.600 392.400 ;
        RECT 89.200 391.700 115.600 392.300 ;
        RECT 89.200 391.600 90.000 391.700 ;
        RECT 97.200 391.600 98.000 391.700 ;
        RECT 108.400 391.600 109.200 391.700 ;
        RECT 114.800 391.600 115.600 391.700 ;
        RECT 158.000 392.300 158.800 392.400 ;
        RECT 170.800 392.300 171.600 392.400 ;
        RECT 177.200 392.300 178.000 392.400 ;
        RECT 194.800 392.300 195.600 392.400 ;
        RECT 204.400 392.300 205.200 392.400 ;
        RECT 158.000 391.700 205.200 392.300 ;
        RECT 158.000 391.600 158.800 391.700 ;
        RECT 170.800 391.600 171.600 391.700 ;
        RECT 177.200 391.600 178.000 391.700 ;
        RECT 194.800 391.600 195.600 391.700 ;
        RECT 204.400 391.600 205.200 391.700 ;
        RECT 226.800 392.300 227.600 392.400 ;
        RECT 242.800 392.300 243.600 392.400 ;
        RECT 226.800 391.700 243.600 392.300 ;
        RECT 226.800 391.600 227.600 391.700 ;
        RECT 242.800 391.600 243.600 391.700 ;
        RECT 254.000 392.300 254.800 392.400 ;
        RECT 271.600 392.300 272.400 392.400 ;
        RECT 254.000 391.700 272.400 392.300 ;
        RECT 254.000 391.600 254.800 391.700 ;
        RECT 271.600 391.600 272.400 391.700 ;
        RECT 276.400 392.300 277.200 392.400 ;
        RECT 279.600 392.300 280.400 392.400 ;
        RECT 276.400 391.700 280.400 392.300 ;
        RECT 276.400 391.600 277.200 391.700 ;
        RECT 279.600 391.600 280.400 391.700 ;
        RECT 308.400 392.300 309.200 392.400 ;
        RECT 311.600 392.300 312.400 392.400 ;
        RECT 308.400 391.700 312.400 392.300 ;
        RECT 308.400 391.600 309.200 391.700 ;
        RECT 311.600 391.600 312.400 391.700 ;
        RECT 313.200 392.300 314.000 392.400 ;
        RECT 326.000 392.300 326.800 392.400 ;
        RECT 313.200 391.700 326.800 392.300 ;
        RECT 313.200 391.600 314.000 391.700 ;
        RECT 326.000 391.600 326.800 391.700 ;
        RECT 15.600 390.300 16.400 390.400 ;
        RECT 47.600 390.300 48.400 390.400 ;
        RECT 52.400 390.300 53.200 390.400 ;
        RECT 15.600 389.700 53.200 390.300 ;
        RECT 15.600 389.600 16.400 389.700 ;
        RECT 47.600 389.600 48.400 389.700 ;
        RECT 52.400 389.600 53.200 389.700 ;
        RECT 62.000 390.300 62.800 390.400 ;
        RECT 92.400 390.300 93.200 390.400 ;
        RECT 105.200 390.300 106.000 390.400 ;
        RECT 62.000 389.700 106.000 390.300 ;
        RECT 62.000 389.600 62.800 389.700 ;
        RECT 92.400 389.600 93.200 389.700 ;
        RECT 105.200 389.600 106.000 389.700 ;
        RECT 126.000 390.300 126.800 390.400 ;
        RECT 140.400 390.300 141.200 390.400 ;
        RECT 126.000 389.700 141.200 390.300 ;
        RECT 126.000 389.600 126.800 389.700 ;
        RECT 140.400 389.600 141.200 389.700 ;
        RECT 162.800 390.300 163.600 390.400 ;
        RECT 166.000 390.300 166.800 390.400 ;
        RECT 162.800 389.700 166.800 390.300 ;
        RECT 162.800 389.600 163.600 389.700 ;
        RECT 166.000 389.600 166.800 389.700 ;
        RECT 167.600 390.300 168.400 390.400 ;
        RECT 172.400 390.300 173.200 390.400 ;
        RECT 167.600 389.700 173.200 390.300 ;
        RECT 167.600 389.600 168.400 389.700 ;
        RECT 172.400 389.600 173.200 389.700 ;
        RECT 188.400 390.300 189.200 390.400 ;
        RECT 196.400 390.300 197.200 390.400 ;
        RECT 188.400 389.700 197.200 390.300 ;
        RECT 188.400 389.600 189.200 389.700 ;
        RECT 196.400 389.600 197.200 389.700 ;
        RECT 198.000 390.300 198.800 390.400 ;
        RECT 228.400 390.300 229.200 390.400 ;
        RECT 198.000 389.700 229.200 390.300 ;
        RECT 198.000 389.600 198.800 389.700 ;
        RECT 228.400 389.600 229.200 389.700 ;
        RECT 270.000 390.300 270.800 390.400 ;
        RECT 281.200 390.300 282.000 390.400 ;
        RECT 270.000 389.700 282.000 390.300 ;
        RECT 270.000 389.600 270.800 389.700 ;
        RECT 281.200 389.600 282.000 389.700 ;
        RECT 292.400 390.300 293.200 390.400 ;
        RECT 313.300 390.300 313.900 391.600 ;
        RECT 292.400 389.700 313.900 390.300 ;
        RECT 321.200 390.300 322.000 390.400 ;
        RECT 327.600 390.300 328.400 390.400 ;
        RECT 321.200 389.700 328.400 390.300 ;
        RECT 292.400 389.600 293.200 389.700 ;
        RECT 321.200 389.600 322.000 389.700 ;
        RECT 327.600 389.600 328.400 389.700 ;
        RECT 348.400 390.300 349.200 390.400 ;
        RECT 353.200 390.300 354.000 390.400 ;
        RECT 361.200 390.300 362.000 390.400 ;
        RECT 348.400 389.700 362.000 390.300 ;
        RECT 348.400 389.600 349.200 389.700 ;
        RECT 353.200 389.600 354.000 389.700 ;
        RECT 361.200 389.600 362.000 389.700 ;
        RECT 377.200 390.300 378.000 390.400 ;
        RECT 396.400 390.300 397.200 390.400 ;
        RECT 377.200 389.700 397.200 390.300 ;
        RECT 377.200 389.600 378.000 389.700 ;
        RECT 396.400 389.600 397.200 389.700 ;
        RECT 402.800 390.300 403.600 390.400 ;
        RECT 414.000 390.300 414.800 390.400 ;
        RECT 423.600 390.300 424.400 390.400 ;
        RECT 428.400 390.300 429.200 390.400 ;
        RECT 402.800 389.700 429.200 390.300 ;
        RECT 402.800 389.600 403.600 389.700 ;
        RECT 414.000 389.600 414.800 389.700 ;
        RECT 423.600 389.600 424.400 389.700 ;
        RECT 428.400 389.600 429.200 389.700 ;
        RECT 473.200 390.300 474.000 390.400 ;
        RECT 481.200 390.300 482.000 390.400 ;
        RECT 473.200 389.700 482.000 390.300 ;
        RECT 473.200 389.600 474.000 389.700 ;
        RECT 481.200 389.600 482.000 389.700 ;
        RECT 498.800 390.300 499.600 390.400 ;
        RECT 505.200 390.300 506.000 390.400 ;
        RECT 498.800 389.700 506.000 390.300 ;
        RECT 498.800 389.600 499.600 389.700 ;
        RECT 505.200 389.600 506.000 389.700 ;
        RECT 1.200 388.300 2.000 388.400 ;
        RECT 7.600 388.300 8.400 388.400 ;
        RECT 1.200 387.700 8.400 388.300 ;
        RECT 1.200 387.600 2.000 387.700 ;
        RECT 7.600 387.600 8.400 387.700 ;
        RECT 10.800 388.300 11.600 388.400 ;
        RECT 22.000 388.300 22.800 388.400 ;
        RECT 10.800 387.700 22.800 388.300 ;
        RECT 10.800 387.600 11.600 387.700 ;
        RECT 22.000 387.600 22.800 387.700 ;
        RECT 54.000 388.300 54.800 388.400 ;
        RECT 63.600 388.300 64.400 388.400 ;
        RECT 54.000 387.700 64.400 388.300 ;
        RECT 54.000 387.600 54.800 387.700 ;
        RECT 63.600 387.600 64.400 387.700 ;
        RECT 74.800 388.300 75.600 388.400 ;
        RECT 82.800 388.300 83.600 388.400 ;
        RECT 74.800 387.700 83.600 388.300 ;
        RECT 74.800 387.600 75.600 387.700 ;
        RECT 82.800 387.600 83.600 387.700 ;
        RECT 92.400 388.300 93.200 388.400 ;
        RECT 98.800 388.300 99.600 388.400 ;
        RECT 100.400 388.300 101.200 388.400 ;
        RECT 92.400 387.700 101.200 388.300 ;
        RECT 92.400 387.600 93.200 387.700 ;
        RECT 98.800 387.600 99.600 387.700 ;
        RECT 100.400 387.600 101.200 387.700 ;
        RECT 103.600 388.300 104.400 388.400 ;
        RECT 108.400 388.300 109.200 388.400 ;
        RECT 111.600 388.300 112.400 388.400 ;
        RECT 124.400 388.300 125.200 388.400 ;
        RECT 103.600 387.700 125.200 388.300 ;
        RECT 103.600 387.600 104.400 387.700 ;
        RECT 108.400 387.600 109.200 387.700 ;
        RECT 111.600 387.600 112.400 387.700 ;
        RECT 124.400 387.600 125.200 387.700 ;
        RECT 161.200 388.300 162.000 388.400 ;
        RECT 166.000 388.300 166.800 388.400 ;
        RECT 161.200 387.700 166.800 388.300 ;
        RECT 161.200 387.600 162.000 387.700 ;
        RECT 166.000 387.600 166.800 387.700 ;
        RECT 178.800 388.300 179.600 388.400 ;
        RECT 190.000 388.300 190.800 388.400 ;
        RECT 178.800 387.700 190.800 388.300 ;
        RECT 178.800 387.600 179.600 387.700 ;
        RECT 190.000 387.600 190.800 387.700 ;
        RECT 202.800 388.300 203.600 388.400 ;
        RECT 212.400 388.300 213.200 388.400 ;
        RECT 202.800 387.700 213.200 388.300 ;
        RECT 202.800 387.600 203.600 387.700 ;
        RECT 212.400 387.600 213.200 387.700 ;
        RECT 220.400 388.300 221.200 388.400 ;
        RECT 223.600 388.300 224.400 388.400 ;
        RECT 220.400 387.700 224.400 388.300 ;
        RECT 220.400 387.600 221.200 387.700 ;
        RECT 223.600 387.600 224.400 387.700 ;
        RECT 228.400 388.300 229.200 388.400 ;
        RECT 238.000 388.300 238.800 388.400 ;
        RECT 228.400 387.700 238.800 388.300 ;
        RECT 228.400 387.600 229.200 387.700 ;
        RECT 238.000 387.600 238.800 387.700 ;
        RECT 265.200 388.300 266.000 388.400 ;
        RECT 274.800 388.300 275.600 388.400 ;
        RECT 265.200 387.700 275.600 388.300 ;
        RECT 265.200 387.600 266.000 387.700 ;
        RECT 274.800 387.600 275.600 387.700 ;
        RECT 298.800 388.300 299.600 388.400 ;
        RECT 303.600 388.300 304.400 388.400 ;
        RECT 298.800 387.700 304.400 388.300 ;
        RECT 298.800 387.600 299.600 387.700 ;
        RECT 303.600 387.600 304.400 387.700 ;
        RECT 342.000 388.300 342.800 388.400 ;
        RECT 348.400 388.300 349.200 388.400 ;
        RECT 342.000 387.700 349.200 388.300 ;
        RECT 342.000 387.600 342.800 387.700 ;
        RECT 348.400 387.600 349.200 387.700 ;
        RECT 354.800 388.300 355.600 388.400 ;
        RECT 358.000 388.300 358.800 388.400 ;
        RECT 369.200 388.300 370.000 388.400 ;
        RECT 374.000 388.300 374.800 388.400 ;
        RECT 354.800 387.700 374.800 388.300 ;
        RECT 354.800 387.600 355.600 387.700 ;
        RECT 358.000 387.600 358.800 387.700 ;
        RECT 369.200 387.600 370.000 387.700 ;
        RECT 374.000 387.600 374.800 387.700 ;
        RECT 410.800 388.300 411.600 388.400 ;
        RECT 418.800 388.300 419.600 388.400 ;
        RECT 410.800 387.700 419.600 388.300 ;
        RECT 410.800 387.600 411.600 387.700 ;
        RECT 418.800 387.600 419.600 387.700 ;
        RECT 474.800 388.300 475.600 388.400 ;
        RECT 478.000 388.300 478.800 388.400 ;
        RECT 474.800 387.700 478.800 388.300 ;
        RECT 474.800 387.600 475.600 387.700 ;
        RECT 478.000 387.600 478.800 387.700 ;
        RECT 545.200 388.300 546.000 388.400 ;
        RECT 559.600 388.300 560.400 388.400 ;
        RECT 545.200 387.700 560.400 388.300 ;
        RECT 545.200 387.600 546.000 387.700 ;
        RECT 559.600 387.600 560.400 387.700 ;
        RECT 30.000 386.300 30.800 386.400 ;
        RECT 33.200 386.300 34.000 386.400 ;
        RECT 30.000 385.700 34.000 386.300 ;
        RECT 30.000 385.600 30.800 385.700 ;
        RECT 33.200 385.600 34.000 385.700 ;
        RECT 36.400 386.300 37.200 386.400 ;
        RECT 41.200 386.300 42.000 386.400 ;
        RECT 36.400 385.700 42.000 386.300 ;
        RECT 36.400 385.600 37.200 385.700 ;
        RECT 41.200 385.600 42.000 385.700 ;
        RECT 137.200 386.300 138.000 386.400 ;
        RECT 162.800 386.300 163.600 386.400 ;
        RECT 137.200 385.700 163.600 386.300 ;
        RECT 137.200 385.600 138.000 385.700 ;
        RECT 162.800 385.600 163.600 385.700 ;
        RECT 169.200 386.300 170.000 386.400 ;
        RECT 186.800 386.300 187.600 386.400 ;
        RECT 169.200 385.700 187.600 386.300 ;
        RECT 169.200 385.600 170.000 385.700 ;
        RECT 186.800 385.600 187.600 385.700 ;
        RECT 190.000 386.300 190.800 386.400 ;
        RECT 191.600 386.300 192.400 386.400 ;
        RECT 190.000 385.700 192.400 386.300 ;
        RECT 190.000 385.600 190.800 385.700 ;
        RECT 191.600 385.600 192.400 385.700 ;
        RECT 196.400 386.300 197.200 386.400 ;
        RECT 254.000 386.300 254.800 386.400 ;
        RECT 196.400 385.700 254.800 386.300 ;
        RECT 196.400 385.600 197.200 385.700 ;
        RECT 254.000 385.600 254.800 385.700 ;
        RECT 255.600 386.300 256.400 386.400 ;
        RECT 271.600 386.300 272.400 386.400 ;
        RECT 255.600 385.700 272.400 386.300 ;
        RECT 255.600 385.600 256.400 385.700 ;
        RECT 271.600 385.600 272.400 385.700 ;
        RECT 302.000 386.300 302.800 386.400 ;
        RECT 322.800 386.300 323.600 386.400 ;
        RECT 302.000 385.700 323.600 386.300 ;
        RECT 302.000 385.600 302.800 385.700 ;
        RECT 322.800 385.600 323.600 385.700 ;
        RECT 474.800 386.300 475.600 386.400 ;
        RECT 479.600 386.300 480.400 386.400 ;
        RECT 474.800 385.700 480.400 386.300 ;
        RECT 474.800 385.600 475.600 385.700 ;
        RECT 479.600 385.600 480.400 385.700 ;
        RECT 487.600 386.300 488.400 386.400 ;
        RECT 495.600 386.300 496.400 386.400 ;
        RECT 487.600 385.700 496.400 386.300 ;
        RECT 487.600 385.600 488.400 385.700 ;
        RECT 495.600 385.600 496.400 385.700 ;
        RECT 15.600 384.300 16.400 384.400 ;
        RECT 113.200 384.300 114.000 384.400 ;
        RECT 15.600 383.700 114.000 384.300 ;
        RECT 15.600 383.600 16.400 383.700 ;
        RECT 113.200 383.600 114.000 383.700 ;
        RECT 148.400 384.300 149.200 384.400 ;
        RECT 246.000 384.300 246.800 384.400 ;
        RECT 148.400 383.700 246.800 384.300 ;
        RECT 148.400 383.600 149.200 383.700 ;
        RECT 246.000 383.600 246.800 383.700 ;
        RECT 249.200 384.300 250.000 384.400 ;
        RECT 286.000 384.300 286.800 384.400 ;
        RECT 249.200 383.700 286.800 384.300 ;
        RECT 249.200 383.600 250.000 383.700 ;
        RECT 286.000 383.600 286.800 383.700 ;
        RECT 287.600 383.600 288.400 384.400 ;
        RECT 502.000 384.300 502.800 384.400 ;
        RECT 514.800 384.300 515.600 384.400 ;
        RECT 502.000 383.700 515.600 384.300 ;
        RECT 502.000 383.600 502.800 383.700 ;
        RECT 514.800 383.600 515.600 383.700 ;
        RECT 127.600 382.300 128.400 382.400 ;
        RECT 214.000 382.300 214.800 382.400 ;
        RECT 246.000 382.300 246.800 382.400 ;
        RECT 127.600 381.700 195.500 382.300 ;
        RECT 127.600 381.600 128.400 381.700 ;
        RECT 63.600 380.300 64.400 380.400 ;
        RECT 151.600 380.300 152.400 380.400 ;
        RECT 63.600 379.700 152.400 380.300 ;
        RECT 194.900 380.300 195.500 381.700 ;
        RECT 214.000 381.700 246.800 382.300 ;
        RECT 214.000 381.600 214.800 381.700 ;
        RECT 246.000 381.600 246.800 381.700 ;
        RECT 254.000 382.300 254.800 382.400 ;
        RECT 287.600 382.300 288.400 382.400 ;
        RECT 254.000 381.700 288.400 382.300 ;
        RECT 254.000 381.600 254.800 381.700 ;
        RECT 287.600 381.600 288.400 381.700 ;
        RECT 258.800 380.300 259.600 380.400 ;
        RECT 194.900 379.700 259.600 380.300 ;
        RECT 63.600 379.600 64.400 379.700 ;
        RECT 151.600 379.600 152.400 379.700 ;
        RECT 258.800 379.600 259.600 379.700 ;
        RECT 262.000 380.300 262.800 380.400 ;
        RECT 266.800 380.300 267.600 380.400 ;
        RECT 262.000 379.700 267.600 380.300 ;
        RECT 262.000 379.600 262.800 379.700 ;
        RECT 266.800 379.600 267.600 379.700 ;
        RECT 305.200 380.300 306.000 380.400 ;
        RECT 311.600 380.300 312.400 380.400 ;
        RECT 322.800 380.300 323.600 380.400 ;
        RECT 305.200 379.700 323.600 380.300 ;
        RECT 305.200 379.600 306.000 379.700 ;
        RECT 311.600 379.600 312.400 379.700 ;
        RECT 322.800 379.600 323.600 379.700 ;
        RECT 434.800 379.600 435.600 380.400 ;
        RECT 439.600 380.300 440.400 380.400 ;
        RECT 444.400 380.300 445.200 380.400 ;
        RECT 439.600 379.700 445.200 380.300 ;
        RECT 439.600 379.600 440.400 379.700 ;
        RECT 444.400 379.600 445.200 379.700 ;
        RECT 510.000 380.300 510.800 380.400 ;
        RECT 511.600 380.300 512.400 380.400 ;
        RECT 510.000 379.700 512.400 380.300 ;
        RECT 510.000 379.600 510.800 379.700 ;
        RECT 511.600 379.600 512.400 379.700 ;
        RECT 524.400 380.300 525.200 380.400 ;
        RECT 530.800 380.300 531.600 380.400 ;
        RECT 524.400 379.700 531.600 380.300 ;
        RECT 524.400 379.600 525.200 379.700 ;
        RECT 530.800 379.600 531.600 379.700 ;
        RECT 34.800 378.300 35.600 378.400 ;
        RECT 89.200 378.300 90.000 378.400 ;
        RECT 34.800 377.700 90.000 378.300 ;
        RECT 34.800 377.600 35.600 377.700 ;
        RECT 89.200 377.600 90.000 377.700 ;
        RECT 153.200 378.300 154.000 378.400 ;
        RECT 233.200 378.300 234.000 378.400 ;
        RECT 153.200 377.700 234.000 378.300 ;
        RECT 153.200 377.600 154.000 377.700 ;
        RECT 233.200 377.600 234.000 377.700 ;
        RECT 242.800 377.600 243.600 378.400 ;
        RECT 252.400 378.300 253.200 378.400 ;
        RECT 270.000 378.300 270.800 378.400 ;
        RECT 276.400 378.300 277.200 378.400 ;
        RECT 252.400 377.700 277.200 378.300 ;
        RECT 252.400 377.600 253.200 377.700 ;
        RECT 270.000 377.600 270.800 377.700 ;
        RECT 276.400 377.600 277.200 377.700 ;
        RECT 287.600 378.300 288.400 378.400 ;
        RECT 311.600 378.300 312.400 378.400 ;
        RECT 287.600 377.700 312.400 378.300 ;
        RECT 287.600 377.600 288.400 377.700 ;
        RECT 311.600 377.600 312.400 377.700 ;
        RECT 372.400 378.300 373.200 378.400 ;
        RECT 393.200 378.300 394.000 378.400 ;
        RECT 420.400 378.300 421.200 378.400 ;
        RECT 428.400 378.300 429.200 378.400 ;
        RECT 460.400 378.300 461.200 378.400 ;
        RECT 372.400 377.700 461.200 378.300 ;
        RECT 372.400 377.600 373.200 377.700 ;
        RECT 393.200 377.600 394.000 377.700 ;
        RECT 420.400 377.600 421.200 377.700 ;
        RECT 428.400 377.600 429.200 377.700 ;
        RECT 460.400 377.600 461.200 377.700 ;
        RECT 31.600 376.300 32.400 376.400 ;
        RECT 36.400 376.300 37.200 376.400 ;
        RECT 73.200 376.300 74.000 376.400 ;
        RECT 31.600 375.700 74.000 376.300 ;
        RECT 31.600 375.600 32.400 375.700 ;
        RECT 36.400 375.600 37.200 375.700 ;
        RECT 73.200 375.600 74.000 375.700 ;
        RECT 175.600 376.300 176.400 376.400 ;
        RECT 178.800 376.300 179.600 376.400 ;
        RECT 175.600 375.700 179.600 376.300 ;
        RECT 175.600 375.600 176.400 375.700 ;
        RECT 178.800 375.600 179.600 375.700 ;
        RECT 180.400 376.300 181.200 376.400 ;
        RECT 191.600 376.300 192.400 376.400 ;
        RECT 180.400 375.700 192.400 376.300 ;
        RECT 180.400 375.600 181.200 375.700 ;
        RECT 191.600 375.600 192.400 375.700 ;
        RECT 194.800 376.300 195.600 376.400 ;
        RECT 202.800 376.300 203.600 376.400 ;
        RECT 194.800 375.700 203.600 376.300 ;
        RECT 194.800 375.600 195.600 375.700 ;
        RECT 202.800 375.600 203.600 375.700 ;
        RECT 204.400 376.300 205.200 376.400 ;
        RECT 207.600 376.300 208.400 376.400 ;
        RECT 204.400 375.700 208.400 376.300 ;
        RECT 204.400 375.600 205.200 375.700 ;
        RECT 207.600 375.600 208.400 375.700 ;
        RECT 210.800 376.300 211.600 376.400 ;
        RECT 230.000 376.300 230.800 376.400 ;
        RECT 210.800 375.700 230.800 376.300 ;
        RECT 210.800 375.600 211.600 375.700 ;
        RECT 230.000 375.600 230.800 375.700 ;
        RECT 239.600 376.300 240.400 376.400 ;
        RECT 255.600 376.300 256.400 376.400 ;
        RECT 239.600 375.700 256.400 376.300 ;
        RECT 239.600 375.600 240.400 375.700 ;
        RECT 255.600 375.600 256.400 375.700 ;
        RECT 274.800 376.300 275.600 376.400 ;
        RECT 287.600 376.300 288.400 376.400 ;
        RECT 318.000 376.300 318.800 376.400 ;
        RECT 274.800 375.700 288.400 376.300 ;
        RECT 274.800 375.600 275.600 375.700 ;
        RECT 287.600 375.600 288.400 375.700 ;
        RECT 289.300 375.700 318.800 376.300 ;
        RECT 289.300 374.400 289.900 375.700 ;
        RECT 318.000 375.600 318.800 375.700 ;
        RECT 351.600 376.300 352.400 376.400 ;
        RECT 362.800 376.300 363.600 376.400 ;
        RECT 367.600 376.300 368.400 376.400 ;
        RECT 351.600 375.700 368.400 376.300 ;
        RECT 351.600 375.600 352.400 375.700 ;
        RECT 362.800 375.600 363.600 375.700 ;
        RECT 367.600 375.600 368.400 375.700 ;
        RECT 374.000 376.300 374.800 376.400 ;
        RECT 382.000 376.300 382.800 376.400 ;
        RECT 390.000 376.300 390.800 376.400 ;
        RECT 374.000 375.700 390.800 376.300 ;
        RECT 374.000 375.600 374.800 375.700 ;
        RECT 382.000 375.600 382.800 375.700 ;
        RECT 390.000 375.600 390.800 375.700 ;
        RECT 450.800 376.300 451.600 376.400 ;
        RECT 455.600 376.300 456.400 376.400 ;
        RECT 487.600 376.300 488.400 376.400 ;
        RECT 450.800 375.700 488.400 376.300 ;
        RECT 450.800 375.600 451.600 375.700 ;
        RECT 455.600 375.600 456.400 375.700 ;
        RECT 487.600 375.600 488.400 375.700 ;
        RECT 497.200 376.300 498.000 376.400 ;
        RECT 502.000 376.300 502.800 376.400 ;
        RECT 497.200 375.700 502.800 376.300 ;
        RECT 497.200 375.600 498.000 375.700 ;
        RECT 502.000 375.600 502.800 375.700 ;
        RECT 2.800 374.300 3.600 374.400 ;
        RECT 6.000 374.300 6.800 374.400 ;
        RECT 2.800 373.700 6.800 374.300 ;
        RECT 2.800 373.600 3.600 373.700 ;
        RECT 6.000 373.600 6.800 373.700 ;
        RECT 10.800 374.300 11.600 374.400 ;
        RECT 12.400 374.300 13.200 374.400 ;
        RECT 17.200 374.300 18.000 374.400 ;
        RECT 10.800 373.700 18.000 374.300 ;
        RECT 10.800 373.600 11.600 373.700 ;
        RECT 12.400 373.600 13.200 373.700 ;
        RECT 17.200 373.600 18.000 373.700 ;
        RECT 31.600 374.300 32.400 374.400 ;
        RECT 47.600 374.300 48.400 374.400 ;
        RECT 31.600 373.700 48.400 374.300 ;
        RECT 31.600 373.600 32.400 373.700 ;
        RECT 47.600 373.600 48.400 373.700 ;
        RECT 65.200 374.300 66.000 374.400 ;
        RECT 84.400 374.300 85.200 374.400 ;
        RECT 65.200 373.700 85.200 374.300 ;
        RECT 65.200 373.600 66.000 373.700 ;
        RECT 84.400 373.600 85.200 373.700 ;
        RECT 129.200 374.300 130.000 374.400 ;
        RECT 150.000 374.300 150.800 374.400 ;
        RECT 129.200 373.700 150.800 374.300 ;
        RECT 129.200 373.600 130.000 373.700 ;
        RECT 150.000 373.600 150.800 373.700 ;
        RECT 196.400 374.300 197.200 374.400 ;
        RECT 199.600 374.300 200.400 374.400 ;
        RECT 196.400 373.700 200.400 374.300 ;
        RECT 196.400 373.600 197.200 373.700 ;
        RECT 199.600 373.600 200.400 373.700 ;
        RECT 212.400 374.300 213.200 374.400 ;
        RECT 225.200 374.300 226.000 374.400 ;
        RECT 212.400 373.700 226.000 374.300 ;
        RECT 212.400 373.600 213.200 373.700 ;
        RECT 225.200 373.600 226.000 373.700 ;
        RECT 226.800 374.300 227.600 374.400 ;
        RECT 228.400 374.300 229.200 374.400 ;
        RECT 226.800 373.700 229.200 374.300 ;
        RECT 226.800 373.600 227.600 373.700 ;
        RECT 228.400 373.600 229.200 373.700 ;
        RECT 230.000 374.300 230.800 374.400 ;
        RECT 250.800 374.300 251.600 374.400 ;
        RECT 279.600 374.300 280.400 374.400 ;
        RECT 289.200 374.300 290.000 374.400 ;
        RECT 230.000 373.700 290.000 374.300 ;
        RECT 230.000 373.600 230.800 373.700 ;
        RECT 250.800 373.600 251.600 373.700 ;
        RECT 279.600 373.600 280.400 373.700 ;
        RECT 289.200 373.600 290.000 373.700 ;
        RECT 302.000 374.300 302.800 374.400 ;
        RECT 305.200 374.300 306.000 374.400 ;
        RECT 302.000 373.700 306.000 374.300 ;
        RECT 302.000 373.600 302.800 373.700 ;
        RECT 305.200 373.600 306.000 373.700 ;
        RECT 343.600 374.300 344.400 374.400 ;
        RECT 361.200 374.300 362.000 374.400 ;
        RECT 343.600 373.700 362.000 374.300 ;
        RECT 343.600 373.600 344.400 373.700 ;
        RECT 361.200 373.600 362.000 373.700 ;
        RECT 362.800 374.300 363.600 374.400 ;
        RECT 364.400 374.300 365.200 374.400 ;
        RECT 385.200 374.300 386.000 374.400 ;
        RECT 362.800 373.700 386.000 374.300 ;
        RECT 362.800 373.600 363.600 373.700 ;
        RECT 364.400 373.600 365.200 373.700 ;
        RECT 385.200 373.600 386.000 373.700 ;
        RECT 561.200 374.300 562.000 374.400 ;
        RECT 578.800 374.300 579.600 374.400 ;
        RECT 561.200 373.700 579.600 374.300 ;
        RECT 561.200 373.600 562.000 373.700 ;
        RECT 578.800 373.600 579.600 373.700 ;
        RECT 6.000 372.300 6.800 372.400 ;
        RECT 23.600 372.300 24.400 372.400 ;
        RECT 31.600 372.300 32.400 372.400 ;
        RECT 6.000 371.700 32.400 372.300 ;
        RECT 6.000 371.600 6.800 371.700 ;
        RECT 23.600 371.600 24.400 371.700 ;
        RECT 31.600 371.600 32.400 371.700 ;
        RECT 62.000 372.300 62.800 372.400 ;
        RECT 63.600 372.300 64.400 372.400 ;
        RECT 62.000 371.700 64.400 372.300 ;
        RECT 62.000 371.600 62.800 371.700 ;
        RECT 63.600 371.600 64.400 371.700 ;
        RECT 71.600 372.300 72.400 372.400 ;
        RECT 76.400 372.300 77.200 372.400 ;
        RECT 71.600 371.700 77.200 372.300 ;
        RECT 71.600 371.600 72.400 371.700 ;
        RECT 76.400 371.600 77.200 371.700 ;
        RECT 90.800 372.300 91.600 372.400 ;
        RECT 94.000 372.300 94.800 372.400 ;
        RECT 90.800 371.700 94.800 372.300 ;
        RECT 90.800 371.600 91.600 371.700 ;
        RECT 94.000 371.600 94.800 371.700 ;
        RECT 146.800 372.300 147.600 372.400 ;
        RECT 183.600 372.300 184.400 372.400 ;
        RECT 199.600 372.300 200.400 372.400 ;
        RECT 207.600 372.300 208.400 372.400 ;
        RECT 209.200 372.300 210.000 372.400 ;
        RECT 210.800 372.300 211.600 372.400 ;
        RECT 146.800 371.700 211.600 372.300 ;
        RECT 146.800 371.600 147.600 371.700 ;
        RECT 183.600 371.600 184.400 371.700 ;
        RECT 199.600 371.600 200.400 371.700 ;
        RECT 207.600 371.600 208.400 371.700 ;
        RECT 209.200 371.600 210.000 371.700 ;
        RECT 210.800 371.600 211.600 371.700 ;
        RECT 217.200 372.300 218.000 372.400 ;
        RECT 218.800 372.300 219.600 372.400 ;
        RECT 244.400 372.300 245.200 372.400 ;
        RECT 257.200 372.300 258.000 372.400 ;
        RECT 217.200 371.700 258.000 372.300 ;
        RECT 217.200 371.600 218.000 371.700 ;
        RECT 218.800 371.600 219.600 371.700 ;
        RECT 244.400 371.600 245.200 371.700 ;
        RECT 257.200 371.600 258.000 371.700 ;
        RECT 262.000 372.300 262.800 372.400 ;
        RECT 266.800 372.300 267.600 372.400 ;
        RECT 276.400 372.300 277.200 372.400 ;
        RECT 262.000 371.700 277.200 372.300 ;
        RECT 262.000 371.600 262.800 371.700 ;
        RECT 266.800 371.600 267.600 371.700 ;
        RECT 276.400 371.600 277.200 371.700 ;
        RECT 350.000 372.300 350.800 372.400 ;
        RECT 377.200 372.300 378.000 372.400 ;
        RECT 350.000 371.700 378.000 372.300 ;
        RECT 350.000 371.600 350.800 371.700 ;
        RECT 377.200 371.600 378.000 371.700 ;
        RECT 399.600 372.300 400.400 372.400 ;
        RECT 406.000 372.300 406.800 372.400 ;
        RECT 418.800 372.300 419.600 372.400 ;
        RECT 399.600 371.700 419.600 372.300 ;
        RECT 399.600 371.600 400.400 371.700 ;
        RECT 406.000 371.600 406.800 371.700 ;
        RECT 418.800 371.600 419.600 371.700 ;
        RECT 434.800 372.300 435.600 372.400 ;
        RECT 438.000 372.300 438.800 372.400 ;
        RECT 434.800 371.700 438.800 372.300 ;
        RECT 434.800 371.600 435.600 371.700 ;
        RECT 438.000 371.600 438.800 371.700 ;
        RECT 441.200 372.300 442.000 372.400 ;
        RECT 446.000 372.300 446.800 372.400 ;
        RECT 441.200 371.700 446.800 372.300 ;
        RECT 441.200 371.600 442.000 371.700 ;
        RECT 446.000 371.600 446.800 371.700 ;
        RECT 487.600 372.300 488.400 372.400 ;
        RECT 492.400 372.300 493.200 372.400 ;
        RECT 487.600 371.700 493.200 372.300 ;
        RECT 487.600 371.600 488.400 371.700 ;
        RECT 492.400 371.600 493.200 371.700 ;
        RECT 511.600 372.300 512.400 372.400 ;
        RECT 514.800 372.300 515.600 372.400 ;
        RECT 527.600 372.300 528.400 372.400 ;
        RECT 511.600 371.700 528.400 372.300 ;
        RECT 511.600 371.600 512.400 371.700 ;
        RECT 514.800 371.600 515.600 371.700 ;
        RECT 527.600 371.600 528.400 371.700 ;
        RECT 20.400 370.300 21.200 370.400 ;
        RECT 28.400 370.300 29.200 370.400 ;
        RECT 20.400 369.700 29.200 370.300 ;
        RECT 20.400 369.600 21.200 369.700 ;
        RECT 28.400 369.600 29.200 369.700 ;
        RECT 34.800 370.300 35.600 370.400 ;
        RECT 36.400 370.300 37.200 370.400 ;
        RECT 46.000 370.300 46.800 370.400 ;
        RECT 68.400 370.300 69.200 370.400 ;
        RECT 34.800 369.700 69.200 370.300 ;
        RECT 34.800 369.600 35.600 369.700 ;
        RECT 36.400 369.600 37.200 369.700 ;
        RECT 46.000 369.600 46.800 369.700 ;
        RECT 68.400 369.600 69.200 369.700 ;
        RECT 110.000 370.300 110.800 370.400 ;
        RECT 162.800 370.300 163.600 370.400 ;
        RECT 110.000 369.700 163.600 370.300 ;
        RECT 110.000 369.600 110.800 369.700 ;
        RECT 162.800 369.600 163.600 369.700 ;
        RECT 186.800 370.300 187.600 370.400 ;
        RECT 204.400 370.300 205.200 370.400 ;
        RECT 222.000 370.300 222.800 370.400 ;
        RECT 239.600 370.300 240.400 370.400 ;
        RECT 186.800 369.700 240.400 370.300 ;
        RECT 186.800 369.600 187.600 369.700 ;
        RECT 204.400 369.600 205.200 369.700 ;
        RECT 222.000 369.600 222.800 369.700 ;
        RECT 239.600 369.600 240.400 369.700 ;
        RECT 255.600 370.300 256.400 370.400 ;
        RECT 278.000 370.300 278.800 370.400 ;
        RECT 255.600 369.700 278.800 370.300 ;
        RECT 255.600 369.600 256.400 369.700 ;
        RECT 278.000 369.600 278.800 369.700 ;
        RECT 286.000 370.300 286.800 370.400 ;
        RECT 302.000 370.300 302.800 370.400 ;
        RECT 286.000 369.700 302.800 370.300 ;
        RECT 286.000 369.600 286.800 369.700 ;
        RECT 302.000 369.600 302.800 369.700 ;
        RECT 324.400 370.300 325.200 370.400 ;
        RECT 353.200 370.300 354.000 370.400 ;
        RECT 324.400 369.700 354.000 370.300 ;
        RECT 324.400 369.600 325.200 369.700 ;
        RECT 353.200 369.600 354.000 369.700 ;
        RECT 375.600 370.300 376.400 370.400 ;
        RECT 380.400 370.300 381.200 370.400 ;
        RECT 375.600 369.700 381.200 370.300 ;
        RECT 375.600 369.600 376.400 369.700 ;
        RECT 380.400 369.600 381.200 369.700 ;
        RECT 14.000 368.300 14.800 368.400 ;
        RECT 42.800 368.300 43.600 368.400 ;
        RECT 14.000 367.700 43.600 368.300 ;
        RECT 14.000 367.600 14.800 367.700 ;
        RECT 42.800 367.600 43.600 367.700 ;
        RECT 73.200 368.300 74.000 368.400 ;
        RECT 97.200 368.300 98.000 368.400 ;
        RECT 73.200 367.700 98.000 368.300 ;
        RECT 73.200 367.600 74.000 367.700 ;
        RECT 97.200 367.600 98.000 367.700 ;
        RECT 172.400 368.300 173.200 368.400 ;
        RECT 190.000 368.300 190.800 368.400 ;
        RECT 172.400 367.700 190.800 368.300 ;
        RECT 172.400 367.600 173.200 367.700 ;
        RECT 190.000 367.600 190.800 367.700 ;
        RECT 193.200 368.300 194.000 368.400 ;
        RECT 207.600 368.300 208.400 368.400 ;
        RECT 193.200 367.700 208.400 368.300 ;
        RECT 193.200 367.600 194.000 367.700 ;
        RECT 207.600 367.600 208.400 367.700 ;
        RECT 215.600 368.300 216.400 368.400 ;
        RECT 225.200 368.300 226.000 368.400 ;
        RECT 241.200 368.300 242.000 368.400 ;
        RECT 250.800 368.300 251.600 368.400 ;
        RECT 215.600 367.700 251.600 368.300 ;
        RECT 215.600 367.600 216.400 367.700 ;
        RECT 225.200 367.600 226.000 367.700 ;
        RECT 241.200 367.600 242.000 367.700 ;
        RECT 250.800 367.600 251.600 367.700 ;
        RECT 255.600 368.300 256.400 368.400 ;
        RECT 263.600 368.300 264.400 368.400 ;
        RECT 255.600 367.700 264.400 368.300 ;
        RECT 255.600 367.600 256.400 367.700 ;
        RECT 263.600 367.600 264.400 367.700 ;
        RECT 354.800 368.300 355.600 368.400 ;
        RECT 366.000 368.300 366.800 368.400 ;
        RECT 380.400 368.300 381.200 368.400 ;
        RECT 354.800 367.700 381.200 368.300 ;
        RECT 354.800 367.600 355.600 367.700 ;
        RECT 366.000 367.600 366.800 367.700 ;
        RECT 380.400 367.600 381.200 367.700 ;
        RECT 6.000 366.300 6.800 366.400 ;
        RECT 22.000 366.300 22.800 366.400 ;
        RECT 6.000 365.700 22.800 366.300 ;
        RECT 6.000 365.600 6.800 365.700 ;
        RECT 22.000 365.600 22.800 365.700 ;
        RECT 38.000 366.300 38.800 366.400 ;
        RECT 74.800 366.300 75.600 366.400 ;
        RECT 38.000 365.700 75.600 366.300 ;
        RECT 38.000 365.600 38.800 365.700 ;
        RECT 74.800 365.600 75.600 365.700 ;
        RECT 76.400 366.300 77.200 366.400 ;
        RECT 116.400 366.300 117.200 366.400 ;
        RECT 76.400 365.700 117.200 366.300 ;
        RECT 76.400 365.600 77.200 365.700 ;
        RECT 116.400 365.600 117.200 365.700 ;
        RECT 191.600 366.300 192.400 366.400 ;
        RECT 223.600 366.300 224.400 366.400 ;
        RECT 191.600 365.700 224.400 366.300 ;
        RECT 191.600 365.600 192.400 365.700 ;
        RECT 223.600 365.600 224.400 365.700 ;
        RECT 18.800 364.300 19.600 364.400 ;
        RECT 22.000 364.300 22.800 364.400 ;
        RECT 30.000 364.300 30.800 364.400 ;
        RECT 49.200 364.300 50.000 364.400 ;
        RECT 18.800 363.700 50.000 364.300 ;
        RECT 18.800 363.600 19.600 363.700 ;
        RECT 22.000 363.600 22.800 363.700 ;
        RECT 30.000 363.600 30.800 363.700 ;
        RECT 49.200 363.600 50.000 363.700 ;
        RECT 78.000 364.300 78.800 364.400 ;
        RECT 98.800 364.300 99.600 364.400 ;
        RECT 78.000 363.700 99.600 364.300 ;
        RECT 78.000 363.600 78.800 363.700 ;
        RECT 98.800 363.600 99.600 363.700 ;
        RECT 130.800 364.300 131.600 364.400 ;
        RECT 140.400 364.300 141.200 364.400 ;
        RECT 130.800 363.700 141.200 364.300 ;
        RECT 130.800 363.600 131.600 363.700 ;
        RECT 140.400 363.600 141.200 363.700 ;
        RECT 177.200 364.300 178.000 364.400 ;
        RECT 201.200 364.300 202.000 364.400 ;
        RECT 177.200 363.700 202.000 364.300 ;
        RECT 177.200 363.600 178.000 363.700 ;
        RECT 201.200 363.600 202.000 363.700 ;
        RECT 412.400 363.600 413.200 364.400 ;
        RECT 498.800 364.300 499.600 364.400 ;
        RECT 518.000 364.300 518.800 364.400 ;
        RECT 535.600 364.300 536.400 364.400 ;
        RECT 542.000 364.300 542.800 364.400 ;
        RECT 498.800 363.700 542.800 364.300 ;
        RECT 498.800 363.600 499.600 363.700 ;
        RECT 518.000 363.600 518.800 363.700 ;
        RECT 535.600 363.600 536.400 363.700 ;
        RECT 542.000 363.600 542.800 363.700 ;
        RECT 9.200 362.300 10.000 362.400 ;
        RECT 20.400 362.300 21.200 362.400 ;
        RECT 26.800 362.300 27.600 362.400 ;
        RECT 9.200 361.700 27.600 362.300 ;
        RECT 9.200 361.600 10.000 361.700 ;
        RECT 20.400 361.600 21.200 361.700 ;
        RECT 26.800 361.600 27.600 361.700 ;
        RECT 34.800 362.300 35.600 362.400 ;
        RECT 39.600 362.300 40.400 362.400 ;
        RECT 34.800 361.700 40.400 362.300 ;
        RECT 34.800 361.600 35.600 361.700 ;
        RECT 39.600 361.600 40.400 361.700 ;
        RECT 47.600 362.300 48.400 362.400 ;
        RECT 54.000 362.300 54.800 362.400 ;
        RECT 47.600 361.700 54.800 362.300 ;
        RECT 47.600 361.600 48.400 361.700 ;
        RECT 54.000 361.600 54.800 361.700 ;
        RECT 244.400 362.300 245.200 362.400 ;
        RECT 334.000 362.300 334.800 362.400 ;
        RECT 244.400 361.700 334.800 362.300 ;
        RECT 244.400 361.600 245.200 361.700 ;
        RECT 334.000 361.600 334.800 361.700 ;
        RECT 25.200 360.300 26.000 360.400 ;
        RECT 57.200 360.300 58.000 360.400 ;
        RECT 60.400 360.300 61.200 360.400 ;
        RECT 25.200 359.700 61.200 360.300 ;
        RECT 25.200 359.600 26.000 359.700 ;
        RECT 57.200 359.600 58.000 359.700 ;
        RECT 60.400 359.600 61.200 359.700 ;
        RECT 159.600 360.300 160.400 360.400 ;
        RECT 194.800 360.300 195.600 360.400 ;
        RECT 287.600 360.300 288.400 360.400 ;
        RECT 159.600 359.700 195.600 360.300 ;
        RECT 159.600 359.600 160.400 359.700 ;
        RECT 194.800 359.600 195.600 359.700 ;
        RECT 196.500 359.700 288.400 360.300 ;
        RECT 166.000 358.300 166.800 358.400 ;
        RECT 196.500 358.300 197.100 359.700 ;
        RECT 287.600 359.600 288.400 359.700 ;
        RECT 166.000 357.700 197.100 358.300 ;
        RECT 223.600 358.300 224.400 358.400 ;
        RECT 244.400 358.300 245.200 358.400 ;
        RECT 223.600 357.700 245.200 358.300 ;
        RECT 166.000 357.600 166.800 357.700 ;
        RECT 223.600 357.600 224.400 357.700 ;
        RECT 244.400 357.600 245.200 357.700 ;
        RECT 249.200 358.300 250.000 358.400 ;
        RECT 262.000 358.300 262.800 358.400 ;
        RECT 289.200 358.300 290.000 358.400 ;
        RECT 249.200 357.700 290.000 358.300 ;
        RECT 249.200 357.600 250.000 357.700 ;
        RECT 262.000 357.600 262.800 357.700 ;
        RECT 289.200 357.600 290.000 357.700 ;
        RECT 369.200 358.300 370.000 358.400 ;
        RECT 378.800 358.300 379.600 358.400 ;
        RECT 369.200 357.700 379.600 358.300 ;
        RECT 369.200 357.600 370.000 357.700 ;
        RECT 378.800 357.600 379.600 357.700 ;
        RECT 473.200 358.300 474.000 358.400 ;
        RECT 481.200 358.300 482.000 358.400 ;
        RECT 473.200 357.700 482.000 358.300 ;
        RECT 473.200 357.600 474.000 357.700 ;
        RECT 481.200 357.600 482.000 357.700 ;
        RECT 185.200 356.300 186.000 356.400 ;
        RECT 268.400 356.300 269.200 356.400 ;
        RECT 185.200 355.700 269.200 356.300 ;
        RECT 185.200 355.600 186.000 355.700 ;
        RECT 268.400 355.600 269.200 355.700 ;
        RECT 270.000 356.300 270.800 356.400 ;
        RECT 326.000 356.300 326.800 356.400 ;
        RECT 270.000 355.700 326.800 356.300 ;
        RECT 270.000 355.600 270.800 355.700 ;
        RECT 326.000 355.600 326.800 355.700 ;
        RECT 15.600 354.300 16.400 354.400 ;
        RECT 18.800 354.300 19.600 354.400 ;
        RECT 15.600 353.700 19.600 354.300 ;
        RECT 15.600 353.600 16.400 353.700 ;
        RECT 18.800 353.600 19.600 353.700 ;
        RECT 42.800 354.300 43.600 354.400 ;
        RECT 63.600 354.300 64.400 354.400 ;
        RECT 42.800 353.700 64.400 354.300 ;
        RECT 42.800 353.600 43.600 353.700 ;
        RECT 63.600 353.600 64.400 353.700 ;
        RECT 150.000 354.300 150.800 354.400 ;
        RECT 159.600 354.300 160.400 354.400 ;
        RECT 178.800 354.300 179.600 354.400 ;
        RECT 198.000 354.300 198.800 354.400 ;
        RECT 150.000 353.700 198.800 354.300 ;
        RECT 150.000 353.600 150.800 353.700 ;
        RECT 159.600 353.600 160.400 353.700 ;
        RECT 178.800 353.600 179.600 353.700 ;
        RECT 198.000 353.600 198.800 353.700 ;
        RECT 201.200 354.300 202.000 354.400 ;
        RECT 215.600 354.300 216.400 354.400 ;
        RECT 266.800 354.300 267.600 354.400 ;
        RECT 276.400 354.300 277.200 354.400 ;
        RECT 292.400 354.300 293.200 354.400 ;
        RECT 201.200 353.700 216.400 354.300 ;
        RECT 201.200 353.600 202.000 353.700 ;
        RECT 215.600 353.600 216.400 353.700 ;
        RECT 217.300 353.700 257.900 354.300 ;
        RECT 28.400 352.300 29.200 352.400 ;
        RECT 49.200 352.300 50.000 352.400 ;
        RECT 28.400 351.700 50.000 352.300 ;
        RECT 28.400 351.600 29.200 351.700 ;
        RECT 49.200 351.600 50.000 351.700 ;
        RECT 60.400 352.300 61.200 352.400 ;
        RECT 65.200 352.300 66.000 352.400 ;
        RECT 60.400 351.700 66.000 352.300 ;
        RECT 60.400 351.600 61.200 351.700 ;
        RECT 65.200 351.600 66.000 351.700 ;
        RECT 87.600 352.300 88.400 352.400 ;
        RECT 113.200 352.300 114.000 352.400 ;
        RECT 118.000 352.300 118.800 352.400 ;
        RECT 87.600 351.700 118.800 352.300 ;
        RECT 87.600 351.600 88.400 351.700 ;
        RECT 113.200 351.600 114.000 351.700 ;
        RECT 118.000 351.600 118.800 351.700 ;
        RECT 130.800 352.300 131.600 352.400 ;
        RECT 135.600 352.300 136.400 352.400 ;
        RECT 130.800 351.700 136.400 352.300 ;
        RECT 130.800 351.600 131.600 351.700 ;
        RECT 135.600 351.600 136.400 351.700 ;
        RECT 137.200 352.300 138.000 352.400 ;
        RECT 199.600 352.300 200.400 352.400 ;
        RECT 137.200 351.700 200.400 352.300 ;
        RECT 137.200 351.600 138.000 351.700 ;
        RECT 199.600 351.600 200.400 351.700 ;
        RECT 207.600 352.300 208.400 352.400 ;
        RECT 217.300 352.300 217.900 353.700 ;
        RECT 207.600 351.700 217.900 352.300 ;
        RECT 207.600 351.600 208.400 351.700 ;
        RECT 233.200 351.600 234.000 352.400 ;
        RECT 247.600 352.300 248.400 352.400 ;
        RECT 255.600 352.300 256.400 352.400 ;
        RECT 247.600 351.700 256.400 352.300 ;
        RECT 257.300 352.300 257.900 353.700 ;
        RECT 266.800 353.700 293.200 354.300 ;
        RECT 266.800 353.600 267.600 353.700 ;
        RECT 276.400 353.600 277.200 353.700 ;
        RECT 292.400 353.600 293.200 353.700 ;
        RECT 410.800 354.300 411.600 354.400 ;
        RECT 425.200 354.300 426.000 354.400 ;
        RECT 431.600 354.300 432.400 354.400 ;
        RECT 410.800 353.700 432.400 354.300 ;
        RECT 410.800 353.600 411.600 353.700 ;
        RECT 425.200 353.600 426.000 353.700 ;
        RECT 431.600 353.600 432.400 353.700 ;
        RECT 474.800 354.300 475.600 354.400 ;
        RECT 484.400 354.300 485.200 354.400 ;
        RECT 474.800 353.700 485.200 354.300 ;
        RECT 474.800 353.600 475.600 353.700 ;
        RECT 484.400 353.600 485.200 353.700 ;
        RECT 268.400 352.300 269.200 352.400 ;
        RECT 278.000 352.300 278.800 352.400 ;
        RECT 257.300 351.700 269.200 352.300 ;
        RECT 247.600 351.600 248.400 351.700 ;
        RECT 255.600 351.600 256.400 351.700 ;
        RECT 268.400 351.600 269.200 351.700 ;
        RECT 270.100 351.700 278.800 352.300 ;
        RECT 4.400 350.300 5.200 350.400 ;
        RECT 6.000 350.300 6.800 350.400 ;
        RECT 4.400 349.700 6.800 350.300 ;
        RECT 4.400 349.600 5.200 349.700 ;
        RECT 6.000 349.600 6.800 349.700 ;
        RECT 17.200 350.300 18.000 350.400 ;
        RECT 41.200 350.300 42.000 350.400 ;
        RECT 62.000 350.300 62.800 350.400 ;
        RECT 17.200 349.700 62.800 350.300 ;
        RECT 17.200 349.600 18.000 349.700 ;
        RECT 41.200 349.600 42.000 349.700 ;
        RECT 62.000 349.600 62.800 349.700 ;
        RECT 68.400 350.300 69.200 350.400 ;
        RECT 74.800 350.300 75.600 350.400 ;
        RECT 68.400 349.700 75.600 350.300 ;
        RECT 68.400 349.600 69.200 349.700 ;
        RECT 74.800 349.600 75.600 349.700 ;
        RECT 116.400 350.300 117.200 350.400 ;
        RECT 121.200 350.300 122.000 350.400 ;
        RECT 132.400 350.300 133.200 350.400 ;
        RECT 116.400 349.700 133.200 350.300 ;
        RECT 116.400 349.600 117.200 349.700 ;
        RECT 121.200 349.600 122.000 349.700 ;
        RECT 132.400 349.600 133.200 349.700 ;
        RECT 196.400 350.300 197.200 350.400 ;
        RECT 209.200 350.300 210.000 350.400 ;
        RECT 196.400 349.700 210.000 350.300 ;
        RECT 196.400 349.600 197.200 349.700 ;
        RECT 209.200 349.600 210.000 349.700 ;
        RECT 214.000 350.300 214.800 350.400 ;
        RECT 228.400 350.300 229.200 350.400 ;
        RECT 214.000 349.700 229.200 350.300 ;
        RECT 214.000 349.600 214.800 349.700 ;
        RECT 228.400 349.600 229.200 349.700 ;
        RECT 231.600 350.300 232.400 350.400 ;
        RECT 236.400 350.300 237.200 350.400 ;
        RECT 249.200 350.300 250.000 350.400 ;
        RECT 231.600 349.700 250.000 350.300 ;
        RECT 231.600 349.600 232.400 349.700 ;
        RECT 236.400 349.600 237.200 349.700 ;
        RECT 249.200 349.600 250.000 349.700 ;
        RECT 265.200 350.300 266.000 350.400 ;
        RECT 270.100 350.300 270.700 351.700 ;
        RECT 278.000 351.600 278.800 351.700 ;
        RECT 294.000 352.300 294.800 352.400 ;
        RECT 303.600 352.300 304.400 352.400 ;
        RECT 294.000 351.700 304.400 352.300 ;
        RECT 294.000 351.600 294.800 351.700 ;
        RECT 303.600 351.600 304.400 351.700 ;
        RECT 412.400 352.300 413.200 352.400 ;
        RECT 417.200 352.300 418.000 352.400 ;
        RECT 412.400 351.700 418.000 352.300 ;
        RECT 412.400 351.600 413.200 351.700 ;
        RECT 417.200 351.600 418.000 351.700 ;
        RECT 426.800 352.300 427.600 352.400 ;
        RECT 441.200 352.300 442.000 352.400 ;
        RECT 426.800 351.700 442.000 352.300 ;
        RECT 426.800 351.600 427.600 351.700 ;
        RECT 441.200 351.600 442.000 351.700 ;
        RECT 450.800 352.300 451.600 352.400 ;
        RECT 463.600 352.300 464.400 352.400 ;
        RECT 468.400 352.300 469.200 352.400 ;
        RECT 450.800 351.700 469.200 352.300 ;
        RECT 450.800 351.600 451.600 351.700 ;
        RECT 463.600 351.600 464.400 351.700 ;
        RECT 468.400 351.600 469.200 351.700 ;
        RECT 265.200 349.700 270.700 350.300 ;
        RECT 274.800 350.300 275.600 350.400 ;
        RECT 294.000 350.300 294.800 350.400 ;
        RECT 274.800 349.700 294.800 350.300 ;
        RECT 265.200 349.600 266.000 349.700 ;
        RECT 274.800 349.600 275.600 349.700 ;
        RECT 294.000 349.600 294.800 349.700 ;
        RECT 298.800 350.300 299.600 350.400 ;
        RECT 314.800 350.300 315.600 350.400 ;
        RECT 298.800 349.700 315.600 350.300 ;
        RECT 298.800 349.600 299.600 349.700 ;
        RECT 314.800 349.600 315.600 349.700 ;
        RECT 345.200 350.300 346.000 350.400 ;
        RECT 351.600 350.300 352.400 350.400 ;
        RECT 345.200 349.700 352.400 350.300 ;
        RECT 345.200 349.600 346.000 349.700 ;
        RECT 351.600 349.600 352.400 349.700 ;
        RECT 364.400 350.300 365.200 350.400 ;
        RECT 374.000 350.300 374.800 350.400 ;
        RECT 364.400 349.700 374.800 350.300 ;
        RECT 364.400 349.600 365.200 349.700 ;
        RECT 374.000 349.600 374.800 349.700 ;
        RECT 406.000 350.300 406.800 350.400 ;
        RECT 412.400 350.300 413.200 350.400 ;
        RECT 406.000 349.700 413.200 350.300 ;
        RECT 406.000 349.600 406.800 349.700 ;
        RECT 412.400 349.600 413.200 349.700 ;
        RECT 415.600 350.300 416.400 350.400 ;
        RECT 430.000 350.300 430.800 350.400 ;
        RECT 415.600 349.700 430.800 350.300 ;
        RECT 415.600 349.600 416.400 349.700 ;
        RECT 430.000 349.600 430.800 349.700 ;
        RECT 434.800 350.300 435.600 350.400 ;
        RECT 452.400 350.300 453.200 350.400 ;
        RECT 457.200 350.300 458.000 350.400 ;
        RECT 434.800 349.700 458.000 350.300 ;
        RECT 434.800 349.600 435.600 349.700 ;
        RECT 452.400 349.600 453.200 349.700 ;
        RECT 457.200 349.600 458.000 349.700 ;
        RECT 514.800 350.300 515.600 350.400 ;
        RECT 518.000 350.300 518.800 350.400 ;
        RECT 514.800 349.700 518.800 350.300 ;
        RECT 514.800 349.600 515.600 349.700 ;
        RECT 518.000 349.600 518.800 349.700 ;
        RECT 18.800 348.300 19.600 348.400 ;
        RECT 33.200 348.300 34.000 348.400 ;
        RECT 46.000 348.300 46.800 348.400 ;
        RECT 47.600 348.300 48.400 348.400 ;
        RECT 18.800 347.700 48.400 348.300 ;
        RECT 18.800 347.600 19.600 347.700 ;
        RECT 33.200 347.600 34.000 347.700 ;
        RECT 46.000 347.600 46.800 347.700 ;
        RECT 47.600 347.600 48.400 347.700 ;
        RECT 50.800 348.300 51.600 348.400 ;
        RECT 55.600 348.300 56.400 348.400 ;
        RECT 50.800 347.700 56.400 348.300 ;
        RECT 50.800 347.600 51.600 347.700 ;
        RECT 55.600 347.600 56.400 347.700 ;
        RECT 62.000 348.300 62.800 348.400 ;
        RECT 78.000 348.300 78.800 348.400 ;
        RECT 79.600 348.300 80.400 348.400 ;
        RECT 62.000 347.700 80.400 348.300 ;
        RECT 62.000 347.600 62.800 347.700 ;
        RECT 78.000 347.600 78.800 347.700 ;
        RECT 79.600 347.600 80.400 347.700 ;
        RECT 89.200 348.300 90.000 348.400 ;
        RECT 102.000 348.300 102.800 348.400 ;
        RECT 119.600 348.300 120.400 348.400 ;
        RECT 142.000 348.300 142.800 348.400 ;
        RECT 172.400 348.300 173.200 348.400 ;
        RECT 183.600 348.300 184.400 348.400 ;
        RECT 89.200 347.700 184.400 348.300 ;
        RECT 89.200 347.600 90.000 347.700 ;
        RECT 102.000 347.600 102.800 347.700 ;
        RECT 119.600 347.600 120.400 347.700 ;
        RECT 142.000 347.600 142.800 347.700 ;
        RECT 172.400 347.600 173.200 347.700 ;
        RECT 183.600 347.600 184.400 347.700 ;
        RECT 196.400 348.300 197.200 348.400 ;
        RECT 209.200 348.300 210.000 348.400 ;
        RECT 196.400 347.700 210.000 348.300 ;
        RECT 196.400 347.600 197.200 347.700 ;
        RECT 209.200 347.600 210.000 347.700 ;
        RECT 222.000 348.300 222.800 348.400 ;
        RECT 238.000 348.300 238.800 348.400 ;
        RECT 321.200 348.300 322.000 348.400 ;
        RECT 326.000 348.300 326.800 348.400 ;
        RECT 222.000 347.700 302.700 348.300 ;
        RECT 222.000 347.600 222.800 347.700 ;
        RECT 238.000 347.600 238.800 347.700 ;
        RECT 302.100 346.400 302.700 347.700 ;
        RECT 321.200 347.700 326.800 348.300 ;
        RECT 321.200 347.600 322.000 347.700 ;
        RECT 326.000 347.600 326.800 347.700 ;
        RECT 348.400 348.300 349.200 348.400 ;
        RECT 370.800 348.300 371.600 348.400 ;
        RECT 402.800 348.300 403.600 348.400 ;
        RECT 348.400 347.700 403.600 348.300 ;
        RECT 348.400 347.600 349.200 347.700 ;
        RECT 370.800 347.600 371.600 347.700 ;
        RECT 402.800 347.600 403.600 347.700 ;
        RECT 417.200 348.300 418.000 348.400 ;
        RECT 426.800 348.300 427.600 348.400 ;
        RECT 417.200 347.700 427.600 348.300 ;
        RECT 417.200 347.600 418.000 347.700 ;
        RECT 426.800 347.600 427.600 347.700 ;
        RECT 438.000 348.300 438.800 348.400 ;
        RECT 449.200 348.300 450.000 348.400 ;
        RECT 454.000 348.300 454.800 348.400 ;
        RECT 438.000 347.700 454.800 348.300 ;
        RECT 438.000 347.600 438.800 347.700 ;
        RECT 449.200 347.600 450.000 347.700 ;
        RECT 454.000 347.600 454.800 347.700 ;
        RECT 458.800 348.300 459.600 348.400 ;
        RECT 468.400 348.300 469.200 348.400 ;
        RECT 458.800 347.700 469.200 348.300 ;
        RECT 458.800 347.600 459.600 347.700 ;
        RECT 468.400 347.600 469.200 347.700 ;
        RECT 521.200 348.300 522.000 348.400 ;
        RECT 527.600 348.300 528.400 348.400 ;
        RECT 521.200 347.700 528.400 348.300 ;
        RECT 521.200 347.600 522.000 347.700 ;
        RECT 527.600 347.600 528.400 347.700 ;
        RECT 546.800 348.300 547.600 348.400 ;
        RECT 562.800 348.300 563.600 348.400 ;
        RECT 546.800 347.700 563.600 348.300 ;
        RECT 546.800 347.600 547.600 347.700 ;
        RECT 562.800 347.600 563.600 347.700 ;
        RECT 6.000 346.300 6.800 346.400 ;
        RECT 7.600 346.300 8.400 346.400 ;
        RECT 22.000 346.300 22.800 346.400 ;
        RECT 6.000 345.700 22.800 346.300 ;
        RECT 6.000 345.600 6.800 345.700 ;
        RECT 7.600 345.600 8.400 345.700 ;
        RECT 22.000 345.600 22.800 345.700 ;
        RECT 33.200 346.300 34.000 346.400 ;
        RECT 38.000 346.300 38.800 346.400 ;
        RECT 33.200 345.700 38.800 346.300 ;
        RECT 33.200 345.600 34.000 345.700 ;
        RECT 38.000 345.600 38.800 345.700 ;
        RECT 44.400 346.300 45.200 346.400 ;
        RECT 47.600 346.300 48.400 346.400 ;
        RECT 44.400 345.700 48.400 346.300 ;
        RECT 44.400 345.600 45.200 345.700 ;
        RECT 47.600 345.600 48.400 345.700 ;
        RECT 60.400 346.300 61.200 346.400 ;
        RECT 76.400 346.300 77.200 346.400 ;
        RECT 82.800 346.300 83.600 346.400 ;
        RECT 60.400 345.700 83.600 346.300 ;
        RECT 60.400 345.600 61.200 345.700 ;
        RECT 76.400 345.600 77.200 345.700 ;
        RECT 82.800 345.600 83.600 345.700 ;
        RECT 106.800 346.300 107.600 346.400 ;
        RECT 137.200 346.300 138.000 346.400 ;
        RECT 106.800 345.700 138.000 346.300 ;
        RECT 106.800 345.600 107.600 345.700 ;
        RECT 137.200 345.600 138.000 345.700 ;
        RECT 218.800 346.300 219.600 346.400 ;
        RECT 231.600 346.300 232.400 346.400 ;
        RECT 218.800 345.700 232.400 346.300 ;
        RECT 218.800 345.600 219.600 345.700 ;
        RECT 231.600 345.600 232.400 345.700 ;
        RECT 244.400 346.300 245.200 346.400 ;
        RECT 247.600 346.300 248.400 346.400 ;
        RECT 244.400 345.700 248.400 346.300 ;
        RECT 244.400 345.600 245.200 345.700 ;
        RECT 247.600 345.600 248.400 345.700 ;
        RECT 255.600 346.300 256.400 346.400 ;
        RECT 274.800 346.300 275.600 346.400 ;
        RECT 255.600 345.700 275.600 346.300 ;
        RECT 255.600 345.600 256.400 345.700 ;
        RECT 274.800 345.600 275.600 345.700 ;
        RECT 284.400 346.300 285.200 346.400 ;
        RECT 295.600 346.300 296.400 346.400 ;
        RECT 284.400 345.700 296.400 346.300 ;
        RECT 284.400 345.600 285.200 345.700 ;
        RECT 295.600 345.600 296.400 345.700 ;
        RECT 302.000 346.300 302.800 346.400 ;
        RECT 310.000 346.300 310.800 346.400 ;
        RECT 330.800 346.300 331.600 346.400 ;
        RECT 302.000 345.700 331.600 346.300 ;
        RECT 302.000 345.600 302.800 345.700 ;
        RECT 310.000 345.600 310.800 345.700 ;
        RECT 330.800 345.600 331.600 345.700 ;
        RECT 423.600 346.300 424.400 346.400 ;
        RECT 450.800 346.300 451.600 346.400 ;
        RECT 423.600 345.700 451.600 346.300 ;
        RECT 423.600 345.600 424.400 345.700 ;
        RECT 450.800 345.600 451.600 345.700 ;
        RECT 511.600 346.300 512.400 346.400 ;
        RECT 530.800 346.300 531.600 346.400 ;
        RECT 511.600 345.700 531.600 346.300 ;
        RECT 511.600 345.600 512.400 345.700 ;
        RECT 530.800 345.600 531.600 345.700 ;
        RECT 36.400 344.300 37.200 344.400 ;
        RECT 42.800 344.300 43.600 344.400 ;
        RECT 52.400 344.300 53.200 344.400 ;
        RECT 36.400 343.700 53.200 344.300 ;
        RECT 36.400 343.600 37.200 343.700 ;
        RECT 42.800 343.600 43.600 343.700 ;
        RECT 52.400 343.600 53.200 343.700 ;
        RECT 68.400 344.300 69.200 344.400 ;
        RECT 122.800 344.300 123.600 344.400 ;
        RECT 68.400 343.700 123.600 344.300 ;
        RECT 68.400 343.600 69.200 343.700 ;
        RECT 122.800 343.600 123.600 343.700 ;
        RECT 148.400 344.300 149.200 344.400 ;
        RECT 154.800 344.300 155.600 344.400 ;
        RECT 148.400 343.700 155.600 344.300 ;
        RECT 148.400 343.600 149.200 343.700 ;
        RECT 154.800 343.600 155.600 343.700 ;
        RECT 194.800 344.300 195.600 344.400 ;
        RECT 225.200 344.300 226.000 344.400 ;
        RECT 194.800 343.700 226.000 344.300 ;
        RECT 194.800 343.600 195.600 343.700 ;
        RECT 225.200 343.600 226.000 343.700 ;
        RECT 249.200 344.300 250.000 344.400 ;
        RECT 298.800 344.300 299.600 344.400 ;
        RECT 327.600 344.300 328.400 344.400 ;
        RECT 354.800 344.300 355.600 344.400 ;
        RECT 249.200 343.700 355.600 344.300 ;
        RECT 249.200 343.600 250.000 343.700 ;
        RECT 298.800 343.600 299.600 343.700 ;
        RECT 327.600 343.600 328.400 343.700 ;
        RECT 354.800 343.600 355.600 343.700 ;
        RECT 442.800 344.300 443.600 344.400 ;
        RECT 455.600 344.300 456.400 344.400 ;
        RECT 442.800 343.700 456.400 344.300 ;
        RECT 442.800 343.600 443.600 343.700 ;
        RECT 455.600 343.600 456.400 343.700 ;
        RECT 578.800 344.300 579.600 344.400 ;
        RECT 582.000 344.300 582.800 344.400 ;
        RECT 578.800 343.700 582.800 344.300 ;
        RECT 578.800 343.600 579.600 343.700 ;
        RECT 582.000 343.600 582.800 343.700 ;
        RECT 18.800 342.300 19.600 342.400 ;
        RECT 79.600 342.300 80.400 342.400 ;
        RECT 18.800 341.700 80.400 342.300 ;
        RECT 18.800 341.600 19.600 341.700 ;
        RECT 79.600 341.600 80.400 341.700 ;
        RECT 116.400 342.300 117.200 342.400 ;
        RECT 119.600 342.300 120.400 342.400 ;
        RECT 151.600 342.300 152.400 342.400 ;
        RECT 116.400 341.700 152.400 342.300 ;
        RECT 116.400 341.600 117.200 341.700 ;
        RECT 119.600 341.600 120.400 341.700 ;
        RECT 151.600 341.600 152.400 341.700 ;
        RECT 262.000 342.300 262.800 342.400 ;
        RECT 271.600 342.300 272.400 342.400 ;
        RECT 262.000 341.700 272.400 342.300 ;
        RECT 262.000 341.600 262.800 341.700 ;
        RECT 271.600 341.600 272.400 341.700 ;
        RECT 311.600 342.300 312.400 342.400 ;
        RECT 318.000 342.300 318.800 342.400 ;
        RECT 311.600 341.700 318.800 342.300 ;
        RECT 311.600 341.600 312.400 341.700 ;
        RECT 318.000 341.600 318.800 341.700 ;
        RECT 38.000 340.300 38.800 340.400 ;
        RECT 54.000 340.300 54.800 340.400 ;
        RECT 58.800 340.300 59.600 340.400 ;
        RECT 74.800 340.300 75.600 340.400 ;
        RECT 38.000 339.700 75.600 340.300 ;
        RECT 38.000 339.600 38.800 339.700 ;
        RECT 54.000 339.600 54.800 339.700 ;
        RECT 58.800 339.600 59.600 339.700 ;
        RECT 74.800 339.600 75.600 339.700 ;
        RECT 153.200 340.300 154.000 340.400 ;
        RECT 174.000 340.300 174.800 340.400 ;
        RECT 153.200 339.700 174.800 340.300 ;
        RECT 153.200 339.600 154.000 339.700 ;
        RECT 174.000 339.600 174.800 339.700 ;
        RECT 262.000 340.300 262.800 340.400 ;
        RECT 266.800 340.300 267.600 340.400 ;
        RECT 262.000 339.700 267.600 340.300 ;
        RECT 262.000 339.600 262.800 339.700 ;
        RECT 266.800 339.600 267.600 339.700 ;
        RECT 308.400 340.300 309.200 340.400 ;
        RECT 311.600 340.300 312.400 340.400 ;
        RECT 308.400 339.700 312.400 340.300 ;
        RECT 308.400 339.600 309.200 339.700 ;
        RECT 311.600 339.600 312.400 339.700 ;
        RECT 313.200 340.300 314.000 340.400 ;
        RECT 332.400 340.300 333.200 340.400 ;
        RECT 356.400 340.300 357.200 340.400 ;
        RECT 313.200 339.700 357.200 340.300 ;
        RECT 313.200 339.600 314.000 339.700 ;
        RECT 332.400 339.600 333.200 339.700 ;
        RECT 356.400 339.600 357.200 339.700 ;
        RECT 375.600 340.300 376.400 340.400 ;
        RECT 391.600 340.300 392.400 340.400 ;
        RECT 375.600 339.700 392.400 340.300 ;
        RECT 375.600 339.600 376.400 339.700 ;
        RECT 391.600 339.600 392.400 339.700 ;
        RECT 393.200 340.300 394.000 340.400 ;
        RECT 396.400 340.300 397.200 340.400 ;
        RECT 393.200 339.700 397.200 340.300 ;
        RECT 393.200 339.600 394.000 339.700 ;
        RECT 396.400 339.600 397.200 339.700 ;
        RECT 418.800 340.300 419.600 340.400 ;
        RECT 449.200 340.300 450.000 340.400 ;
        RECT 450.800 340.300 451.600 340.400 ;
        RECT 470.000 340.300 470.800 340.400 ;
        RECT 418.800 339.700 470.800 340.300 ;
        RECT 418.800 339.600 419.600 339.700 ;
        RECT 449.200 339.600 450.000 339.700 ;
        RECT 450.800 339.600 451.600 339.700 ;
        RECT 470.000 339.600 470.800 339.700 ;
        RECT 530.800 340.300 531.600 340.400 ;
        RECT 537.200 340.300 538.000 340.400 ;
        RECT 566.000 340.300 566.800 340.400 ;
        RECT 530.800 339.700 566.800 340.300 ;
        RECT 530.800 339.600 531.600 339.700 ;
        RECT 537.200 339.600 538.000 339.700 ;
        RECT 566.000 339.600 566.800 339.700 ;
        RECT 78.000 338.300 78.800 338.400 ;
        RECT 81.200 338.300 82.000 338.400 ;
        RECT 78.000 337.700 82.000 338.300 ;
        RECT 78.000 337.600 78.800 337.700 ;
        RECT 81.200 337.600 82.000 337.700 ;
        RECT 102.000 338.300 102.800 338.400 ;
        RECT 108.400 338.300 109.200 338.400 ;
        RECT 102.000 337.700 109.200 338.300 ;
        RECT 102.000 337.600 102.800 337.700 ;
        RECT 108.400 337.600 109.200 337.700 ;
        RECT 113.200 338.300 114.000 338.400 ;
        RECT 124.400 338.300 125.200 338.400 ;
        RECT 113.200 337.700 125.200 338.300 ;
        RECT 113.200 337.600 114.000 337.700 ;
        RECT 124.400 337.600 125.200 337.700 ;
        RECT 140.400 338.300 141.200 338.400 ;
        RECT 162.800 338.300 163.600 338.400 ;
        RECT 172.400 338.300 173.200 338.400 ;
        RECT 140.400 337.700 173.200 338.300 ;
        RECT 140.400 337.600 141.200 337.700 ;
        RECT 162.800 337.600 163.600 337.700 ;
        RECT 172.400 337.600 173.200 337.700 ;
        RECT 206.000 338.300 206.800 338.400 ;
        RECT 218.800 338.300 219.600 338.400 ;
        RECT 233.200 338.300 234.000 338.400 ;
        RECT 206.000 337.700 234.000 338.300 ;
        RECT 206.000 337.600 206.800 337.700 ;
        RECT 218.800 337.600 219.600 337.700 ;
        RECT 233.200 337.600 234.000 337.700 ;
        RECT 241.200 338.300 242.000 338.400 ;
        RECT 250.800 338.300 251.600 338.400 ;
        RECT 241.200 337.700 251.600 338.300 ;
        RECT 241.200 337.600 242.000 337.700 ;
        RECT 250.800 337.600 251.600 337.700 ;
        RECT 254.000 338.300 254.800 338.400 ;
        RECT 270.000 338.300 270.800 338.400 ;
        RECT 254.000 337.700 270.800 338.300 ;
        RECT 254.000 337.600 254.800 337.700 ;
        RECT 270.000 337.600 270.800 337.700 ;
        RECT 282.800 338.300 283.600 338.400 ;
        RECT 314.800 338.300 315.600 338.400 ;
        RECT 282.800 337.700 315.600 338.300 ;
        RECT 282.800 337.600 283.600 337.700 ;
        RECT 314.800 337.600 315.600 337.700 ;
        RECT 407.600 338.300 408.400 338.400 ;
        RECT 473.200 338.300 474.000 338.400 ;
        RECT 407.600 337.700 474.000 338.300 ;
        RECT 407.600 337.600 408.400 337.700 ;
        RECT 473.200 337.600 474.000 337.700 ;
        RECT 511.600 338.300 512.400 338.400 ;
        RECT 513.200 338.300 514.000 338.400 ;
        RECT 511.600 337.700 514.000 338.300 ;
        RECT 511.600 337.600 512.400 337.700 ;
        RECT 513.200 337.600 514.000 337.700 ;
        RECT 10.800 336.300 11.600 336.400 ;
        RECT 25.200 336.300 26.000 336.400 ;
        RECT 10.800 335.700 26.000 336.300 ;
        RECT 10.800 335.600 11.600 335.700 ;
        RECT 25.200 335.600 26.000 335.700 ;
        RECT 26.800 336.300 27.600 336.400 ;
        RECT 31.600 336.300 32.400 336.400 ;
        RECT 26.800 335.700 32.400 336.300 ;
        RECT 26.800 335.600 27.600 335.700 ;
        RECT 31.600 335.600 32.400 335.700 ;
        RECT 71.600 336.300 72.400 336.400 ;
        RECT 81.200 336.300 82.000 336.400 ;
        RECT 89.200 336.300 90.000 336.400 ;
        RECT 71.600 335.700 90.000 336.300 ;
        RECT 71.600 335.600 72.400 335.700 ;
        RECT 81.200 335.600 82.000 335.700 ;
        RECT 89.200 335.600 90.000 335.700 ;
        RECT 95.600 336.300 96.400 336.400 ;
        RECT 102.000 336.300 102.800 336.400 ;
        RECT 95.600 335.700 102.800 336.300 ;
        RECT 95.600 335.600 96.400 335.700 ;
        RECT 102.000 335.600 102.800 335.700 ;
        RECT 103.600 336.300 104.400 336.400 ;
        RECT 118.000 336.300 118.800 336.400 ;
        RECT 159.600 336.300 160.400 336.400 ;
        RECT 164.400 336.300 165.200 336.400 ;
        RECT 103.600 335.700 118.800 336.300 ;
        RECT 103.600 335.600 104.400 335.700 ;
        RECT 118.000 335.600 118.800 335.700 ;
        RECT 124.500 335.700 165.200 336.300 ;
        RECT 31.600 334.300 32.400 334.400 ;
        RECT 41.200 334.300 42.000 334.400 ;
        RECT 31.600 333.700 42.000 334.300 ;
        RECT 31.600 333.600 32.400 333.700 ;
        RECT 41.200 333.600 42.000 333.700 ;
        RECT 89.200 334.300 90.000 334.400 ;
        RECT 97.200 334.300 98.000 334.400 ;
        RECT 89.200 333.700 98.000 334.300 ;
        RECT 89.200 333.600 90.000 333.700 ;
        RECT 97.200 333.600 98.000 333.700 ;
        RECT 106.800 334.300 107.600 334.400 ;
        RECT 124.500 334.300 125.100 335.700 ;
        RECT 159.600 335.600 160.400 335.700 ;
        RECT 164.400 335.600 165.200 335.700 ;
        RECT 239.600 336.300 240.400 336.400 ;
        RECT 242.800 336.300 243.600 336.400 ;
        RECT 246.000 336.300 246.800 336.400 ;
        RECT 254.000 336.300 254.800 336.400 ;
        RECT 239.600 335.700 254.800 336.300 ;
        RECT 239.600 335.600 240.400 335.700 ;
        RECT 242.800 335.600 243.600 335.700 ;
        RECT 246.000 335.600 246.800 335.700 ;
        RECT 254.000 335.600 254.800 335.700 ;
        RECT 263.600 336.300 264.400 336.400 ;
        RECT 268.400 336.300 269.200 336.400 ;
        RECT 263.600 335.700 269.200 336.300 ;
        RECT 263.600 335.600 264.400 335.700 ;
        RECT 268.400 335.600 269.200 335.700 ;
        RECT 273.200 336.300 274.000 336.400 ;
        RECT 281.200 336.300 282.000 336.400 ;
        RECT 273.200 335.700 282.000 336.300 ;
        RECT 273.200 335.600 274.000 335.700 ;
        RECT 281.200 335.600 282.000 335.700 ;
        RECT 284.400 336.300 285.200 336.400 ;
        RECT 302.000 336.300 302.800 336.400 ;
        RECT 284.400 335.700 302.800 336.300 ;
        RECT 284.400 335.600 285.200 335.700 ;
        RECT 302.000 335.600 302.800 335.700 ;
        RECT 306.800 336.300 307.600 336.400 ;
        RECT 311.600 336.300 312.400 336.400 ;
        RECT 319.600 336.300 320.400 336.400 ;
        RECT 306.800 335.700 310.700 336.300 ;
        RECT 306.800 335.600 307.600 335.700 ;
        RECT 106.800 333.700 125.100 334.300 ;
        RECT 126.000 334.300 126.800 334.400 ;
        RECT 130.800 334.300 131.600 334.400 ;
        RECT 126.000 333.700 131.600 334.300 ;
        RECT 106.800 333.600 107.600 333.700 ;
        RECT 126.000 333.600 126.800 333.700 ;
        RECT 130.800 333.600 131.600 333.700 ;
        RECT 134.000 334.300 134.800 334.400 ;
        RECT 143.600 334.300 144.400 334.400 ;
        RECT 134.000 333.700 144.400 334.300 ;
        RECT 134.000 333.600 134.800 333.700 ;
        RECT 143.600 333.600 144.400 333.700 ;
        RECT 156.400 334.300 157.200 334.400 ;
        RECT 159.600 334.300 160.400 334.400 ;
        RECT 156.400 333.700 160.400 334.300 ;
        RECT 156.400 333.600 157.200 333.700 ;
        RECT 159.600 333.600 160.400 333.700 ;
        RECT 244.400 334.300 245.200 334.400 ;
        RECT 265.200 334.300 266.000 334.400 ;
        RECT 273.200 334.300 274.000 334.400 ;
        RECT 244.400 333.700 274.000 334.300 ;
        RECT 244.400 333.600 245.200 333.700 ;
        RECT 265.200 333.600 266.000 333.700 ;
        RECT 273.200 333.600 274.000 333.700 ;
        RECT 276.400 334.300 277.200 334.400 ;
        RECT 300.400 334.300 301.200 334.400 ;
        RECT 306.800 334.300 307.600 334.400 ;
        RECT 276.400 333.700 307.600 334.300 ;
        RECT 310.100 334.300 310.700 335.700 ;
        RECT 311.600 335.700 320.400 336.300 ;
        RECT 311.600 335.600 312.400 335.700 ;
        RECT 319.600 335.600 320.400 335.700 ;
        RECT 386.800 336.300 387.600 336.400 ;
        RECT 390.000 336.300 390.800 336.400 ;
        RECT 463.600 336.300 464.400 336.400 ;
        RECT 386.800 335.700 390.800 336.300 ;
        RECT 386.800 335.600 387.600 335.700 ;
        RECT 390.000 335.600 390.800 335.700 ;
        RECT 454.100 335.700 464.400 336.300 ;
        RECT 454.100 334.400 454.700 335.700 ;
        RECT 463.600 335.600 464.400 335.700 ;
        RECT 540.400 336.300 541.200 336.400 ;
        RECT 550.000 336.300 550.800 336.400 ;
        RECT 540.400 335.700 550.800 336.300 ;
        RECT 540.400 335.600 541.200 335.700 ;
        RECT 550.000 335.600 550.800 335.700 ;
        RECT 322.800 334.300 323.600 334.400 ;
        RECT 310.100 333.700 323.600 334.300 ;
        RECT 276.400 333.600 277.200 333.700 ;
        RECT 300.400 333.600 301.200 333.700 ;
        RECT 306.800 333.600 307.600 333.700 ;
        RECT 322.800 333.600 323.600 333.700 ;
        RECT 382.000 334.300 382.800 334.400 ;
        RECT 386.800 334.300 387.600 334.400 ;
        RECT 382.000 333.700 387.600 334.300 ;
        RECT 382.000 333.600 382.800 333.700 ;
        RECT 386.800 333.600 387.600 333.700 ;
        RECT 410.800 334.300 411.600 334.400 ;
        RECT 423.600 334.300 424.400 334.400 ;
        RECT 410.800 333.700 424.400 334.300 ;
        RECT 410.800 333.600 411.600 333.700 ;
        RECT 423.600 333.600 424.400 333.700 ;
        RECT 430.000 334.300 430.800 334.400 ;
        RECT 433.200 334.300 434.000 334.400 ;
        RECT 430.000 333.700 434.000 334.300 ;
        RECT 430.000 333.600 430.800 333.700 ;
        RECT 433.200 333.600 434.000 333.700 ;
        RECT 438.000 334.300 438.800 334.400 ;
        RECT 447.600 334.300 448.400 334.400 ;
        RECT 454.000 334.300 454.800 334.400 ;
        RECT 438.000 333.700 454.800 334.300 ;
        RECT 438.000 333.600 438.800 333.700 ;
        RECT 447.600 333.600 448.400 333.700 ;
        RECT 454.000 333.600 454.800 333.700 ;
        RECT 460.400 333.600 461.200 334.400 ;
        RECT 537.200 334.300 538.000 334.400 ;
        RECT 553.200 334.300 554.000 334.400 ;
        RECT 537.200 333.700 554.000 334.300 ;
        RECT 537.200 333.600 538.000 333.700 ;
        RECT 553.200 333.600 554.000 333.700 ;
        RECT 14.000 332.300 14.800 332.400 ;
        RECT 25.200 332.300 26.000 332.400 ;
        RECT 30.000 332.300 30.800 332.400 ;
        RECT 14.000 331.700 30.800 332.300 ;
        RECT 14.000 331.600 14.800 331.700 ;
        RECT 25.200 331.600 26.000 331.700 ;
        RECT 30.000 331.600 30.800 331.700 ;
        RECT 57.200 332.300 58.000 332.400 ;
        RECT 70.000 332.300 70.800 332.400 ;
        RECT 57.200 331.700 70.800 332.300 ;
        RECT 57.200 331.600 58.000 331.700 ;
        RECT 70.000 331.600 70.800 331.700 ;
        RECT 84.400 332.300 85.200 332.400 ;
        RECT 89.200 332.300 90.000 332.400 ;
        RECT 94.000 332.300 94.800 332.400 ;
        RECT 84.400 331.700 94.800 332.300 ;
        RECT 84.400 331.600 85.200 331.700 ;
        RECT 89.200 331.600 90.000 331.700 ;
        RECT 94.000 331.600 94.800 331.700 ;
        RECT 95.600 332.300 96.400 332.400 ;
        RECT 102.000 332.300 102.800 332.400 ;
        RECT 95.600 331.700 102.800 332.300 ;
        RECT 95.600 331.600 96.400 331.700 ;
        RECT 102.000 331.600 102.800 331.700 ;
        RECT 110.000 332.300 110.800 332.400 ;
        RECT 113.200 332.300 114.000 332.400 ;
        RECT 110.000 331.700 114.000 332.300 ;
        RECT 110.000 331.600 110.800 331.700 ;
        RECT 113.200 331.600 114.000 331.700 ;
        RECT 130.800 332.300 131.600 332.400 ;
        RECT 137.200 332.300 138.000 332.400 ;
        RECT 130.800 331.700 138.000 332.300 ;
        RECT 130.800 331.600 131.600 331.700 ;
        RECT 137.200 331.600 138.000 331.700 ;
        RECT 138.800 332.300 139.600 332.400 ;
        RECT 156.500 332.300 157.100 333.600 ;
        RECT 138.800 331.700 157.100 332.300 ;
        RECT 212.400 332.300 213.200 332.400 ;
        RECT 218.800 332.300 219.600 332.400 ;
        RECT 212.400 331.700 219.600 332.300 ;
        RECT 138.800 331.600 139.600 331.700 ;
        RECT 212.400 331.600 213.200 331.700 ;
        RECT 218.800 331.600 219.600 331.700 ;
        RECT 234.800 332.300 235.600 332.400 ;
        RECT 250.800 332.300 251.600 332.400 ;
        RECT 234.800 331.700 251.600 332.300 ;
        RECT 234.800 331.600 235.600 331.700 ;
        RECT 250.800 331.600 251.600 331.700 ;
        RECT 252.400 332.300 253.200 332.400 ;
        RECT 263.600 332.300 264.400 332.400 ;
        RECT 252.400 331.700 264.400 332.300 ;
        RECT 252.400 331.600 253.200 331.700 ;
        RECT 263.600 331.600 264.400 331.700 ;
        RECT 274.800 332.300 275.600 332.400 ;
        RECT 295.600 332.300 296.400 332.400 ;
        RECT 274.800 331.700 296.400 332.300 ;
        RECT 274.800 331.600 275.600 331.700 ;
        RECT 295.600 331.600 296.400 331.700 ;
        RECT 346.800 332.300 347.600 332.400 ;
        RECT 353.200 332.300 354.000 332.400 ;
        RECT 346.800 331.700 354.000 332.300 ;
        RECT 346.800 331.600 347.600 331.700 ;
        RECT 353.200 331.600 354.000 331.700 ;
        RECT 354.800 332.300 355.600 332.400 ;
        RECT 369.200 332.300 370.000 332.400 ;
        RECT 383.600 332.300 384.400 332.400 ;
        RECT 354.800 331.700 384.400 332.300 ;
        RECT 354.800 331.600 355.600 331.700 ;
        RECT 369.200 331.600 370.000 331.700 ;
        RECT 383.600 331.600 384.400 331.700 ;
        RECT 426.800 332.300 427.600 332.400 ;
        RECT 436.400 332.300 437.200 332.400 ;
        RECT 426.800 331.700 437.200 332.300 ;
        RECT 426.800 331.600 427.600 331.700 ;
        RECT 436.400 331.600 437.200 331.700 ;
        RECT 455.600 332.300 456.400 332.400 ;
        RECT 460.400 332.300 461.200 332.400 ;
        RECT 455.600 331.700 461.200 332.300 ;
        RECT 455.600 331.600 456.400 331.700 ;
        RECT 460.400 331.600 461.200 331.700 ;
        RECT 506.800 332.300 507.600 332.400 ;
        RECT 511.600 332.300 512.400 332.400 ;
        RECT 506.800 331.700 512.400 332.300 ;
        RECT 506.800 331.600 507.600 331.700 ;
        RECT 511.600 331.600 512.400 331.700 ;
        RECT 566.000 331.600 566.800 332.400 ;
        RECT 28.400 330.300 29.200 330.400 ;
        RECT 36.400 330.300 37.200 330.400 ;
        RECT 28.400 329.700 37.200 330.300 ;
        RECT 28.400 329.600 29.200 329.700 ;
        RECT 36.400 329.600 37.200 329.700 ;
        RECT 54.000 330.300 54.800 330.400 ;
        RECT 60.400 330.300 61.200 330.400 ;
        RECT 54.000 329.700 61.200 330.300 ;
        RECT 54.000 329.600 54.800 329.700 ;
        RECT 60.400 329.600 61.200 329.700 ;
        RECT 71.600 330.300 72.400 330.400 ;
        RECT 74.800 330.300 75.600 330.400 ;
        RECT 71.600 329.700 75.600 330.300 ;
        RECT 71.600 329.600 72.400 329.700 ;
        RECT 74.800 329.600 75.600 329.700 ;
        RECT 113.200 330.300 114.000 330.400 ;
        RECT 119.600 330.300 120.400 330.400 ;
        RECT 113.200 329.700 120.400 330.300 ;
        RECT 113.200 329.600 114.000 329.700 ;
        RECT 119.600 329.600 120.400 329.700 ;
        RECT 239.600 330.300 240.400 330.400 ;
        RECT 255.600 330.300 256.400 330.400 ;
        RECT 239.600 329.700 256.400 330.300 ;
        RECT 239.600 329.600 240.400 329.700 ;
        RECT 255.600 329.600 256.400 329.700 ;
        RECT 266.800 330.300 267.600 330.400 ;
        RECT 276.400 330.300 277.200 330.400 ;
        RECT 266.800 329.700 277.200 330.300 ;
        RECT 266.800 329.600 267.600 329.700 ;
        RECT 276.400 329.600 277.200 329.700 ;
        RECT 279.600 330.300 280.400 330.400 ;
        RECT 310.000 330.300 310.800 330.400 ;
        RECT 279.600 329.700 310.800 330.300 ;
        RECT 279.600 329.600 280.400 329.700 ;
        RECT 310.000 329.600 310.800 329.700 ;
        RECT 378.800 330.300 379.600 330.400 ;
        RECT 383.600 330.300 384.400 330.400 ;
        RECT 378.800 329.700 384.400 330.300 ;
        RECT 378.800 329.600 379.600 329.700 ;
        RECT 383.600 329.600 384.400 329.700 ;
        RECT 468.400 330.300 469.200 330.400 ;
        RECT 474.800 330.300 475.600 330.400 ;
        RECT 468.400 329.700 475.600 330.300 ;
        RECT 468.400 329.600 469.200 329.700 ;
        RECT 474.800 329.600 475.600 329.700 ;
        RECT 47.600 328.300 48.400 328.400 ;
        RECT 52.400 328.300 53.200 328.400 ;
        RECT 47.600 327.700 53.200 328.300 ;
        RECT 47.600 327.600 48.400 327.700 ;
        RECT 52.400 327.600 53.200 327.700 ;
        RECT 65.200 328.300 66.000 328.400 ;
        RECT 70.000 328.300 70.800 328.400 ;
        RECT 65.200 327.700 70.800 328.300 ;
        RECT 65.200 327.600 66.000 327.700 ;
        RECT 70.000 327.600 70.800 327.700 ;
        RECT 228.400 328.300 229.200 328.400 ;
        RECT 302.000 328.300 302.800 328.400 ;
        RECT 228.400 327.700 302.800 328.300 ;
        RECT 228.400 327.600 229.200 327.700 ;
        RECT 302.000 327.600 302.800 327.700 ;
        RECT 351.600 328.300 352.400 328.400 ;
        RECT 377.200 328.300 378.000 328.400 ;
        RECT 351.600 327.700 378.000 328.300 ;
        RECT 351.600 327.600 352.400 327.700 ;
        RECT 377.200 327.600 378.000 327.700 ;
        RECT 463.600 327.600 464.400 328.400 ;
        RECT 41.200 326.300 42.000 326.400 ;
        RECT 66.800 326.300 67.600 326.400 ;
        RECT 81.200 326.300 82.000 326.400 ;
        RECT 41.200 325.700 82.000 326.300 ;
        RECT 41.200 325.600 42.000 325.700 ;
        RECT 66.800 325.600 67.600 325.700 ;
        RECT 81.200 325.600 82.000 325.700 ;
        RECT 255.600 326.300 256.400 326.400 ;
        RECT 276.400 326.300 277.200 326.400 ;
        RECT 255.600 325.700 277.200 326.300 ;
        RECT 255.600 325.600 256.400 325.700 ;
        RECT 276.400 325.600 277.200 325.700 ;
        RECT 426.800 326.300 427.600 326.400 ;
        RECT 457.200 326.300 458.000 326.400 ;
        RECT 476.400 326.300 477.200 326.400 ;
        RECT 426.800 325.700 477.200 326.300 ;
        RECT 426.800 325.600 427.600 325.700 ;
        RECT 457.200 325.600 458.000 325.700 ;
        RECT 476.400 325.600 477.200 325.700 ;
        RECT 7.600 324.300 8.400 324.400 ;
        RECT 26.800 324.300 27.600 324.400 ;
        RECT 7.600 323.700 27.600 324.300 ;
        RECT 7.600 323.600 8.400 323.700 ;
        RECT 26.800 323.600 27.600 323.700 ;
        RECT 146.800 323.600 147.600 324.400 ;
        RECT 172.400 324.300 173.200 324.400 ;
        RECT 199.600 324.300 200.400 324.400 ;
        RECT 172.400 323.700 200.400 324.300 ;
        RECT 172.400 323.600 173.200 323.700 ;
        RECT 199.600 323.600 200.400 323.700 ;
        RECT 380.400 324.300 381.200 324.400 ;
        RECT 388.400 324.300 389.200 324.400 ;
        RECT 391.600 324.300 392.400 324.400 ;
        RECT 380.400 323.700 392.400 324.300 ;
        RECT 380.400 323.600 381.200 323.700 ;
        RECT 388.400 323.600 389.200 323.700 ;
        RECT 391.600 323.600 392.400 323.700 ;
        RECT 553.200 324.300 554.000 324.400 ;
        RECT 554.800 324.300 555.600 324.400 ;
        RECT 553.200 323.700 555.600 324.300 ;
        RECT 553.200 323.600 554.000 323.700 ;
        RECT 554.800 323.600 555.600 323.700 ;
        RECT 382.000 322.300 382.800 322.400 ;
        RECT 390.000 322.300 390.800 322.400 ;
        RECT 394.800 322.300 395.600 322.400 ;
        RECT 382.000 321.700 395.600 322.300 ;
        RECT 382.000 321.600 382.800 321.700 ;
        RECT 390.000 321.600 390.800 321.700 ;
        RECT 394.800 321.600 395.600 321.700 ;
        RECT 74.800 320.300 75.600 320.400 ;
        RECT 79.600 320.300 80.400 320.400 ;
        RECT 122.800 320.300 123.600 320.400 ;
        RECT 130.800 320.300 131.600 320.400 ;
        RECT 74.800 319.700 131.600 320.300 ;
        RECT 74.800 319.600 75.600 319.700 ;
        RECT 79.600 319.600 80.400 319.700 ;
        RECT 122.800 319.600 123.600 319.700 ;
        RECT 130.800 319.600 131.600 319.700 ;
        RECT 212.400 320.300 213.200 320.400 ;
        RECT 326.000 320.300 326.800 320.400 ;
        RECT 212.400 319.700 326.800 320.300 ;
        RECT 212.400 319.600 213.200 319.700 ;
        RECT 326.000 319.600 326.800 319.700 ;
        RECT 47.600 318.300 48.400 318.400 ;
        RECT 52.400 318.300 53.200 318.400 ;
        RECT 47.600 317.700 53.200 318.300 ;
        RECT 47.600 317.600 48.400 317.700 ;
        RECT 52.400 317.600 53.200 317.700 ;
        RECT 233.200 318.300 234.000 318.400 ;
        RECT 234.800 318.300 235.600 318.400 ;
        RECT 268.400 318.300 269.200 318.400 ;
        RECT 273.200 318.300 274.000 318.400 ;
        RECT 233.200 317.700 274.000 318.300 ;
        RECT 233.200 317.600 234.000 317.700 ;
        RECT 234.800 317.600 235.600 317.700 ;
        RECT 268.400 317.600 269.200 317.700 ;
        RECT 273.200 317.600 274.000 317.700 ;
        RECT 364.400 318.300 365.200 318.400 ;
        RECT 385.200 318.300 386.000 318.400 ;
        RECT 364.400 317.700 386.000 318.300 ;
        RECT 364.400 317.600 365.200 317.700 ;
        RECT 385.200 317.600 386.000 317.700 ;
        RECT 417.200 318.300 418.000 318.400 ;
        RECT 468.400 318.300 469.200 318.400 ;
        RECT 417.200 317.700 469.200 318.300 ;
        RECT 417.200 317.600 418.000 317.700 ;
        RECT 468.400 317.600 469.200 317.700 ;
        RECT 497.200 318.300 498.000 318.400 ;
        RECT 500.400 318.300 501.200 318.400 ;
        RECT 497.200 317.700 501.200 318.300 ;
        RECT 497.200 317.600 498.000 317.700 ;
        RECT 500.400 317.600 501.200 317.700 ;
        RECT 68.400 316.300 69.200 316.400 ;
        RECT 90.800 316.300 91.600 316.400 ;
        RECT 68.400 315.700 91.600 316.300 ;
        RECT 68.400 315.600 69.200 315.700 ;
        RECT 90.800 315.600 91.600 315.700 ;
        RECT 127.600 315.600 128.400 316.400 ;
        RECT 228.400 316.300 229.200 316.400 ;
        RECT 260.400 316.300 261.200 316.400 ;
        RECT 228.400 315.700 261.200 316.300 ;
        RECT 228.400 315.600 229.200 315.700 ;
        RECT 260.400 315.600 261.200 315.700 ;
        RECT 337.200 316.300 338.000 316.400 ;
        RECT 342.000 316.300 342.800 316.400 ;
        RECT 377.200 316.300 378.000 316.400 ;
        RECT 337.200 315.700 378.000 316.300 ;
        RECT 337.200 315.600 338.000 315.700 ;
        RECT 342.000 315.600 342.800 315.700 ;
        RECT 377.200 315.600 378.000 315.700 ;
        RECT 412.400 316.300 413.200 316.400 ;
        RECT 428.400 316.300 429.200 316.400 ;
        RECT 412.400 315.700 429.200 316.300 ;
        RECT 412.400 315.600 413.200 315.700 ;
        RECT 428.400 315.600 429.200 315.700 ;
        RECT 1.200 314.300 2.000 314.400 ;
        RECT 18.800 314.300 19.600 314.400 ;
        RECT 1.200 313.700 19.600 314.300 ;
        RECT 1.200 313.600 2.000 313.700 ;
        RECT 18.800 313.600 19.600 313.700 ;
        RECT 20.400 314.300 21.200 314.400 ;
        RECT 31.600 314.300 32.400 314.400 ;
        RECT 20.400 313.700 32.400 314.300 ;
        RECT 20.400 313.600 21.200 313.700 ;
        RECT 31.600 313.600 32.400 313.700 ;
        RECT 41.200 314.300 42.000 314.400 ;
        RECT 44.400 314.300 45.200 314.400 ;
        RECT 41.200 313.700 45.200 314.300 ;
        RECT 41.200 313.600 42.000 313.700 ;
        RECT 44.400 313.600 45.200 313.700 ;
        RECT 54.000 314.300 54.800 314.400 ;
        RECT 63.600 314.300 64.400 314.400 ;
        RECT 54.000 313.700 64.400 314.300 ;
        RECT 54.000 313.600 54.800 313.700 ;
        RECT 63.600 313.600 64.400 313.700 ;
        RECT 66.800 314.300 67.600 314.400 ;
        RECT 73.200 314.300 74.000 314.400 ;
        RECT 66.800 313.700 74.000 314.300 ;
        RECT 66.800 313.600 67.600 313.700 ;
        RECT 73.200 313.600 74.000 313.700 ;
        RECT 119.600 314.300 120.400 314.400 ;
        RECT 137.200 314.300 138.000 314.400 ;
        RECT 119.600 313.700 138.000 314.300 ;
        RECT 119.600 313.600 120.400 313.700 ;
        RECT 137.200 313.600 138.000 313.700 ;
        RECT 241.200 314.300 242.000 314.400 ;
        RECT 244.400 314.300 245.200 314.400 ;
        RECT 241.200 313.700 245.200 314.300 ;
        RECT 241.200 313.600 242.000 313.700 ;
        RECT 244.400 313.600 245.200 313.700 ;
        RECT 249.200 314.300 250.000 314.400 ;
        RECT 263.600 314.300 264.400 314.400 ;
        RECT 289.200 314.300 290.000 314.400 ;
        RECT 249.200 313.700 290.000 314.300 ;
        RECT 249.200 313.600 250.000 313.700 ;
        RECT 263.600 313.600 264.400 313.700 ;
        RECT 289.200 313.600 290.000 313.700 ;
        RECT 310.000 314.300 310.800 314.400 ;
        RECT 353.200 314.300 354.000 314.400 ;
        RECT 310.000 313.700 354.000 314.300 ;
        RECT 310.000 313.600 310.800 313.700 ;
        RECT 353.200 313.600 354.000 313.700 ;
        RECT 354.800 314.300 355.600 314.400 ;
        RECT 404.400 314.300 405.200 314.400 ;
        RECT 354.800 313.700 405.200 314.300 ;
        RECT 354.800 313.600 355.600 313.700 ;
        RECT 404.400 313.600 405.200 313.700 ;
        RECT 444.400 314.300 445.200 314.400 ;
        RECT 458.800 314.300 459.600 314.400 ;
        RECT 460.400 314.300 461.200 314.400 ;
        RECT 444.400 313.700 461.200 314.300 ;
        RECT 444.400 313.600 445.200 313.700 ;
        RECT 458.800 313.600 459.600 313.700 ;
        RECT 460.400 313.600 461.200 313.700 ;
        RECT 22.000 312.300 22.800 312.400 ;
        RECT 25.200 312.300 26.000 312.400 ;
        RECT 22.000 311.700 26.000 312.300 ;
        RECT 22.000 311.600 22.800 311.700 ;
        RECT 25.200 311.600 26.000 311.700 ;
        RECT 30.000 312.300 30.800 312.400 ;
        RECT 71.600 312.300 72.400 312.400 ;
        RECT 92.400 312.300 93.200 312.400 ;
        RECT 30.000 311.700 93.200 312.300 ;
        RECT 30.000 311.600 30.800 311.700 ;
        RECT 71.600 311.600 72.400 311.700 ;
        RECT 92.400 311.600 93.200 311.700 ;
        RECT 124.400 312.300 125.200 312.400 ;
        RECT 127.600 312.300 128.400 312.400 ;
        RECT 124.400 311.700 128.400 312.300 ;
        RECT 124.400 311.600 125.200 311.700 ;
        RECT 127.600 311.600 128.400 311.700 ;
        RECT 143.600 312.300 144.400 312.400 ;
        RECT 151.600 312.300 152.400 312.400 ;
        RECT 143.600 311.700 152.400 312.300 ;
        RECT 143.600 311.600 144.400 311.700 ;
        RECT 151.600 311.600 152.400 311.700 ;
        RECT 153.200 312.300 154.000 312.400 ;
        RECT 167.600 312.300 168.400 312.400 ;
        RECT 153.200 311.700 168.400 312.300 ;
        RECT 153.200 311.600 154.000 311.700 ;
        RECT 167.600 311.600 168.400 311.700 ;
        RECT 193.200 312.300 194.000 312.400 ;
        RECT 231.600 312.300 232.400 312.400 ;
        RECT 193.200 311.700 232.400 312.300 ;
        RECT 193.200 311.600 194.000 311.700 ;
        RECT 231.600 311.600 232.400 311.700 ;
        RECT 244.400 312.300 245.200 312.400 ;
        RECT 247.600 312.300 248.400 312.400 ;
        RECT 244.400 311.700 248.400 312.300 ;
        RECT 244.400 311.600 245.200 311.700 ;
        RECT 247.600 311.600 248.400 311.700 ;
        RECT 271.600 312.300 272.400 312.400 ;
        RECT 316.400 312.300 317.200 312.400 ;
        RECT 271.600 311.700 317.200 312.300 ;
        RECT 271.600 311.600 272.400 311.700 ;
        RECT 316.400 311.600 317.200 311.700 ;
        RECT 322.800 312.300 323.600 312.400 ;
        RECT 330.800 312.300 331.600 312.400 ;
        RECT 322.800 311.700 331.600 312.300 ;
        RECT 322.800 311.600 323.600 311.700 ;
        RECT 330.800 311.600 331.600 311.700 ;
        RECT 338.800 312.300 339.600 312.400 ;
        RECT 343.600 312.300 344.400 312.400 ;
        RECT 338.800 311.700 344.400 312.300 ;
        RECT 338.800 311.600 339.600 311.700 ;
        RECT 343.600 311.600 344.400 311.700 ;
        RECT 345.200 312.300 346.000 312.400 ;
        RECT 375.600 312.300 376.400 312.400 ;
        RECT 345.200 311.700 376.400 312.300 ;
        RECT 345.200 311.600 346.000 311.700 ;
        RECT 375.600 311.600 376.400 311.700 ;
        RECT 425.200 312.300 426.000 312.400 ;
        RECT 434.800 312.300 435.600 312.400 ;
        RECT 425.200 311.700 435.600 312.300 ;
        RECT 425.200 311.600 426.000 311.700 ;
        RECT 434.800 311.600 435.600 311.700 ;
        RECT 438.000 312.300 438.800 312.400 ;
        RECT 454.000 312.300 454.800 312.400 ;
        RECT 438.000 311.700 454.800 312.300 ;
        RECT 438.000 311.600 438.800 311.700 ;
        RECT 454.000 311.600 454.800 311.700 ;
        RECT 529.200 312.300 530.000 312.400 ;
        RECT 535.600 312.300 536.400 312.400 ;
        RECT 529.200 311.700 536.400 312.300 ;
        RECT 529.200 311.600 530.000 311.700 ;
        RECT 535.600 311.600 536.400 311.700 ;
        RECT 562.800 312.300 563.600 312.400 ;
        RECT 569.200 312.300 570.000 312.400 ;
        RECT 562.800 311.700 570.000 312.300 ;
        RECT 562.800 311.600 563.600 311.700 ;
        RECT 569.200 311.600 570.000 311.700 ;
        RECT 12.400 309.600 13.200 310.400 ;
        RECT 20.400 310.300 21.200 310.400 ;
        RECT 36.400 310.300 37.200 310.400 ;
        RECT 20.400 309.700 37.200 310.300 ;
        RECT 20.400 309.600 21.200 309.700 ;
        RECT 36.400 309.600 37.200 309.700 ;
        RECT 49.200 310.300 50.000 310.400 ;
        RECT 89.200 310.300 90.000 310.400 ;
        RECT 95.600 310.300 96.400 310.400 ;
        RECT 49.200 309.700 80.300 310.300 ;
        RECT 49.200 309.600 50.000 309.700 ;
        RECT 79.700 308.400 80.300 309.700 ;
        RECT 89.200 309.700 96.400 310.300 ;
        RECT 89.200 309.600 90.000 309.700 ;
        RECT 95.600 309.600 96.400 309.700 ;
        RECT 106.800 310.300 107.600 310.400 ;
        RECT 132.400 310.300 133.200 310.400 ;
        RECT 106.800 309.700 133.200 310.300 ;
        RECT 106.800 309.600 107.600 309.700 ;
        RECT 132.400 309.600 133.200 309.700 ;
        RECT 134.000 310.300 134.800 310.400 ;
        RECT 150.000 310.300 150.800 310.400 ;
        RECT 169.200 310.300 170.000 310.400 ;
        RECT 175.600 310.300 176.400 310.400 ;
        RECT 199.600 310.300 200.400 310.400 ;
        RECT 134.000 309.700 200.400 310.300 ;
        RECT 134.000 309.600 134.800 309.700 ;
        RECT 150.000 309.600 150.800 309.700 ;
        RECT 169.200 309.600 170.000 309.700 ;
        RECT 175.600 309.600 176.400 309.700 ;
        RECT 199.600 309.600 200.400 309.700 ;
        RECT 231.600 310.300 232.400 310.400 ;
        RECT 242.800 310.300 243.600 310.400 ;
        RECT 231.600 309.700 243.600 310.300 ;
        RECT 231.600 309.600 232.400 309.700 ;
        RECT 242.800 309.600 243.600 309.700 ;
        RECT 246.000 310.300 246.800 310.400 ;
        RECT 250.800 310.300 251.600 310.400 ;
        RECT 246.000 309.700 251.600 310.300 ;
        RECT 246.000 309.600 246.800 309.700 ;
        RECT 250.800 309.600 251.600 309.700 ;
        RECT 286.000 310.300 286.800 310.400 ;
        RECT 327.600 310.300 328.400 310.400 ;
        RECT 335.600 310.300 336.400 310.400 ;
        RECT 286.000 309.700 336.400 310.300 ;
        RECT 286.000 309.600 286.800 309.700 ;
        RECT 327.600 309.600 328.400 309.700 ;
        RECT 335.600 309.600 336.400 309.700 ;
        RECT 348.400 310.300 349.200 310.400 ;
        RECT 380.400 310.300 381.200 310.400 ;
        RECT 348.400 309.700 381.200 310.300 ;
        RECT 348.400 309.600 349.200 309.700 ;
        RECT 380.400 309.600 381.200 309.700 ;
        RECT 385.200 310.300 386.000 310.400 ;
        RECT 388.400 310.300 389.200 310.400 ;
        RECT 396.400 310.300 397.200 310.400 ;
        RECT 385.200 309.700 397.200 310.300 ;
        RECT 385.200 309.600 386.000 309.700 ;
        RECT 388.400 309.600 389.200 309.700 ;
        RECT 396.400 309.600 397.200 309.700 ;
        RECT 430.000 310.300 430.800 310.400 ;
        RECT 439.600 310.300 440.400 310.400 ;
        RECT 430.000 309.700 440.400 310.300 ;
        RECT 430.000 309.600 430.800 309.700 ;
        RECT 439.600 309.600 440.400 309.700 ;
        RECT 457.200 310.300 458.000 310.400 ;
        RECT 474.800 310.300 475.600 310.400 ;
        RECT 457.200 309.700 475.600 310.300 ;
        RECT 457.200 309.600 458.000 309.700 ;
        RECT 474.800 309.600 475.600 309.700 ;
        RECT 481.200 310.300 482.000 310.400 ;
        RECT 484.400 310.300 485.200 310.400 ;
        RECT 481.200 309.700 485.200 310.300 ;
        RECT 481.200 309.600 482.000 309.700 ;
        RECT 484.400 309.600 485.200 309.700 ;
        RECT 529.200 310.300 530.000 310.400 ;
        RECT 537.200 310.300 538.000 310.400 ;
        RECT 529.200 309.700 538.000 310.300 ;
        RECT 529.200 309.600 530.000 309.700 ;
        RECT 537.200 309.600 538.000 309.700 ;
        RECT 4.400 308.300 5.200 308.400 ;
        RECT 10.800 308.300 11.600 308.400 ;
        RECT 17.200 308.300 18.000 308.400 ;
        RECT 30.000 308.300 30.800 308.400 ;
        RECT 4.400 307.700 30.800 308.300 ;
        RECT 4.400 307.600 5.200 307.700 ;
        RECT 10.800 307.600 11.600 307.700 ;
        RECT 17.200 307.600 18.000 307.700 ;
        RECT 30.000 307.600 30.800 307.700 ;
        RECT 33.200 308.300 34.000 308.400 ;
        RECT 41.200 308.300 42.000 308.400 ;
        RECT 50.800 308.300 51.600 308.400 ;
        RECT 33.200 307.700 51.600 308.300 ;
        RECT 33.200 307.600 34.000 307.700 ;
        RECT 41.200 307.600 42.000 307.700 ;
        RECT 50.800 307.600 51.600 307.700 ;
        RECT 60.400 308.300 61.200 308.400 ;
        RECT 76.400 308.300 77.200 308.400 ;
        RECT 60.400 307.700 77.200 308.300 ;
        RECT 60.400 307.600 61.200 307.700 ;
        RECT 76.400 307.600 77.200 307.700 ;
        RECT 79.600 307.600 80.400 308.400 ;
        RECT 84.400 308.300 85.200 308.400 ;
        RECT 97.200 308.300 98.000 308.400 ;
        RECT 103.600 308.300 104.400 308.400 ;
        RECT 84.400 307.700 104.400 308.300 ;
        RECT 84.400 307.600 85.200 307.700 ;
        RECT 97.200 307.600 98.000 307.700 ;
        RECT 103.600 307.600 104.400 307.700 ;
        RECT 130.800 308.300 131.600 308.400 ;
        RECT 145.200 308.300 146.000 308.400 ;
        RECT 130.800 307.700 146.000 308.300 ;
        RECT 130.800 307.600 131.600 307.700 ;
        RECT 145.200 307.600 146.000 307.700 ;
        RECT 153.200 308.300 154.000 308.400 ;
        RECT 156.400 308.300 157.200 308.400 ;
        RECT 153.200 307.700 157.200 308.300 ;
        RECT 153.200 307.600 154.000 307.700 ;
        RECT 156.400 307.600 157.200 307.700 ;
        RECT 158.000 308.300 158.800 308.400 ;
        RECT 161.200 308.300 162.000 308.400 ;
        RECT 158.000 307.700 162.000 308.300 ;
        RECT 158.000 307.600 158.800 307.700 ;
        RECT 161.200 307.600 162.000 307.700 ;
        RECT 230.000 308.300 230.800 308.400 ;
        RECT 239.600 308.300 240.400 308.400 ;
        RECT 252.400 308.300 253.200 308.400 ;
        RECT 230.000 307.700 253.200 308.300 ;
        RECT 230.000 307.600 230.800 307.700 ;
        RECT 239.600 307.600 240.400 307.700 ;
        RECT 252.400 307.600 253.200 307.700 ;
        RECT 292.400 308.300 293.200 308.400 ;
        RECT 303.600 308.300 304.400 308.400 ;
        RECT 292.400 307.700 304.400 308.300 ;
        RECT 292.400 307.600 293.200 307.700 ;
        RECT 303.600 307.600 304.400 307.700 ;
        RECT 330.800 308.300 331.600 308.400 ;
        RECT 338.800 308.300 339.600 308.400 ;
        RECT 330.800 307.700 339.600 308.300 ;
        RECT 330.800 307.600 331.600 307.700 ;
        RECT 338.800 307.600 339.600 307.700 ;
        RECT 366.000 308.300 366.800 308.400 ;
        RECT 366.000 307.700 384.300 308.300 ;
        RECT 366.000 307.600 366.800 307.700 ;
        RECT 12.400 306.300 13.200 306.400 ;
        RECT 15.600 306.300 16.400 306.400 ;
        RECT 20.400 306.300 21.200 306.400 ;
        RECT 12.400 305.700 21.200 306.300 ;
        RECT 12.400 305.600 13.200 305.700 ;
        RECT 15.600 305.600 16.400 305.700 ;
        RECT 20.400 305.600 21.200 305.700 ;
        RECT 23.600 306.300 24.400 306.400 ;
        RECT 28.400 306.300 29.200 306.400 ;
        RECT 23.600 305.700 29.200 306.300 ;
        RECT 23.600 305.600 24.400 305.700 ;
        RECT 28.400 305.600 29.200 305.700 ;
        RECT 34.800 306.300 35.600 306.400 ;
        RECT 39.600 306.300 40.400 306.400 ;
        RECT 34.800 305.700 40.400 306.300 ;
        RECT 34.800 305.600 35.600 305.700 ;
        RECT 39.600 305.600 40.400 305.700 ;
        RECT 82.800 306.300 83.600 306.400 ;
        RECT 84.400 306.300 85.200 306.400 ;
        RECT 87.600 306.300 88.400 306.400 ;
        RECT 82.800 305.700 88.400 306.300 ;
        RECT 82.800 305.600 83.600 305.700 ;
        RECT 84.400 305.600 85.200 305.700 ;
        RECT 87.600 305.600 88.400 305.700 ;
        RECT 92.400 306.300 93.200 306.400 ;
        RECT 100.400 306.300 101.200 306.400 ;
        RECT 102.000 306.300 102.800 306.400 ;
        RECT 105.200 306.300 106.000 306.400 ;
        RECT 146.800 306.300 147.600 306.400 ;
        RECT 172.400 306.300 173.200 306.400 ;
        RECT 92.400 305.700 173.200 306.300 ;
        RECT 92.400 305.600 93.200 305.700 ;
        RECT 100.400 305.600 101.200 305.700 ;
        RECT 102.000 305.600 102.800 305.700 ;
        RECT 105.200 305.600 106.000 305.700 ;
        RECT 146.800 305.600 147.600 305.700 ;
        RECT 172.400 305.600 173.200 305.700 ;
        RECT 332.400 306.300 333.200 306.400 ;
        RECT 343.600 306.300 344.400 306.400 ;
        RECT 332.400 305.700 344.400 306.300 ;
        RECT 332.400 305.600 333.200 305.700 ;
        RECT 343.600 305.600 344.400 305.700 ;
        RECT 375.600 306.300 376.400 306.400 ;
        RECT 382.000 306.300 382.800 306.400 ;
        RECT 375.600 305.700 382.800 306.300 ;
        RECT 383.700 306.300 384.300 307.700 ;
        RECT 386.800 307.600 387.600 308.400 ;
        RECT 393.200 308.300 394.000 308.400 ;
        RECT 396.400 308.300 397.200 308.400 ;
        RECT 401.200 308.300 402.000 308.400 ;
        RECT 414.000 308.300 414.800 308.400 ;
        RECT 393.200 307.700 414.800 308.300 ;
        RECT 393.200 307.600 394.000 307.700 ;
        RECT 396.400 307.600 397.200 307.700 ;
        RECT 401.200 307.600 402.000 307.700 ;
        RECT 414.000 307.600 414.800 307.700 ;
        RECT 423.600 308.300 424.400 308.400 ;
        RECT 450.800 308.300 451.600 308.400 ;
        RECT 452.400 308.300 453.200 308.400 ;
        RECT 460.400 308.300 461.200 308.400 ;
        RECT 423.600 307.700 461.200 308.300 ;
        RECT 423.600 307.600 424.400 307.700 ;
        RECT 450.800 307.600 451.600 307.700 ;
        RECT 452.400 307.600 453.200 307.700 ;
        RECT 460.400 307.600 461.200 307.700 ;
        RECT 487.600 308.300 488.400 308.400 ;
        RECT 516.400 308.300 517.200 308.400 ;
        RECT 487.600 307.700 517.200 308.300 ;
        RECT 487.600 307.600 488.400 307.700 ;
        RECT 516.400 307.600 517.200 307.700 ;
        RECT 551.600 308.300 552.400 308.400 ;
        RECT 566.000 308.300 566.800 308.400 ;
        RECT 551.600 307.700 566.800 308.300 ;
        RECT 551.600 307.600 552.400 307.700 ;
        RECT 566.000 307.600 566.800 307.700 ;
        RECT 388.400 306.300 389.200 306.400 ;
        RECT 383.700 305.700 389.200 306.300 ;
        RECT 375.600 305.600 376.400 305.700 ;
        RECT 382.000 305.600 382.800 305.700 ;
        RECT 388.400 305.600 389.200 305.700 ;
        RECT 441.200 306.300 442.000 306.400 ;
        RECT 462.000 306.300 462.800 306.400 ;
        RECT 441.200 305.700 462.800 306.300 ;
        RECT 441.200 305.600 442.000 305.700 ;
        RECT 462.000 305.600 462.800 305.700 ;
        RECT 478.000 306.300 478.800 306.400 ;
        RECT 500.400 306.300 501.200 306.400 ;
        RECT 478.000 305.700 501.200 306.300 ;
        RECT 478.000 305.600 478.800 305.700 ;
        RECT 500.400 305.600 501.200 305.700 ;
        RECT 543.600 306.300 544.400 306.400 ;
        RECT 546.800 306.300 547.600 306.400 ;
        RECT 578.800 306.300 579.600 306.400 ;
        RECT 543.600 305.700 579.600 306.300 ;
        RECT 543.600 305.600 544.400 305.700 ;
        RECT 546.800 305.600 547.600 305.700 ;
        RECT 578.800 305.600 579.600 305.700 ;
        RECT 65.200 304.300 66.000 304.400 ;
        RECT 71.600 304.300 72.400 304.400 ;
        RECT 65.200 303.700 72.400 304.300 ;
        RECT 65.200 303.600 66.000 303.700 ;
        RECT 71.600 303.600 72.400 303.700 ;
        RECT 102.000 304.300 102.800 304.400 ;
        RECT 118.000 304.300 118.800 304.400 ;
        RECT 121.200 304.300 122.000 304.400 ;
        RECT 102.000 303.700 122.000 304.300 ;
        RECT 102.000 303.600 102.800 303.700 ;
        RECT 118.000 303.600 118.800 303.700 ;
        RECT 121.200 303.600 122.000 303.700 ;
        RECT 127.600 304.300 128.400 304.400 ;
        RECT 183.600 304.300 184.400 304.400 ;
        RECT 127.600 303.700 184.400 304.300 ;
        RECT 127.600 303.600 128.400 303.700 ;
        RECT 183.600 303.600 184.400 303.700 ;
        RECT 391.600 304.300 392.400 304.400 ;
        RECT 398.000 304.300 398.800 304.400 ;
        RECT 391.600 303.700 398.800 304.300 ;
        RECT 391.600 303.600 392.400 303.700 ;
        RECT 398.000 303.600 398.800 303.700 ;
        RECT 455.600 304.300 456.400 304.400 ;
        RECT 481.200 304.300 482.000 304.400 ;
        RECT 455.600 303.700 482.000 304.300 ;
        RECT 455.600 303.600 456.400 303.700 ;
        RECT 481.200 303.600 482.000 303.700 ;
        RECT 532.400 304.300 533.200 304.400 ;
        RECT 550.000 304.300 550.800 304.400 ;
        RECT 532.400 303.700 550.800 304.300 ;
        RECT 532.400 303.600 533.200 303.700 ;
        RECT 550.000 303.600 550.800 303.700 ;
        RECT 582.000 303.600 582.800 304.400 ;
        RECT 33.200 302.300 34.000 302.400 ;
        RECT 44.400 302.300 45.200 302.400 ;
        RECT 33.200 301.700 45.200 302.300 ;
        RECT 33.200 301.600 34.000 301.700 ;
        RECT 44.400 301.600 45.200 301.700 ;
        RECT 68.400 302.300 69.200 302.400 ;
        RECT 90.800 302.300 91.600 302.400 ;
        RECT 68.400 301.700 91.600 302.300 ;
        RECT 68.400 301.600 69.200 301.700 ;
        RECT 90.800 301.600 91.600 301.700 ;
        RECT 129.200 302.300 130.000 302.400 ;
        RECT 145.200 302.300 146.000 302.400 ;
        RECT 129.200 301.700 146.000 302.300 ;
        RECT 129.200 301.600 130.000 301.700 ;
        RECT 145.200 301.600 146.000 301.700 ;
        RECT 150.000 302.300 150.800 302.400 ;
        RECT 154.800 302.300 155.600 302.400 ;
        RECT 150.000 301.700 155.600 302.300 ;
        RECT 150.000 301.600 150.800 301.700 ;
        RECT 154.800 301.600 155.600 301.700 ;
        RECT 156.400 302.300 157.200 302.400 ;
        RECT 159.600 302.300 160.400 302.400 ;
        RECT 156.400 301.700 160.400 302.300 ;
        RECT 156.400 301.600 157.200 301.700 ;
        RECT 159.600 301.600 160.400 301.700 ;
        RECT 377.200 302.300 378.000 302.400 ;
        RECT 414.000 302.300 414.800 302.400 ;
        RECT 377.200 301.700 414.800 302.300 ;
        RECT 377.200 301.600 378.000 301.700 ;
        RECT 414.000 301.600 414.800 301.700 ;
        RECT 22.000 300.300 22.800 300.400 ;
        RECT 46.000 300.300 46.800 300.400 ;
        RECT 22.000 299.700 46.800 300.300 ;
        RECT 22.000 299.600 22.800 299.700 ;
        RECT 46.000 299.600 46.800 299.700 ;
        RECT 47.600 300.300 48.400 300.400 ;
        RECT 82.800 300.300 83.600 300.400 ;
        RECT 47.600 299.700 83.600 300.300 ;
        RECT 47.600 299.600 48.400 299.700 ;
        RECT 82.800 299.600 83.600 299.700 ;
        RECT 108.400 300.300 109.200 300.400 ;
        RECT 114.800 300.300 115.600 300.400 ;
        RECT 108.400 299.700 115.600 300.300 ;
        RECT 108.400 299.600 109.200 299.700 ;
        RECT 114.800 299.600 115.600 299.700 ;
        RECT 118.000 300.300 118.800 300.400 ;
        RECT 156.400 300.300 157.200 300.400 ;
        RECT 118.000 299.700 157.200 300.300 ;
        RECT 118.000 299.600 118.800 299.700 ;
        RECT 156.400 299.600 157.200 299.700 ;
        RECT 343.600 300.300 344.400 300.400 ;
        RECT 367.600 300.300 368.400 300.400 ;
        RECT 343.600 299.700 368.400 300.300 ;
        RECT 343.600 299.600 344.400 299.700 ;
        RECT 367.600 299.600 368.400 299.700 ;
        RECT 6.000 297.600 6.800 298.400 ;
        RECT 31.600 298.300 32.400 298.400 ;
        RECT 36.400 298.300 37.200 298.400 ;
        RECT 41.200 298.300 42.000 298.400 ;
        RECT 31.600 297.700 42.000 298.300 ;
        RECT 31.600 297.600 32.400 297.700 ;
        RECT 36.400 297.600 37.200 297.700 ;
        RECT 41.200 297.600 42.000 297.700 ;
        RECT 47.600 298.300 48.400 298.400 ;
        RECT 50.800 298.300 51.600 298.400 ;
        RECT 63.600 298.300 64.400 298.400 ;
        RECT 66.800 298.300 67.600 298.400 ;
        RECT 73.200 298.300 74.000 298.400 ;
        RECT 47.600 297.700 74.000 298.300 ;
        RECT 47.600 297.600 48.400 297.700 ;
        RECT 50.800 297.600 51.600 297.700 ;
        RECT 63.600 297.600 64.400 297.700 ;
        RECT 66.800 297.600 67.600 297.700 ;
        RECT 73.200 297.600 74.000 297.700 ;
        RECT 76.400 298.300 77.200 298.400 ;
        RECT 78.000 298.300 78.800 298.400 ;
        RECT 76.400 297.700 78.800 298.300 ;
        RECT 76.400 297.600 77.200 297.700 ;
        RECT 78.000 297.600 78.800 297.700 ;
        RECT 98.800 298.300 99.600 298.400 ;
        RECT 102.000 298.300 102.800 298.400 ;
        RECT 98.800 297.700 102.800 298.300 ;
        RECT 98.800 297.600 99.600 297.700 ;
        RECT 102.000 297.600 102.800 297.700 ;
        RECT 110.000 298.300 110.800 298.400 ;
        RECT 113.200 298.300 114.000 298.400 ;
        RECT 137.200 298.300 138.000 298.400 ;
        RECT 110.000 297.700 138.000 298.300 ;
        RECT 110.000 297.600 110.800 297.700 ;
        RECT 113.200 297.600 114.000 297.700 ;
        RECT 137.200 297.600 138.000 297.700 ;
        RECT 150.000 298.300 150.800 298.400 ;
        RECT 167.600 298.300 168.400 298.400 ;
        RECT 150.000 297.700 168.400 298.300 ;
        RECT 150.000 297.600 150.800 297.700 ;
        RECT 167.600 297.600 168.400 297.700 ;
        RECT 169.200 298.300 170.000 298.400 ;
        RECT 175.600 298.300 176.400 298.400 ;
        RECT 178.800 298.300 179.600 298.400 ;
        RECT 182.000 298.300 182.800 298.400 ;
        RECT 254.000 298.300 254.800 298.400 ;
        RECT 169.200 297.700 182.800 298.300 ;
        RECT 169.200 297.600 170.000 297.700 ;
        RECT 175.600 297.600 176.400 297.700 ;
        RECT 178.800 297.600 179.600 297.700 ;
        RECT 182.000 297.600 182.800 297.700 ;
        RECT 246.100 297.700 254.800 298.300 ;
        RECT 246.100 296.400 246.700 297.700 ;
        RECT 254.000 297.600 254.800 297.700 ;
        RECT 386.800 298.300 387.600 298.400 ;
        RECT 394.800 298.300 395.600 298.400 ;
        RECT 386.800 297.700 395.600 298.300 ;
        RECT 386.800 297.600 387.600 297.700 ;
        RECT 394.800 297.600 395.600 297.700 ;
        RECT 6.000 296.300 6.800 296.400 ;
        RECT 12.400 296.300 13.200 296.400 ;
        RECT 6.000 295.700 13.200 296.300 ;
        RECT 6.000 295.600 6.800 295.700 ;
        RECT 12.400 295.600 13.200 295.700 ;
        RECT 14.000 296.300 14.800 296.400 ;
        RECT 20.400 296.300 21.200 296.400 ;
        RECT 14.000 295.700 21.200 296.300 ;
        RECT 14.000 295.600 14.800 295.700 ;
        RECT 20.400 295.600 21.200 295.700 ;
        RECT 34.800 296.300 35.600 296.400 ;
        RECT 38.000 296.300 38.800 296.400 ;
        RECT 39.600 296.300 40.400 296.400 ;
        RECT 50.800 296.300 51.600 296.400 ;
        RECT 54.000 296.300 54.800 296.400 ;
        RECT 34.800 295.700 54.800 296.300 ;
        RECT 34.800 295.600 35.600 295.700 ;
        RECT 38.000 295.600 38.800 295.700 ;
        RECT 39.600 295.600 40.400 295.700 ;
        RECT 50.800 295.600 51.600 295.700 ;
        RECT 54.000 295.600 54.800 295.700 ;
        RECT 62.000 296.300 62.800 296.400 ;
        RECT 74.800 296.300 75.600 296.400 ;
        RECT 62.000 295.700 75.600 296.300 ;
        RECT 62.000 295.600 62.800 295.700 ;
        RECT 74.800 295.600 75.600 295.700 ;
        RECT 76.400 296.300 77.200 296.400 ;
        RECT 118.000 296.300 118.800 296.400 ;
        RECT 76.400 295.700 118.800 296.300 ;
        RECT 76.400 295.600 77.200 295.700 ;
        RECT 118.000 295.600 118.800 295.700 ;
        RECT 119.600 296.300 120.400 296.400 ;
        RECT 130.800 296.300 131.600 296.400 ;
        RECT 119.600 295.700 131.600 296.300 ;
        RECT 119.600 295.600 120.400 295.700 ;
        RECT 130.800 295.600 131.600 295.700 ;
        RECT 132.400 296.300 133.200 296.400 ;
        RECT 151.600 296.300 152.400 296.400 ;
        RECT 132.400 295.700 152.400 296.300 ;
        RECT 132.400 295.600 133.200 295.700 ;
        RECT 151.600 295.600 152.400 295.700 ;
        RECT 154.800 296.300 155.600 296.400 ;
        RECT 159.600 296.300 160.400 296.400 ;
        RECT 154.800 295.700 160.400 296.300 ;
        RECT 154.800 295.600 155.600 295.700 ;
        RECT 159.600 295.600 160.400 295.700 ;
        RECT 170.800 296.300 171.600 296.400 ;
        RECT 178.800 296.300 179.600 296.400 ;
        RECT 170.800 295.700 179.600 296.300 ;
        RECT 170.800 295.600 171.600 295.700 ;
        RECT 178.800 295.600 179.600 295.700 ;
        RECT 246.000 295.600 246.800 296.400 ;
        RECT 574.000 296.300 574.800 296.400 ;
        RECT 578.800 296.300 579.600 296.400 ;
        RECT 574.000 295.700 579.600 296.300 ;
        RECT 574.000 295.600 574.800 295.700 ;
        RECT 578.800 295.600 579.600 295.700 ;
        RECT 18.800 294.300 19.600 294.400 ;
        RECT 25.200 294.300 26.000 294.400 ;
        RECT 36.400 294.300 37.200 294.400 ;
        RECT 68.400 294.300 69.200 294.400 ;
        RECT 18.800 293.700 69.200 294.300 ;
        RECT 18.800 293.600 19.600 293.700 ;
        RECT 25.200 293.600 26.000 293.700 ;
        RECT 36.400 293.600 37.200 293.700 ;
        RECT 68.400 293.600 69.200 293.700 ;
        RECT 86.000 294.300 86.800 294.400 ;
        RECT 89.200 294.300 90.000 294.400 ;
        RECT 102.000 294.300 102.800 294.400 ;
        RECT 105.200 294.300 106.000 294.400 ;
        RECT 86.000 293.700 106.000 294.300 ;
        RECT 86.000 293.600 86.800 293.700 ;
        RECT 89.200 293.600 90.000 293.700 ;
        RECT 102.000 293.600 102.800 293.700 ;
        RECT 105.200 293.600 106.000 293.700 ;
        RECT 108.400 293.600 109.200 294.400 ;
        RECT 113.200 294.300 114.000 294.400 ;
        RECT 119.600 294.300 120.400 294.400 ;
        RECT 113.200 293.700 120.400 294.300 ;
        RECT 113.200 293.600 114.000 293.700 ;
        RECT 119.600 293.600 120.400 293.700 ;
        RECT 121.200 294.300 122.000 294.400 ;
        RECT 122.800 294.300 123.600 294.400 ;
        RECT 121.200 293.700 123.600 294.300 ;
        RECT 121.200 293.600 122.000 293.700 ;
        RECT 122.800 293.600 123.600 293.700 ;
        RECT 124.400 294.300 125.200 294.400 ;
        RECT 146.800 294.300 147.600 294.400 ;
        RECT 185.200 294.300 186.000 294.400 ;
        RECT 124.400 293.700 186.000 294.300 ;
        RECT 124.400 293.600 125.200 293.700 ;
        RECT 146.800 293.600 147.600 293.700 ;
        RECT 185.200 293.600 186.000 293.700 ;
        RECT 270.000 294.300 270.800 294.400 ;
        RECT 322.800 294.300 323.600 294.400 ;
        RECT 270.000 293.700 323.600 294.300 ;
        RECT 270.000 293.600 270.800 293.700 ;
        RECT 322.800 293.600 323.600 293.700 ;
        RECT 361.200 294.300 362.000 294.400 ;
        RECT 369.200 294.300 370.000 294.400 ;
        RECT 361.200 293.700 370.000 294.300 ;
        RECT 361.200 293.600 362.000 293.700 ;
        RECT 369.200 293.600 370.000 293.700 ;
        RECT 386.800 294.300 387.600 294.400 ;
        RECT 402.800 294.300 403.600 294.400 ;
        RECT 386.800 293.700 403.600 294.300 ;
        RECT 386.800 293.600 387.600 293.700 ;
        RECT 402.800 293.600 403.600 293.700 ;
        RECT 442.800 294.300 443.600 294.400 ;
        RECT 457.200 294.300 458.000 294.400 ;
        RECT 442.800 293.700 458.000 294.300 ;
        RECT 442.800 293.600 443.600 293.700 ;
        RECT 457.200 293.600 458.000 293.700 ;
        RECT 458.800 294.300 459.600 294.400 ;
        RECT 462.000 294.300 462.800 294.400 ;
        RECT 458.800 293.700 462.800 294.300 ;
        RECT 458.800 293.600 459.600 293.700 ;
        RECT 462.000 293.600 462.800 293.700 ;
        RECT 508.400 294.300 509.200 294.400 ;
        RECT 511.600 294.300 512.400 294.400 ;
        RECT 508.400 293.700 512.400 294.300 ;
        RECT 508.400 293.600 509.200 293.700 ;
        RECT 511.600 293.600 512.400 293.700 ;
        RECT 17.200 292.300 18.000 292.400 ;
        RECT 23.600 292.300 24.400 292.400 ;
        RECT 17.200 291.700 24.400 292.300 ;
        RECT 17.200 291.600 18.000 291.700 ;
        RECT 23.600 291.600 24.400 291.700 ;
        RECT 30.000 292.300 30.800 292.400 ;
        RECT 55.600 292.300 56.400 292.400 ;
        RECT 30.000 291.700 56.400 292.300 ;
        RECT 30.000 291.600 30.800 291.700 ;
        RECT 55.600 291.600 56.400 291.700 ;
        RECT 57.200 292.300 58.000 292.400 ;
        RECT 62.000 292.300 62.800 292.400 ;
        RECT 57.200 291.700 62.800 292.300 ;
        RECT 57.200 291.600 58.000 291.700 ;
        RECT 62.000 291.600 62.800 291.700 ;
        RECT 65.200 292.300 66.000 292.400 ;
        RECT 76.400 292.300 77.200 292.400 ;
        RECT 65.200 291.700 77.200 292.300 ;
        RECT 65.200 291.600 66.000 291.700 ;
        RECT 76.400 291.600 77.200 291.700 ;
        RECT 78.000 292.300 78.800 292.400 ;
        RECT 87.600 292.300 88.400 292.400 ;
        RECT 89.200 292.300 90.000 292.400 ;
        RECT 90.800 292.300 91.600 292.400 ;
        RECT 78.000 291.700 91.600 292.300 ;
        RECT 78.000 291.600 78.800 291.700 ;
        RECT 87.600 291.600 88.400 291.700 ;
        RECT 89.200 291.600 90.000 291.700 ;
        RECT 90.800 291.600 91.600 291.700 ;
        RECT 95.600 292.300 96.400 292.400 ;
        RECT 180.400 292.300 181.200 292.400 ;
        RECT 95.600 291.700 181.200 292.300 ;
        RECT 95.600 291.600 96.400 291.700 ;
        RECT 180.400 291.600 181.200 291.700 ;
        RECT 186.800 292.300 187.600 292.400 ;
        RECT 204.400 292.300 205.200 292.400 ;
        RECT 186.800 291.700 205.200 292.300 ;
        RECT 186.800 291.600 187.600 291.700 ;
        RECT 204.400 291.600 205.200 291.700 ;
        RECT 210.800 292.300 211.600 292.400 ;
        RECT 246.000 292.300 246.800 292.400 ;
        RECT 210.800 291.700 246.800 292.300 ;
        RECT 210.800 291.600 211.600 291.700 ;
        RECT 246.000 291.600 246.800 291.700 ;
        RECT 263.600 292.300 264.400 292.400 ;
        RECT 282.800 292.300 283.600 292.400 ;
        RECT 263.600 291.700 283.600 292.300 ;
        RECT 263.600 291.600 264.400 291.700 ;
        RECT 282.800 291.600 283.600 291.700 ;
        RECT 289.200 292.300 290.000 292.400 ;
        RECT 303.600 292.300 304.400 292.400 ;
        RECT 289.200 291.700 304.400 292.300 ;
        RECT 289.200 291.600 290.000 291.700 ;
        RECT 303.600 291.600 304.400 291.700 ;
        RECT 340.400 292.300 341.200 292.400 ;
        RECT 354.800 292.300 355.600 292.400 ;
        RECT 374.000 292.300 374.800 292.400 ;
        RECT 340.400 291.700 374.800 292.300 ;
        RECT 340.400 291.600 341.200 291.700 ;
        RECT 354.800 291.600 355.600 291.700 ;
        RECT 374.000 291.600 374.800 291.700 ;
        RECT 401.200 292.300 402.000 292.400 ;
        RECT 407.600 292.300 408.400 292.400 ;
        RECT 401.200 291.700 408.400 292.300 ;
        RECT 401.200 291.600 402.000 291.700 ;
        RECT 407.600 291.600 408.400 291.700 ;
        RECT 454.000 292.300 454.800 292.400 ;
        RECT 460.400 292.300 461.200 292.400 ;
        RECT 454.000 291.700 461.200 292.300 ;
        RECT 454.000 291.600 454.800 291.700 ;
        RECT 460.400 291.600 461.200 291.700 ;
        RECT 462.000 292.300 462.800 292.400 ;
        RECT 470.000 292.300 470.800 292.400 ;
        RECT 462.000 291.700 470.800 292.300 ;
        RECT 462.000 291.600 462.800 291.700 ;
        RECT 470.000 291.600 470.800 291.700 ;
        RECT 490.800 292.300 491.600 292.400 ;
        RECT 494.000 292.300 494.800 292.400 ;
        RECT 490.800 291.700 494.800 292.300 ;
        RECT 490.800 291.600 491.600 291.700 ;
        RECT 494.000 291.600 494.800 291.700 ;
        RECT 564.400 292.300 565.200 292.400 ;
        RECT 574.000 292.300 574.800 292.400 ;
        RECT 564.400 291.700 574.800 292.300 ;
        RECT 564.400 291.600 565.200 291.700 ;
        RECT 574.000 291.600 574.800 291.700 ;
        RECT 2.800 290.300 3.600 290.400 ;
        RECT 7.600 290.300 8.400 290.400 ;
        RECT 2.800 289.700 8.400 290.300 ;
        RECT 2.800 289.600 3.600 289.700 ;
        RECT 7.600 289.600 8.400 289.700 ;
        RECT 33.200 290.300 34.000 290.400 ;
        RECT 52.400 290.300 53.200 290.400 ;
        RECT 33.200 289.700 53.200 290.300 ;
        RECT 33.200 289.600 34.000 289.700 ;
        RECT 52.400 289.600 53.200 289.700 ;
        RECT 74.800 290.300 75.600 290.400 ;
        RECT 90.800 290.300 91.600 290.400 ;
        RECT 74.800 289.700 91.600 290.300 ;
        RECT 74.800 289.600 75.600 289.700 ;
        RECT 90.800 289.600 91.600 289.700 ;
        RECT 114.800 290.300 115.600 290.400 ;
        RECT 132.400 290.300 133.200 290.400 ;
        RECT 114.800 289.700 133.200 290.300 ;
        RECT 114.800 289.600 115.600 289.700 ;
        RECT 132.400 289.600 133.200 289.700 ;
        RECT 143.600 290.300 144.400 290.400 ;
        RECT 148.400 290.300 149.200 290.400 ;
        RECT 143.600 289.700 149.200 290.300 ;
        RECT 143.600 289.600 144.400 289.700 ;
        RECT 148.400 289.600 149.200 289.700 ;
        RECT 153.200 290.300 154.000 290.400 ;
        RECT 156.400 290.300 157.200 290.400 ;
        RECT 153.200 289.700 157.200 290.300 ;
        RECT 153.200 289.600 154.000 289.700 ;
        RECT 156.400 289.600 157.200 289.700 ;
        RECT 158.000 290.300 158.800 290.400 ;
        RECT 161.200 290.300 162.000 290.400 ;
        RECT 158.000 289.700 162.000 290.300 ;
        RECT 158.000 289.600 158.800 289.700 ;
        RECT 161.200 289.600 162.000 289.700 ;
        RECT 282.800 290.300 283.600 290.400 ;
        RECT 297.200 290.300 298.000 290.400 ;
        RECT 282.800 289.700 298.000 290.300 ;
        RECT 282.800 289.600 283.600 289.700 ;
        RECT 297.200 289.600 298.000 289.700 ;
        RECT 302.000 290.300 302.800 290.400 ;
        RECT 316.400 290.300 317.200 290.400 ;
        RECT 302.000 289.700 317.200 290.300 ;
        RECT 302.000 289.600 302.800 289.700 ;
        RECT 316.400 289.600 317.200 289.700 ;
        RECT 383.600 290.300 384.400 290.400 ;
        RECT 396.400 290.300 397.200 290.400 ;
        RECT 404.400 290.300 405.200 290.400 ;
        RECT 383.600 289.700 405.200 290.300 ;
        RECT 383.600 289.600 384.400 289.700 ;
        RECT 396.400 289.600 397.200 289.700 ;
        RECT 404.400 289.600 405.200 289.700 ;
        RECT 452.400 290.300 453.200 290.400 ;
        RECT 463.600 290.300 464.400 290.400 ;
        RECT 452.400 289.700 464.400 290.300 ;
        RECT 452.400 289.600 453.200 289.700 ;
        RECT 463.600 289.600 464.400 289.700 ;
        RECT 564.400 290.300 565.200 290.400 ;
        RECT 569.200 290.300 570.000 290.400 ;
        RECT 564.400 289.700 570.000 290.300 ;
        RECT 564.400 289.600 565.200 289.700 ;
        RECT 569.200 289.600 570.000 289.700 ;
        RECT 30.000 288.300 30.800 288.400 ;
        RECT 49.200 288.300 50.000 288.400 ;
        RECT 30.000 287.700 50.000 288.300 ;
        RECT 30.000 287.600 30.800 287.700 ;
        RECT 49.200 287.600 50.000 287.700 ;
        RECT 76.400 288.300 77.200 288.400 ;
        RECT 81.200 288.300 82.000 288.400 ;
        RECT 76.400 287.700 82.000 288.300 ;
        RECT 76.400 287.600 77.200 287.700 ;
        RECT 81.200 287.600 82.000 287.700 ;
        RECT 82.800 288.300 83.600 288.400 ;
        RECT 116.400 288.300 117.200 288.400 ;
        RECT 132.400 288.300 133.200 288.400 ;
        RECT 82.800 287.700 110.700 288.300 ;
        RECT 82.800 287.600 83.600 287.700 ;
        RECT 7.600 286.300 8.400 286.400 ;
        RECT 10.800 286.300 11.600 286.400 ;
        RECT 7.600 285.700 11.600 286.300 ;
        RECT 7.600 285.600 8.400 285.700 ;
        RECT 10.800 285.600 11.600 285.700 ;
        RECT 12.400 286.300 13.200 286.400 ;
        RECT 60.400 286.300 61.200 286.400 ;
        RECT 12.400 285.700 61.200 286.300 ;
        RECT 12.400 285.600 13.200 285.700 ;
        RECT 60.400 285.600 61.200 285.700 ;
        RECT 70.000 286.300 70.800 286.400 ;
        RECT 108.400 286.300 109.200 286.400 ;
        RECT 70.000 285.700 109.200 286.300 ;
        RECT 110.100 286.300 110.700 287.700 ;
        RECT 116.400 287.700 133.200 288.300 ;
        RECT 116.400 287.600 117.200 287.700 ;
        RECT 132.400 287.600 133.200 287.700 ;
        RECT 146.800 288.300 147.600 288.400 ;
        RECT 153.200 288.300 154.000 288.400 ;
        RECT 146.800 287.700 154.000 288.300 ;
        RECT 146.800 287.600 147.600 287.700 ;
        RECT 153.200 287.600 154.000 287.700 ;
        RECT 162.800 288.300 163.600 288.400 ;
        RECT 185.200 288.300 186.000 288.400 ;
        RECT 190.000 288.300 190.800 288.400 ;
        RECT 162.800 287.700 190.800 288.300 ;
        RECT 162.800 287.600 163.600 287.700 ;
        RECT 185.200 287.600 186.000 287.700 ;
        RECT 190.000 287.600 190.800 287.700 ;
        RECT 342.000 288.300 342.800 288.400 ;
        RECT 390.000 288.300 390.800 288.400 ;
        RECT 342.000 287.700 390.800 288.300 ;
        RECT 342.000 287.600 342.800 287.700 ;
        RECT 390.000 287.600 390.800 287.700 ;
        RECT 457.200 288.300 458.000 288.400 ;
        RECT 460.400 288.300 461.200 288.400 ;
        RECT 457.200 287.700 461.200 288.300 ;
        RECT 457.200 287.600 458.000 287.700 ;
        RECT 460.400 287.600 461.200 287.700 ;
        RECT 482.800 288.300 483.600 288.400 ;
        RECT 514.800 288.300 515.600 288.400 ;
        RECT 482.800 287.700 515.600 288.300 ;
        RECT 482.800 287.600 483.600 287.700 ;
        RECT 514.800 287.600 515.600 287.700 ;
        RECT 527.600 288.300 528.400 288.400 ;
        RECT 580.400 288.300 581.200 288.400 ;
        RECT 527.600 287.700 581.200 288.300 ;
        RECT 527.600 287.600 528.400 287.700 ;
        RECT 580.400 287.600 581.200 287.700 ;
        RECT 121.200 286.300 122.000 286.400 ;
        RECT 110.100 285.700 122.000 286.300 ;
        RECT 70.000 285.600 70.800 285.700 ;
        RECT 108.400 285.600 109.200 285.700 ;
        RECT 121.200 285.600 122.000 285.700 ;
        RECT 129.200 286.300 130.000 286.400 ;
        RECT 198.000 286.300 198.800 286.400 ;
        RECT 129.200 285.700 198.800 286.300 ;
        RECT 129.200 285.600 130.000 285.700 ;
        RECT 198.000 285.600 198.800 285.700 ;
        RECT 380.400 286.300 381.200 286.400 ;
        RECT 436.400 286.300 437.200 286.400 ;
        RECT 380.400 285.700 437.200 286.300 ;
        RECT 380.400 285.600 381.200 285.700 ;
        RECT 436.400 285.600 437.200 285.700 ;
        RECT 10.800 284.300 11.600 284.400 ;
        RECT 15.600 284.300 16.400 284.400 ;
        RECT 10.800 283.700 16.400 284.300 ;
        RECT 10.800 283.600 11.600 283.700 ;
        RECT 15.600 283.600 16.400 283.700 ;
        RECT 92.400 284.300 93.200 284.400 ;
        RECT 111.600 284.300 112.400 284.400 ;
        RECT 92.400 283.700 112.400 284.300 ;
        RECT 92.400 283.600 93.200 283.700 ;
        RECT 111.600 283.600 112.400 283.700 ;
        RECT 116.400 284.300 117.200 284.400 ;
        RECT 122.800 284.300 123.600 284.400 ;
        RECT 116.400 283.700 123.600 284.300 ;
        RECT 116.400 283.600 117.200 283.700 ;
        RECT 122.800 283.600 123.600 283.700 ;
        RECT 130.800 284.300 131.600 284.400 ;
        RECT 135.600 284.300 136.400 284.400 ;
        RECT 156.400 284.300 157.200 284.400 ;
        RECT 174.000 284.300 174.800 284.400 ;
        RECT 130.800 283.700 174.800 284.300 ;
        RECT 130.800 283.600 131.600 283.700 ;
        RECT 135.600 283.600 136.400 283.700 ;
        RECT 156.400 283.600 157.200 283.700 ;
        RECT 174.000 283.600 174.800 283.700 ;
        RECT 228.400 284.300 229.200 284.400 ;
        RECT 257.200 284.300 258.000 284.400 ;
        RECT 228.400 283.700 258.000 284.300 ;
        RECT 228.400 283.600 229.200 283.700 ;
        RECT 257.200 283.600 258.000 283.700 ;
        RECT 260.400 284.300 261.200 284.400 ;
        RECT 276.400 284.300 277.200 284.400 ;
        RECT 260.400 283.700 277.200 284.300 ;
        RECT 260.400 283.600 261.200 283.700 ;
        RECT 276.400 283.600 277.200 283.700 ;
        RECT 318.000 284.300 318.800 284.400 ;
        RECT 329.200 284.300 330.000 284.400 ;
        RECT 318.000 283.700 330.000 284.300 ;
        RECT 318.000 283.600 318.800 283.700 ;
        RECT 329.200 283.600 330.000 283.700 ;
        RECT 34.800 280.300 35.600 280.400 ;
        RECT 70.000 280.300 70.800 280.400 ;
        RECT 34.800 279.700 70.800 280.300 ;
        RECT 34.800 279.600 35.600 279.700 ;
        RECT 70.000 279.600 70.800 279.700 ;
        RECT 98.800 280.300 99.600 280.400 ;
        RECT 108.400 280.300 109.200 280.400 ;
        RECT 98.800 279.700 109.200 280.300 ;
        RECT 98.800 279.600 99.600 279.700 ;
        RECT 108.400 279.600 109.200 279.700 ;
        RECT 18.800 278.300 19.600 278.400 ;
        RECT 79.600 278.300 80.400 278.400 ;
        RECT 18.800 277.700 80.400 278.300 ;
        RECT 18.800 277.600 19.600 277.700 ;
        RECT 79.600 277.600 80.400 277.700 ;
        RECT 126.000 278.300 126.800 278.400 ;
        RECT 143.600 278.300 144.400 278.400 ;
        RECT 126.000 277.700 144.400 278.300 ;
        RECT 126.000 277.600 126.800 277.700 ;
        RECT 143.600 277.600 144.400 277.700 ;
        RECT 386.800 278.300 387.600 278.400 ;
        RECT 398.000 278.300 398.800 278.400 ;
        RECT 386.800 277.700 398.800 278.300 ;
        RECT 386.800 277.600 387.600 277.700 ;
        RECT 398.000 277.600 398.800 277.700 ;
        RECT 561.200 278.300 562.000 278.400 ;
        RECT 562.800 278.300 563.600 278.400 ;
        RECT 561.200 277.700 563.600 278.300 ;
        RECT 561.200 277.600 562.000 277.700 ;
        RECT 562.800 277.600 563.600 277.700 ;
        RECT 47.600 276.300 48.400 276.400 ;
        RECT 55.600 276.300 56.400 276.400 ;
        RECT 58.800 276.300 59.600 276.400 ;
        RECT 95.600 276.300 96.400 276.400 ;
        RECT 47.600 275.700 96.400 276.300 ;
        RECT 47.600 275.600 48.400 275.700 ;
        RECT 55.600 275.600 56.400 275.700 ;
        RECT 58.800 275.600 59.600 275.700 ;
        RECT 95.600 275.600 96.400 275.700 ;
        RECT 127.600 276.300 128.400 276.400 ;
        RECT 145.200 276.300 146.000 276.400 ;
        RECT 127.600 275.700 146.000 276.300 ;
        RECT 127.600 275.600 128.400 275.700 ;
        RECT 145.200 275.600 146.000 275.700 ;
        RECT 22.000 274.300 22.800 274.400 ;
        RECT 28.400 274.300 29.200 274.400 ;
        RECT 22.000 273.700 29.200 274.300 ;
        RECT 22.000 273.600 22.800 273.700 ;
        RECT 28.400 273.600 29.200 273.700 ;
        RECT 42.800 274.300 43.600 274.400 ;
        RECT 52.400 274.300 53.200 274.400 ;
        RECT 124.400 274.300 125.200 274.400 ;
        RECT 42.800 273.700 125.200 274.300 ;
        RECT 42.800 273.600 43.600 273.700 ;
        RECT 52.400 273.600 53.200 273.700 ;
        RECT 124.400 273.600 125.200 273.700 ;
        RECT 130.800 274.300 131.600 274.400 ;
        RECT 137.200 274.300 138.000 274.400 ;
        RECT 130.800 273.700 138.000 274.300 ;
        RECT 130.800 273.600 131.600 273.700 ;
        RECT 137.200 273.600 138.000 273.700 ;
        RECT 148.400 274.300 149.200 274.400 ;
        RECT 169.200 274.300 170.000 274.400 ;
        RECT 148.400 273.700 170.000 274.300 ;
        RECT 148.400 273.600 149.200 273.700 ;
        RECT 169.200 273.600 170.000 273.700 ;
        RECT 191.600 274.300 192.400 274.400 ;
        RECT 220.400 274.300 221.200 274.400 ;
        RECT 191.600 273.700 221.200 274.300 ;
        RECT 191.600 273.600 192.400 273.700 ;
        RECT 220.400 273.600 221.200 273.700 ;
        RECT 262.000 274.300 262.800 274.400 ;
        RECT 268.400 274.300 269.200 274.400 ;
        RECT 262.000 273.700 269.200 274.300 ;
        RECT 262.000 273.600 262.800 273.700 ;
        RECT 268.400 273.600 269.200 273.700 ;
        RECT 305.200 274.300 306.000 274.400 ;
        RECT 313.200 274.300 314.000 274.400 ;
        RECT 348.400 274.300 349.200 274.400 ;
        RECT 305.200 273.700 349.200 274.300 ;
        RECT 305.200 273.600 306.000 273.700 ;
        RECT 313.200 273.600 314.000 273.700 ;
        RECT 348.400 273.600 349.200 273.700 ;
        RECT 382.000 274.300 382.800 274.400 ;
        RECT 402.800 274.300 403.600 274.400 ;
        RECT 382.000 273.700 403.600 274.300 ;
        RECT 382.000 273.600 382.800 273.700 ;
        RECT 402.800 273.600 403.600 273.700 ;
        RECT 422.000 274.300 422.800 274.400 ;
        RECT 433.200 274.300 434.000 274.400 ;
        RECT 479.600 274.300 480.400 274.400 ;
        RECT 484.400 274.300 485.200 274.400 ;
        RECT 422.000 273.700 485.200 274.300 ;
        RECT 422.000 273.600 422.800 273.700 ;
        RECT 433.200 273.600 434.000 273.700 ;
        RECT 479.600 273.600 480.400 273.700 ;
        RECT 484.400 273.600 485.200 273.700 ;
        RECT 14.000 272.300 14.800 272.400 ;
        RECT 15.600 272.300 16.400 272.400 ;
        RECT 14.000 271.700 16.400 272.300 ;
        RECT 14.000 271.600 14.800 271.700 ;
        RECT 15.600 271.600 16.400 271.700 ;
        RECT 23.600 272.300 24.400 272.400 ;
        RECT 26.800 272.300 27.600 272.400 ;
        RECT 23.600 271.700 27.600 272.300 ;
        RECT 23.600 271.600 24.400 271.700 ;
        RECT 26.800 271.600 27.600 271.700 ;
        RECT 31.600 272.300 32.400 272.400 ;
        RECT 36.400 272.300 37.200 272.400 ;
        RECT 31.600 271.700 37.200 272.300 ;
        RECT 31.600 271.600 32.400 271.700 ;
        RECT 36.400 271.600 37.200 271.700 ;
        RECT 68.400 272.300 69.200 272.400 ;
        RECT 118.000 272.300 118.800 272.400 ;
        RECT 121.200 272.300 122.000 272.400 ;
        RECT 68.400 271.700 122.000 272.300 ;
        RECT 68.400 271.600 69.200 271.700 ;
        RECT 118.000 271.600 118.800 271.700 ;
        RECT 121.200 271.600 122.000 271.700 ;
        RECT 150.000 272.300 150.800 272.400 ;
        RECT 156.400 272.300 157.200 272.400 ;
        RECT 166.000 272.300 166.800 272.400 ;
        RECT 172.400 272.300 173.200 272.400 ;
        RECT 178.800 272.300 179.600 272.400 ;
        RECT 150.000 271.700 163.500 272.300 ;
        RECT 150.000 271.600 150.800 271.700 ;
        RECT 156.400 271.600 157.200 271.700 ;
        RECT 162.900 270.400 163.500 271.700 ;
        RECT 166.000 271.700 179.600 272.300 ;
        RECT 166.000 271.600 166.800 271.700 ;
        RECT 172.400 271.600 173.200 271.700 ;
        RECT 178.800 271.600 179.600 271.700 ;
        RECT 217.200 272.300 218.000 272.400 ;
        RECT 241.200 272.300 242.000 272.400 ;
        RECT 217.200 271.700 242.000 272.300 ;
        RECT 217.200 271.600 218.000 271.700 ;
        RECT 241.200 271.600 242.000 271.700 ;
        RECT 249.200 272.300 250.000 272.400 ;
        RECT 258.800 272.300 259.600 272.400 ;
        RECT 311.600 272.300 312.400 272.400 ;
        RECT 249.200 271.700 312.400 272.300 ;
        RECT 249.200 271.600 250.000 271.700 ;
        RECT 258.800 271.600 259.600 271.700 ;
        RECT 311.600 271.600 312.400 271.700 ;
        RECT 354.800 272.300 355.600 272.400 ;
        RECT 364.400 272.300 365.200 272.400 ;
        RECT 354.800 271.700 365.200 272.300 ;
        RECT 354.800 271.600 355.600 271.700 ;
        RECT 364.400 271.600 365.200 271.700 ;
        RECT 385.200 272.300 386.000 272.400 ;
        RECT 388.400 272.300 389.200 272.400 ;
        RECT 394.800 272.300 395.600 272.400 ;
        RECT 385.200 271.700 395.600 272.300 ;
        RECT 385.200 271.600 386.000 271.700 ;
        RECT 388.400 271.600 389.200 271.700 ;
        RECT 394.800 271.600 395.600 271.700 ;
        RECT 398.000 272.300 398.800 272.400 ;
        RECT 404.400 272.300 405.200 272.400 ;
        RECT 398.000 271.700 405.200 272.300 ;
        RECT 398.000 271.600 398.800 271.700 ;
        RECT 404.400 271.600 405.200 271.700 ;
        RECT 438.000 271.600 438.800 272.400 ;
        RECT 482.800 272.300 483.600 272.400 ;
        RECT 489.200 272.300 490.000 272.400 ;
        RECT 482.800 271.700 490.000 272.300 ;
        RECT 482.800 271.600 483.600 271.700 ;
        RECT 489.200 271.600 490.000 271.700 ;
        RECT 521.200 272.300 522.000 272.400 ;
        RECT 527.600 272.300 528.400 272.400 ;
        RECT 521.200 271.700 528.400 272.300 ;
        RECT 521.200 271.600 522.000 271.700 ;
        RECT 527.600 271.600 528.400 271.700 ;
        RECT 559.600 272.300 560.400 272.400 ;
        RECT 566.000 272.300 566.800 272.400 ;
        RECT 559.600 271.700 566.800 272.300 ;
        RECT 559.600 271.600 560.400 271.700 ;
        RECT 566.000 271.600 566.800 271.700 ;
        RECT 17.200 270.300 18.000 270.400 ;
        RECT 20.400 270.300 21.200 270.400 ;
        RECT 17.200 269.700 21.200 270.300 ;
        RECT 17.200 269.600 18.000 269.700 ;
        RECT 20.400 269.600 21.200 269.700 ;
        RECT 26.800 270.300 27.600 270.400 ;
        RECT 34.800 270.300 35.600 270.400 ;
        RECT 26.800 269.700 35.600 270.300 ;
        RECT 26.800 269.600 27.600 269.700 ;
        RECT 34.800 269.600 35.600 269.700 ;
        RECT 60.400 270.300 61.200 270.400 ;
        RECT 65.200 270.300 66.000 270.400 ;
        RECT 60.400 269.700 66.000 270.300 ;
        RECT 60.400 269.600 61.200 269.700 ;
        RECT 65.200 269.600 66.000 269.700 ;
        RECT 76.400 270.300 77.200 270.400 ;
        RECT 97.200 270.300 98.000 270.400 ;
        RECT 76.400 269.700 98.000 270.300 ;
        RECT 76.400 269.600 77.200 269.700 ;
        RECT 97.200 269.600 98.000 269.700 ;
        RECT 106.800 270.300 107.600 270.400 ;
        RECT 121.200 270.300 122.000 270.400 ;
        RECT 106.800 269.700 122.000 270.300 ;
        RECT 106.800 269.600 107.600 269.700 ;
        RECT 121.200 269.600 122.000 269.700 ;
        RECT 124.400 270.300 125.200 270.400 ;
        RECT 146.800 270.300 147.600 270.400 ;
        RECT 124.400 269.700 147.600 270.300 ;
        RECT 124.400 269.600 125.200 269.700 ;
        RECT 146.800 269.600 147.600 269.700 ;
        RECT 158.000 270.300 158.800 270.400 ;
        RECT 161.200 270.300 162.000 270.400 ;
        RECT 158.000 269.700 162.000 270.300 ;
        RECT 158.000 269.600 158.800 269.700 ;
        RECT 161.200 269.600 162.000 269.700 ;
        RECT 162.800 270.300 163.600 270.400 ;
        RECT 169.200 270.300 170.000 270.400 ;
        RECT 162.800 269.700 170.000 270.300 ;
        RECT 162.800 269.600 163.600 269.700 ;
        RECT 169.200 269.600 170.000 269.700 ;
        RECT 210.800 270.300 211.600 270.400 ;
        RECT 233.200 270.300 234.000 270.400 ;
        RECT 210.800 269.700 234.000 270.300 ;
        RECT 210.800 269.600 211.600 269.700 ;
        RECT 233.200 269.600 234.000 269.700 ;
        RECT 238.000 270.300 238.800 270.400 ;
        RECT 242.800 270.300 243.600 270.400 ;
        RECT 250.800 270.300 251.600 270.400 ;
        RECT 238.000 269.700 251.600 270.300 ;
        RECT 238.000 269.600 238.800 269.700 ;
        RECT 242.800 269.600 243.600 269.700 ;
        RECT 250.800 269.600 251.600 269.700 ;
        RECT 257.200 270.300 258.000 270.400 ;
        RECT 265.200 270.300 266.000 270.400 ;
        RECT 295.600 270.300 296.400 270.400 ;
        RECT 257.200 269.700 296.400 270.300 ;
        RECT 257.200 269.600 258.000 269.700 ;
        RECT 265.200 269.600 266.000 269.700 ;
        RECT 295.600 269.600 296.400 269.700 ;
        RECT 300.400 270.300 301.200 270.400 ;
        RECT 303.600 270.300 304.400 270.400 ;
        RECT 300.400 269.700 304.400 270.300 ;
        RECT 300.400 269.600 301.200 269.700 ;
        RECT 303.600 269.600 304.400 269.700 ;
        RECT 316.400 270.300 317.200 270.400 ;
        RECT 321.200 270.300 322.000 270.400 ;
        RECT 327.600 270.300 328.400 270.400 ;
        RECT 334.000 270.300 334.800 270.400 ;
        RECT 316.400 269.700 334.800 270.300 ;
        RECT 316.400 269.600 317.200 269.700 ;
        RECT 321.200 269.600 322.000 269.700 ;
        RECT 327.600 269.600 328.400 269.700 ;
        RECT 334.000 269.600 334.800 269.700 ;
        RECT 361.200 270.300 362.000 270.400 ;
        RECT 370.800 270.300 371.600 270.400 ;
        RECT 361.200 269.700 371.600 270.300 ;
        RECT 361.200 269.600 362.000 269.700 ;
        RECT 370.800 269.600 371.600 269.700 ;
        RECT 377.200 270.300 378.000 270.400 ;
        RECT 386.800 270.300 387.600 270.400 ;
        RECT 390.000 270.300 390.800 270.400 ;
        RECT 377.200 269.700 390.800 270.300 ;
        RECT 377.200 269.600 378.000 269.700 ;
        RECT 386.800 269.600 387.600 269.700 ;
        RECT 390.000 269.600 390.800 269.700 ;
        RECT 439.600 270.300 440.400 270.400 ;
        RECT 460.400 270.300 461.200 270.400 ;
        RECT 439.600 269.700 461.200 270.300 ;
        RECT 439.600 269.600 440.400 269.700 ;
        RECT 460.400 269.600 461.200 269.700 ;
        RECT 495.600 270.300 496.400 270.400 ;
        RECT 511.600 270.300 512.400 270.400 ;
        RECT 495.600 269.700 512.400 270.300 ;
        RECT 495.600 269.600 496.400 269.700 ;
        RECT 511.600 269.600 512.400 269.700 ;
        RECT 521.200 270.300 522.000 270.400 ;
        RECT 546.800 270.300 547.600 270.400 ;
        RECT 521.200 269.700 547.600 270.300 ;
        RECT 521.200 269.600 522.000 269.700 ;
        RECT 546.800 269.600 547.600 269.700 ;
        RECT 17.200 268.300 18.000 268.400 ;
        RECT 33.200 268.300 34.000 268.400 ;
        RECT 17.200 267.700 34.000 268.300 ;
        RECT 17.200 267.600 18.000 267.700 ;
        RECT 33.200 267.600 34.000 267.700 ;
        RECT 36.400 268.300 37.200 268.400 ;
        RECT 41.200 268.300 42.000 268.400 ;
        RECT 36.400 267.700 42.000 268.300 ;
        RECT 36.400 267.600 37.200 267.700 ;
        RECT 41.200 267.600 42.000 267.700 ;
        RECT 54.000 268.300 54.800 268.400 ;
        RECT 68.400 268.300 69.200 268.400 ;
        RECT 54.000 267.700 69.200 268.300 ;
        RECT 54.000 267.600 54.800 267.700 ;
        RECT 68.400 267.600 69.200 267.700 ;
        RECT 76.400 268.300 77.200 268.400 ;
        RECT 84.400 268.300 85.200 268.400 ;
        RECT 76.400 267.700 85.200 268.300 ;
        RECT 76.400 267.600 77.200 267.700 ;
        RECT 84.400 267.600 85.200 267.700 ;
        RECT 98.800 268.300 99.600 268.400 ;
        RECT 102.000 268.300 102.800 268.400 ;
        RECT 98.800 267.700 102.800 268.300 ;
        RECT 98.800 267.600 99.600 267.700 ;
        RECT 102.000 267.600 102.800 267.700 ;
        RECT 110.000 268.300 110.800 268.400 ;
        RECT 119.600 268.300 120.400 268.400 ;
        RECT 122.800 268.300 123.600 268.400 ;
        RECT 110.000 267.700 123.600 268.300 ;
        RECT 110.000 267.600 110.800 267.700 ;
        RECT 119.600 267.600 120.400 267.700 ;
        RECT 122.800 267.600 123.600 267.700 ;
        RECT 126.000 268.300 126.800 268.400 ;
        RECT 129.200 268.300 130.000 268.400 ;
        RECT 126.000 267.700 130.000 268.300 ;
        RECT 126.000 267.600 126.800 267.700 ;
        RECT 129.200 267.600 130.000 267.700 ;
        RECT 130.800 268.300 131.600 268.400 ;
        RECT 151.600 268.300 152.400 268.400 ;
        RECT 130.800 267.700 152.400 268.300 ;
        RECT 130.800 267.600 131.600 267.700 ;
        RECT 151.600 267.600 152.400 267.700 ;
        RECT 153.200 268.300 154.000 268.400 ;
        RECT 177.200 268.300 178.000 268.400 ;
        RECT 153.200 267.700 178.000 268.300 ;
        RECT 153.200 267.600 154.000 267.700 ;
        RECT 177.200 267.600 178.000 267.700 ;
        RECT 230.000 268.300 230.800 268.400 ;
        RECT 239.600 268.300 240.400 268.400 ;
        RECT 246.000 268.300 246.800 268.400 ;
        RECT 230.000 267.700 246.800 268.300 ;
        RECT 230.000 267.600 230.800 267.700 ;
        RECT 239.600 267.600 240.400 267.700 ;
        RECT 246.000 267.600 246.800 267.700 ;
        RECT 250.800 268.300 251.600 268.400 ;
        RECT 255.600 268.300 256.400 268.400 ;
        RECT 281.200 268.300 282.000 268.400 ;
        RECT 250.800 267.700 282.000 268.300 ;
        RECT 250.800 267.600 251.600 267.700 ;
        RECT 255.600 267.600 256.400 267.700 ;
        RECT 281.200 267.600 282.000 267.700 ;
        RECT 294.000 268.300 294.800 268.400 ;
        RECT 308.400 268.300 309.200 268.400 ;
        RECT 294.000 267.700 309.200 268.300 ;
        RECT 294.000 267.600 294.800 267.700 ;
        RECT 305.300 266.400 305.900 267.700 ;
        RECT 308.400 267.600 309.200 267.700 ;
        RECT 311.600 268.300 312.400 268.400 ;
        RECT 318.000 268.300 318.800 268.400 ;
        RECT 311.600 267.700 318.800 268.300 ;
        RECT 311.600 267.600 312.400 267.700 ;
        RECT 318.000 267.600 318.800 267.700 ;
        RECT 329.200 268.300 330.000 268.400 ;
        RECT 334.000 268.300 334.800 268.400 ;
        RECT 338.800 268.300 339.600 268.400 ;
        RECT 342.000 268.300 342.800 268.400 ;
        RECT 329.200 267.700 342.800 268.300 ;
        RECT 329.200 267.600 330.000 267.700 ;
        RECT 334.000 267.600 334.800 267.700 ;
        RECT 338.800 267.600 339.600 267.700 ;
        RECT 342.000 267.600 342.800 267.700 ;
        RECT 358.000 268.300 358.800 268.400 ;
        RECT 374.000 268.300 374.800 268.400 ;
        RECT 358.000 267.700 374.800 268.300 ;
        RECT 358.000 267.600 358.800 267.700 ;
        RECT 374.000 267.600 374.800 267.700 ;
        RECT 377.200 268.300 378.000 268.400 ;
        RECT 382.000 268.300 382.800 268.400 ;
        RECT 377.200 267.700 382.800 268.300 ;
        RECT 377.200 267.600 378.000 267.700 ;
        RECT 382.000 267.600 382.800 267.700 ;
        RECT 430.000 268.300 430.800 268.400 ;
        RECT 466.800 268.300 467.600 268.400 ;
        RECT 430.000 267.700 467.600 268.300 ;
        RECT 430.000 267.600 430.800 267.700 ;
        RECT 466.800 267.600 467.600 267.700 ;
        RECT 534.000 268.300 534.800 268.400 ;
        RECT 543.600 268.300 544.400 268.400 ;
        RECT 562.800 268.300 563.600 268.400 ;
        RECT 534.000 267.700 563.600 268.300 ;
        RECT 534.000 267.600 534.800 267.700 ;
        RECT 543.600 267.600 544.400 267.700 ;
        RECT 562.800 267.600 563.600 267.700 ;
        RECT 28.400 266.300 29.200 266.400 ;
        RECT 41.200 266.300 42.000 266.400 ;
        RECT 28.400 265.700 42.000 266.300 ;
        RECT 28.400 265.600 29.200 265.700 ;
        RECT 41.200 265.600 42.000 265.700 ;
        RECT 47.600 266.300 48.400 266.400 ;
        RECT 55.600 266.300 56.400 266.400 ;
        RECT 47.600 265.700 56.400 266.300 ;
        RECT 47.600 265.600 48.400 265.700 ;
        RECT 55.600 265.600 56.400 265.700 ;
        RECT 82.800 266.300 83.600 266.400 ;
        RECT 100.400 266.300 101.200 266.400 ;
        RECT 82.800 265.700 101.200 266.300 ;
        RECT 82.800 265.600 83.600 265.700 ;
        RECT 100.400 265.600 101.200 265.700 ;
        RECT 116.400 266.300 117.200 266.400 ;
        RECT 132.400 266.300 133.200 266.400 ;
        RECT 154.800 266.300 155.600 266.400 ;
        RECT 159.600 266.300 160.400 266.400 ;
        RECT 164.400 266.300 165.200 266.400 ;
        RECT 116.400 265.700 165.200 266.300 ;
        RECT 116.400 265.600 117.200 265.700 ;
        RECT 132.400 265.600 133.200 265.700 ;
        RECT 154.800 265.600 155.600 265.700 ;
        RECT 159.600 265.600 160.400 265.700 ;
        RECT 164.400 265.600 165.200 265.700 ;
        RECT 234.800 266.300 235.600 266.400 ;
        RECT 244.400 266.300 245.200 266.400 ;
        RECT 262.000 266.300 262.800 266.400 ;
        RECT 234.800 265.700 262.800 266.300 ;
        RECT 234.800 265.600 235.600 265.700 ;
        RECT 244.400 265.600 245.200 265.700 ;
        RECT 262.000 265.600 262.800 265.700 ;
        RECT 279.600 266.300 280.400 266.400 ;
        RECT 282.800 266.300 283.600 266.400 ;
        RECT 279.600 265.700 283.600 266.300 ;
        RECT 279.600 265.600 280.400 265.700 ;
        RECT 282.800 265.600 283.600 265.700 ;
        RECT 284.400 266.300 285.200 266.400 ;
        RECT 303.600 266.300 304.400 266.400 ;
        RECT 284.400 265.700 304.400 266.300 ;
        RECT 284.400 265.600 285.200 265.700 ;
        RECT 303.600 265.600 304.400 265.700 ;
        RECT 305.200 265.600 306.000 266.400 ;
        RECT 306.800 266.300 307.600 266.400 ;
        RECT 321.200 266.300 322.000 266.400 ;
        RECT 306.800 265.700 322.000 266.300 ;
        RECT 306.800 265.600 307.600 265.700 ;
        RECT 321.200 265.600 322.000 265.700 ;
        RECT 334.000 266.300 334.800 266.400 ;
        RECT 340.400 266.300 341.200 266.400 ;
        RECT 345.200 266.300 346.000 266.400 ;
        RECT 334.000 265.700 346.000 266.300 ;
        RECT 334.000 265.600 334.800 265.700 ;
        RECT 340.400 265.600 341.200 265.700 ;
        RECT 345.200 265.600 346.000 265.700 ;
        RECT 380.400 266.300 381.200 266.400 ;
        RECT 402.800 266.300 403.600 266.400 ;
        RECT 412.400 266.300 413.200 266.400 ;
        RECT 380.400 265.700 389.100 266.300 ;
        RECT 380.400 265.600 381.200 265.700 ;
        RECT 388.500 264.400 389.100 265.700 ;
        RECT 402.800 265.700 413.200 266.300 ;
        RECT 402.800 265.600 403.600 265.700 ;
        RECT 412.400 265.600 413.200 265.700 ;
        RECT 6.000 264.300 6.800 264.400 ;
        RECT 33.200 264.300 34.000 264.400 ;
        RECT 6.000 263.700 34.000 264.300 ;
        RECT 6.000 263.600 6.800 263.700 ;
        RECT 33.200 263.600 34.000 263.700 ;
        RECT 46.000 264.300 46.800 264.400 ;
        RECT 49.200 264.300 50.000 264.400 ;
        RECT 62.000 264.300 62.800 264.400 ;
        RECT 46.000 263.700 62.800 264.300 ;
        RECT 46.000 263.600 46.800 263.700 ;
        RECT 49.200 263.600 50.000 263.700 ;
        RECT 62.000 263.600 62.800 263.700 ;
        RECT 134.000 264.300 134.800 264.400 ;
        RECT 137.200 264.300 138.000 264.400 ;
        RECT 175.600 264.300 176.400 264.400 ;
        RECT 134.000 263.700 176.400 264.300 ;
        RECT 134.000 263.600 134.800 263.700 ;
        RECT 137.200 263.600 138.000 263.700 ;
        RECT 175.600 263.600 176.400 263.700 ;
        RECT 182.000 264.300 182.800 264.400 ;
        RECT 198.000 264.300 198.800 264.400 ;
        RECT 182.000 263.700 198.800 264.300 ;
        RECT 182.000 263.600 182.800 263.700 ;
        RECT 198.000 263.600 198.800 263.700 ;
        RECT 215.600 264.300 216.400 264.400 ;
        RECT 287.600 264.300 288.400 264.400 ;
        RECT 215.600 263.700 288.400 264.300 ;
        RECT 215.600 263.600 216.400 263.700 ;
        RECT 287.600 263.600 288.400 263.700 ;
        RECT 310.000 264.300 310.800 264.400 ;
        RECT 332.400 264.300 333.200 264.400 ;
        RECT 310.000 263.700 333.200 264.300 ;
        RECT 310.000 263.600 310.800 263.700 ;
        RECT 332.400 263.600 333.200 263.700 ;
        RECT 370.800 264.300 371.600 264.400 ;
        RECT 383.600 264.300 384.400 264.400 ;
        RECT 370.800 263.700 384.400 264.300 ;
        RECT 370.800 263.600 371.600 263.700 ;
        RECT 383.600 263.600 384.400 263.700 ;
        RECT 388.400 264.300 389.200 264.400 ;
        RECT 393.200 264.300 394.000 264.400 ;
        RECT 396.400 264.300 397.200 264.400 ;
        RECT 388.400 263.700 397.200 264.300 ;
        RECT 388.400 263.600 389.200 263.700 ;
        RECT 393.200 263.600 394.000 263.700 ;
        RECT 396.400 263.600 397.200 263.700 ;
        RECT 444.400 264.300 445.200 264.400 ;
        RECT 457.200 264.300 458.000 264.400 ;
        RECT 444.400 263.700 458.000 264.300 ;
        RECT 444.400 263.600 445.200 263.700 ;
        RECT 457.200 263.600 458.000 263.700 ;
        RECT 540.400 264.300 541.200 264.400 ;
        RECT 577.200 264.300 578.000 264.400 ;
        RECT 540.400 263.700 578.000 264.300 ;
        RECT 540.400 263.600 541.200 263.700 ;
        RECT 577.200 263.600 578.000 263.700 ;
        RECT 6.000 262.300 6.800 262.400 ;
        RECT 18.800 262.300 19.600 262.400 ;
        RECT 92.400 262.300 93.200 262.400 ;
        RECT 6.000 261.700 93.200 262.300 ;
        RECT 6.000 261.600 6.800 261.700 ;
        RECT 18.800 261.600 19.600 261.700 ;
        RECT 92.400 261.600 93.200 261.700 ;
        RECT 324.400 262.300 325.200 262.400 ;
        RECT 329.200 262.300 330.000 262.400 ;
        RECT 358.000 262.300 358.800 262.400 ;
        RECT 324.400 261.700 358.800 262.300 ;
        RECT 324.400 261.600 325.200 261.700 ;
        RECT 329.200 261.600 330.000 261.700 ;
        RECT 358.000 261.600 358.800 261.700 ;
        RECT 438.000 262.300 438.800 262.400 ;
        RECT 487.600 262.300 488.400 262.400 ;
        RECT 438.000 261.700 488.400 262.300 ;
        RECT 438.000 261.600 438.800 261.700 ;
        RECT 487.600 261.600 488.400 261.700 ;
        RECT 502.000 262.300 502.800 262.400 ;
        RECT 556.400 262.300 557.200 262.400 ;
        RECT 502.000 261.700 557.200 262.300 ;
        RECT 502.000 261.600 502.800 261.700 ;
        RECT 556.400 261.600 557.200 261.700 ;
        RECT 14.000 260.300 14.800 260.400 ;
        RECT 54.000 260.300 54.800 260.400 ;
        RECT 14.000 259.700 54.800 260.300 ;
        RECT 14.000 259.600 14.800 259.700 ;
        RECT 54.000 259.600 54.800 259.700 ;
        RECT 102.000 260.300 102.800 260.400 ;
        RECT 110.000 260.300 110.800 260.400 ;
        RECT 118.000 260.300 118.800 260.400 ;
        RECT 102.000 259.700 118.800 260.300 ;
        RECT 102.000 259.600 102.800 259.700 ;
        RECT 110.000 259.600 110.800 259.700 ;
        RECT 118.000 259.600 118.800 259.700 ;
        RECT 167.600 260.300 168.400 260.400 ;
        RECT 170.800 260.300 171.600 260.400 ;
        RECT 167.600 259.700 171.600 260.300 ;
        RECT 167.600 259.600 168.400 259.700 ;
        RECT 170.800 259.600 171.600 259.700 ;
        RECT 190.000 260.300 190.800 260.400 ;
        RECT 198.000 260.300 198.800 260.400 ;
        RECT 260.400 260.300 261.200 260.400 ;
        RECT 190.000 259.700 261.200 260.300 ;
        RECT 190.000 259.600 190.800 259.700 ;
        RECT 198.000 259.600 198.800 259.700 ;
        RECT 260.400 259.600 261.200 259.700 ;
        RECT 372.400 260.300 373.200 260.400 ;
        RECT 393.200 260.300 394.000 260.400 ;
        RECT 398.000 260.300 398.800 260.400 ;
        RECT 372.400 259.700 398.800 260.300 ;
        RECT 372.400 259.600 373.200 259.700 ;
        RECT 393.200 259.600 394.000 259.700 ;
        RECT 398.000 259.600 398.800 259.700 ;
        RECT 434.800 260.300 435.600 260.400 ;
        RECT 439.600 260.300 440.400 260.400 ;
        RECT 452.400 260.300 453.200 260.400 ;
        RECT 434.800 259.700 453.200 260.300 ;
        RECT 434.800 259.600 435.600 259.700 ;
        RECT 439.600 259.600 440.400 259.700 ;
        RECT 452.400 259.600 453.200 259.700 ;
        RECT 458.800 260.300 459.600 260.400 ;
        RECT 463.600 260.300 464.400 260.400 ;
        RECT 481.200 260.300 482.000 260.400 ;
        RECT 494.000 260.300 494.800 260.400 ;
        RECT 458.800 259.700 494.800 260.300 ;
        RECT 458.800 259.600 459.600 259.700 ;
        RECT 463.600 259.600 464.400 259.700 ;
        RECT 481.200 259.600 482.000 259.700 ;
        RECT 494.000 259.600 494.800 259.700 ;
        RECT 10.800 258.300 11.600 258.400 ;
        RECT 20.400 258.300 21.200 258.400 ;
        RECT 10.800 257.700 21.200 258.300 ;
        RECT 10.800 257.600 11.600 257.700 ;
        RECT 20.400 257.600 21.200 257.700 ;
        RECT 78.000 258.300 78.800 258.400 ;
        RECT 90.800 258.300 91.600 258.400 ;
        RECT 118.000 258.300 118.800 258.400 ;
        RECT 78.000 257.700 118.800 258.300 ;
        RECT 78.000 257.600 78.800 257.700 ;
        RECT 90.800 257.600 91.600 257.700 ;
        RECT 118.000 257.600 118.800 257.700 ;
        RECT 169.200 258.300 170.000 258.400 ;
        RECT 218.800 258.300 219.600 258.400 ;
        RECT 169.200 257.700 219.600 258.300 ;
        RECT 169.200 257.600 170.000 257.700 ;
        RECT 218.800 257.600 219.600 257.700 ;
        RECT 241.200 258.300 242.000 258.400 ;
        RECT 262.000 258.300 262.800 258.400 ;
        RECT 241.200 257.700 262.800 258.300 ;
        RECT 241.200 257.600 242.000 257.700 ;
        RECT 262.000 257.600 262.800 257.700 ;
        RECT 319.600 258.300 320.400 258.400 ;
        RECT 327.600 258.300 328.400 258.400 ;
        RECT 330.800 258.300 331.600 258.400 ;
        RECT 340.400 258.300 341.200 258.400 ;
        RECT 319.600 257.700 341.200 258.300 ;
        RECT 319.600 257.600 320.400 257.700 ;
        RECT 327.600 257.600 328.400 257.700 ;
        RECT 330.800 257.600 331.600 257.700 ;
        RECT 340.400 257.600 341.200 257.700 ;
        RECT 366.000 258.300 366.800 258.400 ;
        RECT 399.600 258.300 400.400 258.400 ;
        RECT 366.000 257.700 400.400 258.300 ;
        RECT 366.000 257.600 366.800 257.700 ;
        RECT 399.600 257.600 400.400 257.700 ;
        RECT 406.000 258.300 406.800 258.400 ;
        RECT 418.800 258.300 419.600 258.400 ;
        RECT 406.000 257.700 419.600 258.300 ;
        RECT 406.000 257.600 406.800 257.700 ;
        RECT 418.800 257.600 419.600 257.700 ;
        RECT 431.600 258.300 432.400 258.400 ;
        RECT 529.200 258.300 530.000 258.400 ;
        RECT 431.600 257.700 530.000 258.300 ;
        RECT 431.600 257.600 432.400 257.700 ;
        RECT 529.200 257.600 530.000 257.700 ;
        RECT 15.600 255.600 16.400 256.400 ;
        RECT 18.800 256.300 19.600 256.400 ;
        RECT 22.000 256.300 22.800 256.400 ;
        RECT 26.800 256.300 27.600 256.400 ;
        RECT 18.800 255.700 27.600 256.300 ;
        RECT 18.800 255.600 19.600 255.700 ;
        RECT 22.000 255.600 22.800 255.700 ;
        RECT 26.800 255.600 27.600 255.700 ;
        RECT 33.200 256.300 34.000 256.400 ;
        RECT 50.800 256.300 51.600 256.400 ;
        RECT 33.200 255.700 51.600 256.300 ;
        RECT 33.200 255.600 34.000 255.700 ;
        RECT 50.800 255.600 51.600 255.700 ;
        RECT 89.200 256.300 90.000 256.400 ;
        RECT 94.000 256.300 94.800 256.400 ;
        RECT 89.200 255.700 94.800 256.300 ;
        RECT 89.200 255.600 90.000 255.700 ;
        RECT 94.000 255.600 94.800 255.700 ;
        RECT 114.800 256.300 115.600 256.400 ;
        RECT 122.800 256.300 123.600 256.400 ;
        RECT 114.800 255.700 123.600 256.300 ;
        RECT 114.800 255.600 115.600 255.700 ;
        RECT 122.800 255.600 123.600 255.700 ;
        RECT 180.400 256.300 181.200 256.400 ;
        RECT 186.800 256.300 187.600 256.400 ;
        RECT 180.400 255.700 187.600 256.300 ;
        RECT 180.400 255.600 181.200 255.700 ;
        RECT 186.800 255.600 187.600 255.700 ;
        RECT 193.200 256.300 194.000 256.400 ;
        RECT 199.600 256.300 200.400 256.400 ;
        RECT 193.200 255.700 200.400 256.300 ;
        RECT 193.200 255.600 194.000 255.700 ;
        RECT 199.600 255.600 200.400 255.700 ;
        RECT 230.000 256.300 230.800 256.400 ;
        RECT 273.200 256.300 274.000 256.400 ;
        RECT 230.000 255.700 274.000 256.300 ;
        RECT 230.000 255.600 230.800 255.700 ;
        RECT 273.200 255.600 274.000 255.700 ;
        RECT 319.600 256.300 320.400 256.400 ;
        RECT 326.000 256.300 326.800 256.400 ;
        RECT 319.600 255.700 326.800 256.300 ;
        RECT 319.600 255.600 320.400 255.700 ;
        RECT 326.000 255.600 326.800 255.700 ;
        RECT 350.000 256.300 350.800 256.400 ;
        RECT 353.200 256.300 354.000 256.400 ;
        RECT 350.000 255.700 354.000 256.300 ;
        RECT 350.000 255.600 350.800 255.700 ;
        RECT 353.200 255.600 354.000 255.700 ;
        RECT 394.800 256.300 395.600 256.400 ;
        RECT 410.800 256.300 411.600 256.400 ;
        RECT 394.800 255.700 411.600 256.300 ;
        RECT 394.800 255.600 395.600 255.700 ;
        RECT 410.800 255.600 411.600 255.700 ;
        RECT 498.800 256.300 499.600 256.400 ;
        RECT 502.000 256.300 502.800 256.400 ;
        RECT 498.800 255.700 502.800 256.300 ;
        RECT 498.800 255.600 499.600 255.700 ;
        RECT 502.000 255.600 502.800 255.700 ;
        RECT 1.200 254.300 2.000 254.400 ;
        RECT 22.000 254.300 22.800 254.400 ;
        RECT 1.200 253.700 22.800 254.300 ;
        RECT 1.200 253.600 2.000 253.700 ;
        RECT 22.000 253.600 22.800 253.700 ;
        RECT 39.600 254.300 40.400 254.400 ;
        RECT 47.600 254.300 48.400 254.400 ;
        RECT 39.600 253.700 48.400 254.300 ;
        RECT 39.600 253.600 40.400 253.700 ;
        RECT 47.600 253.600 48.400 253.700 ;
        RECT 60.400 253.600 61.200 254.400 ;
        RECT 62.000 254.300 62.800 254.400 ;
        RECT 73.200 254.300 74.000 254.400 ;
        RECT 62.000 253.700 74.000 254.300 ;
        RECT 62.000 253.600 62.800 253.700 ;
        RECT 73.200 253.600 74.000 253.700 ;
        RECT 74.800 254.300 75.600 254.400 ;
        RECT 78.000 254.300 78.800 254.400 ;
        RECT 74.800 253.700 78.800 254.300 ;
        RECT 74.800 253.600 75.600 253.700 ;
        RECT 78.000 253.600 78.800 253.700 ;
        RECT 87.600 254.300 88.400 254.400 ;
        RECT 97.200 254.300 98.000 254.400 ;
        RECT 87.600 253.700 98.000 254.300 ;
        RECT 87.600 253.600 88.400 253.700 ;
        RECT 97.200 253.600 98.000 253.700 ;
        RECT 102.000 254.300 102.800 254.400 ;
        RECT 105.200 254.300 106.000 254.400 ;
        RECT 111.600 254.300 112.400 254.400 ;
        RECT 102.000 253.700 112.400 254.300 ;
        RECT 102.000 253.600 102.800 253.700 ;
        RECT 105.200 253.600 106.000 253.700 ;
        RECT 111.600 253.600 112.400 253.700 ;
        RECT 153.200 254.300 154.000 254.400 ;
        RECT 156.400 254.300 157.200 254.400 ;
        RECT 153.200 253.700 157.200 254.300 ;
        RECT 153.200 253.600 154.000 253.700 ;
        RECT 156.400 253.600 157.200 253.700 ;
        RECT 175.600 254.300 176.400 254.400 ;
        RECT 182.000 254.300 182.800 254.400 ;
        RECT 175.600 253.700 182.800 254.300 ;
        RECT 175.600 253.600 176.400 253.700 ;
        RECT 182.000 253.600 182.800 253.700 ;
        RECT 255.600 254.300 256.400 254.400 ;
        RECT 281.200 254.300 282.000 254.400 ;
        RECT 255.600 253.700 282.000 254.300 ;
        RECT 255.600 253.600 256.400 253.700 ;
        RECT 281.200 253.600 282.000 253.700 ;
        RECT 310.000 254.300 310.800 254.400 ;
        RECT 321.200 254.300 322.000 254.400 ;
        RECT 310.000 253.700 322.000 254.300 ;
        RECT 310.000 253.600 310.800 253.700 ;
        RECT 321.200 253.600 322.000 253.700 ;
        RECT 322.800 254.300 323.600 254.400 ;
        RECT 324.400 254.300 325.200 254.400 ;
        RECT 322.800 253.700 325.200 254.300 ;
        RECT 322.800 253.600 323.600 253.700 ;
        RECT 324.400 253.600 325.200 253.700 ;
        RECT 332.400 254.300 333.200 254.400 ;
        RECT 343.600 254.300 344.400 254.400 ;
        RECT 350.000 254.300 350.800 254.400 ;
        RECT 332.400 253.700 350.800 254.300 ;
        RECT 332.400 253.600 333.200 253.700 ;
        RECT 343.600 253.600 344.400 253.700 ;
        RECT 350.000 253.600 350.800 253.700 ;
        RECT 356.400 254.300 357.200 254.400 ;
        RECT 362.800 254.300 363.600 254.400 ;
        RECT 367.600 254.300 368.400 254.400 ;
        RECT 356.400 253.700 368.400 254.300 ;
        RECT 356.400 253.600 357.200 253.700 ;
        RECT 362.800 253.600 363.600 253.700 ;
        RECT 367.600 253.600 368.400 253.700 ;
        RECT 383.600 254.300 384.400 254.400 ;
        RECT 415.600 254.300 416.400 254.400 ;
        RECT 430.000 254.300 430.800 254.400 ;
        RECT 383.600 253.700 430.800 254.300 ;
        RECT 383.600 253.600 384.400 253.700 ;
        RECT 415.600 253.600 416.400 253.700 ;
        RECT 430.000 253.600 430.800 253.700 ;
        RECT 462.000 254.300 462.800 254.400 ;
        RECT 468.400 254.300 469.200 254.400 ;
        RECT 462.000 253.700 469.200 254.300 ;
        RECT 462.000 253.600 462.800 253.700 ;
        RECT 468.400 253.600 469.200 253.700 ;
        RECT 502.000 254.300 502.800 254.400 ;
        RECT 513.200 254.300 514.000 254.400 ;
        RECT 502.000 253.700 514.000 254.300 ;
        RECT 502.000 253.600 502.800 253.700 ;
        RECT 513.200 253.600 514.000 253.700 ;
        RECT 31.600 252.300 32.400 252.400 ;
        RECT 34.800 252.300 35.600 252.400 ;
        RECT 31.600 251.700 35.600 252.300 ;
        RECT 31.600 251.600 32.400 251.700 ;
        RECT 34.800 251.600 35.600 251.700 ;
        RECT 82.800 252.300 83.600 252.400 ;
        RECT 113.200 252.300 114.000 252.400 ;
        RECT 82.800 251.700 114.000 252.300 ;
        RECT 82.800 251.600 83.600 251.700 ;
        RECT 113.200 251.600 114.000 251.700 ;
        RECT 150.000 252.300 150.800 252.400 ;
        RECT 154.800 252.300 155.600 252.400 ;
        RECT 169.200 252.300 170.000 252.400 ;
        RECT 150.000 251.700 170.000 252.300 ;
        RECT 150.000 251.600 150.800 251.700 ;
        RECT 154.800 251.600 155.600 251.700 ;
        RECT 169.200 251.600 170.000 251.700 ;
        RECT 177.200 252.300 178.000 252.400 ;
        RECT 178.800 252.300 179.600 252.400 ;
        RECT 186.800 252.300 187.600 252.400 ;
        RECT 190.000 252.300 190.800 252.400 ;
        RECT 177.200 251.700 190.800 252.300 ;
        RECT 177.200 251.600 178.000 251.700 ;
        RECT 178.800 251.600 179.600 251.700 ;
        RECT 186.800 251.600 187.600 251.700 ;
        RECT 190.000 251.600 190.800 251.700 ;
        RECT 212.400 252.300 213.200 252.400 ;
        RECT 215.600 252.300 216.400 252.400 ;
        RECT 212.400 251.700 216.400 252.300 ;
        RECT 212.400 251.600 213.200 251.700 ;
        RECT 215.600 251.600 216.400 251.700 ;
        RECT 258.800 252.300 259.600 252.400 ;
        RECT 263.600 252.300 264.400 252.400 ;
        RECT 268.400 252.300 269.200 252.400 ;
        RECT 297.200 252.300 298.000 252.400 ;
        RECT 258.800 251.700 298.000 252.300 ;
        RECT 258.800 251.600 259.600 251.700 ;
        RECT 263.600 251.600 264.400 251.700 ;
        RECT 268.400 251.600 269.200 251.700 ;
        RECT 297.200 251.600 298.000 251.700 ;
        RECT 303.600 252.300 304.400 252.400 ;
        RECT 322.800 252.300 323.600 252.400 ;
        RECT 303.600 251.700 323.600 252.300 ;
        RECT 303.600 251.600 304.400 251.700 ;
        RECT 322.800 251.600 323.600 251.700 ;
        RECT 324.400 252.300 325.200 252.400 ;
        RECT 334.000 252.300 334.800 252.400 ;
        RECT 324.400 251.700 334.800 252.300 ;
        RECT 324.400 251.600 325.200 251.700 ;
        RECT 334.000 251.600 334.800 251.700 ;
        RECT 337.200 252.300 338.000 252.400 ;
        RECT 356.400 252.300 357.200 252.400 ;
        RECT 337.200 251.700 357.200 252.300 ;
        RECT 337.200 251.600 338.000 251.700 ;
        RECT 356.400 251.600 357.200 251.700 ;
        RECT 361.200 252.300 362.000 252.400 ;
        RECT 366.000 252.300 366.800 252.400 ;
        RECT 361.200 251.700 366.800 252.300 ;
        RECT 361.200 251.600 362.000 251.700 ;
        RECT 366.000 251.600 366.800 251.700 ;
        RECT 380.400 252.300 381.200 252.400 ;
        RECT 390.000 252.300 390.800 252.400 ;
        RECT 380.400 251.700 390.800 252.300 ;
        RECT 380.400 251.600 381.200 251.700 ;
        RECT 390.000 251.600 390.800 251.700 ;
        RECT 398.000 252.300 398.800 252.400 ;
        RECT 409.200 252.300 410.000 252.400 ;
        RECT 398.000 251.700 410.000 252.300 ;
        RECT 398.000 251.600 398.800 251.700 ;
        RECT 409.200 251.600 410.000 251.700 ;
        RECT 438.000 252.300 438.800 252.400 ;
        RECT 441.200 252.300 442.000 252.400 ;
        RECT 450.800 252.300 451.600 252.400 ;
        RECT 438.000 251.700 451.600 252.300 ;
        RECT 438.000 251.600 438.800 251.700 ;
        RECT 441.200 251.600 442.000 251.700 ;
        RECT 450.800 251.600 451.600 251.700 ;
        RECT 466.800 252.300 467.600 252.400 ;
        RECT 471.600 252.300 472.400 252.400 ;
        RECT 466.800 251.700 472.400 252.300 ;
        RECT 466.800 251.600 467.600 251.700 ;
        RECT 471.600 251.600 472.400 251.700 ;
        RECT 474.800 252.300 475.600 252.400 ;
        RECT 486.000 252.300 486.800 252.400 ;
        RECT 474.800 251.700 486.800 252.300 ;
        RECT 474.800 251.600 475.600 251.700 ;
        RECT 486.000 251.600 486.800 251.700 ;
        RECT 508.400 252.300 509.200 252.400 ;
        RECT 514.800 252.300 515.600 252.400 ;
        RECT 508.400 251.700 515.600 252.300 ;
        RECT 508.400 251.600 509.200 251.700 ;
        RECT 514.800 251.600 515.600 251.700 ;
        RECT 15.600 250.300 16.400 250.400 ;
        RECT 31.600 250.300 32.400 250.400 ;
        RECT 41.200 250.300 42.000 250.400 ;
        RECT 46.000 250.300 46.800 250.400 ;
        RECT 15.600 249.700 46.800 250.300 ;
        RECT 15.600 249.600 16.400 249.700 ;
        RECT 31.600 249.600 32.400 249.700 ;
        RECT 41.200 249.600 42.000 249.700 ;
        RECT 46.000 249.600 46.800 249.700 ;
        RECT 161.200 250.300 162.000 250.400 ;
        RECT 177.200 250.300 178.000 250.400 ;
        RECT 161.200 249.700 178.000 250.300 ;
        RECT 161.200 249.600 162.000 249.700 ;
        RECT 177.200 249.600 178.000 249.700 ;
        RECT 274.800 250.300 275.600 250.400 ;
        RECT 313.200 250.300 314.000 250.400 ;
        RECT 274.800 249.700 314.000 250.300 ;
        RECT 274.800 249.600 275.600 249.700 ;
        RECT 313.200 249.600 314.000 249.700 ;
        RECT 321.200 250.300 322.000 250.400 ;
        RECT 322.800 250.300 323.600 250.400 ;
        RECT 321.200 249.700 323.600 250.300 ;
        RECT 321.200 249.600 322.000 249.700 ;
        RECT 322.800 249.600 323.600 249.700 ;
        RECT 324.400 250.300 325.200 250.400 ;
        RECT 334.000 250.300 334.800 250.400 ;
        RECT 324.400 249.700 334.800 250.300 ;
        RECT 324.400 249.600 325.200 249.700 ;
        RECT 334.000 249.600 334.800 249.700 ;
        RECT 345.200 250.300 346.000 250.400 ;
        RECT 353.200 250.300 354.000 250.400 ;
        RECT 364.400 250.300 365.200 250.400 ;
        RECT 345.200 249.700 365.200 250.300 ;
        RECT 345.200 249.600 346.000 249.700 ;
        RECT 353.200 249.600 354.000 249.700 ;
        RECT 364.400 249.600 365.200 249.700 ;
        RECT 442.800 250.300 443.600 250.400 ;
        RECT 454.000 250.300 454.800 250.400 ;
        RECT 468.400 250.300 469.200 250.400 ;
        RECT 442.800 249.700 469.200 250.300 ;
        RECT 442.800 249.600 443.600 249.700 ;
        RECT 454.000 249.600 454.800 249.700 ;
        RECT 468.400 249.600 469.200 249.700 ;
        RECT 486.000 250.300 486.800 250.400 ;
        RECT 489.200 250.300 490.000 250.400 ;
        RECT 486.000 249.700 490.000 250.300 ;
        RECT 486.000 249.600 486.800 249.700 ;
        RECT 489.200 249.600 490.000 249.700 ;
        RECT 98.800 248.300 99.600 248.400 ;
        RECT 103.600 248.300 104.400 248.400 ;
        RECT 98.800 247.700 104.400 248.300 ;
        RECT 98.800 247.600 99.600 247.700 ;
        RECT 103.600 247.600 104.400 247.700 ;
        RECT 143.600 248.300 144.400 248.400 ;
        RECT 146.800 248.300 147.600 248.400 ;
        RECT 143.600 247.700 147.600 248.300 ;
        RECT 143.600 247.600 144.400 247.700 ;
        RECT 146.800 247.600 147.600 247.700 ;
        RECT 159.600 248.300 160.400 248.400 ;
        RECT 175.600 248.300 176.400 248.400 ;
        RECT 193.200 248.300 194.000 248.400 ;
        RECT 159.600 247.700 194.000 248.300 ;
        RECT 159.600 247.600 160.400 247.700 ;
        RECT 175.600 247.600 176.400 247.700 ;
        RECT 193.200 247.600 194.000 247.700 ;
        RECT 452.400 248.300 453.200 248.400 ;
        RECT 455.600 248.300 456.400 248.400 ;
        RECT 452.400 247.700 456.400 248.300 ;
        RECT 452.400 247.600 453.200 247.700 ;
        RECT 455.600 247.600 456.400 247.700 ;
        RECT 457.200 248.300 458.000 248.400 ;
        RECT 460.400 248.300 461.200 248.400 ;
        RECT 457.200 247.700 461.200 248.300 ;
        RECT 457.200 247.600 458.000 247.700 ;
        RECT 460.400 247.600 461.200 247.700 ;
        RECT 554.800 248.300 555.600 248.400 ;
        RECT 566.000 248.300 566.800 248.400 ;
        RECT 554.800 247.700 566.800 248.300 ;
        RECT 554.800 247.600 555.600 247.700 ;
        RECT 566.000 247.600 566.800 247.700 ;
        RECT 180.400 246.300 181.200 246.400 ;
        RECT 185.200 246.300 186.000 246.400 ;
        RECT 180.400 245.700 186.000 246.300 ;
        RECT 180.400 245.600 181.200 245.700 ;
        RECT 185.200 245.600 186.000 245.700 ;
        RECT 449.200 246.300 450.000 246.400 ;
        RECT 468.400 246.300 469.200 246.400 ;
        RECT 449.200 245.700 469.200 246.300 ;
        RECT 449.200 245.600 450.000 245.700 ;
        RECT 468.400 245.600 469.200 245.700 ;
        RECT 146.800 243.600 147.600 244.400 ;
        RECT 439.600 244.300 440.400 244.400 ;
        RECT 482.800 244.300 483.600 244.400 ;
        RECT 439.600 243.700 483.600 244.300 ;
        RECT 439.600 243.600 440.400 243.700 ;
        RECT 482.800 243.600 483.600 243.700 ;
        RECT 151.600 242.300 152.400 242.400 ;
        RECT 182.000 242.300 182.800 242.400 ;
        RECT 151.600 241.700 182.800 242.300 ;
        RECT 151.600 241.600 152.400 241.700 ;
        RECT 182.000 241.600 182.800 241.700 ;
        RECT 450.800 242.300 451.600 242.400 ;
        RECT 474.800 242.300 475.600 242.400 ;
        RECT 450.800 241.700 475.600 242.300 ;
        RECT 450.800 241.600 451.600 241.700 ;
        RECT 474.800 241.600 475.600 241.700 ;
        RECT 455.600 240.300 456.400 240.400 ;
        RECT 466.800 240.300 467.600 240.400 ;
        RECT 455.600 239.700 467.600 240.300 ;
        RECT 455.600 239.600 456.400 239.700 ;
        RECT 466.800 239.600 467.600 239.700 ;
        RECT 110.000 238.300 110.800 238.400 ;
        RECT 130.800 238.300 131.600 238.400 ;
        RECT 110.000 237.700 131.600 238.300 ;
        RECT 110.000 237.600 110.800 237.700 ;
        RECT 130.800 237.600 131.600 237.700 ;
        RECT 433.200 238.300 434.000 238.400 ;
        RECT 465.200 238.300 466.000 238.400 ;
        RECT 433.200 237.700 466.000 238.300 ;
        RECT 433.200 237.600 434.000 237.700 ;
        RECT 465.200 237.600 466.000 237.700 ;
        RECT 401.200 236.300 402.000 236.400 ;
        RECT 425.200 236.300 426.000 236.400 ;
        RECT 462.000 236.300 462.800 236.400 ;
        RECT 401.200 235.700 462.800 236.300 ;
        RECT 401.200 235.600 402.000 235.700 ;
        RECT 425.200 235.600 426.000 235.700 ;
        RECT 462.000 235.600 462.800 235.700 ;
        RECT 55.600 234.300 56.400 234.400 ;
        RECT 84.400 234.300 85.200 234.400 ;
        RECT 55.600 233.700 85.200 234.300 ;
        RECT 55.600 233.600 56.400 233.700 ;
        RECT 84.400 233.600 85.200 233.700 ;
        RECT 129.200 234.300 130.000 234.400 ;
        RECT 156.400 234.300 157.200 234.400 ;
        RECT 129.200 233.700 157.200 234.300 ;
        RECT 129.200 233.600 130.000 233.700 ;
        RECT 156.400 233.600 157.200 233.700 ;
        RECT 210.800 234.300 211.600 234.400 ;
        RECT 238.000 234.300 238.800 234.400 ;
        RECT 210.800 233.700 238.800 234.300 ;
        RECT 210.800 233.600 211.600 233.700 ;
        RECT 238.000 233.600 238.800 233.700 ;
        RECT 297.200 234.300 298.000 234.400 ;
        RECT 327.600 234.300 328.400 234.400 ;
        RECT 297.200 233.700 328.400 234.300 ;
        RECT 297.200 233.600 298.000 233.700 ;
        RECT 327.600 233.600 328.400 233.700 ;
        RECT 430.000 234.300 430.800 234.400 ;
        RECT 442.800 234.300 443.600 234.400 ;
        RECT 430.000 233.700 443.600 234.300 ;
        RECT 430.000 233.600 430.800 233.700 ;
        RECT 442.800 233.600 443.600 233.700 ;
        RECT 455.600 234.300 456.400 234.400 ;
        RECT 476.400 234.300 477.200 234.400 ;
        RECT 498.800 234.300 499.600 234.400 ;
        RECT 455.600 233.700 499.600 234.300 ;
        RECT 455.600 233.600 456.400 233.700 ;
        RECT 476.400 233.600 477.200 233.700 ;
        RECT 498.800 233.600 499.600 233.700 ;
        RECT 79.600 232.300 80.400 232.400 ;
        RECT 92.400 232.300 93.200 232.400 ;
        RECT 79.600 231.700 93.200 232.300 ;
        RECT 79.600 231.600 80.400 231.700 ;
        RECT 92.400 231.600 93.200 231.700 ;
        RECT 140.400 232.300 141.200 232.400 ;
        RECT 153.200 232.300 154.000 232.400 ;
        RECT 140.400 231.700 154.000 232.300 ;
        RECT 140.400 231.600 141.200 231.700 ;
        RECT 153.200 231.600 154.000 231.700 ;
        RECT 230.000 232.300 230.800 232.400 ;
        RECT 239.600 232.300 240.400 232.400 ;
        RECT 230.000 231.700 240.400 232.300 ;
        RECT 230.000 231.600 230.800 231.700 ;
        RECT 239.600 231.600 240.400 231.700 ;
        RECT 305.200 232.300 306.000 232.400 ;
        RECT 338.800 232.300 339.600 232.400 ;
        RECT 305.200 231.700 339.600 232.300 ;
        RECT 305.200 231.600 306.000 231.700 ;
        RECT 338.800 231.600 339.600 231.700 ;
        RECT 438.000 232.300 438.800 232.400 ;
        RECT 442.800 232.300 443.600 232.400 ;
        RECT 452.400 232.300 453.200 232.400 ;
        RECT 458.800 232.300 459.600 232.400 ;
        RECT 438.000 231.700 459.600 232.300 ;
        RECT 438.000 231.600 438.800 231.700 ;
        RECT 442.800 231.600 443.600 231.700 ;
        RECT 452.400 231.600 453.200 231.700 ;
        RECT 458.800 231.600 459.600 231.700 ;
        RECT 465.200 232.300 466.000 232.400 ;
        RECT 470.000 232.300 470.800 232.400 ;
        RECT 465.200 231.700 470.800 232.300 ;
        RECT 465.200 231.600 466.000 231.700 ;
        RECT 470.000 231.600 470.800 231.700 ;
        RECT 486.000 232.300 486.800 232.400 ;
        RECT 495.600 232.300 496.400 232.400 ;
        RECT 486.000 231.700 496.400 232.300 ;
        RECT 486.000 231.600 486.800 231.700 ;
        RECT 495.600 231.600 496.400 231.700 ;
        RECT 508.400 232.300 509.200 232.400 ;
        RECT 514.800 232.300 515.600 232.400 ;
        RECT 508.400 231.700 515.600 232.300 ;
        RECT 508.400 231.600 509.200 231.700 ;
        RECT 514.800 231.600 515.600 231.700 ;
        RECT 551.600 232.300 552.400 232.400 ;
        RECT 558.000 232.300 558.800 232.400 ;
        RECT 551.600 231.700 558.800 232.300 ;
        RECT 551.600 231.600 552.400 231.700 ;
        RECT 558.000 231.600 558.800 231.700 ;
        RECT 38.000 230.300 38.800 230.400 ;
        RECT 41.200 230.300 42.000 230.400 ;
        RECT 38.000 229.700 42.000 230.300 ;
        RECT 38.000 229.600 38.800 229.700 ;
        RECT 41.200 229.600 42.000 229.700 ;
        RECT 153.200 230.300 154.000 230.400 ;
        RECT 158.000 230.300 158.800 230.400 ;
        RECT 153.200 229.700 158.800 230.300 ;
        RECT 153.200 229.600 154.000 229.700 ;
        RECT 158.000 229.600 158.800 229.700 ;
        RECT 159.600 230.300 160.400 230.400 ;
        RECT 185.200 230.300 186.000 230.400 ;
        RECT 159.600 229.700 186.000 230.300 ;
        RECT 159.600 229.600 160.400 229.700 ;
        RECT 185.200 229.600 186.000 229.700 ;
        RECT 196.400 230.300 197.200 230.400 ;
        RECT 204.400 230.300 205.200 230.400 ;
        RECT 223.600 230.300 224.400 230.400 ;
        RECT 246.000 230.300 246.800 230.400 ;
        RECT 196.400 229.700 246.800 230.300 ;
        RECT 196.400 229.600 197.200 229.700 ;
        RECT 204.400 229.600 205.200 229.700 ;
        RECT 223.600 229.600 224.400 229.700 ;
        RECT 246.000 229.600 246.800 229.700 ;
        RECT 284.400 230.300 285.200 230.400 ;
        RECT 294.000 230.300 294.800 230.400 ;
        RECT 284.400 229.700 294.800 230.300 ;
        RECT 284.400 229.600 285.200 229.700 ;
        RECT 294.000 229.600 294.800 229.700 ;
        RECT 295.600 230.300 296.400 230.400 ;
        RECT 306.800 230.300 307.600 230.400 ;
        RECT 295.600 229.700 307.600 230.300 ;
        RECT 295.600 229.600 296.400 229.700 ;
        RECT 306.800 229.600 307.600 229.700 ;
        RECT 362.800 230.300 363.600 230.400 ;
        RECT 375.600 230.300 376.400 230.400 ;
        RECT 362.800 229.700 376.400 230.300 ;
        RECT 362.800 229.600 363.600 229.700 ;
        RECT 375.600 229.600 376.400 229.700 ;
        RECT 394.800 230.300 395.600 230.400 ;
        RECT 404.400 230.300 405.200 230.400 ;
        RECT 394.800 229.700 405.200 230.300 ;
        RECT 394.800 229.600 395.600 229.700 ;
        RECT 404.400 229.600 405.200 229.700 ;
        RECT 436.400 230.300 437.200 230.400 ;
        RECT 449.200 230.300 450.000 230.400 ;
        RECT 497.200 230.300 498.000 230.400 ;
        RECT 436.400 229.700 498.000 230.300 ;
        RECT 436.400 229.600 437.200 229.700 ;
        RECT 449.200 229.600 450.000 229.700 ;
        RECT 497.200 229.600 498.000 229.700 ;
        RECT 521.200 230.300 522.000 230.400 ;
        RECT 538.800 230.300 539.600 230.400 ;
        RECT 521.200 229.700 539.600 230.300 ;
        RECT 521.200 229.600 522.000 229.700 ;
        RECT 538.800 229.600 539.600 229.700 ;
        RECT 76.400 228.300 77.200 228.400 ;
        RECT 81.200 228.300 82.000 228.400 ;
        RECT 76.400 227.700 82.000 228.300 ;
        RECT 76.400 227.600 77.200 227.700 ;
        RECT 81.200 227.600 82.000 227.700 ;
        RECT 121.200 228.300 122.000 228.400 ;
        RECT 151.600 228.300 152.400 228.400 ;
        RECT 121.200 227.700 152.400 228.300 ;
        RECT 121.200 227.600 122.000 227.700 ;
        RECT 151.600 227.600 152.400 227.700 ;
        RECT 238.000 228.300 238.800 228.400 ;
        RECT 249.200 228.300 250.000 228.400 ;
        RECT 238.000 227.700 250.000 228.300 ;
        RECT 238.000 227.600 238.800 227.700 ;
        RECT 249.200 227.600 250.000 227.700 ;
        RECT 463.600 227.600 464.400 228.400 ;
        RECT 492.400 228.300 493.200 228.400 ;
        RECT 511.600 228.300 512.400 228.400 ;
        RECT 554.800 228.300 555.600 228.400 ;
        RECT 492.400 227.700 555.600 228.300 ;
        RECT 492.400 227.600 493.200 227.700 ;
        RECT 511.600 227.600 512.400 227.700 ;
        RECT 554.800 227.600 555.600 227.700 ;
        RECT 281.200 226.300 282.000 226.400 ;
        RECT 302.000 226.300 302.800 226.400 ;
        RECT 281.200 225.700 302.800 226.300 ;
        RECT 281.200 225.600 282.000 225.700 ;
        RECT 302.000 225.600 302.800 225.700 ;
        RECT 434.800 226.300 435.600 226.400 ;
        RECT 438.000 226.300 438.800 226.400 ;
        RECT 444.400 226.300 445.200 226.400 ;
        RECT 434.800 225.700 445.200 226.300 ;
        RECT 434.800 225.600 435.600 225.700 ;
        RECT 438.000 225.600 438.800 225.700 ;
        RECT 444.400 225.600 445.200 225.700 ;
        RECT 457.200 225.600 458.000 226.400 ;
        RECT 458.800 226.300 459.600 226.400 ;
        RECT 479.600 226.300 480.400 226.400 ;
        RECT 458.800 225.700 480.400 226.300 ;
        RECT 458.800 225.600 459.600 225.700 ;
        RECT 479.600 225.600 480.400 225.700 ;
        RECT 495.600 226.300 496.400 226.400 ;
        RECT 502.000 226.300 502.800 226.400 ;
        RECT 495.600 225.700 502.800 226.300 ;
        RECT 495.600 225.600 496.400 225.700 ;
        RECT 502.000 225.600 502.800 225.700 ;
        RECT 1.200 224.300 2.000 224.400 ;
        RECT 2.800 224.300 3.600 224.400 ;
        RECT 1.200 223.700 3.600 224.300 ;
        RECT 1.200 223.600 2.000 223.700 ;
        RECT 2.800 223.600 3.600 223.700 ;
        RECT 79.600 224.300 80.400 224.400 ;
        RECT 92.400 224.300 93.200 224.400 ;
        RECT 79.600 223.700 93.200 224.300 ;
        RECT 79.600 223.600 80.400 223.700 ;
        RECT 92.400 223.600 93.200 223.700 ;
        RECT 191.600 224.300 192.400 224.400 ;
        RECT 198.000 224.300 198.800 224.400 ;
        RECT 191.600 223.700 198.800 224.300 ;
        RECT 191.600 223.600 192.400 223.700 ;
        RECT 198.000 223.600 198.800 223.700 ;
        RECT 217.200 224.300 218.000 224.400 ;
        RECT 236.400 224.300 237.200 224.400 ;
        RECT 217.200 223.700 237.200 224.300 ;
        RECT 217.200 223.600 218.000 223.700 ;
        RECT 236.400 223.600 237.200 223.700 ;
        RECT 262.000 224.300 262.800 224.400 ;
        RECT 273.200 224.300 274.000 224.400 ;
        RECT 284.400 224.300 285.200 224.400 ;
        RECT 262.000 223.700 285.200 224.300 ;
        RECT 262.000 223.600 262.800 223.700 ;
        RECT 273.200 223.600 274.000 223.700 ;
        RECT 284.400 223.600 285.200 223.700 ;
        RECT 326.000 224.300 326.800 224.400 ;
        RECT 332.400 224.300 333.200 224.400 ;
        RECT 326.000 223.700 333.200 224.300 ;
        RECT 326.000 223.600 326.800 223.700 ;
        RECT 332.400 223.600 333.200 223.700 ;
        RECT 345.200 224.300 346.000 224.400 ;
        RECT 364.400 224.300 365.200 224.400 ;
        RECT 345.200 223.700 365.200 224.300 ;
        RECT 345.200 223.600 346.000 223.700 ;
        RECT 364.400 223.600 365.200 223.700 ;
        RECT 428.400 224.300 429.200 224.400 ;
        RECT 473.200 224.300 474.000 224.400 ;
        RECT 428.400 223.700 474.000 224.300 ;
        RECT 428.400 223.600 429.200 223.700 ;
        RECT 473.200 223.600 474.000 223.700 ;
        RECT 486.000 224.300 486.800 224.400 ;
        RECT 489.200 224.300 490.000 224.400 ;
        RECT 486.000 223.700 490.000 224.300 ;
        RECT 486.000 223.600 486.800 223.700 ;
        RECT 489.200 223.600 490.000 223.700 ;
        RECT 510.000 224.300 510.800 224.400 ;
        RECT 524.400 224.300 525.200 224.400 ;
        RECT 510.000 223.700 525.200 224.300 ;
        RECT 510.000 223.600 510.800 223.700 ;
        RECT 524.400 223.600 525.200 223.700 ;
        RECT 54.000 222.300 54.800 222.400 ;
        RECT 65.200 222.300 66.000 222.400 ;
        RECT 54.000 221.700 66.000 222.300 ;
        RECT 54.000 221.600 54.800 221.700 ;
        RECT 65.200 221.600 66.000 221.700 ;
        RECT 89.200 222.300 90.000 222.400 ;
        RECT 97.200 222.300 98.000 222.400 ;
        RECT 89.200 221.700 98.000 222.300 ;
        RECT 89.200 221.600 90.000 221.700 ;
        RECT 97.200 221.600 98.000 221.700 ;
        RECT 103.600 222.300 104.400 222.400 ;
        RECT 116.400 222.300 117.200 222.400 ;
        RECT 103.600 221.700 117.200 222.300 ;
        RECT 103.600 221.600 104.400 221.700 ;
        RECT 116.400 221.600 117.200 221.700 ;
        RECT 314.800 222.300 315.600 222.400 ;
        RECT 326.000 222.300 326.800 222.400 ;
        RECT 314.800 221.700 326.800 222.300 ;
        RECT 314.800 221.600 315.600 221.700 ;
        RECT 326.000 221.600 326.800 221.700 ;
        RECT 474.800 222.300 475.600 222.400 ;
        RECT 497.200 222.300 498.000 222.400 ;
        RECT 474.800 221.700 498.000 222.300 ;
        RECT 474.800 221.600 475.600 221.700 ;
        RECT 497.200 221.600 498.000 221.700 ;
        RECT 52.400 220.300 53.200 220.400 ;
        RECT 57.200 220.300 58.000 220.400 ;
        RECT 52.400 219.700 58.000 220.300 ;
        RECT 52.400 219.600 53.200 219.700 ;
        RECT 57.200 219.600 58.000 219.700 ;
        RECT 442.800 220.300 443.600 220.400 ;
        RECT 452.400 220.300 453.200 220.400 ;
        RECT 458.800 220.300 459.600 220.400 ;
        RECT 442.800 219.700 459.600 220.300 ;
        RECT 442.800 219.600 443.600 219.700 ;
        RECT 452.400 219.600 453.200 219.700 ;
        RECT 458.800 219.600 459.600 219.700 ;
        RECT 470.000 220.300 470.800 220.400 ;
        RECT 494.000 220.300 494.800 220.400 ;
        RECT 470.000 219.700 494.800 220.300 ;
        RECT 470.000 219.600 470.800 219.700 ;
        RECT 494.000 219.600 494.800 219.700 ;
        RECT 180.400 218.300 181.200 218.400 ;
        RECT 204.400 218.300 205.200 218.400 ;
        RECT 180.400 217.700 205.200 218.300 ;
        RECT 180.400 217.600 181.200 217.700 ;
        RECT 204.400 217.600 205.200 217.700 ;
        RECT 220.400 218.300 221.200 218.400 ;
        RECT 225.200 218.300 226.000 218.400 ;
        RECT 220.400 217.700 226.000 218.300 ;
        RECT 220.400 217.600 221.200 217.700 ;
        RECT 225.200 217.600 226.000 217.700 ;
        RECT 271.600 218.300 272.400 218.400 ;
        RECT 282.800 218.300 283.600 218.400 ;
        RECT 271.600 217.700 283.600 218.300 ;
        RECT 271.600 217.600 272.400 217.700 ;
        RECT 282.800 217.600 283.600 217.700 ;
        RECT 284.400 218.300 285.200 218.400 ;
        RECT 294.000 218.300 294.800 218.400 ;
        RECT 284.400 217.700 294.800 218.300 ;
        RECT 284.400 217.600 285.200 217.700 ;
        RECT 294.000 217.600 294.800 217.700 ;
        RECT 329.200 218.300 330.000 218.400 ;
        RECT 370.800 218.300 371.600 218.400 ;
        RECT 329.200 217.700 371.600 218.300 ;
        RECT 329.200 217.600 330.000 217.700 ;
        RECT 370.800 217.600 371.600 217.700 ;
        RECT 26.800 216.300 27.600 216.400 ;
        RECT 34.800 216.300 35.600 216.400 ;
        RECT 26.800 215.700 35.600 216.300 ;
        RECT 26.800 215.600 27.600 215.700 ;
        RECT 34.800 215.600 35.600 215.700 ;
        RECT 164.400 216.300 165.200 216.400 ;
        RECT 174.000 216.300 174.800 216.400 ;
        RECT 188.400 216.300 189.200 216.400 ;
        RECT 164.400 215.700 189.200 216.300 ;
        RECT 164.400 215.600 165.200 215.700 ;
        RECT 174.000 215.600 174.800 215.700 ;
        RECT 188.400 215.600 189.200 215.700 ;
        RECT 292.400 216.300 293.200 216.400 ;
        RECT 298.800 216.300 299.600 216.400 ;
        RECT 292.400 215.700 299.600 216.300 ;
        RECT 292.400 215.600 293.200 215.700 ;
        RECT 298.800 215.600 299.600 215.700 ;
        RECT 335.600 216.300 336.400 216.400 ;
        RECT 342.000 216.300 342.800 216.400 ;
        RECT 335.600 215.700 342.800 216.300 ;
        RECT 335.600 215.600 336.400 215.700 ;
        RECT 342.000 215.600 342.800 215.700 ;
        RECT 380.400 216.300 381.200 216.400 ;
        RECT 393.200 216.300 394.000 216.400 ;
        RECT 380.400 215.700 394.000 216.300 ;
        RECT 380.400 215.600 381.200 215.700 ;
        RECT 393.200 215.600 394.000 215.700 ;
        RECT 457.200 216.300 458.000 216.400 ;
        RECT 465.200 216.300 466.000 216.400 ;
        RECT 476.400 216.300 477.200 216.400 ;
        RECT 487.600 216.300 488.400 216.400 ;
        RECT 457.200 215.700 488.400 216.300 ;
        RECT 457.200 215.600 458.000 215.700 ;
        RECT 465.200 215.600 466.000 215.700 ;
        RECT 476.400 215.600 477.200 215.700 ;
        RECT 487.600 215.600 488.400 215.700 ;
        RECT 490.800 216.300 491.600 216.400 ;
        RECT 498.800 216.300 499.600 216.400 ;
        RECT 490.800 215.700 499.600 216.300 ;
        RECT 490.800 215.600 491.600 215.700 ;
        RECT 498.800 215.600 499.600 215.700 ;
        RECT 524.400 216.300 525.200 216.400 ;
        RECT 529.200 216.300 530.000 216.400 ;
        RECT 524.400 215.700 530.000 216.300 ;
        RECT 524.400 215.600 525.200 215.700 ;
        RECT 529.200 215.600 530.000 215.700 ;
        RECT 12.400 214.300 13.200 214.400 ;
        RECT 31.600 214.300 32.400 214.400 ;
        RECT 55.600 214.300 56.400 214.400 ;
        RECT 70.000 214.300 70.800 214.400 ;
        RECT 94.000 214.300 94.800 214.400 ;
        RECT 97.200 214.300 98.000 214.400 ;
        RECT 106.800 214.300 107.600 214.400 ;
        RECT 118.000 214.300 118.800 214.400 ;
        RECT 12.400 213.700 118.800 214.300 ;
        RECT 12.400 213.600 13.200 213.700 ;
        RECT 31.600 213.600 32.400 213.700 ;
        RECT 55.600 213.600 56.400 213.700 ;
        RECT 70.000 213.600 70.800 213.700 ;
        RECT 94.000 213.600 94.800 213.700 ;
        RECT 97.200 213.600 98.000 213.700 ;
        RECT 106.800 213.600 107.600 213.700 ;
        RECT 118.000 213.600 118.800 213.700 ;
        RECT 177.200 214.300 178.000 214.400 ;
        RECT 182.000 214.300 182.800 214.400 ;
        RECT 177.200 213.700 182.800 214.300 ;
        RECT 177.200 213.600 178.000 213.700 ;
        RECT 182.000 213.600 182.800 213.700 ;
        RECT 183.600 214.300 184.400 214.400 ;
        RECT 193.200 214.300 194.000 214.400 ;
        RECT 207.600 214.300 208.400 214.400 ;
        RECT 183.600 213.700 208.400 214.300 ;
        RECT 183.600 213.600 184.400 213.700 ;
        RECT 193.200 213.600 194.000 213.700 ;
        RECT 207.600 213.600 208.400 213.700 ;
        RECT 230.000 214.300 230.800 214.400 ;
        RECT 234.800 214.300 235.600 214.400 ;
        RECT 230.000 213.700 235.600 214.300 ;
        RECT 230.000 213.600 230.800 213.700 ;
        RECT 234.800 213.600 235.600 213.700 ;
        RECT 246.000 214.300 246.800 214.400 ;
        RECT 258.800 214.300 259.600 214.400 ;
        RECT 246.000 213.700 259.600 214.300 ;
        RECT 246.000 213.600 246.800 213.700 ;
        RECT 258.800 213.600 259.600 213.700 ;
        RECT 310.000 214.300 310.800 214.400 ;
        RECT 329.200 214.300 330.000 214.400 ;
        RECT 348.400 214.300 349.200 214.400 ;
        RECT 310.000 213.700 349.200 214.300 ;
        RECT 310.000 213.600 310.800 213.700 ;
        RECT 329.200 213.600 330.000 213.700 ;
        RECT 348.400 213.600 349.200 213.700 ;
        RECT 366.000 214.300 366.800 214.400 ;
        RECT 375.600 214.300 376.400 214.400 ;
        RECT 366.000 213.700 376.400 214.300 ;
        RECT 366.000 213.600 366.800 213.700 ;
        RECT 375.600 213.600 376.400 213.700 ;
        RECT 457.200 213.600 458.000 214.400 ;
        RECT 465.200 214.300 466.000 214.400 ;
        RECT 482.800 214.300 483.600 214.400 ;
        RECT 465.200 213.700 483.600 214.300 ;
        RECT 465.200 213.600 466.000 213.700 ;
        RECT 482.800 213.600 483.600 213.700 ;
        RECT 489.200 214.300 490.000 214.400 ;
        RECT 495.600 214.300 496.400 214.400 ;
        RECT 489.200 213.700 496.400 214.300 ;
        RECT 489.200 213.600 490.000 213.700 ;
        RECT 495.600 213.600 496.400 213.700 ;
        RECT 497.200 214.300 498.000 214.400 ;
        RECT 500.400 214.300 501.200 214.400 ;
        RECT 497.200 213.700 501.200 214.300 ;
        RECT 497.200 213.600 498.000 213.700 ;
        RECT 500.400 213.600 501.200 213.700 ;
        RECT 513.200 214.300 514.000 214.400 ;
        RECT 530.800 214.300 531.600 214.400 ;
        RECT 537.200 214.300 538.000 214.400 ;
        RECT 513.200 213.700 538.000 214.300 ;
        RECT 513.200 213.600 514.000 213.700 ;
        RECT 530.800 213.600 531.600 213.700 ;
        RECT 537.200 213.600 538.000 213.700 ;
        RECT 6.000 211.600 6.800 212.400 ;
        RECT 124.400 212.300 125.200 212.400 ;
        RECT 127.600 212.300 128.400 212.400 ;
        RECT 124.400 211.700 128.400 212.300 ;
        RECT 124.400 211.600 125.200 211.700 ;
        RECT 127.600 211.600 128.400 211.700 ;
        RECT 146.800 212.300 147.600 212.400 ;
        RECT 156.400 212.300 157.200 212.400 ;
        RECT 166.000 212.300 166.800 212.400 ;
        RECT 170.800 212.300 171.600 212.400 ;
        RECT 146.800 211.700 171.600 212.300 ;
        RECT 146.800 211.600 147.600 211.700 ;
        RECT 156.400 211.600 157.200 211.700 ;
        RECT 166.000 211.600 166.800 211.700 ;
        RECT 170.800 211.600 171.600 211.700 ;
        RECT 193.200 212.300 194.000 212.400 ;
        RECT 198.000 212.300 198.800 212.400 ;
        RECT 193.200 211.700 198.800 212.300 ;
        RECT 193.200 211.600 194.000 211.700 ;
        RECT 198.000 211.600 198.800 211.700 ;
        RECT 217.200 212.300 218.000 212.400 ;
        RECT 222.000 212.300 222.800 212.400 ;
        RECT 217.200 211.700 222.800 212.300 ;
        RECT 217.200 211.600 218.000 211.700 ;
        RECT 222.000 211.600 222.800 211.700 ;
        RECT 226.800 212.300 227.600 212.400 ;
        RECT 241.200 212.300 242.000 212.400 ;
        RECT 247.600 212.300 248.400 212.400 ;
        RECT 226.800 211.700 248.400 212.300 ;
        RECT 226.800 211.600 227.600 211.700 ;
        RECT 241.200 211.600 242.000 211.700 ;
        RECT 247.600 211.600 248.400 211.700 ;
        RECT 265.200 212.300 266.000 212.400 ;
        RECT 276.400 212.300 277.200 212.400 ;
        RECT 265.200 211.700 277.200 212.300 ;
        RECT 265.200 211.600 266.000 211.700 ;
        RECT 276.400 211.600 277.200 211.700 ;
        RECT 279.600 212.300 280.400 212.400 ;
        RECT 284.400 212.300 285.200 212.400 ;
        RECT 279.600 211.700 285.200 212.300 ;
        RECT 279.600 211.600 280.400 211.700 ;
        RECT 284.400 211.600 285.200 211.700 ;
        RECT 311.600 212.300 312.400 212.400 ;
        RECT 318.000 212.300 318.800 212.400 ;
        RECT 311.600 211.700 318.800 212.300 ;
        RECT 311.600 211.600 312.400 211.700 ;
        RECT 318.000 211.600 318.800 211.700 ;
        RECT 338.800 212.300 339.600 212.400 ;
        RECT 377.200 212.300 378.000 212.400 ;
        RECT 338.800 211.700 378.000 212.300 ;
        RECT 338.800 211.600 339.600 211.700 ;
        RECT 377.200 211.600 378.000 211.700 ;
        RECT 396.400 212.300 397.200 212.400 ;
        RECT 399.600 212.300 400.400 212.400 ;
        RECT 396.400 211.700 400.400 212.300 ;
        RECT 396.400 211.600 397.200 211.700 ;
        RECT 399.600 211.600 400.400 211.700 ;
        RECT 412.400 212.300 413.200 212.400 ;
        RECT 415.600 212.300 416.400 212.400 ;
        RECT 412.400 211.700 416.400 212.300 ;
        RECT 412.400 211.600 413.200 211.700 ;
        RECT 415.600 211.600 416.400 211.700 ;
        RECT 433.200 212.300 434.000 212.400 ;
        RECT 439.600 212.300 440.400 212.400 ;
        RECT 458.800 212.300 459.600 212.400 ;
        RECT 433.200 211.700 459.600 212.300 ;
        RECT 433.200 211.600 434.000 211.700 ;
        RECT 439.600 211.600 440.400 211.700 ;
        RECT 458.800 211.600 459.600 211.700 ;
        RECT 463.600 212.300 464.400 212.400 ;
        RECT 474.800 212.300 475.600 212.400 ;
        RECT 463.600 211.700 475.600 212.300 ;
        RECT 463.600 211.600 464.400 211.700 ;
        RECT 474.800 211.600 475.600 211.700 ;
        RECT 476.400 212.300 477.200 212.400 ;
        RECT 492.400 212.300 493.200 212.400 ;
        RECT 476.400 211.700 493.200 212.300 ;
        RECT 476.400 211.600 477.200 211.700 ;
        RECT 492.400 211.600 493.200 211.700 ;
        RECT 497.200 212.300 498.000 212.400 ;
        RECT 508.400 212.300 509.200 212.400 ;
        RECT 497.200 211.700 509.200 212.300 ;
        RECT 497.200 211.600 498.000 211.700 ;
        RECT 508.400 211.600 509.200 211.700 ;
        RECT 521.200 212.300 522.000 212.400 ;
        RECT 527.600 212.300 528.400 212.400 ;
        RECT 534.000 212.300 534.800 212.400 ;
        RECT 521.200 211.700 534.800 212.300 ;
        RECT 521.200 211.600 522.000 211.700 ;
        RECT 527.600 211.600 528.400 211.700 ;
        RECT 534.000 211.600 534.800 211.700 ;
        RECT 186.800 210.300 187.600 210.400 ;
        RECT 196.400 210.300 197.200 210.400 ;
        RECT 186.800 209.700 197.200 210.300 ;
        RECT 186.800 209.600 187.600 209.700 ;
        RECT 196.400 209.600 197.200 209.700 ;
        RECT 233.200 210.300 234.000 210.400 ;
        RECT 249.200 210.300 250.000 210.400 ;
        RECT 273.200 210.300 274.000 210.400 ;
        RECT 233.200 209.700 274.000 210.300 ;
        RECT 233.200 209.600 234.000 209.700 ;
        RECT 249.200 209.600 250.000 209.700 ;
        RECT 273.200 209.600 274.000 209.700 ;
        RECT 281.200 210.300 282.000 210.400 ;
        RECT 284.400 210.300 285.200 210.400 ;
        RECT 281.200 209.700 285.200 210.300 ;
        RECT 281.200 209.600 282.000 209.700 ;
        RECT 284.400 209.600 285.200 209.700 ;
        RECT 380.400 210.300 381.200 210.400 ;
        RECT 399.600 210.300 400.400 210.400 ;
        RECT 418.800 210.300 419.600 210.400 ;
        RECT 380.400 209.700 398.700 210.300 ;
        RECT 380.400 209.600 381.200 209.700 ;
        RECT 188.400 208.300 189.200 208.400 ;
        RECT 201.200 208.300 202.000 208.400 ;
        RECT 188.400 207.700 202.000 208.300 ;
        RECT 188.400 207.600 189.200 207.700 ;
        RECT 201.200 207.600 202.000 207.700 ;
        RECT 246.000 208.300 246.800 208.400 ;
        RECT 249.200 208.300 250.000 208.400 ;
        RECT 246.000 207.700 250.000 208.300 ;
        RECT 246.000 207.600 246.800 207.700 ;
        RECT 249.200 207.600 250.000 207.700 ;
        RECT 265.200 208.300 266.000 208.400 ;
        RECT 270.000 208.300 270.800 208.400 ;
        RECT 265.200 207.700 270.800 208.300 ;
        RECT 265.200 207.600 266.000 207.700 ;
        RECT 270.000 207.600 270.800 207.700 ;
        RECT 370.800 208.300 371.600 208.400 ;
        RECT 396.400 208.300 397.200 208.400 ;
        RECT 370.800 207.700 397.200 208.300 ;
        RECT 398.100 208.300 398.700 209.700 ;
        RECT 399.600 209.700 419.600 210.300 ;
        RECT 399.600 209.600 400.400 209.700 ;
        RECT 418.800 209.600 419.600 209.700 ;
        RECT 444.400 210.300 445.200 210.400 ;
        RECT 463.600 210.300 464.400 210.400 ;
        RECT 444.400 209.700 464.400 210.300 ;
        RECT 444.400 209.600 445.200 209.700 ;
        RECT 463.600 209.600 464.400 209.700 ;
        RECT 482.800 210.300 483.600 210.400 ;
        RECT 486.000 210.300 486.800 210.400 ;
        RECT 482.800 209.700 486.800 210.300 ;
        RECT 482.800 209.600 483.600 209.700 ;
        RECT 486.000 209.600 486.800 209.700 ;
        RECT 538.800 210.300 539.600 210.400 ;
        RECT 542.000 210.300 542.800 210.400 ;
        RECT 538.800 209.700 542.800 210.300 ;
        RECT 538.800 209.600 539.600 209.700 ;
        RECT 542.000 209.600 542.800 209.700 ;
        RECT 410.800 208.300 411.600 208.400 ;
        RECT 398.100 207.700 411.600 208.300 ;
        RECT 370.800 207.600 371.600 207.700 ;
        RECT 396.400 207.600 397.200 207.700 ;
        RECT 410.800 207.600 411.600 207.700 ;
        RECT 431.600 208.300 432.400 208.400 ;
        RECT 466.800 208.300 467.600 208.400 ;
        RECT 431.600 207.700 467.600 208.300 ;
        RECT 431.600 207.600 432.400 207.700 ;
        RECT 466.800 207.600 467.600 207.700 ;
        RECT 474.800 208.300 475.600 208.400 ;
        RECT 479.600 208.300 480.400 208.400 ;
        RECT 502.000 208.300 502.800 208.400 ;
        RECT 474.800 207.700 502.800 208.300 ;
        RECT 474.800 207.600 475.600 207.700 ;
        RECT 479.600 207.600 480.400 207.700 ;
        RECT 502.000 207.600 502.800 207.700 ;
        RECT 505.200 208.300 506.000 208.400 ;
        RECT 548.400 208.300 549.200 208.400 ;
        RECT 505.200 207.700 549.200 208.300 ;
        RECT 505.200 207.600 506.000 207.700 ;
        RECT 548.400 207.600 549.200 207.700 ;
        RECT 561.200 208.300 562.000 208.400 ;
        RECT 569.200 208.300 570.000 208.400 ;
        RECT 561.200 207.700 570.000 208.300 ;
        RECT 561.200 207.600 562.000 207.700 ;
        RECT 569.200 207.600 570.000 207.700 ;
        RECT 239.600 206.300 240.400 206.400 ;
        RECT 249.200 206.300 250.000 206.400 ;
        RECT 239.600 205.700 250.000 206.300 ;
        RECT 239.600 205.600 240.400 205.700 ;
        RECT 249.200 205.600 250.000 205.700 ;
        RECT 466.800 206.300 467.600 206.400 ;
        RECT 481.200 206.300 482.000 206.400 ;
        RECT 466.800 205.700 482.000 206.300 ;
        RECT 466.800 205.600 467.600 205.700 ;
        RECT 481.200 205.600 482.000 205.700 ;
        RECT 39.600 204.300 40.400 204.400 ;
        RECT 44.400 204.300 45.200 204.400 ;
        RECT 39.600 203.700 45.200 204.300 ;
        RECT 39.600 203.600 40.400 203.700 ;
        RECT 44.400 203.600 45.200 203.700 ;
        RECT 111.600 203.600 112.400 204.400 ;
        RECT 252.400 204.300 253.200 204.400 ;
        RECT 298.800 204.300 299.600 204.400 ;
        RECT 252.400 203.700 299.600 204.300 ;
        RECT 252.400 203.600 253.200 203.700 ;
        RECT 298.800 203.600 299.600 203.700 ;
        RECT 436.400 204.300 437.200 204.400 ;
        RECT 439.600 204.300 440.400 204.400 ;
        RECT 465.200 204.300 466.000 204.400 ;
        RECT 470.000 204.300 470.800 204.400 ;
        RECT 474.800 204.300 475.600 204.400 ;
        RECT 436.400 203.700 475.600 204.300 ;
        RECT 436.400 203.600 437.200 203.700 ;
        RECT 439.600 203.600 440.400 203.700 ;
        RECT 465.200 203.600 466.000 203.700 ;
        RECT 470.000 203.600 470.800 203.700 ;
        RECT 474.800 203.600 475.600 203.700 ;
        RECT 462.000 200.300 462.800 200.400 ;
        RECT 468.400 200.300 469.200 200.400 ;
        RECT 462.000 199.700 469.200 200.300 ;
        RECT 462.000 199.600 462.800 199.700 ;
        RECT 468.400 199.600 469.200 199.700 ;
        RECT 481.200 200.300 482.000 200.400 ;
        RECT 486.000 200.300 486.800 200.400 ;
        RECT 498.800 200.300 499.600 200.400 ;
        RECT 527.600 200.300 528.400 200.400 ;
        RECT 481.200 199.700 528.400 200.300 ;
        RECT 481.200 199.600 482.000 199.700 ;
        RECT 486.000 199.600 486.800 199.700 ;
        RECT 498.800 199.600 499.600 199.700 ;
        RECT 527.600 199.600 528.400 199.700 ;
        RECT 401.200 198.300 402.000 198.400 ;
        RECT 409.200 198.300 410.000 198.400 ;
        RECT 401.200 197.700 410.000 198.300 ;
        RECT 401.200 197.600 402.000 197.700 ;
        RECT 409.200 197.600 410.000 197.700 ;
        RECT 76.400 196.300 77.200 196.400 ;
        RECT 87.600 196.300 88.400 196.400 ;
        RECT 121.200 196.300 122.000 196.400 ;
        RECT 76.400 195.700 122.000 196.300 ;
        RECT 76.400 195.600 77.200 195.700 ;
        RECT 87.600 195.600 88.400 195.700 ;
        RECT 121.200 195.600 122.000 195.700 ;
        RECT 186.800 196.300 187.600 196.400 ;
        RECT 190.000 196.300 190.800 196.400 ;
        RECT 186.800 195.700 190.800 196.300 ;
        RECT 186.800 195.600 187.600 195.700 ;
        RECT 190.000 195.600 190.800 195.700 ;
        RECT 198.000 196.300 198.800 196.400 ;
        RECT 223.600 196.300 224.400 196.400 ;
        RECT 198.000 195.700 224.400 196.300 ;
        RECT 198.000 195.600 198.800 195.700 ;
        RECT 223.600 195.600 224.400 195.700 ;
        RECT 34.800 194.300 35.600 194.400 ;
        RECT 42.800 194.300 43.600 194.400 ;
        RECT 34.800 193.700 43.600 194.300 ;
        RECT 34.800 193.600 35.600 193.700 ;
        RECT 42.800 193.600 43.600 193.700 ;
        RECT 202.800 194.300 203.600 194.400 ;
        RECT 230.000 194.300 230.800 194.400 ;
        RECT 202.800 193.700 230.800 194.300 ;
        RECT 202.800 193.600 203.600 193.700 ;
        RECT 230.000 193.600 230.800 193.700 ;
        RECT 306.800 194.300 307.600 194.400 ;
        RECT 321.200 194.300 322.000 194.400 ;
        RECT 306.800 193.700 322.000 194.300 ;
        RECT 306.800 193.600 307.600 193.700 ;
        RECT 321.200 193.600 322.000 193.700 ;
        RECT 42.800 192.300 43.600 192.400 ;
        RECT 49.200 192.300 50.000 192.400 ;
        RECT 55.600 192.300 56.400 192.400 ;
        RECT 42.800 191.700 56.400 192.300 ;
        RECT 42.800 191.600 43.600 191.700 ;
        RECT 49.200 191.600 50.000 191.700 ;
        RECT 55.600 191.600 56.400 191.700 ;
        RECT 68.400 192.300 69.200 192.400 ;
        RECT 78.000 192.300 78.800 192.400 ;
        RECT 68.400 191.700 78.800 192.300 ;
        RECT 68.400 191.600 69.200 191.700 ;
        RECT 78.000 191.600 78.800 191.700 ;
        RECT 86.000 192.300 86.800 192.400 ;
        RECT 110.000 192.300 110.800 192.400 ;
        RECT 86.000 191.700 110.800 192.300 ;
        RECT 86.000 191.600 86.800 191.700 ;
        RECT 110.000 191.600 110.800 191.700 ;
        RECT 191.600 192.300 192.400 192.400 ;
        RECT 199.600 192.300 200.400 192.400 ;
        RECT 191.600 191.700 200.400 192.300 ;
        RECT 191.600 191.600 192.400 191.700 ;
        RECT 199.600 191.600 200.400 191.700 ;
        RECT 217.200 192.300 218.000 192.400 ;
        RECT 226.800 192.300 227.600 192.400 ;
        RECT 217.200 191.700 227.600 192.300 ;
        RECT 217.200 191.600 218.000 191.700 ;
        RECT 226.800 191.600 227.600 191.700 ;
        RECT 255.600 192.300 256.400 192.400 ;
        RECT 302.000 192.300 302.800 192.400 ;
        RECT 255.600 191.700 302.800 192.300 ;
        RECT 255.600 191.600 256.400 191.700 ;
        RECT 302.000 191.600 302.800 191.700 ;
        RECT 303.600 192.300 304.400 192.400 ;
        RECT 311.600 192.300 312.400 192.400 ;
        RECT 303.600 191.700 312.400 192.300 ;
        RECT 303.600 191.600 304.400 191.700 ;
        RECT 311.600 191.600 312.400 191.700 ;
        RECT 452.400 192.300 453.200 192.400 ;
        RECT 454.000 192.300 454.800 192.400 ;
        RECT 452.400 191.700 454.800 192.300 ;
        RECT 452.400 191.600 453.200 191.700 ;
        RECT 454.000 191.600 454.800 191.700 ;
        RECT 511.600 192.300 512.400 192.400 ;
        RECT 514.800 192.300 515.600 192.400 ;
        RECT 518.000 192.300 518.800 192.400 ;
        RECT 511.600 191.700 518.800 192.300 ;
        RECT 511.600 191.600 512.400 191.700 ;
        RECT 514.800 191.600 515.600 191.700 ;
        RECT 518.000 191.600 518.800 191.700 ;
        RECT 519.600 192.300 520.400 192.400 ;
        RECT 548.400 192.300 549.200 192.400 ;
        RECT 519.600 191.700 549.200 192.300 ;
        RECT 519.600 191.600 520.400 191.700 ;
        RECT 548.400 191.600 549.200 191.700 ;
        RECT 39.600 190.300 40.400 190.400 ;
        RECT 63.600 190.300 64.400 190.400 ;
        RECT 39.600 189.700 64.400 190.300 ;
        RECT 39.600 189.600 40.400 189.700 ;
        RECT 63.600 189.600 64.400 189.700 ;
        RECT 65.200 190.300 66.000 190.400 ;
        RECT 66.800 190.300 67.600 190.400 ;
        RECT 94.000 190.300 94.800 190.400 ;
        RECT 65.200 189.700 94.800 190.300 ;
        RECT 65.200 189.600 66.000 189.700 ;
        RECT 66.800 189.600 67.600 189.700 ;
        RECT 94.000 189.600 94.800 189.700 ;
        RECT 129.200 190.300 130.000 190.400 ;
        RECT 143.600 190.300 144.400 190.400 ;
        RECT 129.200 189.700 144.400 190.300 ;
        RECT 129.200 189.600 130.000 189.700 ;
        RECT 143.600 189.600 144.400 189.700 ;
        RECT 146.800 190.300 147.600 190.400 ;
        RECT 151.600 190.300 152.400 190.400 ;
        RECT 146.800 189.700 152.400 190.300 ;
        RECT 146.800 189.600 147.600 189.700 ;
        RECT 151.600 189.600 152.400 189.700 ;
        RECT 180.400 190.300 181.200 190.400 ;
        RECT 191.600 190.300 192.400 190.400 ;
        RECT 180.400 189.700 192.400 190.300 ;
        RECT 180.400 189.600 181.200 189.700 ;
        RECT 191.600 189.600 192.400 189.700 ;
        RECT 217.200 190.300 218.000 190.400 ;
        RECT 279.600 190.300 280.400 190.400 ;
        RECT 217.200 189.700 280.400 190.300 ;
        RECT 217.200 189.600 218.000 189.700 ;
        RECT 279.600 189.600 280.400 189.700 ;
        RECT 372.400 190.300 373.200 190.400 ;
        RECT 377.200 190.300 378.000 190.400 ;
        RECT 372.400 189.700 378.000 190.300 ;
        RECT 372.400 189.600 373.200 189.700 ;
        RECT 377.200 189.600 378.000 189.700 ;
        RECT 382.000 190.300 382.800 190.400 ;
        RECT 385.200 190.300 386.000 190.400 ;
        RECT 382.000 189.700 386.000 190.300 ;
        RECT 382.000 189.600 382.800 189.700 ;
        RECT 385.200 189.600 386.000 189.700 ;
        RECT 393.200 190.300 394.000 190.400 ;
        RECT 407.600 190.300 408.400 190.400 ;
        RECT 393.200 189.700 408.400 190.300 ;
        RECT 393.200 189.600 394.000 189.700 ;
        RECT 407.600 189.600 408.400 189.700 ;
        RECT 430.000 190.300 430.800 190.400 ;
        RECT 433.200 190.300 434.000 190.400 ;
        RECT 430.000 189.700 434.000 190.300 ;
        RECT 430.000 189.600 430.800 189.700 ;
        RECT 433.200 189.600 434.000 189.700 ;
        RECT 438.000 190.300 438.800 190.400 ;
        RECT 454.000 190.300 454.800 190.400 ;
        RECT 462.000 190.300 462.800 190.400 ;
        RECT 438.000 189.700 462.800 190.300 ;
        RECT 438.000 189.600 438.800 189.700 ;
        RECT 454.000 189.600 454.800 189.700 ;
        RECT 462.000 189.600 462.800 189.700 ;
        RECT 478.000 190.300 478.800 190.400 ;
        RECT 487.600 190.300 488.400 190.400 ;
        RECT 478.000 189.700 488.400 190.300 ;
        RECT 478.000 189.600 478.800 189.700 ;
        RECT 487.600 189.600 488.400 189.700 ;
        RECT 516.400 190.300 517.200 190.400 ;
        RECT 538.800 190.300 539.600 190.400 ;
        RECT 516.400 189.700 539.600 190.300 ;
        RECT 516.400 189.600 517.200 189.700 ;
        RECT 538.800 189.600 539.600 189.700 ;
        RECT 558.000 190.300 558.800 190.400 ;
        RECT 570.800 190.300 571.600 190.400 ;
        RECT 558.000 189.700 571.600 190.300 ;
        RECT 558.000 189.600 558.800 189.700 ;
        RECT 570.800 189.600 571.600 189.700 ;
        RECT 44.400 188.300 45.200 188.400 ;
        RECT 63.600 188.300 64.400 188.400 ;
        RECT 71.600 188.300 72.400 188.400 ;
        RECT 44.400 187.700 72.400 188.300 ;
        RECT 44.400 187.600 45.200 187.700 ;
        RECT 63.600 187.600 64.400 187.700 ;
        RECT 71.600 187.600 72.400 187.700 ;
        RECT 97.200 188.300 98.000 188.400 ;
        RECT 98.800 188.300 99.600 188.400 ;
        RECT 103.600 188.300 104.400 188.400 ;
        RECT 97.200 187.700 104.400 188.300 ;
        RECT 97.200 187.600 98.000 187.700 ;
        RECT 98.800 187.600 99.600 187.700 ;
        RECT 103.600 187.600 104.400 187.700 ;
        RECT 108.400 188.300 109.200 188.400 ;
        RECT 113.200 188.300 114.000 188.400 ;
        RECT 108.400 187.700 114.000 188.300 ;
        RECT 108.400 187.600 109.200 187.700 ;
        RECT 113.200 187.600 114.000 187.700 ;
        RECT 193.200 188.300 194.000 188.400 ;
        RECT 204.400 188.300 205.200 188.400 ;
        RECT 193.200 187.700 205.200 188.300 ;
        RECT 193.200 187.600 194.000 187.700 ;
        RECT 204.400 187.600 205.200 187.700 ;
        RECT 246.000 188.300 246.800 188.400 ;
        RECT 258.800 188.300 259.600 188.400 ;
        RECT 246.000 187.700 259.600 188.300 ;
        RECT 246.000 187.600 246.800 187.700 ;
        RECT 258.800 187.600 259.600 187.700 ;
        RECT 308.400 188.300 309.200 188.400 ;
        RECT 332.400 188.300 333.200 188.400 ;
        RECT 308.400 187.700 333.200 188.300 ;
        RECT 308.400 187.600 309.200 187.700 ;
        RECT 332.400 187.600 333.200 187.700 ;
        RECT 342.000 188.300 342.800 188.400 ;
        RECT 354.800 188.300 355.600 188.400 ;
        RECT 342.000 187.700 355.600 188.300 ;
        RECT 342.000 187.600 342.800 187.700 ;
        RECT 354.800 187.600 355.600 187.700 ;
        RECT 388.400 188.300 389.200 188.400 ;
        RECT 406.000 188.300 406.800 188.400 ;
        RECT 388.400 187.700 406.800 188.300 ;
        RECT 388.400 187.600 389.200 187.700 ;
        RECT 406.000 187.600 406.800 187.700 ;
        RECT 452.400 188.300 453.200 188.400 ;
        RECT 463.600 188.300 464.400 188.400 ;
        RECT 476.400 188.300 477.200 188.400 ;
        RECT 452.400 187.700 477.200 188.300 ;
        RECT 452.400 187.600 453.200 187.700 ;
        RECT 463.600 187.600 464.400 187.700 ;
        RECT 476.400 187.600 477.200 187.700 ;
        RECT 481.200 188.300 482.000 188.400 ;
        RECT 492.400 188.300 493.200 188.400 ;
        RECT 481.200 187.700 493.200 188.300 ;
        RECT 481.200 187.600 482.000 187.700 ;
        RECT 492.400 187.600 493.200 187.700 ;
        RECT 494.000 188.300 494.800 188.400 ;
        RECT 497.200 188.300 498.000 188.400 ;
        RECT 508.400 188.300 509.200 188.400 ;
        RECT 494.000 187.700 509.200 188.300 ;
        RECT 494.000 187.600 494.800 187.700 ;
        RECT 497.200 187.600 498.000 187.700 ;
        RECT 508.400 187.600 509.200 187.700 ;
        RECT 532.400 188.300 533.200 188.400 ;
        RECT 542.000 188.300 542.800 188.400 ;
        RECT 532.400 187.700 542.800 188.300 ;
        RECT 532.400 187.600 533.200 187.700 ;
        RECT 542.000 187.600 542.800 187.700 ;
        RECT 548.400 188.300 549.200 188.400 ;
        RECT 564.400 188.300 565.200 188.400 ;
        RECT 548.400 187.700 565.200 188.300 ;
        RECT 548.400 187.600 549.200 187.700 ;
        RECT 564.400 187.600 565.200 187.700 ;
        RECT 18.800 186.300 19.600 186.400 ;
        RECT 25.200 186.300 26.000 186.400 ;
        RECT 18.800 185.700 26.000 186.300 ;
        RECT 18.800 185.600 19.600 185.700 ;
        RECT 25.200 185.600 26.000 185.700 ;
        RECT 38.000 186.300 38.800 186.400 ;
        RECT 46.000 186.300 46.800 186.400 ;
        RECT 50.800 186.300 51.600 186.400 ;
        RECT 60.400 186.300 61.200 186.400 ;
        RECT 73.200 186.300 74.000 186.400 ;
        RECT 74.800 186.300 75.600 186.400 ;
        RECT 78.000 186.300 78.800 186.400 ;
        RECT 38.000 185.700 78.800 186.300 ;
        RECT 38.000 185.600 38.800 185.700 ;
        RECT 46.000 185.600 46.800 185.700 ;
        RECT 50.800 185.600 51.600 185.700 ;
        RECT 60.400 185.600 61.200 185.700 ;
        RECT 73.200 185.600 74.000 185.700 ;
        RECT 74.800 185.600 75.600 185.700 ;
        RECT 78.000 185.600 78.800 185.700 ;
        RECT 92.400 186.300 93.200 186.400 ;
        RECT 108.500 186.300 109.100 187.600 ;
        RECT 92.400 185.700 109.100 186.300 ;
        RECT 172.400 186.300 173.200 186.400 ;
        RECT 198.000 186.300 198.800 186.400 ;
        RECT 212.400 186.300 213.200 186.400 ;
        RECT 172.400 185.700 213.200 186.300 ;
        RECT 92.400 185.600 93.200 185.700 ;
        RECT 172.400 185.600 173.200 185.700 ;
        RECT 198.000 185.600 198.800 185.700 ;
        RECT 212.400 185.600 213.200 185.700 ;
        RECT 242.800 186.300 243.600 186.400 ;
        RECT 257.200 186.300 258.000 186.400 ;
        RECT 268.400 186.300 269.200 186.400 ;
        RECT 242.800 185.700 269.200 186.300 ;
        RECT 242.800 185.600 243.600 185.700 ;
        RECT 257.200 185.600 258.000 185.700 ;
        RECT 268.400 185.600 269.200 185.700 ;
        RECT 292.400 186.300 293.200 186.400 ;
        RECT 310.000 186.300 310.800 186.400 ;
        RECT 292.400 185.700 310.800 186.300 ;
        RECT 292.400 185.600 293.200 185.700 ;
        RECT 310.000 185.600 310.800 185.700 ;
        RECT 313.200 186.300 314.000 186.400 ;
        RECT 322.800 186.300 323.600 186.400 ;
        RECT 313.200 185.700 323.600 186.300 ;
        RECT 313.200 185.600 314.000 185.700 ;
        RECT 322.800 185.600 323.600 185.700 ;
        RECT 332.400 186.300 333.200 186.400 ;
        RECT 343.600 186.300 344.400 186.400 ;
        RECT 332.400 185.700 344.400 186.300 ;
        RECT 332.400 185.600 333.200 185.700 ;
        RECT 343.600 185.600 344.400 185.700 ;
        RECT 378.800 186.300 379.600 186.400 ;
        RECT 391.600 186.300 392.400 186.400 ;
        RECT 378.800 185.700 392.400 186.300 ;
        RECT 378.800 185.600 379.600 185.700 ;
        RECT 391.600 185.600 392.400 185.700 ;
        RECT 460.400 186.300 461.200 186.400 ;
        RECT 465.200 186.300 466.000 186.400 ;
        RECT 460.400 185.700 466.000 186.300 ;
        RECT 460.400 185.600 461.200 185.700 ;
        RECT 465.200 185.600 466.000 185.700 ;
        RECT 476.400 186.300 477.200 186.400 ;
        RECT 494.000 186.300 494.800 186.400 ;
        RECT 513.200 186.300 514.000 186.400 ;
        RECT 521.200 186.300 522.000 186.400 ;
        RECT 524.400 186.300 525.200 186.400 ;
        RECT 476.400 185.700 525.200 186.300 ;
        RECT 476.400 185.600 477.200 185.700 ;
        RECT 494.000 185.600 494.800 185.700 ;
        RECT 513.200 185.600 514.000 185.700 ;
        RECT 521.200 185.600 522.000 185.700 ;
        RECT 524.400 185.600 525.200 185.700 ;
        RECT 526.000 186.300 526.800 186.400 ;
        RECT 532.400 186.300 533.200 186.400 ;
        RECT 535.600 186.300 536.400 186.400 ;
        RECT 526.000 185.700 536.400 186.300 ;
        RECT 526.000 185.600 526.800 185.700 ;
        RECT 532.400 185.600 533.200 185.700 ;
        RECT 535.600 185.600 536.400 185.700 ;
        RECT 2.800 184.300 3.600 184.400 ;
        RECT 18.800 184.300 19.600 184.400 ;
        RECT 2.800 183.700 19.600 184.300 ;
        RECT 2.800 183.600 3.600 183.700 ;
        RECT 18.800 183.600 19.600 183.700 ;
        RECT 26.800 184.300 27.600 184.400 ;
        RECT 38.000 184.300 38.800 184.400 ;
        RECT 26.800 183.700 38.800 184.300 ;
        RECT 26.800 183.600 27.600 183.700 ;
        RECT 38.000 183.600 38.800 183.700 ;
        RECT 145.200 184.300 146.000 184.400 ;
        RECT 150.000 184.300 150.800 184.400 ;
        RECT 145.200 183.700 150.800 184.300 ;
        RECT 145.200 183.600 146.000 183.700 ;
        RECT 150.000 183.600 150.800 183.700 ;
        RECT 183.600 184.300 184.400 184.400 ;
        RECT 210.800 184.300 211.600 184.400 ;
        RECT 183.600 183.700 211.600 184.300 ;
        RECT 183.600 183.600 184.400 183.700 ;
        RECT 210.800 183.600 211.600 183.700 ;
        RECT 273.200 184.300 274.000 184.400 ;
        RECT 314.800 184.300 315.600 184.400 ;
        RECT 335.600 184.300 336.400 184.400 ;
        RECT 273.200 183.700 336.400 184.300 ;
        RECT 273.200 183.600 274.000 183.700 ;
        RECT 314.800 183.600 315.600 183.700 ;
        RECT 335.600 183.600 336.400 183.700 ;
        RECT 351.600 184.300 352.400 184.400 ;
        RECT 420.400 184.300 421.200 184.400 ;
        RECT 351.600 183.700 421.200 184.300 ;
        RECT 351.600 183.600 352.400 183.700 ;
        RECT 420.400 183.600 421.200 183.700 ;
        RECT 474.800 184.300 475.600 184.400 ;
        RECT 484.400 184.300 485.200 184.400 ;
        RECT 489.200 184.300 490.000 184.400 ;
        RECT 474.800 183.700 490.000 184.300 ;
        RECT 474.800 183.600 475.600 183.700 ;
        RECT 484.400 183.600 485.200 183.700 ;
        RECT 489.200 183.600 490.000 183.700 ;
        RECT 492.400 184.300 493.200 184.400 ;
        RECT 516.400 184.300 517.200 184.400 ;
        RECT 492.400 183.700 517.200 184.300 ;
        RECT 492.400 183.600 493.200 183.700 ;
        RECT 516.400 183.600 517.200 183.700 ;
        RECT 559.600 184.300 560.400 184.400 ;
        RECT 566.000 184.300 566.800 184.400 ;
        RECT 559.600 183.700 566.800 184.300 ;
        RECT 559.600 183.600 560.400 183.700 ;
        RECT 566.000 183.600 566.800 183.700 ;
        RECT 153.200 182.300 154.000 182.400 ;
        RECT 172.400 182.300 173.200 182.400 ;
        RECT 185.200 182.300 186.000 182.400 ;
        RECT 153.200 181.700 186.000 182.300 ;
        RECT 153.200 181.600 154.000 181.700 ;
        RECT 172.400 181.600 173.200 181.700 ;
        RECT 185.200 181.600 186.000 181.700 ;
        RECT 391.600 182.300 392.400 182.400 ;
        RECT 399.600 182.300 400.400 182.400 ;
        RECT 391.600 181.700 400.400 182.300 ;
        RECT 391.600 181.600 392.400 181.700 ;
        RECT 399.600 181.600 400.400 181.700 ;
        RECT 425.200 182.300 426.000 182.400 ;
        RECT 458.800 182.300 459.600 182.400 ;
        RECT 425.200 181.700 459.600 182.300 ;
        RECT 425.200 181.600 426.000 181.700 ;
        RECT 458.800 181.600 459.600 181.700 ;
        RECT 486.000 182.300 486.800 182.400 ;
        RECT 498.800 182.300 499.600 182.400 ;
        RECT 486.000 181.700 499.600 182.300 ;
        RECT 486.000 181.600 486.800 181.700 ;
        RECT 498.800 181.600 499.600 181.700 ;
        RECT 508.400 182.300 509.200 182.400 ;
        RECT 534.000 182.300 534.800 182.400 ;
        RECT 508.400 181.700 534.800 182.300 ;
        RECT 508.400 181.600 509.200 181.700 ;
        RECT 534.000 181.600 534.800 181.700 ;
        RECT 566.000 182.300 566.800 182.400 ;
        RECT 583.600 182.300 584.400 182.400 ;
        RECT 566.000 181.700 584.400 182.300 ;
        RECT 566.000 181.600 566.800 181.700 ;
        RECT 583.600 181.600 584.400 181.700 ;
        RECT 326.000 180.300 326.800 180.400 ;
        RECT 343.600 180.300 344.400 180.400 ;
        RECT 361.200 180.300 362.000 180.400 ;
        RECT 326.000 179.700 362.000 180.300 ;
        RECT 326.000 179.600 326.800 179.700 ;
        RECT 343.600 179.600 344.400 179.700 ;
        RECT 361.200 179.600 362.000 179.700 ;
        RECT 374.000 180.300 374.800 180.400 ;
        RECT 414.000 180.300 414.800 180.400 ;
        RECT 374.000 179.700 414.800 180.300 ;
        RECT 374.000 179.600 374.800 179.700 ;
        RECT 414.000 179.600 414.800 179.700 ;
        RECT 457.200 180.300 458.000 180.400 ;
        RECT 476.400 180.300 477.200 180.400 ;
        RECT 457.200 179.700 477.200 180.300 ;
        RECT 457.200 179.600 458.000 179.700 ;
        RECT 476.400 179.600 477.200 179.700 ;
        RECT 503.600 180.300 504.400 180.400 ;
        RECT 532.400 180.300 533.200 180.400 ;
        RECT 540.400 180.300 541.200 180.400 ;
        RECT 503.600 179.700 541.200 180.300 ;
        RECT 503.600 179.600 504.400 179.700 ;
        RECT 532.400 179.600 533.200 179.700 ;
        RECT 540.400 179.600 541.200 179.700 ;
        RECT 23.600 178.300 24.400 178.400 ;
        RECT 39.600 178.300 40.400 178.400 ;
        RECT 23.600 177.700 40.400 178.300 ;
        RECT 23.600 177.600 24.400 177.700 ;
        RECT 39.600 177.600 40.400 177.700 ;
        RECT 92.400 178.300 93.200 178.400 ;
        RECT 102.000 178.300 102.800 178.400 ;
        RECT 92.400 177.700 102.800 178.300 ;
        RECT 92.400 177.600 93.200 177.700 ;
        RECT 102.000 177.600 102.800 177.700 ;
        RECT 186.800 178.300 187.600 178.400 ;
        RECT 193.200 178.300 194.000 178.400 ;
        RECT 204.400 178.300 205.200 178.400 ;
        RECT 186.800 177.700 205.200 178.300 ;
        RECT 186.800 177.600 187.600 177.700 ;
        RECT 193.200 177.600 194.000 177.700 ;
        RECT 204.400 177.600 205.200 177.700 ;
        RECT 308.400 178.300 309.200 178.400 ;
        RECT 313.200 178.300 314.000 178.400 ;
        RECT 374.000 178.300 374.800 178.400 ;
        RECT 390.000 178.300 390.800 178.400 ;
        RECT 401.200 178.300 402.000 178.400 ;
        RECT 404.400 178.300 405.200 178.400 ;
        RECT 308.400 177.700 341.100 178.300 ;
        RECT 308.400 177.600 309.200 177.700 ;
        RECT 313.200 177.600 314.000 177.700 ;
        RECT 340.500 176.400 341.100 177.700 ;
        RECT 374.000 177.700 405.200 178.300 ;
        RECT 374.000 177.600 374.800 177.700 ;
        RECT 390.000 177.600 390.800 177.700 ;
        RECT 401.200 177.600 402.000 177.700 ;
        RECT 404.400 177.600 405.200 177.700 ;
        RECT 500.400 178.300 501.200 178.400 ;
        RECT 506.800 178.300 507.600 178.400 ;
        RECT 500.400 177.700 507.600 178.300 ;
        RECT 500.400 177.600 501.200 177.700 ;
        RECT 506.800 177.600 507.600 177.700 ;
        RECT 530.800 178.300 531.600 178.400 ;
        RECT 556.400 178.300 557.200 178.400 ;
        RECT 530.800 177.700 557.200 178.300 ;
        RECT 530.800 177.600 531.600 177.700 ;
        RECT 556.400 177.600 557.200 177.700 ;
        RECT 12.400 176.300 13.200 176.400 ;
        RECT 14.000 176.300 14.800 176.400 ;
        RECT 12.400 175.700 14.800 176.300 ;
        RECT 12.400 175.600 13.200 175.700 ;
        RECT 14.000 175.600 14.800 175.700 ;
        RECT 25.200 176.300 26.000 176.400 ;
        RECT 30.000 176.300 30.800 176.400 ;
        RECT 25.200 175.700 30.800 176.300 ;
        RECT 25.200 175.600 26.000 175.700 ;
        RECT 30.000 175.600 30.800 175.700 ;
        RECT 52.400 176.300 53.200 176.400 ;
        RECT 55.600 176.300 56.400 176.400 ;
        RECT 52.400 175.700 56.400 176.300 ;
        RECT 52.400 175.600 53.200 175.700 ;
        RECT 55.600 175.600 56.400 175.700 ;
        RECT 60.400 176.300 61.200 176.400 ;
        RECT 82.800 176.300 83.600 176.400 ;
        RECT 60.400 175.700 83.600 176.300 ;
        RECT 60.400 175.600 61.200 175.700 ;
        RECT 82.800 175.600 83.600 175.700 ;
        RECT 185.200 176.300 186.000 176.400 ;
        RECT 207.600 176.300 208.400 176.400 ;
        RECT 185.200 175.700 208.400 176.300 ;
        RECT 185.200 175.600 186.000 175.700 ;
        RECT 207.600 175.600 208.400 175.700 ;
        RECT 210.800 176.300 211.600 176.400 ;
        RECT 217.200 176.300 218.000 176.400 ;
        RECT 210.800 175.700 218.000 176.300 ;
        RECT 210.800 175.600 211.600 175.700 ;
        RECT 217.200 175.600 218.000 175.700 ;
        RECT 321.200 176.300 322.000 176.400 ;
        RECT 332.400 176.300 333.200 176.400 ;
        RECT 321.200 175.700 333.200 176.300 ;
        RECT 321.200 175.600 322.000 175.700 ;
        RECT 332.400 175.600 333.200 175.700 ;
        RECT 340.400 176.300 341.200 176.400 ;
        RECT 345.200 176.300 346.000 176.400 ;
        RECT 340.400 175.700 346.000 176.300 ;
        RECT 340.400 175.600 341.200 175.700 ;
        RECT 345.200 175.600 346.000 175.700 ;
        RECT 362.800 176.300 363.600 176.400 ;
        RECT 396.400 176.300 397.200 176.400 ;
        RECT 362.800 175.700 397.200 176.300 ;
        RECT 362.800 175.600 363.600 175.700 ;
        RECT 396.400 175.600 397.200 175.700 ;
        RECT 502.000 176.300 502.800 176.400 ;
        RECT 510.000 176.300 510.800 176.400 ;
        RECT 502.000 175.700 510.800 176.300 ;
        RECT 502.000 175.600 502.800 175.700 ;
        RECT 510.000 175.600 510.800 175.700 ;
        RECT 511.600 176.300 512.400 176.400 ;
        RECT 514.800 176.300 515.600 176.400 ;
        RECT 511.600 175.700 515.600 176.300 ;
        RECT 511.600 175.600 512.400 175.700 ;
        RECT 514.800 175.600 515.600 175.700 ;
        RECT 518.000 176.300 518.800 176.400 ;
        RECT 522.800 176.300 523.600 176.400 ;
        RECT 518.000 175.700 523.600 176.300 ;
        RECT 518.000 175.600 518.800 175.700 ;
        RECT 522.800 175.600 523.600 175.700 ;
        RECT 524.400 176.300 525.200 176.400 ;
        RECT 529.200 176.300 530.000 176.400 ;
        RECT 524.400 175.700 530.000 176.300 ;
        RECT 524.400 175.600 525.200 175.700 ;
        RECT 529.200 175.600 530.000 175.700 ;
        RECT 534.000 176.300 534.800 176.400 ;
        RECT 543.600 176.300 544.400 176.400 ;
        RECT 534.000 175.700 544.400 176.300 ;
        RECT 534.000 175.600 534.800 175.700 ;
        RECT 543.600 175.600 544.400 175.700 ;
        RECT 47.600 173.600 48.400 174.400 ;
        RECT 54.000 174.300 54.800 174.400 ;
        RECT 70.000 174.300 70.800 174.400 ;
        RECT 54.000 173.700 70.800 174.300 ;
        RECT 54.000 173.600 54.800 173.700 ;
        RECT 70.000 173.600 70.800 173.700 ;
        RECT 74.800 174.300 75.600 174.400 ;
        RECT 94.000 174.300 94.800 174.400 ;
        RECT 74.800 173.700 94.800 174.300 ;
        RECT 74.800 173.600 75.600 173.700 ;
        RECT 94.000 173.600 94.800 173.700 ;
        RECT 111.600 174.300 112.400 174.400 ;
        RECT 124.400 174.300 125.200 174.400 ;
        RECT 111.600 173.700 125.200 174.300 ;
        RECT 111.600 173.600 112.400 173.700 ;
        RECT 124.400 173.600 125.200 173.700 ;
        RECT 145.200 174.300 146.000 174.400 ;
        RECT 154.800 174.300 155.600 174.400 ;
        RECT 145.200 173.700 155.600 174.300 ;
        RECT 145.200 173.600 146.000 173.700 ;
        RECT 154.800 173.600 155.600 173.700 ;
        RECT 183.600 174.300 184.400 174.400 ;
        RECT 190.000 174.300 190.800 174.400 ;
        RECT 199.600 174.300 200.400 174.400 ;
        RECT 201.200 174.300 202.000 174.400 ;
        RECT 222.000 174.300 222.800 174.400 ;
        RECT 183.600 173.700 202.000 174.300 ;
        RECT 183.600 173.600 184.400 173.700 ;
        RECT 190.000 173.600 190.800 173.700 ;
        RECT 199.600 173.600 200.400 173.700 ;
        RECT 201.200 173.600 202.000 173.700 ;
        RECT 212.500 173.700 222.800 174.300 ;
        RECT 33.200 172.300 34.000 172.400 ;
        RECT 38.000 172.300 38.800 172.400 ;
        RECT 33.200 171.700 38.800 172.300 ;
        RECT 33.200 171.600 34.000 171.700 ;
        RECT 38.000 171.600 38.800 171.700 ;
        RECT 41.200 172.300 42.000 172.400 ;
        RECT 47.700 172.300 48.300 173.600 ;
        RECT 212.500 172.400 213.100 173.700 ;
        RECT 222.000 173.600 222.800 173.700 ;
        RECT 265.200 174.300 266.000 174.400 ;
        RECT 268.400 174.300 269.200 174.400 ;
        RECT 292.400 174.300 293.200 174.400 ;
        RECT 265.200 173.700 293.200 174.300 ;
        RECT 265.200 173.600 266.000 173.700 ;
        RECT 268.400 173.600 269.200 173.700 ;
        RECT 292.400 173.600 293.200 173.700 ;
        RECT 324.400 174.300 325.200 174.400 ;
        RECT 348.400 174.300 349.200 174.400 ;
        RECT 324.400 173.700 349.200 174.300 ;
        RECT 324.400 173.600 325.200 173.700 ;
        RECT 348.400 173.600 349.200 173.700 ;
        RECT 356.400 174.300 357.200 174.400 ;
        RECT 358.000 174.300 358.800 174.400 ;
        RECT 356.400 173.700 358.800 174.300 ;
        RECT 356.400 173.600 357.200 173.700 ;
        RECT 358.000 173.600 358.800 173.700 ;
        RECT 361.200 174.300 362.000 174.400 ;
        RECT 366.000 174.300 366.800 174.400 ;
        RECT 361.200 173.700 366.800 174.300 ;
        RECT 361.200 173.600 362.000 173.700 ;
        RECT 366.000 173.600 366.800 173.700 ;
        RECT 372.400 174.300 373.200 174.400 ;
        RECT 377.200 174.300 378.000 174.400 ;
        RECT 372.400 173.700 378.000 174.300 ;
        RECT 372.400 173.600 373.200 173.700 ;
        RECT 377.200 173.600 378.000 173.700 ;
        RECT 418.800 174.300 419.600 174.400 ;
        RECT 446.000 174.300 446.800 174.400 ;
        RECT 418.800 173.700 446.800 174.300 ;
        RECT 418.800 173.600 419.600 173.700 ;
        RECT 446.000 173.600 446.800 173.700 ;
        RECT 490.800 174.300 491.600 174.400 ;
        RECT 530.800 174.300 531.600 174.400 ;
        RECT 490.800 173.700 531.600 174.300 ;
        RECT 490.800 173.600 491.600 173.700 ;
        RECT 530.800 173.600 531.600 173.700 ;
        RECT 538.800 174.300 539.600 174.400 ;
        RECT 543.600 174.300 544.400 174.400 ;
        RECT 538.800 173.700 544.400 174.300 ;
        RECT 538.800 173.600 539.600 173.700 ;
        RECT 543.600 173.600 544.400 173.700 ;
        RECT 545.200 173.600 546.000 174.400 ;
        RECT 41.200 171.700 48.300 172.300 ;
        RECT 57.200 172.300 58.000 172.400 ;
        RECT 60.400 172.300 61.200 172.400 ;
        RECT 57.200 171.700 61.200 172.300 ;
        RECT 41.200 171.600 42.000 171.700 ;
        RECT 57.200 171.600 58.000 171.700 ;
        RECT 60.400 171.600 61.200 171.700 ;
        RECT 65.200 172.300 66.000 172.400 ;
        RECT 70.000 172.300 70.800 172.400 ;
        RECT 65.200 171.700 70.800 172.300 ;
        RECT 65.200 171.600 66.000 171.700 ;
        RECT 70.000 171.600 70.800 171.700 ;
        RECT 87.600 172.300 88.400 172.400 ;
        RECT 110.000 172.300 110.800 172.400 ;
        RECT 87.600 171.700 110.800 172.300 ;
        RECT 87.600 171.600 88.400 171.700 ;
        RECT 110.000 171.600 110.800 171.700 ;
        RECT 132.400 172.300 133.200 172.400 ;
        RECT 158.000 172.300 158.800 172.400 ;
        RECT 132.400 171.700 158.800 172.300 ;
        RECT 132.400 171.600 133.200 171.700 ;
        RECT 158.000 171.600 158.800 171.700 ;
        RECT 182.000 172.300 182.800 172.400 ;
        RECT 186.800 172.300 187.600 172.400 ;
        RECT 182.000 171.700 187.600 172.300 ;
        RECT 182.000 171.600 182.800 171.700 ;
        RECT 186.800 171.600 187.600 171.700 ;
        RECT 202.800 172.300 203.600 172.400 ;
        RECT 212.400 172.300 213.200 172.400 ;
        RECT 202.800 171.700 213.200 172.300 ;
        RECT 202.800 171.600 203.600 171.700 ;
        RECT 212.400 171.600 213.200 171.700 ;
        RECT 215.600 172.300 216.400 172.400 ;
        RECT 220.400 172.300 221.200 172.400 ;
        RECT 226.800 172.300 227.600 172.400 ;
        RECT 238.000 172.300 238.800 172.400 ;
        RECT 215.600 171.700 238.800 172.300 ;
        RECT 215.600 171.600 216.400 171.700 ;
        RECT 220.400 171.600 221.200 171.700 ;
        RECT 226.800 171.600 227.600 171.700 ;
        RECT 238.000 171.600 238.800 171.700 ;
        RECT 319.600 172.300 320.400 172.400 ;
        RECT 337.200 172.300 338.000 172.400 ;
        RECT 319.600 171.700 338.000 172.300 ;
        RECT 319.600 171.600 320.400 171.700 ;
        RECT 337.200 171.600 338.000 171.700 ;
        RECT 353.200 172.300 354.000 172.400 ;
        RECT 364.400 172.300 365.200 172.400 ;
        RECT 382.000 172.300 382.800 172.400 ;
        RECT 386.800 172.300 387.600 172.400 ;
        RECT 353.200 171.700 387.600 172.300 ;
        RECT 353.200 171.600 354.000 171.700 ;
        RECT 364.400 171.600 365.200 171.700 ;
        RECT 382.000 171.600 382.800 171.700 ;
        RECT 386.800 171.600 387.600 171.700 ;
        RECT 390.000 172.300 390.800 172.400 ;
        RECT 401.200 172.300 402.000 172.400 ;
        RECT 390.000 171.700 402.000 172.300 ;
        RECT 390.000 171.600 390.800 171.700 ;
        RECT 401.200 171.600 402.000 171.700 ;
        RECT 406.000 172.300 406.800 172.400 ;
        RECT 409.200 172.300 410.000 172.400 ;
        RECT 406.000 171.700 410.000 172.300 ;
        RECT 406.000 171.600 406.800 171.700 ;
        RECT 409.200 171.600 410.000 171.700 ;
        RECT 410.800 172.300 411.600 172.400 ;
        RECT 420.400 172.300 421.200 172.400 ;
        RECT 410.800 171.700 421.200 172.300 ;
        RECT 410.800 171.600 411.600 171.700 ;
        RECT 420.400 171.600 421.200 171.700 ;
        RECT 452.400 172.300 453.200 172.400 ;
        RECT 462.000 172.300 462.800 172.400 ;
        RECT 452.400 171.700 462.800 172.300 ;
        RECT 452.400 171.600 453.200 171.700 ;
        RECT 462.000 171.600 462.800 171.700 ;
        RECT 503.600 172.300 504.400 172.400 ;
        RECT 508.400 172.300 509.200 172.400 ;
        RECT 518.000 172.300 518.800 172.400 ;
        RECT 503.600 171.700 518.800 172.300 ;
        RECT 503.600 171.600 504.400 171.700 ;
        RECT 508.400 171.600 509.200 171.700 ;
        RECT 518.000 171.600 518.800 171.700 ;
        RECT 530.800 172.300 531.600 172.400 ;
        RECT 545.300 172.300 545.900 173.600 ;
        RECT 530.800 171.700 545.900 172.300 ;
        RECT 530.800 171.600 531.600 171.700 ;
        RECT 58.800 170.300 59.600 170.400 ;
        RECT 81.200 170.300 82.000 170.400 ;
        RECT 119.600 170.300 120.400 170.400 ;
        RECT 127.600 170.300 128.400 170.400 ;
        RECT 58.800 169.700 128.400 170.300 ;
        RECT 58.800 169.600 59.600 169.700 ;
        RECT 81.200 169.600 82.000 169.700 ;
        RECT 119.600 169.600 120.400 169.700 ;
        RECT 127.600 169.600 128.400 169.700 ;
        RECT 198.000 170.300 198.800 170.400 ;
        RECT 215.600 170.300 216.400 170.400 ;
        RECT 223.600 170.300 224.400 170.400 ;
        RECT 198.000 169.700 224.400 170.300 ;
        RECT 198.000 169.600 198.800 169.700 ;
        RECT 215.600 169.600 216.400 169.700 ;
        RECT 223.600 169.600 224.400 169.700 ;
        RECT 230.000 170.300 230.800 170.400 ;
        RECT 271.600 170.300 272.400 170.400 ;
        RECT 230.000 169.700 272.400 170.300 ;
        RECT 230.000 169.600 230.800 169.700 ;
        RECT 271.600 169.600 272.400 169.700 ;
        RECT 298.800 170.300 299.600 170.400 ;
        RECT 306.800 170.300 307.600 170.400 ;
        RECT 318.000 170.300 318.800 170.400 ;
        RECT 298.800 169.700 318.800 170.300 ;
        RECT 298.800 169.600 299.600 169.700 ;
        RECT 306.800 169.600 307.600 169.700 ;
        RECT 318.000 169.600 318.800 169.700 ;
        RECT 321.200 170.300 322.000 170.400 ;
        RECT 326.000 170.300 326.800 170.400 ;
        RECT 321.200 169.700 326.800 170.300 ;
        RECT 321.200 169.600 322.000 169.700 ;
        RECT 326.000 169.600 326.800 169.700 ;
        RECT 335.600 170.300 336.400 170.400 ;
        RECT 342.000 170.300 342.800 170.400 ;
        RECT 335.600 169.700 342.800 170.300 ;
        RECT 335.600 169.600 336.400 169.700 ;
        RECT 342.000 169.600 342.800 169.700 ;
        RECT 348.400 170.300 349.200 170.400 ;
        RECT 351.600 170.300 352.400 170.400 ;
        RECT 348.400 169.700 352.400 170.300 ;
        RECT 348.400 169.600 349.200 169.700 ;
        RECT 351.600 169.600 352.400 169.700 ;
        RECT 361.200 170.300 362.000 170.400 ;
        RECT 374.000 170.300 374.800 170.400 ;
        RECT 361.200 169.700 374.800 170.300 ;
        RECT 361.200 169.600 362.000 169.700 ;
        RECT 374.000 169.600 374.800 169.700 ;
        RECT 380.400 170.300 381.200 170.400 ;
        RECT 388.400 170.300 389.200 170.400 ;
        RECT 393.200 170.300 394.000 170.400 ;
        RECT 380.400 169.700 394.000 170.300 ;
        RECT 380.400 169.600 381.200 169.700 ;
        RECT 388.400 169.600 389.200 169.700 ;
        RECT 393.200 169.600 394.000 169.700 ;
        RECT 396.400 170.300 397.200 170.400 ;
        RECT 399.600 170.300 400.400 170.400 ;
        RECT 396.400 169.700 400.400 170.300 ;
        RECT 396.400 169.600 397.200 169.700 ;
        RECT 399.600 169.600 400.400 169.700 ;
        RECT 431.600 169.600 432.400 170.400 ;
        RECT 498.800 170.300 499.600 170.400 ;
        RECT 505.200 170.300 506.000 170.400 ;
        RECT 508.400 170.300 509.200 170.400 ;
        RECT 498.800 169.700 509.200 170.300 ;
        RECT 498.800 169.600 499.600 169.700 ;
        RECT 505.200 169.600 506.000 169.700 ;
        RECT 508.400 169.600 509.200 169.700 ;
        RECT 511.600 170.300 512.400 170.400 ;
        RECT 519.600 170.300 520.400 170.400 ;
        RECT 511.600 169.700 520.400 170.300 ;
        RECT 511.600 169.600 512.400 169.700 ;
        RECT 519.600 169.600 520.400 169.700 ;
        RECT 527.600 170.300 528.400 170.400 ;
        RECT 530.800 170.300 531.600 170.400 ;
        RECT 546.800 170.300 547.600 170.400 ;
        RECT 527.600 169.700 547.600 170.300 ;
        RECT 527.600 169.600 528.400 169.700 ;
        RECT 530.800 169.600 531.600 169.700 ;
        RECT 546.800 169.600 547.600 169.700 ;
        RECT 49.200 168.300 50.000 168.400 ;
        RECT 78.000 168.300 78.800 168.400 ;
        RECT 49.200 167.700 78.800 168.300 ;
        RECT 49.200 167.600 50.000 167.700 ;
        RECT 78.000 167.600 78.800 167.700 ;
        RECT 220.400 168.300 221.200 168.400 ;
        RECT 231.600 168.300 232.400 168.400 ;
        RECT 220.400 167.700 232.400 168.300 ;
        RECT 220.400 167.600 221.200 167.700 ;
        RECT 231.600 167.600 232.400 167.700 ;
        RECT 284.400 168.300 285.200 168.400 ;
        RECT 330.800 168.300 331.600 168.400 ;
        RECT 346.800 168.300 347.600 168.400 ;
        RECT 284.400 167.700 347.600 168.300 ;
        RECT 284.400 167.600 285.200 167.700 ;
        RECT 330.800 167.600 331.600 167.700 ;
        RECT 346.800 167.600 347.600 167.700 ;
        RECT 369.200 168.300 370.000 168.400 ;
        RECT 377.200 168.300 378.000 168.400 ;
        RECT 385.200 168.300 386.000 168.400 ;
        RECT 391.600 168.300 392.400 168.400 ;
        RECT 406.000 168.300 406.800 168.400 ;
        RECT 369.200 167.700 406.800 168.300 ;
        RECT 369.200 167.600 370.000 167.700 ;
        RECT 377.200 167.600 378.000 167.700 ;
        RECT 385.200 167.600 386.000 167.700 ;
        RECT 391.600 167.600 392.400 167.700 ;
        RECT 406.000 167.600 406.800 167.700 ;
        RECT 510.000 168.300 510.800 168.400 ;
        RECT 513.200 168.300 514.000 168.400 ;
        RECT 510.000 167.700 514.000 168.300 ;
        RECT 510.000 167.600 510.800 167.700 ;
        RECT 513.200 167.600 514.000 167.700 ;
        RECT 516.400 168.300 517.200 168.400 ;
        RECT 529.200 168.300 530.000 168.400 ;
        RECT 516.400 167.700 530.000 168.300 ;
        RECT 516.400 167.600 517.200 167.700 ;
        RECT 529.200 167.600 530.000 167.700 ;
        RECT 537.200 168.300 538.000 168.400 ;
        RECT 550.000 168.300 550.800 168.400 ;
        RECT 537.200 167.700 550.800 168.300 ;
        RECT 537.200 167.600 538.000 167.700 ;
        RECT 550.000 167.600 550.800 167.700 ;
        RECT 44.400 166.300 45.200 166.400 ;
        RECT 138.800 166.300 139.600 166.400 ;
        RECT 44.400 165.700 139.600 166.300 ;
        RECT 44.400 165.600 45.200 165.700 ;
        RECT 138.800 165.600 139.600 165.700 ;
        RECT 178.800 166.300 179.600 166.400 ;
        RECT 295.600 166.300 296.400 166.400 ;
        RECT 178.800 165.700 296.400 166.300 ;
        RECT 178.800 165.600 179.600 165.700 ;
        RECT 295.600 165.600 296.400 165.700 ;
        RECT 356.400 166.300 357.200 166.400 ;
        RECT 375.600 166.300 376.400 166.400 ;
        RECT 356.400 165.700 376.400 166.300 ;
        RECT 356.400 165.600 357.200 165.700 ;
        RECT 375.600 165.600 376.400 165.700 ;
        RECT 527.600 166.300 528.400 166.400 ;
        RECT 537.200 166.300 538.000 166.400 ;
        RECT 527.600 165.700 538.000 166.300 ;
        RECT 527.600 165.600 528.400 165.700 ;
        RECT 537.200 165.600 538.000 165.700 ;
        RECT 538.800 166.300 539.600 166.400 ;
        RECT 545.200 166.300 546.000 166.400 ;
        RECT 538.800 165.700 546.000 166.300 ;
        RECT 538.800 165.600 539.600 165.700 ;
        RECT 545.200 165.600 546.000 165.700 ;
        RECT 100.400 164.300 101.200 164.400 ;
        RECT 110.000 164.300 110.800 164.400 ;
        RECT 100.400 163.700 110.800 164.300 ;
        RECT 100.400 163.600 101.200 163.700 ;
        RECT 110.000 163.600 110.800 163.700 ;
        RECT 247.600 164.300 248.400 164.400 ;
        RECT 250.800 164.300 251.600 164.400 ;
        RECT 247.600 163.700 251.600 164.300 ;
        RECT 247.600 163.600 248.400 163.700 ;
        RECT 250.800 163.600 251.600 163.700 ;
        RECT 514.800 164.300 515.600 164.400 ;
        RECT 535.600 164.300 536.400 164.400 ;
        RECT 514.800 163.700 536.400 164.300 ;
        RECT 514.800 163.600 515.600 163.700 ;
        RECT 535.600 163.600 536.400 163.700 ;
        RECT 546.800 164.300 547.600 164.400 ;
        RECT 551.600 164.300 552.400 164.400 ;
        RECT 546.800 163.700 552.400 164.300 ;
        RECT 546.800 163.600 547.600 163.700 ;
        RECT 551.600 163.600 552.400 163.700 ;
        RECT 553.200 164.300 554.000 164.400 ;
        RECT 570.800 164.300 571.600 164.400 ;
        RECT 553.200 163.700 571.600 164.300 ;
        RECT 553.200 163.600 554.000 163.700 ;
        RECT 570.800 163.600 571.600 163.700 ;
        RECT 103.600 162.300 104.400 162.400 ;
        RECT 111.600 162.300 112.400 162.400 ;
        RECT 103.600 161.700 112.400 162.300 ;
        RECT 103.600 161.600 104.400 161.700 ;
        RECT 111.600 161.600 112.400 161.700 ;
        RECT 170.800 162.300 171.600 162.400 ;
        RECT 268.400 162.300 269.200 162.400 ;
        RECT 170.800 161.700 269.200 162.300 ;
        RECT 170.800 161.600 171.600 161.700 ;
        RECT 268.400 161.600 269.200 161.700 ;
        RECT 524.400 162.300 525.200 162.400 ;
        RECT 537.200 162.300 538.000 162.400 ;
        RECT 524.400 161.700 538.000 162.300 ;
        RECT 524.400 161.600 525.200 161.700 ;
        RECT 537.200 161.600 538.000 161.700 ;
        RECT 540.400 162.300 541.200 162.400 ;
        RECT 553.200 162.300 554.000 162.400 ;
        RECT 540.400 161.700 554.000 162.300 ;
        RECT 540.400 161.600 541.200 161.700 ;
        RECT 553.200 161.600 554.000 161.700 ;
        RECT 398.000 160.300 398.800 160.400 ;
        RECT 402.800 160.300 403.600 160.400 ;
        RECT 398.000 159.700 403.600 160.300 ;
        RECT 398.000 159.600 398.800 159.700 ;
        RECT 402.800 159.600 403.600 159.700 ;
        RECT 513.200 160.300 514.000 160.400 ;
        RECT 551.600 160.300 552.400 160.400 ;
        RECT 513.200 159.700 552.400 160.300 ;
        RECT 513.200 159.600 514.000 159.700 ;
        RECT 551.600 159.600 552.400 159.700 ;
        RECT 18.800 158.300 19.600 158.400 ;
        RECT 33.200 158.300 34.000 158.400 ;
        RECT 18.800 157.700 34.000 158.300 ;
        RECT 18.800 157.600 19.600 157.700 ;
        RECT 33.200 157.600 34.000 157.700 ;
        RECT 122.800 158.300 123.600 158.400 ;
        RECT 244.400 158.300 245.200 158.400 ;
        RECT 122.800 157.700 245.200 158.300 ;
        RECT 122.800 157.600 123.600 157.700 ;
        RECT 244.400 157.600 245.200 157.700 ;
        RECT 375.600 158.300 376.400 158.400 ;
        RECT 398.000 158.300 398.800 158.400 ;
        RECT 417.200 158.300 418.000 158.400 ;
        RECT 375.600 157.700 418.000 158.300 ;
        RECT 375.600 157.600 376.400 157.700 ;
        RECT 398.000 157.600 398.800 157.700 ;
        RECT 417.200 157.600 418.000 157.700 ;
        RECT 447.600 158.300 448.400 158.400 ;
        RECT 455.600 158.300 456.400 158.400 ;
        RECT 447.600 157.700 456.400 158.300 ;
        RECT 447.600 157.600 448.400 157.700 ;
        RECT 455.600 157.600 456.400 157.700 ;
        RECT 486.000 158.300 486.800 158.400 ;
        RECT 490.800 158.300 491.600 158.400 ;
        RECT 486.000 157.700 491.600 158.300 ;
        RECT 486.000 157.600 486.800 157.700 ;
        RECT 490.800 157.600 491.600 157.700 ;
        RECT 530.800 158.300 531.600 158.400 ;
        RECT 534.000 158.300 534.800 158.400 ;
        RECT 530.800 157.700 534.800 158.300 ;
        RECT 530.800 157.600 531.600 157.700 ;
        RECT 534.000 157.600 534.800 157.700 ;
        RECT 23.600 156.300 24.400 156.400 ;
        RECT 26.800 156.300 27.600 156.400 ;
        RECT 23.600 155.700 27.600 156.300 ;
        RECT 23.600 155.600 24.400 155.700 ;
        RECT 26.800 155.600 27.600 155.700 ;
        RECT 108.400 156.300 109.200 156.400 ;
        RECT 188.400 156.300 189.200 156.400 ;
        RECT 108.400 155.700 189.200 156.300 ;
        RECT 108.400 155.600 109.200 155.700 ;
        RECT 188.400 155.600 189.200 155.700 ;
        RECT 324.400 156.300 325.200 156.400 ;
        RECT 370.800 156.300 371.600 156.400 ;
        RECT 375.600 156.300 376.400 156.400 ;
        RECT 380.400 156.300 381.200 156.400 ;
        RECT 324.400 155.700 381.200 156.300 ;
        RECT 324.400 155.600 325.200 155.700 ;
        RECT 370.800 155.600 371.600 155.700 ;
        RECT 375.600 155.600 376.400 155.700 ;
        RECT 380.400 155.600 381.200 155.700 ;
        RECT 420.400 156.300 421.200 156.400 ;
        RECT 463.600 156.300 464.400 156.400 ;
        RECT 420.400 155.700 464.400 156.300 ;
        RECT 420.400 155.600 421.200 155.700 ;
        RECT 463.600 155.600 464.400 155.700 ;
        RECT 505.200 156.300 506.000 156.400 ;
        RECT 519.600 156.300 520.400 156.400 ;
        RECT 526.000 156.300 526.800 156.400 ;
        RECT 505.200 155.700 526.800 156.300 ;
        RECT 505.200 155.600 506.000 155.700 ;
        RECT 519.600 155.600 520.400 155.700 ;
        RECT 526.000 155.600 526.800 155.700 ;
        RECT 12.400 154.300 13.200 154.400 ;
        RECT 22.000 154.300 22.800 154.400 ;
        RECT 12.400 153.700 22.800 154.300 ;
        RECT 12.400 153.600 13.200 153.700 ;
        RECT 22.000 153.600 22.800 153.700 ;
        RECT 49.200 154.300 50.000 154.400 ;
        RECT 63.600 154.300 64.400 154.400 ;
        RECT 49.200 153.700 64.400 154.300 ;
        RECT 49.200 153.600 50.000 153.700 ;
        RECT 63.600 153.600 64.400 153.700 ;
        RECT 103.600 154.300 104.400 154.400 ;
        RECT 106.800 154.300 107.600 154.400 ;
        RECT 103.600 153.700 107.600 154.300 ;
        RECT 103.600 153.600 104.400 153.700 ;
        RECT 106.800 153.600 107.600 153.700 ;
        RECT 110.000 154.300 110.800 154.400 ;
        RECT 142.000 154.300 142.800 154.400 ;
        RECT 110.000 153.700 142.800 154.300 ;
        RECT 110.000 153.600 110.800 153.700 ;
        RECT 142.000 153.600 142.800 153.700 ;
        RECT 239.600 154.300 240.400 154.400 ;
        RECT 298.800 154.300 299.600 154.400 ;
        RECT 239.600 153.700 299.600 154.300 ;
        RECT 239.600 153.600 240.400 153.700 ;
        RECT 298.800 153.600 299.600 153.700 ;
        RECT 345.200 154.300 346.000 154.400 ;
        RECT 364.400 154.300 365.200 154.400 ;
        RECT 369.200 154.300 370.000 154.400 ;
        RECT 345.200 153.700 370.000 154.300 ;
        RECT 345.200 153.600 346.000 153.700 ;
        RECT 364.400 153.600 365.200 153.700 ;
        RECT 369.200 153.600 370.000 153.700 ;
        RECT 374.000 154.300 374.800 154.400 ;
        RECT 380.400 154.300 381.200 154.400 ;
        RECT 374.000 153.700 381.200 154.300 ;
        RECT 374.000 153.600 374.800 153.700 ;
        RECT 380.400 153.600 381.200 153.700 ;
        RECT 404.400 154.300 405.200 154.400 ;
        RECT 439.600 154.300 440.400 154.400 ;
        RECT 404.400 153.700 440.400 154.300 ;
        RECT 404.400 153.600 405.200 153.700 ;
        RECT 439.600 153.600 440.400 153.700 ;
        RECT 532.400 154.300 533.200 154.400 ;
        RECT 538.800 154.300 539.600 154.400 ;
        RECT 532.400 153.700 539.600 154.300 ;
        RECT 532.400 153.600 533.200 153.700 ;
        RECT 538.800 153.600 539.600 153.700 ;
        RECT 12.400 152.300 13.200 152.400 ;
        RECT 31.600 152.300 32.400 152.400 ;
        RECT 12.400 151.700 32.400 152.300 ;
        RECT 12.400 151.600 13.200 151.700 ;
        RECT 31.600 151.600 32.400 151.700 ;
        RECT 36.400 152.300 37.200 152.400 ;
        RECT 55.600 152.300 56.400 152.400 ;
        RECT 36.400 151.700 56.400 152.300 ;
        RECT 36.400 151.600 37.200 151.700 ;
        RECT 55.600 151.600 56.400 151.700 ;
        RECT 74.800 152.300 75.600 152.400 ;
        RECT 158.000 152.300 158.800 152.400 ;
        RECT 74.800 151.700 158.800 152.300 ;
        RECT 74.800 151.600 75.600 151.700 ;
        RECT 158.000 151.600 158.800 151.700 ;
        RECT 209.200 152.300 210.000 152.400 ;
        RECT 225.200 152.300 226.000 152.400 ;
        RECT 209.200 151.700 226.000 152.300 ;
        RECT 209.200 151.600 210.000 151.700 ;
        RECT 225.200 151.600 226.000 151.700 ;
        RECT 351.600 152.300 352.400 152.400 ;
        RECT 374.000 152.300 374.800 152.400 ;
        RECT 351.600 151.700 374.800 152.300 ;
        RECT 351.600 151.600 352.400 151.700 ;
        RECT 374.000 151.600 374.800 151.700 ;
        RECT 385.200 152.300 386.000 152.400 ;
        RECT 415.600 152.300 416.400 152.400 ;
        RECT 450.800 152.300 451.600 152.400 ;
        RECT 385.200 151.700 451.600 152.300 ;
        RECT 385.200 151.600 386.000 151.700 ;
        RECT 415.600 151.600 416.400 151.700 ;
        RECT 450.800 151.600 451.600 151.700 ;
        RECT 462.000 152.300 462.800 152.400 ;
        RECT 473.200 152.300 474.000 152.400 ;
        RECT 462.000 151.700 474.000 152.300 ;
        RECT 462.000 151.600 462.800 151.700 ;
        RECT 473.200 151.600 474.000 151.700 ;
        RECT 513.200 152.300 514.000 152.400 ;
        RECT 522.800 152.300 523.600 152.400 ;
        RECT 527.600 152.300 528.400 152.400 ;
        RECT 513.200 151.700 528.400 152.300 ;
        RECT 513.200 151.600 514.000 151.700 ;
        RECT 522.800 151.600 523.600 151.700 ;
        RECT 527.600 151.600 528.400 151.700 ;
        RECT 530.800 151.600 531.600 152.400 ;
        RECT 7.600 150.300 8.400 150.400 ;
        RECT 10.800 150.300 11.600 150.400 ;
        RECT 15.600 150.300 16.400 150.400 ;
        RECT 20.400 150.300 21.200 150.400 ;
        RECT 7.600 149.700 21.200 150.300 ;
        RECT 7.600 149.600 8.400 149.700 ;
        RECT 10.800 149.600 11.600 149.700 ;
        RECT 15.600 149.600 16.400 149.700 ;
        RECT 20.400 149.600 21.200 149.700 ;
        RECT 28.400 150.300 29.200 150.400 ;
        RECT 33.200 150.300 34.000 150.400 ;
        RECT 28.400 149.700 34.000 150.300 ;
        RECT 28.400 149.600 29.200 149.700 ;
        RECT 33.200 149.600 34.000 149.700 ;
        RECT 41.200 150.300 42.000 150.400 ;
        RECT 47.600 150.300 48.400 150.400 ;
        RECT 41.200 149.700 48.400 150.300 ;
        RECT 41.200 149.600 42.000 149.700 ;
        RECT 47.600 149.600 48.400 149.700 ;
        RECT 49.200 150.300 50.000 150.400 ;
        RECT 60.400 150.300 61.200 150.400 ;
        RECT 49.200 149.700 61.200 150.300 ;
        RECT 49.200 149.600 50.000 149.700 ;
        RECT 60.400 149.600 61.200 149.700 ;
        RECT 86.000 150.300 86.800 150.400 ;
        RECT 97.200 150.300 98.000 150.400 ;
        RECT 86.000 149.700 98.000 150.300 ;
        RECT 86.000 149.600 86.800 149.700 ;
        RECT 97.200 149.600 98.000 149.700 ;
        RECT 98.800 150.300 99.600 150.400 ;
        RECT 106.800 150.300 107.600 150.400 ;
        RECT 114.800 150.300 115.600 150.400 ;
        RECT 126.000 150.300 126.800 150.400 ;
        RECT 98.800 149.700 126.800 150.300 ;
        RECT 98.800 149.600 99.600 149.700 ;
        RECT 106.800 149.600 107.600 149.700 ;
        RECT 114.800 149.600 115.600 149.700 ;
        RECT 126.000 149.600 126.800 149.700 ;
        RECT 164.400 150.300 165.200 150.400 ;
        RECT 172.400 150.300 173.200 150.400 ;
        RECT 164.400 149.700 173.200 150.300 ;
        RECT 164.400 149.600 165.200 149.700 ;
        RECT 172.400 149.600 173.200 149.700 ;
        RECT 214.000 149.600 214.800 150.400 ;
        RECT 246.000 150.300 246.800 150.400 ;
        RECT 255.600 150.300 256.400 150.400 ;
        RECT 263.600 150.300 264.400 150.400 ;
        RECT 266.800 150.300 267.600 150.400 ;
        RECT 246.000 149.700 267.600 150.300 ;
        RECT 246.000 149.600 246.800 149.700 ;
        RECT 255.600 149.600 256.400 149.700 ;
        RECT 263.600 149.600 264.400 149.700 ;
        RECT 266.800 149.600 267.600 149.700 ;
        RECT 281.200 150.300 282.000 150.400 ;
        RECT 318.000 150.300 318.800 150.400 ;
        RECT 281.200 149.700 318.800 150.300 ;
        RECT 281.200 149.600 282.000 149.700 ;
        RECT 318.000 149.600 318.800 149.700 ;
        RECT 348.400 150.300 349.200 150.400 ;
        RECT 364.400 150.300 365.200 150.400 ;
        RECT 348.400 149.700 365.200 150.300 ;
        RECT 348.400 149.600 349.200 149.700 ;
        RECT 364.400 149.600 365.200 149.700 ;
        RECT 367.600 150.300 368.400 150.400 ;
        RECT 388.400 150.300 389.200 150.400 ;
        RECT 367.600 149.700 389.200 150.300 ;
        RECT 367.600 149.600 368.400 149.700 ;
        RECT 388.400 149.600 389.200 149.700 ;
        RECT 409.200 150.300 410.000 150.400 ;
        RECT 412.400 150.300 413.200 150.400 ;
        RECT 409.200 149.700 413.200 150.300 ;
        RECT 409.200 149.600 410.000 149.700 ;
        RECT 412.400 149.600 413.200 149.700 ;
        RECT 428.400 150.300 429.200 150.400 ;
        RECT 458.800 150.300 459.600 150.400 ;
        RECT 428.400 149.700 459.600 150.300 ;
        RECT 428.400 149.600 429.200 149.700 ;
        RECT 458.800 149.600 459.600 149.700 ;
        RECT 466.800 150.300 467.600 150.400 ;
        RECT 473.200 150.300 474.000 150.400 ;
        RECT 466.800 149.700 474.000 150.300 ;
        RECT 466.800 149.600 467.600 149.700 ;
        RECT 473.200 149.600 474.000 149.700 ;
        RECT 478.000 150.300 478.800 150.400 ;
        RECT 487.600 150.300 488.400 150.400 ;
        RECT 492.400 150.300 493.200 150.400 ;
        RECT 478.000 149.700 493.200 150.300 ;
        RECT 478.000 149.600 478.800 149.700 ;
        RECT 487.600 149.600 488.400 149.700 ;
        RECT 492.400 149.600 493.200 149.700 ;
        RECT 506.800 150.300 507.600 150.400 ;
        RECT 516.400 150.300 517.200 150.400 ;
        RECT 506.800 149.700 517.200 150.300 ;
        RECT 506.800 149.600 507.600 149.700 ;
        RECT 516.400 149.600 517.200 149.700 ;
        RECT 524.400 150.300 525.200 150.400 ;
        RECT 529.200 150.300 530.000 150.400 ;
        RECT 524.400 149.700 530.000 150.300 ;
        RECT 524.400 149.600 525.200 149.700 ;
        RECT 529.200 149.600 530.000 149.700 ;
        RECT 534.000 150.300 534.800 150.400 ;
        RECT 540.400 150.300 541.200 150.400 ;
        RECT 534.000 149.700 541.200 150.300 ;
        RECT 534.000 149.600 534.800 149.700 ;
        RECT 540.400 149.600 541.200 149.700 ;
        RECT 543.600 150.300 544.400 150.400 ;
        RECT 548.400 150.300 549.200 150.400 ;
        RECT 543.600 149.700 549.200 150.300 ;
        RECT 543.600 149.600 544.400 149.700 ;
        RECT 548.400 149.600 549.200 149.700 ;
        RECT 9.200 148.300 10.000 148.400 ;
        RECT 14.000 148.300 14.800 148.400 ;
        RECT 9.200 147.700 14.800 148.300 ;
        RECT 9.200 147.600 10.000 147.700 ;
        RECT 14.000 147.600 14.800 147.700 ;
        RECT 31.600 148.300 32.400 148.400 ;
        RECT 68.400 148.300 69.200 148.400 ;
        RECT 31.600 147.700 69.200 148.300 ;
        RECT 31.600 147.600 32.400 147.700 ;
        RECT 68.400 147.600 69.200 147.700 ;
        RECT 82.800 148.300 83.600 148.400 ;
        RECT 89.200 148.300 90.000 148.400 ;
        RECT 134.000 148.300 134.800 148.400 ;
        RECT 82.800 147.700 90.000 148.300 ;
        RECT 82.800 147.600 83.600 147.700 ;
        RECT 89.200 147.600 90.000 147.700 ;
        RECT 132.500 147.700 134.800 148.300 ;
        RECT 18.800 146.300 19.600 146.400 ;
        RECT 38.000 146.300 38.800 146.400 ;
        RECT 18.800 145.700 38.800 146.300 ;
        RECT 18.800 145.600 19.600 145.700 ;
        RECT 38.000 145.600 38.800 145.700 ;
        RECT 39.600 146.300 40.400 146.400 ;
        RECT 46.000 146.300 46.800 146.400 ;
        RECT 58.800 146.300 59.600 146.400 ;
        RECT 62.000 146.300 62.800 146.400 ;
        RECT 39.600 145.700 62.800 146.300 ;
        RECT 39.600 145.600 40.400 145.700 ;
        RECT 46.000 145.600 46.800 145.700 ;
        RECT 58.800 145.600 59.600 145.700 ;
        RECT 62.000 145.600 62.800 145.700 ;
        RECT 66.800 146.300 67.600 146.400 ;
        RECT 78.000 146.300 78.800 146.400 ;
        RECT 66.800 145.700 78.800 146.300 ;
        RECT 66.800 145.600 67.600 145.700 ;
        RECT 78.000 145.600 78.800 145.700 ;
        RECT 97.200 146.300 98.000 146.400 ;
        RECT 103.600 146.300 104.400 146.400 ;
        RECT 97.200 145.700 104.400 146.300 ;
        RECT 97.200 145.600 98.000 145.700 ;
        RECT 103.600 145.600 104.400 145.700 ;
        RECT 121.200 146.300 122.000 146.400 ;
        RECT 132.500 146.300 133.100 147.700 ;
        RECT 134.000 147.600 134.800 147.700 ;
        RECT 196.400 148.300 197.200 148.400 ;
        RECT 207.600 148.300 208.400 148.400 ;
        RECT 223.600 148.300 224.400 148.400 ;
        RECT 196.400 147.700 224.400 148.300 ;
        RECT 196.400 147.600 197.200 147.700 ;
        RECT 207.600 147.600 208.400 147.700 ;
        RECT 223.600 147.600 224.400 147.700 ;
        RECT 228.400 148.300 229.200 148.400 ;
        RECT 231.600 148.300 232.400 148.400 ;
        RECT 228.400 147.700 232.400 148.300 ;
        RECT 228.400 147.600 229.200 147.700 ;
        RECT 231.600 147.600 232.400 147.700 ;
        RECT 257.200 148.300 258.000 148.400 ;
        RECT 271.600 148.300 272.400 148.400 ;
        RECT 257.200 147.700 272.400 148.300 ;
        RECT 257.200 147.600 258.000 147.700 ;
        RECT 271.600 147.600 272.400 147.700 ;
        RECT 354.800 148.300 355.600 148.400 ;
        RECT 372.400 148.300 373.200 148.400 ;
        RECT 375.600 148.300 376.400 148.400 ;
        RECT 354.800 147.700 376.400 148.300 ;
        RECT 354.800 147.600 355.600 147.700 ;
        RECT 372.400 147.600 373.200 147.700 ;
        RECT 375.600 147.600 376.400 147.700 ;
        RECT 380.400 148.300 381.200 148.400 ;
        RECT 386.800 148.300 387.600 148.400 ;
        RECT 380.400 147.700 387.600 148.300 ;
        RECT 380.400 147.600 381.200 147.700 ;
        RECT 386.800 147.600 387.600 147.700 ;
        RECT 390.000 148.300 390.800 148.400 ;
        RECT 410.800 148.300 411.600 148.400 ;
        RECT 390.000 147.700 411.600 148.300 ;
        RECT 390.000 147.600 390.800 147.700 ;
        RECT 410.800 147.600 411.600 147.700 ;
        RECT 425.200 148.300 426.000 148.400 ;
        RECT 428.400 148.300 429.200 148.400 ;
        RECT 425.200 147.700 429.200 148.300 ;
        RECT 425.200 147.600 426.000 147.700 ;
        RECT 428.400 147.600 429.200 147.700 ;
        RECT 466.800 148.300 467.600 148.400 ;
        RECT 474.800 148.300 475.600 148.400 ;
        RECT 466.800 147.700 475.600 148.300 ;
        RECT 466.800 147.600 467.600 147.700 ;
        RECT 474.800 147.600 475.600 147.700 ;
        RECT 526.000 148.300 526.800 148.400 ;
        RECT 534.000 148.300 534.800 148.400 ;
        RECT 526.000 147.700 534.800 148.300 ;
        RECT 526.000 147.600 526.800 147.700 ;
        RECT 534.000 147.600 534.800 147.700 ;
        RECT 540.400 148.300 541.200 148.400 ;
        RECT 543.600 148.300 544.400 148.400 ;
        RECT 540.400 147.700 544.400 148.300 ;
        RECT 540.400 147.600 541.200 147.700 ;
        RECT 543.600 147.600 544.400 147.700 ;
        RECT 562.800 148.300 563.600 148.400 ;
        RECT 570.800 148.300 571.600 148.400 ;
        RECT 562.800 147.700 571.600 148.300 ;
        RECT 562.800 147.600 563.600 147.700 ;
        RECT 570.800 147.600 571.600 147.700 ;
        RECT 121.200 145.700 133.100 146.300 ;
        RECT 134.000 146.300 134.800 146.400 ;
        RECT 146.800 146.300 147.600 146.400 ;
        RECT 134.000 145.700 147.600 146.300 ;
        RECT 121.200 145.600 122.000 145.700 ;
        RECT 134.000 145.600 134.800 145.700 ;
        RECT 146.800 145.600 147.600 145.700 ;
        RECT 151.600 146.300 152.400 146.400 ;
        RECT 193.200 146.300 194.000 146.400 ;
        RECT 198.000 146.300 198.800 146.400 ;
        RECT 214.000 146.300 214.800 146.400 ;
        RECT 231.600 146.300 232.400 146.400 ;
        RECT 151.600 145.700 232.400 146.300 ;
        RECT 151.600 145.600 152.400 145.700 ;
        RECT 193.200 145.600 194.000 145.700 ;
        RECT 198.000 145.600 198.800 145.700 ;
        RECT 214.000 145.600 214.800 145.700 ;
        RECT 231.600 145.600 232.400 145.700 ;
        RECT 244.400 146.300 245.200 146.400 ;
        RECT 258.800 146.300 259.600 146.400 ;
        RECT 244.400 145.700 259.600 146.300 ;
        RECT 244.400 145.600 245.200 145.700 ;
        RECT 258.800 145.600 259.600 145.700 ;
        RECT 263.600 146.300 264.400 146.400 ;
        RECT 270.000 146.300 270.800 146.400 ;
        RECT 274.800 146.300 275.600 146.400 ;
        RECT 263.600 145.700 275.600 146.300 ;
        RECT 263.600 145.600 264.400 145.700 ;
        RECT 270.000 145.600 270.800 145.700 ;
        RECT 274.800 145.600 275.600 145.700 ;
        RECT 330.800 146.300 331.600 146.400 ;
        RECT 337.200 146.300 338.000 146.400 ;
        RECT 346.800 146.300 347.600 146.400 ;
        RECT 358.000 146.300 358.800 146.400 ;
        RECT 362.800 146.300 363.600 146.400 ;
        RECT 330.800 145.700 363.600 146.300 ;
        RECT 330.800 145.600 331.600 145.700 ;
        RECT 337.200 145.600 338.000 145.700 ;
        RECT 346.800 145.600 347.600 145.700 ;
        RECT 358.000 145.600 358.800 145.700 ;
        RECT 362.800 145.600 363.600 145.700 ;
        RECT 374.000 146.300 374.800 146.400 ;
        RECT 382.000 146.300 382.800 146.400 ;
        RECT 374.000 145.700 382.800 146.300 ;
        RECT 386.900 146.300 387.500 147.600 ;
        RECT 394.800 146.300 395.600 146.400 ;
        RECT 386.900 145.700 395.600 146.300 ;
        RECT 374.000 145.600 374.800 145.700 ;
        RECT 382.000 145.600 382.800 145.700 ;
        RECT 394.800 145.600 395.600 145.700 ;
        RECT 410.800 146.300 411.600 146.400 ;
        RECT 420.400 146.300 421.200 146.400 ;
        RECT 410.800 145.700 421.200 146.300 ;
        RECT 410.800 145.600 411.600 145.700 ;
        RECT 420.400 145.600 421.200 145.700 ;
        RECT 431.600 146.300 432.400 146.400 ;
        RECT 444.400 146.300 445.200 146.400 ;
        RECT 431.600 145.700 445.200 146.300 ;
        RECT 431.600 145.600 432.400 145.700 ;
        RECT 444.400 145.600 445.200 145.700 ;
        RECT 516.400 146.300 517.200 146.400 ;
        RECT 532.400 146.300 533.200 146.400 ;
        RECT 516.400 145.700 533.200 146.300 ;
        RECT 516.400 145.600 517.200 145.700 ;
        RECT 532.400 145.600 533.200 145.700 ;
        RECT 535.600 146.300 536.400 146.400 ;
        RECT 540.400 146.300 541.200 146.400 ;
        RECT 535.600 145.700 541.200 146.300 ;
        RECT 535.600 145.600 536.400 145.700 ;
        RECT 540.400 145.600 541.200 145.700 ;
        RECT 542.000 146.300 542.800 146.400 ;
        RECT 551.600 146.300 552.400 146.400 ;
        RECT 553.200 146.300 554.000 146.400 ;
        RECT 542.000 145.700 554.000 146.300 ;
        RECT 542.000 145.600 542.800 145.700 ;
        RECT 551.600 145.600 552.400 145.700 ;
        RECT 553.200 145.600 554.000 145.700 ;
        RECT 18.800 144.300 19.600 144.400 ;
        RECT 41.200 144.300 42.000 144.400 ;
        RECT 18.800 143.700 42.000 144.300 ;
        RECT 18.800 143.600 19.600 143.700 ;
        RECT 41.200 143.600 42.000 143.700 ;
        RECT 44.400 144.300 45.200 144.400 ;
        RECT 55.600 144.300 56.400 144.400 ;
        RECT 44.400 143.700 56.400 144.300 ;
        RECT 44.400 143.600 45.200 143.700 ;
        RECT 55.600 143.600 56.400 143.700 ;
        RECT 60.400 144.300 61.200 144.400 ;
        RECT 65.200 144.300 66.000 144.400 ;
        RECT 60.400 143.700 66.000 144.300 ;
        RECT 60.400 143.600 61.200 143.700 ;
        RECT 65.200 143.600 66.000 143.700 ;
        RECT 89.200 144.300 90.000 144.400 ;
        RECT 122.800 144.300 123.600 144.400 ;
        RECT 89.200 143.700 123.600 144.300 ;
        RECT 89.200 143.600 90.000 143.700 ;
        RECT 122.800 143.600 123.600 143.700 ;
        RECT 158.000 144.300 158.800 144.400 ;
        RECT 162.800 144.300 163.600 144.400 ;
        RECT 158.000 143.700 163.600 144.300 ;
        RECT 158.000 143.600 158.800 143.700 ;
        RECT 162.800 143.600 163.600 143.700 ;
        RECT 220.400 144.300 221.200 144.400 ;
        RECT 228.400 144.300 229.200 144.400 ;
        RECT 220.400 143.700 229.200 144.300 ;
        RECT 220.400 143.600 221.200 143.700 ;
        RECT 228.400 143.600 229.200 143.700 ;
        RECT 258.800 144.300 259.600 144.400 ;
        RECT 265.200 144.300 266.000 144.400 ;
        RECT 258.800 143.700 266.000 144.300 ;
        RECT 258.800 143.600 259.600 143.700 ;
        RECT 265.200 143.600 266.000 143.700 ;
        RECT 279.600 144.300 280.400 144.400 ;
        RECT 287.600 144.300 288.400 144.400 ;
        RECT 279.600 143.700 288.400 144.300 ;
        RECT 279.600 143.600 280.400 143.700 ;
        RECT 287.600 143.600 288.400 143.700 ;
        RECT 356.400 144.300 357.200 144.400 ;
        RECT 380.400 144.300 381.200 144.400 ;
        RECT 356.400 143.700 381.200 144.300 ;
        RECT 356.400 143.600 357.200 143.700 ;
        RECT 380.400 143.600 381.200 143.700 ;
        RECT 385.200 144.300 386.000 144.400 ;
        RECT 401.200 144.300 402.000 144.400 ;
        RECT 385.200 143.700 402.000 144.300 ;
        RECT 385.200 143.600 386.000 143.700 ;
        RECT 401.200 143.600 402.000 143.700 ;
        RECT 409.200 144.300 410.000 144.400 ;
        RECT 410.800 144.300 411.600 144.400 ;
        RECT 409.200 143.700 411.600 144.300 ;
        RECT 409.200 143.600 410.000 143.700 ;
        RECT 410.800 143.600 411.600 143.700 ;
        RECT 428.400 144.300 429.200 144.400 ;
        RECT 433.200 144.300 434.000 144.400 ;
        RECT 428.400 143.700 434.000 144.300 ;
        RECT 428.400 143.600 429.200 143.700 ;
        RECT 433.200 143.600 434.000 143.700 ;
        RECT 25.200 142.300 26.000 142.400 ;
        RECT 34.800 142.300 35.600 142.400 ;
        RECT 47.600 142.300 48.400 142.400 ;
        RECT 25.200 141.700 48.400 142.300 ;
        RECT 25.200 141.600 26.000 141.700 ;
        RECT 34.800 141.600 35.600 141.700 ;
        RECT 47.600 141.600 48.400 141.700 ;
        RECT 74.800 142.300 75.600 142.400 ;
        RECT 98.800 142.300 99.600 142.400 ;
        RECT 127.600 142.300 128.400 142.400 ;
        RECT 135.600 142.300 136.400 142.400 ;
        RECT 183.600 142.300 184.400 142.400 ;
        RECT 74.800 141.700 184.400 142.300 ;
        RECT 74.800 141.600 75.600 141.700 ;
        RECT 98.800 141.600 99.600 141.700 ;
        RECT 127.600 141.600 128.400 141.700 ;
        RECT 135.600 141.600 136.400 141.700 ;
        RECT 183.600 141.600 184.400 141.700 ;
        RECT 206.000 142.300 206.800 142.400 ;
        RECT 278.000 142.300 278.800 142.400 ;
        RECT 206.000 141.700 278.800 142.300 ;
        RECT 206.000 141.600 206.800 141.700 ;
        RECT 278.000 141.600 278.800 141.700 ;
        RECT 311.600 142.300 312.400 142.400 ;
        RECT 326.000 142.300 326.800 142.400 ;
        RECT 348.400 142.300 349.200 142.400 ;
        RECT 311.600 141.700 349.200 142.300 ;
        RECT 311.600 141.600 312.400 141.700 ;
        RECT 326.000 141.600 326.800 141.700 ;
        RECT 348.400 141.600 349.200 141.700 ;
        RECT 351.600 142.300 352.400 142.400 ;
        RECT 362.800 142.300 363.600 142.400 ;
        RECT 351.600 141.700 363.600 142.300 ;
        RECT 351.600 141.600 352.400 141.700 ;
        RECT 362.800 141.600 363.600 141.700 ;
        RECT 414.000 142.300 414.800 142.400 ;
        RECT 431.600 142.300 432.400 142.400 ;
        RECT 414.000 141.700 432.400 142.300 ;
        RECT 414.000 141.600 414.800 141.700 ;
        RECT 431.600 141.600 432.400 141.700 ;
        RECT 455.600 142.300 456.400 142.400 ;
        RECT 462.000 142.300 462.800 142.400 ;
        RECT 455.600 141.700 462.800 142.300 ;
        RECT 455.600 141.600 456.400 141.700 ;
        RECT 462.000 141.600 462.800 141.700 ;
        RECT 522.800 142.300 523.600 142.400 ;
        RECT 548.400 142.300 549.200 142.400 ;
        RECT 522.800 141.700 549.200 142.300 ;
        RECT 522.800 141.600 523.600 141.700 ;
        RECT 548.400 141.600 549.200 141.700 ;
        RECT 550.000 142.300 550.800 142.400 ;
        RECT 553.200 142.300 554.000 142.400 ;
        RECT 550.000 141.700 554.000 142.300 ;
        RECT 550.000 141.600 550.800 141.700 ;
        RECT 553.200 141.600 554.000 141.700 ;
        RECT 28.400 140.300 29.200 140.400 ;
        RECT 33.200 140.300 34.000 140.400 ;
        RECT 28.400 139.700 34.000 140.300 ;
        RECT 28.400 139.600 29.200 139.700 ;
        RECT 33.200 139.600 34.000 139.700 ;
        RECT 62.000 140.300 62.800 140.400 ;
        RECT 90.800 140.300 91.600 140.400 ;
        RECT 62.000 139.700 91.600 140.300 ;
        RECT 62.000 139.600 62.800 139.700 ;
        RECT 90.800 139.600 91.600 139.700 ;
        RECT 223.600 140.300 224.400 140.400 ;
        RECT 226.800 140.300 227.600 140.400 ;
        RECT 223.600 139.700 227.600 140.300 ;
        RECT 223.600 139.600 224.400 139.700 ;
        RECT 226.800 139.600 227.600 139.700 ;
        RECT 374.000 140.300 374.800 140.400 ;
        RECT 426.800 140.300 427.600 140.400 ;
        RECT 374.000 139.700 427.600 140.300 ;
        RECT 374.000 139.600 374.800 139.700 ;
        RECT 426.800 139.600 427.600 139.700 ;
        RECT 438.000 140.300 438.800 140.400 ;
        RECT 450.800 140.300 451.600 140.400 ;
        RECT 438.000 139.700 451.600 140.300 ;
        RECT 438.000 139.600 438.800 139.700 ;
        RECT 450.800 139.600 451.600 139.700 ;
        RECT 510.000 140.300 510.800 140.400 ;
        RECT 566.000 140.300 566.800 140.400 ;
        RECT 510.000 139.700 566.800 140.300 ;
        RECT 510.000 139.600 510.800 139.700 ;
        RECT 566.000 139.600 566.800 139.700 ;
        RECT 14.000 138.300 14.800 138.400 ;
        RECT 30.000 138.300 30.800 138.400 ;
        RECT 14.000 137.700 30.800 138.300 ;
        RECT 14.000 137.600 14.800 137.700 ;
        RECT 30.000 137.600 30.800 137.700 ;
        RECT 86.000 138.300 86.800 138.400 ;
        RECT 90.800 138.300 91.600 138.400 ;
        RECT 86.000 137.700 91.600 138.300 ;
        RECT 86.000 137.600 86.800 137.700 ;
        RECT 90.800 137.600 91.600 137.700 ;
        RECT 92.400 138.300 93.200 138.400 ;
        RECT 118.000 138.300 118.800 138.400 ;
        RECT 92.400 137.700 118.800 138.300 ;
        RECT 92.400 137.600 93.200 137.700 ;
        RECT 118.000 137.600 118.800 137.700 ;
        RECT 201.200 138.300 202.000 138.400 ;
        RECT 225.200 138.300 226.000 138.400 ;
        RECT 201.200 137.700 226.000 138.300 ;
        RECT 201.200 137.600 202.000 137.700 ;
        RECT 225.200 137.600 226.000 137.700 ;
        RECT 276.400 138.300 277.200 138.400 ;
        RECT 281.200 138.300 282.000 138.400 ;
        RECT 276.400 137.700 282.000 138.300 ;
        RECT 276.400 137.600 277.200 137.700 ;
        RECT 281.200 137.600 282.000 137.700 ;
        RECT 342.000 138.300 342.800 138.400 ;
        RECT 343.600 138.300 344.400 138.400 ;
        RECT 342.000 137.700 344.400 138.300 ;
        RECT 342.000 137.600 342.800 137.700 ;
        RECT 343.600 137.600 344.400 137.700 ;
        RECT 364.400 138.300 365.200 138.400 ;
        RECT 369.200 138.300 370.000 138.400 ;
        RECT 364.400 137.700 370.000 138.300 ;
        RECT 364.400 137.600 365.200 137.700 ;
        RECT 369.200 137.600 370.000 137.700 ;
        RECT 370.800 138.300 371.600 138.400 ;
        RECT 383.600 138.300 384.400 138.400 ;
        RECT 370.800 137.700 384.400 138.300 ;
        RECT 370.800 137.600 371.600 137.700 ;
        RECT 383.600 137.600 384.400 137.700 ;
        RECT 386.800 138.300 387.600 138.400 ;
        RECT 404.400 138.300 405.200 138.400 ;
        RECT 386.800 137.700 405.200 138.300 ;
        RECT 386.800 137.600 387.600 137.700 ;
        RECT 404.400 137.600 405.200 137.700 ;
        RECT 426.800 138.300 427.600 138.400 ;
        RECT 430.000 138.300 430.800 138.400 ;
        RECT 426.800 137.700 430.800 138.300 ;
        RECT 426.800 137.600 427.600 137.700 ;
        RECT 430.000 137.600 430.800 137.700 ;
        RECT 444.400 138.300 445.200 138.400 ;
        RECT 454.000 138.300 454.800 138.400 ;
        RECT 444.400 137.700 454.800 138.300 ;
        RECT 444.400 137.600 445.200 137.700 ;
        RECT 454.000 137.600 454.800 137.700 ;
        RECT 521.200 138.300 522.000 138.400 ;
        RECT 556.400 138.300 557.200 138.400 ;
        RECT 521.200 137.700 557.200 138.300 ;
        RECT 521.200 137.600 522.000 137.700 ;
        RECT 556.400 137.600 557.200 137.700 ;
        RECT 1.200 136.300 2.000 136.400 ;
        RECT 7.600 136.300 8.400 136.400 ;
        RECT 1.200 135.700 8.400 136.300 ;
        RECT 1.200 135.600 2.000 135.700 ;
        RECT 7.600 135.600 8.400 135.700 ;
        RECT 23.600 136.300 24.400 136.400 ;
        RECT 33.200 136.300 34.000 136.400 ;
        RECT 38.000 136.300 38.800 136.400 ;
        RECT 23.600 135.700 38.800 136.300 ;
        RECT 23.600 135.600 24.400 135.700 ;
        RECT 33.200 135.600 34.000 135.700 ;
        RECT 38.000 135.600 38.800 135.700 ;
        RECT 68.400 136.300 69.200 136.400 ;
        RECT 70.000 136.300 70.800 136.400 ;
        RECT 82.800 136.300 83.600 136.400 ;
        RECT 68.400 135.700 83.600 136.300 ;
        RECT 68.400 135.600 69.200 135.700 ;
        RECT 70.000 135.600 70.800 135.700 ;
        RECT 82.800 135.600 83.600 135.700 ;
        RECT 110.000 136.300 110.800 136.400 ;
        RECT 146.800 136.300 147.600 136.400 ;
        RECT 110.000 135.700 147.600 136.300 ;
        RECT 110.000 135.600 110.800 135.700 ;
        RECT 146.800 135.600 147.600 135.700 ;
        RECT 148.400 136.300 149.200 136.400 ;
        RECT 156.400 136.300 157.200 136.400 ;
        RECT 148.400 135.700 157.200 136.300 ;
        RECT 148.400 135.600 149.200 135.700 ;
        RECT 156.400 135.600 157.200 135.700 ;
        RECT 193.200 136.300 194.000 136.400 ;
        RECT 198.000 136.300 198.800 136.400 ;
        RECT 206.000 136.300 206.800 136.400 ;
        RECT 193.200 135.700 206.800 136.300 ;
        RECT 193.200 135.600 194.000 135.700 ;
        RECT 198.000 135.600 198.800 135.700 ;
        RECT 206.000 135.600 206.800 135.700 ;
        RECT 226.800 136.300 227.600 136.400 ;
        RECT 230.000 136.300 230.800 136.400 ;
        RECT 226.800 135.700 230.800 136.300 ;
        RECT 226.800 135.600 227.600 135.700 ;
        RECT 230.000 135.600 230.800 135.700 ;
        RECT 250.800 136.300 251.600 136.400 ;
        RECT 295.600 136.300 296.400 136.400 ;
        RECT 250.800 135.700 296.400 136.300 ;
        RECT 250.800 135.600 251.600 135.700 ;
        RECT 295.600 135.600 296.400 135.700 ;
        RECT 358.000 136.300 358.800 136.400 ;
        RECT 367.600 136.300 368.400 136.400 ;
        RECT 377.200 136.300 378.000 136.400 ;
        RECT 358.000 135.700 378.000 136.300 ;
        RECT 358.000 135.600 358.800 135.700 ;
        RECT 367.600 135.600 368.400 135.700 ;
        RECT 377.200 135.600 378.000 135.700 ;
        RECT 378.800 136.300 379.600 136.400 ;
        RECT 386.800 136.300 387.600 136.400 ;
        RECT 388.400 136.300 389.200 136.400 ;
        RECT 378.800 135.700 389.200 136.300 ;
        RECT 378.800 135.600 379.600 135.700 ;
        RECT 386.800 135.600 387.600 135.700 ;
        RECT 388.400 135.600 389.200 135.700 ;
        RECT 399.600 136.300 400.400 136.400 ;
        RECT 449.200 136.300 450.000 136.400 ;
        RECT 466.800 136.300 467.600 136.400 ;
        RECT 577.200 136.300 578.000 136.400 ;
        RECT 399.600 135.700 448.300 136.300 ;
        RECT 399.600 135.600 400.400 135.700 ;
        RECT 4.400 134.300 5.200 134.400 ;
        RECT 28.400 134.300 29.200 134.400 ;
        RECT 4.400 133.700 29.200 134.300 ;
        RECT 4.400 133.600 5.200 133.700 ;
        RECT 28.400 133.600 29.200 133.700 ;
        RECT 76.400 134.300 77.200 134.400 ;
        RECT 92.400 134.300 93.200 134.400 ;
        RECT 116.400 134.300 117.200 134.400 ;
        RECT 76.400 133.700 117.200 134.300 ;
        RECT 76.400 133.600 77.200 133.700 ;
        RECT 92.400 133.600 93.200 133.700 ;
        RECT 116.400 133.600 117.200 133.700 ;
        RECT 126.000 134.300 126.800 134.400 ;
        RECT 130.800 134.300 131.600 134.400 ;
        RECT 126.000 133.700 131.600 134.300 ;
        RECT 126.000 133.600 126.800 133.700 ;
        RECT 130.800 133.600 131.600 133.700 ;
        RECT 178.800 134.300 179.600 134.400 ;
        RECT 183.600 134.300 184.400 134.400 ;
        RECT 196.400 134.300 197.200 134.400 ;
        RECT 178.800 133.700 197.200 134.300 ;
        RECT 178.800 133.600 179.600 133.700 ;
        RECT 183.600 133.600 184.400 133.700 ;
        RECT 196.400 133.600 197.200 133.700 ;
        RECT 214.000 134.300 214.800 134.400 ;
        RECT 215.600 134.300 216.400 134.400 ;
        RECT 214.000 133.700 216.400 134.300 ;
        RECT 214.000 133.600 214.800 133.700 ;
        RECT 215.600 133.600 216.400 133.700 ;
        RECT 223.600 134.300 224.400 134.400 ;
        RECT 228.400 134.300 229.200 134.400 ;
        RECT 223.600 133.700 229.200 134.300 ;
        RECT 223.600 133.600 224.400 133.700 ;
        RECT 228.400 133.600 229.200 133.700 ;
        RECT 231.600 134.300 232.400 134.400 ;
        RECT 238.000 134.300 238.800 134.400 ;
        RECT 231.600 133.700 238.800 134.300 ;
        RECT 231.600 133.600 232.400 133.700 ;
        RECT 238.000 133.600 238.800 133.700 ;
        RECT 255.600 134.300 256.400 134.400 ;
        RECT 262.000 134.300 262.800 134.400 ;
        RECT 265.200 134.300 266.000 134.400 ;
        RECT 255.600 133.700 266.000 134.300 ;
        RECT 255.600 133.600 256.400 133.700 ;
        RECT 262.000 133.600 262.800 133.700 ;
        RECT 265.200 133.600 266.000 133.700 ;
        RECT 268.400 134.300 269.200 134.400 ;
        RECT 281.200 134.300 282.000 134.400 ;
        RECT 268.400 133.700 282.000 134.300 ;
        RECT 268.400 133.600 269.200 133.700 ;
        RECT 281.200 133.600 282.000 133.700 ;
        RECT 294.000 134.300 294.800 134.400 ;
        RECT 305.200 134.300 306.000 134.400 ;
        RECT 294.000 133.700 306.000 134.300 ;
        RECT 294.000 133.600 294.800 133.700 ;
        RECT 305.200 133.600 306.000 133.700 ;
        RECT 335.600 134.300 336.400 134.400 ;
        RECT 348.400 134.300 349.200 134.400 ;
        RECT 335.600 133.700 349.200 134.300 ;
        RECT 335.600 133.600 336.400 133.700 ;
        RECT 348.400 133.600 349.200 133.700 ;
        RECT 361.200 134.300 362.000 134.400 ;
        RECT 367.600 134.300 368.400 134.400 ;
        RECT 372.400 134.300 373.200 134.400 ;
        RECT 390.000 134.300 390.800 134.400 ;
        RECT 398.000 134.300 398.800 134.400 ;
        RECT 420.400 134.300 421.200 134.400 ;
        RECT 361.200 133.700 373.200 134.300 ;
        RECT 361.200 133.600 362.000 133.700 ;
        RECT 367.600 133.600 368.400 133.700 ;
        RECT 372.400 133.600 373.200 133.700 ;
        RECT 375.700 133.700 421.200 134.300 ;
        RECT 447.700 134.300 448.300 135.700 ;
        RECT 449.200 135.700 467.600 136.300 ;
        RECT 449.200 135.600 450.000 135.700 ;
        RECT 466.800 135.600 467.600 135.700 ;
        RECT 532.500 135.700 578.000 136.300 ;
        RECT 532.500 134.400 533.100 135.700 ;
        RECT 577.200 135.600 578.000 135.700 ;
        RECT 468.400 134.300 469.200 134.400 ;
        RECT 447.700 133.700 469.200 134.300 ;
        RECT 23.600 132.300 24.400 132.400 ;
        RECT 44.400 132.300 45.200 132.400 ;
        RECT 23.600 131.700 45.200 132.300 ;
        RECT 23.600 131.600 24.400 131.700 ;
        RECT 44.400 131.600 45.200 131.700 ;
        RECT 57.200 132.300 58.000 132.400 ;
        RECT 62.000 132.300 62.800 132.400 ;
        RECT 57.200 131.700 62.800 132.300 ;
        RECT 57.200 131.600 58.000 131.700 ;
        RECT 62.000 131.600 62.800 131.700 ;
        RECT 78.000 132.300 78.800 132.400 ;
        RECT 94.000 132.300 94.800 132.400 ;
        RECT 78.000 131.700 94.800 132.300 ;
        RECT 78.000 131.600 78.800 131.700 ;
        RECT 94.000 131.600 94.800 131.700 ;
        RECT 108.400 132.300 109.200 132.400 ;
        RECT 113.200 132.300 114.000 132.400 ;
        RECT 108.400 131.700 114.000 132.300 ;
        RECT 108.400 131.600 109.200 131.700 ;
        RECT 113.200 131.600 114.000 131.700 ;
        RECT 114.800 132.300 115.600 132.400 ;
        RECT 126.000 132.300 126.800 132.400 ;
        RECT 114.800 131.700 126.800 132.300 ;
        RECT 114.800 131.600 115.600 131.700 ;
        RECT 126.000 131.600 126.800 131.700 ;
        RECT 156.400 132.300 157.200 132.400 ;
        RECT 164.400 132.300 165.200 132.400 ;
        RECT 156.400 131.700 165.200 132.300 ;
        RECT 156.400 131.600 157.200 131.700 ;
        RECT 164.400 131.600 165.200 131.700 ;
        RECT 170.800 132.300 171.600 132.400 ;
        RECT 182.000 132.300 182.800 132.400 ;
        RECT 188.400 132.300 189.200 132.400 ;
        RECT 193.200 132.300 194.000 132.400 ;
        RECT 215.600 132.300 216.400 132.400 ;
        RECT 234.800 132.300 235.600 132.400 ;
        RECT 170.800 131.700 216.400 132.300 ;
        RECT 170.800 131.600 171.600 131.700 ;
        RECT 182.000 131.600 182.800 131.700 ;
        RECT 188.400 131.600 189.200 131.700 ;
        RECT 193.200 131.600 194.000 131.700 ;
        RECT 215.600 131.600 216.400 131.700 ;
        RECT 222.100 131.700 235.600 132.300 ;
        RECT 222.100 130.400 222.700 131.700 ;
        RECT 234.800 131.600 235.600 131.700 ;
        RECT 244.400 132.300 245.200 132.400 ;
        RECT 247.600 132.300 248.400 132.400 ;
        RECT 284.400 132.300 285.200 132.400 ;
        RECT 298.800 132.300 299.600 132.400 ;
        RECT 318.000 132.300 318.800 132.400 ;
        RECT 244.400 131.700 318.800 132.300 ;
        RECT 244.400 131.600 245.200 131.700 ;
        RECT 247.600 131.600 248.400 131.700 ;
        RECT 284.400 131.600 285.200 131.700 ;
        RECT 298.800 131.600 299.600 131.700 ;
        RECT 318.000 131.600 318.800 131.700 ;
        RECT 354.800 132.300 355.600 132.400 ;
        RECT 375.700 132.300 376.300 133.700 ;
        RECT 390.000 133.600 390.800 133.700 ;
        RECT 398.000 133.600 398.800 133.700 ;
        RECT 420.400 133.600 421.200 133.700 ;
        RECT 468.400 133.600 469.200 133.700 ;
        RECT 490.800 134.300 491.600 134.400 ;
        RECT 513.200 134.300 514.000 134.400 ;
        RECT 532.400 134.300 533.200 134.400 ;
        RECT 490.800 133.700 533.200 134.300 ;
        RECT 490.800 133.600 491.600 133.700 ;
        RECT 513.200 133.600 514.000 133.700 ;
        RECT 532.400 133.600 533.200 133.700 ;
        RECT 538.800 134.300 539.600 134.400 ;
        RECT 543.600 134.300 544.400 134.400 ;
        RECT 550.000 134.300 550.800 134.400 ;
        RECT 538.800 133.700 550.800 134.300 ;
        RECT 538.800 133.600 539.600 133.700 ;
        RECT 543.600 133.600 544.400 133.700 ;
        RECT 550.000 133.600 550.800 133.700 ;
        RECT 354.800 131.700 376.300 132.300 ;
        RECT 385.200 132.300 386.000 132.400 ;
        RECT 399.600 132.300 400.400 132.400 ;
        RECT 385.200 131.700 400.400 132.300 ;
        RECT 354.800 131.600 355.600 131.700 ;
        RECT 385.200 131.600 386.000 131.700 ;
        RECT 399.600 131.600 400.400 131.700 ;
        RECT 417.200 132.300 418.000 132.400 ;
        RECT 430.000 132.300 430.800 132.400 ;
        RECT 417.200 131.700 430.800 132.300 ;
        RECT 417.200 131.600 418.000 131.700 ;
        RECT 430.000 131.600 430.800 131.700 ;
        RECT 434.800 132.300 435.600 132.400 ;
        RECT 441.200 132.300 442.000 132.400 ;
        RECT 457.200 132.300 458.000 132.400 ;
        RECT 434.800 131.700 458.000 132.300 ;
        RECT 434.800 131.600 435.600 131.700 ;
        RECT 441.200 131.600 442.000 131.700 ;
        RECT 457.200 131.600 458.000 131.700 ;
        RECT 471.600 132.300 472.400 132.400 ;
        RECT 474.800 132.300 475.600 132.400 ;
        RECT 471.600 131.700 475.600 132.300 ;
        RECT 471.600 131.600 472.400 131.700 ;
        RECT 474.800 131.600 475.600 131.700 ;
        RECT 30.000 130.300 30.800 130.400 ;
        RECT 38.000 130.300 38.800 130.400 ;
        RECT 41.200 130.300 42.000 130.400 ;
        RECT 52.400 130.300 53.200 130.400 ;
        RECT 30.000 129.700 53.200 130.300 ;
        RECT 30.000 129.600 30.800 129.700 ;
        RECT 38.000 129.600 38.800 129.700 ;
        RECT 41.200 129.600 42.000 129.700 ;
        RECT 52.400 129.600 53.200 129.700 ;
        RECT 54.000 130.300 54.800 130.400 ;
        RECT 57.200 130.300 58.000 130.400 ;
        RECT 54.000 129.700 58.000 130.300 ;
        RECT 54.000 129.600 54.800 129.700 ;
        RECT 57.200 129.600 58.000 129.700 ;
        RECT 65.200 130.300 66.000 130.400 ;
        RECT 79.600 130.300 80.400 130.400 ;
        RECT 81.200 130.300 82.000 130.400 ;
        RECT 111.600 130.300 112.400 130.400 ;
        RECT 119.600 130.300 120.400 130.400 ;
        RECT 148.400 130.300 149.200 130.400 ;
        RECT 65.200 129.700 149.200 130.300 ;
        RECT 65.200 129.600 66.000 129.700 ;
        RECT 79.600 129.600 80.400 129.700 ;
        RECT 81.200 129.600 82.000 129.700 ;
        RECT 111.600 129.600 112.400 129.700 ;
        RECT 119.600 129.600 120.400 129.700 ;
        RECT 148.400 129.600 149.200 129.700 ;
        RECT 185.200 130.300 186.000 130.400 ;
        RECT 201.200 130.300 202.000 130.400 ;
        RECT 185.200 129.700 202.000 130.300 ;
        RECT 185.200 129.600 186.000 129.700 ;
        RECT 201.200 129.600 202.000 129.700 ;
        RECT 210.800 130.300 211.600 130.400 ;
        RECT 218.800 130.300 219.600 130.400 ;
        RECT 222.000 130.300 222.800 130.400 ;
        RECT 210.800 129.700 222.800 130.300 ;
        RECT 210.800 129.600 211.600 129.700 ;
        RECT 218.800 129.600 219.600 129.700 ;
        RECT 222.000 129.600 222.800 129.700 ;
        RECT 223.600 130.300 224.400 130.400 ;
        RECT 231.600 130.300 232.400 130.400 ;
        RECT 252.400 130.300 253.200 130.400 ;
        RECT 223.600 129.700 253.200 130.300 ;
        RECT 223.600 129.600 224.400 129.700 ;
        RECT 231.600 129.600 232.400 129.700 ;
        RECT 252.400 129.600 253.200 129.700 ;
        RECT 268.400 130.300 269.200 130.400 ;
        RECT 271.600 130.300 272.400 130.400 ;
        RECT 268.400 129.700 272.400 130.300 ;
        RECT 268.400 129.600 269.200 129.700 ;
        RECT 271.600 129.600 272.400 129.700 ;
        RECT 287.600 130.300 288.400 130.400 ;
        RECT 289.200 130.300 290.000 130.400 ;
        RECT 287.600 129.700 290.000 130.300 ;
        RECT 287.600 129.600 288.400 129.700 ;
        RECT 289.200 129.600 290.000 129.700 ;
        RECT 343.600 130.300 344.400 130.400 ;
        RECT 380.400 130.300 381.200 130.400 ;
        RECT 415.600 130.300 416.400 130.400 ;
        RECT 343.600 129.700 416.400 130.300 ;
        RECT 343.600 129.600 344.400 129.700 ;
        RECT 380.400 129.600 381.200 129.700 ;
        RECT 415.600 129.600 416.400 129.700 ;
        RECT 465.200 130.300 466.000 130.400 ;
        RECT 471.600 130.300 472.400 130.400 ;
        RECT 465.200 129.700 472.400 130.300 ;
        RECT 465.200 129.600 466.000 129.700 ;
        RECT 471.600 129.600 472.400 129.700 ;
        RECT 526.000 130.300 526.800 130.400 ;
        RECT 535.600 130.300 536.400 130.400 ;
        RECT 526.000 129.700 536.400 130.300 ;
        RECT 526.000 129.600 526.800 129.700 ;
        RECT 535.600 129.600 536.400 129.700 ;
        RECT 537.200 130.300 538.000 130.400 ;
        RECT 543.600 130.300 544.400 130.400 ;
        RECT 537.200 129.700 544.400 130.300 ;
        RECT 537.200 129.600 538.000 129.700 ;
        RECT 543.600 129.600 544.400 129.700 ;
        RECT 1.200 128.300 2.000 128.400 ;
        RECT 25.200 128.300 26.000 128.400 ;
        RECT 1.200 127.700 26.000 128.300 ;
        RECT 1.200 127.600 2.000 127.700 ;
        RECT 25.200 127.600 26.000 127.700 ;
        RECT 63.600 128.300 64.400 128.400 ;
        RECT 89.200 128.300 90.000 128.400 ;
        RECT 97.200 128.300 98.000 128.400 ;
        RECT 63.600 127.700 98.000 128.300 ;
        RECT 63.600 127.600 64.400 127.700 ;
        RECT 89.200 127.600 90.000 127.700 ;
        RECT 97.200 127.600 98.000 127.700 ;
        RECT 118.000 128.300 118.800 128.400 ;
        RECT 127.600 128.300 128.400 128.400 ;
        RECT 118.000 127.700 128.400 128.300 ;
        RECT 118.000 127.600 118.800 127.700 ;
        RECT 127.600 127.600 128.400 127.700 ;
        RECT 210.800 128.300 211.600 128.400 ;
        RECT 246.000 128.300 246.800 128.400 ;
        RECT 210.800 127.700 246.800 128.300 ;
        RECT 210.800 127.600 211.600 127.700 ;
        RECT 246.000 127.600 246.800 127.700 ;
        RECT 252.400 128.300 253.200 128.400 ;
        RECT 311.600 128.300 312.400 128.400 ;
        RECT 252.400 127.700 312.400 128.300 ;
        RECT 252.400 127.600 253.200 127.700 ;
        RECT 311.600 127.600 312.400 127.700 ;
        RECT 345.200 127.600 346.000 128.400 ;
        RECT 356.400 128.300 357.200 128.400 ;
        RECT 358.000 128.300 358.800 128.400 ;
        RECT 356.400 127.700 358.800 128.300 ;
        RECT 356.400 127.600 357.200 127.700 ;
        RECT 358.000 127.600 358.800 127.700 ;
        RECT 366.000 128.300 366.800 128.400 ;
        RECT 393.200 128.300 394.000 128.400 ;
        RECT 366.000 127.700 394.000 128.300 ;
        RECT 366.000 127.600 366.800 127.700 ;
        RECT 393.200 127.600 394.000 127.700 ;
        RECT 396.400 128.300 397.200 128.400 ;
        RECT 407.600 128.300 408.400 128.400 ;
        RECT 434.800 128.300 435.600 128.400 ;
        RECT 396.400 127.700 435.600 128.300 ;
        RECT 396.400 127.600 397.200 127.700 ;
        RECT 407.600 127.600 408.400 127.700 ;
        RECT 434.800 127.600 435.600 127.700 ;
        RECT 436.400 128.300 437.200 128.400 ;
        RECT 476.400 128.300 477.200 128.400 ;
        RECT 436.400 127.700 477.200 128.300 ;
        RECT 436.400 127.600 437.200 127.700 ;
        RECT 476.400 127.600 477.200 127.700 ;
        RECT 511.600 128.300 512.400 128.400 ;
        RECT 516.400 128.300 517.200 128.400 ;
        RECT 538.800 128.300 539.600 128.400 ;
        RECT 511.600 127.700 539.600 128.300 ;
        RECT 511.600 127.600 512.400 127.700 ;
        RECT 516.400 127.600 517.200 127.700 ;
        RECT 538.800 127.600 539.600 127.700 ;
        RECT 14.000 126.300 14.800 126.400 ;
        RECT 22.000 126.300 22.800 126.400 ;
        RECT 14.000 125.700 22.800 126.300 ;
        RECT 14.000 125.600 14.800 125.700 ;
        RECT 22.000 125.600 22.800 125.700 ;
        RECT 95.600 126.300 96.400 126.400 ;
        RECT 111.600 126.300 112.400 126.400 ;
        RECT 95.600 125.700 112.400 126.300 ;
        RECT 95.600 125.600 96.400 125.700 ;
        RECT 111.600 125.600 112.400 125.700 ;
        RECT 306.800 125.600 307.600 126.400 ;
        RECT 332.400 126.300 333.200 126.400 ;
        RECT 418.800 126.300 419.600 126.400 ;
        RECT 332.400 125.700 419.600 126.300 ;
        RECT 332.400 125.600 333.200 125.700 ;
        RECT 418.800 125.600 419.600 125.700 ;
        RECT 87.600 124.300 88.400 124.400 ;
        RECT 114.800 124.300 115.600 124.400 ;
        RECT 87.600 123.700 115.600 124.300 ;
        RECT 87.600 123.600 88.400 123.700 ;
        RECT 114.800 123.600 115.600 123.700 ;
        RECT 302.000 124.300 302.800 124.400 ;
        RECT 313.200 124.300 314.000 124.400 ;
        RECT 302.000 123.700 314.000 124.300 ;
        RECT 302.000 123.600 302.800 123.700 ;
        RECT 313.200 123.600 314.000 123.700 ;
        RECT 532.400 124.300 533.200 124.400 ;
        RECT 540.400 124.300 541.200 124.400 ;
        RECT 548.400 124.300 549.200 124.400 ;
        RECT 532.400 123.700 549.200 124.300 ;
        RECT 532.400 123.600 533.200 123.700 ;
        RECT 540.400 123.600 541.200 123.700 ;
        RECT 548.400 123.600 549.200 123.700 ;
        RECT 102.000 122.300 102.800 122.400 ;
        RECT 105.200 122.300 106.000 122.400 ;
        RECT 102.000 121.700 106.000 122.300 ;
        RECT 102.000 121.600 102.800 121.700 ;
        RECT 105.200 121.600 106.000 121.700 ;
        RECT 214.000 122.300 214.800 122.400 ;
        RECT 226.800 122.300 227.600 122.400 ;
        RECT 214.000 121.700 227.600 122.300 ;
        RECT 214.000 121.600 214.800 121.700 ;
        RECT 226.800 121.600 227.600 121.700 ;
        RECT 250.800 122.300 251.600 122.400 ;
        RECT 270.000 122.300 270.800 122.400 ;
        RECT 274.800 122.300 275.600 122.400 ;
        RECT 310.000 122.300 310.800 122.400 ;
        RECT 250.800 121.700 310.800 122.300 ;
        RECT 250.800 121.600 251.600 121.700 ;
        RECT 270.000 121.600 270.800 121.700 ;
        RECT 274.800 121.600 275.600 121.700 ;
        RECT 310.000 121.600 310.800 121.700 ;
        RECT 70.000 120.300 70.800 120.400 ;
        RECT 73.200 120.300 74.000 120.400 ;
        RECT 102.000 120.300 102.800 120.400 ;
        RECT 70.000 119.700 102.800 120.300 ;
        RECT 70.000 119.600 70.800 119.700 ;
        RECT 73.200 119.600 74.000 119.700 ;
        RECT 102.000 119.600 102.800 119.700 ;
        RECT 177.200 120.300 178.000 120.400 ;
        RECT 274.800 120.300 275.600 120.400 ;
        RECT 276.400 120.300 277.200 120.400 ;
        RECT 177.200 119.700 277.200 120.300 ;
        RECT 177.200 119.600 178.000 119.700 ;
        RECT 274.800 119.600 275.600 119.700 ;
        RECT 276.400 119.600 277.200 119.700 ;
        RECT 399.600 120.300 400.400 120.400 ;
        RECT 406.000 120.300 406.800 120.400 ;
        RECT 399.600 119.700 406.800 120.300 ;
        RECT 399.600 119.600 400.400 119.700 ;
        RECT 406.000 119.600 406.800 119.700 ;
        RECT 431.600 120.300 432.400 120.400 ;
        RECT 433.200 120.300 434.000 120.400 ;
        RECT 431.600 119.700 434.000 120.300 ;
        RECT 431.600 119.600 432.400 119.700 ;
        RECT 433.200 119.600 434.000 119.700 ;
        RECT 47.600 118.300 48.400 118.400 ;
        RECT 50.800 118.300 51.600 118.400 ;
        RECT 47.600 117.700 51.600 118.300 ;
        RECT 47.600 117.600 48.400 117.700 ;
        RECT 50.800 117.600 51.600 117.700 ;
        RECT 52.400 118.300 53.200 118.400 ;
        RECT 82.800 118.300 83.600 118.400 ;
        RECT 52.400 117.700 83.600 118.300 ;
        RECT 52.400 117.600 53.200 117.700 ;
        RECT 82.800 117.600 83.600 117.700 ;
        RECT 114.800 118.300 115.600 118.400 ;
        RECT 130.800 118.300 131.600 118.400 ;
        RECT 151.600 118.300 152.400 118.400 ;
        RECT 114.800 117.700 152.400 118.300 ;
        RECT 114.800 117.600 115.600 117.700 ;
        RECT 130.800 117.600 131.600 117.700 ;
        RECT 151.600 117.600 152.400 117.700 ;
        RECT 201.200 118.300 202.000 118.400 ;
        RECT 207.600 118.300 208.400 118.400 ;
        RECT 201.200 117.700 208.400 118.300 ;
        RECT 201.200 117.600 202.000 117.700 ;
        RECT 207.600 117.600 208.400 117.700 ;
        RECT 223.600 118.300 224.400 118.400 ;
        RECT 226.800 118.300 227.600 118.400 ;
        RECT 223.600 117.700 227.600 118.300 ;
        RECT 223.600 117.600 224.400 117.700 ;
        RECT 226.800 117.600 227.600 117.700 ;
        RECT 228.400 118.300 229.200 118.400 ;
        RECT 265.200 118.300 266.000 118.400 ;
        RECT 228.400 117.700 266.000 118.300 ;
        RECT 228.400 117.600 229.200 117.700 ;
        RECT 265.200 117.600 266.000 117.700 ;
        RECT 380.400 118.300 381.200 118.400 ;
        RECT 431.600 118.300 432.400 118.400 ;
        RECT 380.400 117.700 432.400 118.300 ;
        RECT 380.400 117.600 381.200 117.700 ;
        RECT 431.600 117.600 432.400 117.700 ;
        RECT 449.200 118.300 450.000 118.400 ;
        RECT 454.000 118.300 454.800 118.400 ;
        RECT 449.200 117.700 454.800 118.300 ;
        RECT 449.200 117.600 450.000 117.700 ;
        RECT 454.000 117.600 454.800 117.700 ;
        RECT 508.400 118.300 509.200 118.400 ;
        RECT 513.200 118.300 514.000 118.400 ;
        RECT 567.600 118.300 568.400 118.400 ;
        RECT 508.400 117.700 568.400 118.300 ;
        RECT 508.400 117.600 509.200 117.700 ;
        RECT 513.200 117.600 514.000 117.700 ;
        RECT 567.600 117.600 568.400 117.700 ;
        RECT 578.800 118.300 579.600 118.400 ;
        RECT 582.000 118.300 582.800 118.400 ;
        RECT 578.800 117.700 582.800 118.300 ;
        RECT 578.800 117.600 579.600 117.700 ;
        RECT 582.000 117.600 582.800 117.700 ;
        RECT 12.400 116.300 13.200 116.400 ;
        RECT 54.000 116.300 54.800 116.400 ;
        RECT 12.400 115.700 54.800 116.300 ;
        RECT 12.400 115.600 13.200 115.700 ;
        RECT 54.000 115.600 54.800 115.700 ;
        RECT 108.400 116.300 109.200 116.400 ;
        RECT 137.200 116.300 138.000 116.400 ;
        RECT 108.400 115.700 138.000 116.300 ;
        RECT 108.400 115.600 109.200 115.700 ;
        RECT 137.200 115.600 138.000 115.700 ;
        RECT 209.200 116.300 210.000 116.400 ;
        RECT 212.400 116.300 213.200 116.400 ;
        RECT 273.200 116.300 274.000 116.400 ;
        RECT 209.200 115.700 274.000 116.300 ;
        RECT 209.200 115.600 210.000 115.700 ;
        RECT 212.400 115.600 213.200 115.700 ;
        RECT 273.200 115.600 274.000 115.700 ;
        RECT 414.000 116.300 414.800 116.400 ;
        RECT 417.200 116.300 418.000 116.400 ;
        RECT 414.000 115.700 418.000 116.300 ;
        RECT 414.000 115.600 414.800 115.700 ;
        RECT 417.200 115.600 418.000 115.700 ;
        RECT 431.600 116.300 432.400 116.400 ;
        RECT 479.600 116.300 480.400 116.400 ;
        RECT 431.600 115.700 480.400 116.300 ;
        RECT 431.600 115.600 432.400 115.700 ;
        RECT 479.600 115.600 480.400 115.700 ;
        RECT 527.600 116.300 528.400 116.400 ;
        RECT 537.200 116.300 538.000 116.400 ;
        RECT 527.600 115.700 538.000 116.300 ;
        RECT 527.600 115.600 528.400 115.700 ;
        RECT 537.200 115.600 538.000 115.700 ;
        RECT 41.200 114.300 42.000 114.400 ;
        RECT 65.200 114.300 66.000 114.400 ;
        RECT 41.200 113.700 66.000 114.300 ;
        RECT 41.200 113.600 42.000 113.700 ;
        RECT 65.200 113.600 66.000 113.700 ;
        RECT 78.000 114.300 78.800 114.400 ;
        RECT 169.200 114.300 170.000 114.400 ;
        RECT 78.000 113.700 170.000 114.300 ;
        RECT 78.000 113.600 78.800 113.700 ;
        RECT 169.200 113.600 170.000 113.700 ;
        RECT 182.000 114.300 182.800 114.400 ;
        RECT 262.000 114.300 262.800 114.400 ;
        RECT 182.000 113.700 262.800 114.300 ;
        RECT 182.000 113.600 182.800 113.700 ;
        RECT 262.000 113.600 262.800 113.700 ;
        RECT 289.200 114.300 290.000 114.400 ;
        RECT 332.400 114.300 333.200 114.400 ;
        RECT 289.200 113.700 333.200 114.300 ;
        RECT 289.200 113.600 290.000 113.700 ;
        RECT 332.400 113.600 333.200 113.700 ;
        RECT 362.800 114.300 363.600 114.400 ;
        RECT 388.400 114.300 389.200 114.400 ;
        RECT 394.800 114.300 395.600 114.400 ;
        RECT 406.000 114.300 406.800 114.400 ;
        RECT 362.800 113.700 406.800 114.300 ;
        RECT 362.800 113.600 363.600 113.700 ;
        RECT 388.400 113.600 389.200 113.700 ;
        RECT 394.800 113.600 395.600 113.700 ;
        RECT 406.000 113.600 406.800 113.700 ;
        RECT 473.200 114.300 474.000 114.400 ;
        RECT 476.400 114.300 477.200 114.400 ;
        RECT 473.200 113.700 477.200 114.300 ;
        RECT 473.200 113.600 474.000 113.700 ;
        RECT 476.400 113.600 477.200 113.700 ;
        RECT 534.000 114.300 534.800 114.400 ;
        RECT 545.200 114.300 546.000 114.400 ;
        RECT 534.000 113.700 546.000 114.300 ;
        RECT 534.000 113.600 534.800 113.700 ;
        RECT 545.200 113.600 546.000 113.700 ;
        RECT 6.000 112.300 6.800 112.400 ;
        RECT 10.800 112.300 11.600 112.400 ;
        RECT 6.000 111.700 11.600 112.300 ;
        RECT 6.000 111.600 6.800 111.700 ;
        RECT 10.800 111.600 11.600 111.700 ;
        RECT 36.400 112.300 37.200 112.400 ;
        RECT 49.200 112.300 50.000 112.400 ;
        RECT 36.400 111.700 50.000 112.300 ;
        RECT 36.400 111.600 37.200 111.700 ;
        RECT 49.200 111.600 50.000 111.700 ;
        RECT 74.800 112.300 75.600 112.400 ;
        RECT 76.400 112.300 77.200 112.400 ;
        RECT 74.800 111.700 77.200 112.300 ;
        RECT 74.800 111.600 75.600 111.700 ;
        RECT 76.400 111.600 77.200 111.700 ;
        RECT 84.400 112.300 85.200 112.400 ;
        RECT 89.200 112.300 90.000 112.400 ;
        RECT 92.400 112.300 93.200 112.400 ;
        RECT 97.200 112.300 98.000 112.400 ;
        RECT 111.600 112.300 112.400 112.400 ;
        RECT 84.400 111.700 98.000 112.300 ;
        RECT 84.400 111.600 85.200 111.700 ;
        RECT 89.200 111.600 90.000 111.700 ;
        RECT 92.400 111.600 93.200 111.700 ;
        RECT 97.200 111.600 98.000 111.700 ;
        RECT 98.900 111.700 112.400 112.300 ;
        RECT 98.900 110.400 99.500 111.700 ;
        RECT 111.600 111.600 112.400 111.700 ;
        RECT 121.200 112.300 122.000 112.400 ;
        RECT 134.000 112.300 134.800 112.400 ;
        RECT 121.200 111.700 134.800 112.300 ;
        RECT 121.200 111.600 122.000 111.700 ;
        RECT 134.000 111.600 134.800 111.700 ;
        RECT 193.200 112.300 194.000 112.400 ;
        RECT 196.400 112.300 197.200 112.400 ;
        RECT 193.200 111.700 197.200 112.300 ;
        RECT 193.200 111.600 194.000 111.700 ;
        RECT 196.400 111.600 197.200 111.700 ;
        RECT 204.400 112.300 205.200 112.400 ;
        RECT 207.600 112.300 208.400 112.400 ;
        RECT 204.400 111.700 208.400 112.300 ;
        RECT 204.400 111.600 205.200 111.700 ;
        RECT 207.600 111.600 208.400 111.700 ;
        RECT 217.200 112.300 218.000 112.400 ;
        RECT 242.800 112.300 243.600 112.400 ;
        RECT 217.200 111.700 243.600 112.300 ;
        RECT 217.200 111.600 218.000 111.700 ;
        RECT 242.800 111.600 243.600 111.700 ;
        RECT 265.200 112.300 266.000 112.400 ;
        RECT 278.000 112.300 278.800 112.400 ;
        RECT 265.200 111.700 278.800 112.300 ;
        RECT 265.200 111.600 266.000 111.700 ;
        RECT 278.000 111.600 278.800 111.700 ;
        RECT 367.600 111.600 368.400 112.400 ;
        RECT 370.800 112.300 371.600 112.400 ;
        RECT 390.000 112.300 390.800 112.400 ;
        RECT 370.800 111.700 390.800 112.300 ;
        RECT 370.800 111.600 371.600 111.700 ;
        RECT 390.000 111.600 390.800 111.700 ;
        RECT 407.600 112.300 408.400 112.400 ;
        RECT 412.400 112.300 413.200 112.400 ;
        RECT 407.600 111.700 413.200 112.300 ;
        RECT 407.600 111.600 408.400 111.700 ;
        RECT 412.400 111.600 413.200 111.700 ;
        RECT 458.800 112.300 459.600 112.400 ;
        RECT 460.400 112.300 461.200 112.400 ;
        RECT 458.800 111.700 461.200 112.300 ;
        RECT 458.800 111.600 459.600 111.700 ;
        RECT 460.400 111.600 461.200 111.700 ;
        RECT 486.000 112.300 486.800 112.400 ;
        RECT 529.200 112.300 530.000 112.400 ;
        RECT 486.000 111.700 530.000 112.300 ;
        RECT 486.000 111.600 486.800 111.700 ;
        RECT 529.200 111.600 530.000 111.700 ;
        RECT 562.800 112.300 563.600 112.400 ;
        RECT 569.200 112.300 570.000 112.400 ;
        RECT 562.800 111.700 570.000 112.300 ;
        RECT 562.800 111.600 563.600 111.700 ;
        RECT 569.200 111.600 570.000 111.700 ;
        RECT 1.200 110.300 2.000 110.400 ;
        RECT 7.600 110.300 8.400 110.400 ;
        RECT 1.200 109.700 8.400 110.300 ;
        RECT 1.200 109.600 2.000 109.700 ;
        RECT 7.600 109.600 8.400 109.700 ;
        RECT 33.200 110.300 34.000 110.400 ;
        RECT 38.000 110.300 38.800 110.400 ;
        RECT 33.200 109.700 38.800 110.300 ;
        RECT 33.200 109.600 34.000 109.700 ;
        RECT 38.000 109.600 38.800 109.700 ;
        RECT 44.400 110.300 45.200 110.400 ;
        RECT 50.800 110.300 51.600 110.400 ;
        RECT 63.600 110.300 64.400 110.400 ;
        RECT 44.400 109.700 49.900 110.300 ;
        RECT 44.400 109.600 45.200 109.700 ;
        RECT 2.800 108.300 3.600 108.400 ;
        RECT 22.000 108.300 22.800 108.400 ;
        RECT 2.800 107.700 22.800 108.300 ;
        RECT 2.800 107.600 3.600 107.700 ;
        RECT 22.000 107.600 22.800 107.700 ;
        RECT 33.200 108.300 34.000 108.400 ;
        RECT 36.400 108.300 37.200 108.400 ;
        RECT 41.200 108.300 42.000 108.400 ;
        RECT 33.200 107.700 42.000 108.300 ;
        RECT 33.200 107.600 34.000 107.700 ;
        RECT 36.400 107.600 37.200 107.700 ;
        RECT 41.200 107.600 42.000 107.700 ;
        RECT 42.800 108.300 43.600 108.400 ;
        RECT 47.600 108.300 48.400 108.400 ;
        RECT 42.800 107.700 48.400 108.300 ;
        RECT 49.300 108.300 49.900 109.700 ;
        RECT 50.800 109.700 64.400 110.300 ;
        RECT 50.800 109.600 51.600 109.700 ;
        RECT 63.600 109.600 64.400 109.700 ;
        RECT 89.200 110.300 90.000 110.400 ;
        RECT 98.800 110.300 99.600 110.400 ;
        RECT 89.200 109.700 99.600 110.300 ;
        RECT 89.200 109.600 90.000 109.700 ;
        RECT 98.800 109.600 99.600 109.700 ;
        RECT 105.200 110.300 106.000 110.400 ;
        RECT 108.400 110.300 109.200 110.400 ;
        RECT 105.200 109.700 109.200 110.300 ;
        RECT 105.200 109.600 106.000 109.700 ;
        RECT 108.400 109.600 109.200 109.700 ;
        RECT 127.600 110.300 128.400 110.400 ;
        RECT 148.400 110.300 149.200 110.400 ;
        RECT 156.400 110.300 157.200 110.400 ;
        RECT 127.600 109.700 157.200 110.300 ;
        RECT 127.600 109.600 128.400 109.700 ;
        RECT 148.400 109.600 149.200 109.700 ;
        RECT 156.400 109.600 157.200 109.700 ;
        RECT 191.600 110.300 192.400 110.400 ;
        RECT 210.800 110.300 211.600 110.400 ;
        RECT 191.600 109.700 211.600 110.300 ;
        RECT 191.600 109.600 192.400 109.700 ;
        RECT 210.800 109.600 211.600 109.700 ;
        RECT 223.600 110.300 224.400 110.400 ;
        RECT 241.200 110.300 242.000 110.400 ;
        RECT 268.400 110.300 269.200 110.400 ;
        RECT 223.600 109.700 269.200 110.300 ;
        RECT 223.600 109.600 224.400 109.700 ;
        RECT 241.200 109.600 242.000 109.700 ;
        RECT 268.400 109.600 269.200 109.700 ;
        RECT 274.800 110.300 275.600 110.400 ;
        RECT 282.800 110.300 283.600 110.400 ;
        RECT 297.200 110.300 298.000 110.400 ;
        RECT 274.800 109.700 298.000 110.300 ;
        RECT 274.800 109.600 275.600 109.700 ;
        RECT 282.800 109.600 283.600 109.700 ;
        RECT 297.200 109.600 298.000 109.700 ;
        RECT 351.600 110.300 352.400 110.400 ;
        RECT 359.600 110.300 360.400 110.400 ;
        RECT 351.600 109.700 360.400 110.300 ;
        RECT 351.600 109.600 352.400 109.700 ;
        RECT 359.600 109.600 360.400 109.700 ;
        RECT 375.600 110.300 376.400 110.400 ;
        RECT 409.200 110.300 410.000 110.400 ;
        RECT 375.600 109.700 410.000 110.300 ;
        RECT 375.600 109.600 376.400 109.700 ;
        RECT 409.200 109.600 410.000 109.700 ;
        RECT 412.400 110.300 413.200 110.400 ;
        RECT 417.200 110.300 418.000 110.400 ;
        RECT 412.400 109.700 418.000 110.300 ;
        RECT 412.400 109.600 413.200 109.700 ;
        RECT 417.200 109.600 418.000 109.700 ;
        RECT 423.600 110.300 424.400 110.400 ;
        RECT 436.400 110.300 437.200 110.400 ;
        RECT 423.600 109.700 437.200 110.300 ;
        RECT 423.600 109.600 424.400 109.700 ;
        RECT 436.400 109.600 437.200 109.700 ;
        RECT 438.000 110.300 438.800 110.400 ;
        RECT 462.000 110.300 462.800 110.400 ;
        RECT 438.000 109.700 462.800 110.300 ;
        RECT 438.000 109.600 438.800 109.700 ;
        RECT 462.000 109.600 462.800 109.700 ;
        RECT 473.200 110.300 474.000 110.400 ;
        RECT 508.400 110.300 509.200 110.400 ;
        RECT 473.200 109.700 509.200 110.300 ;
        RECT 473.200 109.600 474.000 109.700 ;
        RECT 508.400 109.600 509.200 109.700 ;
        RECT 521.200 110.300 522.000 110.400 ;
        RECT 527.600 110.300 528.400 110.400 ;
        RECT 521.200 109.700 528.400 110.300 ;
        RECT 521.200 109.600 522.000 109.700 ;
        RECT 527.600 109.600 528.400 109.700 ;
        RECT 551.600 110.300 552.400 110.400 ;
        RECT 559.600 110.300 560.400 110.400 ;
        RECT 551.600 109.700 560.400 110.300 ;
        RECT 551.600 109.600 552.400 109.700 ;
        RECT 559.600 109.600 560.400 109.700 ;
        RECT 54.000 108.300 54.800 108.400 ;
        RECT 65.200 108.300 66.000 108.400 ;
        RECT 68.400 108.300 69.200 108.400 ;
        RECT 49.300 107.700 64.300 108.300 ;
        RECT 42.800 107.600 43.600 107.700 ;
        RECT 47.600 107.600 48.400 107.700 ;
        RECT 54.000 107.600 54.800 107.700 ;
        RECT 6.000 106.300 6.800 106.400 ;
        RECT 15.600 106.300 16.400 106.400 ;
        RECT 6.000 105.700 16.400 106.300 ;
        RECT 6.000 105.600 6.800 105.700 ;
        RECT 15.600 105.600 16.400 105.700 ;
        RECT 34.800 106.300 35.600 106.400 ;
        RECT 60.400 106.300 61.200 106.400 ;
        RECT 34.800 105.700 61.200 106.300 ;
        RECT 63.700 106.300 64.300 107.700 ;
        RECT 65.200 107.700 69.200 108.300 ;
        RECT 65.200 107.600 66.000 107.700 ;
        RECT 68.400 107.600 69.200 107.700 ;
        RECT 71.600 108.300 72.400 108.400 ;
        RECT 81.200 108.300 82.000 108.400 ;
        RECT 71.600 107.700 82.000 108.300 ;
        RECT 71.600 107.600 72.400 107.700 ;
        RECT 81.200 107.600 82.000 107.700 ;
        RECT 87.600 108.300 88.400 108.400 ;
        RECT 103.600 108.300 104.400 108.400 ;
        RECT 127.600 108.300 128.400 108.400 ;
        RECT 87.600 107.700 128.400 108.300 ;
        RECT 87.600 107.600 88.400 107.700 ;
        RECT 103.600 107.600 104.400 107.700 ;
        RECT 127.600 107.600 128.400 107.700 ;
        RECT 194.800 108.300 195.600 108.400 ;
        RECT 201.200 108.300 202.000 108.400 ;
        RECT 194.800 107.700 202.000 108.300 ;
        RECT 194.800 107.600 195.600 107.700 ;
        RECT 201.200 107.600 202.000 107.700 ;
        RECT 204.400 108.300 205.200 108.400 ;
        RECT 209.200 108.300 210.000 108.400 ;
        RECT 223.600 108.300 224.400 108.400 ;
        RECT 204.400 107.700 224.400 108.300 ;
        RECT 204.400 107.600 205.200 107.700 ;
        RECT 209.200 107.600 210.000 107.700 ;
        RECT 223.600 107.600 224.400 107.700 ;
        RECT 225.200 108.300 226.000 108.400 ;
        RECT 233.200 108.300 234.000 108.400 ;
        RECT 225.200 107.700 234.000 108.300 ;
        RECT 225.200 107.600 226.000 107.700 ;
        RECT 233.200 107.600 234.000 107.700 ;
        RECT 239.600 108.300 240.400 108.400 ;
        RECT 255.600 108.300 256.400 108.400 ;
        RECT 239.600 107.700 256.400 108.300 ;
        RECT 239.600 107.600 240.400 107.700 ;
        RECT 255.600 107.600 256.400 107.700 ;
        RECT 263.600 108.300 264.400 108.400 ;
        RECT 271.600 108.300 272.400 108.400 ;
        RECT 276.400 108.300 277.200 108.400 ;
        RECT 263.600 107.700 277.200 108.300 ;
        RECT 263.600 107.600 264.400 107.700 ;
        RECT 271.600 107.600 272.400 107.700 ;
        RECT 276.400 107.600 277.200 107.700 ;
        RECT 314.800 108.300 315.600 108.400 ;
        RECT 329.200 108.300 330.000 108.400 ;
        RECT 314.800 107.700 330.000 108.300 ;
        RECT 314.800 107.600 315.600 107.700 ;
        RECT 329.200 107.600 330.000 107.700 ;
        RECT 366.000 108.300 366.800 108.400 ;
        RECT 386.800 108.300 387.600 108.400 ;
        RECT 396.400 108.300 397.200 108.400 ;
        RECT 366.000 107.700 397.200 108.300 ;
        RECT 366.000 107.600 366.800 107.700 ;
        RECT 386.800 107.600 387.600 107.700 ;
        RECT 396.400 107.600 397.200 107.700 ;
        RECT 410.800 108.300 411.600 108.400 ;
        RECT 414.000 108.300 414.800 108.400 ;
        RECT 410.800 107.700 414.800 108.300 ;
        RECT 410.800 107.600 411.600 107.700 ;
        RECT 414.000 107.600 414.800 107.700 ;
        RECT 543.600 108.300 544.400 108.400 ;
        RECT 546.800 108.300 547.600 108.400 ;
        RECT 550.000 108.300 550.800 108.400 ;
        RECT 543.600 107.700 550.800 108.300 ;
        RECT 543.600 107.600 544.400 107.700 ;
        RECT 546.800 107.600 547.600 107.700 ;
        RECT 550.000 107.600 550.800 107.700 ;
        RECT 554.800 108.300 555.600 108.400 ;
        RECT 562.800 108.300 563.600 108.400 ;
        RECT 566.000 108.300 566.800 108.400 ;
        RECT 554.800 107.700 566.800 108.300 ;
        RECT 554.800 107.600 555.600 107.700 ;
        RECT 562.800 107.600 563.600 107.700 ;
        RECT 566.000 107.600 566.800 107.700 ;
        RECT 65.200 106.300 66.000 106.400 ;
        RECT 63.700 105.700 66.000 106.300 ;
        RECT 34.800 105.600 35.600 105.700 ;
        RECT 60.400 105.600 61.200 105.700 ;
        RECT 65.200 105.600 66.000 105.700 ;
        RECT 82.800 106.300 83.600 106.400 ;
        RECT 89.200 106.300 90.000 106.400 ;
        RECT 92.400 106.300 93.200 106.400 ;
        RECT 94.000 106.300 94.800 106.400 ;
        RECT 82.800 105.700 94.800 106.300 ;
        RECT 82.800 105.600 83.600 105.700 ;
        RECT 89.200 105.600 90.000 105.700 ;
        RECT 92.400 105.600 93.200 105.700 ;
        RECT 94.000 105.600 94.800 105.700 ;
        RECT 98.800 106.300 99.600 106.400 ;
        RECT 102.000 106.300 102.800 106.400 ;
        RECT 110.000 106.300 110.800 106.400 ;
        RECT 98.800 105.700 110.800 106.300 ;
        RECT 98.800 105.600 99.600 105.700 ;
        RECT 102.000 105.600 102.800 105.700 ;
        RECT 110.000 105.600 110.800 105.700 ;
        RECT 135.600 106.300 136.400 106.400 ;
        RECT 143.600 106.300 144.400 106.400 ;
        RECT 135.600 105.700 144.400 106.300 ;
        RECT 135.600 105.600 136.400 105.700 ;
        RECT 143.600 105.600 144.400 105.700 ;
        RECT 145.200 106.300 146.000 106.400 ;
        RECT 150.000 106.300 150.800 106.400 ;
        RECT 145.200 105.700 150.800 106.300 ;
        RECT 145.200 105.600 146.000 105.700 ;
        RECT 150.000 105.600 150.800 105.700 ;
        RECT 159.600 106.300 160.400 106.400 ;
        RECT 162.800 106.300 163.600 106.400 ;
        RECT 159.600 105.700 163.600 106.300 ;
        RECT 159.600 105.600 160.400 105.700 ;
        RECT 162.800 105.600 163.600 105.700 ;
        RECT 223.600 106.300 224.400 106.400 ;
        RECT 230.000 106.300 230.800 106.400 ;
        RECT 223.600 105.700 230.800 106.300 ;
        RECT 223.600 105.600 224.400 105.700 ;
        RECT 230.000 105.600 230.800 105.700 ;
        RECT 273.200 106.300 274.000 106.400 ;
        RECT 281.200 106.300 282.000 106.400 ;
        RECT 273.200 105.700 282.000 106.300 ;
        RECT 273.200 105.600 274.000 105.700 ;
        RECT 281.200 105.600 282.000 105.700 ;
        RECT 378.800 106.300 379.600 106.400 ;
        RECT 382.000 106.300 382.800 106.400 ;
        RECT 378.800 105.700 382.800 106.300 ;
        RECT 378.800 105.600 379.600 105.700 ;
        RECT 382.000 105.600 382.800 105.700 ;
        RECT 409.200 106.300 410.000 106.400 ;
        RECT 430.000 106.300 430.800 106.400 ;
        RECT 409.200 105.700 430.800 106.300 ;
        RECT 409.200 105.600 410.000 105.700 ;
        RECT 430.000 105.600 430.800 105.700 ;
        RECT 462.000 106.300 462.800 106.400 ;
        RECT 478.000 106.300 478.800 106.400 ;
        RECT 462.000 105.700 478.800 106.300 ;
        RECT 462.000 105.600 462.800 105.700 ;
        RECT 478.000 105.600 478.800 105.700 ;
        RECT 28.400 104.300 29.200 104.400 ;
        RECT 33.200 104.300 34.000 104.400 ;
        RECT 28.400 103.700 34.000 104.300 ;
        RECT 28.400 103.600 29.200 103.700 ;
        RECT 33.200 103.600 34.000 103.700 ;
        RECT 102.000 104.300 102.800 104.400 ;
        RECT 105.200 104.300 106.000 104.400 ;
        RECT 102.000 103.700 106.000 104.300 ;
        RECT 102.000 103.600 102.800 103.700 ;
        RECT 105.200 103.600 106.000 103.700 ;
        RECT 201.200 104.300 202.000 104.400 ;
        RECT 218.800 104.300 219.600 104.400 ;
        RECT 234.800 104.300 235.600 104.400 ;
        RECT 242.800 104.300 243.600 104.400 ;
        RECT 257.200 104.300 258.000 104.400 ;
        RECT 201.200 103.700 258.000 104.300 ;
        RECT 201.200 103.600 202.000 103.700 ;
        RECT 218.800 103.600 219.600 103.700 ;
        RECT 234.800 103.600 235.600 103.700 ;
        RECT 242.800 103.600 243.600 103.700 ;
        RECT 257.200 103.600 258.000 103.700 ;
        RECT 258.800 104.300 259.600 104.400 ;
        RECT 282.800 104.300 283.600 104.400 ;
        RECT 292.400 104.300 293.200 104.400 ;
        RECT 258.800 103.700 283.600 104.300 ;
        RECT 258.800 103.600 259.600 103.700 ;
        RECT 282.800 103.600 283.600 103.700 ;
        RECT 286.100 103.700 293.200 104.300 ;
        RECT 2.800 102.300 3.600 102.400 ;
        RECT 9.200 102.300 10.000 102.400 ;
        RECT 18.800 102.300 19.600 102.400 ;
        RECT 2.800 101.700 19.600 102.300 ;
        RECT 2.800 101.600 3.600 101.700 ;
        RECT 9.200 101.600 10.000 101.700 ;
        RECT 18.800 101.600 19.600 101.700 ;
        RECT 22.000 102.300 22.800 102.400 ;
        RECT 46.000 102.300 46.800 102.400 ;
        RECT 22.000 101.700 46.800 102.300 ;
        RECT 22.000 101.600 22.800 101.700 ;
        RECT 46.000 101.600 46.800 101.700 ;
        RECT 86.000 102.300 86.800 102.400 ;
        RECT 146.800 102.300 147.600 102.400 ;
        RECT 86.000 101.700 147.600 102.300 ;
        RECT 86.000 101.600 86.800 101.700 ;
        RECT 146.800 101.600 147.600 101.700 ;
        RECT 220.400 102.300 221.200 102.400 ;
        RECT 260.400 102.300 261.200 102.400 ;
        RECT 220.400 101.700 261.200 102.300 ;
        RECT 220.400 101.600 221.200 101.700 ;
        RECT 260.400 101.600 261.200 101.700 ;
        RECT 265.200 102.300 266.000 102.400 ;
        RECT 286.100 102.300 286.700 103.700 ;
        RECT 292.400 103.600 293.200 103.700 ;
        RECT 356.400 104.300 357.200 104.400 ;
        RECT 382.000 104.300 382.800 104.400 ;
        RECT 356.400 103.700 382.800 104.300 ;
        RECT 356.400 103.600 357.200 103.700 ;
        RECT 382.000 103.600 382.800 103.700 ;
        RECT 417.200 104.300 418.000 104.400 ;
        RECT 466.800 104.300 467.600 104.400 ;
        RECT 481.200 104.300 482.000 104.400 ;
        RECT 535.600 104.300 536.400 104.400 ;
        RECT 417.200 103.700 536.400 104.300 ;
        RECT 417.200 103.600 418.000 103.700 ;
        RECT 466.800 103.600 467.600 103.700 ;
        RECT 481.200 103.600 482.000 103.700 ;
        RECT 535.600 103.600 536.400 103.700 ;
        RECT 540.400 104.300 541.200 104.400 ;
        RECT 546.800 104.300 547.600 104.400 ;
        RECT 540.400 103.700 547.600 104.300 ;
        RECT 540.400 103.600 541.200 103.700 ;
        RECT 546.800 103.600 547.600 103.700 ;
        RECT 265.200 101.700 286.700 102.300 ;
        RECT 265.200 101.600 266.000 101.700 ;
        RECT 287.600 101.600 288.400 102.400 ;
        RECT 326.000 102.300 326.800 102.400 ;
        RECT 356.400 102.300 357.200 102.400 ;
        RECT 326.000 101.700 357.200 102.300 ;
        RECT 326.000 101.600 326.800 101.700 ;
        RECT 356.400 101.600 357.200 101.700 ;
        RECT 378.800 102.300 379.600 102.400 ;
        RECT 396.400 102.300 397.200 102.400 ;
        RECT 398.000 102.300 398.800 102.400 ;
        RECT 406.000 102.300 406.800 102.400 ;
        RECT 378.800 101.700 406.800 102.300 ;
        RECT 378.800 101.600 379.600 101.700 ;
        RECT 396.400 101.600 397.200 101.700 ;
        RECT 398.000 101.600 398.800 101.700 ;
        RECT 406.000 101.600 406.800 101.700 ;
        RECT 462.000 102.300 462.800 102.400 ;
        RECT 489.200 102.300 490.000 102.400 ;
        RECT 462.000 101.700 490.000 102.300 ;
        RECT 462.000 101.600 462.800 101.700 ;
        RECT 489.200 101.600 490.000 101.700 ;
        RECT 529.200 102.300 530.000 102.400 ;
        RECT 537.200 102.300 538.000 102.400 ;
        RECT 529.200 101.700 538.000 102.300 ;
        RECT 529.200 101.600 530.000 101.700 ;
        RECT 537.200 101.600 538.000 101.700 ;
        RECT 577.200 102.300 578.000 102.400 ;
        RECT 583.600 102.300 584.400 102.400 ;
        RECT 577.200 101.700 584.400 102.300 ;
        RECT 577.200 101.600 578.000 101.700 ;
        RECT 583.600 101.600 584.400 101.700 ;
        RECT 2.800 100.300 3.600 100.400 ;
        RECT 14.000 100.300 14.800 100.400 ;
        RECT 2.800 99.700 14.800 100.300 ;
        RECT 2.800 99.600 3.600 99.700 ;
        RECT 14.000 99.600 14.800 99.700 ;
        RECT 114.800 100.300 115.600 100.400 ;
        RECT 124.400 100.300 125.200 100.400 ;
        RECT 114.800 99.700 125.200 100.300 ;
        RECT 114.800 99.600 115.600 99.700 ;
        RECT 124.400 99.600 125.200 99.700 ;
        RECT 196.400 100.300 197.200 100.400 ;
        RECT 212.400 100.300 213.200 100.400 ;
        RECT 220.400 100.300 221.200 100.400 ;
        RECT 196.400 99.700 221.200 100.300 ;
        RECT 196.400 99.600 197.200 99.700 ;
        RECT 212.400 99.600 213.200 99.700 ;
        RECT 220.400 99.600 221.200 99.700 ;
        RECT 382.000 100.300 382.800 100.400 ;
        RECT 452.400 100.300 453.200 100.400 ;
        RECT 458.800 100.300 459.600 100.400 ;
        RECT 466.800 100.300 467.600 100.400 ;
        RECT 382.000 99.700 467.600 100.300 ;
        RECT 382.000 99.600 382.800 99.700 ;
        RECT 452.400 99.600 453.200 99.700 ;
        RECT 458.800 99.600 459.600 99.700 ;
        RECT 466.800 99.600 467.600 99.700 ;
        RECT 479.600 99.600 480.400 100.400 ;
        RECT 100.400 98.300 101.200 98.400 ;
        RECT 102.000 98.300 102.800 98.400 ;
        RECT 100.400 97.700 102.800 98.300 ;
        RECT 100.400 97.600 101.200 97.700 ;
        RECT 102.000 97.600 102.800 97.700 ;
        RECT 105.200 98.300 106.000 98.400 ;
        RECT 134.000 98.300 134.800 98.400 ;
        RECT 145.200 98.300 146.000 98.400 ;
        RECT 105.200 97.700 146.000 98.300 ;
        RECT 105.200 97.600 106.000 97.700 ;
        RECT 134.000 97.600 134.800 97.700 ;
        RECT 145.200 97.600 146.000 97.700 ;
        RECT 183.600 98.300 184.400 98.400 ;
        RECT 190.000 98.300 190.800 98.400 ;
        RECT 196.400 98.300 197.200 98.400 ;
        RECT 202.800 98.300 203.600 98.400 ;
        RECT 217.200 98.300 218.000 98.400 ;
        RECT 218.800 98.300 219.600 98.400 ;
        RECT 183.600 97.700 219.600 98.300 ;
        RECT 183.600 97.600 184.400 97.700 ;
        RECT 190.000 97.600 190.800 97.700 ;
        RECT 196.400 97.600 197.200 97.700 ;
        RECT 202.800 97.600 203.600 97.700 ;
        RECT 217.200 97.600 218.000 97.700 ;
        RECT 218.800 97.600 219.600 97.700 ;
        RECT 230.000 98.300 230.800 98.400 ;
        RECT 233.200 98.300 234.000 98.400 ;
        RECT 230.000 97.700 234.000 98.300 ;
        RECT 230.000 97.600 230.800 97.700 ;
        RECT 233.200 97.600 234.000 97.700 ;
        RECT 268.400 98.300 269.200 98.400 ;
        RECT 274.800 98.300 275.600 98.400 ;
        RECT 303.600 98.300 304.400 98.400 ;
        RECT 268.400 97.700 304.400 98.300 ;
        RECT 268.400 97.600 269.200 97.700 ;
        RECT 274.800 97.600 275.600 97.700 ;
        RECT 303.600 97.600 304.400 97.700 ;
        RECT 366.000 98.300 366.800 98.400 ;
        RECT 388.400 98.300 389.200 98.400 ;
        RECT 394.800 98.300 395.600 98.400 ;
        RECT 366.000 97.700 395.600 98.300 ;
        RECT 366.000 97.600 366.800 97.700 ;
        RECT 388.400 97.600 389.200 97.700 ;
        RECT 394.800 97.600 395.600 97.700 ;
        RECT 423.600 98.300 424.400 98.400 ;
        RECT 463.600 98.300 464.400 98.400 ;
        RECT 468.400 98.300 469.200 98.400 ;
        RECT 423.600 97.700 469.200 98.300 ;
        RECT 423.600 97.600 424.400 97.700 ;
        RECT 463.600 97.600 464.400 97.700 ;
        RECT 468.400 97.600 469.200 97.700 ;
        RECT 476.400 98.300 477.200 98.400 ;
        RECT 478.000 98.300 478.800 98.400 ;
        RECT 476.400 97.700 478.800 98.300 ;
        RECT 476.400 97.600 477.200 97.700 ;
        RECT 478.000 97.600 478.800 97.700 ;
        RECT 52.400 96.300 53.200 96.400 ;
        RECT 57.200 96.300 58.000 96.400 ;
        RECT 52.400 95.700 58.000 96.300 ;
        RECT 52.400 95.600 53.200 95.700 ;
        RECT 57.200 95.600 58.000 95.700 ;
        RECT 58.800 96.300 59.600 96.400 ;
        RECT 73.200 96.300 74.000 96.400 ;
        RECT 58.800 95.700 74.000 96.300 ;
        RECT 58.800 95.600 59.600 95.700 ;
        RECT 73.200 95.600 74.000 95.700 ;
        RECT 94.000 96.300 94.800 96.400 ;
        RECT 98.800 96.300 99.600 96.400 ;
        RECT 94.000 95.700 99.600 96.300 ;
        RECT 94.000 95.600 94.800 95.700 ;
        RECT 98.800 95.600 99.600 95.700 ;
        RECT 100.400 96.300 101.200 96.400 ;
        RECT 108.400 96.300 109.200 96.400 ;
        RECT 100.400 95.700 109.200 96.300 ;
        RECT 100.400 95.600 101.200 95.700 ;
        RECT 108.400 95.600 109.200 95.700 ;
        RECT 121.200 96.300 122.000 96.400 ;
        RECT 130.800 96.300 131.600 96.400 ;
        RECT 121.200 95.700 131.600 96.300 ;
        RECT 121.200 95.600 122.000 95.700 ;
        RECT 130.800 95.600 131.600 95.700 ;
        RECT 175.600 96.300 176.400 96.400 ;
        RECT 180.400 96.300 181.200 96.400 ;
        RECT 183.600 96.300 184.400 96.400 ;
        RECT 175.600 95.700 184.400 96.300 ;
        RECT 175.600 95.600 176.400 95.700 ;
        RECT 180.400 95.600 181.200 95.700 ;
        RECT 183.600 95.600 184.400 95.700 ;
        RECT 186.800 96.300 187.600 96.400 ;
        RECT 246.000 96.300 246.800 96.400 ;
        RECT 186.800 95.700 246.800 96.300 ;
        RECT 186.800 95.600 187.600 95.700 ;
        RECT 246.000 95.600 246.800 95.700 ;
        RECT 278.000 96.300 278.800 96.400 ;
        RECT 282.800 96.300 283.600 96.400 ;
        RECT 300.400 96.300 301.200 96.400 ;
        RECT 329.200 96.300 330.000 96.400 ;
        RECT 278.000 95.700 330.000 96.300 ;
        RECT 278.000 95.600 278.800 95.700 ;
        RECT 282.800 95.600 283.600 95.700 ;
        RECT 300.400 95.600 301.200 95.700 ;
        RECT 329.200 95.600 330.000 95.700 ;
        RECT 356.400 96.300 357.200 96.400 ;
        RECT 378.800 96.300 379.600 96.400 ;
        RECT 356.400 95.700 379.600 96.300 ;
        RECT 356.400 95.600 357.200 95.700 ;
        RECT 378.800 95.600 379.600 95.700 ;
        RECT 385.200 96.300 386.000 96.400 ;
        RECT 390.000 96.300 390.800 96.400 ;
        RECT 409.200 96.300 410.000 96.400 ;
        RECT 385.200 95.700 410.000 96.300 ;
        RECT 385.200 95.600 386.000 95.700 ;
        RECT 390.000 95.600 390.800 95.700 ;
        RECT 409.200 95.600 410.000 95.700 ;
        RECT 426.800 96.300 427.600 96.400 ;
        RECT 465.200 96.300 466.000 96.400 ;
        RECT 426.800 95.700 466.000 96.300 ;
        RECT 426.800 95.600 427.600 95.700 ;
        RECT 465.200 95.600 466.000 95.700 ;
        RECT 473.200 96.300 474.000 96.400 ;
        RECT 479.600 96.300 480.400 96.400 ;
        RECT 473.200 95.700 480.400 96.300 ;
        RECT 473.200 95.600 474.000 95.700 ;
        RECT 479.600 95.600 480.400 95.700 ;
        RECT 26.800 94.300 27.600 94.400 ;
        RECT 34.800 94.300 35.600 94.400 ;
        RECT 38.000 94.300 38.800 94.400 ;
        RECT 26.800 93.700 38.800 94.300 ;
        RECT 26.800 93.600 27.600 93.700 ;
        RECT 34.800 93.600 35.600 93.700 ;
        RECT 38.000 93.600 38.800 93.700 ;
        RECT 41.200 94.300 42.000 94.400 ;
        RECT 60.400 94.300 61.200 94.400 ;
        RECT 41.200 93.700 61.200 94.300 ;
        RECT 41.200 93.600 42.000 93.700 ;
        RECT 60.400 93.600 61.200 93.700 ;
        RECT 63.600 93.600 64.400 94.400 ;
        RECT 65.200 94.300 66.000 94.400 ;
        RECT 70.000 94.300 70.800 94.400 ;
        RECT 65.200 93.700 70.800 94.300 ;
        RECT 65.200 93.600 66.000 93.700 ;
        RECT 70.000 93.600 70.800 93.700 ;
        RECT 84.400 94.300 85.200 94.400 ;
        RECT 89.200 94.300 90.000 94.400 ;
        RECT 84.400 93.700 90.000 94.300 ;
        RECT 84.400 93.600 85.200 93.700 ;
        RECT 89.200 93.600 90.000 93.700 ;
        RECT 90.800 94.300 91.600 94.400 ;
        RECT 97.200 94.300 98.000 94.400 ;
        RECT 122.800 94.300 123.600 94.400 ;
        RECT 140.400 94.300 141.200 94.400 ;
        RECT 90.800 93.700 141.200 94.300 ;
        RECT 90.800 93.600 91.600 93.700 ;
        RECT 97.200 93.600 98.000 93.700 ;
        RECT 122.800 93.600 123.600 93.700 ;
        RECT 140.400 93.600 141.200 93.700 ;
        RECT 143.600 94.300 144.400 94.400 ;
        RECT 162.800 94.300 163.600 94.400 ;
        RECT 143.600 93.700 163.600 94.300 ;
        RECT 143.600 93.600 144.400 93.700 ;
        RECT 162.800 93.600 163.600 93.700 ;
        RECT 194.800 94.300 195.600 94.400 ;
        RECT 201.200 94.300 202.000 94.400 ;
        RECT 194.800 93.700 202.000 94.300 ;
        RECT 194.800 93.600 195.600 93.700 ;
        RECT 201.200 93.600 202.000 93.700 ;
        RECT 202.800 94.300 203.600 94.400 ;
        RECT 207.600 94.300 208.400 94.400 ;
        RECT 202.800 93.700 208.400 94.300 ;
        RECT 202.800 93.600 203.600 93.700 ;
        RECT 207.600 93.600 208.400 93.700 ;
        RECT 217.200 94.300 218.000 94.400 ;
        RECT 236.400 94.300 237.200 94.400 ;
        RECT 217.200 93.700 237.200 94.300 ;
        RECT 217.200 93.600 218.000 93.700 ;
        RECT 236.400 93.600 237.200 93.700 ;
        RECT 255.600 94.300 256.400 94.400 ;
        RECT 266.800 94.300 267.600 94.400 ;
        RECT 255.600 93.700 267.600 94.300 ;
        RECT 255.600 93.600 256.400 93.700 ;
        RECT 266.800 93.600 267.600 93.700 ;
        RECT 292.400 94.300 293.200 94.400 ;
        RECT 297.200 94.300 298.000 94.400 ;
        RECT 298.800 94.300 299.600 94.400 ;
        RECT 292.400 93.700 299.600 94.300 ;
        RECT 292.400 93.600 293.200 93.700 ;
        RECT 297.200 93.600 298.000 93.700 ;
        RECT 298.800 93.600 299.600 93.700 ;
        RECT 302.000 94.300 302.800 94.400 ;
        RECT 306.800 94.300 307.600 94.400 ;
        RECT 302.000 93.700 307.600 94.300 ;
        RECT 302.000 93.600 302.800 93.700 ;
        RECT 306.800 93.600 307.600 93.700 ;
        RECT 358.000 94.300 358.800 94.400 ;
        RECT 398.000 94.300 398.800 94.400 ;
        RECT 358.000 93.700 398.800 94.300 ;
        RECT 358.000 93.600 358.800 93.700 ;
        RECT 398.000 93.600 398.800 93.700 ;
        RECT 418.800 94.300 419.600 94.400 ;
        RECT 430.000 94.300 430.800 94.400 ;
        RECT 418.800 93.700 430.800 94.300 ;
        RECT 418.800 93.600 419.600 93.700 ;
        RECT 430.000 93.600 430.800 93.700 ;
        RECT 542.000 94.300 542.800 94.400 ;
        RECT 554.800 94.300 555.600 94.400 ;
        RECT 542.000 93.700 555.600 94.300 ;
        RECT 542.000 93.600 542.800 93.700 ;
        RECT 554.800 93.600 555.600 93.700 ;
        RECT 10.800 92.300 11.600 92.400 ;
        RECT 12.400 92.300 13.200 92.400 ;
        RECT 10.800 91.700 13.200 92.300 ;
        RECT 10.800 91.600 11.600 91.700 ;
        RECT 12.400 91.600 13.200 91.700 ;
        RECT 30.000 92.300 30.800 92.400 ;
        RECT 36.400 92.300 37.200 92.400 ;
        RECT 30.000 91.700 37.200 92.300 ;
        RECT 30.000 91.600 30.800 91.700 ;
        RECT 36.400 91.600 37.200 91.700 ;
        RECT 62.000 92.300 62.800 92.400 ;
        RECT 68.400 92.300 69.200 92.400 ;
        RECT 62.000 91.700 69.200 92.300 ;
        RECT 62.000 91.600 62.800 91.700 ;
        RECT 68.400 91.600 69.200 91.700 ;
        RECT 81.200 92.300 82.000 92.400 ;
        RECT 95.600 92.300 96.400 92.400 ;
        RECT 81.200 91.700 96.400 92.300 ;
        RECT 81.200 91.600 82.000 91.700 ;
        RECT 95.600 91.600 96.400 91.700 ;
        RECT 98.800 92.300 99.600 92.400 ;
        RECT 105.200 92.300 106.000 92.400 ;
        RECT 98.800 91.700 106.000 92.300 ;
        RECT 98.800 91.600 99.600 91.700 ;
        RECT 105.200 91.600 106.000 91.700 ;
        RECT 108.400 92.300 109.200 92.400 ;
        RECT 124.400 92.300 125.200 92.400 ;
        RECT 153.200 92.300 154.000 92.400 ;
        RECT 108.400 91.700 154.000 92.300 ;
        RECT 108.400 91.600 109.200 91.700 ;
        RECT 124.400 91.600 125.200 91.700 ;
        RECT 153.200 91.600 154.000 91.700 ;
        RECT 177.200 92.300 178.000 92.400 ;
        RECT 198.000 92.300 198.800 92.400 ;
        RECT 177.200 91.700 198.800 92.300 ;
        RECT 177.200 91.600 178.000 91.700 ;
        RECT 198.000 91.600 198.800 91.700 ;
        RECT 233.200 92.300 234.000 92.400 ;
        RECT 241.200 92.300 242.000 92.400 ;
        RECT 233.200 91.700 242.000 92.300 ;
        RECT 233.200 91.600 234.000 91.700 ;
        RECT 241.200 91.600 242.000 91.700 ;
        RECT 244.400 92.300 245.200 92.400 ;
        RECT 247.600 92.300 248.400 92.400 ;
        RECT 244.400 91.700 248.400 92.300 ;
        RECT 244.400 91.600 245.200 91.700 ;
        RECT 247.600 91.600 248.400 91.700 ;
        RECT 295.600 92.300 296.400 92.400 ;
        RECT 302.000 92.300 302.800 92.400 ;
        RECT 303.600 92.300 304.400 92.400 ;
        RECT 295.600 91.700 304.400 92.300 ;
        RECT 295.600 91.600 296.400 91.700 ;
        RECT 302.000 91.600 302.800 91.700 ;
        RECT 303.600 91.600 304.400 91.700 ;
        RECT 322.800 92.300 323.600 92.400 ;
        RECT 342.000 92.300 342.800 92.400 ;
        RECT 322.800 91.700 342.800 92.300 ;
        RECT 322.800 91.600 323.600 91.700 ;
        RECT 342.000 91.600 342.800 91.700 ;
        RECT 367.600 92.300 368.400 92.400 ;
        RECT 390.000 92.300 390.800 92.400 ;
        RECT 367.600 91.700 390.800 92.300 ;
        RECT 367.600 91.600 368.400 91.700 ;
        RECT 390.000 91.600 390.800 91.700 ;
        RECT 391.600 92.300 392.400 92.400 ;
        RECT 407.600 92.300 408.400 92.400 ;
        RECT 391.600 91.700 408.400 92.300 ;
        RECT 391.600 91.600 392.400 91.700 ;
        RECT 407.600 91.600 408.400 91.700 ;
        RECT 422.000 92.300 422.800 92.400 ;
        RECT 460.400 92.300 461.200 92.400 ;
        RECT 422.000 91.700 461.200 92.300 ;
        RECT 422.000 91.600 422.800 91.700 ;
        RECT 460.400 91.600 461.200 91.700 ;
        RECT 503.600 92.300 504.400 92.400 ;
        RECT 518.000 92.300 518.800 92.400 ;
        RECT 503.600 91.700 518.800 92.300 ;
        RECT 503.600 91.600 504.400 91.700 ;
        RECT 518.000 91.600 518.800 91.700 ;
        RECT 31.600 90.300 32.400 90.400 ;
        RECT 50.800 90.300 51.600 90.400 ;
        RECT 71.600 90.300 72.400 90.400 ;
        RECT 31.600 89.700 72.400 90.300 ;
        RECT 31.600 89.600 32.400 89.700 ;
        RECT 50.800 89.600 51.600 89.700 ;
        RECT 71.600 89.600 72.400 89.700 ;
        RECT 73.200 90.300 74.000 90.400 ;
        RECT 76.400 90.300 77.200 90.400 ;
        RECT 73.200 89.700 77.200 90.300 ;
        RECT 73.200 89.600 74.000 89.700 ;
        RECT 76.400 89.600 77.200 89.700 ;
        RECT 78.000 90.300 78.800 90.400 ;
        RECT 84.400 90.300 85.200 90.400 ;
        RECT 143.600 90.300 144.400 90.400 ;
        RECT 78.000 89.700 85.200 90.300 ;
        RECT 78.000 89.600 78.800 89.700 ;
        RECT 84.400 89.600 85.200 89.700 ;
        RECT 113.300 89.700 144.400 90.300 ;
        RECT 33.200 88.300 34.000 88.400 ;
        RECT 38.000 88.300 38.800 88.400 ;
        RECT 54.000 88.300 54.800 88.400 ;
        RECT 33.200 87.700 54.800 88.300 ;
        RECT 33.200 87.600 34.000 87.700 ;
        RECT 38.000 87.600 38.800 87.700 ;
        RECT 54.000 87.600 54.800 87.700 ;
        RECT 74.800 88.300 75.600 88.400 ;
        RECT 113.300 88.300 113.900 89.700 ;
        RECT 143.600 89.600 144.400 89.700 ;
        RECT 145.200 90.300 146.000 90.400 ;
        RECT 146.800 90.300 147.600 90.400 ;
        RECT 150.000 90.300 150.800 90.400 ;
        RECT 145.200 89.700 150.800 90.300 ;
        RECT 145.200 89.600 146.000 89.700 ;
        RECT 146.800 89.600 147.600 89.700 ;
        RECT 150.000 89.600 150.800 89.700 ;
        RECT 194.800 90.300 195.600 90.400 ;
        RECT 215.600 90.300 216.400 90.400 ;
        RECT 194.800 89.700 216.400 90.300 ;
        RECT 194.800 89.600 195.600 89.700 ;
        RECT 215.600 89.600 216.400 89.700 ;
        RECT 223.600 90.300 224.400 90.400 ;
        RECT 234.800 90.300 235.600 90.400 ;
        RECT 223.600 89.700 235.600 90.300 ;
        RECT 223.600 89.600 224.400 89.700 ;
        RECT 234.800 89.600 235.600 89.700 ;
        RECT 239.600 90.300 240.400 90.400 ;
        RECT 254.000 90.300 254.800 90.400 ;
        RECT 239.600 89.700 254.800 90.300 ;
        RECT 239.600 89.600 240.400 89.700 ;
        RECT 254.000 89.600 254.800 89.700 ;
        RECT 260.400 90.300 261.200 90.400 ;
        RECT 316.400 90.300 317.200 90.400 ;
        RECT 260.400 89.700 317.200 90.300 ;
        RECT 260.400 89.600 261.200 89.700 ;
        RECT 316.400 89.600 317.200 89.700 ;
        RECT 382.000 90.300 382.800 90.400 ;
        RECT 385.200 90.300 386.000 90.400 ;
        RECT 402.800 90.300 403.600 90.400 ;
        RECT 382.000 89.700 403.600 90.300 ;
        RECT 382.000 89.600 382.800 89.700 ;
        RECT 385.200 89.600 386.000 89.700 ;
        RECT 402.800 89.600 403.600 89.700 ;
        RECT 414.000 90.300 414.800 90.400 ;
        RECT 418.800 90.300 419.600 90.400 ;
        RECT 414.000 89.700 419.600 90.300 ;
        RECT 414.000 89.600 414.800 89.700 ;
        RECT 418.800 89.600 419.600 89.700 ;
        RECT 422.000 90.300 422.800 90.400 ;
        RECT 425.200 90.300 426.000 90.400 ;
        RECT 422.000 89.700 426.000 90.300 ;
        RECT 422.000 89.600 422.800 89.700 ;
        RECT 425.200 89.600 426.000 89.700 ;
        RECT 74.800 87.700 113.900 88.300 ;
        RECT 114.800 88.300 115.600 88.400 ;
        RECT 146.800 88.300 147.600 88.400 ;
        RECT 114.800 87.700 147.600 88.300 ;
        RECT 74.800 87.600 75.600 87.700 ;
        RECT 114.800 87.600 115.600 87.700 ;
        RECT 146.800 87.600 147.600 87.700 ;
        RECT 175.600 88.300 176.400 88.400 ;
        RECT 202.800 88.300 203.600 88.400 ;
        RECT 175.600 87.700 203.600 88.300 ;
        RECT 175.600 87.600 176.400 87.700 ;
        RECT 202.800 87.600 203.600 87.700 ;
        RECT 222.000 88.300 222.800 88.400 ;
        RECT 257.200 88.300 258.000 88.400 ;
        RECT 222.000 87.700 258.000 88.300 ;
        RECT 222.000 87.600 222.800 87.700 ;
        RECT 257.200 87.600 258.000 87.700 ;
        RECT 276.400 88.300 277.200 88.400 ;
        RECT 282.800 88.300 283.600 88.400 ;
        RECT 276.400 87.700 283.600 88.300 ;
        RECT 276.400 87.600 277.200 87.700 ;
        RECT 282.800 87.600 283.600 87.700 ;
        RECT 290.800 88.300 291.600 88.400 ;
        RECT 335.600 88.300 336.400 88.400 ;
        RECT 290.800 87.700 336.400 88.300 ;
        RECT 290.800 87.600 291.600 87.700 ;
        RECT 335.600 87.600 336.400 87.700 ;
        RECT 377.200 88.300 378.000 88.400 ;
        RECT 391.600 88.300 392.400 88.400 ;
        RECT 377.200 87.700 392.400 88.300 ;
        RECT 377.200 87.600 378.000 87.700 ;
        RECT 391.600 87.600 392.400 87.700 ;
        RECT 394.800 88.300 395.600 88.400 ;
        RECT 401.200 88.300 402.000 88.400 ;
        RECT 394.800 87.700 402.000 88.300 ;
        RECT 394.800 87.600 395.600 87.700 ;
        RECT 401.200 87.600 402.000 87.700 ;
        RECT 412.400 88.300 413.200 88.400 ;
        RECT 436.400 88.300 437.200 88.400 ;
        RECT 412.400 87.700 437.200 88.300 ;
        RECT 412.400 87.600 413.200 87.700 ;
        RECT 436.400 87.600 437.200 87.700 ;
        RECT 468.400 88.300 469.200 88.400 ;
        RECT 497.200 88.300 498.000 88.400 ;
        RECT 468.400 87.700 498.000 88.300 ;
        RECT 468.400 87.600 469.200 87.700 ;
        RECT 497.200 87.600 498.000 87.700 ;
        RECT 524.400 88.300 525.200 88.400 ;
        RECT 529.200 88.300 530.000 88.400 ;
        RECT 524.400 87.700 530.000 88.300 ;
        RECT 524.400 87.600 525.200 87.700 ;
        RECT 529.200 87.600 530.000 87.700 ;
        RECT 548.400 88.300 549.200 88.400 ;
        RECT 558.000 88.300 558.800 88.400 ;
        RECT 548.400 87.700 558.800 88.300 ;
        RECT 548.400 87.600 549.200 87.700 ;
        RECT 558.000 87.600 558.800 87.700 ;
        RECT 47.600 86.300 48.400 86.400 ;
        RECT 57.200 86.300 58.000 86.400 ;
        RECT 47.600 85.700 58.000 86.300 ;
        RECT 47.600 85.600 48.400 85.700 ;
        RECT 57.200 85.600 58.000 85.700 ;
        RECT 121.200 86.300 122.000 86.400 ;
        RECT 156.400 86.300 157.200 86.400 ;
        RECT 121.200 85.700 157.200 86.300 ;
        RECT 121.200 85.600 122.000 85.700 ;
        RECT 156.400 85.600 157.200 85.700 ;
        RECT 218.800 86.300 219.600 86.400 ;
        RECT 249.200 86.300 250.000 86.400 ;
        RECT 218.800 85.700 250.000 86.300 ;
        RECT 218.800 85.600 219.600 85.700 ;
        RECT 249.200 85.600 250.000 85.700 ;
        RECT 484.400 86.300 485.200 86.400 ;
        RECT 487.600 86.300 488.400 86.400 ;
        RECT 484.400 85.700 488.400 86.300 ;
        RECT 484.400 85.600 485.200 85.700 ;
        RECT 487.600 85.600 488.400 85.700 ;
        RECT 199.600 84.300 200.400 84.400 ;
        RECT 225.200 84.300 226.000 84.400 ;
        RECT 199.600 83.700 226.000 84.300 ;
        RECT 199.600 83.600 200.400 83.700 ;
        RECT 225.200 83.600 226.000 83.700 ;
        RECT 482.800 84.300 483.600 84.400 ;
        RECT 503.600 84.300 504.400 84.400 ;
        RECT 482.800 83.700 504.400 84.300 ;
        RECT 482.800 83.600 483.600 83.700 ;
        RECT 503.600 83.600 504.400 83.700 ;
        RECT 17.200 82.300 18.000 82.400 ;
        RECT 30.000 82.300 30.800 82.400 ;
        RECT 17.200 81.700 30.800 82.300 ;
        RECT 17.200 81.600 18.000 81.700 ;
        RECT 30.000 81.600 30.800 81.700 ;
        RECT 102.000 82.300 102.800 82.400 ;
        RECT 121.200 82.300 122.000 82.400 ;
        RECT 102.000 81.700 122.000 82.300 ;
        RECT 102.000 81.600 102.800 81.700 ;
        RECT 121.200 81.600 122.000 81.700 ;
        RECT 190.000 82.300 190.800 82.400 ;
        RECT 217.200 82.300 218.000 82.400 ;
        RECT 190.000 81.700 218.000 82.300 ;
        RECT 190.000 81.600 190.800 81.700 ;
        RECT 217.200 81.600 218.000 81.700 ;
        RECT 409.200 82.300 410.000 82.400 ;
        RECT 433.200 82.300 434.000 82.400 ;
        RECT 409.200 81.700 434.000 82.300 ;
        RECT 409.200 81.600 410.000 81.700 ;
        RECT 433.200 81.600 434.000 81.700 ;
        RECT 14.000 80.300 14.800 80.400 ;
        RECT 34.800 80.300 35.600 80.400 ;
        RECT 103.600 80.300 104.400 80.400 ;
        RECT 14.000 79.700 104.400 80.300 ;
        RECT 14.000 79.600 14.800 79.700 ;
        RECT 34.800 79.600 35.600 79.700 ;
        RECT 103.600 79.600 104.400 79.700 ;
        RECT 20.400 78.300 21.200 78.400 ;
        RECT 28.400 78.300 29.200 78.400 ;
        RECT 20.400 77.700 29.200 78.300 ;
        RECT 20.400 77.600 21.200 77.700 ;
        RECT 28.400 77.600 29.200 77.700 ;
        RECT 41.200 78.300 42.000 78.400 ;
        RECT 78.000 78.300 78.800 78.400 ;
        RECT 41.200 77.700 78.800 78.300 ;
        RECT 41.200 77.600 42.000 77.700 ;
        RECT 78.000 77.600 78.800 77.700 ;
        RECT 361.200 78.300 362.000 78.400 ;
        RECT 423.600 78.300 424.400 78.400 ;
        RECT 426.800 78.300 427.600 78.400 ;
        RECT 361.200 77.700 427.600 78.300 ;
        RECT 361.200 77.600 362.000 77.700 ;
        RECT 423.600 77.600 424.400 77.700 ;
        RECT 426.800 77.600 427.600 77.700 ;
        RECT 9.200 76.300 10.000 76.400 ;
        RECT 26.800 76.300 27.600 76.400 ;
        RECT 9.200 75.700 27.600 76.300 ;
        RECT 9.200 75.600 10.000 75.700 ;
        RECT 26.800 75.600 27.600 75.700 ;
        RECT 39.600 76.300 40.400 76.400 ;
        RECT 66.800 76.300 67.600 76.400 ;
        RECT 39.600 75.700 67.600 76.300 ;
        RECT 39.600 75.600 40.400 75.700 ;
        RECT 66.800 75.600 67.600 75.700 ;
        RECT 76.400 76.300 77.200 76.400 ;
        RECT 82.800 76.300 83.600 76.400 ;
        RECT 76.400 75.700 83.600 76.300 ;
        RECT 76.400 75.600 77.200 75.700 ;
        RECT 82.800 75.600 83.600 75.700 ;
        RECT 414.000 76.300 414.800 76.400 ;
        RECT 479.600 76.300 480.400 76.400 ;
        RECT 414.000 75.700 480.400 76.300 ;
        RECT 414.000 75.600 414.800 75.700 ;
        RECT 479.600 75.600 480.400 75.700 ;
        RECT 12.400 74.300 13.200 74.400 ;
        RECT 23.600 74.300 24.400 74.400 ;
        RECT 12.400 73.700 24.400 74.300 ;
        RECT 12.400 73.600 13.200 73.700 ;
        RECT 23.600 73.600 24.400 73.700 ;
        RECT 25.200 74.300 26.000 74.400 ;
        RECT 73.200 74.300 74.000 74.400 ;
        RECT 79.600 74.300 80.400 74.400 ;
        RECT 25.200 73.700 80.400 74.300 ;
        RECT 25.200 73.600 26.000 73.700 ;
        RECT 73.200 73.600 74.000 73.700 ;
        RECT 79.600 73.600 80.400 73.700 ;
        RECT 82.800 74.300 83.600 74.400 ;
        RECT 113.200 74.300 114.000 74.400 ;
        RECT 130.800 74.300 131.600 74.400 ;
        RECT 137.200 74.300 138.000 74.400 ;
        RECT 82.800 73.700 138.000 74.300 ;
        RECT 82.800 73.600 83.600 73.700 ;
        RECT 113.200 73.600 114.000 73.700 ;
        RECT 130.800 73.600 131.600 73.700 ;
        RECT 137.200 73.600 138.000 73.700 ;
        RECT 174.000 74.300 174.800 74.400 ;
        RECT 186.800 74.300 187.600 74.400 ;
        RECT 220.400 74.300 221.200 74.400 ;
        RECT 174.000 73.700 221.200 74.300 ;
        RECT 174.000 73.600 174.800 73.700 ;
        RECT 186.800 73.600 187.600 73.700 ;
        RECT 220.400 73.600 221.200 73.700 ;
        RECT 228.400 74.300 229.200 74.400 ;
        RECT 244.400 74.300 245.200 74.400 ;
        RECT 228.400 73.700 245.200 74.300 ;
        RECT 228.400 73.600 229.200 73.700 ;
        RECT 244.400 73.600 245.200 73.700 ;
        RECT 270.000 74.300 270.800 74.400 ;
        RECT 316.400 74.300 317.200 74.400 ;
        RECT 270.000 73.700 317.200 74.300 ;
        RECT 270.000 73.600 270.800 73.700 ;
        RECT 316.400 73.600 317.200 73.700 ;
        RECT 329.200 74.300 330.000 74.400 ;
        RECT 423.600 74.300 424.400 74.400 ;
        RECT 438.000 74.300 438.800 74.400 ;
        RECT 329.200 73.700 438.800 74.300 ;
        RECT 329.200 73.600 330.000 73.700 ;
        RECT 423.600 73.600 424.400 73.700 ;
        RECT 438.000 73.600 438.800 73.700 ;
        RECT 460.400 74.300 461.200 74.400 ;
        RECT 463.600 74.300 464.400 74.400 ;
        RECT 460.400 73.700 464.400 74.300 ;
        RECT 460.400 73.600 461.200 73.700 ;
        RECT 463.600 73.600 464.400 73.700 ;
        RECT 478.000 74.300 478.800 74.400 ;
        RECT 494.000 74.300 494.800 74.400 ;
        RECT 478.000 73.700 494.800 74.300 ;
        RECT 478.000 73.600 478.800 73.700 ;
        RECT 494.000 73.600 494.800 73.700 ;
        RECT 12.400 72.300 13.200 72.400 ;
        RECT 15.600 72.300 16.400 72.400 ;
        RECT 17.200 72.300 18.000 72.400 ;
        RECT 12.400 71.700 18.000 72.300 ;
        RECT 12.400 71.600 13.200 71.700 ;
        RECT 15.600 71.600 16.400 71.700 ;
        RECT 17.200 71.600 18.000 71.700 ;
        RECT 31.600 72.300 32.400 72.400 ;
        RECT 44.400 72.300 45.200 72.400 ;
        RECT 31.600 71.700 45.200 72.300 ;
        RECT 31.600 71.600 32.400 71.700 ;
        RECT 44.400 71.600 45.200 71.700 ;
        RECT 66.800 72.300 67.600 72.400 ;
        RECT 74.800 72.300 75.600 72.400 ;
        RECT 76.400 72.300 77.200 72.400 ;
        RECT 66.800 71.700 77.200 72.300 ;
        RECT 66.800 71.600 67.600 71.700 ;
        RECT 74.800 71.600 75.600 71.700 ;
        RECT 76.400 71.600 77.200 71.700 ;
        RECT 102.000 72.300 102.800 72.400 ;
        RECT 105.200 72.300 106.000 72.400 ;
        RECT 102.000 71.700 106.000 72.300 ;
        RECT 102.000 71.600 102.800 71.700 ;
        RECT 105.200 71.600 106.000 71.700 ;
        RECT 210.800 72.300 211.600 72.400 ;
        RECT 244.400 72.300 245.200 72.400 ;
        RECT 250.800 72.300 251.600 72.400 ;
        RECT 210.800 71.700 243.500 72.300 ;
        RECT 210.800 71.600 211.600 71.700 ;
        RECT 12.400 70.300 13.200 70.400 ;
        RECT 14.000 70.300 14.800 70.400 ;
        RECT 18.800 70.300 19.600 70.400 ;
        RECT 12.400 69.700 19.600 70.300 ;
        RECT 12.400 69.600 13.200 69.700 ;
        RECT 14.000 69.600 14.800 69.700 ;
        RECT 18.800 69.600 19.600 69.700 ;
        RECT 42.800 70.300 43.600 70.400 ;
        RECT 50.800 70.300 51.600 70.400 ;
        RECT 42.800 69.700 51.600 70.300 ;
        RECT 42.800 69.600 43.600 69.700 ;
        RECT 50.800 69.600 51.600 69.700 ;
        RECT 55.600 70.300 56.400 70.400 ;
        RECT 62.000 70.300 62.800 70.400 ;
        RECT 55.600 69.700 62.800 70.300 ;
        RECT 55.600 69.600 56.400 69.700 ;
        RECT 62.000 69.600 62.800 69.700 ;
        RECT 116.400 70.300 117.200 70.400 ;
        RECT 122.800 70.300 123.600 70.400 ;
        RECT 116.400 69.700 123.600 70.300 ;
        RECT 116.400 69.600 117.200 69.700 ;
        RECT 122.800 69.600 123.600 69.700 ;
        RECT 142.000 70.300 142.800 70.400 ;
        RECT 159.600 70.300 160.400 70.400 ;
        RECT 142.000 69.700 160.400 70.300 ;
        RECT 142.000 69.600 142.800 69.700 ;
        RECT 159.600 69.600 160.400 69.700 ;
        RECT 182.000 70.300 182.800 70.400 ;
        RECT 188.400 70.300 189.200 70.400 ;
        RECT 193.200 70.300 194.000 70.400 ;
        RECT 182.000 69.700 194.000 70.300 ;
        RECT 182.000 69.600 182.800 69.700 ;
        RECT 188.400 69.600 189.200 69.700 ;
        RECT 193.200 69.600 194.000 69.700 ;
        RECT 206.000 70.300 206.800 70.400 ;
        RECT 218.800 70.300 219.600 70.400 ;
        RECT 206.000 69.700 219.600 70.300 ;
        RECT 242.900 70.300 243.500 71.700 ;
        RECT 244.400 71.700 251.600 72.300 ;
        RECT 244.400 71.600 245.200 71.700 ;
        RECT 250.800 71.600 251.600 71.700 ;
        RECT 254.000 72.300 254.800 72.400 ;
        RECT 260.400 72.300 261.200 72.400 ;
        RECT 284.400 72.300 285.200 72.400 ;
        RECT 254.000 71.700 285.200 72.300 ;
        RECT 254.000 71.600 254.800 71.700 ;
        RECT 260.400 71.600 261.200 71.700 ;
        RECT 284.400 71.600 285.200 71.700 ;
        RECT 286.000 72.300 286.800 72.400 ;
        RECT 306.800 72.300 307.600 72.400 ;
        RECT 286.000 71.700 307.600 72.300 ;
        RECT 286.000 71.600 286.800 71.700 ;
        RECT 306.800 71.600 307.600 71.700 ;
        RECT 308.400 72.300 309.200 72.400 ;
        RECT 367.600 72.300 368.400 72.400 ;
        RECT 308.400 71.700 368.400 72.300 ;
        RECT 308.400 71.600 309.200 71.700 ;
        RECT 367.600 71.600 368.400 71.700 ;
        RECT 399.600 72.300 400.400 72.400 ;
        RECT 406.000 72.300 406.800 72.400 ;
        RECT 414.000 72.300 414.800 72.400 ;
        RECT 399.600 71.700 414.800 72.300 ;
        RECT 399.600 71.600 400.400 71.700 ;
        RECT 406.000 71.600 406.800 71.700 ;
        RECT 414.000 71.600 414.800 71.700 ;
        RECT 428.400 72.300 429.200 72.400 ;
        RECT 474.800 72.300 475.600 72.400 ;
        RECT 428.400 71.700 475.600 72.300 ;
        RECT 428.400 71.600 429.200 71.700 ;
        RECT 474.800 71.600 475.600 71.700 ;
        RECT 478.000 72.300 478.800 72.400 ;
        RECT 479.600 72.300 480.400 72.400 ;
        RECT 478.000 71.700 480.400 72.300 ;
        RECT 478.000 71.600 478.800 71.700 ;
        RECT 479.600 71.600 480.400 71.700 ;
        RECT 495.600 72.300 496.400 72.400 ;
        RECT 524.400 72.300 525.200 72.400 ;
        RECT 532.400 72.300 533.200 72.400 ;
        RECT 495.600 71.700 533.200 72.300 ;
        RECT 495.600 71.600 496.400 71.700 ;
        RECT 524.400 71.600 525.200 71.700 ;
        RECT 532.400 71.600 533.200 71.700 ;
        RECT 559.600 72.300 560.400 72.400 ;
        RECT 566.000 72.300 566.800 72.400 ;
        RECT 559.600 71.700 566.800 72.300 ;
        RECT 559.600 71.600 560.400 71.700 ;
        RECT 566.000 71.600 566.800 71.700 ;
        RECT 246.000 70.300 246.800 70.400 ;
        RECT 242.900 69.700 246.800 70.300 ;
        RECT 206.000 69.600 206.800 69.700 ;
        RECT 218.800 69.600 219.600 69.700 ;
        RECT 246.000 69.600 246.800 69.700 ;
        RECT 254.000 70.300 254.800 70.400 ;
        RECT 258.800 70.300 259.600 70.400 ;
        RECT 254.000 69.700 259.600 70.300 ;
        RECT 254.000 69.600 254.800 69.700 ;
        RECT 258.800 69.600 259.600 69.700 ;
        RECT 287.600 70.300 288.400 70.400 ;
        RECT 298.800 70.300 299.600 70.400 ;
        RECT 287.600 69.700 299.600 70.300 ;
        RECT 287.600 69.600 288.400 69.700 ;
        RECT 298.800 69.600 299.600 69.700 ;
        RECT 303.600 70.300 304.400 70.400 ;
        RECT 306.800 70.300 307.600 70.400 ;
        RECT 303.600 69.700 307.600 70.300 ;
        RECT 303.600 69.600 304.400 69.700 ;
        RECT 306.800 69.600 307.600 69.700 ;
        RECT 308.400 70.300 309.200 70.400 ;
        RECT 311.600 70.300 312.400 70.400 ;
        RECT 308.400 69.700 312.400 70.300 ;
        RECT 308.400 69.600 309.200 69.700 ;
        RECT 311.600 69.600 312.400 69.700 ;
        RECT 322.800 70.300 323.600 70.400 ;
        RECT 329.200 70.300 330.000 70.400 ;
        RECT 322.800 69.700 330.000 70.300 ;
        RECT 322.800 69.600 323.600 69.700 ;
        RECT 329.200 69.600 330.000 69.700 ;
        RECT 394.800 70.300 395.600 70.400 ;
        RECT 407.600 70.300 408.400 70.400 ;
        RECT 410.800 70.300 411.600 70.400 ;
        RECT 394.800 69.700 411.600 70.300 ;
        RECT 394.800 69.600 395.600 69.700 ;
        RECT 407.600 69.600 408.400 69.700 ;
        RECT 410.800 69.600 411.600 69.700 ;
        RECT 431.600 70.300 432.400 70.400 ;
        RECT 438.000 70.300 438.800 70.400 ;
        RECT 452.400 70.300 453.200 70.400 ;
        RECT 431.600 69.700 453.200 70.300 ;
        RECT 431.600 69.600 432.400 69.700 ;
        RECT 438.000 69.600 438.800 69.700 ;
        RECT 452.400 69.600 453.200 69.700 ;
        RECT 458.800 70.300 459.600 70.400 ;
        RECT 460.400 70.300 461.200 70.400 ;
        RECT 458.800 69.700 461.200 70.300 ;
        RECT 458.800 69.600 459.600 69.700 ;
        RECT 460.400 69.600 461.200 69.700 ;
        RECT 497.200 70.300 498.000 70.400 ;
        RECT 498.800 70.300 499.600 70.400 ;
        RECT 497.200 69.700 499.600 70.300 ;
        RECT 497.200 69.600 498.000 69.700 ;
        RECT 498.800 69.600 499.600 69.700 ;
        RECT 506.800 70.300 507.600 70.400 ;
        RECT 518.000 70.300 518.800 70.400 ;
        RECT 506.800 69.700 518.800 70.300 ;
        RECT 506.800 69.600 507.600 69.700 ;
        RECT 518.000 69.600 518.800 69.700 ;
        RECT 17.200 68.300 18.000 68.400 ;
        RECT 36.400 68.300 37.200 68.400 ;
        RECT 17.200 67.700 37.200 68.300 ;
        RECT 50.900 68.300 51.500 69.600 ;
        RECT 60.400 68.300 61.200 68.400 ;
        RECT 50.900 67.700 61.200 68.300 ;
        RECT 17.200 67.600 18.000 67.700 ;
        RECT 36.400 67.600 37.200 67.700 ;
        RECT 60.400 67.600 61.200 67.700 ;
        RECT 62.000 68.300 62.800 68.400 ;
        RECT 76.400 68.300 77.200 68.400 ;
        RECT 62.000 67.700 77.200 68.300 ;
        RECT 62.000 67.600 62.800 67.700 ;
        RECT 76.400 67.600 77.200 67.700 ;
        RECT 92.400 68.300 93.200 68.400 ;
        RECT 95.600 68.300 96.400 68.400 ;
        RECT 97.200 68.300 98.000 68.400 ;
        RECT 92.400 67.700 98.000 68.300 ;
        RECT 92.400 67.600 93.200 67.700 ;
        RECT 95.600 67.600 96.400 67.700 ;
        RECT 97.200 67.600 98.000 67.700 ;
        RECT 98.800 67.600 99.600 68.400 ;
        RECT 102.000 68.300 102.800 68.400 ;
        RECT 174.000 68.300 174.800 68.400 ;
        RECT 102.000 67.700 174.800 68.300 ;
        RECT 102.000 67.600 102.800 67.700 ;
        RECT 174.000 67.600 174.800 67.700 ;
        RECT 186.800 68.300 187.600 68.400 ;
        RECT 196.400 68.300 197.200 68.400 ;
        RECT 202.800 68.300 203.600 68.400 ;
        RECT 186.800 67.700 203.600 68.300 ;
        RECT 186.800 67.600 187.600 67.700 ;
        RECT 196.400 67.600 197.200 67.700 ;
        RECT 202.800 67.600 203.600 67.700 ;
        RECT 223.600 68.300 224.400 68.400 ;
        RECT 226.800 68.300 227.600 68.400 ;
        RECT 223.600 67.700 227.600 68.300 ;
        RECT 223.600 67.600 224.400 67.700 ;
        RECT 226.800 67.600 227.600 67.700 ;
        RECT 228.400 68.300 229.200 68.400 ;
        RECT 239.600 68.300 240.400 68.400 ;
        RECT 249.200 68.300 250.000 68.400 ;
        RECT 228.400 67.700 240.400 68.300 ;
        RECT 228.400 67.600 229.200 67.700 ;
        RECT 239.600 67.600 240.400 67.700 ;
        RECT 244.500 67.700 250.000 68.300 ;
        RECT 7.600 66.300 8.400 66.400 ;
        RECT 15.600 66.300 16.400 66.400 ;
        RECT 22.000 66.300 22.800 66.400 ;
        RECT 31.600 66.300 32.400 66.400 ;
        RECT 7.600 65.700 32.400 66.300 ;
        RECT 36.500 66.300 37.100 67.600 ;
        RECT 86.000 66.300 86.800 66.400 ;
        RECT 94.000 66.300 94.800 66.400 ;
        RECT 36.500 65.700 94.800 66.300 ;
        RECT 7.600 65.600 8.400 65.700 ;
        RECT 15.600 65.600 16.400 65.700 ;
        RECT 22.000 65.600 22.800 65.700 ;
        RECT 31.600 65.600 32.400 65.700 ;
        RECT 86.000 65.600 86.800 65.700 ;
        RECT 94.000 65.600 94.800 65.700 ;
        RECT 103.600 66.300 104.400 66.400 ;
        RECT 106.800 66.300 107.600 66.400 ;
        RECT 113.200 66.300 114.000 66.400 ;
        RECT 153.200 66.300 154.000 66.400 ;
        RECT 164.400 66.300 165.200 66.400 ;
        RECT 103.600 65.700 165.200 66.300 ;
        RECT 174.100 66.300 174.700 67.600 ;
        RECT 180.400 66.300 181.200 66.400 ;
        RECT 198.000 66.300 198.800 66.400 ;
        RECT 174.100 65.700 198.800 66.300 ;
        RECT 103.600 65.600 104.400 65.700 ;
        RECT 106.800 65.600 107.600 65.700 ;
        RECT 113.200 65.600 114.000 65.700 ;
        RECT 153.200 65.600 154.000 65.700 ;
        RECT 164.400 65.600 165.200 65.700 ;
        RECT 180.400 65.600 181.200 65.700 ;
        RECT 198.000 65.600 198.800 65.700 ;
        RECT 206.000 66.300 206.800 66.400 ;
        RECT 214.000 66.300 214.800 66.400 ;
        RECT 206.000 65.700 214.800 66.300 ;
        RECT 206.000 65.600 206.800 65.700 ;
        RECT 214.000 65.600 214.800 65.700 ;
        RECT 215.600 66.300 216.400 66.400 ;
        RECT 244.500 66.300 245.100 67.700 ;
        RECT 249.200 67.600 250.000 67.700 ;
        RECT 268.400 68.300 269.200 68.400 ;
        RECT 281.200 68.300 282.000 68.400 ;
        RECT 268.400 67.700 282.000 68.300 ;
        RECT 268.400 67.600 269.200 67.700 ;
        RECT 281.200 67.600 282.000 67.700 ;
        RECT 282.800 68.300 283.600 68.400 ;
        RECT 308.400 68.300 309.200 68.400 ;
        RECT 332.400 68.300 333.200 68.400 ;
        RECT 282.800 67.700 333.200 68.300 ;
        RECT 282.800 67.600 283.600 67.700 ;
        RECT 308.400 67.600 309.200 67.700 ;
        RECT 332.400 67.600 333.200 67.700 ;
        RECT 353.200 68.300 354.000 68.400 ;
        RECT 364.400 68.300 365.200 68.400 ;
        RECT 353.200 67.700 365.200 68.300 ;
        RECT 353.200 67.600 354.000 67.700 ;
        RECT 364.400 67.600 365.200 67.700 ;
        RECT 380.400 68.300 381.200 68.400 ;
        RECT 390.000 68.300 390.800 68.400 ;
        RECT 396.400 68.300 397.200 68.400 ;
        RECT 380.400 67.700 397.200 68.300 ;
        RECT 380.400 67.600 381.200 67.700 ;
        RECT 390.000 67.600 390.800 67.700 ;
        RECT 396.400 67.600 397.200 67.700 ;
        RECT 438.000 68.300 438.800 68.400 ;
        RECT 455.600 68.300 456.400 68.400 ;
        RECT 438.000 67.700 456.400 68.300 ;
        RECT 438.000 67.600 438.800 67.700 ;
        RECT 455.600 67.600 456.400 67.700 ;
        RECT 458.800 68.300 459.600 68.400 ;
        RECT 478.000 68.300 478.800 68.400 ;
        RECT 458.800 67.700 478.800 68.300 ;
        RECT 458.800 67.600 459.600 67.700 ;
        RECT 478.000 67.600 478.800 67.700 ;
        RECT 484.400 68.300 485.200 68.400 ;
        RECT 492.400 68.300 493.200 68.400 ;
        RECT 484.400 67.700 493.200 68.300 ;
        RECT 484.400 67.600 485.200 67.700 ;
        RECT 492.400 67.600 493.200 67.700 ;
        RECT 498.800 68.300 499.600 68.400 ;
        RECT 505.200 68.300 506.000 68.400 ;
        RECT 498.800 67.700 506.000 68.300 ;
        RECT 498.800 67.600 499.600 67.700 ;
        RECT 505.200 67.600 506.000 67.700 ;
        RECT 508.400 68.300 509.200 68.400 ;
        RECT 510.000 68.300 510.800 68.400 ;
        RECT 508.400 67.700 510.800 68.300 ;
        RECT 508.400 67.600 509.200 67.700 ;
        RECT 510.000 67.600 510.800 67.700 ;
        RECT 514.800 68.300 515.600 68.400 ;
        RECT 519.600 68.300 520.400 68.400 ;
        RECT 514.800 67.700 520.400 68.300 ;
        RECT 514.800 67.600 515.600 67.700 ;
        RECT 519.600 67.600 520.400 67.700 ;
        RECT 530.800 68.300 531.600 68.400 ;
        RECT 540.400 68.300 541.200 68.400 ;
        RECT 553.200 68.300 554.000 68.400 ;
        RECT 530.800 67.700 554.000 68.300 ;
        RECT 530.800 67.600 531.600 67.700 ;
        RECT 540.400 67.600 541.200 67.700 ;
        RECT 553.200 67.600 554.000 67.700 ;
        RECT 215.600 65.700 245.100 66.300 ;
        RECT 246.000 66.300 246.800 66.400 ;
        RECT 255.600 66.300 256.400 66.400 ;
        RECT 246.000 65.700 256.400 66.300 ;
        RECT 215.600 65.600 216.400 65.700 ;
        RECT 246.000 65.600 246.800 65.700 ;
        RECT 255.600 65.600 256.400 65.700 ;
        RECT 262.000 66.300 262.800 66.400 ;
        RECT 263.600 66.300 264.400 66.400 ;
        RECT 282.800 66.300 283.600 66.400 ;
        RECT 262.000 65.700 283.600 66.300 ;
        RECT 262.000 65.600 262.800 65.700 ;
        RECT 263.600 65.600 264.400 65.700 ;
        RECT 282.800 65.600 283.600 65.700 ;
        RECT 284.400 66.300 285.200 66.400 ;
        RECT 303.600 66.300 304.400 66.400 ;
        RECT 306.800 66.300 307.600 66.400 ;
        RECT 319.600 66.300 320.400 66.400 ;
        RECT 284.400 65.700 307.600 66.300 ;
        RECT 284.400 65.600 285.200 65.700 ;
        RECT 303.600 65.600 304.400 65.700 ;
        RECT 306.800 65.600 307.600 65.700 ;
        RECT 308.500 65.700 320.400 66.300 ;
        RECT 31.600 64.300 32.400 64.400 ;
        RECT 38.000 64.300 38.800 64.400 ;
        RECT 31.600 63.700 38.800 64.300 ;
        RECT 31.600 63.600 32.400 63.700 ;
        RECT 38.000 63.600 38.800 63.700 ;
        RECT 50.800 64.300 51.600 64.400 ;
        RECT 63.600 64.300 64.400 64.400 ;
        RECT 50.800 63.700 64.400 64.300 ;
        RECT 50.800 63.600 51.600 63.700 ;
        RECT 63.600 63.600 64.400 63.700 ;
        RECT 105.200 64.300 106.000 64.400 ;
        RECT 110.000 64.300 110.800 64.400 ;
        RECT 121.200 64.300 122.000 64.400 ;
        RECT 105.200 63.700 122.000 64.300 ;
        RECT 105.200 63.600 106.000 63.700 ;
        RECT 110.000 63.600 110.800 63.700 ;
        RECT 121.200 63.600 122.000 63.700 ;
        RECT 122.800 64.300 123.600 64.400 ;
        RECT 143.600 64.300 144.400 64.400 ;
        RECT 150.000 64.300 150.800 64.400 ;
        RECT 153.200 64.300 154.000 64.400 ;
        RECT 122.800 63.700 154.000 64.300 ;
        RECT 122.800 63.600 123.600 63.700 ;
        RECT 143.600 63.600 144.400 63.700 ;
        RECT 150.000 63.600 150.800 63.700 ;
        RECT 153.200 63.600 154.000 63.700 ;
        RECT 172.400 63.600 173.200 64.400 ;
        RECT 183.600 64.300 184.400 64.400 ;
        RECT 191.600 64.300 192.400 64.400 ;
        RECT 196.400 64.300 197.200 64.400 ;
        RECT 183.600 63.700 197.200 64.300 ;
        RECT 183.600 63.600 184.400 63.700 ;
        RECT 191.600 63.600 192.400 63.700 ;
        RECT 196.400 63.600 197.200 63.700 ;
        RECT 212.400 64.300 213.200 64.400 ;
        RECT 220.400 64.300 221.200 64.400 ;
        RECT 226.800 64.300 227.600 64.400 ;
        RECT 212.400 63.700 227.600 64.300 ;
        RECT 212.400 63.600 213.200 63.700 ;
        RECT 220.400 63.600 221.200 63.700 ;
        RECT 226.800 63.600 227.600 63.700 ;
        RECT 238.000 64.300 238.800 64.400 ;
        RECT 244.400 64.300 245.200 64.400 ;
        RECT 238.000 63.700 245.200 64.300 ;
        RECT 238.000 63.600 238.800 63.700 ;
        RECT 244.400 63.600 245.200 63.700 ;
        RECT 247.600 64.300 248.400 64.400 ;
        RECT 262.000 64.300 262.800 64.400 ;
        RECT 273.200 64.300 274.000 64.400 ;
        RECT 247.600 63.700 274.000 64.300 ;
        RECT 247.600 63.600 248.400 63.700 ;
        RECT 262.000 63.600 262.800 63.700 ;
        RECT 273.200 63.600 274.000 63.700 ;
        RECT 281.200 64.300 282.000 64.400 ;
        RECT 286.000 64.300 286.800 64.400 ;
        RECT 300.400 64.300 301.200 64.400 ;
        RECT 302.000 64.300 302.800 64.400 ;
        RECT 281.200 63.700 286.800 64.300 ;
        RECT 281.200 63.600 282.000 63.700 ;
        RECT 286.000 63.600 286.800 63.700 ;
        RECT 287.700 63.700 299.500 64.300 ;
        RECT 20.400 62.300 21.200 62.400 ;
        RECT 42.800 62.300 43.600 62.400 ;
        RECT 55.600 62.300 56.400 62.400 ;
        RECT 79.600 62.300 80.400 62.400 ;
        RECT 20.400 61.700 80.400 62.300 ;
        RECT 20.400 61.600 21.200 61.700 ;
        RECT 42.800 61.600 43.600 61.700 ;
        RECT 55.600 61.600 56.400 61.700 ;
        RECT 79.600 61.600 80.400 61.700 ;
        RECT 108.400 62.300 109.200 62.400 ;
        RECT 113.200 62.300 114.000 62.400 ;
        RECT 108.400 61.700 114.000 62.300 ;
        RECT 108.400 61.600 109.200 61.700 ;
        RECT 113.200 61.600 114.000 61.700 ;
        RECT 114.800 62.300 115.600 62.400 ;
        RECT 118.000 62.300 118.800 62.400 ;
        RECT 114.800 61.700 118.800 62.300 ;
        RECT 114.800 61.600 115.600 61.700 ;
        RECT 118.000 61.600 118.800 61.700 ;
        RECT 119.600 62.300 120.400 62.400 ;
        RECT 140.400 62.300 141.200 62.400 ;
        RECT 146.800 62.300 147.600 62.400 ;
        RECT 119.600 61.700 147.600 62.300 ;
        RECT 119.600 61.600 120.400 61.700 ;
        RECT 140.400 61.600 141.200 61.700 ;
        RECT 146.800 61.600 147.600 61.700 ;
        RECT 148.400 62.300 149.200 62.400 ;
        RECT 166.000 62.300 166.800 62.400 ;
        RECT 178.800 62.300 179.600 62.400 ;
        RECT 148.400 61.700 179.600 62.300 ;
        RECT 148.400 61.600 149.200 61.700 ;
        RECT 166.000 61.600 166.800 61.700 ;
        RECT 178.800 61.600 179.600 61.700 ;
        RECT 206.000 62.300 206.800 62.400 ;
        RECT 287.700 62.300 288.300 63.700 ;
        RECT 206.000 61.700 288.300 62.300 ;
        RECT 298.900 62.300 299.500 63.700 ;
        RECT 300.400 63.700 302.800 64.300 ;
        RECT 300.400 63.600 301.200 63.700 ;
        RECT 302.000 63.600 302.800 63.700 ;
        RECT 303.600 64.300 304.400 64.400 ;
        RECT 308.500 64.300 309.100 65.700 ;
        RECT 319.600 65.600 320.400 65.700 ;
        RECT 321.200 66.300 322.000 66.400 ;
        RECT 327.600 66.300 328.400 66.400 ;
        RECT 321.200 65.700 328.400 66.300 ;
        RECT 321.200 65.600 322.000 65.700 ;
        RECT 327.600 65.600 328.400 65.700 ;
        RECT 426.800 66.300 427.600 66.400 ;
        RECT 430.000 66.300 430.800 66.400 ;
        RECT 434.800 66.300 435.600 66.400 ;
        RECT 426.800 65.700 435.600 66.300 ;
        RECT 426.800 65.600 427.600 65.700 ;
        RECT 430.000 65.600 430.800 65.700 ;
        RECT 434.800 65.600 435.600 65.700 ;
        RECT 454.000 66.300 454.800 66.400 ;
        RECT 462.000 66.300 462.800 66.400 ;
        RECT 454.000 65.700 462.800 66.300 ;
        RECT 454.000 65.600 454.800 65.700 ;
        RECT 462.000 65.600 462.800 65.700 ;
        RECT 471.600 66.300 472.400 66.400 ;
        RECT 476.400 66.300 477.200 66.400 ;
        RECT 471.600 65.700 477.200 66.300 ;
        RECT 471.600 65.600 472.400 65.700 ;
        RECT 476.400 65.600 477.200 65.700 ;
        RECT 478.000 66.300 478.800 66.400 ;
        RECT 484.400 66.300 485.200 66.400 ;
        RECT 497.200 66.300 498.000 66.400 ;
        RECT 478.000 65.700 498.000 66.300 ;
        RECT 478.000 65.600 478.800 65.700 ;
        RECT 484.400 65.600 485.200 65.700 ;
        RECT 497.200 65.600 498.000 65.700 ;
        RECT 498.800 65.600 499.600 66.400 ;
        RECT 510.000 66.300 510.800 66.400 ;
        RECT 514.800 66.300 515.600 66.400 ;
        RECT 510.000 65.700 515.600 66.300 ;
        RECT 510.000 65.600 510.800 65.700 ;
        RECT 514.800 65.600 515.600 65.700 ;
        RECT 519.600 66.300 520.400 66.400 ;
        RECT 529.200 66.300 530.000 66.400 ;
        RECT 519.600 65.700 530.000 66.300 ;
        RECT 519.600 65.600 520.400 65.700 ;
        RECT 529.200 65.600 530.000 65.700 ;
        RECT 303.600 63.700 309.100 64.300 ;
        RECT 310.000 64.300 310.800 64.400 ;
        RECT 324.400 64.300 325.200 64.400 ;
        RECT 310.000 63.700 325.200 64.300 ;
        RECT 303.600 63.600 304.400 63.700 ;
        RECT 310.000 63.600 310.800 63.700 ;
        RECT 324.400 63.600 325.200 63.700 ;
        RECT 329.200 64.300 330.000 64.400 ;
        RECT 334.000 64.300 334.800 64.400 ;
        RECT 329.200 63.700 334.800 64.300 ;
        RECT 329.200 63.600 330.000 63.700 ;
        RECT 334.000 63.600 334.800 63.700 ;
        RECT 420.400 64.300 421.200 64.400 ;
        RECT 436.400 64.300 437.200 64.400 ;
        RECT 441.200 64.300 442.000 64.400 ;
        RECT 420.400 63.700 442.000 64.300 ;
        RECT 420.400 63.600 421.200 63.700 ;
        RECT 436.400 63.600 437.200 63.700 ;
        RECT 441.200 63.600 442.000 63.700 ;
        RECT 492.400 64.300 493.200 64.400 ;
        RECT 500.400 64.300 501.200 64.400 ;
        RECT 503.600 64.300 504.400 64.400 ;
        RECT 492.400 63.700 504.400 64.300 ;
        RECT 492.400 63.600 493.200 63.700 ;
        RECT 500.400 63.600 501.200 63.700 ;
        RECT 503.600 63.600 504.400 63.700 ;
        RECT 540.400 64.300 541.200 64.400 ;
        RECT 542.000 64.300 542.800 64.400 ;
        RECT 540.400 63.700 542.800 64.300 ;
        RECT 540.400 63.600 541.200 63.700 ;
        RECT 542.000 63.600 542.800 63.700 ;
        RECT 348.400 62.300 349.200 62.400 ;
        RECT 298.900 61.700 349.200 62.300 ;
        RECT 206.000 61.600 206.800 61.700 ;
        RECT 348.400 61.600 349.200 61.700 ;
        RECT 412.400 62.300 413.200 62.400 ;
        RECT 473.200 62.300 474.000 62.400 ;
        RECT 478.000 62.300 478.800 62.400 ;
        RECT 412.400 61.700 478.800 62.300 ;
        RECT 412.400 61.600 413.200 61.700 ;
        RECT 473.200 61.600 474.000 61.700 ;
        RECT 478.000 61.600 478.800 61.700 ;
        RECT 9.200 60.300 10.000 60.400 ;
        RECT 33.200 60.300 34.000 60.400 ;
        RECT 9.200 59.700 34.000 60.300 ;
        RECT 9.200 59.600 10.000 59.700 ;
        RECT 33.200 59.600 34.000 59.700 ;
        RECT 127.600 60.300 128.400 60.400 ;
        RECT 129.200 60.300 130.000 60.400 ;
        RECT 146.800 60.300 147.600 60.400 ;
        RECT 150.000 60.300 150.800 60.400 ;
        RECT 127.600 59.700 134.700 60.300 ;
        RECT 127.600 59.600 128.400 59.700 ;
        RECT 129.200 59.600 130.000 59.700 ;
        RECT 2.800 58.300 3.600 58.400 ;
        RECT 10.800 58.300 11.600 58.400 ;
        RECT 25.200 58.300 26.000 58.400 ;
        RECT 2.800 57.700 26.000 58.300 ;
        RECT 2.800 57.600 3.600 57.700 ;
        RECT 10.800 57.600 11.600 57.700 ;
        RECT 25.200 57.600 26.000 57.700 ;
        RECT 30.000 58.300 30.800 58.400 ;
        RECT 41.200 58.300 42.000 58.400 ;
        RECT 86.000 58.300 86.800 58.400 ;
        RECT 30.000 57.700 86.800 58.300 ;
        RECT 30.000 57.600 30.800 57.700 ;
        RECT 41.200 57.600 42.000 57.700 ;
        RECT 86.000 57.600 86.800 57.700 ;
        RECT 97.200 58.300 98.000 58.400 ;
        RECT 132.400 58.300 133.200 58.400 ;
        RECT 97.200 57.700 133.200 58.300 ;
        RECT 134.100 58.300 134.700 59.700 ;
        RECT 146.800 59.700 150.800 60.300 ;
        RECT 146.800 59.600 147.600 59.700 ;
        RECT 150.000 59.600 150.800 59.700 ;
        RECT 156.400 60.300 157.200 60.400 ;
        RECT 166.000 60.300 166.800 60.400 ;
        RECT 156.400 59.700 166.800 60.300 ;
        RECT 156.400 59.600 157.200 59.700 ;
        RECT 166.000 59.600 166.800 59.700 ;
        RECT 273.200 60.300 274.000 60.400 ;
        RECT 278.000 60.300 278.800 60.400 ;
        RECT 273.200 59.700 278.800 60.300 ;
        RECT 273.200 59.600 274.000 59.700 ;
        RECT 278.000 59.600 278.800 59.700 ;
        RECT 281.200 60.300 282.000 60.400 ;
        RECT 287.600 60.300 288.400 60.400 ;
        RECT 281.200 59.700 288.400 60.300 ;
        RECT 281.200 59.600 282.000 59.700 ;
        RECT 287.600 59.600 288.400 59.700 ;
        RECT 300.400 60.300 301.200 60.400 ;
        RECT 342.000 60.300 342.800 60.400 ;
        RECT 300.400 59.700 342.800 60.300 ;
        RECT 300.400 59.600 301.200 59.700 ;
        RECT 342.000 59.600 342.800 59.700 ;
        RECT 380.400 60.300 381.200 60.400 ;
        RECT 390.000 60.300 390.800 60.400 ;
        RECT 401.200 60.300 402.000 60.400 ;
        RECT 380.400 59.700 402.000 60.300 ;
        RECT 380.400 59.600 381.200 59.700 ;
        RECT 390.000 59.600 390.800 59.700 ;
        RECT 401.200 59.600 402.000 59.700 ;
        RECT 422.000 60.300 422.800 60.400 ;
        RECT 423.600 60.300 424.400 60.400 ;
        RECT 450.800 60.300 451.600 60.400 ;
        RECT 422.000 59.700 451.600 60.300 ;
        RECT 422.000 59.600 422.800 59.700 ;
        RECT 423.600 59.600 424.400 59.700 ;
        RECT 450.800 59.600 451.600 59.700 ;
        RECT 143.600 58.300 144.400 58.400 ;
        RECT 134.100 57.700 144.400 58.300 ;
        RECT 97.200 57.600 98.000 57.700 ;
        RECT 132.400 57.600 133.200 57.700 ;
        RECT 143.600 57.600 144.400 57.700 ;
        RECT 202.800 58.300 203.600 58.400 ;
        RECT 215.600 58.300 216.400 58.400 ;
        RECT 233.200 58.300 234.000 58.400 ;
        RECT 202.800 57.700 234.000 58.300 ;
        RECT 202.800 57.600 203.600 57.700 ;
        RECT 215.600 57.600 216.400 57.700 ;
        RECT 233.200 57.600 234.000 57.700 ;
        RECT 239.600 58.300 240.400 58.400 ;
        RECT 242.800 58.300 243.600 58.400 ;
        RECT 260.400 58.300 261.200 58.400 ;
        RECT 239.600 57.700 261.200 58.300 ;
        RECT 239.600 57.600 240.400 57.700 ;
        RECT 242.800 57.600 243.600 57.700 ;
        RECT 260.400 57.600 261.200 57.700 ;
        RECT 266.800 58.300 267.600 58.400 ;
        RECT 278.000 58.300 278.800 58.400 ;
        RECT 266.800 57.700 278.800 58.300 ;
        RECT 266.800 57.600 267.600 57.700 ;
        RECT 278.000 57.600 278.800 57.700 ;
        RECT 281.200 58.300 282.000 58.400 ;
        RECT 375.600 58.300 376.400 58.400 ;
        RECT 281.200 57.700 376.400 58.300 ;
        RECT 281.200 57.600 282.000 57.700 ;
        RECT 375.600 57.600 376.400 57.700 ;
        RECT 434.800 58.300 435.600 58.400 ;
        RECT 439.600 58.300 440.400 58.400 ;
        RECT 452.400 58.300 453.200 58.400 ;
        RECT 434.800 57.700 453.200 58.300 ;
        RECT 434.800 57.600 435.600 57.700 ;
        RECT 439.600 57.600 440.400 57.700 ;
        RECT 452.400 57.600 453.200 57.700 ;
        RECT 455.600 58.300 456.400 58.400 ;
        RECT 460.400 58.300 461.200 58.400 ;
        RECT 455.600 57.700 461.200 58.300 ;
        RECT 455.600 57.600 456.400 57.700 ;
        RECT 460.400 57.600 461.200 57.700 ;
        RECT 479.600 58.300 480.400 58.400 ;
        RECT 489.200 58.300 490.000 58.400 ;
        RECT 479.600 57.700 490.000 58.300 ;
        RECT 479.600 57.600 480.400 57.700 ;
        RECT 489.200 57.600 490.000 57.700 ;
        RECT 490.800 58.300 491.600 58.400 ;
        RECT 495.600 58.300 496.400 58.400 ;
        RECT 522.800 58.300 523.600 58.400 ;
        RECT 490.800 57.700 523.600 58.300 ;
        RECT 490.800 57.600 491.600 57.700 ;
        RECT 495.600 57.600 496.400 57.700 ;
        RECT 522.800 57.600 523.600 57.700 ;
        RECT 551.600 58.300 552.400 58.400 ;
        RECT 562.800 58.300 563.600 58.400 ;
        RECT 551.600 57.700 563.600 58.300 ;
        RECT 551.600 57.600 552.400 57.700 ;
        RECT 562.800 57.600 563.600 57.700 ;
        RECT 28.400 56.300 29.200 56.400 ;
        RECT 36.400 56.300 37.200 56.400 ;
        RECT 28.400 55.700 37.200 56.300 ;
        RECT 28.400 55.600 29.200 55.700 ;
        RECT 36.400 55.600 37.200 55.700 ;
        RECT 38.000 56.300 38.800 56.400 ;
        RECT 54.000 56.300 54.800 56.400 ;
        RECT 38.000 55.700 54.800 56.300 ;
        RECT 38.000 55.600 38.800 55.700 ;
        RECT 54.000 55.600 54.800 55.700 ;
        RECT 62.000 56.300 62.800 56.400 ;
        RECT 66.800 56.300 67.600 56.400 ;
        RECT 62.000 55.700 67.600 56.300 ;
        RECT 62.000 55.600 62.800 55.700 ;
        RECT 66.800 55.600 67.600 55.700 ;
        RECT 78.000 56.300 78.800 56.400 ;
        RECT 81.200 56.300 82.000 56.400 ;
        RECT 78.000 55.700 82.000 56.300 ;
        RECT 78.000 55.600 78.800 55.700 ;
        RECT 81.200 55.600 82.000 55.700 ;
        RECT 86.000 56.300 86.800 56.400 ;
        RECT 110.000 56.300 110.800 56.400 ;
        RECT 116.400 56.300 117.200 56.400 ;
        RECT 86.000 55.700 117.200 56.300 ;
        RECT 86.000 55.600 86.800 55.700 ;
        RECT 110.000 55.600 110.800 55.700 ;
        RECT 116.400 55.600 117.200 55.700 ;
        RECT 130.800 56.300 131.600 56.400 ;
        RECT 151.600 56.300 152.400 56.400 ;
        RECT 130.800 55.700 152.400 56.300 ;
        RECT 130.800 55.600 131.600 55.700 ;
        RECT 151.600 55.600 152.400 55.700 ;
        RECT 217.200 56.300 218.000 56.400 ;
        RECT 223.600 56.300 224.400 56.400 ;
        RECT 241.200 56.300 242.000 56.400 ;
        RECT 217.200 55.700 242.000 56.300 ;
        RECT 217.200 55.600 218.000 55.700 ;
        RECT 223.600 55.600 224.400 55.700 ;
        RECT 241.200 55.600 242.000 55.700 ;
        RECT 276.400 56.300 277.200 56.400 ;
        RECT 300.400 56.300 301.200 56.400 ;
        RECT 276.400 55.700 301.200 56.300 ;
        RECT 276.400 55.600 277.200 55.700 ;
        RECT 300.400 55.600 301.200 55.700 ;
        RECT 306.800 56.300 307.600 56.400 ;
        RECT 316.400 56.300 317.200 56.400 ;
        RECT 306.800 55.700 317.200 56.300 ;
        RECT 306.800 55.600 307.600 55.700 ;
        RECT 316.400 55.600 317.200 55.700 ;
        RECT 326.000 56.300 326.800 56.400 ;
        RECT 338.800 56.300 339.600 56.400 ;
        RECT 348.400 56.300 349.200 56.400 ;
        RECT 326.000 55.700 337.900 56.300 ;
        RECT 326.000 55.600 326.800 55.700 ;
        RECT 12.400 54.300 13.200 54.400 ;
        RECT 23.600 54.300 24.400 54.400 ;
        RECT 12.400 53.700 24.400 54.300 ;
        RECT 12.400 53.600 13.200 53.700 ;
        RECT 23.600 53.600 24.400 53.700 ;
        RECT 34.800 54.300 35.600 54.400 ;
        RECT 89.200 54.300 90.000 54.400 ;
        RECT 95.600 54.300 96.400 54.400 ;
        RECT 102.000 54.300 102.800 54.400 ;
        RECT 34.800 53.700 102.800 54.300 ;
        RECT 34.800 53.600 35.600 53.700 ;
        RECT 89.200 53.600 90.000 53.700 ;
        RECT 95.600 53.600 96.400 53.700 ;
        RECT 102.000 53.600 102.800 53.700 ;
        RECT 111.600 54.300 112.400 54.400 ;
        RECT 122.800 54.300 123.600 54.400 ;
        RECT 111.600 53.700 123.600 54.300 ;
        RECT 111.600 53.600 112.400 53.700 ;
        RECT 122.800 53.600 123.600 53.700 ;
        RECT 126.000 54.300 126.800 54.400 ;
        RECT 175.600 54.300 176.400 54.400 ;
        RECT 126.000 53.700 176.400 54.300 ;
        RECT 126.000 53.600 126.800 53.700 ;
        RECT 175.600 53.600 176.400 53.700 ;
        RECT 198.000 54.300 198.800 54.400 ;
        RECT 209.200 54.300 210.000 54.400 ;
        RECT 198.000 53.700 210.000 54.300 ;
        RECT 198.000 53.600 198.800 53.700 ;
        RECT 209.200 53.600 210.000 53.700 ;
        RECT 220.400 54.300 221.200 54.400 ;
        RECT 250.800 54.300 251.600 54.400 ;
        RECT 255.600 54.300 256.400 54.400 ;
        RECT 220.400 53.700 256.400 54.300 ;
        RECT 220.400 53.600 221.200 53.700 ;
        RECT 250.800 53.600 251.600 53.700 ;
        RECT 255.600 53.600 256.400 53.700 ;
        RECT 258.800 54.300 259.600 54.400 ;
        RECT 281.200 54.300 282.000 54.400 ;
        RECT 258.800 53.700 282.000 54.300 ;
        RECT 258.800 53.600 259.600 53.700 ;
        RECT 281.200 53.600 282.000 53.700 ;
        RECT 282.800 54.300 283.600 54.400 ;
        RECT 292.400 54.300 293.200 54.400 ;
        RECT 282.800 53.700 293.200 54.300 ;
        RECT 282.800 53.600 283.600 53.700 ;
        RECT 292.400 53.600 293.200 53.700 ;
        RECT 300.400 53.600 301.200 54.400 ;
        RECT 303.600 54.300 304.400 54.400 ;
        RECT 305.200 54.300 306.000 54.400 ;
        RECT 303.600 53.700 306.000 54.300 ;
        RECT 303.600 53.600 304.400 53.700 ;
        RECT 305.200 53.600 306.000 53.700 ;
        RECT 308.400 54.300 309.200 54.400 ;
        RECT 314.800 54.300 315.600 54.400 ;
        RECT 322.800 54.300 323.600 54.400 ;
        RECT 308.400 53.700 323.600 54.300 ;
        RECT 337.300 54.300 337.900 55.700 ;
        RECT 338.800 55.700 349.200 56.300 ;
        RECT 338.800 55.600 339.600 55.700 ;
        RECT 348.400 55.600 349.200 55.700 ;
        RECT 369.200 56.300 370.000 56.400 ;
        RECT 385.200 56.300 386.000 56.400 ;
        RECT 396.400 56.300 397.200 56.400 ;
        RECT 412.400 56.300 413.200 56.400 ;
        RECT 369.200 55.700 413.200 56.300 ;
        RECT 369.200 55.600 370.000 55.700 ;
        RECT 385.200 55.600 386.000 55.700 ;
        RECT 396.400 55.600 397.200 55.700 ;
        RECT 412.400 55.600 413.200 55.700 ;
        RECT 415.600 56.300 416.400 56.400 ;
        RECT 433.200 56.300 434.000 56.400 ;
        RECT 438.000 56.300 438.800 56.400 ;
        RECT 415.600 55.700 438.800 56.300 ;
        RECT 415.600 55.600 416.400 55.700 ;
        RECT 433.200 55.600 434.000 55.700 ;
        RECT 438.000 55.600 438.800 55.700 ;
        RECT 457.200 56.300 458.000 56.400 ;
        RECT 470.000 56.300 470.800 56.400 ;
        RECT 457.200 55.700 470.800 56.300 ;
        RECT 457.200 55.600 458.000 55.700 ;
        RECT 470.000 55.600 470.800 55.700 ;
        RECT 486.000 56.300 486.800 56.400 ;
        RECT 508.400 56.300 509.200 56.400 ;
        RECT 511.600 56.300 512.400 56.400 ;
        RECT 486.000 55.700 512.400 56.300 ;
        RECT 486.000 55.600 486.800 55.700 ;
        RECT 508.400 55.600 509.200 55.700 ;
        RECT 511.600 55.600 512.400 55.700 ;
        RECT 340.400 54.300 341.200 54.400 ;
        RECT 337.300 53.700 341.200 54.300 ;
        RECT 308.400 53.600 309.200 53.700 ;
        RECT 314.800 53.600 315.600 53.700 ;
        RECT 322.800 53.600 323.600 53.700 ;
        RECT 340.400 53.600 341.200 53.700 ;
        RECT 385.200 54.300 386.000 54.400 ;
        RECT 399.600 54.300 400.400 54.400 ;
        RECT 385.200 53.700 400.400 54.300 ;
        RECT 385.200 53.600 386.000 53.700 ;
        RECT 399.600 53.600 400.400 53.700 ;
        RECT 434.800 53.600 435.600 54.400 ;
        RECT 449.200 54.300 450.000 54.400 ;
        RECT 458.800 54.300 459.600 54.400 ;
        RECT 449.200 53.700 459.600 54.300 ;
        RECT 449.200 53.600 450.000 53.700 ;
        RECT 458.800 53.600 459.600 53.700 ;
        RECT 463.600 54.300 464.400 54.400 ;
        RECT 468.400 54.300 469.200 54.400 ;
        RECT 471.600 54.300 472.400 54.400 ;
        RECT 463.600 53.700 472.400 54.300 ;
        RECT 463.600 53.600 464.400 53.700 ;
        RECT 468.400 53.600 469.200 53.700 ;
        RECT 471.600 53.600 472.400 53.700 ;
        RECT 486.000 54.300 486.800 54.400 ;
        RECT 494.000 54.300 494.800 54.400 ;
        RECT 486.000 53.700 494.800 54.300 ;
        RECT 486.000 53.600 486.800 53.700 ;
        RECT 494.000 53.600 494.800 53.700 ;
        RECT 497.200 54.300 498.000 54.400 ;
        RECT 500.400 54.300 501.200 54.400 ;
        RECT 497.200 53.700 501.200 54.300 ;
        RECT 497.200 53.600 498.000 53.700 ;
        RECT 500.400 53.600 501.200 53.700 ;
        RECT 508.400 53.600 509.200 54.400 ;
        RECT 559.600 54.300 560.400 54.400 ;
        RECT 572.400 54.300 573.200 54.400 ;
        RECT 559.600 53.700 573.200 54.300 ;
        RECT 559.600 53.600 560.400 53.700 ;
        RECT 572.400 53.600 573.200 53.700 ;
        RECT 1.200 52.300 2.000 52.400 ;
        RECT 9.200 52.300 10.000 52.400 ;
        RECT 1.200 51.700 10.000 52.300 ;
        RECT 1.200 51.600 2.000 51.700 ;
        RECT 9.200 51.600 10.000 51.700 ;
        RECT 14.000 52.300 14.800 52.400 ;
        RECT 20.400 52.300 21.200 52.400 ;
        RECT 14.000 51.700 21.200 52.300 ;
        RECT 14.000 51.600 14.800 51.700 ;
        RECT 20.400 51.600 21.200 51.700 ;
        RECT 28.400 52.300 29.200 52.400 ;
        RECT 38.000 52.300 38.800 52.400 ;
        RECT 28.400 51.700 38.800 52.300 ;
        RECT 28.400 51.600 29.200 51.700 ;
        RECT 38.000 51.600 38.800 51.700 ;
        RECT 39.600 52.300 40.400 52.400 ;
        RECT 68.400 52.300 69.200 52.400 ;
        RECT 39.600 51.700 69.200 52.300 ;
        RECT 39.600 51.600 40.400 51.700 ;
        RECT 68.400 51.600 69.200 51.700 ;
        RECT 74.800 52.300 75.600 52.400 ;
        RECT 78.000 52.300 78.800 52.400 ;
        RECT 74.800 51.700 78.800 52.300 ;
        RECT 74.800 51.600 75.600 51.700 ;
        RECT 78.000 51.600 78.800 51.700 ;
        RECT 90.800 52.300 91.600 52.400 ;
        RECT 114.800 52.300 115.600 52.400 ;
        RECT 90.800 51.700 115.600 52.300 ;
        RECT 90.800 51.600 91.600 51.700 ;
        RECT 114.800 51.600 115.600 51.700 ;
        RECT 118.000 52.300 118.800 52.400 ;
        RECT 146.800 52.300 147.600 52.400 ;
        RECT 118.000 51.700 147.600 52.300 ;
        RECT 118.000 51.600 118.800 51.700 ;
        RECT 146.800 51.600 147.600 51.700 ;
        RECT 172.400 52.300 173.200 52.400 ;
        RECT 182.000 52.300 182.800 52.400 ;
        RECT 172.400 51.700 182.800 52.300 ;
        RECT 172.400 51.600 173.200 51.700 ;
        RECT 182.000 51.600 182.800 51.700 ;
        RECT 217.200 52.300 218.000 52.400 ;
        RECT 230.000 52.300 230.800 52.400 ;
        RECT 234.800 52.300 235.600 52.400 ;
        RECT 217.200 51.700 235.600 52.300 ;
        RECT 217.200 51.600 218.000 51.700 ;
        RECT 230.000 51.600 230.800 51.700 ;
        RECT 234.800 51.600 235.600 51.700 ;
        RECT 252.400 52.300 253.200 52.400 ;
        RECT 258.800 52.300 259.600 52.400 ;
        RECT 263.600 52.300 264.400 52.400 ;
        RECT 252.400 51.700 264.400 52.300 ;
        RECT 252.400 51.600 253.200 51.700 ;
        RECT 258.800 51.600 259.600 51.700 ;
        RECT 263.600 51.600 264.400 51.700 ;
        RECT 276.400 52.300 277.200 52.400 ;
        RECT 282.800 52.300 283.600 52.400 ;
        RECT 321.200 52.300 322.000 52.400 ;
        RECT 330.800 52.300 331.600 52.400 ;
        RECT 276.400 51.700 331.600 52.300 ;
        RECT 276.400 51.600 277.200 51.700 ;
        RECT 282.800 51.600 283.600 51.700 ;
        RECT 321.200 51.600 322.000 51.700 ;
        RECT 330.800 51.600 331.600 51.700 ;
        RECT 332.400 52.300 333.200 52.400 ;
        RECT 338.800 52.300 339.600 52.400 ;
        RECT 332.400 51.700 339.600 52.300 ;
        RECT 332.400 51.600 333.200 51.700 ;
        RECT 338.800 51.600 339.600 51.700 ;
        RECT 346.800 52.300 347.600 52.400 ;
        RECT 356.400 52.300 357.200 52.400 ;
        RECT 346.800 51.700 357.200 52.300 ;
        RECT 346.800 51.600 347.600 51.700 ;
        RECT 356.400 51.600 357.200 51.700 ;
        RECT 438.000 52.300 438.800 52.400 ;
        RECT 481.200 52.300 482.000 52.400 ;
        RECT 487.600 52.300 488.400 52.400 ;
        RECT 511.600 52.300 512.400 52.400 ;
        RECT 521.200 52.300 522.000 52.400 ;
        RECT 438.000 51.700 522.000 52.300 ;
        RECT 438.000 51.600 438.800 51.700 ;
        RECT 481.200 51.600 482.000 51.700 ;
        RECT 487.600 51.600 488.400 51.700 ;
        RECT 511.600 51.600 512.400 51.700 ;
        RECT 521.200 51.600 522.000 51.700 ;
        RECT 535.600 52.300 536.400 52.400 ;
        RECT 550.000 52.300 550.800 52.400 ;
        RECT 535.600 51.700 550.800 52.300 ;
        RECT 535.600 51.600 536.400 51.700 ;
        RECT 550.000 51.600 550.800 51.700 ;
        RECT 556.400 52.300 557.200 52.400 ;
        RECT 569.200 52.300 570.000 52.400 ;
        RECT 556.400 51.700 570.000 52.300 ;
        RECT 556.400 51.600 557.200 51.700 ;
        RECT 569.200 51.600 570.000 51.700 ;
        RECT 575.600 51.600 576.400 52.400 ;
        RECT 18.800 50.300 19.600 50.400 ;
        RECT 23.600 50.300 24.400 50.400 ;
        RECT 34.800 50.300 35.600 50.400 ;
        RECT 18.800 49.700 35.600 50.300 ;
        RECT 18.800 49.600 19.600 49.700 ;
        RECT 23.600 49.600 24.400 49.700 ;
        RECT 34.800 49.600 35.600 49.700 ;
        RECT 49.200 50.300 50.000 50.400 ;
        RECT 50.800 50.300 51.600 50.400 ;
        RECT 49.200 49.700 51.600 50.300 ;
        RECT 49.200 49.600 50.000 49.700 ;
        RECT 50.800 49.600 51.600 49.700 ;
        RECT 55.600 50.300 56.400 50.400 ;
        RECT 84.400 50.300 85.200 50.400 ;
        RECT 98.800 50.300 99.600 50.400 ;
        RECT 105.200 50.300 106.000 50.400 ;
        RECT 129.200 50.300 130.000 50.400 ;
        RECT 55.600 49.700 130.000 50.300 ;
        RECT 55.600 49.600 56.400 49.700 ;
        RECT 84.400 49.600 85.200 49.700 ;
        RECT 98.800 49.600 99.600 49.700 ;
        RECT 105.200 49.600 106.000 49.700 ;
        RECT 129.200 49.600 130.000 49.700 ;
        RECT 255.600 50.300 256.400 50.400 ;
        RECT 278.000 50.300 278.800 50.400 ;
        RECT 255.600 49.700 278.800 50.300 ;
        RECT 255.600 49.600 256.400 49.700 ;
        RECT 278.000 49.600 278.800 49.700 ;
        RECT 297.200 49.600 298.000 50.400 ;
        RECT 337.200 50.300 338.000 50.400 ;
        RECT 343.600 50.300 344.400 50.400 ;
        RECT 350.000 50.300 350.800 50.400 ;
        RECT 337.200 49.700 350.800 50.300 ;
        RECT 337.200 49.600 338.000 49.700 ;
        RECT 343.600 49.600 344.400 49.700 ;
        RECT 350.000 49.600 350.800 49.700 ;
        RECT 430.000 50.300 430.800 50.400 ;
        RECT 457.200 50.300 458.000 50.400 ;
        RECT 465.200 50.300 466.000 50.400 ;
        RECT 430.000 49.700 466.000 50.300 ;
        RECT 430.000 49.600 430.800 49.700 ;
        RECT 457.200 49.600 458.000 49.700 ;
        RECT 465.200 49.600 466.000 49.700 ;
        RECT 468.400 50.300 469.200 50.400 ;
        RECT 476.400 50.300 477.200 50.400 ;
        RECT 468.400 49.700 477.200 50.300 ;
        RECT 468.400 49.600 469.200 49.700 ;
        RECT 476.400 49.600 477.200 49.700 ;
        RECT 492.400 50.300 493.200 50.400 ;
        RECT 495.600 50.300 496.400 50.400 ;
        RECT 503.600 50.300 504.400 50.400 ;
        RECT 492.400 49.700 504.400 50.300 ;
        RECT 492.400 49.600 493.200 49.700 ;
        RECT 495.600 49.600 496.400 49.700 ;
        RECT 503.600 49.600 504.400 49.700 ;
        RECT 516.400 50.300 517.200 50.400 ;
        RECT 527.600 50.300 528.400 50.400 ;
        RECT 516.400 49.700 528.400 50.300 ;
        RECT 516.400 49.600 517.200 49.700 ;
        RECT 527.600 49.600 528.400 49.700 ;
        RECT 550.000 50.300 550.800 50.400 ;
        RECT 556.400 50.300 557.200 50.400 ;
        RECT 550.000 49.700 557.200 50.300 ;
        RECT 550.000 49.600 550.800 49.700 ;
        RECT 556.400 49.600 557.200 49.700 ;
        RECT 42.800 48.300 43.600 48.400 ;
        RECT 76.400 48.300 77.200 48.400 ;
        RECT 42.800 47.700 77.200 48.300 ;
        RECT 42.800 47.600 43.600 47.700 ;
        RECT 76.400 47.600 77.200 47.700 ;
        RECT 100.400 48.300 101.200 48.400 ;
        RECT 124.400 48.300 125.200 48.400 ;
        RECT 100.400 47.700 125.200 48.300 ;
        RECT 100.400 47.600 101.200 47.700 ;
        RECT 124.400 47.600 125.200 47.700 ;
        RECT 193.200 48.300 194.000 48.400 ;
        RECT 265.200 48.300 266.000 48.400 ;
        RECT 193.200 47.700 266.000 48.300 ;
        RECT 193.200 47.600 194.000 47.700 ;
        RECT 265.200 47.600 266.000 47.700 ;
        RECT 268.400 48.300 269.200 48.400 ;
        RECT 327.600 48.300 328.400 48.400 ;
        RECT 348.400 48.300 349.200 48.400 ;
        RECT 268.400 47.700 349.200 48.300 ;
        RECT 268.400 47.600 269.200 47.700 ;
        RECT 327.600 47.600 328.400 47.700 ;
        RECT 348.400 47.600 349.200 47.700 ;
        RECT 388.400 48.300 389.200 48.400 ;
        RECT 394.800 48.300 395.600 48.400 ;
        RECT 417.200 48.300 418.000 48.400 ;
        RECT 388.400 47.700 418.000 48.300 ;
        RECT 388.400 47.600 389.200 47.700 ;
        RECT 394.800 47.600 395.600 47.700 ;
        RECT 417.200 47.600 418.000 47.700 ;
        RECT 452.400 48.300 453.200 48.400 ;
        RECT 463.600 48.300 464.400 48.400 ;
        RECT 484.400 48.300 485.200 48.400 ;
        RECT 452.400 47.700 485.200 48.300 ;
        RECT 452.400 47.600 453.200 47.700 ;
        RECT 463.600 47.600 464.400 47.700 ;
        RECT 484.400 47.600 485.200 47.700 ;
        RECT 502.000 48.300 502.800 48.400 ;
        RECT 510.000 48.300 510.800 48.400 ;
        RECT 502.000 47.700 510.800 48.300 ;
        RECT 502.000 47.600 502.800 47.700 ;
        RECT 510.000 47.600 510.800 47.700 ;
        RECT 87.600 46.300 88.400 46.400 ;
        RECT 156.400 46.300 157.200 46.400 ;
        RECT 174.000 46.300 174.800 46.400 ;
        RECT 199.600 46.300 200.400 46.400 ;
        RECT 87.600 45.700 200.400 46.300 ;
        RECT 87.600 45.600 88.400 45.700 ;
        RECT 156.400 45.600 157.200 45.700 ;
        RECT 174.000 45.600 174.800 45.700 ;
        RECT 199.600 45.600 200.400 45.700 ;
        RECT 207.600 46.300 208.400 46.400 ;
        RECT 210.800 46.300 211.600 46.400 ;
        RECT 270.000 46.300 270.800 46.400 ;
        RECT 207.600 45.700 270.800 46.300 ;
        RECT 207.600 45.600 208.400 45.700 ;
        RECT 210.800 45.600 211.600 45.700 ;
        RECT 270.000 45.600 270.800 45.700 ;
        RECT 278.000 46.300 278.800 46.400 ;
        RECT 313.200 46.300 314.000 46.400 ;
        RECT 278.000 45.700 314.000 46.300 ;
        RECT 278.000 45.600 278.800 45.700 ;
        RECT 313.200 45.600 314.000 45.700 ;
        RECT 447.600 46.300 448.400 46.400 ;
        RECT 450.800 46.300 451.600 46.400 ;
        RECT 447.600 45.700 451.600 46.300 ;
        RECT 447.600 45.600 448.400 45.700 ;
        RECT 450.800 45.600 451.600 45.700 ;
        RECT 177.200 44.300 178.000 44.400 ;
        RECT 252.400 44.300 253.200 44.400 ;
        RECT 177.200 43.700 253.200 44.300 ;
        RECT 177.200 43.600 178.000 43.700 ;
        RECT 252.400 43.600 253.200 43.700 ;
        RECT 265.200 44.300 266.000 44.400 ;
        RECT 402.800 44.300 403.600 44.400 ;
        RECT 265.200 43.700 403.600 44.300 ;
        RECT 265.200 43.600 266.000 43.700 ;
        RECT 402.800 43.600 403.600 43.700 ;
        RECT 436.400 44.300 437.200 44.400 ;
        RECT 470.000 44.300 470.800 44.400 ;
        RECT 436.400 43.700 470.800 44.300 ;
        RECT 436.400 43.600 437.200 43.700 ;
        RECT 470.000 43.600 470.800 43.700 ;
        RECT 543.600 44.300 544.400 44.400 ;
        RECT 553.200 44.300 554.000 44.400 ;
        RECT 558.000 44.300 558.800 44.400 ;
        RECT 543.600 43.700 558.800 44.300 ;
        RECT 543.600 43.600 544.400 43.700 ;
        RECT 553.200 43.600 554.000 43.700 ;
        RECT 558.000 43.600 558.800 43.700 ;
        RECT 153.200 42.300 154.000 42.400 ;
        RECT 198.000 42.300 198.800 42.400 ;
        RECT 153.200 41.700 198.800 42.300 ;
        RECT 153.200 41.600 154.000 41.700 ;
        RECT 198.000 41.600 198.800 41.700 ;
        RECT 287.600 42.300 288.400 42.400 ;
        RECT 318.000 42.300 318.800 42.400 ;
        RECT 356.400 42.300 357.200 42.400 ;
        RECT 287.600 41.700 357.200 42.300 ;
        RECT 287.600 41.600 288.400 41.700 ;
        RECT 318.000 41.600 318.800 41.700 ;
        RECT 356.400 41.600 357.200 41.700 ;
        RECT 175.600 40.300 176.400 40.400 ;
        RECT 183.600 40.300 184.400 40.400 ;
        RECT 175.600 39.700 184.400 40.300 ;
        RECT 175.600 39.600 176.400 39.700 ;
        RECT 183.600 39.600 184.400 39.700 ;
        RECT 254.000 40.300 254.800 40.400 ;
        RECT 316.400 40.300 317.200 40.400 ;
        RECT 254.000 39.700 317.200 40.300 ;
        RECT 254.000 39.600 254.800 39.700 ;
        RECT 316.400 39.600 317.200 39.700 ;
        RECT 318.000 40.300 318.800 40.400 ;
        RECT 329.200 40.300 330.000 40.400 ;
        RECT 318.000 39.700 330.000 40.300 ;
        RECT 318.000 39.600 318.800 39.700 ;
        RECT 329.200 39.600 330.000 39.700 ;
        RECT 418.800 40.300 419.600 40.400 ;
        RECT 471.600 40.300 472.400 40.400 ;
        RECT 494.000 40.300 494.800 40.400 ;
        RECT 418.800 39.700 441.900 40.300 ;
        RECT 418.800 39.600 419.600 39.700 ;
        RECT 68.400 38.300 69.200 38.400 ;
        RECT 73.200 38.300 74.000 38.400 ;
        RECT 68.400 37.700 74.000 38.300 ;
        RECT 68.400 37.600 69.200 37.700 ;
        RECT 73.200 37.600 74.000 37.700 ;
        RECT 98.800 38.300 99.600 38.400 ;
        RECT 158.000 38.300 158.800 38.400 ;
        RECT 98.800 37.700 158.800 38.300 ;
        RECT 98.800 37.600 99.600 37.700 ;
        RECT 158.000 37.600 158.800 37.700 ;
        RECT 164.400 38.300 165.200 38.400 ;
        RECT 218.800 38.300 219.600 38.400 ;
        RECT 164.400 37.700 219.600 38.300 ;
        RECT 164.400 37.600 165.200 37.700 ;
        RECT 218.800 37.600 219.600 37.700 ;
        RECT 247.600 38.300 248.400 38.400 ;
        RECT 266.800 38.300 267.600 38.400 ;
        RECT 303.600 38.300 304.400 38.400 ;
        RECT 247.600 37.700 304.400 38.300 ;
        RECT 247.600 37.600 248.400 37.700 ;
        RECT 266.800 37.600 267.600 37.700 ;
        RECT 303.600 37.600 304.400 37.700 ;
        RECT 350.000 38.300 350.800 38.400 ;
        RECT 354.800 38.300 355.600 38.400 ;
        RECT 350.000 37.700 355.600 38.300 ;
        RECT 350.000 37.600 350.800 37.700 ;
        RECT 354.800 37.600 355.600 37.700 ;
        RECT 425.200 38.300 426.000 38.400 ;
        RECT 431.600 38.300 432.400 38.400 ;
        RECT 425.200 37.700 432.400 38.300 ;
        RECT 441.300 38.300 441.900 39.700 ;
        RECT 471.600 39.700 494.800 40.300 ;
        RECT 471.600 39.600 472.400 39.700 ;
        RECT 494.000 39.600 494.800 39.700 ;
        RECT 506.800 40.300 507.600 40.400 ;
        RECT 519.600 40.300 520.400 40.400 ;
        RECT 506.800 39.700 520.400 40.300 ;
        RECT 506.800 39.600 507.600 39.700 ;
        RECT 519.600 39.600 520.400 39.700 ;
        RECT 458.800 38.300 459.600 38.400 ;
        RECT 441.300 37.700 459.600 38.300 ;
        RECT 425.200 37.600 426.000 37.700 ;
        RECT 431.600 37.600 432.400 37.700 ;
        RECT 458.800 37.600 459.600 37.700 ;
        RECT 460.400 38.300 461.200 38.400 ;
        RECT 473.200 38.300 474.000 38.400 ;
        RECT 460.400 37.700 474.000 38.300 ;
        RECT 460.400 37.600 461.200 37.700 ;
        RECT 473.200 37.600 474.000 37.700 ;
        RECT 476.400 38.300 477.200 38.400 ;
        RECT 479.600 38.300 480.400 38.400 ;
        RECT 486.000 38.300 486.800 38.400 ;
        RECT 476.400 37.700 486.800 38.300 ;
        RECT 476.400 37.600 477.200 37.700 ;
        RECT 479.600 37.600 480.400 37.700 ;
        RECT 486.000 37.600 486.800 37.700 ;
        RECT 487.600 38.300 488.400 38.400 ;
        RECT 498.800 38.300 499.600 38.400 ;
        RECT 487.600 37.700 499.600 38.300 ;
        RECT 487.600 37.600 488.400 37.700 ;
        RECT 498.800 37.600 499.600 37.700 ;
        RECT 30.000 36.300 30.800 36.400 ;
        RECT 140.400 36.300 141.200 36.400 ;
        RECT 151.600 36.300 152.400 36.400 ;
        RECT 217.200 36.300 218.000 36.400 ;
        RECT 30.000 35.700 53.100 36.300 ;
        RECT 30.000 35.600 30.800 35.700 ;
        RECT 52.500 34.400 53.100 35.700 ;
        RECT 140.400 35.700 218.000 36.300 ;
        RECT 140.400 35.600 141.200 35.700 ;
        RECT 151.600 35.600 152.400 35.700 ;
        RECT 217.200 35.600 218.000 35.700 ;
        RECT 218.800 36.300 219.600 36.400 ;
        RECT 226.800 36.300 227.600 36.400 ;
        RECT 218.800 35.700 227.600 36.300 ;
        RECT 218.800 35.600 219.600 35.700 ;
        RECT 226.800 35.600 227.600 35.700 ;
        RECT 233.200 36.300 234.000 36.400 ;
        RECT 268.400 36.300 269.200 36.400 ;
        RECT 233.200 35.700 269.200 36.300 ;
        RECT 233.200 35.600 234.000 35.700 ;
        RECT 268.400 35.600 269.200 35.700 ;
        RECT 425.200 36.300 426.000 36.400 ;
        RECT 428.400 36.300 429.200 36.400 ;
        RECT 425.200 35.700 429.200 36.300 ;
        RECT 425.200 35.600 426.000 35.700 ;
        RECT 428.400 35.600 429.200 35.700 ;
        RECT 436.400 36.300 437.200 36.400 ;
        RECT 458.800 36.300 459.600 36.400 ;
        RECT 436.400 35.700 459.600 36.300 ;
        RECT 436.400 35.600 437.200 35.700 ;
        RECT 458.800 35.600 459.600 35.700 ;
        RECT 460.400 36.300 461.200 36.400 ;
        RECT 487.600 36.300 488.400 36.400 ;
        RECT 460.400 35.700 488.400 36.300 ;
        RECT 460.400 35.600 461.200 35.700 ;
        RECT 487.600 35.600 488.400 35.700 ;
        RECT 489.200 36.300 490.000 36.400 ;
        RECT 508.400 36.300 509.200 36.400 ;
        RECT 489.200 35.700 509.200 36.300 ;
        RECT 489.200 35.600 490.000 35.700 ;
        RECT 508.400 35.600 509.200 35.700 ;
        RECT 10.800 34.300 11.600 34.400 ;
        RECT 20.400 34.300 21.200 34.400 ;
        RECT 10.800 33.700 21.200 34.300 ;
        RECT 10.800 33.600 11.600 33.700 ;
        RECT 20.400 33.600 21.200 33.700 ;
        RECT 26.800 34.300 27.600 34.400 ;
        RECT 42.800 34.300 43.600 34.400 ;
        RECT 26.800 33.700 43.600 34.300 ;
        RECT 26.800 33.600 27.600 33.700 ;
        RECT 42.800 33.600 43.600 33.700 ;
        RECT 52.400 34.300 53.200 34.400 ;
        RECT 70.000 34.300 70.800 34.400 ;
        RECT 52.400 33.700 70.800 34.300 ;
        RECT 52.400 33.600 53.200 33.700 ;
        RECT 70.000 33.600 70.800 33.700 ;
        RECT 103.600 34.300 104.400 34.400 ;
        RECT 130.800 34.300 131.600 34.400 ;
        RECT 103.600 33.700 131.600 34.300 ;
        RECT 103.600 33.600 104.400 33.700 ;
        RECT 130.800 33.600 131.600 33.700 ;
        RECT 158.000 34.300 158.800 34.400 ;
        RECT 242.800 34.300 243.600 34.400 ;
        RECT 158.000 33.700 243.600 34.300 ;
        RECT 158.000 33.600 158.800 33.700 ;
        RECT 242.800 33.600 243.600 33.700 ;
        RECT 246.000 34.300 246.800 34.400 ;
        RECT 249.200 34.300 250.000 34.400 ;
        RECT 262.000 34.300 262.800 34.400 ;
        RECT 284.400 34.300 285.200 34.400 ;
        RECT 294.000 34.300 294.800 34.400 ;
        RECT 298.800 34.300 299.600 34.400 ;
        RECT 246.000 33.700 248.300 34.300 ;
        RECT 246.000 33.600 246.800 33.700 ;
        RECT 7.600 32.300 8.400 32.400 ;
        RECT 12.400 32.300 13.200 32.400 ;
        RECT 7.600 31.700 13.200 32.300 ;
        RECT 7.600 31.600 8.400 31.700 ;
        RECT 12.400 31.600 13.200 31.700 ;
        RECT 36.400 32.300 37.200 32.400 ;
        RECT 38.000 32.300 38.800 32.400 ;
        RECT 36.400 31.700 38.800 32.300 ;
        RECT 36.400 31.600 37.200 31.700 ;
        RECT 38.000 31.600 38.800 31.700 ;
        RECT 39.600 32.300 40.400 32.400 ;
        RECT 63.600 32.300 64.400 32.400 ;
        RECT 39.600 31.700 64.400 32.300 ;
        RECT 39.600 31.600 40.400 31.700 ;
        RECT 63.600 31.600 64.400 31.700 ;
        RECT 76.400 32.300 77.200 32.400 ;
        RECT 92.400 32.300 93.200 32.400 ;
        RECT 76.400 31.700 93.200 32.300 ;
        RECT 76.400 31.600 77.200 31.700 ;
        RECT 92.400 31.600 93.200 31.700 ;
        RECT 118.000 32.300 118.800 32.400 ;
        RECT 148.400 32.300 149.200 32.400 ;
        RECT 118.000 31.700 149.200 32.300 ;
        RECT 118.000 31.600 118.800 31.700 ;
        RECT 148.400 31.600 149.200 31.700 ;
        RECT 170.800 32.300 171.600 32.400 ;
        RECT 199.600 32.300 200.400 32.400 ;
        RECT 204.400 32.300 205.200 32.400 ;
        RECT 170.800 31.700 205.200 32.300 ;
        RECT 170.800 31.600 171.600 31.700 ;
        RECT 199.600 31.600 200.400 31.700 ;
        RECT 204.400 31.600 205.200 31.700 ;
        RECT 215.600 32.300 216.400 32.400 ;
        RECT 218.800 32.300 219.600 32.400 ;
        RECT 215.600 31.700 219.600 32.300 ;
        RECT 215.600 31.600 216.400 31.700 ;
        RECT 218.800 31.600 219.600 31.700 ;
        RECT 226.800 32.300 227.600 32.400 ;
        RECT 234.800 32.300 235.600 32.400 ;
        RECT 226.800 31.700 235.600 32.300 ;
        RECT 226.800 31.600 227.600 31.700 ;
        RECT 234.800 31.600 235.600 31.700 ;
        RECT 239.600 32.300 240.400 32.400 ;
        RECT 246.000 32.300 246.800 32.400 ;
        RECT 239.600 31.700 246.800 32.300 ;
        RECT 247.700 32.300 248.300 33.700 ;
        RECT 249.200 33.700 299.600 34.300 ;
        RECT 249.200 33.600 250.000 33.700 ;
        RECT 262.000 33.600 262.800 33.700 ;
        RECT 284.400 33.600 285.200 33.700 ;
        RECT 294.000 33.600 294.800 33.700 ;
        RECT 298.800 33.600 299.600 33.700 ;
        RECT 313.200 34.300 314.000 34.400 ;
        RECT 330.800 34.300 331.600 34.400 ;
        RECT 313.200 33.700 331.600 34.300 ;
        RECT 313.200 33.600 314.000 33.700 ;
        RECT 330.800 33.600 331.600 33.700 ;
        RECT 417.200 34.300 418.000 34.400 ;
        RECT 434.800 34.300 435.600 34.400 ;
        RECT 417.200 33.700 435.600 34.300 ;
        RECT 417.200 33.600 418.000 33.700 ;
        RECT 434.800 33.600 435.600 33.700 ;
        RECT 455.600 34.300 456.400 34.400 ;
        RECT 465.200 34.300 466.000 34.400 ;
        RECT 529.200 34.300 530.000 34.400 ;
        RECT 455.600 33.700 530.000 34.300 ;
        RECT 455.600 33.600 456.400 33.700 ;
        RECT 465.200 33.600 466.000 33.700 ;
        RECT 529.200 33.600 530.000 33.700 ;
        RECT 250.800 32.300 251.600 32.400 ;
        RECT 247.700 31.700 251.600 32.300 ;
        RECT 239.600 31.600 240.400 31.700 ;
        RECT 246.000 31.600 246.800 31.700 ;
        RECT 250.800 31.600 251.600 31.700 ;
        RECT 252.400 32.300 253.200 32.400 ;
        RECT 257.200 32.300 258.000 32.400 ;
        RECT 252.400 31.700 258.000 32.300 ;
        RECT 252.400 31.600 253.200 31.700 ;
        RECT 257.200 31.600 258.000 31.700 ;
        RECT 258.800 32.300 259.600 32.400 ;
        RECT 284.400 32.300 285.200 32.400 ;
        RECT 258.800 31.700 285.200 32.300 ;
        RECT 258.800 31.600 259.600 31.700 ;
        RECT 284.400 31.600 285.200 31.700 ;
        RECT 286.000 32.300 286.800 32.400 ;
        RECT 290.800 32.300 291.600 32.400 ;
        RECT 286.000 31.700 291.600 32.300 ;
        RECT 286.000 31.600 286.800 31.700 ;
        RECT 290.800 31.600 291.600 31.700 ;
        RECT 302.000 32.300 302.800 32.400 ;
        RECT 322.800 32.300 323.600 32.400 ;
        RECT 334.000 32.300 334.800 32.400 ;
        RECT 302.000 31.700 334.800 32.300 ;
        RECT 302.000 31.600 302.800 31.700 ;
        RECT 322.800 31.600 323.600 31.700 ;
        RECT 334.000 31.600 334.800 31.700 ;
        RECT 353.200 32.300 354.000 32.400 ;
        RECT 359.600 32.300 360.400 32.400 ;
        RECT 353.200 31.700 360.400 32.300 ;
        RECT 353.200 31.600 354.000 31.700 ;
        RECT 359.600 31.600 360.400 31.700 ;
        RECT 422.000 32.300 422.800 32.400 ;
        RECT 447.600 32.300 448.400 32.400 ;
        RECT 422.000 31.700 448.400 32.300 ;
        RECT 422.000 31.600 422.800 31.700 ;
        RECT 447.600 31.600 448.400 31.700 ;
        RECT 449.200 32.300 450.000 32.400 ;
        RECT 502.000 32.300 502.800 32.400 ;
        RECT 449.200 31.700 502.800 32.300 ;
        RECT 449.200 31.600 450.000 31.700 ;
        RECT 502.000 31.600 502.800 31.700 ;
        RECT 508.400 32.300 509.200 32.400 ;
        RECT 540.400 32.300 541.200 32.400 ;
        RECT 508.400 31.700 541.200 32.300 ;
        RECT 508.400 31.600 509.200 31.700 ;
        RECT 540.400 31.600 541.200 31.700 ;
        RECT 554.800 32.300 555.600 32.400 ;
        RECT 559.600 32.300 560.400 32.400 ;
        RECT 554.800 31.700 560.400 32.300 ;
        RECT 554.800 31.600 555.600 31.700 ;
        RECT 559.600 31.600 560.400 31.700 ;
        RECT 14.000 30.300 14.800 30.400 ;
        RECT 17.200 30.300 18.000 30.400 ;
        RECT 14.000 29.700 18.000 30.300 ;
        RECT 14.000 29.600 14.800 29.700 ;
        RECT 17.200 29.600 18.000 29.700 ;
        RECT 18.800 30.300 19.600 30.400 ;
        RECT 23.600 30.300 24.400 30.400 ;
        RECT 28.400 30.300 29.200 30.400 ;
        RECT 18.800 29.700 29.200 30.300 ;
        RECT 18.800 29.600 19.600 29.700 ;
        RECT 23.600 29.600 24.400 29.700 ;
        RECT 28.400 29.600 29.200 29.700 ;
        RECT 31.600 30.300 32.400 30.400 ;
        RECT 44.400 30.300 45.200 30.400 ;
        RECT 31.600 29.700 45.200 30.300 ;
        RECT 31.600 29.600 32.400 29.700 ;
        RECT 44.400 29.600 45.200 29.700 ;
        RECT 49.200 30.300 50.000 30.400 ;
        RECT 81.200 30.300 82.000 30.400 ;
        RECT 49.200 29.700 82.000 30.300 ;
        RECT 49.200 29.600 50.000 29.700 ;
        RECT 81.200 29.600 82.000 29.700 ;
        RECT 100.400 30.300 101.200 30.400 ;
        RECT 111.600 30.300 112.400 30.400 ;
        RECT 100.400 29.700 112.400 30.300 ;
        RECT 100.400 29.600 101.200 29.700 ;
        RECT 111.600 29.600 112.400 29.700 ;
        RECT 132.400 30.300 133.200 30.400 ;
        RECT 135.600 30.300 136.400 30.400 ;
        RECT 167.600 30.300 168.400 30.400 ;
        RECT 132.400 29.700 136.400 30.300 ;
        RECT 132.400 29.600 133.200 29.700 ;
        RECT 135.600 29.600 136.400 29.700 ;
        RECT 161.300 29.700 168.400 30.300 ;
        RECT 161.300 28.400 161.900 29.700 ;
        RECT 167.600 29.600 168.400 29.700 ;
        RECT 172.400 30.300 173.200 30.400 ;
        RECT 183.600 30.300 184.400 30.400 ;
        RECT 172.400 29.700 184.400 30.300 ;
        RECT 172.400 29.600 173.200 29.700 ;
        RECT 183.600 29.600 184.400 29.700 ;
        RECT 196.400 30.300 197.200 30.400 ;
        RECT 198.000 30.300 198.800 30.400 ;
        RECT 210.800 30.300 211.600 30.400 ;
        RECT 218.800 30.300 219.600 30.400 ;
        RECT 196.400 29.700 219.600 30.300 ;
        RECT 196.400 29.600 197.200 29.700 ;
        RECT 198.000 29.600 198.800 29.700 ;
        RECT 210.800 29.600 211.600 29.700 ;
        RECT 218.800 29.600 219.600 29.700 ;
        RECT 223.600 30.300 224.400 30.400 ;
        RECT 249.200 30.300 250.000 30.400 ;
        RECT 262.000 30.300 262.800 30.400 ;
        RECT 273.200 30.300 274.000 30.400 ;
        RECT 223.600 29.700 274.000 30.300 ;
        RECT 223.600 29.600 224.400 29.700 ;
        RECT 249.200 29.600 250.000 29.700 ;
        RECT 262.000 29.600 262.800 29.700 ;
        RECT 273.200 29.600 274.000 29.700 ;
        RECT 281.200 30.300 282.000 30.400 ;
        RECT 295.600 30.300 296.400 30.400 ;
        RECT 281.200 29.700 296.400 30.300 ;
        RECT 281.200 29.600 282.000 29.700 ;
        RECT 295.600 29.600 296.400 29.700 ;
        RECT 311.600 30.300 312.400 30.400 ;
        RECT 327.600 30.300 328.400 30.400 ;
        RECT 311.600 29.700 328.400 30.300 ;
        RECT 311.600 29.600 312.400 29.700 ;
        RECT 327.600 29.600 328.400 29.700 ;
        RECT 329.200 30.300 330.000 30.400 ;
        RECT 335.600 30.300 336.400 30.400 ;
        RECT 329.200 29.700 336.400 30.300 ;
        RECT 329.200 29.600 330.000 29.700 ;
        RECT 335.600 29.600 336.400 29.700 ;
        RECT 367.600 30.300 368.400 30.400 ;
        RECT 380.400 30.300 381.200 30.400 ;
        RECT 367.600 29.700 381.200 30.300 ;
        RECT 367.600 29.600 368.400 29.700 ;
        RECT 380.400 29.600 381.200 29.700 ;
        RECT 412.400 30.300 413.200 30.400 ;
        RECT 422.000 30.300 422.800 30.400 ;
        RECT 425.200 30.300 426.000 30.400 ;
        RECT 412.400 29.700 426.000 30.300 ;
        RECT 412.400 29.600 413.200 29.700 ;
        RECT 422.000 29.600 422.800 29.700 ;
        RECT 425.200 29.600 426.000 29.700 ;
        RECT 426.800 30.300 427.600 30.400 ;
        RECT 468.400 30.300 469.200 30.400 ;
        RECT 426.800 29.700 469.200 30.300 ;
        RECT 426.800 29.600 427.600 29.700 ;
        RECT 468.400 29.600 469.200 29.700 ;
        RECT 470.000 30.300 470.800 30.400 ;
        RECT 473.200 30.300 474.000 30.400 ;
        RECT 470.000 29.700 474.000 30.300 ;
        RECT 470.000 29.600 470.800 29.700 ;
        RECT 473.200 29.600 474.000 29.700 ;
        RECT 484.400 30.300 485.200 30.400 ;
        RECT 511.600 30.300 512.400 30.400 ;
        RECT 514.800 30.300 515.600 30.400 ;
        RECT 543.600 30.300 544.400 30.400 ;
        RECT 484.400 29.700 544.400 30.300 ;
        RECT 484.400 29.600 485.200 29.700 ;
        RECT 511.600 29.600 512.400 29.700 ;
        RECT 514.800 29.600 515.600 29.700 ;
        RECT 543.600 29.600 544.400 29.700 ;
        RECT 550.000 30.300 550.800 30.400 ;
        RECT 562.800 30.300 563.600 30.400 ;
        RECT 550.000 29.700 563.600 30.300 ;
        RECT 550.000 29.600 550.800 29.700 ;
        RECT 562.800 29.600 563.600 29.700 ;
        RECT 569.200 30.300 570.000 30.400 ;
        RECT 578.800 30.300 579.600 30.400 ;
        RECT 569.200 29.700 579.600 30.300 ;
        RECT 569.200 29.600 570.000 29.700 ;
        RECT 578.800 29.600 579.600 29.700 ;
        RECT 9.200 28.300 10.000 28.400 ;
        RECT 25.200 28.300 26.000 28.400 ;
        RECT 9.200 27.700 26.000 28.300 ;
        RECT 9.200 27.600 10.000 27.700 ;
        RECT 25.200 27.600 26.000 27.700 ;
        RECT 44.400 28.300 45.200 28.400 ;
        RECT 58.800 28.300 59.600 28.400 ;
        RECT 44.400 27.700 59.600 28.300 ;
        RECT 44.400 27.600 45.200 27.700 ;
        RECT 58.800 27.600 59.600 27.700 ;
        RECT 89.200 28.300 90.000 28.400 ;
        RECT 100.400 28.300 101.200 28.400 ;
        RECT 89.200 27.700 101.200 28.300 ;
        RECT 89.200 27.600 90.000 27.700 ;
        RECT 100.400 27.600 101.200 27.700 ;
        RECT 142.000 28.300 142.800 28.400 ;
        RECT 161.200 28.300 162.000 28.400 ;
        RECT 142.000 27.700 162.000 28.300 ;
        RECT 142.000 27.600 142.800 27.700 ;
        RECT 161.200 27.600 162.000 27.700 ;
        RECT 162.800 28.300 163.600 28.400 ;
        RECT 198.000 28.300 198.800 28.400 ;
        RECT 206.000 28.300 206.800 28.400 ;
        RECT 162.800 27.700 206.800 28.300 ;
        RECT 162.800 27.600 163.600 27.700 ;
        RECT 198.000 27.600 198.800 27.700 ;
        RECT 206.000 27.600 206.800 27.700 ;
        RECT 214.000 28.300 214.800 28.400 ;
        RECT 220.400 28.300 221.200 28.400 ;
        RECT 214.000 27.700 221.200 28.300 ;
        RECT 214.000 27.600 214.800 27.700 ;
        RECT 220.400 27.600 221.200 27.700 ;
        RECT 226.800 28.300 227.600 28.400 ;
        RECT 255.600 28.300 256.400 28.400 ;
        RECT 266.800 28.300 267.600 28.400 ;
        RECT 226.800 27.700 267.600 28.300 ;
        RECT 226.800 27.600 227.600 27.700 ;
        RECT 255.600 27.600 256.400 27.700 ;
        RECT 266.800 27.600 267.600 27.700 ;
        RECT 284.400 28.300 285.200 28.400 ;
        RECT 286.000 28.300 286.800 28.400 ;
        RECT 284.400 27.700 286.800 28.300 ;
        RECT 284.400 27.600 285.200 27.700 ;
        RECT 286.000 27.600 286.800 27.700 ;
        RECT 297.200 28.300 298.000 28.400 ;
        RECT 306.800 28.300 307.600 28.400 ;
        RECT 308.400 28.300 309.200 28.400 ;
        RECT 297.200 27.700 309.200 28.300 ;
        RECT 297.200 27.600 298.000 27.700 ;
        RECT 306.800 27.600 307.600 27.700 ;
        RECT 308.400 27.600 309.200 27.700 ;
        RECT 314.800 28.300 315.600 28.400 ;
        RECT 319.600 28.300 320.400 28.400 ;
        RECT 324.400 28.300 325.200 28.400 ;
        RECT 314.800 27.700 325.200 28.300 ;
        RECT 314.800 27.600 315.600 27.700 ;
        RECT 319.600 27.600 320.400 27.700 ;
        RECT 324.400 27.600 325.200 27.700 ;
        RECT 343.600 28.300 344.400 28.400 ;
        RECT 346.800 28.300 347.600 28.400 ;
        RECT 343.600 27.700 347.600 28.300 ;
        RECT 343.600 27.600 344.400 27.700 ;
        RECT 346.800 27.600 347.600 27.700 ;
        RECT 361.200 28.300 362.000 28.400 ;
        RECT 374.000 28.300 374.800 28.400 ;
        RECT 361.200 27.700 374.800 28.300 ;
        RECT 361.200 27.600 362.000 27.700 ;
        RECT 374.000 27.600 374.800 27.700 ;
        RECT 414.000 28.300 414.800 28.400 ;
        RECT 428.400 28.300 429.200 28.400 ;
        RECT 431.600 28.300 432.400 28.400 ;
        RECT 414.000 27.700 432.400 28.300 ;
        RECT 414.000 27.600 414.800 27.700 ;
        RECT 428.400 27.600 429.200 27.700 ;
        RECT 431.600 27.600 432.400 27.700 ;
        RECT 433.200 28.300 434.000 28.400 ;
        RECT 438.000 28.300 438.800 28.400 ;
        RECT 433.200 27.700 438.800 28.300 ;
        RECT 433.200 27.600 434.000 27.700 ;
        RECT 438.000 27.600 438.800 27.700 ;
        RECT 439.600 28.300 440.400 28.400 ;
        RECT 462.000 28.300 462.800 28.400 ;
        RECT 439.600 27.700 462.800 28.300 ;
        RECT 439.600 27.600 440.400 27.700 ;
        RECT 462.000 27.600 462.800 27.700 ;
        RECT 463.600 28.300 464.400 28.400 ;
        RECT 510.000 28.300 510.800 28.400 ;
        RECT 550.000 28.300 550.800 28.400 ;
        RECT 463.600 27.700 550.800 28.300 ;
        RECT 463.600 27.600 464.400 27.700 ;
        RECT 510.000 27.600 510.800 27.700 ;
        RECT 550.000 27.600 550.800 27.700 ;
        RECT 554.800 28.300 555.600 28.400 ;
        RECT 564.400 28.300 565.200 28.400 ;
        RECT 554.800 27.700 565.200 28.300 ;
        RECT 554.800 27.600 555.600 27.700 ;
        RECT 564.400 27.600 565.200 27.700 ;
        RECT 578.800 28.300 579.600 28.400 ;
        RECT 582.000 28.300 582.800 28.400 ;
        RECT 578.800 27.700 582.800 28.300 ;
        RECT 578.800 27.600 579.600 27.700 ;
        RECT 582.000 27.600 582.800 27.700 ;
        RECT 1.200 26.300 2.000 26.400 ;
        RECT 17.200 26.300 18.000 26.400 ;
        RECT 28.400 26.300 29.200 26.400 ;
        RECT 1.200 25.700 29.200 26.300 ;
        RECT 1.200 25.600 2.000 25.700 ;
        RECT 17.200 25.600 18.000 25.700 ;
        RECT 28.400 25.600 29.200 25.700 ;
        RECT 41.200 26.300 42.000 26.400 ;
        RECT 46.000 26.300 46.800 26.400 ;
        RECT 41.200 25.700 46.800 26.300 ;
        RECT 41.200 25.600 42.000 25.700 ;
        RECT 46.000 25.600 46.800 25.700 ;
        RECT 57.200 26.300 58.000 26.400 ;
        RECT 153.200 26.300 154.000 26.400 ;
        RECT 57.200 25.700 154.000 26.300 ;
        RECT 57.200 25.600 58.000 25.700 ;
        RECT 153.200 25.600 154.000 25.700 ;
        RECT 182.000 26.300 182.800 26.400 ;
        RECT 196.400 26.300 197.200 26.400 ;
        RECT 182.000 25.700 197.200 26.300 ;
        RECT 182.000 25.600 182.800 25.700 ;
        RECT 196.400 25.600 197.200 25.700 ;
        RECT 209.200 26.300 210.000 26.400 ;
        RECT 217.200 26.300 218.000 26.400 ;
        RECT 209.200 25.700 218.000 26.300 ;
        RECT 209.200 25.600 210.000 25.700 ;
        RECT 217.200 25.600 218.000 25.700 ;
        RECT 218.800 26.300 219.600 26.400 ;
        RECT 278.000 26.300 278.800 26.400 ;
        RECT 218.800 25.700 278.800 26.300 ;
        RECT 218.800 25.600 219.600 25.700 ;
        RECT 278.000 25.600 278.800 25.700 ;
        RECT 316.400 26.300 317.200 26.400 ;
        RECT 346.900 26.300 347.500 27.600 ;
        RECT 361.200 26.300 362.000 26.400 ;
        RECT 316.400 25.700 362.000 26.300 ;
        RECT 316.400 25.600 317.200 25.700 ;
        RECT 361.200 25.600 362.000 25.700 ;
        RECT 407.600 26.300 408.400 26.400 ;
        RECT 412.400 26.300 413.200 26.400 ;
        RECT 450.800 26.300 451.600 26.400 ;
        RECT 476.400 26.300 477.200 26.400 ;
        RECT 505.200 26.300 506.000 26.400 ;
        RECT 407.600 25.700 506.000 26.300 ;
        RECT 407.600 25.600 408.400 25.700 ;
        RECT 412.400 25.600 413.200 25.700 ;
        RECT 450.800 25.600 451.600 25.700 ;
        RECT 476.400 25.600 477.200 25.700 ;
        RECT 505.200 25.600 506.000 25.700 ;
        RECT 506.800 26.300 507.600 26.400 ;
        RECT 508.400 26.300 509.200 26.400 ;
        RECT 518.000 26.300 518.800 26.400 ;
        RECT 506.800 25.700 518.800 26.300 ;
        RECT 506.800 25.600 507.600 25.700 ;
        RECT 508.400 25.600 509.200 25.700 ;
        RECT 518.000 25.600 518.800 25.700 ;
        RECT 561.200 26.300 562.000 26.400 ;
        RECT 575.600 26.300 576.400 26.400 ;
        RECT 561.200 25.700 576.400 26.300 ;
        RECT 561.200 25.600 562.000 25.700 ;
        RECT 575.600 25.600 576.400 25.700 ;
        RECT 65.200 24.300 66.000 24.400 ;
        RECT 102.000 24.300 102.800 24.400 ;
        RECT 65.200 23.700 102.800 24.300 ;
        RECT 65.200 23.600 66.000 23.700 ;
        RECT 102.000 23.600 102.800 23.700 ;
        RECT 122.800 24.300 123.600 24.400 ;
        RECT 129.200 24.300 130.000 24.400 ;
        RECT 122.800 23.700 130.000 24.300 ;
        RECT 122.800 23.600 123.600 23.700 ;
        RECT 129.200 23.600 130.000 23.700 ;
        RECT 134.000 24.300 134.800 24.400 ;
        RECT 230.000 24.300 230.800 24.400 ;
        RECT 231.600 24.300 232.400 24.400 ;
        RECT 265.200 24.300 266.000 24.400 ;
        RECT 276.400 24.300 277.200 24.400 ;
        RECT 300.400 24.300 301.200 24.400 ;
        RECT 134.000 23.700 277.200 24.300 ;
        RECT 134.000 23.600 134.800 23.700 ;
        RECT 230.000 23.600 230.800 23.700 ;
        RECT 231.600 23.600 232.400 23.700 ;
        RECT 265.200 23.600 266.000 23.700 ;
        RECT 276.400 23.600 277.200 23.700 ;
        RECT 287.700 23.700 301.200 24.300 ;
        RECT 124.400 22.300 125.200 22.400 ;
        RECT 142.000 22.300 142.800 22.400 ;
        RECT 124.400 21.700 142.800 22.300 ;
        RECT 124.400 21.600 125.200 21.700 ;
        RECT 142.000 21.600 142.800 21.700 ;
        RECT 159.600 22.300 160.400 22.400 ;
        RECT 172.400 22.300 173.200 22.400 ;
        RECT 159.600 21.700 173.200 22.300 ;
        RECT 159.600 21.600 160.400 21.700 ;
        RECT 172.400 21.600 173.200 21.700 ;
        RECT 178.800 22.300 179.600 22.400 ;
        RECT 185.200 22.300 186.000 22.400 ;
        RECT 178.800 21.700 186.000 22.300 ;
        RECT 178.800 21.600 179.600 21.700 ;
        RECT 185.200 21.600 186.000 21.700 ;
        RECT 193.200 22.300 194.000 22.400 ;
        RECT 217.200 22.300 218.000 22.400 ;
        RECT 233.200 22.300 234.000 22.400 ;
        RECT 239.600 22.300 240.400 22.400 ;
        RECT 193.200 21.700 240.400 22.300 ;
        RECT 193.200 21.600 194.000 21.700 ;
        RECT 217.200 21.600 218.000 21.700 ;
        RECT 233.200 21.600 234.000 21.700 ;
        RECT 239.600 21.600 240.400 21.700 ;
        RECT 244.400 22.300 245.200 22.400 ;
        RECT 254.000 22.300 254.800 22.400 ;
        RECT 244.400 21.700 254.800 22.300 ;
        RECT 244.400 21.600 245.200 21.700 ;
        RECT 254.000 21.600 254.800 21.700 ;
        RECT 265.200 22.300 266.000 22.400 ;
        RECT 287.700 22.300 288.300 23.700 ;
        RECT 300.400 23.600 301.200 23.700 ;
        RECT 305.200 24.300 306.000 24.400 ;
        RECT 337.200 24.300 338.000 24.400 ;
        RECT 342.000 24.300 342.800 24.400 ;
        RECT 305.200 23.700 342.800 24.300 ;
        RECT 305.200 23.600 306.000 23.700 ;
        RECT 337.200 23.600 338.000 23.700 ;
        RECT 342.000 23.600 342.800 23.700 ;
        RECT 393.200 24.300 394.000 24.400 ;
        RECT 466.800 24.300 467.600 24.400 ;
        RECT 478.000 24.300 478.800 24.400 ;
        RECT 393.200 23.700 464.300 24.300 ;
        RECT 393.200 23.600 394.000 23.700 ;
        RECT 463.700 22.400 464.300 23.700 ;
        RECT 466.800 23.700 478.800 24.300 ;
        RECT 466.800 23.600 467.600 23.700 ;
        RECT 478.000 23.600 478.800 23.700 ;
        RECT 481.200 24.300 482.000 24.400 ;
        RECT 490.800 24.300 491.600 24.400 ;
        RECT 481.200 23.700 491.600 24.300 ;
        RECT 481.200 23.600 482.000 23.700 ;
        RECT 490.800 23.600 491.600 23.700 ;
        RECT 497.200 24.300 498.000 24.400 ;
        RECT 514.800 24.300 515.600 24.400 ;
        RECT 526.000 24.300 526.800 24.400 ;
        RECT 497.200 23.700 526.800 24.300 ;
        RECT 497.200 23.600 498.000 23.700 ;
        RECT 514.800 23.600 515.600 23.700 ;
        RECT 526.000 23.600 526.800 23.700 ;
        RECT 551.600 24.300 552.400 24.400 ;
        RECT 577.200 24.300 578.000 24.400 ;
        RECT 551.600 23.700 578.000 24.300 ;
        RECT 551.600 23.600 552.400 23.700 ;
        RECT 577.200 23.600 578.000 23.700 ;
        RECT 265.200 21.700 288.300 22.300 ;
        RECT 356.400 22.300 357.200 22.400 ;
        RECT 410.800 22.300 411.600 22.400 ;
        RECT 418.800 22.300 419.600 22.400 ;
        RECT 452.400 22.300 453.200 22.400 ;
        RECT 457.200 22.300 458.000 22.400 ;
        RECT 356.400 21.700 441.900 22.300 ;
        RECT 265.200 21.600 266.000 21.700 ;
        RECT 356.400 21.600 357.200 21.700 ;
        RECT 410.800 21.600 411.600 21.700 ;
        RECT 418.800 21.600 419.600 21.700 ;
        RECT 441.300 20.400 441.900 21.700 ;
        RECT 452.400 21.700 458.000 22.300 ;
        RECT 452.400 21.600 453.200 21.700 ;
        RECT 457.200 21.600 458.000 21.700 ;
        RECT 463.600 22.300 464.400 22.400 ;
        RECT 481.200 22.300 482.000 22.400 ;
        RECT 505.200 22.300 506.000 22.400 ;
        RECT 508.400 22.300 509.200 22.400 ;
        RECT 463.600 21.700 501.100 22.300 ;
        RECT 463.600 21.600 464.400 21.700 ;
        RECT 481.200 21.600 482.000 21.700 ;
        RECT 500.500 20.400 501.100 21.700 ;
        RECT 505.200 21.700 509.200 22.300 ;
        RECT 505.200 21.600 506.000 21.700 ;
        RECT 508.400 21.600 509.200 21.700 ;
        RECT 518.000 22.300 518.800 22.400 ;
        RECT 519.600 22.300 520.400 22.400 ;
        RECT 518.000 21.700 520.400 22.300 ;
        RECT 518.000 21.600 518.800 21.700 ;
        RECT 519.600 21.600 520.400 21.700 ;
        RECT 527.600 22.300 528.400 22.400 ;
        RECT 542.000 22.300 542.800 22.400 ;
        RECT 548.400 22.300 549.200 22.400 ;
        RECT 566.000 22.300 566.800 22.400 ;
        RECT 527.600 21.700 566.800 22.300 ;
        RECT 527.600 21.600 528.400 21.700 ;
        RECT 542.000 21.600 542.800 21.700 ;
        RECT 548.400 21.600 549.200 21.700 ;
        RECT 566.000 21.600 566.800 21.700 ;
        RECT 575.600 22.300 576.400 22.400 ;
        RECT 577.200 22.300 578.000 22.400 ;
        RECT 575.600 21.700 578.000 22.300 ;
        RECT 575.600 21.600 576.400 21.700 ;
        RECT 577.200 21.600 578.000 21.700 ;
        RECT 1.200 20.300 2.000 20.400 ;
        RECT 4.400 20.300 5.200 20.400 ;
        RECT 1.200 19.700 5.200 20.300 ;
        RECT 1.200 19.600 2.000 19.700 ;
        RECT 4.400 19.600 5.200 19.700 ;
        RECT 34.800 20.300 35.600 20.400 ;
        RECT 63.600 20.300 64.400 20.400 ;
        RECT 34.800 19.700 64.400 20.300 ;
        RECT 34.800 19.600 35.600 19.700 ;
        RECT 63.600 19.600 64.400 19.700 ;
        RECT 76.400 20.300 77.200 20.400 ;
        RECT 177.200 20.300 178.000 20.400 ;
        RECT 76.400 19.700 178.000 20.300 ;
        RECT 76.400 19.600 77.200 19.700 ;
        RECT 177.200 19.600 178.000 19.700 ;
        RECT 188.400 20.300 189.200 20.400 ;
        RECT 202.800 20.300 203.600 20.400 ;
        RECT 249.200 20.300 250.000 20.400 ;
        RECT 265.200 20.300 266.000 20.400 ;
        RECT 188.400 19.700 266.000 20.300 ;
        RECT 188.400 19.600 189.200 19.700 ;
        RECT 202.800 19.600 203.600 19.700 ;
        RECT 249.200 19.600 250.000 19.700 ;
        RECT 265.200 19.600 266.000 19.700 ;
        RECT 302.000 20.300 302.800 20.400 ;
        RECT 310.000 20.300 310.800 20.400 ;
        RECT 302.000 19.700 310.800 20.300 ;
        RECT 302.000 19.600 302.800 19.700 ;
        RECT 310.000 19.600 310.800 19.700 ;
        RECT 324.400 20.300 325.200 20.400 ;
        RECT 345.200 20.300 346.000 20.400 ;
        RECT 324.400 19.700 346.000 20.300 ;
        RECT 324.400 19.600 325.200 19.700 ;
        RECT 345.200 19.600 346.000 19.700 ;
        RECT 409.200 20.300 410.000 20.400 ;
        RECT 426.800 20.300 427.600 20.400 ;
        RECT 409.200 19.700 427.600 20.300 ;
        RECT 409.200 19.600 410.000 19.700 ;
        RECT 426.800 19.600 427.600 19.700 ;
        RECT 428.400 20.300 429.200 20.400 ;
        RECT 433.200 20.300 434.000 20.400 ;
        RECT 428.400 19.700 434.000 20.300 ;
        RECT 428.400 19.600 429.200 19.700 ;
        RECT 433.200 19.600 434.000 19.700 ;
        RECT 434.800 19.600 435.600 20.400 ;
        RECT 438.000 19.600 438.800 20.400 ;
        RECT 441.200 20.300 442.000 20.400 ;
        RECT 444.400 20.300 445.200 20.400 ;
        RECT 441.200 19.700 445.200 20.300 ;
        RECT 441.200 19.600 442.000 19.700 ;
        RECT 444.400 19.600 445.200 19.700 ;
        RECT 455.600 20.300 456.400 20.400 ;
        RECT 474.800 20.300 475.600 20.400 ;
        RECT 482.800 20.300 483.600 20.400 ;
        RECT 455.600 19.700 483.600 20.300 ;
        RECT 455.600 19.600 456.400 19.700 ;
        RECT 474.800 19.600 475.600 19.700 ;
        RECT 482.800 19.600 483.600 19.700 ;
        RECT 500.400 20.300 501.200 20.400 ;
        RECT 506.800 20.300 507.600 20.400 ;
        RECT 500.400 19.700 507.600 20.300 ;
        RECT 500.400 19.600 501.200 19.700 ;
        RECT 506.800 19.600 507.600 19.700 ;
        RECT 513.200 20.300 514.000 20.400 ;
        RECT 538.800 20.300 539.600 20.400 ;
        RECT 513.200 19.700 539.600 20.300 ;
        RECT 513.200 19.600 514.000 19.700 ;
        RECT 538.800 19.600 539.600 19.700 ;
        RECT 559.600 20.300 560.400 20.400 ;
        RECT 569.200 20.300 570.000 20.400 ;
        RECT 559.600 19.700 570.000 20.300 ;
        RECT 559.600 19.600 560.400 19.700 ;
        RECT 569.200 19.600 570.000 19.700 ;
        RECT 20.400 18.300 21.200 18.400 ;
        RECT 38.000 18.300 38.800 18.400 ;
        RECT 20.400 17.700 38.800 18.300 ;
        RECT 20.400 17.600 21.200 17.700 ;
        RECT 38.000 17.600 38.800 17.700 ;
        RECT 95.600 18.300 96.400 18.400 ;
        RECT 102.000 18.300 102.800 18.400 ;
        RECT 95.600 17.700 102.800 18.300 ;
        RECT 95.600 17.600 96.400 17.700 ;
        RECT 102.000 17.600 102.800 17.700 ;
        RECT 114.800 18.300 115.600 18.400 ;
        RECT 140.400 18.300 141.200 18.400 ;
        RECT 114.800 17.700 141.200 18.300 ;
        RECT 114.800 17.600 115.600 17.700 ;
        RECT 140.400 17.600 141.200 17.700 ;
        RECT 148.400 18.300 149.200 18.400 ;
        RECT 174.000 18.300 174.800 18.400 ;
        RECT 186.800 18.300 187.600 18.400 ;
        RECT 148.400 17.700 187.600 18.300 ;
        RECT 148.400 17.600 149.200 17.700 ;
        RECT 174.000 17.600 174.800 17.700 ;
        RECT 186.800 17.600 187.600 17.700 ;
        RECT 191.600 18.300 192.400 18.400 ;
        RECT 198.000 18.300 198.800 18.400 ;
        RECT 191.600 17.700 198.800 18.300 ;
        RECT 191.600 17.600 192.400 17.700 ;
        RECT 198.000 17.600 198.800 17.700 ;
        RECT 199.600 18.300 200.400 18.400 ;
        RECT 210.800 18.300 211.600 18.400 ;
        RECT 199.600 17.700 211.600 18.300 ;
        RECT 199.600 17.600 200.400 17.700 ;
        RECT 210.800 17.600 211.600 17.700 ;
        RECT 215.600 18.300 216.400 18.400 ;
        RECT 220.400 18.300 221.200 18.400 ;
        RECT 215.600 17.700 221.200 18.300 ;
        RECT 215.600 17.600 216.400 17.700 ;
        RECT 220.400 17.600 221.200 17.700 ;
        RECT 225.200 18.300 226.000 18.400 ;
        RECT 244.400 18.300 245.200 18.400 ;
        RECT 225.200 17.700 245.200 18.300 ;
        RECT 225.200 17.600 226.000 17.700 ;
        RECT 244.400 17.600 245.200 17.700 ;
        RECT 246.000 18.300 246.800 18.400 ;
        RECT 252.400 18.300 253.200 18.400 ;
        RECT 246.000 17.700 253.200 18.300 ;
        RECT 246.000 17.600 246.800 17.700 ;
        RECT 252.400 17.600 253.200 17.700 ;
        RECT 254.000 18.300 254.800 18.400 ;
        RECT 265.200 18.300 266.000 18.400 ;
        RECT 287.600 18.300 288.400 18.400 ;
        RECT 254.000 17.700 266.000 18.300 ;
        RECT 254.000 17.600 254.800 17.700 ;
        RECT 265.200 17.600 266.000 17.700 ;
        RECT 266.900 17.700 288.400 18.300 ;
        RECT 151.600 16.300 152.400 16.400 ;
        RECT 154.800 16.300 155.600 16.400 ;
        RECT 151.600 15.700 155.600 16.300 ;
        RECT 151.600 15.600 152.400 15.700 ;
        RECT 154.800 15.600 155.600 15.700 ;
        RECT 159.600 16.300 160.400 16.400 ;
        RECT 164.400 16.300 165.200 16.400 ;
        RECT 159.600 15.700 165.200 16.300 ;
        RECT 159.600 15.600 160.400 15.700 ;
        RECT 164.400 15.600 165.200 15.700 ;
        RECT 170.800 16.300 171.600 16.400 ;
        RECT 194.800 16.300 195.600 16.400 ;
        RECT 263.600 16.300 264.400 16.400 ;
        RECT 266.900 16.300 267.500 17.700 ;
        RECT 287.600 17.600 288.400 17.700 ;
        RECT 289.200 18.300 290.000 18.400 ;
        RECT 310.000 18.300 310.800 18.400 ;
        RECT 332.400 18.300 333.200 18.400 ;
        RECT 337.200 18.300 338.000 18.400 ;
        RECT 289.200 17.700 338.000 18.300 ;
        RECT 289.200 17.600 290.000 17.700 ;
        RECT 310.000 17.600 310.800 17.700 ;
        RECT 332.400 17.600 333.200 17.700 ;
        RECT 337.200 17.600 338.000 17.700 ;
        RECT 423.600 18.300 424.400 18.400 ;
        RECT 522.800 18.300 523.600 18.400 ;
        RECT 548.400 18.300 549.200 18.400 ;
        RECT 423.600 17.700 549.200 18.300 ;
        RECT 423.600 17.600 424.400 17.700 ;
        RECT 522.800 17.600 523.600 17.700 ;
        RECT 548.400 17.600 549.200 17.700 ;
        RECT 564.400 18.300 565.200 18.400 ;
        RECT 572.400 18.300 573.200 18.400 ;
        RECT 582.000 18.300 582.800 18.400 ;
        RECT 564.400 17.700 582.800 18.300 ;
        RECT 564.400 17.600 565.200 17.700 ;
        RECT 572.400 17.600 573.200 17.700 ;
        RECT 582.000 17.600 582.800 17.700 ;
        RECT 170.800 15.700 267.500 16.300 ;
        RECT 268.400 16.300 269.200 16.400 ;
        RECT 274.800 16.300 275.600 16.400 ;
        RECT 268.400 15.700 275.600 16.300 ;
        RECT 170.800 15.600 171.600 15.700 ;
        RECT 194.800 15.600 195.600 15.700 ;
        RECT 263.600 15.600 264.400 15.700 ;
        RECT 268.400 15.600 269.200 15.700 ;
        RECT 274.800 15.600 275.600 15.700 ;
        RECT 276.400 16.300 277.200 16.400 ;
        RECT 297.200 16.300 298.000 16.400 ;
        RECT 276.400 15.700 298.000 16.300 ;
        RECT 276.400 15.600 277.200 15.700 ;
        RECT 297.200 15.600 298.000 15.700 ;
        RECT 300.400 16.300 301.200 16.400 ;
        RECT 306.800 16.300 307.600 16.400 ;
        RECT 300.400 15.700 307.600 16.300 ;
        RECT 300.400 15.600 301.200 15.700 ;
        RECT 306.800 15.600 307.600 15.700 ;
        RECT 308.400 16.300 309.200 16.400 ;
        RECT 316.400 16.300 317.200 16.400 ;
        RECT 308.400 15.700 317.200 16.300 ;
        RECT 308.400 15.600 309.200 15.700 ;
        RECT 316.400 15.600 317.200 15.700 ;
        RECT 322.800 16.300 323.600 16.400 ;
        RECT 327.600 16.300 328.400 16.400 ;
        RECT 322.800 15.700 328.400 16.300 ;
        RECT 322.800 15.600 323.600 15.700 ;
        RECT 327.600 15.600 328.400 15.700 ;
        RECT 375.600 16.300 376.400 16.400 ;
        RECT 402.800 16.300 403.600 16.400 ;
        RECT 414.000 16.300 414.800 16.400 ;
        RECT 375.600 15.700 414.800 16.300 ;
        RECT 375.600 15.600 376.400 15.700 ;
        RECT 402.800 15.600 403.600 15.700 ;
        RECT 414.000 15.600 414.800 15.700 ;
        RECT 415.600 16.300 416.400 16.400 ;
        RECT 433.200 16.300 434.000 16.400 ;
        RECT 457.200 16.300 458.000 16.400 ;
        RECT 415.600 15.700 458.000 16.300 ;
        RECT 415.600 15.600 416.400 15.700 ;
        RECT 433.200 15.600 434.000 15.700 ;
        RECT 457.200 15.600 458.000 15.700 ;
        RECT 458.800 16.300 459.600 16.400 ;
        RECT 466.800 16.300 467.600 16.400 ;
        RECT 458.800 15.700 467.600 16.300 ;
        RECT 458.800 15.600 459.600 15.700 ;
        RECT 466.800 15.600 467.600 15.700 ;
        RECT 468.400 16.300 469.200 16.400 ;
        RECT 492.400 16.300 493.200 16.400 ;
        RECT 468.400 15.700 493.200 16.300 ;
        RECT 468.400 15.600 469.200 15.700 ;
        RECT 492.400 15.600 493.200 15.700 ;
        RECT 506.800 16.300 507.600 16.400 ;
        RECT 510.000 16.300 510.800 16.400 ;
        RECT 506.800 15.700 510.800 16.300 ;
        RECT 506.800 15.600 507.600 15.700 ;
        RECT 510.000 15.600 510.800 15.700 ;
        RECT 511.600 16.300 512.400 16.400 ;
        RECT 535.600 16.300 536.400 16.400 ;
        RECT 511.600 15.700 536.400 16.300 ;
        RECT 511.600 15.600 512.400 15.700 ;
        RECT 535.600 15.600 536.400 15.700 ;
        RECT 546.800 16.300 547.600 16.400 ;
        RECT 570.800 16.300 571.600 16.400 ;
        RECT 546.800 15.700 571.600 16.300 ;
        RECT 546.800 15.600 547.600 15.700 ;
        RECT 570.800 15.600 571.600 15.700 ;
        RECT 2.800 14.300 3.600 14.400 ;
        RECT 17.200 14.300 18.000 14.400 ;
        RECT 2.800 13.700 18.000 14.300 ;
        RECT 2.800 13.600 3.600 13.700 ;
        RECT 17.200 13.600 18.000 13.700 ;
        RECT 150.000 14.300 150.800 14.400 ;
        RECT 161.200 14.300 162.000 14.400 ;
        RECT 150.000 13.700 162.000 14.300 ;
        RECT 150.000 13.600 150.800 13.700 ;
        RECT 161.200 13.600 162.000 13.700 ;
        RECT 182.000 14.300 182.800 14.400 ;
        RECT 212.400 14.300 213.200 14.400 ;
        RECT 182.000 13.700 213.200 14.300 ;
        RECT 182.000 13.600 182.800 13.700 ;
        RECT 212.400 13.600 213.200 13.700 ;
        RECT 223.600 13.600 224.400 14.400 ;
        RECT 231.600 14.300 232.400 14.400 ;
        RECT 244.400 14.300 245.200 14.400 ;
        RECT 231.600 13.700 245.200 14.300 ;
        RECT 231.600 13.600 232.400 13.700 ;
        RECT 244.400 13.600 245.200 13.700 ;
        RECT 246.000 13.600 246.800 14.400 ;
        RECT 247.600 14.300 248.400 14.400 ;
        RECT 249.200 14.300 250.000 14.400 ;
        RECT 247.600 13.700 250.000 14.300 ;
        RECT 247.600 13.600 248.400 13.700 ;
        RECT 249.200 13.600 250.000 13.700 ;
        RECT 254.000 14.300 254.800 14.400 ;
        RECT 260.400 14.300 261.200 14.400 ;
        RECT 326.000 14.300 326.800 14.400 ;
        RECT 254.000 13.700 326.800 14.300 ;
        RECT 254.000 13.600 254.800 13.700 ;
        RECT 260.400 13.600 261.200 13.700 ;
        RECT 326.000 13.600 326.800 13.700 ;
        RECT 350.000 14.300 350.800 14.400 ;
        RECT 369.200 14.300 370.000 14.400 ;
        RECT 385.200 14.300 386.000 14.400 ;
        RECT 350.000 13.700 386.000 14.300 ;
        RECT 350.000 13.600 350.800 13.700 ;
        RECT 369.200 13.600 370.000 13.700 ;
        RECT 385.200 13.600 386.000 13.700 ;
        RECT 401.200 14.300 402.000 14.400 ;
        RECT 412.400 14.300 413.200 14.400 ;
        RECT 401.200 13.700 413.200 14.300 ;
        RECT 414.100 14.300 414.700 15.600 ;
        RECT 417.200 14.300 418.000 14.400 ;
        RECT 414.100 13.700 418.000 14.300 ;
        RECT 401.200 13.600 402.000 13.700 ;
        RECT 412.400 13.600 413.200 13.700 ;
        RECT 417.200 13.600 418.000 13.700 ;
        RECT 422.000 14.300 422.800 14.400 ;
        RECT 430.000 14.300 430.800 14.400 ;
        RECT 422.000 13.700 430.800 14.300 ;
        RECT 422.000 13.600 422.800 13.700 ;
        RECT 430.000 13.600 430.800 13.700 ;
        RECT 446.000 14.300 446.800 14.400 ;
        RECT 452.400 14.300 453.200 14.400 ;
        RECT 495.600 14.300 496.400 14.400 ;
        RECT 502.000 14.300 502.800 14.400 ;
        RECT 516.400 14.300 517.200 14.400 ;
        RECT 527.600 14.300 528.400 14.400 ;
        RECT 446.000 13.700 453.200 14.300 ;
        RECT 446.000 13.600 446.800 13.700 ;
        RECT 452.400 13.600 453.200 13.700 ;
        RECT 479.700 13.700 502.800 14.300 ;
        RECT 12.400 12.300 13.200 12.400 ;
        RECT 26.800 12.300 27.600 12.400 ;
        RECT 12.400 11.700 27.600 12.300 ;
        RECT 12.400 11.600 13.200 11.700 ;
        RECT 26.800 11.600 27.600 11.700 ;
        RECT 50.800 12.300 51.600 12.400 ;
        RECT 60.400 12.300 61.200 12.400 ;
        RECT 50.800 11.700 61.200 12.300 ;
        RECT 50.800 11.600 51.600 11.700 ;
        RECT 60.400 11.600 61.200 11.700 ;
        RECT 63.600 11.600 64.400 12.400 ;
        RECT 70.000 12.300 70.800 12.400 ;
        RECT 89.200 12.300 90.000 12.400 ;
        RECT 98.800 12.300 99.600 12.400 ;
        RECT 70.000 11.700 99.600 12.300 ;
        RECT 70.000 11.600 70.800 11.700 ;
        RECT 89.200 11.600 90.000 11.700 ;
        RECT 98.800 11.600 99.600 11.700 ;
        RECT 178.800 12.300 179.600 12.400 ;
        RECT 199.600 12.300 200.400 12.400 ;
        RECT 206.000 12.300 206.800 12.400 ;
        RECT 178.800 11.700 206.800 12.300 ;
        RECT 212.500 12.300 213.100 13.600 ;
        RECT 479.700 12.400 480.300 13.700 ;
        RECT 495.600 13.600 496.400 13.700 ;
        RECT 502.000 13.600 502.800 13.700 ;
        RECT 503.700 13.700 515.500 14.300 ;
        RECT 281.200 12.300 282.000 12.400 ;
        RECT 212.500 11.700 282.000 12.300 ;
        RECT 178.800 11.600 179.600 11.700 ;
        RECT 199.600 11.600 200.400 11.700 ;
        RECT 206.000 11.600 206.800 11.700 ;
        RECT 281.200 11.600 282.000 11.700 ;
        RECT 305.200 12.300 306.000 12.400 ;
        RECT 319.600 12.300 320.400 12.400 ;
        RECT 305.200 11.700 320.400 12.300 ;
        RECT 305.200 11.600 306.000 11.700 ;
        RECT 319.600 11.600 320.400 11.700 ;
        RECT 337.200 12.300 338.000 12.400 ;
        RECT 382.000 12.300 382.800 12.400 ;
        RECT 337.200 11.700 382.800 12.300 ;
        RECT 337.200 11.600 338.000 11.700 ;
        RECT 382.000 11.600 382.800 11.700 ;
        RECT 394.800 12.300 395.600 12.400 ;
        RECT 465.200 12.300 466.000 12.400 ;
        RECT 479.600 12.300 480.400 12.400 ;
        RECT 394.800 11.700 480.400 12.300 ;
        RECT 394.800 11.600 395.600 11.700 ;
        RECT 465.200 11.600 466.000 11.700 ;
        RECT 479.600 11.600 480.400 11.700 ;
        RECT 486.000 12.300 486.800 12.400 ;
        RECT 494.000 12.300 494.800 12.400 ;
        RECT 486.000 11.700 494.800 12.300 ;
        RECT 486.000 11.600 486.800 11.700 ;
        RECT 494.000 11.600 494.800 11.700 ;
        RECT 498.800 12.300 499.600 12.400 ;
        RECT 503.700 12.300 504.300 13.700 ;
        RECT 498.800 11.700 504.300 12.300 ;
        RECT 510.000 12.300 510.800 12.400 ;
        RECT 511.600 12.300 512.400 12.400 ;
        RECT 510.000 11.700 512.400 12.300 ;
        RECT 514.900 12.300 515.500 13.700 ;
        RECT 516.400 13.700 528.400 14.300 ;
        RECT 516.400 13.600 517.200 13.700 ;
        RECT 527.600 13.600 528.400 13.700 ;
        RECT 529.200 14.300 530.000 14.400 ;
        RECT 534.000 14.300 534.800 14.400 ;
        RECT 543.600 14.300 544.400 14.400 ;
        RECT 529.200 13.700 544.400 14.300 ;
        RECT 529.200 13.600 530.000 13.700 ;
        RECT 534.000 13.600 534.800 13.700 ;
        RECT 543.600 13.600 544.400 13.700 ;
        RECT 545.200 14.300 546.000 14.400 ;
        RECT 550.000 14.300 550.800 14.400 ;
        RECT 554.800 14.300 555.600 14.400 ;
        RECT 545.200 13.700 555.600 14.300 ;
        RECT 545.200 13.600 546.000 13.700 ;
        RECT 550.000 13.600 550.800 13.700 ;
        RECT 554.800 13.600 555.600 13.700 ;
        RECT 535.600 12.300 536.400 12.400 ;
        RECT 540.400 12.300 541.200 12.400 ;
        RECT 546.800 12.300 547.600 12.400 ;
        RECT 514.900 11.700 547.600 12.300 ;
        RECT 498.800 11.600 499.600 11.700 ;
        RECT 510.000 11.600 510.800 11.700 ;
        RECT 511.600 11.600 512.400 11.700 ;
        RECT 535.600 11.600 536.400 11.700 ;
        RECT 540.400 11.600 541.200 11.700 ;
        RECT 546.800 11.600 547.600 11.700 ;
        RECT 564.400 12.300 565.200 12.400 ;
        RECT 574.000 12.300 574.800 12.400 ;
        RECT 564.400 11.700 574.800 12.300 ;
        RECT 564.400 11.600 565.200 11.700 ;
        RECT 574.000 11.600 574.800 11.700 ;
        RECT 9.200 10.300 10.000 10.400 ;
        RECT 15.600 10.300 16.400 10.400 ;
        RECT 9.200 9.700 16.400 10.300 ;
        RECT 9.200 9.600 10.000 9.700 ;
        RECT 15.600 9.600 16.400 9.700 ;
        RECT 34.800 10.300 35.600 10.400 ;
        RECT 82.800 10.300 83.600 10.400 ;
        RECT 34.800 9.700 83.600 10.300 ;
        RECT 34.800 9.600 35.600 9.700 ;
        RECT 82.800 9.600 83.600 9.700 ;
        RECT 172.400 10.300 173.200 10.400 ;
        RECT 278.000 10.300 278.800 10.400 ;
        RECT 302.000 10.300 302.800 10.400 ;
        RECT 172.400 9.700 302.800 10.300 ;
        RECT 172.400 9.600 173.200 9.700 ;
        RECT 278.000 9.600 278.800 9.700 ;
        RECT 302.000 9.600 302.800 9.700 ;
        RECT 412.400 10.300 413.200 10.400 ;
        RECT 462.000 10.300 462.800 10.400 ;
        RECT 468.400 10.300 469.200 10.400 ;
        RECT 412.400 9.700 469.200 10.300 ;
        RECT 412.400 9.600 413.200 9.700 ;
        RECT 462.000 9.600 462.800 9.700 ;
        RECT 468.400 9.600 469.200 9.700 ;
        RECT 476.400 10.300 477.200 10.400 ;
        RECT 521.200 10.300 522.000 10.400 ;
        RECT 553.200 10.300 554.000 10.400 ;
        RECT 556.400 10.300 557.200 10.400 ;
        RECT 561.200 10.300 562.000 10.400 ;
        RECT 476.400 9.700 562.000 10.300 ;
        RECT 476.400 9.600 477.200 9.700 ;
        RECT 521.200 9.600 522.000 9.700 ;
        RECT 553.200 9.600 554.000 9.700 ;
        RECT 556.400 9.600 557.200 9.700 ;
        RECT 561.200 9.600 562.000 9.700 ;
        RECT 577.200 10.300 578.000 10.400 ;
        RECT 580.400 10.300 581.200 10.400 ;
        RECT 577.200 9.700 581.200 10.300 ;
        RECT 577.200 9.600 578.000 9.700 ;
        RECT 580.400 9.600 581.200 9.700 ;
        RECT 7.600 8.300 8.400 8.400 ;
        RECT 10.800 8.300 11.600 8.400 ;
        RECT 7.600 7.700 11.600 8.300 ;
        RECT 7.600 7.600 8.400 7.700 ;
        RECT 10.800 7.600 11.600 7.700 ;
        RECT 23.600 8.300 24.400 8.400 ;
        RECT 44.400 8.300 45.200 8.400 ;
        RECT 23.600 7.700 45.200 8.300 ;
        RECT 23.600 7.600 24.400 7.700 ;
        RECT 44.400 7.600 45.200 7.700 ;
        RECT 201.200 8.300 202.000 8.400 ;
        RECT 209.200 8.300 210.000 8.400 ;
        RECT 225.200 8.300 226.000 8.400 ;
        RECT 201.200 7.700 226.000 8.300 ;
        RECT 201.200 7.600 202.000 7.700 ;
        RECT 209.200 7.600 210.000 7.700 ;
        RECT 225.200 7.600 226.000 7.700 ;
        RECT 226.800 8.300 227.600 8.400 ;
        RECT 239.600 8.300 240.400 8.400 ;
        RECT 226.800 7.700 240.400 8.300 ;
        RECT 226.800 7.600 227.600 7.700 ;
        RECT 239.600 7.600 240.400 7.700 ;
        RECT 242.800 8.300 243.600 8.400 ;
        RECT 252.400 8.300 253.200 8.400 ;
        RECT 242.800 7.700 253.200 8.300 ;
        RECT 242.800 7.600 243.600 7.700 ;
        RECT 252.400 7.600 253.200 7.700 ;
        RECT 255.600 8.300 256.400 8.400 ;
        RECT 265.200 8.300 266.000 8.400 ;
        RECT 255.600 7.700 266.000 8.300 ;
        RECT 255.600 7.600 256.400 7.700 ;
        RECT 265.200 7.600 266.000 7.700 ;
        RECT 271.600 8.300 272.400 8.400 ;
        RECT 362.800 8.300 363.600 8.400 ;
        RECT 271.600 7.700 363.600 8.300 ;
        RECT 271.600 7.600 272.400 7.700 ;
        RECT 362.800 7.600 363.600 7.700 ;
        RECT 425.200 8.300 426.000 8.400 ;
        RECT 430.000 8.300 430.800 8.400 ;
        RECT 425.200 7.700 430.800 8.300 ;
        RECT 425.200 7.600 426.000 7.700 ;
        RECT 430.000 7.600 430.800 7.700 ;
        RECT 201.200 6.300 202.000 6.400 ;
        RECT 233.200 6.300 234.000 6.400 ;
        RECT 201.200 5.700 234.000 6.300 ;
        RECT 201.200 5.600 202.000 5.700 ;
        RECT 233.200 5.600 234.000 5.700 ;
        RECT 239.600 6.300 240.400 6.400 ;
        RECT 343.600 6.300 344.400 6.400 ;
        RECT 239.600 5.700 344.400 6.300 ;
        RECT 239.600 5.600 240.400 5.700 ;
        RECT 343.600 5.600 344.400 5.700 ;
      LAYER metal4 ;
        RECT 5.800 349.400 7.000 366.600 ;
        RECT 31.400 335.400 32.600 376.600 ;
        RECT 2.600 99.400 3.800 224.600 ;
        RECT 5.800 211.400 7.000 298.600 ;
        RECT 12.200 175.400 13.400 310.600 ;
        RECT 18.600 293.400 19.800 314.600 ;
        RECT 37.800 295.400 39.000 412.600 ;
        RECT 201.000 397.400 202.200 402.600 ;
        RECT 63.400 371.400 64.600 380.600 ;
        RECT 47.400 317.400 48.600 348.600 ;
        RECT 15.400 255.400 16.600 272.600 ;
        RECT 47.400 253.400 48.600 298.600 ;
        RECT 53.800 267.400 55.000 296.600 ;
        RECT 57.000 219.400 58.200 332.600 ;
        RECT 60.200 307.400 61.400 330.600 ;
        RECT 79.400 307.400 80.600 348.600 ;
        RECT 89.000 309.400 90.200 378.600 ;
        RECT 60.200 253.400 61.400 270.600 ;
        RECT 76.200 227.400 77.400 298.600 ;
        RECT 89.000 255.400 90.200 292.600 ;
        RECT 92.200 283.400 93.400 312.600 ;
        RECT 98.600 279.400 99.800 364.600 ;
        RECT 108.200 293.400 109.400 300.600 ;
        RECT 114.600 289.400 115.800 392.600 ;
        RECT 117.800 295.400 119.000 300.600 ;
        RECT 121.000 285.400 122.200 294.600 ;
        RECT 124.200 293.400 125.400 388.600 ;
        RECT 191.400 365.400 192.600 386.600 ;
        RECT 197.800 353.400 199.000 390.600 ;
        RECT 226.600 373.400 227.800 392.600 ;
        RECT 242.600 377.400 243.800 404.600 ;
        RECT 287.400 359.400 288.600 384.600 ;
        RECT 434.600 371.400 435.800 380.600 ;
        RECT 268.200 355.400 271.000 356.600 ;
        RECT 121.000 227.400 122.200 272.600 ;
        RECT 12.200 91.400 13.400 154.600 ;
        RECT 28.200 29.400 29.400 140.600 ;
        RECT 34.600 79.400 35.800 194.600 ;
        RECT 57.000 95.400 64.600 96.600 ;
        RECT 63.400 93.400 64.600 95.400 ;
        RECT 69.800 93.400 71.000 136.600 ;
        RECT 37.800 31.400 39.000 88.600 ;
        RECT 50.600 49.400 51.800 90.600 ;
        RECT 76.200 71.400 77.400 112.600 ;
        RECT 89.000 111.400 90.200 222.600 ;
        RECT 92.200 105.400 93.400 224.600 ;
        RECT 127.400 211.400 128.600 316.600 ;
        RECT 130.600 273.400 131.800 284.600 ;
        RECT 98.600 141.400 99.800 188.600 ;
        RECT 95.400 67.400 96.600 126.600 ;
        RECT 111.400 125.400 112.600 204.600 ;
        RECT 143.400 189.400 144.600 248.600 ;
        RECT 146.600 247.400 147.800 324.600 ;
        RECT 233.000 317.400 234.200 352.600 ;
        RECT 268.200 351.400 269.400 355.400 ;
        RECT 153.000 287.400 154.200 308.600 ;
        RECT 156.200 289.400 157.400 302.600 ;
        RECT 386.600 293.400 387.800 336.600 ;
        RECT 396.200 289.400 397.400 340.600 ;
        RECT 412.200 315.400 413.400 364.600 ;
        RECT 437.800 333.400 439.000 400.600 ;
        RECT 460.200 313.400 461.400 334.600 ;
        RECT 463.400 327.400 464.600 404.600 ;
        RECT 473.000 357.400 474.200 400.600 ;
        RECT 511.400 337.400 512.600 380.600 ;
        RECT 514.600 349.400 515.800 384.600 ;
        RECT 146.600 189.400 147.800 244.600 ;
        RECT 156.200 233.400 157.400 272.600 ;
        RECT 303.400 267.400 307.800 268.600 ;
        RECT 303.400 265.400 304.600 267.400 ;
        RECT 306.600 265.400 307.800 267.400 ;
        RECT 322.600 249.400 323.800 254.600 ;
        RECT 437.800 225.400 439.000 272.600 ;
        RECT 284.200 217.400 285.400 224.600 ;
        RECT 457.000 213.400 458.200 248.600 ;
        RECT 463.400 211.400 464.600 260.600 ;
        RECT 101.800 103.400 103.000 122.600 ;
        RECT 101.800 81.400 103.000 98.600 ;
        RECT 105.000 91.400 106.200 98.600 ;
        RECT 143.400 89.400 144.600 94.600 ;
        RECT 98.600 49.400 99.800 68.600 ;
        RECT 63.400 11.400 64.600 20.600 ;
        RECT 101.800 17.400 103.000 68.600 ;
        RECT 146.600 59.400 147.800 90.600 ;
        RECT 149.800 63.400 151.000 184.600 ;
        RECT 156.200 131.400 157.400 136.600 ;
        RECT 213.800 133.400 215.000 150.600 ;
        RECT 223.400 117.400 224.600 140.600 ;
        RECT 172.200 9.400 173.400 64.600 ;
        RECT 217.000 55.400 218.200 98.600 ;
        RECT 261.800 65.400 263.000 134.600 ;
        RECT 268.200 133.400 269.400 162.600 ;
        RECT 274.600 97.400 275.800 120.600 ;
        RECT 287.400 101.400 288.600 130.600 ;
        RECT 306.600 125.400 307.800 170.600 ;
        RECT 277.800 59.400 279.000 96.600 ;
        RECT 281.000 63.400 282.200 68.600 ;
        RECT 281.000 53.400 282.200 58.600 ;
        RECT 297.000 49.400 298.200 94.600 ;
        RECT 300.200 53.400 301.400 64.600 ;
        RECT 303.400 53.400 304.600 92.600 ;
        RECT 197.800 17.400 199.000 30.600 ;
        RECT 223.400 13.400 224.600 30.600 ;
        RECT 226.600 27.400 227.800 36.600 ;
        RECT 239.400 7.400 240.600 32.600 ;
        RECT 245.800 13.400 247.000 34.600 ;
        RECT 249.000 13.400 250.200 34.600 ;
        RECT 252.200 17.400 253.400 32.600 ;
        RECT 284.200 27.400 285.400 32.600 ;
        RECT 306.600 27.400 307.800 70.600 ;
        RECT 329.000 63.400 330.200 96.600 ;
        RECT 341.800 91.400 343.000 138.600 ;
        RECT 345.000 127.400 346.200 154.600 ;
        RECT 357.800 127.400 359.000 174.600 ;
        RECT 409.000 143.400 410.200 172.600 ;
        RECT 367.400 111.400 368.600 136.600 ;
        RECT 431.400 119.400 432.600 170.600 ;
        RECT 453.800 117.400 455.000 192.600 ;
        RECT 409.000 105.400 410.200 110.600 ;
        RECT 460.200 69.400 461.400 112.600 ;
        RECT 463.400 73.400 464.600 98.600 ;
        RECT 473.000 95.400 474.200 152.600 ;
        RECT 492.200 149.400 493.400 228.600 ;
        RECT 508.200 211.400 509.400 252.600 ;
        RECT 508.200 117.400 509.400 170.600 ;
        RECT 476.200 97.400 477.400 114.600 ;
        RECT 479.400 71.400 480.600 100.600 ;
        RECT 434.600 53.400 435.800 66.600 ;
        RECT 265.000 17.400 266.200 22.600 ;
        RECT 268.200 12.600 269.400 16.600 ;
        RECT 265.000 11.400 269.400 12.600 ;
        RECT 265.000 7.400 266.200 11.400 ;
        RECT 425.000 7.400 426.200 38.600 ;
        RECT 428.200 19.400 429.400 36.600 ;
        RECT 434.600 19.400 435.800 34.600 ;
        RECT 437.800 19.400 439.000 52.600 ;
        RECT 495.400 49.400 496.600 72.600 ;
        RECT 498.600 65.400 499.800 70.600 ;
        RECT 508.200 53.400 509.400 68.600 ;
        RECT 450.600 25.400 451.800 46.600 ;
        RECT 460.200 36.600 461.400 38.600 ;
        RECT 458.600 35.400 461.400 36.600 ;
        RECT 473.000 29.400 474.200 38.600 ;
        RECT 508.200 21.400 509.400 26.600 ;
        RECT 511.400 11.400 512.600 30.600 ;
        RECT 517.800 21.400 519.000 364.600 ;
        RECT 530.600 151.400 531.800 170.600 ;
        RECT 521.000 51.400 522.200 110.600 ;
        RECT 527.400 49.400 528.600 116.600 ;
        RECT 537.000 115.400 538.200 334.600 ;
        RECT 553.000 163.400 554.200 324.600 ;
        RECT 540.200 63.400 541.400 124.600 ;
        RECT 549.800 49.400 551.000 142.600 ;
        RECT 553.000 43.400 554.200 146.600 ;
        RECT 562.600 107.400 563.800 278.600 ;
        RECT 565.800 183.400 567.000 332.600 ;
        RECT 578.600 117.400 579.800 296.600 ;
        RECT 569.000 19.400 570.200 30.600 ;
        RECT 575.400 21.400 576.600 52.600 ;
        RECT 581.800 27.400 583.000 304.600 ;
  END
END sincos
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cordic
  CLASS BLOCK ;
  FOREIGN cordic ;
  ORIGIN 1.900 4.000 ;
  SIZE 224.600 BY 208.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.400 200.400 220.400 201.600 ;
        RECT 2.800 193.000 3.600 200.400 ;
        RECT 7.800 199.800 8.600 200.400 ;
        RECT 7.600 193.200 8.600 199.800 ;
        RECT 13.800 193.200 14.800 200.400 ;
        RECT 17.200 195.800 18.000 200.400 ;
        RECT 30.000 193.800 30.800 200.400 ;
        RECT 33.200 191.800 34.000 200.400 ;
        RECT 37.400 195.800 38.200 200.400 ;
        RECT 41.200 193.000 42.000 200.400 ;
        RECT 44.400 195.800 45.200 200.400 ;
        RECT 47.600 195.800 48.400 200.400 ;
        RECT 50.800 196.200 51.600 200.400 ;
        RECT 55.600 195.800 56.400 200.400 ;
        RECT 57.200 195.800 58.000 200.400 ;
        RECT 60.400 195.800 61.200 200.400 ;
        RECT 66.800 195.800 67.600 200.400 ;
        RECT 70.000 195.800 70.800 200.400 ;
        RECT 73.200 195.800 74.000 200.400 ;
        RECT 76.400 195.800 77.200 200.400 ;
        RECT 84.400 195.800 85.200 200.400 ;
        RECT 87.600 195.800 88.400 200.400 ;
        RECT 94.000 195.800 94.800 200.400 ;
        RECT 97.200 195.800 98.000 200.400 ;
        RECT 100.400 195.800 101.200 200.400 ;
        RECT 103.600 193.000 104.400 200.400 ;
        RECT 106.800 195.800 107.600 200.400 ;
        RECT 110.000 195.800 110.800 200.400 ;
        RECT 113.200 195.800 114.000 200.400 ;
        RECT 119.600 195.800 120.400 200.400 ;
        RECT 122.800 195.800 123.600 200.400 ;
        RECT 130.800 195.800 131.600 200.400 ;
        RECT 134.000 195.800 134.800 200.400 ;
        RECT 137.200 195.800 138.000 200.400 ;
        RECT 140.400 195.800 141.200 200.400 ;
        RECT 143.600 193.000 144.400 200.400 ;
        RECT 148.400 193.200 149.400 200.400 ;
        RECT 154.600 199.800 155.400 200.400 ;
        RECT 154.600 193.200 155.600 199.800 ;
        RECT 164.400 193.000 165.200 200.400 ;
        RECT 167.600 195.800 168.400 200.400 ;
        RECT 93.800 191.800 94.600 192.000 ;
        RECT 97.200 191.800 98.000 192.400 ;
        RECT 71.000 191.200 98.000 191.800 ;
        RECT 110.000 191.800 110.800 192.400 ;
        RECT 113.200 191.800 114.200 192.000 ;
        RECT 170.800 191.800 171.600 200.400 ;
        RECT 175.600 195.800 176.400 200.400 ;
        RECT 178.800 192.200 179.600 200.400 ;
        RECT 182.000 195.800 182.800 200.400 ;
        RECT 185.200 195.800 186.000 200.400 ;
        RECT 188.400 195.800 189.200 200.400 ;
        RECT 194.800 195.800 195.600 200.400 ;
        RECT 198.000 195.800 198.800 200.400 ;
        RECT 206.000 195.800 206.800 200.400 ;
        RECT 209.200 195.800 210.000 200.400 ;
        RECT 212.400 195.800 213.200 200.400 ;
        RECT 215.600 195.800 216.400 200.400 ;
        RECT 185.200 191.800 186.000 192.400 ;
        RECT 188.400 191.800 189.400 192.000 ;
        RECT 110.000 191.200 137.000 191.800 ;
        RECT 185.200 191.200 212.200 191.800 ;
        RECT 71.000 191.000 71.800 191.200 ;
        RECT 136.200 191.000 137.000 191.200 ;
        RECT 211.400 191.000 212.200 191.200 ;
        RECT 10.800 172.000 11.600 172.600 ;
        RECT 28.400 172.000 29.200 172.400 ;
        RECT 33.400 172.000 34.200 172.200 ;
        RECT 10.800 171.400 34.200 172.000 ;
        RECT 133.000 170.800 133.800 171.000 ;
        RECT 106.800 170.200 133.800 170.800 ;
        RECT 1.200 161.600 2.000 166.200 ;
        RECT 4.400 161.600 5.200 166.200 ;
        RECT 7.600 161.600 8.400 166.200 ;
        RECT 10.800 161.600 11.600 166.200 ;
        RECT 18.800 161.600 19.600 166.200 ;
        RECT 22.000 161.600 22.800 166.200 ;
        RECT 28.400 161.600 29.200 166.200 ;
        RECT 31.600 161.600 32.400 166.200 ;
        RECT 34.800 161.600 35.600 166.200 ;
        RECT 38.000 161.600 38.800 169.000 ;
        RECT 42.800 161.600 43.600 165.800 ;
        RECT 46.000 161.600 46.800 166.200 ;
        RECT 49.200 161.600 50.000 166.200 ;
        RECT 52.400 161.600 53.200 166.200 ;
        RECT 54.600 161.600 55.400 166.200 ;
        RECT 58.800 161.600 59.600 170.200 ;
        RECT 66.800 161.600 67.600 168.200 ;
        RECT 79.600 162.200 80.600 168.800 ;
        RECT 79.800 161.600 80.600 162.200 ;
        RECT 85.800 161.600 86.800 168.800 ;
        RECT 89.200 161.600 90.000 170.200 ;
        RECT 92.400 161.600 93.200 170.200 ;
        RECT 95.600 161.600 96.400 170.200 ;
        RECT 98.800 161.600 99.600 170.200 ;
        RECT 102.000 161.600 102.800 170.200 ;
        RECT 106.800 169.600 107.600 170.200 ;
        RECT 110.200 170.000 111.000 170.200 ;
        RECT 103.600 161.600 104.400 166.200 ;
        RECT 106.800 161.600 107.600 166.200 ;
        RECT 110.000 161.600 110.800 166.200 ;
        RECT 116.400 161.600 117.200 166.200 ;
        RECT 119.600 161.600 120.400 166.200 ;
        RECT 127.600 161.600 128.400 166.200 ;
        RECT 130.800 161.600 131.600 166.200 ;
        RECT 134.000 161.600 134.800 166.200 ;
        RECT 137.200 161.600 138.000 166.200 ;
        RECT 140.400 161.600 141.200 169.000 ;
        RECT 145.200 162.200 146.200 168.800 ;
        RECT 145.400 161.600 146.200 162.200 ;
        RECT 151.400 161.600 152.400 168.800 ;
        RECT 159.600 161.600 160.400 166.200 ;
        RECT 162.800 161.600 163.600 166.200 ;
        RECT 166.000 161.600 166.800 166.200 ;
        RECT 169.200 161.600 170.200 168.800 ;
        RECT 175.400 162.200 176.400 168.800 ;
        RECT 175.400 161.600 176.200 162.200 ;
        RECT 178.800 161.600 179.600 166.200 ;
        RECT 182.000 161.600 182.800 166.200 ;
        RECT 186.800 161.600 187.600 170.200 ;
        RECT 190.000 161.600 190.800 166.200 ;
        RECT 193.200 162.200 194.200 168.800 ;
        RECT 193.400 161.600 194.200 162.200 ;
        RECT 199.400 161.600 200.400 168.800 ;
        RECT 204.400 161.600 205.200 169.800 ;
        RECT 207.600 161.600 208.400 166.200 ;
        RECT 210.800 161.600 211.600 169.000 ;
        RECT 215.600 161.600 216.400 169.000 ;
        RECT 0.400 160.400 220.400 161.600 ;
        RECT 2.800 153.000 3.600 160.400 ;
        RECT 7.600 153.000 8.400 160.400 ;
        RECT 10.800 155.800 11.600 160.400 ;
        RECT 14.000 155.800 14.800 160.400 ;
        RECT 17.200 155.800 18.000 160.400 ;
        RECT 20.400 156.200 21.200 160.400 ;
        RECT 23.600 155.800 24.400 160.400 ;
        RECT 26.800 155.800 27.600 160.400 ;
        RECT 29.000 155.800 29.800 160.400 ;
        RECT 33.200 151.800 34.000 160.400 ;
        RECT 34.800 155.800 35.600 160.400 ;
        RECT 38.000 155.800 38.800 160.400 ;
        RECT 39.600 155.800 40.400 160.400 ;
        RECT 42.800 155.800 43.600 160.400 ;
        RECT 46.000 155.800 46.800 160.400 ;
        RECT 52.400 155.600 53.200 160.400 ;
        RECT 55.600 155.800 56.400 160.400 ;
        RECT 63.600 155.800 64.400 160.400 ;
        RECT 66.800 155.800 67.600 160.400 ;
        RECT 70.000 155.800 70.800 160.400 ;
        RECT 73.200 155.800 74.000 160.400 ;
        RECT 79.600 155.800 80.400 160.400 ;
        RECT 82.800 155.800 83.600 160.400 ;
        RECT 86.000 155.800 86.800 160.400 ;
        RECT 92.400 155.600 93.200 160.400 ;
        RECT 95.600 155.800 96.400 160.400 ;
        RECT 103.600 155.800 104.400 160.400 ;
        RECT 106.800 155.800 107.600 160.400 ;
        RECT 110.000 155.800 110.800 160.400 ;
        RECT 113.200 155.800 114.000 160.400 ;
        RECT 114.800 151.800 115.600 160.400 ;
        RECT 118.000 151.800 118.800 160.400 ;
        RECT 121.200 151.800 122.000 160.400 ;
        RECT 124.400 151.800 125.200 160.400 ;
        RECT 127.600 151.800 128.400 160.400 ;
        RECT 129.200 155.800 130.000 160.400 ;
        RECT 132.400 155.800 133.200 160.400 ;
        RECT 135.600 155.800 136.400 160.400 ;
        RECT 142.000 155.800 142.800 160.400 ;
        RECT 145.200 155.800 146.000 160.400 ;
        RECT 153.200 155.800 154.000 160.400 ;
        RECT 156.400 155.800 157.200 160.400 ;
        RECT 159.600 155.800 160.400 160.400 ;
        RECT 162.800 155.800 163.600 160.400 ;
        RECT 169.200 155.800 170.000 160.400 ;
        RECT 172.400 155.800 173.200 160.400 ;
        RECT 174.000 155.800 174.800 160.400 ;
        RECT 177.200 155.800 178.000 160.400 ;
        RECT 180.400 155.800 181.200 160.400 ;
        RECT 186.800 155.800 187.600 160.400 ;
        RECT 190.000 155.800 190.800 160.400 ;
        RECT 198.000 155.800 198.800 160.400 ;
        RECT 201.200 155.800 202.000 160.400 ;
        RECT 204.400 155.800 205.200 160.400 ;
        RECT 207.600 155.800 208.400 160.400 ;
        RECT 210.800 153.000 211.600 160.400 ;
        RECT 215.600 153.000 216.400 160.400 ;
        RECT 132.400 151.800 133.200 152.400 ;
        RECT 135.600 151.800 136.600 152.000 ;
        RECT 177.200 151.800 178.000 152.400 ;
        RECT 180.400 151.800 181.400 152.000 ;
        RECT 132.400 151.200 159.400 151.800 ;
        RECT 177.200 151.200 204.200 151.800 ;
        RECT 158.600 151.000 159.400 151.200 ;
        RECT 203.400 151.000 204.200 151.200 ;
        RECT 41.000 150.000 64.400 150.600 ;
        RECT 41.000 149.800 41.800 150.000 ;
        RECT 46.000 149.600 46.800 150.000 ;
        RECT 52.400 149.600 53.200 150.000 ;
        RECT 63.600 149.400 64.400 150.000 ;
        RECT 81.000 150.000 104.400 150.600 ;
        RECT 81.000 149.800 81.800 150.000 ;
        RECT 86.000 149.600 86.800 150.000 ;
        RECT 92.400 149.600 93.200 150.000 ;
        RECT 103.600 149.400 104.400 150.000 ;
        RECT 74.800 132.000 75.600 132.600 ;
        RECT 92.400 132.000 93.200 132.400 ;
        RECT 97.400 132.000 98.200 132.200 ;
        RECT 74.800 131.400 98.200 132.000 ;
        RECT 5.400 130.800 6.200 131.000 ;
        RECT 163.400 130.800 164.200 131.000 ;
        RECT 5.400 130.200 32.400 130.800 ;
        RECT 137.200 130.200 164.200 130.800 ;
        RECT 28.200 130.000 29.000 130.200 ;
        RECT 31.600 129.600 32.400 130.200 ;
        RECT 1.200 121.600 2.000 126.200 ;
        RECT 4.400 121.600 5.200 126.200 ;
        RECT 7.600 121.600 8.400 126.200 ;
        RECT 10.800 121.600 11.600 126.200 ;
        RECT 18.800 121.600 19.600 126.200 ;
        RECT 22.000 121.600 22.800 126.200 ;
        RECT 28.400 121.600 29.200 126.200 ;
        RECT 31.600 121.600 32.400 126.200 ;
        RECT 34.800 121.600 35.600 126.200 ;
        RECT 38.000 121.600 38.800 128.200 ;
        RECT 50.800 122.200 51.800 128.800 ;
        RECT 51.000 121.600 51.800 122.200 ;
        RECT 57.000 121.600 58.000 128.800 ;
        RECT 65.200 121.600 66.000 126.200 ;
        RECT 68.400 121.600 69.200 126.200 ;
        RECT 71.600 121.600 72.400 126.200 ;
        RECT 74.800 121.600 75.600 126.200 ;
        RECT 82.800 121.600 83.600 126.200 ;
        RECT 86.000 121.600 86.800 126.200 ;
        RECT 92.400 121.600 93.200 126.200 ;
        RECT 95.600 121.600 96.400 126.200 ;
        RECT 98.800 121.600 99.600 126.200 ;
        RECT 102.000 121.600 103.000 128.800 ;
        RECT 108.200 122.200 109.200 128.800 ;
        RECT 108.200 121.600 109.000 122.200 ;
        RECT 111.600 121.600 112.400 130.200 ;
        RECT 137.200 129.600 138.000 130.200 ;
        RECT 140.400 130.000 141.400 130.200 ;
        RECT 114.800 121.600 115.600 129.000 ;
        RECT 118.000 121.600 118.800 126.200 ;
        RECT 121.200 121.600 122.000 126.200 ;
        RECT 124.400 121.600 125.400 128.800 ;
        RECT 130.600 122.200 131.600 128.800 ;
        RECT 130.600 121.600 131.400 122.200 ;
        RECT 134.000 121.600 134.800 126.200 ;
        RECT 137.200 121.600 138.000 126.200 ;
        RECT 140.400 121.600 141.200 126.200 ;
        RECT 146.800 121.600 147.600 126.200 ;
        RECT 150.000 121.600 150.800 126.200 ;
        RECT 158.000 121.600 158.800 126.200 ;
        RECT 161.200 121.600 162.000 126.200 ;
        RECT 164.400 121.600 165.200 126.200 ;
        RECT 167.600 121.600 168.400 126.200 ;
        RECT 175.600 121.600 176.600 128.800 ;
        RECT 181.800 122.200 182.800 128.800 ;
        RECT 181.800 121.600 182.600 122.200 ;
        RECT 188.400 121.600 189.200 130.200 ;
        RECT 191.600 121.600 192.400 125.800 ;
        RECT 194.800 121.600 195.600 126.200 ;
        RECT 198.000 122.200 199.000 128.800 ;
        RECT 198.200 121.600 199.000 122.200 ;
        RECT 204.200 121.600 205.200 128.800 ;
        RECT 207.600 121.600 208.400 126.200 ;
        RECT 210.800 121.600 211.600 126.200 ;
        RECT 214.000 121.600 214.800 129.000 ;
        RECT 0.400 120.400 220.400 121.600 ;
        RECT 2.800 113.000 3.600 120.400 ;
        RECT 7.600 113.000 8.400 120.400 ;
        RECT 12.400 113.200 13.400 120.400 ;
        RECT 18.600 119.800 19.400 120.400 ;
        RECT 18.600 113.200 19.600 119.800 ;
        RECT 22.000 115.800 22.800 120.400 ;
        RECT 25.200 115.800 26.000 120.400 ;
        RECT 28.400 115.800 29.200 120.400 ;
        RECT 31.600 116.200 32.400 120.400 ;
        RECT 36.400 113.000 37.200 120.400 ;
        RECT 39.600 111.800 40.400 120.400 ;
        RECT 42.800 111.800 43.600 120.400 ;
        RECT 46.000 111.800 46.800 120.400 ;
        RECT 49.200 113.000 50.000 120.400 ;
        RECT 52.400 111.800 53.200 120.400 ;
        RECT 58.800 115.800 59.600 120.400 ;
        RECT 62.000 115.800 62.800 120.400 ;
        RECT 65.200 115.800 66.000 120.400 ;
        RECT 68.400 115.800 69.200 120.400 ;
        RECT 76.400 115.800 77.200 120.400 ;
        RECT 79.600 115.800 80.400 120.400 ;
        RECT 86.000 115.800 86.800 120.400 ;
        RECT 89.200 115.800 90.000 120.400 ;
        RECT 92.400 115.800 93.200 120.400 ;
        RECT 94.000 115.800 94.800 120.400 ;
        RECT 97.200 115.800 98.000 120.400 ;
        RECT 100.400 115.800 101.200 120.400 ;
        RECT 103.600 115.800 104.400 120.400 ;
        RECT 111.600 115.800 112.400 120.400 ;
        RECT 114.800 115.800 115.600 120.400 ;
        RECT 121.200 115.800 122.000 120.400 ;
        RECT 124.400 115.800 125.200 120.400 ;
        RECT 127.600 115.800 128.400 120.400 ;
        RECT 130.800 113.000 131.600 120.400 ;
        RECT 85.800 111.800 86.600 112.000 ;
        RECT 89.200 111.800 90.000 112.400 ;
        RECT 121.000 111.800 122.000 112.000 ;
        RECT 124.400 111.800 125.200 112.400 ;
        RECT 134.000 111.800 134.800 120.400 ;
        RECT 135.600 115.800 136.400 120.400 ;
        RECT 138.800 115.800 139.600 120.400 ;
        RECT 142.000 115.800 142.800 120.400 ;
        RECT 148.400 115.800 149.200 120.400 ;
        RECT 151.600 115.800 152.400 120.400 ;
        RECT 159.600 115.800 160.400 120.400 ;
        RECT 162.800 115.800 163.600 120.400 ;
        RECT 166.000 115.800 166.800 120.400 ;
        RECT 169.200 115.800 170.000 120.400 ;
        RECT 175.600 115.800 176.400 120.400 ;
        RECT 178.800 115.800 179.600 120.400 ;
        RECT 182.000 115.800 182.800 120.400 ;
        RECT 188.400 115.800 189.200 120.400 ;
        RECT 191.600 115.800 192.400 120.400 ;
        RECT 199.600 115.800 200.400 120.400 ;
        RECT 202.800 115.800 203.600 120.400 ;
        RECT 206.000 115.800 206.800 120.400 ;
        RECT 209.200 115.800 210.000 120.400 ;
        RECT 212.400 113.000 213.200 120.400 ;
        RECT 138.800 111.800 139.600 112.400 ;
        RECT 142.200 111.800 143.000 112.000 ;
        RECT 178.800 111.800 179.600 112.400 ;
        RECT 182.200 111.800 183.000 112.000 ;
        RECT 63.000 111.200 90.000 111.800 ;
        RECT 98.200 111.200 125.200 111.800 ;
        RECT 138.800 111.200 165.800 111.800 ;
        RECT 178.800 111.200 205.800 111.800 ;
        RECT 63.000 111.000 63.800 111.200 ;
        RECT 98.200 111.000 99.000 111.200 ;
        RECT 165.000 111.000 165.800 111.200 ;
        RECT 205.000 111.000 205.800 111.200 ;
        RECT 10.800 92.000 11.600 92.600 ;
        RECT 28.400 92.000 29.200 92.400 ;
        RECT 33.400 92.000 34.200 92.200 ;
        RECT 10.800 91.400 34.200 92.000 ;
        RECT 46.000 92.000 46.800 92.600 ;
        RECT 63.600 92.000 64.400 92.400 ;
        RECT 68.600 92.000 69.400 92.200 ;
        RECT 46.000 91.400 69.400 92.000 ;
        RECT 112.600 90.800 113.400 91.000 ;
        RECT 177.800 90.800 178.600 91.000 ;
        RECT 112.600 90.200 139.600 90.800 ;
        RECT 1.200 81.600 2.000 86.200 ;
        RECT 4.400 81.600 5.200 86.200 ;
        RECT 7.600 81.600 8.400 86.200 ;
        RECT 10.800 81.600 11.600 86.200 ;
        RECT 18.800 81.600 19.600 86.200 ;
        RECT 22.000 81.600 22.800 86.200 ;
        RECT 28.400 81.600 29.200 86.200 ;
        RECT 31.600 81.600 32.400 86.200 ;
        RECT 34.800 81.600 35.600 86.200 ;
        RECT 36.400 81.600 37.200 86.200 ;
        RECT 39.600 81.600 40.400 86.200 ;
        RECT 42.800 81.600 43.600 86.200 ;
        RECT 46.000 81.600 46.800 86.200 ;
        RECT 54.000 81.600 54.800 86.200 ;
        RECT 57.200 81.600 58.000 86.200 ;
        RECT 63.600 81.600 64.400 86.200 ;
        RECT 66.800 81.600 67.600 86.200 ;
        RECT 70.000 81.600 70.800 86.200 ;
        RECT 76.400 81.600 77.200 90.200 ;
        RECT 79.600 81.600 80.400 89.000 ;
        RECT 84.400 82.200 85.400 88.800 ;
        RECT 84.600 81.600 85.400 82.200 ;
        RECT 90.600 81.600 91.600 88.800 ;
        RECT 94.000 81.600 94.800 90.200 ;
        RECT 135.400 90.000 136.400 90.200 ;
        RECT 138.800 89.600 139.600 90.200 ;
        RECT 151.600 90.200 178.600 90.800 ;
        RECT 151.600 89.600 152.400 90.200 ;
        RECT 155.000 90.000 155.800 90.200 ;
        RECT 98.200 81.600 99.000 86.200 ;
        RECT 100.400 81.600 101.200 86.200 ;
        RECT 103.600 81.600 104.400 86.200 ;
        RECT 106.800 81.600 107.600 86.200 ;
        RECT 108.400 81.600 109.200 86.200 ;
        RECT 111.600 81.600 112.400 86.200 ;
        RECT 114.800 81.600 115.600 86.200 ;
        RECT 118.000 81.600 118.800 86.200 ;
        RECT 126.000 81.600 126.800 86.200 ;
        RECT 129.200 81.600 130.000 86.200 ;
        RECT 135.600 81.600 136.400 86.200 ;
        RECT 138.800 81.600 139.600 86.200 ;
        RECT 142.000 81.600 142.800 86.200 ;
        RECT 148.400 81.600 149.200 86.200 ;
        RECT 151.600 81.600 152.400 86.200 ;
        RECT 154.800 81.600 155.600 86.200 ;
        RECT 161.200 81.600 162.000 86.200 ;
        RECT 164.400 81.600 165.200 86.200 ;
        RECT 172.400 81.600 173.200 86.200 ;
        RECT 175.600 81.600 176.400 86.200 ;
        RECT 178.800 81.600 179.600 86.200 ;
        RECT 182.000 81.600 182.800 86.200 ;
        RECT 185.200 81.600 186.200 88.800 ;
        RECT 191.400 82.200 192.400 88.800 ;
        RECT 191.400 81.600 192.200 82.200 ;
        RECT 194.800 81.600 195.600 86.200 ;
        RECT 198.000 81.600 198.800 86.200 ;
        RECT 199.600 81.600 200.400 86.200 ;
        RECT 202.800 81.600 203.600 86.200 ;
        RECT 206.000 82.200 207.000 88.800 ;
        RECT 206.200 81.600 207.000 82.200 ;
        RECT 212.200 81.600 213.200 88.800 ;
        RECT 217.200 81.600 218.000 89.000 ;
        RECT 0.400 80.400 220.400 81.600 ;
        RECT 2.800 73.000 3.600 80.400 ;
        RECT 7.600 73.000 8.400 80.400 ;
        RECT 12.400 73.800 13.200 80.400 ;
        RECT 23.600 71.800 24.400 80.400 ;
        RECT 27.800 75.800 28.600 80.400 ;
        RECT 30.000 75.800 30.800 80.400 ;
        RECT 33.200 75.800 34.000 80.400 ;
        RECT 36.600 79.800 37.400 80.400 ;
        RECT 36.400 73.200 37.400 79.800 ;
        RECT 42.600 73.200 43.600 80.400 ;
        RECT 50.800 75.800 51.600 80.400 ;
        RECT 54.000 75.800 54.800 80.400 ;
        RECT 57.200 75.800 58.000 80.400 ;
        RECT 60.400 75.800 61.200 80.400 ;
        RECT 68.400 75.800 69.200 80.400 ;
        RECT 71.600 75.600 72.400 80.400 ;
        RECT 78.000 75.800 78.800 80.400 ;
        RECT 81.200 75.800 82.000 80.400 ;
        RECT 84.400 75.800 85.200 80.400 ;
        RECT 87.600 75.800 88.400 80.400 ;
        RECT 89.200 71.800 90.000 80.400 ;
        RECT 92.400 71.800 93.200 80.400 ;
        RECT 95.600 71.800 96.400 80.400 ;
        RECT 98.800 71.800 99.600 80.400 ;
        RECT 102.000 71.800 102.800 80.400 ;
        RECT 103.600 75.800 104.400 80.400 ;
        RECT 106.800 76.200 107.600 80.400 ;
        RECT 110.000 75.800 110.800 80.400 ;
        RECT 113.200 71.800 114.000 80.400 ;
        RECT 116.400 71.800 117.200 80.400 ;
        RECT 119.600 71.800 120.400 80.400 ;
        RECT 122.800 71.800 123.600 80.400 ;
        RECT 126.000 71.800 126.800 80.400 ;
        RECT 129.200 73.000 130.000 80.400 ;
        RECT 132.400 71.800 133.200 80.400 ;
        RECT 134.000 71.800 134.800 80.400 ;
        RECT 137.200 71.800 138.000 80.400 ;
        RECT 140.400 71.800 141.200 80.400 ;
        RECT 143.600 71.800 144.400 80.400 ;
        RECT 146.800 71.800 147.600 80.400 ;
        RECT 148.400 71.800 149.200 80.400 ;
        RECT 161.200 71.800 162.000 80.400 ;
        RECT 162.800 75.800 163.600 80.400 ;
        RECT 166.000 72.200 166.800 80.400 ;
        RECT 170.800 73.000 171.600 80.400 ;
        RECT 175.800 79.800 176.600 80.400 ;
        RECT 175.600 73.200 176.600 79.800 ;
        RECT 181.800 73.200 182.800 80.400 ;
        RECT 185.200 75.800 186.000 80.400 ;
        RECT 188.400 72.200 189.200 80.400 ;
        RECT 193.200 72.200 194.000 80.400 ;
        RECT 196.400 75.800 197.200 80.400 ;
        RECT 201.200 71.800 202.000 80.400 ;
        RECT 202.800 71.800 203.600 80.400 ;
        RECT 209.200 75.800 210.000 80.400 ;
        RECT 212.400 73.000 213.200 80.400 ;
        RECT 60.400 70.000 83.800 70.600 ;
        RECT 60.400 69.400 61.200 70.000 ;
        RECT 71.600 69.600 72.400 70.000 ;
        RECT 78.000 69.600 78.800 70.000 ;
        RECT 83.000 69.800 83.800 70.000 ;
        RECT 10.800 52.000 11.600 52.600 ;
        RECT 28.400 52.000 29.200 52.400 ;
        RECT 33.400 52.000 34.200 52.200 ;
        RECT 10.800 51.400 34.200 52.000 ;
        RECT 153.800 50.800 154.600 51.000 ;
        RECT 193.800 50.800 194.600 51.000 ;
        RECT 127.600 50.200 154.600 50.800 ;
        RECT 167.600 50.200 194.600 50.800 ;
        RECT 1.200 41.600 2.000 46.200 ;
        RECT 4.400 41.600 5.200 46.200 ;
        RECT 7.600 41.600 8.400 46.200 ;
        RECT 10.800 41.600 11.600 46.200 ;
        RECT 18.800 41.600 19.600 46.200 ;
        RECT 22.000 41.600 22.800 46.200 ;
        RECT 28.400 41.600 29.200 46.200 ;
        RECT 31.600 41.600 32.400 46.200 ;
        RECT 34.800 41.600 35.600 46.200 ;
        RECT 36.400 41.600 37.200 46.200 ;
        RECT 39.600 41.600 40.400 46.200 ;
        RECT 41.200 41.600 42.000 46.200 ;
        RECT 44.400 41.600 45.200 46.200 ;
        RECT 47.600 41.600 48.400 45.800 ;
        RECT 51.400 41.600 52.200 46.200 ;
        RECT 55.600 41.600 56.400 50.200 ;
        RECT 63.600 41.600 64.400 48.200 ;
        RECT 74.800 41.600 75.600 46.200 ;
        RECT 78.000 41.600 78.800 46.200 ;
        RECT 81.200 41.600 82.000 45.800 ;
        RECT 94.000 41.600 94.800 48.200 ;
        RECT 97.200 41.600 98.000 50.200 ;
        RECT 101.400 41.600 102.200 46.200 ;
        RECT 103.600 41.600 104.400 46.200 ;
        RECT 106.800 41.600 107.600 46.200 ;
        RECT 108.400 41.600 109.200 50.200 ;
        RECT 113.200 41.600 114.000 46.200 ;
        RECT 116.400 41.600 117.200 49.800 ;
        RECT 119.600 41.600 120.400 50.200 ;
        RECT 127.600 49.600 128.400 50.200 ;
        RECT 131.000 50.000 131.800 50.200 ;
        RECT 167.600 49.600 168.400 50.200 ;
        RECT 171.000 50.000 171.800 50.200 ;
        RECT 124.400 41.600 125.200 46.200 ;
        RECT 127.600 41.600 128.400 46.200 ;
        RECT 130.800 41.600 131.600 46.200 ;
        RECT 137.200 41.600 138.000 46.200 ;
        RECT 140.400 41.600 141.200 46.200 ;
        RECT 148.400 41.600 149.200 46.200 ;
        RECT 151.600 41.600 152.400 46.200 ;
        RECT 154.800 41.600 155.600 46.200 ;
        RECT 158.000 41.600 158.800 46.200 ;
        RECT 164.400 41.600 165.200 46.200 ;
        RECT 167.600 41.600 168.400 46.200 ;
        RECT 170.800 41.600 171.600 46.200 ;
        RECT 177.200 41.600 178.000 46.200 ;
        RECT 180.400 41.600 181.200 46.200 ;
        RECT 188.400 41.600 189.200 46.200 ;
        RECT 191.600 41.600 192.400 46.200 ;
        RECT 194.800 41.600 195.600 46.200 ;
        RECT 198.000 41.600 198.800 46.200 ;
        RECT 202.800 41.600 203.600 50.200 ;
        RECT 204.400 41.600 205.200 46.200 ;
        RECT 207.600 41.600 208.400 46.200 ;
        RECT 210.800 41.600 211.600 49.000 ;
        RECT 217.200 41.600 218.000 49.000 ;
        RECT 0.400 40.400 220.400 41.600 ;
        RECT 2.800 33.000 3.600 40.400 ;
        RECT 6.000 35.800 6.800 40.400 ;
        RECT 10.800 36.200 11.600 40.400 ;
        RECT 14.000 35.800 14.800 40.400 ;
        RECT 17.200 35.800 18.000 40.400 ;
        RECT 20.400 33.200 21.400 40.400 ;
        RECT 26.600 39.800 27.400 40.400 ;
        RECT 26.600 33.200 27.600 39.800 ;
        RECT 30.000 31.800 30.800 40.400 ;
        RECT 34.200 35.800 35.000 40.400 ;
        RECT 38.000 33.800 38.800 40.400 ;
        RECT 50.800 35.800 51.600 40.400 ;
        RECT 52.400 35.800 53.200 40.400 ;
        RECT 55.600 35.800 56.400 40.400 ;
        RECT 63.800 39.800 64.600 40.400 ;
        RECT 63.600 33.200 64.600 39.800 ;
        RECT 69.800 33.200 70.800 40.400 ;
        RECT 73.200 35.800 74.000 40.400 ;
        RECT 76.400 35.800 77.200 40.400 ;
        RECT 79.600 35.800 80.400 40.400 ;
        RECT 86.000 35.800 86.800 40.400 ;
        RECT 89.200 35.800 90.000 40.400 ;
        RECT 97.200 35.800 98.000 40.400 ;
        RECT 100.400 35.800 101.200 40.400 ;
        RECT 103.600 35.800 104.400 40.400 ;
        RECT 106.800 35.800 107.600 40.400 ;
        RECT 108.400 35.800 109.200 40.400 ;
        RECT 111.600 35.800 112.400 40.400 ;
        RECT 114.800 35.800 115.600 40.400 ;
        RECT 118.000 35.800 118.800 40.400 ;
        RECT 126.000 35.800 126.800 40.400 ;
        RECT 129.200 35.800 130.000 40.400 ;
        RECT 135.600 35.800 136.400 40.400 ;
        RECT 138.800 35.800 139.600 40.400 ;
        RECT 142.000 35.800 142.800 40.400 ;
        RECT 143.600 35.800 144.400 40.400 ;
        RECT 146.800 35.800 147.600 40.400 ;
        RECT 76.400 31.800 77.200 32.400 ;
        RECT 79.600 31.800 80.600 32.000 ;
        RECT 151.600 31.800 152.400 40.400 ;
        RECT 158.000 35.800 158.800 40.400 ;
        RECT 164.400 31.800 165.200 40.400 ;
        RECT 166.000 35.800 166.800 40.400 ;
        RECT 169.200 35.800 170.000 40.400 ;
        RECT 172.400 35.800 173.200 40.400 ;
        RECT 178.800 35.800 179.600 40.400 ;
        RECT 182.000 35.800 182.800 40.400 ;
        RECT 190.000 35.800 190.800 40.400 ;
        RECT 193.200 35.800 194.000 40.400 ;
        RECT 196.400 35.800 197.200 40.400 ;
        RECT 199.600 35.800 200.400 40.400 ;
        RECT 203.000 39.800 203.800 40.400 ;
        RECT 202.800 33.200 203.800 39.800 ;
        RECT 209.000 33.200 210.000 40.400 ;
        RECT 214.000 33.000 214.800 40.400 ;
        RECT 169.200 31.800 170.000 32.400 ;
        RECT 172.400 31.800 173.400 32.000 ;
        RECT 76.400 31.200 103.400 31.800 ;
        RECT 169.200 31.200 196.200 31.800 ;
        RECT 102.600 31.000 103.400 31.200 ;
        RECT 195.400 31.000 196.200 31.200 ;
        RECT 118.000 30.000 141.400 30.600 ;
        RECT 118.000 29.400 118.800 30.000 ;
        RECT 135.600 29.600 136.400 30.000 ;
        RECT 140.600 29.800 141.400 30.000 ;
        RECT 10.200 10.800 11.000 11.000 ;
        RECT 55.000 10.800 55.800 11.000 ;
        RECT 109.400 10.800 110.200 11.000 ;
        RECT 149.400 10.800 150.200 11.000 ;
        RECT 209.800 10.800 210.600 11.000 ;
        RECT 10.200 10.200 37.200 10.800 ;
        RECT 55.000 10.200 82.000 10.800 ;
        RECT 109.400 10.200 136.400 10.800 ;
        RECT 149.400 10.200 176.400 10.800 ;
        RECT 33.000 10.000 33.800 10.200 ;
        RECT 36.400 9.600 37.200 10.200 ;
        RECT 77.800 10.000 78.600 10.200 ;
        RECT 81.200 9.600 82.000 10.200 ;
        RECT 132.200 10.000 133.000 10.200 ;
        RECT 135.600 9.600 136.400 10.200 ;
        RECT 172.200 10.000 173.200 10.200 ;
        RECT 175.600 9.600 176.400 10.200 ;
        RECT 183.600 10.200 210.600 10.800 ;
        RECT 183.600 9.600 184.400 10.200 ;
        RECT 186.800 10.000 187.800 10.200 ;
        RECT 2.800 1.600 3.600 9.000 ;
        RECT 6.000 1.600 6.800 6.200 ;
        RECT 9.200 1.600 10.000 6.200 ;
        RECT 12.400 1.600 13.200 6.200 ;
        RECT 15.600 1.600 16.400 6.200 ;
        RECT 23.600 1.600 24.400 6.200 ;
        RECT 26.800 1.600 27.600 6.200 ;
        RECT 33.200 1.600 34.000 6.200 ;
        RECT 36.400 1.600 37.200 6.200 ;
        RECT 39.600 1.600 40.400 6.200 ;
        RECT 42.800 1.600 43.600 9.000 ;
        RECT 50.800 1.600 51.600 6.200 ;
        RECT 54.000 1.600 54.800 6.200 ;
        RECT 57.200 1.600 58.000 6.200 ;
        RECT 60.400 1.600 61.200 6.200 ;
        RECT 68.400 1.600 69.200 6.200 ;
        RECT 71.600 1.600 72.400 6.200 ;
        RECT 78.000 1.600 78.800 6.200 ;
        RECT 81.200 1.600 82.000 6.200 ;
        RECT 84.400 1.600 85.200 6.200 ;
        RECT 87.600 1.600 88.400 9.000 ;
        RECT 92.400 1.600 93.200 9.000 ;
        RECT 97.200 1.600 98.000 9.000 ;
        RECT 102.000 1.600 102.800 9.000 ;
        RECT 105.200 1.600 106.000 6.200 ;
        RECT 108.400 1.600 109.200 6.200 ;
        RECT 111.600 1.600 112.400 6.200 ;
        RECT 114.800 1.600 115.600 6.200 ;
        RECT 122.800 1.600 123.600 6.200 ;
        RECT 126.000 1.600 126.800 6.200 ;
        RECT 132.400 1.600 133.200 6.200 ;
        RECT 135.600 1.600 136.400 6.200 ;
        RECT 138.800 1.600 139.600 6.200 ;
        RECT 145.200 1.600 146.000 6.200 ;
        RECT 148.400 1.600 149.200 6.200 ;
        RECT 151.600 1.600 152.400 6.200 ;
        RECT 154.800 1.600 155.600 6.200 ;
        RECT 162.800 1.600 163.600 6.200 ;
        RECT 166.000 1.600 166.800 6.200 ;
        RECT 172.400 1.600 173.200 6.200 ;
        RECT 175.600 1.600 176.400 6.200 ;
        RECT 178.800 1.600 179.600 6.200 ;
        RECT 180.400 1.600 181.200 6.200 ;
        RECT 183.600 1.600 184.400 6.200 ;
        RECT 186.800 1.600 187.600 6.200 ;
        RECT 193.200 1.600 194.000 6.200 ;
        RECT 196.400 1.600 197.200 6.200 ;
        RECT 204.400 1.600 205.200 6.200 ;
        RECT 207.600 1.600 208.400 6.200 ;
        RECT 210.800 1.600 211.600 6.200 ;
        RECT 214.000 1.600 214.800 6.200 ;
        RECT 0.400 0.400 220.400 1.600 ;
      LAYER via1 ;
        RECT 59.000 200.600 59.800 201.400 ;
        RECT 60.400 200.600 61.200 201.400 ;
        RECT 61.800 200.600 62.600 201.400 ;
        RECT 97.200 197.600 98.000 198.400 ;
        RECT 97.200 191.600 98.000 192.400 ;
        RECT 113.200 191.200 114.000 192.000 ;
        RECT 188.400 191.200 189.200 192.000 ;
        RECT 10.800 171.600 11.600 172.400 ;
        RECT 10.800 165.400 11.600 166.200 ;
        RECT 106.800 163.600 107.600 164.400 ;
        RECT 59.000 160.600 59.800 161.400 ;
        RECT 60.400 160.600 61.200 161.400 ;
        RECT 61.800 160.600 62.600 161.400 ;
        RECT 135.600 151.200 136.400 152.000 ;
        RECT 180.400 151.200 181.200 152.000 ;
        RECT 74.800 131.600 75.600 132.400 ;
        RECT 31.600 123.600 32.400 124.400 ;
        RECT 74.800 125.400 75.600 126.200 ;
        RECT 140.400 125.400 141.200 126.200 ;
        RECT 59.000 120.600 59.800 121.400 ;
        RECT 60.400 120.600 61.200 121.400 ;
        RECT 61.800 120.600 62.600 121.400 ;
        RECT 89.200 117.600 90.000 118.400 ;
        RECT 89.200 111.600 90.000 112.400 ;
        RECT 121.200 111.200 122.000 112.000 ;
        RECT 138.800 117.600 139.600 118.400 ;
        RECT 178.800 117.600 179.600 118.400 ;
        RECT 138.800 111.600 139.600 112.400 ;
        RECT 178.800 111.600 179.600 112.400 ;
        RECT 10.800 91.600 11.600 92.400 ;
        RECT 46.000 91.600 46.800 92.400 ;
        RECT 10.800 85.400 11.600 86.200 ;
        RECT 46.000 85.400 46.800 86.200 ;
        RECT 135.600 90.000 136.400 90.800 ;
        RECT 135.600 83.600 136.400 84.400 ;
        RECT 151.600 83.600 152.400 84.400 ;
        RECT 59.000 80.600 59.800 81.400 ;
        RECT 60.400 80.600 61.200 81.400 ;
        RECT 61.800 80.600 62.600 81.400 ;
        RECT 10.800 51.600 11.600 52.400 ;
        RECT 10.800 45.400 11.600 46.200 ;
        RECT 127.600 43.600 128.400 44.400 ;
        RECT 167.600 43.600 168.400 44.400 ;
        RECT 59.000 40.600 59.800 41.400 ;
        RECT 60.400 40.600 61.200 41.400 ;
        RECT 61.800 40.600 62.600 41.400 ;
        RECT 79.600 31.200 80.400 32.000 ;
        RECT 172.400 31.200 173.200 32.000 ;
        RECT 118.000 29.600 118.800 30.400 ;
        RECT 172.400 10.000 173.200 10.800 ;
        RECT 36.400 3.600 37.200 4.400 ;
        RECT 81.200 3.600 82.000 4.400 ;
        RECT 135.600 3.600 136.400 4.400 ;
        RECT 172.400 3.600 173.200 4.400 ;
        RECT 186.800 3.600 187.600 4.400 ;
        RECT 59.000 0.600 59.800 1.400 ;
        RECT 60.400 0.600 61.200 1.400 ;
        RECT 61.800 0.600 62.600 1.400 ;
      LAYER metal2 ;
        RECT 58.400 200.600 63.200 201.400 ;
        RECT 97.200 197.600 98.000 198.400 ;
        RECT 97.300 192.400 97.900 197.600 ;
        RECT 113.200 195.800 114.000 196.600 ;
        RECT 188.400 195.800 189.200 196.600 ;
        RECT 97.200 191.600 98.000 192.400 ;
        RECT 113.300 192.000 113.900 195.800 ;
        RECT 188.500 192.000 189.100 195.800 ;
        RECT 113.200 191.200 114.000 192.000 ;
        RECT 188.400 191.200 189.200 192.000 ;
        RECT 10.800 171.600 11.600 172.400 ;
        RECT 10.900 166.200 11.500 171.600 ;
        RECT 106.800 169.600 107.600 170.400 ;
        RECT 10.800 165.400 11.600 166.200 ;
        RECT 106.900 164.400 107.500 169.600 ;
        RECT 106.800 163.600 107.600 164.400 ;
        RECT 58.400 160.600 63.200 161.400 ;
        RECT 52.400 155.600 53.200 156.400 ;
        RECT 92.400 155.600 93.200 156.400 ;
        RECT 135.600 155.800 136.400 156.600 ;
        RECT 180.400 155.800 181.200 156.600 ;
        RECT 52.500 150.400 53.100 155.600 ;
        RECT 92.500 150.400 93.100 155.600 ;
        RECT 135.700 152.000 136.300 155.800 ;
        RECT 180.500 152.000 181.100 155.800 ;
        RECT 135.600 151.200 136.400 152.000 ;
        RECT 180.400 151.200 181.200 152.000 ;
        RECT 52.400 149.600 53.200 150.400 ;
        RECT 92.400 149.600 93.200 150.400 ;
        RECT 74.800 131.600 75.600 132.400 ;
        RECT 31.600 129.600 32.400 130.400 ;
        RECT 31.700 124.400 32.300 129.600 ;
        RECT 74.900 126.200 75.500 131.600 ;
        RECT 140.400 130.000 141.200 130.800 ;
        RECT 140.500 126.200 141.100 130.000 ;
        RECT 74.800 125.400 75.600 126.200 ;
        RECT 140.400 125.400 141.200 126.200 ;
        RECT 31.600 123.600 32.400 124.400 ;
        RECT 58.400 120.600 63.200 121.400 ;
        RECT 89.200 117.600 90.000 118.400 ;
        RECT 138.800 117.600 139.600 118.400 ;
        RECT 178.800 117.600 179.600 118.400 ;
        RECT 89.300 112.400 89.900 117.600 ;
        RECT 121.200 115.800 122.000 116.600 ;
        RECT 89.200 111.600 90.000 112.400 ;
        RECT 121.300 112.000 121.900 115.800 ;
        RECT 138.900 112.400 139.500 117.600 ;
        RECT 178.900 112.400 179.500 117.600 ;
        RECT 121.200 111.200 122.000 112.000 ;
        RECT 138.800 111.600 139.600 112.400 ;
        RECT 178.800 111.600 179.600 112.400 ;
        RECT 10.800 91.600 11.600 92.400 ;
        RECT 46.000 91.600 46.800 92.400 ;
        RECT 10.900 86.200 11.500 91.600 ;
        RECT 46.100 86.200 46.700 91.600 ;
        RECT 135.600 90.000 136.400 90.800 ;
        RECT 10.800 85.400 11.600 86.200 ;
        RECT 46.000 85.400 46.800 86.200 ;
        RECT 135.700 84.400 136.300 90.000 ;
        RECT 151.600 89.600 152.400 90.400 ;
        RECT 151.700 84.400 152.300 89.600 ;
        RECT 135.600 83.600 136.400 84.400 ;
        RECT 151.600 83.600 152.400 84.400 ;
        RECT 58.400 80.600 63.200 81.400 ;
        RECT 71.600 75.600 72.400 76.400 ;
        RECT 71.700 70.400 72.300 75.600 ;
        RECT 71.600 69.600 72.400 70.400 ;
        RECT 10.800 51.600 11.600 52.400 ;
        RECT 10.900 46.200 11.500 51.600 ;
        RECT 127.600 49.600 128.400 50.400 ;
        RECT 167.600 49.600 168.400 50.400 ;
        RECT 10.800 45.400 11.600 46.200 ;
        RECT 127.700 44.400 128.300 49.600 ;
        RECT 167.700 44.400 168.300 49.600 ;
        RECT 127.600 43.600 128.400 44.400 ;
        RECT 167.600 43.600 168.400 44.400 ;
        RECT 58.400 40.600 63.200 41.400 ;
        RECT 79.600 35.800 80.400 36.600 ;
        RECT 118.000 35.800 118.800 36.600 ;
        RECT 172.400 35.800 173.200 36.600 ;
        RECT 79.700 32.000 80.300 35.800 ;
        RECT 79.600 31.200 80.400 32.000 ;
        RECT 118.100 30.400 118.700 35.800 ;
        RECT 172.500 32.000 173.100 35.800 ;
        RECT 172.400 31.200 173.200 32.000 ;
        RECT 118.000 29.600 118.800 30.400 ;
        RECT 36.400 9.600 37.200 10.400 ;
        RECT 81.200 9.600 82.000 10.400 ;
        RECT 135.600 9.600 136.400 10.400 ;
        RECT 172.400 10.000 173.200 10.800 ;
        RECT 186.800 10.000 187.600 10.800 ;
        RECT 36.500 4.400 37.100 9.600 ;
        RECT 81.300 4.400 81.900 9.600 ;
        RECT 135.700 4.400 136.300 9.600 ;
        RECT 172.500 4.400 173.100 10.000 ;
        RECT 186.900 4.400 187.500 10.000 ;
        RECT 36.400 3.600 37.200 4.400 ;
        RECT 81.200 3.600 82.000 4.400 ;
        RECT 135.600 3.600 136.400 4.400 ;
        RECT 172.400 3.600 173.200 4.400 ;
        RECT 186.800 3.600 187.600 4.400 ;
        RECT 58.400 0.600 63.200 1.400 ;
      LAYER via2 ;
        RECT 59.000 200.600 59.800 201.400 ;
        RECT 60.400 200.600 61.200 201.400 ;
        RECT 61.800 200.600 62.600 201.400 ;
        RECT 59.000 160.600 59.800 161.400 ;
        RECT 60.400 160.600 61.200 161.400 ;
        RECT 61.800 160.600 62.600 161.400 ;
        RECT 59.000 120.600 59.800 121.400 ;
        RECT 60.400 120.600 61.200 121.400 ;
        RECT 61.800 120.600 62.600 121.400 ;
        RECT 59.000 80.600 59.800 81.400 ;
        RECT 60.400 80.600 61.200 81.400 ;
        RECT 61.800 80.600 62.600 81.400 ;
        RECT 59.000 40.600 59.800 41.400 ;
        RECT 60.400 40.600 61.200 41.400 ;
        RECT 61.800 40.600 62.600 41.400 ;
        RECT 59.000 0.600 59.800 1.400 ;
        RECT 60.400 0.600 61.200 1.400 ;
        RECT 61.800 0.600 62.600 1.400 ;
      LAYER metal3 ;
        RECT 58.400 200.400 63.200 201.600 ;
        RECT 58.400 160.400 63.200 161.600 ;
        RECT 58.400 120.400 63.200 121.600 ;
        RECT 58.400 80.400 63.200 81.600 ;
        RECT 58.400 40.400 63.200 41.600 ;
        RECT 58.400 0.400 63.200 1.600 ;
      LAYER via3 ;
        RECT 58.800 200.600 59.600 201.400 ;
        RECT 60.400 200.600 61.200 201.400 ;
        RECT 62.000 200.600 62.800 201.400 ;
        RECT 58.800 160.600 59.600 161.400 ;
        RECT 60.400 160.600 61.200 161.400 ;
        RECT 62.000 160.600 62.800 161.400 ;
        RECT 58.800 120.600 59.600 121.400 ;
        RECT 60.400 120.600 61.200 121.400 ;
        RECT 62.000 120.600 62.800 121.400 ;
        RECT 58.800 80.600 59.600 81.400 ;
        RECT 60.400 80.600 61.200 81.400 ;
        RECT 62.000 80.600 62.800 81.400 ;
        RECT 58.800 40.600 59.600 41.400 ;
        RECT 60.400 40.600 61.200 41.400 ;
        RECT 62.000 40.600 62.800 41.400 ;
        RECT 58.800 0.600 59.600 1.400 ;
        RECT 60.400 0.600 61.200 1.400 ;
        RECT 62.000 0.600 62.800 1.400 ;
      LAYER metal4 ;
        RECT 58.400 -4.000 63.200 204.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 2.800 181.600 3.600 186.200 ;
        RECT 7.600 182.200 8.600 185.600 ;
        RECT 7.800 181.600 8.600 182.200 ;
        RECT 13.800 181.600 14.800 185.600 ;
        RECT 17.200 181.600 18.000 184.200 ;
        RECT 26.800 181.600 27.600 183.800 ;
        RECT 30.000 181.600 30.800 184.200 ;
        RECT 34.800 181.600 35.600 185.400 ;
        RECT 41.200 181.600 42.000 186.200 ;
        RECT 44.400 181.600 45.200 184.200 ;
        RECT 47.600 181.600 48.400 188.200 ;
        RECT 55.600 181.600 56.400 184.200 ;
        RECT 57.200 181.600 58.000 186.200 ;
        RECT 66.800 181.600 67.600 184.200 ;
        RECT 73.200 181.600 74.000 186.200 ;
        RECT 84.400 181.600 85.200 184.200 ;
        RECT 87.600 181.600 88.400 184.200 ;
        RECT 97.200 181.600 98.000 186.200 ;
        RECT 103.600 181.600 104.400 186.200 ;
        RECT 110.000 181.600 110.800 186.200 ;
        RECT 119.600 181.600 120.400 184.200 ;
        RECT 122.800 181.600 123.600 184.200 ;
        RECT 134.000 181.600 134.800 186.200 ;
        RECT 140.400 181.600 141.200 184.200 ;
        RECT 143.600 181.600 144.400 186.200 ;
        RECT 148.400 181.600 149.400 185.600 ;
        RECT 154.600 182.200 155.600 185.600 ;
        RECT 154.600 181.600 155.400 182.200 ;
        RECT 164.400 181.600 165.200 186.200 ;
        RECT 167.600 181.600 168.400 184.200 ;
        RECT 170.800 181.600 171.600 184.200 ;
        RECT 174.000 181.600 174.800 184.200 ;
        RECT 178.200 181.600 179.000 186.000 ;
        RECT 185.200 181.600 186.000 186.200 ;
        RECT 194.800 181.600 195.600 184.200 ;
        RECT 198.000 181.600 198.800 184.200 ;
        RECT 209.200 181.600 210.000 186.200 ;
        RECT 215.600 181.600 216.400 184.200 ;
        RECT 0.400 180.400 220.400 181.600 ;
        RECT 1.200 177.800 2.000 180.400 ;
        RECT 7.600 175.800 8.400 180.400 ;
        RECT 18.800 177.800 19.600 180.400 ;
        RECT 22.000 177.800 22.800 180.400 ;
        RECT 31.600 175.800 32.400 180.400 ;
        RECT 38.000 175.800 38.800 180.400 ;
        RECT 46.000 173.800 46.800 180.400 ;
        RECT 49.200 177.800 50.000 180.400 ;
        RECT 52.400 177.800 53.200 180.400 ;
        RECT 57.200 176.600 58.000 180.400 ;
        RECT 66.800 177.800 67.600 180.400 ;
        RECT 70.000 178.200 70.800 180.400 ;
        RECT 79.800 179.800 80.600 180.400 ;
        RECT 79.600 176.400 80.600 179.800 ;
        RECT 85.800 176.400 86.800 180.400 ;
        RECT 89.200 175.800 90.000 180.400 ;
        RECT 92.400 175.800 93.200 180.400 ;
        RECT 95.600 175.800 96.400 180.400 ;
        RECT 98.800 175.800 99.600 180.400 ;
        RECT 102.000 175.800 102.800 180.400 ;
        RECT 106.800 175.800 107.600 180.400 ;
        RECT 116.400 177.800 117.200 180.400 ;
        RECT 119.600 177.800 120.400 180.400 ;
        RECT 130.800 175.800 131.600 180.400 ;
        RECT 137.200 177.800 138.000 180.400 ;
        RECT 140.400 175.800 141.200 180.400 ;
        RECT 145.400 179.800 146.200 180.400 ;
        RECT 145.200 176.400 146.200 179.800 ;
        RECT 151.400 176.400 152.400 180.400 ;
        RECT 159.600 177.800 160.400 180.400 ;
        RECT 166.000 175.800 166.800 180.400 ;
        RECT 169.200 176.400 170.200 180.400 ;
        RECT 175.400 179.800 176.200 180.400 ;
        RECT 175.400 176.400 176.400 179.800 ;
        RECT 178.800 175.800 179.600 180.400 ;
        RECT 183.600 177.800 184.400 180.400 ;
        RECT 186.800 177.800 187.600 180.400 ;
        RECT 190.000 177.800 190.800 180.400 ;
        RECT 193.400 179.800 194.200 180.400 ;
        RECT 193.200 176.400 194.200 179.800 ;
        RECT 199.400 176.400 200.400 180.400 ;
        RECT 205.000 176.000 205.800 180.400 ;
        RECT 210.800 175.800 211.600 180.400 ;
        RECT 215.600 175.800 216.400 180.400 ;
        RECT 2.800 141.600 3.600 146.200 ;
        RECT 7.600 141.600 8.400 146.200 ;
        RECT 10.800 141.600 11.600 144.200 ;
        RECT 14.000 141.600 14.800 144.200 ;
        RECT 17.200 141.600 18.000 148.200 ;
        RECT 23.600 141.600 24.400 146.200 ;
        RECT 31.600 141.600 32.400 145.400 ;
        RECT 38.000 141.600 38.800 146.200 ;
        RECT 42.800 141.600 43.600 146.200 ;
        RECT 52.400 141.600 53.200 144.200 ;
        RECT 55.600 141.600 56.400 144.200 ;
        RECT 66.800 141.600 67.600 146.200 ;
        RECT 73.200 141.600 74.000 144.200 ;
        RECT 82.800 141.600 83.600 146.200 ;
        RECT 92.400 141.600 93.200 144.200 ;
        RECT 95.600 141.600 96.400 144.200 ;
        RECT 106.800 141.600 107.600 146.200 ;
        RECT 113.200 141.600 114.000 144.200 ;
        RECT 114.800 141.600 115.600 146.200 ;
        RECT 118.000 141.600 118.800 146.200 ;
        RECT 121.200 141.600 122.000 146.200 ;
        RECT 124.400 141.600 125.200 146.200 ;
        RECT 127.600 141.600 128.400 146.200 ;
        RECT 132.400 141.600 133.200 146.200 ;
        RECT 142.000 141.600 142.800 144.200 ;
        RECT 145.200 141.600 146.000 144.200 ;
        RECT 156.400 141.600 157.200 146.200 ;
        RECT 162.800 141.600 163.600 144.200 ;
        RECT 172.400 141.600 173.200 146.200 ;
        RECT 177.200 141.600 178.000 146.200 ;
        RECT 186.800 141.600 187.600 144.200 ;
        RECT 190.000 141.600 190.800 144.200 ;
        RECT 201.200 141.600 202.000 146.200 ;
        RECT 207.600 141.600 208.400 144.200 ;
        RECT 210.800 141.600 211.600 146.200 ;
        RECT 215.600 141.600 216.400 146.200 ;
        RECT 0.400 140.400 220.400 141.600 ;
        RECT 1.200 137.800 2.000 140.400 ;
        RECT 7.600 135.800 8.400 140.400 ;
        RECT 18.800 137.800 19.600 140.400 ;
        RECT 22.000 137.800 22.800 140.400 ;
        RECT 31.600 135.800 32.400 140.400 ;
        RECT 38.000 137.800 38.800 140.400 ;
        RECT 41.200 138.200 42.000 140.400 ;
        RECT 51.000 139.800 51.800 140.400 ;
        RECT 50.800 136.400 51.800 139.800 ;
        RECT 57.000 136.400 58.000 140.400 ;
        RECT 65.200 137.800 66.000 140.400 ;
        RECT 71.600 135.800 72.400 140.400 ;
        RECT 82.800 137.800 83.600 140.400 ;
        RECT 86.000 137.800 86.800 140.400 ;
        RECT 95.600 135.800 96.400 140.400 ;
        RECT 102.000 136.400 103.000 140.400 ;
        RECT 108.200 139.800 109.000 140.400 ;
        RECT 108.200 136.400 109.200 139.800 ;
        RECT 111.600 135.800 112.400 140.400 ;
        RECT 114.800 135.800 115.600 140.400 ;
        RECT 121.200 135.800 122.000 140.400 ;
        RECT 124.400 136.400 125.400 140.400 ;
        RECT 130.600 139.800 131.400 140.400 ;
        RECT 130.600 136.400 131.600 139.800 ;
        RECT 137.200 135.800 138.000 140.400 ;
        RECT 146.800 137.800 147.600 140.400 ;
        RECT 150.000 137.800 150.800 140.400 ;
        RECT 161.200 135.800 162.000 140.400 ;
        RECT 167.600 137.800 168.400 140.400 ;
        RECT 175.600 136.400 176.600 140.400 ;
        RECT 181.800 139.800 182.600 140.400 ;
        RECT 181.800 136.400 182.800 139.800 ;
        RECT 185.200 137.800 186.000 140.400 ;
        RECT 188.400 137.800 189.200 140.400 ;
        RECT 194.800 133.800 195.600 140.400 ;
        RECT 198.200 139.800 199.000 140.400 ;
        RECT 198.000 136.400 199.000 139.800 ;
        RECT 204.200 136.400 205.200 140.400 ;
        RECT 210.800 135.800 211.600 140.400 ;
        RECT 214.000 135.800 214.800 140.400 ;
        RECT 2.800 101.600 3.600 106.200 ;
        RECT 7.600 101.600 8.400 106.200 ;
        RECT 12.400 101.600 13.400 105.600 ;
        RECT 18.600 102.200 19.600 105.600 ;
        RECT 18.600 101.600 19.400 102.200 ;
        RECT 22.000 101.600 22.800 104.200 ;
        RECT 25.200 101.600 26.000 104.200 ;
        RECT 28.400 101.600 29.200 108.200 ;
        RECT 36.400 101.600 37.200 106.200 ;
        RECT 39.600 101.600 40.400 106.200 ;
        RECT 42.800 101.600 43.600 106.200 ;
        RECT 46.000 101.600 46.800 106.200 ;
        RECT 49.200 101.600 50.000 106.200 ;
        RECT 52.400 101.600 53.200 106.200 ;
        RECT 58.800 101.600 59.600 104.200 ;
        RECT 65.200 101.600 66.000 106.200 ;
        RECT 76.400 101.600 77.200 104.200 ;
        RECT 79.600 101.600 80.400 104.200 ;
        RECT 89.200 101.600 90.000 106.200 ;
        RECT 94.000 101.600 94.800 104.200 ;
        RECT 100.400 101.600 101.200 106.200 ;
        RECT 111.600 101.600 112.400 104.200 ;
        RECT 114.800 101.600 115.600 104.200 ;
        RECT 124.400 101.600 125.200 106.200 ;
        RECT 130.800 101.600 131.600 106.200 ;
        RECT 134.000 101.600 134.800 106.200 ;
        RECT 138.800 101.600 139.600 106.200 ;
        RECT 148.400 101.600 149.200 104.200 ;
        RECT 151.600 101.600 152.400 104.200 ;
        RECT 162.800 101.600 163.600 106.200 ;
        RECT 169.200 101.600 170.000 104.200 ;
        RECT 178.800 101.600 179.600 106.200 ;
        RECT 188.400 101.600 189.200 104.200 ;
        RECT 191.600 101.600 192.400 104.200 ;
        RECT 202.800 101.600 203.600 106.200 ;
        RECT 209.200 101.600 210.000 104.200 ;
        RECT 212.400 101.600 213.200 106.200 ;
        RECT 0.400 100.400 220.400 101.600 ;
        RECT 1.200 97.800 2.000 100.400 ;
        RECT 7.600 95.800 8.400 100.400 ;
        RECT 18.800 97.800 19.600 100.400 ;
        RECT 22.000 97.800 22.800 100.400 ;
        RECT 31.600 95.800 32.400 100.400 ;
        RECT 36.400 97.800 37.200 100.400 ;
        RECT 42.800 95.800 43.600 100.400 ;
        RECT 54.000 97.800 54.800 100.400 ;
        RECT 57.200 97.800 58.000 100.400 ;
        RECT 66.800 95.800 67.600 100.400 ;
        RECT 76.400 95.800 77.200 100.400 ;
        RECT 79.600 95.800 80.400 100.400 ;
        RECT 84.600 99.800 85.400 100.400 ;
        RECT 84.400 96.400 85.400 99.800 ;
        RECT 90.600 96.400 91.600 100.400 ;
        RECT 95.600 96.600 96.400 100.400 ;
        RECT 100.400 97.800 101.200 100.400 ;
        RECT 103.600 95.800 104.400 100.400 ;
        RECT 108.400 97.800 109.200 100.400 ;
        RECT 114.800 95.800 115.600 100.400 ;
        RECT 126.000 97.800 126.800 100.400 ;
        RECT 129.200 97.800 130.000 100.400 ;
        RECT 138.800 95.800 139.600 100.400 ;
        RECT 151.600 95.800 152.400 100.400 ;
        RECT 161.200 97.800 162.000 100.400 ;
        RECT 164.400 97.800 165.200 100.400 ;
        RECT 175.600 95.800 176.400 100.400 ;
        RECT 182.000 97.800 182.800 100.400 ;
        RECT 185.200 96.400 186.200 100.400 ;
        RECT 191.400 99.800 192.200 100.400 ;
        RECT 191.400 96.400 192.400 99.800 ;
        RECT 198.000 95.800 198.800 100.400 ;
        RECT 202.800 95.800 203.600 100.400 ;
        RECT 206.200 99.800 207.000 100.400 ;
        RECT 206.000 96.400 207.000 99.800 ;
        RECT 212.200 96.400 213.200 100.400 ;
        RECT 217.200 95.800 218.000 100.400 ;
        RECT 2.800 61.600 3.600 66.200 ;
        RECT 7.600 61.600 8.400 66.200 ;
        RECT 12.400 61.600 13.200 64.200 ;
        RECT 15.600 61.600 16.400 63.800 ;
        RECT 25.200 61.600 26.000 65.400 ;
        RECT 30.000 61.600 30.800 66.200 ;
        RECT 36.400 62.200 37.400 65.600 ;
        RECT 36.600 61.600 37.400 62.200 ;
        RECT 42.600 61.600 43.600 65.600 ;
        RECT 50.800 61.600 51.600 64.200 ;
        RECT 57.200 61.600 58.000 66.200 ;
        RECT 68.400 61.600 69.200 64.200 ;
        RECT 71.600 61.600 72.400 64.200 ;
        RECT 81.200 61.600 82.000 66.200 ;
        RECT 87.600 61.600 88.400 64.200 ;
        RECT 89.200 61.600 90.000 66.200 ;
        RECT 92.400 61.600 93.200 66.200 ;
        RECT 95.600 61.600 96.400 66.200 ;
        RECT 98.800 61.600 99.600 66.200 ;
        RECT 102.000 61.600 102.800 66.200 ;
        RECT 103.600 61.600 104.400 68.200 ;
        RECT 110.000 61.600 110.800 64.200 ;
        RECT 113.200 61.600 114.000 66.200 ;
        RECT 116.400 61.600 117.200 66.200 ;
        RECT 119.600 61.600 120.400 66.200 ;
        RECT 122.800 61.600 123.600 66.200 ;
        RECT 126.000 61.600 126.800 66.200 ;
        RECT 129.200 61.600 130.000 66.200 ;
        RECT 132.400 61.600 133.200 66.200 ;
        RECT 134.000 61.600 134.800 66.200 ;
        RECT 137.200 61.600 138.000 66.200 ;
        RECT 140.400 61.600 141.200 66.200 ;
        RECT 143.600 61.600 144.400 66.200 ;
        RECT 146.800 61.600 147.600 66.200 ;
        RECT 148.400 61.600 149.200 64.200 ;
        RECT 151.600 61.600 152.400 64.200 ;
        RECT 158.000 61.600 158.800 64.200 ;
        RECT 161.200 61.600 162.000 64.200 ;
        RECT 165.400 61.600 166.200 66.000 ;
        RECT 170.800 61.600 171.600 66.200 ;
        RECT 175.600 62.200 176.600 65.600 ;
        RECT 175.800 61.600 176.600 62.200 ;
        RECT 181.800 61.600 182.800 65.600 ;
        RECT 187.800 61.600 188.600 66.000 ;
        RECT 193.800 61.600 194.600 66.000 ;
        RECT 198.000 61.600 198.800 64.200 ;
        RECT 201.200 61.600 202.000 64.200 ;
        RECT 202.800 61.600 203.600 64.200 ;
        RECT 206.000 61.600 206.800 64.200 ;
        RECT 209.200 61.600 210.000 64.200 ;
        RECT 212.400 61.600 213.200 66.200 ;
        RECT 0.400 60.400 220.400 61.600 ;
        RECT 1.200 57.800 2.000 60.400 ;
        RECT 7.600 55.800 8.400 60.400 ;
        RECT 18.800 57.800 19.600 60.400 ;
        RECT 22.000 57.800 22.800 60.400 ;
        RECT 31.600 55.800 32.400 60.400 ;
        RECT 39.600 55.800 40.400 60.400 ;
        RECT 41.200 57.800 42.000 60.400 ;
        RECT 44.400 53.800 45.200 60.400 ;
        RECT 54.000 56.600 54.800 60.400 ;
        RECT 63.600 57.800 64.400 60.400 ;
        RECT 66.800 58.200 67.600 60.400 ;
        RECT 74.800 57.800 75.600 60.400 ;
        RECT 78.000 53.800 78.800 60.400 ;
        RECT 90.800 58.200 91.600 60.400 ;
        RECT 94.000 57.800 94.800 60.400 ;
        RECT 98.800 56.600 99.600 60.400 ;
        RECT 103.600 55.800 104.400 60.400 ;
        RECT 108.400 57.800 109.200 60.400 ;
        RECT 111.600 57.800 112.400 60.400 ;
        RECT 115.800 56.000 116.600 60.400 ;
        RECT 119.600 57.800 120.400 60.400 ;
        RECT 122.800 57.800 123.600 60.400 ;
        RECT 127.600 55.800 128.400 60.400 ;
        RECT 137.200 57.800 138.000 60.400 ;
        RECT 140.400 57.800 141.200 60.400 ;
        RECT 151.600 55.800 152.400 60.400 ;
        RECT 158.000 57.800 158.800 60.400 ;
        RECT 167.600 55.800 168.400 60.400 ;
        RECT 177.200 57.800 178.000 60.400 ;
        RECT 180.400 57.800 181.200 60.400 ;
        RECT 191.600 55.800 192.400 60.400 ;
        RECT 198.000 57.800 198.800 60.400 ;
        RECT 199.600 57.800 200.400 60.400 ;
        RECT 202.800 57.800 203.600 60.400 ;
        RECT 207.600 55.800 208.400 60.400 ;
        RECT 209.800 55.800 210.600 60.400 ;
        RECT 214.000 57.800 214.800 60.400 ;
        RECT 217.200 55.800 218.000 60.400 ;
        RECT 2.800 21.600 3.600 26.200 ;
        RECT 6.000 21.600 6.800 24.200 ;
        RECT 14.000 21.600 14.800 28.200 ;
        RECT 17.200 21.600 18.000 24.200 ;
        RECT 20.400 21.600 21.400 25.600 ;
        RECT 26.600 22.200 27.600 25.600 ;
        RECT 26.600 21.600 27.400 22.200 ;
        RECT 31.600 21.600 32.400 25.400 ;
        RECT 38.000 21.600 38.800 24.200 ;
        RECT 41.200 21.600 42.000 23.800 ;
        RECT 50.800 21.600 51.600 24.200 ;
        RECT 52.400 21.600 53.200 26.200 ;
        RECT 63.600 22.200 64.600 25.600 ;
        RECT 63.800 21.600 64.600 22.200 ;
        RECT 69.800 21.600 70.800 25.600 ;
        RECT 76.400 21.600 77.200 26.200 ;
        RECT 86.000 21.600 86.800 24.200 ;
        RECT 89.200 21.600 90.000 24.200 ;
        RECT 100.400 21.600 101.200 26.200 ;
        RECT 106.800 21.600 107.600 24.200 ;
        RECT 108.400 21.600 109.200 24.200 ;
        RECT 114.800 21.600 115.600 26.200 ;
        RECT 126.000 21.600 126.800 24.200 ;
        RECT 129.200 21.600 130.000 24.200 ;
        RECT 138.800 21.600 139.600 26.200 ;
        RECT 143.600 21.600 144.400 26.200 ;
        RECT 148.400 21.600 149.200 24.200 ;
        RECT 151.600 21.600 152.400 24.200 ;
        RECT 158.000 21.600 158.800 24.200 ;
        RECT 161.200 21.600 162.000 24.200 ;
        RECT 164.400 21.600 165.200 24.200 ;
        RECT 169.200 21.600 170.000 26.200 ;
        RECT 178.800 21.600 179.600 24.200 ;
        RECT 182.000 21.600 182.800 24.200 ;
        RECT 193.200 21.600 194.000 26.200 ;
        RECT 199.600 21.600 200.400 24.200 ;
        RECT 202.800 22.200 203.800 25.600 ;
        RECT 203.000 21.600 203.800 22.200 ;
        RECT 209.000 21.600 210.000 25.600 ;
        RECT 214.000 21.600 214.800 26.200 ;
        RECT 0.400 20.400 220.400 21.600 ;
        RECT 2.800 15.800 3.600 20.400 ;
        RECT 6.000 17.800 6.800 20.400 ;
        RECT 12.400 15.800 13.200 20.400 ;
        RECT 23.600 17.800 24.400 20.400 ;
        RECT 26.800 17.800 27.600 20.400 ;
        RECT 36.400 15.800 37.200 20.400 ;
        RECT 42.800 15.800 43.600 20.400 ;
        RECT 50.800 17.800 51.600 20.400 ;
        RECT 57.200 15.800 58.000 20.400 ;
        RECT 68.400 17.800 69.200 20.400 ;
        RECT 71.600 17.800 72.400 20.400 ;
        RECT 81.200 15.800 82.000 20.400 ;
        RECT 87.600 15.800 88.400 20.400 ;
        RECT 92.400 15.800 93.200 20.400 ;
        RECT 97.200 15.800 98.000 20.400 ;
        RECT 102.000 15.800 102.800 20.400 ;
        RECT 105.200 17.800 106.000 20.400 ;
        RECT 111.600 15.800 112.400 20.400 ;
        RECT 122.800 17.800 123.600 20.400 ;
        RECT 126.000 17.800 126.800 20.400 ;
        RECT 135.600 15.800 136.400 20.400 ;
        RECT 145.200 17.800 146.000 20.400 ;
        RECT 151.600 15.800 152.400 20.400 ;
        RECT 162.800 17.800 163.600 20.400 ;
        RECT 166.000 17.800 166.800 20.400 ;
        RECT 175.600 15.800 176.400 20.400 ;
        RECT 183.600 15.800 184.400 20.400 ;
        RECT 193.200 17.800 194.000 20.400 ;
        RECT 196.400 17.800 197.200 20.400 ;
        RECT 207.600 15.800 208.400 20.400 ;
        RECT 214.000 17.800 214.800 20.400 ;
      LAYER via1 ;
        RECT 156.600 180.600 157.400 181.400 ;
        RECT 158.000 180.600 158.800 181.400 ;
        RECT 159.400 180.600 160.200 181.400 ;
        RECT 156.600 140.600 157.400 141.400 ;
        RECT 158.000 140.600 158.800 141.400 ;
        RECT 159.400 140.600 160.200 141.400 ;
        RECT 156.600 100.600 157.400 101.400 ;
        RECT 158.000 100.600 158.800 101.400 ;
        RECT 159.400 100.600 160.200 101.400 ;
        RECT 156.600 60.600 157.400 61.400 ;
        RECT 158.000 60.600 158.800 61.400 ;
        RECT 159.400 60.600 160.200 61.400 ;
        RECT 156.600 20.600 157.400 21.400 ;
        RECT 158.000 20.600 158.800 21.400 ;
        RECT 159.400 20.600 160.200 21.400 ;
      LAYER metal2 ;
        RECT 156.000 180.600 160.800 181.400 ;
        RECT 156.000 140.600 160.800 141.400 ;
        RECT 156.000 100.600 160.800 101.400 ;
        RECT 156.000 60.600 160.800 61.400 ;
        RECT 156.000 20.600 160.800 21.400 ;
      LAYER via2 ;
        RECT 156.600 180.600 157.400 181.400 ;
        RECT 158.000 180.600 158.800 181.400 ;
        RECT 159.400 180.600 160.200 181.400 ;
        RECT 156.600 140.600 157.400 141.400 ;
        RECT 158.000 140.600 158.800 141.400 ;
        RECT 159.400 140.600 160.200 141.400 ;
        RECT 156.600 100.600 157.400 101.400 ;
        RECT 158.000 100.600 158.800 101.400 ;
        RECT 159.400 100.600 160.200 101.400 ;
        RECT 156.600 60.600 157.400 61.400 ;
        RECT 158.000 60.600 158.800 61.400 ;
        RECT 159.400 60.600 160.200 61.400 ;
        RECT 156.600 20.600 157.400 21.400 ;
        RECT 158.000 20.600 158.800 21.400 ;
        RECT 159.400 20.600 160.200 21.400 ;
      LAYER metal3 ;
        RECT 156.000 180.400 160.800 181.600 ;
        RECT 156.000 140.400 160.800 141.600 ;
        RECT 156.000 100.400 160.800 101.600 ;
        RECT 156.000 60.400 160.800 61.600 ;
        RECT 156.000 20.400 160.800 21.600 ;
      LAYER via3 ;
        RECT 156.400 180.600 157.200 181.400 ;
        RECT 158.000 180.600 158.800 181.400 ;
        RECT 159.600 180.600 160.400 181.400 ;
        RECT 156.400 140.600 157.200 141.400 ;
        RECT 158.000 140.600 158.800 141.400 ;
        RECT 159.600 140.600 160.400 141.400 ;
        RECT 156.400 100.600 157.200 101.400 ;
        RECT 158.000 100.600 158.800 101.400 ;
        RECT 159.600 100.600 160.400 101.400 ;
        RECT 156.400 60.600 157.200 61.400 ;
        RECT 158.000 60.600 158.800 61.400 ;
        RECT 159.600 60.600 160.400 61.400 ;
        RECT 156.400 20.600 157.200 21.400 ;
        RECT 158.000 20.600 158.800 21.400 ;
        RECT 159.600 20.600 160.400 21.400 ;
      LAYER metal4 ;
        RECT 156.000 -4.000 160.800 204.000 ;
    END
  END gnd
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 102.000 173.800 102.800 174.400 ;
        RECT 101.000 173.000 102.800 173.800 ;
        RECT 114.800 148.200 116.600 149.000 ;
        RECT 114.800 147.600 115.600 148.200 ;
        RECT 101.000 68.200 102.800 69.000 ;
        RECT 125.000 68.200 126.800 69.000 ;
        RECT 102.000 67.600 102.800 68.200 ;
        RECT 126.000 67.600 126.800 68.200 ;
        RECT 132.400 68.300 133.200 68.400 ;
        RECT 134.000 68.300 135.800 69.000 ;
        RECT 132.400 68.200 135.800 68.300 ;
        RECT 132.400 67.700 134.800 68.200 ;
        RECT 132.400 67.600 133.200 67.700 ;
        RECT 134.000 67.600 134.800 67.700 ;
      LAYER via1 ;
        RECT 102.000 173.600 102.800 174.400 ;
      LAYER metal2 ;
        RECT 102.100 203.700 104.300 204.300 ;
        RECT 102.000 174.300 102.800 174.400 ;
        RECT 103.700 174.300 104.300 203.700 ;
        RECT 102.000 173.700 104.300 174.300 ;
        RECT 102.000 173.600 102.800 173.700 ;
        RECT 102.100 164.400 102.700 173.600 ;
        RECT 102.000 163.600 102.800 164.400 ;
        RECT 114.800 163.600 115.600 164.400 ;
        RECT 114.900 148.400 115.500 163.600 ;
        RECT 114.800 147.600 115.600 148.400 ;
        RECT 114.900 142.400 115.500 147.600 ;
        RECT 114.800 141.600 115.600 142.400 ;
        RECT 102.000 67.600 102.800 68.400 ;
        RECT 126.000 67.600 126.800 68.400 ;
        RECT 132.400 67.600 133.200 68.400 ;
      LAYER metal3 ;
        RECT 102.000 164.300 102.800 164.400 ;
        RECT 114.800 164.300 115.600 164.400 ;
        RECT 102.000 163.700 115.600 164.300 ;
        RECT 102.000 163.600 102.800 163.700 ;
        RECT 114.800 163.600 115.600 163.700 ;
        RECT 113.200 142.300 114.000 142.400 ;
        RECT 114.800 142.300 115.600 142.400 ;
        RECT 113.200 141.700 115.600 142.300 ;
        RECT 113.200 141.600 114.000 141.700 ;
        RECT 114.800 141.600 115.600 141.700 ;
        RECT 102.000 68.300 102.800 68.400 ;
        RECT 113.200 68.300 114.000 68.400 ;
        RECT 126.000 68.300 126.800 68.400 ;
        RECT 132.400 68.300 133.200 68.400 ;
        RECT 102.000 67.700 133.200 68.300 ;
        RECT 102.000 67.600 102.800 67.700 ;
        RECT 113.200 67.600 114.000 67.700 ;
        RECT 126.000 67.600 126.800 67.700 ;
        RECT 132.400 67.600 133.200 67.700 ;
      LAYER metal4 ;
        RECT 113.000 67.400 114.200 142.600 ;
    END
  END clk
  PIN rst
    PORT
      LAYER metal1 ;
        RECT 46.000 106.800 46.800 108.400 ;
      LAYER via1 ;
        RECT 46.000 107.600 46.800 108.400 ;
      LAYER metal2 ;
        RECT 46.000 107.600 46.800 108.400 ;
      LAYER metal3 ;
        RECT 26.800 126.300 27.600 126.400 ;
        RECT -1.900 125.700 27.600 126.300 ;
        RECT 26.800 125.600 27.600 125.700 ;
        RECT 26.800 108.300 27.600 108.400 ;
        RECT 46.000 108.300 46.800 108.400 ;
        RECT 26.800 107.700 46.800 108.300 ;
        RECT 26.800 107.600 27.600 107.700 ;
        RECT 46.000 107.600 46.800 107.700 ;
      LAYER metal4 ;
        RECT 26.600 107.400 27.800 126.600 ;
    END
  END rst
  PIN theta[0]
    PORT
      LAYER metal3 ;
        RECT -1.900 51.700 -1.300 52.300 ;
    END
  END theta[0]
  PIN theta[1]
    PORT
      LAYER metal3 ;
        RECT -1.900 29.700 -1.300 30.300 ;
    END
  END theta[1]
  PIN theta[2]
    PORT
      LAYER metal3 ;
        RECT 222.100 11.700 222.700 12.300 ;
    END
  END theta[2]
  PIN theta[3]
    PORT
      LAYER metal3 ;
        RECT -1.900 141.700 -1.300 142.300 ;
    END
  END theta[3]
  PIN theta[4]
    PORT
      LAYER metal3 ;
        RECT -1.900 135.700 -1.300 136.300 ;
    END
  END theta[4]
  PIN theta[5]
    PORT
      LAYER metal3 ;
        RECT 222.100 117.700 222.700 118.300 ;
    END
  END theta[5]
  PIN theta[6]
    PORT
      LAYER metal2 ;
        RECT 172.500 203.700 173.100 204.300 ;
    END
  END theta[6]
  PIN theta[7]
    PORT
      LAYER metal2 ;
        RECT 201.300 203.700 201.900 204.300 ;
    END
  END theta[7]
  PIN theta[8]
    PORT
      LAYER metal2 ;
        RECT 47.700 -2.300 48.300 -1.700 ;
    END
  END theta[8]
  PIN theta[9]
    PORT
      LAYER metal3 ;
        RECT -1.900 15.700 -1.300 16.300 ;
    END
  END theta[9]
  PIN theta[10]
    PORT
      LAYER metal3 ;
        RECT -1.900 109.700 -1.300 110.300 ;
    END
  END theta[10]
  PIN theta[11]
    PORT
      LAYER metal2 ;
        RECT 145.300 -2.300 145.900 -1.700 ;
    END
  END theta[11]
  PIN theta[12]
    PORT
      LAYER metal3 ;
        RECT -1.900 147.700 -1.300 148.300 ;
    END
  END theta[12]
  PIN theta[13]
    PORT
      LAYER metal2 ;
        RECT 167.700 203.700 168.300 204.300 ;
    END
  END theta[13]
  PIN theta[14]
    PORT
      LAYER metal3 ;
        RECT 222.100 179.700 222.700 180.300 ;
    END
  END theta[14]
  PIN theta[15]
    PORT
      LAYER metal3 ;
        RECT 222.100 95.700 222.700 96.300 ;
    END
  END theta[15]
  PIN sine[0]
    PORT
      LAYER metal1 ;
        RECT 103.600 12.400 104.400 19.800 ;
        RECT 103.800 10.200 104.400 12.400 ;
        RECT 103.600 2.200 104.400 10.200 ;
      LAYER via1 ;
        RECT 103.600 3.600 104.400 4.400 ;
      LAYER metal2 ;
        RECT 103.600 3.600 104.400 4.400 ;
        RECT 103.700 -1.700 104.300 3.600 ;
        RECT 102.100 -2.300 104.300 -1.700 ;
    END
  END sine[0]
  PIN sine[1]
    PORT
      LAYER metal1 ;
        RECT 138.800 172.400 139.600 179.800 ;
        RECT 138.800 170.200 139.400 172.400 ;
        RECT 138.800 162.200 139.600 170.200 ;
      LAYER via1 ;
        RECT 138.800 163.600 139.600 164.400 ;
      LAYER metal2 ;
        RECT 138.800 163.600 139.600 164.400 ;
        RECT 138.900 160.400 139.500 163.600 ;
        RECT 138.800 159.600 139.600 160.400 ;
        RECT 140.400 1.600 141.200 2.400 ;
        RECT 140.500 -2.300 141.100 1.600 ;
      LAYER metal3 ;
        RECT 138.800 159.600 139.600 160.400 ;
        RECT 138.800 2.300 139.600 2.400 ;
        RECT 140.400 2.300 141.200 2.400 ;
        RECT 138.800 1.700 141.200 2.300 ;
        RECT 138.800 1.600 139.600 1.700 ;
        RECT 140.400 1.600 141.200 1.700 ;
      LAYER metal4 ;
        RECT 138.600 1.400 139.800 160.600 ;
    END
  END sine[1]
  PIN sine[2]
    PORT
      LAYER metal1 ;
        RECT 172.400 71.800 173.200 79.800 ;
        RECT 172.600 69.600 173.200 71.800 ;
        RECT 172.400 62.200 173.200 69.600 ;
      LAYER via1 ;
        RECT 172.400 73.600 173.200 74.400 ;
      LAYER metal2 ;
        RECT 172.400 73.600 173.200 74.400 ;
      LAYER metal3 ;
        RECT 172.400 74.300 173.200 74.400 ;
        RECT 172.400 73.700 222.700 74.300 ;
        RECT 172.400 73.600 173.200 73.700 ;
    END
  END sine[2]
  PIN sine[3]
    PORT
      LAYER metal1 ;
        RECT 214.000 71.800 214.800 79.800 ;
        RECT 214.200 69.600 214.800 71.800 ;
        RECT 214.000 68.300 214.800 69.600 ;
        RECT 218.800 68.300 219.600 68.400 ;
        RECT 214.000 67.700 219.600 68.300 ;
        RECT 214.000 62.200 214.800 67.700 ;
        RECT 218.800 67.600 219.600 67.700 ;
      LAYER metal2 ;
        RECT 218.800 69.600 219.600 70.400 ;
        RECT 218.900 68.400 219.500 69.600 ;
        RECT 218.800 67.600 219.600 68.400 ;
      LAYER metal3 ;
        RECT 218.800 70.300 219.600 70.400 ;
        RECT 218.800 69.700 222.700 70.300 ;
        RECT 218.800 69.600 219.600 69.700 ;
    END
  END sine[3]
  PIN sine[4]
    PORT
      LAYER metal1 ;
        RECT 215.600 31.800 216.400 39.800 ;
        RECT 215.800 29.600 216.400 31.800 ;
        RECT 215.600 28.300 216.400 29.600 ;
        RECT 218.800 28.300 219.600 28.400 ;
        RECT 215.600 27.700 219.600 28.300 ;
        RECT 215.600 22.200 216.400 27.700 ;
        RECT 218.800 27.600 219.600 27.700 ;
      LAYER metal2 ;
        RECT 218.800 29.600 219.600 30.400 ;
        RECT 218.900 28.400 219.500 29.600 ;
        RECT 218.800 27.600 219.600 28.400 ;
      LAYER metal3 ;
        RECT 218.800 30.300 219.600 30.400 ;
        RECT 218.800 29.700 222.700 30.300 ;
        RECT 218.800 29.600 219.600 29.700 ;
    END
  END sine[4]
  PIN sine[5]
    PORT
      LAYER metal1 ;
        RECT 218.800 52.400 219.600 59.800 ;
        RECT 219.000 50.200 219.600 52.400 ;
        RECT 218.800 42.200 219.600 50.200 ;
      LAYER via1 ;
        RECT 218.800 47.600 219.600 48.400 ;
      LAYER metal2 ;
        RECT 218.800 49.600 219.600 50.400 ;
        RECT 218.900 48.400 219.500 49.600 ;
        RECT 218.800 47.600 219.600 48.400 ;
      LAYER metal3 ;
        RECT 218.800 50.300 219.600 50.400 ;
        RECT 218.800 49.700 222.700 50.300 ;
        RECT 218.800 49.600 219.600 49.700 ;
    END
  END sine[5]
  PIN sine[6]
    PORT
      LAYER metal1 ;
        RECT 214.000 111.800 214.800 119.800 ;
        RECT 214.200 109.600 214.800 111.800 ;
        RECT 214.000 108.300 214.800 109.600 ;
        RECT 218.800 108.300 219.600 108.400 ;
        RECT 214.000 107.700 219.600 108.300 ;
        RECT 214.000 102.200 214.800 107.700 ;
        RECT 218.800 107.600 219.600 107.700 ;
      LAYER metal2 ;
        RECT 218.800 109.600 219.600 110.400 ;
        RECT 218.900 108.400 219.500 109.600 ;
        RECT 218.800 107.600 219.600 108.400 ;
      LAYER metal3 ;
        RECT 218.800 110.300 219.600 110.400 ;
        RECT 218.800 109.700 222.700 110.300 ;
        RECT 218.800 109.600 219.600 109.700 ;
    END
  END sine[6]
  PIN sine[7]
    PORT
      LAYER metal1 ;
        RECT 218.800 92.400 219.600 99.800 ;
        RECT 219.000 90.200 219.600 92.400 ;
        RECT 218.800 82.200 219.600 90.200 ;
      LAYER via1 ;
        RECT 218.800 87.600 219.600 88.400 ;
      LAYER metal2 ;
        RECT 218.800 89.600 219.600 90.400 ;
        RECT 218.900 88.400 219.500 89.600 ;
        RECT 218.800 87.600 219.600 88.400 ;
      LAYER metal3 ;
        RECT 218.800 90.300 219.600 90.400 ;
        RECT 218.800 89.700 222.700 90.300 ;
        RECT 218.800 89.600 219.600 89.700 ;
    END
  END sine[7]
  PIN sine[8]
    PORT
      LAYER metal1 ;
        RECT 166.000 191.800 166.800 199.800 ;
        RECT 166.200 189.600 166.800 191.800 ;
        RECT 166.000 182.200 166.800 189.600 ;
      LAYER via1 ;
        RECT 166.000 197.600 166.800 198.400 ;
      LAYER metal2 ;
        RECT 164.500 203.700 166.700 204.300 ;
        RECT 166.100 198.400 166.700 203.700 ;
        RECT 166.000 197.600 166.800 198.400 ;
    END
  END sine[8]
  PIN sine[9]
    PORT
      LAYER metal1 ;
        RECT 142.000 191.800 142.800 199.800 ;
        RECT 142.000 189.600 142.600 191.800 ;
        RECT 142.000 182.200 142.800 189.600 ;
      LAYER via1 ;
        RECT 142.000 197.600 142.800 198.400 ;
      LAYER metal2 ;
        RECT 142.100 203.700 144.300 204.300 ;
        RECT 142.100 198.400 142.700 203.700 ;
        RECT 142.000 197.600 142.800 198.400 ;
    END
  END sine[9]
  PIN sine[10]
    PORT
      LAYER metal1 ;
        RECT 212.400 172.400 213.200 179.800 ;
        RECT 212.600 170.200 213.200 172.400 ;
        RECT 212.400 162.200 213.200 170.200 ;
      LAYER via1 ;
        RECT 212.400 173.600 213.200 174.400 ;
      LAYER metal2 ;
        RECT 212.400 173.600 213.200 174.400 ;
      LAYER metal3 ;
        RECT 212.400 174.300 213.200 174.400 ;
        RECT 212.400 173.700 222.700 174.300 ;
        RECT 212.400 173.600 213.200 173.700 ;
    END
  END sine[10]
  PIN sine[11]
    PORT
      LAYER metal1 ;
        RECT 217.200 172.400 218.000 179.800 ;
        RECT 217.400 170.200 218.000 172.400 ;
        RECT 217.200 168.300 218.000 170.200 ;
        RECT 218.800 168.300 219.600 168.400 ;
        RECT 217.200 167.700 219.600 168.300 ;
        RECT 217.200 162.200 218.000 167.700 ;
        RECT 218.800 167.600 219.600 167.700 ;
      LAYER metal2 ;
        RECT 218.800 169.600 219.600 170.400 ;
        RECT 218.900 168.400 219.500 169.600 ;
        RECT 218.800 167.600 219.600 168.400 ;
      LAYER metal3 ;
        RECT 218.800 170.300 219.600 170.400 ;
        RECT 218.800 169.700 222.700 170.300 ;
        RECT 218.800 169.600 219.600 169.700 ;
    END
  END sine[11]
  PIN sine[12]
    PORT
      LAYER metal1 ;
        RECT 215.600 132.400 216.400 139.800 ;
        RECT 215.800 130.200 216.400 132.400 ;
        RECT 215.600 128.300 216.400 130.200 ;
        RECT 218.800 128.300 219.600 128.400 ;
        RECT 215.600 127.700 219.600 128.300 ;
        RECT 215.600 122.200 216.400 127.700 ;
        RECT 218.800 127.600 219.600 127.700 ;
      LAYER metal2 ;
        RECT 218.800 129.600 219.600 130.400 ;
        RECT 218.900 128.400 219.500 129.600 ;
        RECT 218.800 127.600 219.600 128.400 ;
      LAYER metal3 ;
        RECT 218.800 130.300 219.600 130.400 ;
        RECT 218.800 129.700 222.700 130.300 ;
        RECT 218.800 129.600 219.600 129.700 ;
    END
  END sine[12]
  PIN sine[13]
    PORT
      LAYER metal1 ;
        RECT 212.400 151.800 213.200 159.800 ;
        RECT 212.600 149.600 213.200 151.800 ;
        RECT 212.400 142.200 213.200 149.600 ;
      LAYER via1 ;
        RECT 212.400 153.600 213.200 154.400 ;
      LAYER metal2 ;
        RECT 212.400 153.600 213.200 154.400 ;
      LAYER metal3 ;
        RECT 212.400 154.300 213.200 154.400 ;
        RECT 212.400 153.700 222.700 154.300 ;
        RECT 212.400 153.600 213.200 153.700 ;
    END
  END sine[13]
  PIN sine[14]
    PORT
      LAYER metal1 ;
        RECT 217.200 151.800 218.000 159.800 ;
        RECT 217.400 149.600 218.000 151.800 ;
        RECT 217.200 148.300 218.000 149.600 ;
        RECT 218.800 148.300 219.600 148.400 ;
        RECT 217.200 147.700 219.600 148.300 ;
        RECT 217.200 142.200 218.000 147.700 ;
        RECT 218.800 147.600 219.600 147.700 ;
      LAYER metal2 ;
        RECT 218.800 149.600 219.600 150.400 ;
        RECT 218.900 148.400 219.500 149.600 ;
        RECT 218.800 147.600 219.600 148.400 ;
      LAYER metal3 ;
        RECT 218.800 150.300 219.600 150.400 ;
        RECT 218.800 149.700 222.700 150.300 ;
        RECT 218.800 149.600 219.600 149.700 ;
    END
  END sine[14]
  PIN sine[15]
    PORT
      LAYER metal1 ;
        RECT 6.000 111.800 6.800 119.800 ;
        RECT 6.000 109.600 6.600 111.800 ;
        RECT 6.000 102.200 6.800 109.600 ;
      LAYER via1 ;
        RECT 6.000 117.600 6.800 118.400 ;
      LAYER metal2 ;
        RECT 6.000 117.600 6.800 118.400 ;
      LAYER metal3 ;
        RECT 6.000 118.300 6.800 118.400 ;
        RECT -1.900 117.700 6.800 118.300 ;
        RECT 6.000 117.600 6.800 117.700 ;
    END
  END sine[15]
  PIN cosine[0]
    PORT
      LAYER metal1 ;
        RECT 1.200 191.800 2.000 199.800 ;
        RECT 1.200 189.600 1.800 191.800 ;
        RECT 1.200 182.200 2.000 189.600 ;
      LAYER via1 ;
        RECT 1.200 187.600 2.000 188.400 ;
      LAYER metal2 ;
        RECT 1.200 189.600 2.000 190.400 ;
        RECT 1.300 188.400 1.900 189.600 ;
        RECT 1.200 187.600 2.000 188.400 ;
      LAYER metal3 ;
        RECT 1.200 190.300 2.000 190.400 ;
        RECT -1.900 189.700 2.000 190.300 ;
        RECT 1.200 189.600 2.000 189.700 ;
    END
  END cosine[0]
  PIN cosine[1]
    PORT
      LAYER metal1 ;
        RECT 42.800 191.800 43.600 199.800 ;
        RECT 43.000 189.600 43.600 191.800 ;
        RECT 42.800 182.200 43.600 189.600 ;
      LAYER via1 ;
        RECT 42.800 197.600 43.600 198.400 ;
      LAYER metal2 ;
        RECT 41.300 203.700 43.500 204.300 ;
        RECT 42.900 198.400 43.500 203.700 ;
        RECT 42.800 197.600 43.600 198.400 ;
    END
  END cosine[1]
  PIN cosine[2]
    PORT
      LAYER metal1 ;
        RECT 105.200 191.800 106.000 199.800 ;
        RECT 105.400 189.600 106.000 191.800 ;
        RECT 105.200 182.200 106.000 189.600 ;
      LAYER via1 ;
        RECT 105.200 197.600 106.000 198.400 ;
      LAYER metal2 ;
        RECT 105.300 198.400 105.900 204.300 ;
        RECT 105.200 197.600 106.000 198.400 ;
    END
  END cosine[2]
  PIN cosine[3]
    PORT
      LAYER metal1 ;
        RECT 36.400 172.400 37.200 179.800 ;
        RECT 36.400 170.200 37.000 172.400 ;
        RECT 36.400 162.200 37.200 170.200 ;
      LAYER via1 ;
        RECT 36.400 177.600 37.200 178.400 ;
      LAYER metal2 ;
        RECT 36.500 203.700 38.700 204.300 ;
        RECT 36.500 178.400 37.100 203.700 ;
        RECT 36.400 177.600 37.200 178.400 ;
    END
  END cosine[3]
  PIN cosine[4]
    PORT
      LAYER metal1 ;
        RECT 6.000 151.800 6.800 159.800 ;
        RECT 6.000 149.600 6.600 151.800 ;
        RECT 6.000 142.200 6.800 149.600 ;
      LAYER via1 ;
        RECT 6.000 155.600 6.800 156.400 ;
      LAYER metal2 ;
        RECT 6.000 155.600 6.800 156.400 ;
      LAYER metal3 ;
        RECT 6.000 156.300 6.800 156.400 ;
        RECT -1.900 155.700 6.800 156.300 ;
        RECT 6.000 155.600 6.800 155.700 ;
    END
  END cosine[4]
  PIN cosine[5]
    PORT
      LAYER metal1 ;
        RECT 1.200 151.800 2.000 159.800 ;
        RECT 1.200 149.600 1.800 151.800 ;
        RECT 1.200 142.200 2.000 149.600 ;
      LAYER via1 ;
        RECT 1.200 153.600 2.000 154.400 ;
      LAYER metal2 ;
        RECT 1.200 153.600 2.000 154.400 ;
        RECT 1.300 152.400 1.900 153.600 ;
        RECT 1.200 151.600 2.000 152.400 ;
      LAYER metal3 ;
        RECT 1.200 152.300 2.000 152.400 ;
        RECT -1.900 151.700 2.000 152.300 ;
        RECT 1.200 151.600 2.000 151.700 ;
    END
  END cosine[5]
  PIN cosine[6]
    PORT
      LAYER metal1 ;
        RECT 1.200 111.800 2.000 119.800 ;
        RECT 1.200 109.600 1.800 111.800 ;
        RECT 1.200 102.200 2.000 109.600 ;
      LAYER via1 ;
        RECT 1.200 113.600 2.000 114.400 ;
      LAYER metal2 ;
        RECT 1.200 113.600 2.000 114.400 ;
      LAYER metal3 ;
        RECT 1.200 114.300 2.000 114.400 ;
        RECT -1.900 113.700 2.000 114.300 ;
        RECT 1.200 113.600 2.000 113.700 ;
    END
  END cosine[6]
  PIN cosine[7]
    PORT
      LAYER metal1 ;
        RECT 1.200 71.800 2.000 79.800 ;
        RECT 1.200 69.600 1.800 71.800 ;
        RECT 1.200 62.200 2.000 69.600 ;
      LAYER via1 ;
        RECT 1.200 73.600 2.000 74.400 ;
      LAYER metal2 ;
        RECT 1.200 73.600 2.000 74.400 ;
      LAYER metal3 ;
        RECT 1.200 74.300 2.000 74.400 ;
        RECT -1.900 73.700 2.000 74.300 ;
        RECT 1.200 73.600 2.000 73.700 ;
    END
  END cosine[7]
  PIN cosine[8]
    PORT
      LAYER metal1 ;
        RECT 1.200 12.400 2.000 19.800 ;
        RECT 1.200 10.200 1.800 12.400 ;
        RECT 1.200 2.200 2.000 10.200 ;
      LAYER via1 ;
        RECT 1.200 7.600 2.000 8.400 ;
      LAYER metal2 ;
        RECT 1.200 9.600 2.000 10.400 ;
        RECT 1.300 8.400 1.900 9.600 ;
        RECT 1.200 7.600 2.000 8.400 ;
      LAYER metal3 ;
        RECT 1.200 10.300 2.000 10.400 ;
        RECT -1.900 9.700 2.000 10.300 ;
        RECT 1.200 9.600 2.000 9.700 ;
    END
  END cosine[8]
  PIN cosine[9]
    PORT
      LAYER metal1 ;
        RECT 1.200 31.800 2.000 39.800 ;
        RECT 1.200 29.600 1.800 31.800 ;
        RECT 1.200 22.200 2.000 29.600 ;
      LAYER via1 ;
        RECT 1.200 33.600 2.000 34.400 ;
      LAYER metal2 ;
        RECT 1.200 33.600 2.000 34.400 ;
      LAYER metal3 ;
        RECT 1.200 34.300 2.000 34.400 ;
        RECT -1.900 33.700 2.000 34.300 ;
        RECT 1.200 33.600 2.000 33.700 ;
    END
  END cosine[9]
  PIN cosine[10]
    PORT
      LAYER metal1 ;
        RECT 6.000 71.800 6.800 79.800 ;
        RECT 6.000 69.600 6.600 71.800 ;
        RECT 6.000 62.200 6.800 69.600 ;
      LAYER via1 ;
        RECT 6.000 67.600 6.800 68.400 ;
      LAYER metal2 ;
        RECT 6.000 69.600 6.800 70.400 ;
        RECT 6.100 68.400 6.700 69.600 ;
        RECT 6.000 67.600 6.800 68.400 ;
      LAYER metal3 ;
        RECT 6.000 70.300 6.800 70.400 ;
        RECT -1.900 69.700 6.800 70.300 ;
        RECT 6.000 69.600 6.800 69.700 ;
    END
  END cosine[10]
  PIN cosine[11]
    PORT
      LAYER metal1 ;
        RECT 41.200 12.400 42.000 19.800 ;
        RECT 41.200 10.200 41.800 12.400 ;
        RECT 41.200 2.200 42.000 10.200 ;
      LAYER via1 ;
        RECT 41.200 3.600 42.000 4.400 ;
      LAYER metal2 ;
        RECT 41.200 3.600 42.000 4.400 ;
        RECT 41.300 -1.700 41.900 3.600 ;
        RECT 41.300 -2.300 43.500 -1.700 ;
    END
  END cosine[11]
  PIN cosine[12]
    PORT
      LAYER metal1 ;
        RECT 86.000 12.400 86.800 19.800 ;
        RECT 86.000 10.200 86.600 12.400 ;
        RECT 86.000 2.200 86.800 10.200 ;
      LAYER via1 ;
        RECT 86.000 3.600 86.800 4.400 ;
      LAYER metal2 ;
        RECT 86.000 3.600 86.800 4.400 ;
        RECT 86.100 -1.700 86.700 3.600 ;
        RECT 86.100 -2.300 88.300 -1.700 ;
    END
  END cosine[12]
  PIN cosine[13]
    PORT
      LAYER metal1 ;
        RECT 94.000 12.400 94.800 19.800 ;
        RECT 94.200 10.200 94.800 12.400 ;
        RECT 94.000 2.200 94.800 10.200 ;
      LAYER via1 ;
        RECT 94.000 3.600 94.800 4.400 ;
      LAYER metal2 ;
        RECT 94.000 3.600 94.800 4.400 ;
        RECT 94.100 -1.700 94.700 3.600 ;
        RECT 92.500 -2.300 94.700 -1.700 ;
    END
  END cosine[13]
  PIN cosine[14]
    PORT
      LAYER metal1 ;
        RECT 34.800 111.800 35.600 119.800 ;
        RECT 34.800 109.600 35.400 111.800 ;
        RECT 34.800 102.200 35.600 109.600 ;
      LAYER via1 ;
        RECT 34.800 117.600 35.600 118.400 ;
      LAYER metal2 ;
        RECT 34.800 121.600 35.600 122.400 ;
        RECT 34.900 118.400 35.500 121.600 ;
        RECT 34.800 117.600 35.600 118.400 ;
      LAYER metal3 ;
        RECT 34.800 122.300 35.600 122.400 ;
        RECT -1.900 121.700 35.600 122.300 ;
        RECT 34.800 121.600 35.600 121.700 ;
    END
  END cosine[14]
  PIN cosine[15]
    PORT
      LAYER metal1 ;
        RECT 98.800 12.400 99.600 19.800 ;
        RECT 99.000 10.200 99.600 12.400 ;
        RECT 98.800 2.200 99.600 10.200 ;
      LAYER via1 ;
        RECT 98.800 3.600 99.600 4.400 ;
      LAYER metal2 ;
        RECT 98.800 3.600 99.600 4.400 ;
        RECT 98.900 -1.700 99.500 3.600 ;
        RECT 97.300 -2.300 99.500 -1.700 ;
    END
  END cosine[15]
  OBS
      LAYER metal1 ;
        RECT 4.400 192.400 5.200 199.800 ;
        RECT 3.000 191.800 5.200 192.400 ;
        RECT 6.000 192.400 6.800 199.800 ;
        RECT 7.800 192.400 8.600 192.600 ;
        RECT 6.000 191.800 8.600 192.400 ;
        RECT 10.400 191.800 12.000 199.800 ;
        RECT 14.000 192.400 14.800 192.600 ;
        RECT 15.600 192.400 16.400 199.800 ;
        RECT 14.000 191.800 16.400 192.400 ;
        RECT 3.000 191.200 3.600 191.800 ;
        RECT 2.400 190.400 3.600 191.200 ;
        RECT 9.000 190.400 9.800 190.600 ;
        RECT 11.000 190.400 11.600 191.800 ;
        RECT 3.000 187.400 3.600 190.400 ;
        RECT 4.400 190.300 5.200 190.400 ;
        RECT 4.400 189.700 6.700 190.300 ;
        RECT 4.400 188.800 5.200 189.700 ;
        RECT 6.100 188.400 6.700 189.700 ;
        RECT 8.200 189.800 9.800 190.400 ;
        RECT 8.200 189.600 9.000 189.800 ;
        RECT 10.800 189.600 11.600 190.400 ;
        RECT 9.600 188.600 10.400 188.800 ;
        RECT 7.600 188.400 10.400 188.600 ;
        RECT 6.000 188.000 10.400 188.400 ;
        RECT 11.000 188.400 11.600 189.600 ;
        RECT 18.800 190.300 19.600 199.800 ;
        RECT 20.600 199.200 24.200 199.800 ;
        RECT 20.600 199.000 21.200 199.200 ;
        RECT 20.400 193.000 21.200 199.000 ;
        RECT 23.600 199.000 24.200 199.200 ;
        RECT 25.200 199.200 29.200 199.800 ;
        RECT 22.000 193.000 22.800 198.600 ;
        RECT 23.600 193.400 24.400 199.000 ;
        RECT 25.200 194.000 26.000 199.200 ;
        RECT 26.800 193.800 27.600 198.600 ;
        RECT 28.400 193.800 29.200 199.200 ;
        RECT 26.800 193.400 27.400 193.800 ;
        RECT 23.600 193.000 27.400 193.400 ;
        RECT 22.200 192.400 22.800 193.000 ;
        RECT 23.800 192.800 27.400 193.000 ;
        RECT 28.600 193.200 29.200 193.800 ;
        RECT 31.600 193.800 32.400 199.800 ;
        RECT 31.600 193.200 32.200 193.800 ;
        RECT 28.600 192.600 32.200 193.200 ;
        RECT 35.800 192.400 36.600 199.800 ;
        RECT 37.200 193.600 38.000 194.400 ;
        RECT 37.400 192.400 38.000 193.600 ;
        RECT 39.600 192.400 40.400 199.800 ;
        RECT 22.000 192.200 22.800 192.400 ;
        RECT 22.000 191.600 25.400 192.200 ;
        RECT 34.800 191.600 36.800 192.400 ;
        RECT 37.400 191.800 38.800 192.400 ;
        RECT 39.600 191.800 41.800 192.400 ;
        RECT 38.000 191.600 38.800 191.800 ;
        RECT 22.000 190.300 22.800 190.400 ;
        RECT 18.800 189.700 22.800 190.300 ;
        RECT 6.000 187.800 8.200 188.000 ;
        RECT 11.000 187.800 12.000 188.400 ;
        RECT 6.000 187.600 7.600 187.800 ;
        RECT 3.000 186.800 5.200 187.400 ;
        RECT 7.800 186.800 8.600 187.000 ;
        RECT 4.400 182.200 5.200 186.800 ;
        RECT 6.000 186.200 8.600 186.800 ;
        RECT 9.200 186.400 10.800 187.200 ;
        RECT 6.000 182.200 6.800 186.200 ;
        RECT 11.400 185.800 12.000 187.800 ;
        RECT 12.800 187.600 13.600 188.400 ;
        RECT 14.800 188.300 16.400 188.400 ;
        RECT 14.800 187.700 17.900 188.300 ;
        RECT 14.800 187.600 16.400 187.700 ;
        RECT 12.800 187.200 13.400 187.600 ;
        RECT 12.600 186.400 13.400 187.200 ;
        RECT 14.000 186.800 14.800 187.000 ;
        RECT 14.000 186.200 16.400 186.800 ;
        RECT 17.300 186.400 17.900 187.700 ;
        RECT 10.400 182.200 12.000 185.800 ;
        RECT 15.600 182.200 16.400 186.200 ;
        RECT 17.200 184.800 18.000 186.400 ;
        RECT 18.800 182.200 19.600 189.700 ;
        RECT 22.000 189.600 22.800 189.700 ;
        RECT 24.800 185.000 25.400 191.600 ;
        RECT 26.000 190.300 27.600 190.400 ;
        RECT 34.800 190.300 35.600 190.400 ;
        RECT 26.000 189.700 35.600 190.300 ;
        RECT 26.000 189.600 27.600 189.700 ;
        RECT 34.800 188.800 35.600 189.700 ;
        RECT 36.200 188.400 36.800 191.600 ;
        RECT 38.100 190.400 38.700 191.600 ;
        RECT 41.200 191.200 41.800 191.800 ;
        RECT 41.200 190.400 42.400 191.200 ;
        RECT 38.000 190.300 38.800 190.400 ;
        RECT 39.600 190.300 40.400 190.400 ;
        RECT 38.000 189.700 40.400 190.300 ;
        RECT 38.000 189.600 38.800 189.700 ;
        RECT 39.600 188.800 40.400 189.700 ;
        RECT 27.600 187.600 29.200 188.400 ;
        RECT 33.200 188.300 34.000 188.400 ;
        RECT 31.700 188.200 34.000 188.300 ;
        RECT 31.700 187.700 34.800 188.200 ;
        RECT 28.400 186.300 30.800 186.400 ;
        RECT 31.700 186.300 32.300 187.700 ;
        RECT 33.200 187.600 34.800 187.700 ;
        RECT 36.200 187.600 38.800 188.400 ;
        RECT 34.000 187.200 34.800 187.600 ;
        RECT 28.400 185.700 32.300 186.300 ;
        RECT 33.400 186.200 37.000 186.600 ;
        RECT 38.000 186.200 38.600 187.600 ;
        RECT 41.200 187.400 41.800 190.400 ;
        RECT 39.600 186.800 41.800 187.400 ;
        RECT 33.200 186.000 37.200 186.200 ;
        RECT 28.400 185.600 30.800 185.700 ;
        RECT 24.800 184.400 28.800 185.000 ;
        RECT 24.800 184.200 26.000 184.400 ;
        RECT 25.200 182.200 26.000 184.200 ;
        RECT 28.200 183.600 29.200 184.400 ;
        RECT 28.400 182.200 29.200 183.600 ;
        RECT 33.200 182.200 34.000 186.000 ;
        RECT 36.400 182.200 37.200 186.000 ;
        RECT 38.000 182.200 38.800 186.200 ;
        RECT 39.600 182.200 40.400 186.800 ;
        RECT 44.400 184.800 45.200 186.400 ;
        RECT 46.000 182.200 46.800 199.800 ;
        RECT 49.200 195.800 50.000 199.800 ;
        RECT 49.400 195.600 50.000 195.800 ;
        RECT 52.400 195.800 53.200 199.800 ;
        RECT 52.400 195.600 53.000 195.800 ;
        RECT 49.400 195.000 53.000 195.600 ;
        RECT 50.800 192.800 51.600 194.400 ;
        RECT 52.400 192.400 53.000 195.000 ;
        RECT 47.600 190.800 48.400 192.400 ;
        RECT 52.400 191.600 53.200 192.400 ;
        RECT 49.200 189.600 50.800 190.400 ;
        RECT 52.400 188.400 53.000 191.600 ;
        RECT 51.400 188.200 53.200 188.400 ;
        RECT 51.200 187.600 53.200 188.200 ;
        RECT 51.200 182.200 52.000 187.600 ;
        RECT 54.000 182.200 54.800 199.800 ;
        RECT 57.200 186.800 58.000 188.400 ;
        RECT 55.600 184.800 56.400 186.400 ;
        RECT 58.800 186.200 59.600 199.800 ;
        RECT 60.400 191.600 61.200 193.200 ;
        RECT 68.400 192.000 69.200 199.800 ;
        RECT 71.600 195.200 72.400 199.800 ;
        RECT 68.200 191.200 69.200 192.000 ;
        RECT 69.800 194.600 72.400 195.200 ;
        RECT 69.800 193.000 70.400 194.600 ;
        RECT 74.800 194.400 75.600 199.800 ;
        RECT 78.000 197.000 78.800 199.800 ;
        RECT 79.600 197.000 80.400 199.800 ;
        RECT 81.200 197.000 82.000 199.800 ;
        RECT 76.200 194.400 80.400 195.200 ;
        RECT 73.000 193.600 75.600 194.400 ;
        RECT 82.800 193.600 83.600 199.800 ;
        RECT 86.000 195.000 86.800 199.800 ;
        RECT 89.200 195.000 90.000 199.800 ;
        RECT 90.800 197.000 91.600 199.800 ;
        RECT 92.400 197.000 93.200 199.800 ;
        RECT 95.600 195.200 96.400 199.800 ;
        RECT 98.800 196.400 99.600 199.800 ;
        RECT 98.800 195.800 99.800 196.400 ;
        RECT 99.200 195.200 99.800 195.800 ;
        RECT 94.400 194.400 98.600 195.200 ;
        RECT 99.200 194.600 101.200 195.200 ;
        RECT 86.000 193.600 88.600 194.400 ;
        RECT 89.200 193.800 95.000 194.400 ;
        RECT 98.000 194.000 98.600 194.400 ;
        RECT 78.000 193.000 78.800 193.200 ;
        RECT 69.800 192.400 78.800 193.000 ;
        RECT 81.200 193.000 82.000 193.200 ;
        RECT 89.200 193.000 89.800 193.800 ;
        RECT 95.600 193.200 97.000 193.800 ;
        RECT 98.000 193.200 99.600 194.000 ;
        RECT 81.200 192.400 89.800 193.000 ;
        RECT 90.800 193.000 97.000 193.200 ;
        RECT 90.800 192.600 96.200 193.000 ;
        RECT 90.800 192.400 91.600 192.600 ;
        RECT 68.200 186.800 69.000 191.200 ;
        RECT 69.800 190.600 70.400 192.400 ;
        RECT 69.600 190.000 70.400 190.600 ;
        RECT 76.400 190.000 99.800 190.600 ;
        RECT 69.600 188.000 70.200 190.000 ;
        RECT 76.400 189.400 77.200 190.000 ;
        RECT 94.000 189.600 94.800 190.000 ;
        RECT 97.200 189.600 98.000 190.000 ;
        RECT 99.000 189.800 99.800 190.000 ;
        RECT 70.800 188.600 74.600 189.400 ;
        RECT 69.600 187.400 70.800 188.000 ;
        RECT 58.800 185.600 60.600 186.200 ;
        RECT 68.200 186.000 69.200 186.800 ;
        RECT 59.800 182.200 60.600 185.600 ;
        RECT 68.400 182.200 69.200 186.000 ;
        RECT 70.000 182.200 70.800 187.400 ;
        RECT 73.800 187.400 74.600 188.600 ;
        RECT 73.800 186.800 75.600 187.400 ;
        RECT 74.800 186.200 75.600 186.800 ;
        RECT 79.600 186.400 80.400 189.200 ;
        RECT 82.800 188.600 86.000 189.400 ;
        RECT 89.800 188.600 91.800 189.400 ;
        RECT 100.400 189.000 101.200 194.600 ;
        RECT 102.000 192.400 102.800 199.800 ;
        RECT 108.400 196.400 109.200 199.800 ;
        RECT 108.200 195.800 109.200 196.400 ;
        RECT 108.200 195.200 108.800 195.800 ;
        RECT 111.600 195.200 112.400 199.800 ;
        RECT 114.800 197.000 115.600 199.800 ;
        RECT 116.400 197.000 117.200 199.800 ;
        RECT 106.800 194.600 108.800 195.200 ;
        RECT 102.000 191.800 104.200 192.400 ;
        RECT 103.600 191.200 104.200 191.800 ;
        RECT 103.600 190.400 104.800 191.200 ;
        RECT 82.400 187.800 83.200 188.000 ;
        RECT 82.400 187.200 86.800 187.800 ;
        RECT 86.000 187.000 86.800 187.200 ;
        RECT 87.600 186.800 88.400 188.400 ;
        RECT 74.800 185.400 77.200 186.200 ;
        RECT 79.600 185.600 80.600 186.400 ;
        RECT 83.600 185.600 85.200 186.400 ;
        RECT 86.000 186.200 86.800 186.400 ;
        RECT 89.800 186.200 90.600 188.600 ;
        RECT 92.400 188.200 101.200 189.000 ;
        RECT 102.000 188.800 102.800 190.400 ;
        RECT 95.800 186.800 98.800 187.600 ;
        RECT 95.800 186.200 96.600 186.800 ;
        RECT 86.000 185.600 90.600 186.200 ;
        RECT 76.400 182.200 77.200 185.400 ;
        RECT 94.000 185.400 96.600 186.200 ;
        RECT 78.000 182.200 78.800 185.000 ;
        RECT 79.600 182.200 80.400 185.000 ;
        RECT 81.200 182.200 82.000 185.000 ;
        RECT 82.800 182.200 83.600 185.000 ;
        RECT 86.000 182.200 86.800 185.000 ;
        RECT 89.200 182.200 90.000 185.000 ;
        RECT 90.800 182.200 91.600 185.000 ;
        RECT 92.400 182.200 93.200 185.000 ;
        RECT 94.000 182.200 94.800 185.400 ;
        RECT 100.400 182.200 101.200 188.200 ;
        RECT 103.600 187.400 104.200 190.400 ;
        RECT 102.000 186.800 104.200 187.400 ;
        RECT 106.800 189.000 107.600 194.600 ;
        RECT 109.400 194.400 113.600 195.200 ;
        RECT 118.000 195.000 118.800 199.800 ;
        RECT 121.200 195.000 122.000 199.800 ;
        RECT 109.400 194.000 110.000 194.400 ;
        RECT 108.400 193.200 110.000 194.000 ;
        RECT 113.000 193.800 118.800 194.400 ;
        RECT 111.000 193.200 112.400 193.800 ;
        RECT 111.000 193.000 117.200 193.200 ;
        RECT 111.800 192.600 117.200 193.000 ;
        RECT 116.400 192.400 117.200 192.600 ;
        RECT 118.200 193.000 118.800 193.800 ;
        RECT 119.400 193.600 122.000 194.400 ;
        RECT 124.400 193.600 125.200 199.800 ;
        RECT 126.000 197.000 126.800 199.800 ;
        RECT 127.600 197.000 128.400 199.800 ;
        RECT 129.200 197.000 130.000 199.800 ;
        RECT 127.600 194.400 131.800 195.200 ;
        RECT 132.400 194.400 133.200 199.800 ;
        RECT 135.600 195.200 136.400 199.800 ;
        RECT 135.600 194.600 138.200 195.200 ;
        RECT 132.400 193.600 135.000 194.400 ;
        RECT 126.000 193.000 126.800 193.200 ;
        RECT 118.200 192.400 126.800 193.000 ;
        RECT 129.200 193.000 130.000 193.200 ;
        RECT 137.600 193.000 138.200 194.600 ;
        RECT 129.200 192.400 138.200 193.000 ;
        RECT 137.600 190.600 138.200 192.400 ;
        RECT 138.800 192.000 139.600 199.800 ;
        RECT 145.200 192.400 146.000 199.800 ;
        RECT 138.800 191.200 139.800 192.000 ;
        RECT 143.800 191.800 146.000 192.400 ;
        RECT 146.800 192.400 147.600 199.800 ;
        RECT 148.400 192.400 149.200 192.600 ;
        RECT 151.200 192.400 152.800 199.800 ;
        RECT 146.800 191.800 149.200 192.400 ;
        RECT 150.000 191.800 152.800 192.400 ;
        RECT 155.000 192.400 155.800 192.600 ;
        RECT 156.400 192.400 157.200 199.800 ;
        RECT 155.000 191.800 157.200 192.400 ;
        RECT 162.800 192.400 163.600 199.800 ;
        RECT 162.800 191.800 165.000 192.400 ;
        RECT 143.800 191.200 144.400 191.800 ;
        RECT 150.000 191.600 151.400 191.800 ;
        RECT 108.200 190.000 131.600 190.600 ;
        RECT 137.600 190.000 138.400 190.600 ;
        RECT 108.200 189.800 109.000 190.000 ;
        RECT 110.000 189.600 110.800 190.000 ;
        RECT 113.200 189.600 114.000 190.000 ;
        RECT 130.800 189.400 131.600 190.000 ;
        RECT 106.800 188.200 115.600 189.000 ;
        RECT 116.200 188.600 118.200 189.400 ;
        RECT 122.000 188.600 125.200 189.400 ;
        RECT 102.000 182.200 102.800 186.800 ;
        RECT 106.800 182.200 107.600 188.200 ;
        RECT 109.200 186.800 112.200 187.600 ;
        RECT 111.400 186.200 112.200 186.800 ;
        RECT 117.400 186.200 118.200 188.600 ;
        RECT 119.600 186.800 120.400 188.400 ;
        RECT 124.800 187.800 125.600 188.000 ;
        RECT 121.200 187.200 125.600 187.800 ;
        RECT 121.200 187.000 122.000 187.200 ;
        RECT 127.600 186.400 128.400 189.200 ;
        RECT 133.400 188.600 137.200 189.400 ;
        RECT 133.400 187.400 134.200 188.600 ;
        RECT 137.800 188.000 138.400 190.000 ;
        RECT 121.200 186.200 122.000 186.400 ;
        RECT 111.400 185.400 114.000 186.200 ;
        RECT 117.400 185.600 122.000 186.200 ;
        RECT 122.800 185.600 124.400 186.400 ;
        RECT 127.400 185.600 128.400 186.400 ;
        RECT 132.400 186.800 134.200 187.400 ;
        RECT 137.200 187.400 138.400 188.000 ;
        RECT 132.400 186.200 133.200 186.800 ;
        RECT 113.200 182.200 114.000 185.400 ;
        RECT 130.800 185.400 133.200 186.200 ;
        RECT 114.800 182.200 115.600 185.000 ;
        RECT 116.400 182.200 117.200 185.000 ;
        RECT 118.000 182.200 118.800 185.000 ;
        RECT 121.200 182.200 122.000 185.000 ;
        RECT 124.400 182.200 125.200 185.000 ;
        RECT 126.000 182.200 126.800 185.000 ;
        RECT 127.600 182.200 128.400 185.000 ;
        RECT 129.200 182.200 130.000 185.000 ;
        RECT 130.800 182.200 131.600 185.400 ;
        RECT 137.200 182.200 138.000 187.400 ;
        RECT 139.000 186.800 139.800 191.200 ;
        RECT 143.200 190.400 144.400 191.200 ;
        RECT 150.800 190.400 151.400 191.600 ;
        RECT 155.000 191.200 155.600 191.800 ;
        RECT 152.200 190.600 155.600 191.200 ;
        RECT 164.400 191.200 165.000 191.800 ;
        RECT 152.200 190.400 153.000 190.600 ;
        RECT 164.400 190.400 165.600 191.200 ;
        RECT 143.800 187.400 144.400 190.400 ;
        RECT 145.200 190.300 146.000 190.400 ;
        RECT 145.200 189.700 147.500 190.300 ;
        RECT 145.200 188.800 146.000 189.700 ;
        RECT 146.900 188.400 147.500 189.700 ;
        RECT 150.000 189.800 151.400 190.400 ;
        RECT 154.400 189.800 155.200 190.000 ;
        RECT 150.000 189.600 151.800 189.800 ;
        RECT 150.800 189.200 151.800 189.600 ;
        RECT 146.800 187.600 148.400 188.400 ;
        RECT 149.600 187.600 150.400 188.400 ;
        RECT 143.800 186.800 146.000 187.400 ;
        RECT 149.800 187.200 150.400 187.600 ;
        RECT 148.400 186.800 149.200 187.000 ;
        RECT 138.800 186.000 139.800 186.800 ;
        RECT 138.800 182.200 139.600 186.000 ;
        RECT 145.200 182.200 146.000 186.800 ;
        RECT 146.800 186.200 149.200 186.800 ;
        RECT 149.800 186.400 150.600 187.200 ;
        RECT 146.800 182.200 147.600 186.200 ;
        RECT 151.200 185.800 151.800 189.200 ;
        RECT 152.600 189.200 155.200 189.800 ;
        RECT 152.600 188.600 153.200 189.200 ;
        RECT 162.800 188.800 163.600 190.400 ;
        RECT 152.400 187.800 153.200 188.600 ;
        RECT 155.600 188.200 157.200 188.400 ;
        RECT 153.800 187.600 157.200 188.200 ;
        RECT 153.800 187.200 154.400 187.600 ;
        RECT 164.400 187.400 165.000 190.400 ;
        RECT 152.400 186.600 154.400 187.200 ;
        RECT 155.000 186.800 155.800 187.000 ;
        RECT 162.800 186.800 165.000 187.400 ;
        RECT 169.200 190.300 170.000 199.800 ;
        RECT 173.400 192.600 174.200 199.800 ;
        RECT 177.200 195.800 178.000 199.800 ;
        RECT 172.400 191.800 174.200 192.600 ;
        RECT 170.800 190.300 171.600 190.400 ;
        RECT 169.200 189.700 171.600 190.300 ;
        RECT 152.400 186.400 154.000 186.600 ;
        RECT 155.000 186.200 157.200 186.800 ;
        RECT 151.200 182.200 152.800 185.800 ;
        RECT 156.400 182.200 157.200 186.200 ;
        RECT 162.800 182.200 163.600 186.800 ;
        RECT 167.600 184.800 168.400 186.400 ;
        RECT 169.200 182.200 170.000 189.700 ;
        RECT 170.800 189.600 171.600 189.700 ;
        RECT 172.600 188.400 173.200 191.800 ;
        RECT 177.400 191.600 178.000 195.800 ;
        RECT 180.400 191.800 181.200 199.800 ;
        RECT 183.600 196.400 184.400 199.800 ;
        RECT 183.400 195.800 184.400 196.400 ;
        RECT 183.400 195.200 184.000 195.800 ;
        RECT 186.800 195.200 187.600 199.800 ;
        RECT 190.000 197.000 190.800 199.800 ;
        RECT 191.600 197.000 192.400 199.800 ;
        RECT 174.000 189.600 174.800 191.200 ;
        RECT 177.400 191.000 179.800 191.600 ;
        RECT 177.200 189.600 178.000 190.400 ;
        RECT 172.400 188.300 173.200 188.400 ;
        RECT 175.600 188.300 176.400 189.200 ;
        RECT 177.400 188.800 178.000 189.600 ;
        RECT 172.400 187.700 176.400 188.300 ;
        RECT 177.200 188.000 178.400 188.800 ;
        RECT 172.400 187.600 173.200 187.700 ;
        RECT 175.600 187.600 176.400 187.700 ;
        RECT 179.200 187.600 179.800 191.000 ;
        RECT 180.600 190.400 181.200 191.800 ;
        RECT 180.400 189.600 181.200 190.400 ;
        RECT 170.800 184.800 171.600 186.400 ;
        RECT 172.600 184.400 173.200 187.600 ;
        RECT 179.200 187.400 180.000 187.600 ;
        RECT 177.000 187.000 180.000 187.400 ;
        RECT 175.800 186.800 180.000 187.000 ;
        RECT 175.800 186.400 177.600 186.800 ;
        RECT 175.800 186.200 176.400 186.400 ;
        RECT 180.600 186.200 181.200 189.600 ;
        RECT 172.400 182.200 173.200 184.400 ;
        RECT 175.600 182.200 176.400 186.200 ;
        RECT 179.800 185.200 181.200 186.200 ;
        RECT 182.000 194.600 184.000 195.200 ;
        RECT 182.000 189.000 182.800 194.600 ;
        RECT 184.600 194.400 188.800 195.200 ;
        RECT 193.200 195.000 194.000 199.800 ;
        RECT 196.400 195.000 197.200 199.800 ;
        RECT 184.600 194.000 185.200 194.400 ;
        RECT 183.600 193.200 185.200 194.000 ;
        RECT 188.200 193.800 194.000 194.400 ;
        RECT 186.200 193.200 187.600 193.800 ;
        RECT 186.200 193.000 192.400 193.200 ;
        RECT 187.000 192.600 192.400 193.000 ;
        RECT 191.600 192.400 192.400 192.600 ;
        RECT 193.400 193.000 194.000 193.800 ;
        RECT 194.600 193.600 197.200 194.400 ;
        RECT 199.600 193.600 200.400 199.800 ;
        RECT 201.200 197.000 202.000 199.800 ;
        RECT 202.800 197.000 203.600 199.800 ;
        RECT 204.400 197.000 205.200 199.800 ;
        RECT 202.800 194.400 207.000 195.200 ;
        RECT 207.600 194.400 208.400 199.800 ;
        RECT 210.800 195.200 211.600 199.800 ;
        RECT 210.800 194.600 213.400 195.200 ;
        RECT 207.600 193.600 210.200 194.400 ;
        RECT 201.200 193.000 202.000 193.200 ;
        RECT 193.400 192.400 202.000 193.000 ;
        RECT 204.400 193.000 205.200 193.200 ;
        RECT 212.800 193.000 213.400 194.600 ;
        RECT 204.400 192.400 213.400 193.000 ;
        RECT 212.800 190.600 213.400 192.400 ;
        RECT 214.000 192.000 214.800 199.800 ;
        RECT 214.000 191.200 215.000 192.000 ;
        RECT 183.400 190.000 206.800 190.600 ;
        RECT 212.800 190.000 213.600 190.600 ;
        RECT 183.400 189.800 184.200 190.000 ;
        RECT 185.200 189.600 186.000 190.000 ;
        RECT 188.400 189.600 189.200 190.000 ;
        RECT 206.000 189.400 206.800 190.000 ;
        RECT 182.000 188.200 190.800 189.000 ;
        RECT 191.400 188.600 193.400 189.400 ;
        RECT 197.200 188.600 200.400 189.400 ;
        RECT 179.800 184.400 180.600 185.200 ;
        RECT 179.800 183.600 181.200 184.400 ;
        RECT 179.800 182.200 180.600 183.600 ;
        RECT 182.000 182.200 182.800 188.200 ;
        RECT 184.400 186.800 187.400 187.600 ;
        RECT 186.600 186.200 187.400 186.800 ;
        RECT 192.600 186.200 193.400 188.600 ;
        RECT 194.800 186.800 195.600 188.400 ;
        RECT 200.000 187.800 200.800 188.000 ;
        RECT 196.400 187.200 200.800 187.800 ;
        RECT 196.400 187.000 197.200 187.200 ;
        RECT 202.800 186.400 203.600 189.200 ;
        RECT 208.600 188.600 212.400 189.400 ;
        RECT 208.600 187.400 209.400 188.600 ;
        RECT 213.000 188.000 213.600 190.000 ;
        RECT 196.400 186.200 197.200 186.400 ;
        RECT 186.600 185.400 189.200 186.200 ;
        RECT 192.600 185.600 197.200 186.200 ;
        RECT 198.000 185.600 199.600 186.400 ;
        RECT 202.600 185.600 203.600 186.400 ;
        RECT 207.600 186.800 209.400 187.400 ;
        RECT 212.400 187.400 213.600 188.000 ;
        RECT 207.600 186.200 208.400 186.800 ;
        RECT 188.400 182.200 189.200 185.400 ;
        RECT 206.000 185.400 208.400 186.200 ;
        RECT 190.000 182.200 190.800 185.000 ;
        RECT 191.600 182.200 192.400 185.000 ;
        RECT 193.200 182.200 194.000 185.000 ;
        RECT 196.400 182.200 197.200 185.000 ;
        RECT 199.600 182.200 200.400 185.000 ;
        RECT 201.200 182.200 202.000 185.000 ;
        RECT 202.800 182.200 203.600 185.000 ;
        RECT 204.400 182.200 205.200 185.000 ;
        RECT 206.000 182.200 206.800 185.400 ;
        RECT 212.400 182.200 213.200 187.400 ;
        RECT 214.200 186.800 215.000 191.200 ;
        RECT 214.000 186.000 215.000 186.800 ;
        RECT 214.000 182.200 214.800 186.000 ;
        RECT 2.800 176.000 3.600 179.800 ;
        RECT 2.600 175.200 3.600 176.000 ;
        RECT 2.600 170.800 3.400 175.200 ;
        RECT 4.400 174.600 5.200 179.800 ;
        RECT 10.800 176.600 11.600 179.800 ;
        RECT 12.400 177.000 13.200 179.800 ;
        RECT 14.000 177.000 14.800 179.800 ;
        RECT 15.600 177.000 16.400 179.800 ;
        RECT 17.200 177.000 18.000 179.800 ;
        RECT 20.400 177.000 21.200 179.800 ;
        RECT 23.600 177.000 24.400 179.800 ;
        RECT 25.200 177.000 26.000 179.800 ;
        RECT 26.800 177.000 27.600 179.800 ;
        RECT 9.200 175.800 11.600 176.600 ;
        RECT 28.400 176.600 29.200 179.800 ;
        RECT 9.200 175.200 10.000 175.800 ;
        RECT 4.000 174.000 5.200 174.600 ;
        RECT 8.200 174.600 10.000 175.200 ;
        RECT 14.000 175.600 15.000 176.400 ;
        RECT 18.000 175.600 19.600 176.400 ;
        RECT 20.400 175.800 25.000 176.400 ;
        RECT 28.400 175.800 31.000 176.600 ;
        RECT 20.400 175.600 21.200 175.800 ;
        RECT 4.000 172.000 4.600 174.000 ;
        RECT 8.200 173.400 9.000 174.600 ;
        RECT 5.200 172.600 9.000 173.400 ;
        RECT 14.000 172.800 14.800 175.600 ;
        RECT 20.400 174.800 21.200 175.000 ;
        RECT 16.800 174.200 21.200 174.800 ;
        RECT 16.800 174.000 17.600 174.200 ;
        RECT 22.000 173.600 22.800 175.200 ;
        RECT 24.200 173.400 25.000 175.800 ;
        RECT 30.200 175.200 31.000 175.800 ;
        RECT 30.200 174.400 33.200 175.200 ;
        RECT 34.800 173.800 35.600 179.800 ;
        RECT 39.600 175.200 40.400 179.800 ;
        RECT 17.200 172.600 20.400 173.400 ;
        RECT 24.200 172.600 26.200 173.400 ;
        RECT 26.800 173.000 35.600 173.800 ;
        RECT 4.000 171.400 4.800 172.000 ;
        RECT 2.600 170.000 3.600 170.800 ;
        RECT 2.800 162.200 3.600 170.000 ;
        RECT 4.200 169.600 4.800 171.400 ;
        RECT 5.400 170.800 6.200 171.000 ;
        RECT 5.400 170.200 32.400 170.800 ;
        RECT 28.200 170.000 29.000 170.200 ;
        RECT 31.600 169.600 32.400 170.200 ;
        RECT 4.200 169.000 13.200 169.600 ;
        RECT 4.200 167.400 4.800 169.000 ;
        RECT 12.400 168.800 13.200 169.000 ;
        RECT 15.600 169.000 24.200 169.600 ;
        RECT 15.600 168.800 16.400 169.000 ;
        RECT 7.400 167.600 10.000 168.400 ;
        RECT 4.200 166.800 6.800 167.400 ;
        RECT 6.000 162.200 6.800 166.800 ;
        RECT 9.200 162.200 10.000 167.600 ;
        RECT 10.600 166.800 14.800 167.600 ;
        RECT 12.400 162.200 13.200 165.000 ;
        RECT 14.000 162.200 14.800 165.000 ;
        RECT 15.600 162.200 16.400 165.000 ;
        RECT 17.200 162.200 18.000 168.400 ;
        RECT 20.400 167.600 23.000 168.400 ;
        RECT 23.600 168.200 24.200 169.000 ;
        RECT 25.200 169.400 26.000 169.600 ;
        RECT 25.200 169.000 30.600 169.400 ;
        RECT 25.200 168.800 31.400 169.000 ;
        RECT 30.000 168.200 31.400 168.800 ;
        RECT 23.600 167.600 29.400 168.200 ;
        RECT 32.400 168.000 34.000 168.800 ;
        RECT 32.400 167.600 33.000 168.000 ;
        RECT 20.400 162.200 21.200 167.000 ;
        RECT 23.600 162.200 24.400 167.000 ;
        RECT 28.800 166.800 33.000 167.600 ;
        RECT 34.800 167.400 35.600 173.000 ;
        RECT 38.200 174.600 40.400 175.200 ;
        RECT 38.200 171.600 38.800 174.600 ;
        RECT 42.400 174.200 43.200 179.800 ;
        RECT 41.400 173.800 43.200 174.200 ;
        RECT 41.400 173.600 43.000 173.800 ;
        RECT 39.600 171.600 40.400 173.200 ;
        RECT 37.600 170.800 38.800 171.600 ;
        RECT 38.200 170.200 38.800 170.800 ;
        RECT 41.400 170.400 42.000 173.600 ;
        RECT 43.600 171.600 45.200 172.400 ;
        RECT 38.200 169.600 40.400 170.200 ;
        RECT 41.200 169.600 42.000 170.400 ;
        RECT 46.000 169.600 46.800 171.200 ;
        RECT 33.600 166.800 35.600 167.400 ;
        RECT 25.200 162.200 26.000 165.000 ;
        RECT 26.800 162.200 27.600 165.000 ;
        RECT 30.000 162.200 30.800 166.800 ;
        RECT 33.600 166.200 34.200 166.800 ;
        RECT 33.200 165.600 34.200 166.200 ;
        RECT 33.200 162.200 34.000 165.600 ;
        RECT 39.600 162.200 40.400 169.600 ;
        RECT 41.400 167.000 42.000 169.600 ;
        RECT 42.800 167.600 43.600 169.200 ;
        RECT 41.400 166.400 45.000 167.000 ;
        RECT 41.400 166.200 42.000 166.400 ;
        RECT 41.200 162.200 42.000 166.200 ;
        RECT 44.400 166.200 45.000 166.400 ;
        RECT 44.400 162.200 45.200 166.200 ;
        RECT 47.600 162.200 48.400 179.800 ;
        RECT 49.200 175.600 50.000 177.200 ;
        RECT 49.200 168.300 50.000 168.400 ;
        RECT 50.800 168.300 51.600 179.800 ;
        RECT 52.400 175.600 53.200 177.200 ;
        RECT 54.000 175.800 54.800 179.800 ;
        RECT 55.600 176.000 56.400 179.800 ;
        RECT 58.800 176.000 59.600 179.800 ;
        RECT 68.400 178.400 69.200 179.800 ;
        RECT 68.400 177.600 69.400 178.400 ;
        RECT 71.600 177.800 72.400 179.800 ;
        RECT 71.600 177.600 72.800 177.800 ;
        RECT 68.800 177.000 72.800 177.600 ;
        RECT 66.800 176.300 69.200 176.400 ;
        RECT 55.600 175.800 59.600 176.000 ;
        RECT 54.200 174.400 54.800 175.800 ;
        RECT 55.800 175.400 59.400 175.800 ;
        RECT 60.500 175.700 69.200 176.300 ;
        RECT 58.000 174.400 58.800 174.800 ;
        RECT 54.000 173.600 56.600 174.400 ;
        RECT 58.000 174.300 59.600 174.400 ;
        RECT 60.500 174.300 61.100 175.700 ;
        RECT 66.800 175.600 69.200 175.700 ;
        RECT 58.000 173.800 61.100 174.300 ;
        RECT 58.800 173.700 61.100 173.800 ;
        RECT 58.800 173.600 59.600 173.700 ;
        RECT 68.400 173.600 70.000 174.400 ;
        RECT 56.000 172.400 56.600 173.600 ;
        RECT 55.600 171.600 56.600 172.400 ;
        RECT 57.200 172.300 58.000 173.200 ;
        RECT 70.000 172.300 71.600 172.400 ;
        RECT 57.200 171.700 71.600 172.300 ;
        RECT 57.200 171.600 58.000 171.700 ;
        RECT 70.000 171.600 71.600 171.700 ;
        RECT 54.000 170.200 54.800 170.400 ;
        RECT 56.000 170.200 56.600 171.600 ;
        RECT 72.200 170.400 72.800 177.000 ;
        RECT 78.000 175.800 78.800 179.800 ;
        RECT 82.400 176.200 84.000 179.800 ;
        RECT 78.000 175.200 80.200 175.800 ;
        RECT 81.200 175.400 82.800 175.600 ;
        RECT 79.400 175.000 80.200 175.200 ;
        RECT 80.800 174.800 82.800 175.400 ;
        RECT 80.800 174.400 81.400 174.800 ;
        RECT 78.000 173.800 81.400 174.400 ;
        RECT 78.000 173.600 79.600 173.800 ;
        RECT 82.000 173.400 82.800 174.200 ;
        RECT 82.000 172.800 82.600 173.400 ;
        RECT 80.000 172.200 82.600 172.800 ;
        RECT 83.400 172.800 84.000 176.200 ;
        RECT 87.600 175.800 88.400 179.800 ;
        RECT 84.600 174.800 85.400 175.600 ;
        RECT 86.000 175.200 88.400 175.800 ;
        RECT 90.800 175.200 91.600 179.800 ;
        RECT 94.000 175.200 94.800 179.800 ;
        RECT 97.200 175.200 98.000 179.800 ;
        RECT 100.400 175.200 101.200 179.800 ;
        RECT 86.000 175.000 86.800 175.200 ;
        RECT 84.800 174.400 85.400 174.800 ;
        RECT 89.200 174.400 91.600 175.200 ;
        RECT 92.600 174.400 94.800 175.200 ;
        RECT 95.800 174.400 98.000 175.200 ;
        RECT 99.400 174.400 101.200 175.200 ;
        RECT 84.800 173.600 85.600 174.400 ;
        RECT 86.800 173.600 88.400 174.400 ;
        RECT 83.400 172.400 84.400 172.800 ;
        RECT 83.400 172.200 85.200 172.400 ;
        RECT 80.000 172.000 80.800 172.200 ;
        RECT 83.800 171.600 85.200 172.200 ;
        RECT 89.200 171.600 90.000 174.400 ;
        RECT 92.600 173.800 93.400 174.400 ;
        RECT 95.800 173.800 96.600 174.400 ;
        RECT 99.400 173.800 100.200 174.400 ;
        RECT 90.800 173.000 93.400 173.800 ;
        RECT 94.200 173.000 96.600 173.800 ;
        RECT 97.600 173.000 100.200 173.800 ;
        RECT 92.600 171.600 93.400 173.000 ;
        RECT 95.800 171.600 96.600 173.000 ;
        RECT 99.400 171.600 100.200 173.000 ;
        RECT 103.600 173.800 104.400 179.800 ;
        RECT 110.000 176.600 110.800 179.800 ;
        RECT 111.600 177.000 112.400 179.800 ;
        RECT 113.200 177.000 114.000 179.800 ;
        RECT 114.800 177.000 115.600 179.800 ;
        RECT 118.000 177.000 118.800 179.800 ;
        RECT 121.200 177.000 122.000 179.800 ;
        RECT 122.800 177.000 123.600 179.800 ;
        RECT 124.400 177.000 125.200 179.800 ;
        RECT 126.000 177.000 126.800 179.800 ;
        RECT 108.200 175.800 110.800 176.600 ;
        RECT 127.600 176.600 128.400 179.800 ;
        RECT 114.200 175.800 118.800 176.400 ;
        RECT 108.200 175.200 109.000 175.800 ;
        RECT 106.000 174.400 109.000 175.200 ;
        RECT 103.600 173.000 112.400 173.800 ;
        RECT 114.200 173.400 115.000 175.800 ;
        RECT 118.000 175.600 118.800 175.800 ;
        RECT 119.600 175.600 121.200 176.400 ;
        RECT 124.200 175.600 125.200 176.400 ;
        RECT 127.600 175.800 130.000 176.600 ;
        RECT 116.400 173.600 117.200 175.200 ;
        RECT 118.000 174.800 118.800 175.000 ;
        RECT 118.000 174.200 122.400 174.800 ;
        RECT 121.600 174.000 122.400 174.200 ;
        RECT 82.200 171.400 83.000 171.600 ;
        RECT 79.600 170.800 83.000 171.400 ;
        RECT 54.000 169.600 55.400 170.200 ;
        RECT 56.000 169.600 57.000 170.200 ;
        RECT 72.200 169.800 75.600 170.400 ;
        RECT 79.600 170.200 80.200 170.800 ;
        RECT 83.800 170.200 84.400 171.600 ;
        RECT 89.200 170.800 91.600 171.600 ;
        RECT 92.600 170.800 94.800 171.600 ;
        RECT 95.800 170.800 98.000 171.600 ;
        RECT 99.400 170.800 101.200 171.600 ;
        RECT 49.200 167.700 51.600 168.300 ;
        RECT 49.200 167.600 50.000 167.700 ;
        RECT 50.800 162.200 51.600 167.700 ;
        RECT 54.800 168.400 55.400 169.600 ;
        RECT 54.800 167.600 55.600 168.400 ;
        RECT 56.200 162.200 57.000 169.600 ;
        RECT 74.800 169.600 75.600 169.800 ;
        RECT 78.000 169.600 80.200 170.200 ;
        RECT 65.400 168.800 69.000 169.400 ;
        RECT 65.400 168.200 66.000 168.800 ;
        RECT 65.200 162.200 66.000 168.200 ;
        RECT 68.400 168.200 69.000 168.800 ;
        RECT 70.200 169.000 73.800 169.200 ;
        RECT 74.800 169.000 75.400 169.600 ;
        RECT 70.200 168.600 74.000 169.000 ;
        RECT 70.200 168.200 70.800 168.600 ;
        RECT 68.400 162.800 69.200 168.200 ;
        RECT 70.000 163.400 70.800 168.200 ;
        RECT 71.600 162.800 72.400 168.000 ;
        RECT 73.200 163.000 74.000 168.600 ;
        RECT 74.800 163.400 75.600 169.000 ;
        RECT 68.400 162.200 72.400 162.800 ;
        RECT 73.400 162.800 74.000 163.000 ;
        RECT 76.400 163.000 77.200 169.000 ;
        RECT 76.400 162.800 77.000 163.000 ;
        RECT 73.400 162.200 77.000 162.800 ;
        RECT 78.000 162.200 78.800 169.600 ;
        RECT 79.400 169.400 80.200 169.600 ;
        RECT 82.400 169.600 84.400 170.200 ;
        RECT 86.000 169.600 88.400 170.200 ;
        RECT 82.400 162.200 84.000 169.600 ;
        RECT 86.000 169.400 86.800 169.600 ;
        RECT 87.600 162.200 88.400 169.600 ;
        RECT 90.800 162.200 91.600 170.800 ;
        RECT 94.000 162.200 94.800 170.800 ;
        RECT 97.200 162.200 98.000 170.800 ;
        RECT 100.400 162.200 101.200 170.800 ;
        RECT 103.600 167.400 104.400 173.000 ;
        RECT 113.000 172.600 115.000 173.400 ;
        RECT 118.800 172.600 122.000 173.400 ;
        RECT 124.400 172.800 125.200 175.600 ;
        RECT 129.200 175.200 130.000 175.800 ;
        RECT 129.200 174.600 131.000 175.200 ;
        RECT 130.200 173.400 131.000 174.600 ;
        RECT 134.000 174.600 134.800 179.800 ;
        RECT 135.600 176.000 136.400 179.800 ;
        RECT 135.600 175.200 136.600 176.000 ;
        RECT 142.000 175.200 142.800 179.800 ;
        RECT 143.600 175.800 144.400 179.800 ;
        RECT 148.000 176.200 149.600 179.800 ;
        RECT 143.600 175.200 145.800 175.800 ;
        RECT 146.800 175.400 148.400 175.600 ;
        RECT 134.000 174.000 135.200 174.600 ;
        RECT 130.200 172.600 134.000 173.400 ;
        RECT 105.000 172.000 105.800 172.200 ;
        RECT 110.000 172.000 110.800 172.400 ;
        RECT 127.600 172.000 128.400 172.600 ;
        RECT 134.600 172.000 135.200 174.000 ;
        RECT 105.000 171.400 128.400 172.000 ;
        RECT 134.400 171.400 135.200 172.000 ;
        RECT 134.400 169.600 135.000 171.400 ;
        RECT 135.800 170.800 136.600 175.200 ;
        RECT 140.600 174.600 142.800 175.200 ;
        RECT 145.000 175.000 145.800 175.200 ;
        RECT 146.400 174.800 148.400 175.400 ;
        RECT 140.600 171.600 141.200 174.600 ;
        RECT 146.400 174.400 147.000 174.800 ;
        RECT 143.600 173.800 147.000 174.400 ;
        RECT 143.600 173.600 145.200 173.800 ;
        RECT 147.600 173.400 148.400 174.200 ;
        RECT 142.000 171.600 142.800 173.200 ;
        RECT 147.600 172.800 148.200 173.400 ;
        RECT 145.600 172.200 148.200 172.800 ;
        RECT 149.000 172.800 149.600 176.200 ;
        RECT 153.200 175.800 154.000 179.800 ;
        RECT 150.200 174.800 151.000 175.600 ;
        RECT 151.600 175.200 154.000 175.800 ;
        RECT 159.600 175.600 160.400 177.200 ;
        RECT 151.600 175.000 152.400 175.200 ;
        RECT 150.400 174.400 151.000 174.800 ;
        RECT 150.400 173.600 151.200 174.400 ;
        RECT 152.400 174.300 154.000 174.400 ;
        RECT 161.200 174.300 162.000 179.800 ;
        RECT 163.400 178.400 164.200 179.800 ;
        RECT 163.400 177.600 165.200 178.400 ;
        RECT 163.400 176.400 164.200 177.600 ;
        RECT 163.400 175.800 165.200 176.400 ;
        RECT 152.400 173.700 162.000 174.300 ;
        RECT 152.400 173.600 154.000 173.700 ;
        RECT 149.000 172.400 150.000 172.800 ;
        RECT 149.000 172.200 150.800 172.400 ;
        RECT 145.600 172.000 146.400 172.200 ;
        RECT 149.400 171.600 150.800 172.200 ;
        RECT 140.000 170.800 141.200 171.600 ;
        RECT 147.800 171.400 148.600 171.600 ;
        RECT 113.200 169.400 114.000 169.600 ;
        RECT 108.600 169.000 114.000 169.400 ;
        RECT 107.800 168.800 114.000 169.000 ;
        RECT 115.000 169.000 123.600 169.600 ;
        RECT 105.200 168.000 106.800 168.800 ;
        RECT 107.800 168.200 109.200 168.800 ;
        RECT 115.000 168.200 115.600 169.000 ;
        RECT 122.800 168.800 123.600 169.000 ;
        RECT 126.000 169.000 135.000 169.600 ;
        RECT 126.000 168.800 126.800 169.000 ;
        RECT 106.200 167.600 106.800 168.000 ;
        RECT 109.800 167.600 115.600 168.200 ;
        RECT 116.200 167.600 118.800 168.400 ;
        RECT 103.600 166.800 105.600 167.400 ;
        RECT 106.200 166.800 110.400 167.600 ;
        RECT 105.000 166.200 105.600 166.800 ;
        RECT 105.000 165.600 106.000 166.200 ;
        RECT 105.200 162.200 106.000 165.600 ;
        RECT 108.400 162.200 109.200 166.800 ;
        RECT 111.600 162.200 112.400 165.000 ;
        RECT 113.200 162.200 114.000 165.000 ;
        RECT 114.800 162.200 115.600 167.000 ;
        RECT 118.000 162.200 118.800 167.000 ;
        RECT 121.200 162.200 122.000 168.400 ;
        RECT 129.200 167.600 131.800 168.400 ;
        RECT 124.400 166.800 128.600 167.600 ;
        RECT 122.800 162.200 123.600 165.000 ;
        RECT 124.400 162.200 125.200 165.000 ;
        RECT 126.000 162.200 126.800 165.000 ;
        RECT 129.200 162.200 130.000 167.600 ;
        RECT 134.400 167.400 135.000 169.000 ;
        RECT 132.400 166.800 135.000 167.400 ;
        RECT 135.600 170.000 136.600 170.800 ;
        RECT 140.600 170.200 141.200 170.800 ;
        RECT 145.200 170.800 148.600 171.400 ;
        RECT 145.200 170.200 145.800 170.800 ;
        RECT 149.400 170.200 150.000 171.600 ;
        RECT 132.400 162.200 133.200 166.800 ;
        RECT 135.600 162.200 136.400 170.000 ;
        RECT 140.600 169.600 142.800 170.200 ;
        RECT 142.000 162.200 142.800 169.600 ;
        RECT 143.600 169.600 145.800 170.200 ;
        RECT 143.600 162.200 144.400 169.600 ;
        RECT 145.000 169.400 145.800 169.600 ;
        RECT 148.000 169.600 150.000 170.200 ;
        RECT 151.600 169.600 154.000 170.200 ;
        RECT 148.000 168.400 149.600 169.600 ;
        RECT 151.600 169.400 152.400 169.600 ;
        RECT 146.800 167.600 149.600 168.400 ;
        RECT 148.000 162.200 149.600 167.600 ;
        RECT 153.200 162.200 154.000 169.600 ;
        RECT 161.200 162.200 162.000 173.700 ;
        RECT 162.800 168.800 163.600 170.400 ;
        RECT 164.400 162.200 165.200 175.800 ;
        RECT 167.600 175.800 168.400 179.800 ;
        RECT 172.000 176.200 173.600 179.800 ;
        RECT 167.600 175.200 170.000 175.800 ;
        RECT 166.000 173.600 166.800 175.200 ;
        RECT 169.200 175.000 170.000 175.200 ;
        RECT 170.600 174.800 171.400 175.600 ;
        RECT 170.600 174.400 171.200 174.800 ;
        RECT 167.600 173.600 169.200 174.400 ;
        RECT 170.400 173.600 171.200 174.400 ;
        RECT 172.000 172.800 172.600 176.200 ;
        RECT 177.200 175.800 178.000 179.800 ;
        RECT 181.400 176.400 182.200 179.800 ;
        RECT 173.200 175.400 174.800 175.600 ;
        RECT 173.200 174.800 175.200 175.400 ;
        RECT 175.800 175.200 178.000 175.800 ;
        RECT 180.400 175.800 182.200 176.400 ;
        RECT 185.200 177.800 186.000 179.800 ;
        RECT 175.800 175.000 176.600 175.200 ;
        RECT 174.600 174.400 175.200 174.800 ;
        RECT 173.200 173.400 174.000 174.200 ;
        RECT 174.600 173.800 178.000 174.400 ;
        RECT 176.400 173.600 178.000 173.800 ;
        RECT 178.800 173.600 179.600 175.200 ;
        RECT 171.600 172.400 172.600 172.800 ;
        RECT 170.800 172.200 172.600 172.400 ;
        RECT 173.400 172.800 174.000 173.400 ;
        RECT 173.400 172.200 176.000 172.800 ;
        RECT 170.800 171.600 172.200 172.200 ;
        RECT 175.200 172.000 176.000 172.200 ;
        RECT 177.300 172.300 177.900 173.600 ;
        RECT 180.400 172.300 181.200 175.800 ;
        RECT 185.200 174.400 185.800 177.800 ;
        RECT 186.800 176.300 187.600 177.200 ;
        RECT 188.400 176.300 189.200 179.800 ;
        RECT 186.800 175.700 189.200 176.300 ;
        RECT 186.800 175.600 187.600 175.700 ;
        RECT 185.200 174.300 186.000 174.400 ;
        RECT 186.800 174.300 187.600 174.400 ;
        RECT 185.200 173.700 187.600 174.300 ;
        RECT 185.200 173.600 186.000 173.700 ;
        RECT 186.800 173.600 187.600 173.700 ;
        RECT 183.600 172.300 184.400 172.400 ;
        RECT 177.300 171.700 184.400 172.300 ;
        RECT 171.600 170.200 172.200 171.600 ;
        RECT 173.000 171.400 173.800 171.600 ;
        RECT 173.000 170.800 176.400 171.400 ;
        RECT 175.800 170.200 176.400 170.800 ;
        RECT 167.600 169.600 170.000 170.200 ;
        RECT 171.600 169.600 173.600 170.200 ;
        RECT 167.600 162.200 168.400 169.600 ;
        RECT 169.200 169.400 170.000 169.600 ;
        RECT 172.000 164.400 173.600 169.600 ;
        RECT 175.800 169.600 178.000 170.200 ;
        RECT 175.800 169.400 176.600 169.600 ;
        RECT 170.800 163.600 173.600 164.400 ;
        RECT 172.000 162.200 173.600 163.600 ;
        RECT 177.200 162.200 178.000 169.600 ;
        RECT 180.400 162.200 181.200 171.700 ;
        RECT 183.600 170.800 184.400 171.700 ;
        RECT 182.000 168.800 182.800 170.400 ;
        RECT 185.200 170.200 185.800 173.600 ;
        RECT 184.200 169.400 186.000 170.200 ;
        RECT 184.200 162.200 185.000 169.400 ;
        RECT 188.400 162.200 189.200 175.700 ;
        RECT 190.000 175.600 190.800 177.200 ;
        RECT 191.600 175.800 192.400 179.800 ;
        RECT 196.000 178.400 197.600 179.800 ;
        RECT 194.800 177.600 197.600 178.400 ;
        RECT 196.000 176.200 197.600 177.600 ;
        RECT 191.600 175.200 194.200 175.800 ;
        RECT 193.400 175.000 194.200 175.200 ;
        RECT 194.800 174.800 196.400 175.600 ;
        RECT 191.600 174.200 193.200 174.400 ;
        RECT 197.000 174.200 197.600 176.200 ;
        RECT 201.200 175.800 202.000 179.800 ;
        RECT 203.400 178.400 204.200 179.800 ;
        RECT 202.800 177.600 204.200 178.400 ;
        RECT 203.400 176.800 204.200 177.600 ;
        RECT 198.200 174.800 199.000 175.600 ;
        RECT 199.600 175.200 202.000 175.800 ;
        RECT 202.800 175.800 204.200 176.800 ;
        RECT 207.600 175.800 208.400 179.800 ;
        RECT 199.600 175.000 200.400 175.200 ;
        RECT 191.600 174.000 193.800 174.200 ;
        RECT 191.600 173.600 196.000 174.000 ;
        RECT 193.200 173.400 196.000 173.600 ;
        RECT 195.200 173.200 196.000 173.400 ;
        RECT 196.600 173.600 197.600 174.200 ;
        RECT 198.400 174.400 199.000 174.800 ;
        RECT 198.400 173.600 199.200 174.400 ;
        RECT 200.400 173.600 202.000 174.400 ;
        RECT 196.600 172.400 197.200 173.600 ;
        RECT 193.800 172.200 194.600 172.400 ;
        RECT 193.800 171.600 195.400 172.200 ;
        RECT 196.400 171.600 197.200 172.400 ;
        RECT 194.600 171.400 195.400 171.600 ;
        RECT 196.600 170.200 197.200 171.600 ;
        RECT 202.800 172.400 203.400 175.800 ;
        RECT 207.600 175.600 208.200 175.800 ;
        RECT 206.400 175.200 208.200 175.600 ;
        RECT 204.000 175.000 208.200 175.200 ;
        RECT 209.200 175.200 210.000 179.800 ;
        RECT 214.000 175.200 214.800 179.800 ;
        RECT 204.000 174.600 207.000 175.000 ;
        RECT 209.200 174.600 211.400 175.200 ;
        RECT 214.000 174.600 216.200 175.200 ;
        RECT 204.000 174.400 204.800 174.600 ;
        RECT 202.800 171.600 203.600 172.400 ;
        RECT 202.800 170.200 203.400 171.600 ;
        RECT 204.200 171.000 204.800 174.400 ;
        RECT 205.600 173.800 206.400 174.000 ;
        RECT 205.600 173.200 206.600 173.800 ;
        RECT 206.000 172.400 206.600 173.200 ;
        RECT 206.000 171.600 206.800 172.400 ;
        RECT 207.600 172.300 208.400 174.400 ;
        RECT 209.200 172.300 210.000 173.200 ;
        RECT 207.600 171.700 210.000 172.300 ;
        RECT 209.200 171.600 210.000 171.700 ;
        RECT 210.800 171.600 211.400 174.600 ;
        RECT 214.000 171.600 214.800 173.200 ;
        RECT 215.600 171.600 216.200 174.600 ;
        RECT 204.200 170.400 206.600 171.000 ;
        RECT 191.600 169.600 194.200 170.200 ;
        RECT 191.600 162.200 192.400 169.600 ;
        RECT 193.400 169.400 194.200 169.600 ;
        RECT 196.000 162.200 197.600 170.200 ;
        RECT 199.600 169.600 202.000 170.200 ;
        RECT 199.600 169.400 200.400 169.600 ;
        RECT 201.200 162.200 202.000 169.600 ;
        RECT 202.800 162.200 203.600 170.200 ;
        RECT 206.000 166.200 206.600 170.400 ;
        RECT 210.800 170.800 212.000 171.600 ;
        RECT 215.600 170.800 216.800 171.600 ;
        RECT 210.800 170.200 211.400 170.800 ;
        RECT 215.600 170.200 216.200 170.800 ;
        RECT 209.200 169.600 211.400 170.200 ;
        RECT 214.000 169.600 216.200 170.200 ;
        RECT 206.000 162.200 206.800 166.200 ;
        RECT 209.200 162.200 210.000 169.600 ;
        RECT 214.000 162.200 214.800 169.600 ;
        RECT 4.400 152.400 5.200 159.800 ;
        RECT 9.200 152.400 10.000 159.800 ;
        RECT 3.000 151.800 5.200 152.400 ;
        RECT 7.800 151.800 10.000 152.400 ;
        RECT 3.000 151.200 3.600 151.800 ;
        RECT 7.800 151.200 8.400 151.800 ;
        RECT 2.400 150.400 3.600 151.200 ;
        RECT 7.200 150.400 8.400 151.200 ;
        RECT 3.000 147.400 3.600 150.400 ;
        RECT 4.400 148.800 5.200 150.400 ;
        RECT 7.800 147.400 8.400 150.400 ;
        RECT 9.200 148.800 10.000 150.400 ;
        RECT 12.400 150.300 13.200 159.800 ;
        RECT 15.600 152.300 16.400 159.800 ;
        RECT 18.800 155.800 19.600 159.800 ;
        RECT 19.000 155.600 19.600 155.800 ;
        RECT 22.000 155.800 22.800 159.800 ;
        RECT 22.000 155.600 22.600 155.800 ;
        RECT 19.000 155.000 22.600 155.600 ;
        RECT 20.400 152.800 21.200 154.400 ;
        RECT 22.000 152.400 22.600 155.000 ;
        RECT 17.200 152.300 18.000 152.400 ;
        RECT 15.600 151.700 18.000 152.300 ;
        RECT 14.000 150.300 14.800 150.400 ;
        RECT 12.400 149.700 14.800 150.300 ;
        RECT 3.000 146.800 5.200 147.400 ;
        RECT 7.800 146.800 10.000 147.400 ;
        RECT 4.400 142.200 5.200 146.800 ;
        RECT 9.200 142.200 10.000 146.800 ;
        RECT 10.800 144.800 11.600 146.400 ;
        RECT 12.400 142.200 13.200 149.700 ;
        RECT 14.000 149.600 14.800 149.700 ;
        RECT 14.000 144.800 14.800 146.400 ;
        RECT 15.600 142.200 16.400 151.700 ;
        RECT 17.200 150.800 18.000 151.700 ;
        RECT 22.000 151.600 22.800 152.400 ;
        RECT 18.800 149.600 20.400 150.400 ;
        RECT 22.000 148.400 22.600 151.600 ;
        RECT 21.000 148.300 22.600 148.400 ;
        RECT 23.600 148.300 24.400 148.400 ;
        RECT 21.000 148.200 24.400 148.300 ;
        RECT 20.800 147.700 24.400 148.200 ;
        RECT 20.800 144.400 21.600 147.700 ;
        RECT 23.600 146.800 24.400 147.700 ;
        RECT 25.200 146.200 26.000 159.800 ;
        RECT 29.200 153.600 30.000 154.400 ;
        RECT 26.800 151.600 27.600 153.200 ;
        RECT 29.200 152.400 29.800 153.600 ;
        RECT 30.600 152.400 31.400 159.800 ;
        RECT 28.400 151.800 29.800 152.400 ;
        RECT 30.400 151.800 31.400 152.400 ;
        RECT 28.400 151.600 29.200 151.800 ;
        RECT 26.900 150.300 27.500 151.600 ;
        RECT 30.400 150.300 31.000 151.800 ;
        RECT 34.800 151.600 35.600 153.200 ;
        RECT 26.900 149.700 31.000 150.300 ;
        RECT 30.400 148.400 31.000 149.700 ;
        RECT 31.600 150.300 32.400 150.400 ;
        RECT 34.900 150.300 35.500 151.600 ;
        RECT 31.600 149.700 35.500 150.300 ;
        RECT 31.600 148.800 32.400 149.700 ;
        RECT 28.400 147.600 31.000 148.400 ;
        RECT 33.200 148.300 34.000 148.400 ;
        RECT 34.800 148.300 35.600 148.400 ;
        RECT 33.200 148.200 35.600 148.300 ;
        RECT 32.400 147.700 35.600 148.200 ;
        RECT 32.400 147.600 34.000 147.700 ;
        RECT 34.800 147.600 35.600 147.700 ;
        RECT 28.600 146.200 29.200 147.600 ;
        RECT 32.400 147.200 33.200 147.600 ;
        RECT 30.200 146.200 33.800 146.600 ;
        RECT 36.400 146.200 37.200 159.800 ;
        RECT 41.200 156.400 42.000 159.800 ;
        RECT 41.000 155.800 42.000 156.400 ;
        RECT 41.000 155.200 41.600 155.800 ;
        RECT 44.400 155.200 45.200 159.800 ;
        RECT 47.600 157.000 48.400 159.800 ;
        RECT 49.200 157.000 50.000 159.800 ;
        RECT 39.600 154.600 41.600 155.200 ;
        RECT 39.600 149.000 40.400 154.600 ;
        RECT 42.200 154.400 46.400 155.200 ;
        RECT 50.800 155.000 51.600 159.800 ;
        RECT 54.000 155.000 54.800 159.800 ;
        RECT 42.200 154.000 42.800 154.400 ;
        RECT 41.200 153.200 42.800 154.000 ;
        RECT 45.800 153.800 51.600 154.400 ;
        RECT 43.800 153.200 45.200 153.800 ;
        RECT 43.800 153.000 50.000 153.200 ;
        RECT 44.600 152.600 50.000 153.000 ;
        RECT 49.200 152.400 50.000 152.600 ;
        RECT 51.000 153.000 51.600 153.800 ;
        RECT 52.200 153.600 54.800 154.400 ;
        RECT 57.200 153.600 58.000 159.800 ;
        RECT 58.800 157.000 59.600 159.800 ;
        RECT 60.400 157.000 61.200 159.800 ;
        RECT 62.000 157.000 62.800 159.800 ;
        RECT 60.400 154.400 64.600 155.200 ;
        RECT 65.200 154.400 66.000 159.800 ;
        RECT 68.400 155.200 69.200 159.800 ;
        RECT 68.400 154.600 71.000 155.200 ;
        RECT 65.200 153.600 67.800 154.400 ;
        RECT 58.800 153.000 59.600 153.200 ;
        RECT 51.000 152.400 59.600 153.000 ;
        RECT 62.000 153.000 62.800 153.200 ;
        RECT 70.400 153.000 71.000 154.600 ;
        RECT 62.000 152.400 71.000 153.000 ;
        RECT 42.800 151.800 43.600 152.400 ;
        RECT 46.000 151.800 47.000 152.000 ;
        RECT 42.800 151.200 69.800 151.800 ;
        RECT 69.000 151.000 69.800 151.200 ;
        RECT 70.400 150.600 71.000 152.400 ;
        RECT 71.600 152.000 72.400 159.800 ;
        RECT 81.200 156.400 82.000 159.800 ;
        RECT 81.000 155.800 82.000 156.400 ;
        RECT 81.000 155.200 81.600 155.800 ;
        RECT 84.400 155.200 85.200 159.800 ;
        RECT 87.600 157.000 88.400 159.800 ;
        RECT 89.200 157.000 90.000 159.800 ;
        RECT 79.600 154.600 81.600 155.200 ;
        RECT 71.600 151.200 72.600 152.000 ;
        RECT 70.400 150.000 71.200 150.600 ;
        RECT 38.000 146.800 38.800 148.400 ;
        RECT 39.600 148.200 48.400 149.000 ;
        RECT 49.000 148.600 51.000 149.400 ;
        RECT 54.800 148.600 58.000 149.400 ;
        RECT 25.200 145.600 27.000 146.200 ;
        RECT 20.400 143.600 21.600 144.400 ;
        RECT 20.800 142.200 21.600 143.600 ;
        RECT 26.200 142.200 27.000 145.600 ;
        RECT 28.400 142.200 29.200 146.200 ;
        RECT 30.000 146.000 34.000 146.200 ;
        RECT 30.000 142.200 30.800 146.000 ;
        RECT 33.200 142.200 34.000 146.000 ;
        RECT 35.400 145.600 37.200 146.200 ;
        RECT 35.400 142.200 36.200 145.600 ;
        RECT 39.600 142.200 40.400 148.200 ;
        RECT 42.000 146.800 45.000 147.600 ;
        RECT 44.200 146.200 45.000 146.800 ;
        RECT 50.200 146.200 51.000 148.600 ;
        RECT 52.400 146.800 53.200 148.400 ;
        RECT 57.600 147.800 58.400 148.000 ;
        RECT 54.000 147.200 58.400 147.800 ;
        RECT 54.000 147.000 54.800 147.200 ;
        RECT 60.400 146.400 61.200 149.200 ;
        RECT 66.200 148.600 70.000 149.400 ;
        RECT 66.200 147.400 67.000 148.600 ;
        RECT 70.600 148.000 71.200 150.000 ;
        RECT 54.000 146.200 54.800 146.400 ;
        RECT 44.200 145.400 46.800 146.200 ;
        RECT 50.200 145.600 54.800 146.200 ;
        RECT 55.600 145.600 57.200 146.400 ;
        RECT 60.200 145.600 61.200 146.400 ;
        RECT 65.200 146.800 67.000 147.400 ;
        RECT 70.000 147.400 71.200 148.000 ;
        RECT 65.200 146.200 66.000 146.800 ;
        RECT 46.000 142.200 46.800 145.400 ;
        RECT 63.600 145.400 66.000 146.200 ;
        RECT 47.600 142.200 48.400 145.000 ;
        RECT 49.200 142.200 50.000 145.000 ;
        RECT 50.800 142.200 51.600 145.000 ;
        RECT 54.000 142.200 54.800 145.000 ;
        RECT 57.200 142.200 58.000 145.000 ;
        RECT 58.800 142.200 59.600 145.000 ;
        RECT 60.400 142.200 61.200 145.000 ;
        RECT 62.000 142.200 62.800 145.000 ;
        RECT 63.600 142.200 64.400 145.400 ;
        RECT 70.000 142.200 70.800 147.400 ;
        RECT 71.800 146.800 72.600 151.200 ;
        RECT 71.600 146.000 72.600 146.800 ;
        RECT 79.600 149.000 80.400 154.600 ;
        RECT 82.200 154.400 86.400 155.200 ;
        RECT 90.800 155.000 91.600 159.800 ;
        RECT 94.000 155.000 94.800 159.800 ;
        RECT 82.200 154.000 82.800 154.400 ;
        RECT 81.200 153.200 82.800 154.000 ;
        RECT 85.800 153.800 91.600 154.400 ;
        RECT 83.800 153.200 85.200 153.800 ;
        RECT 83.800 153.000 90.000 153.200 ;
        RECT 84.600 152.600 90.000 153.000 ;
        RECT 89.200 152.400 90.000 152.600 ;
        RECT 91.000 153.000 91.600 153.800 ;
        RECT 92.200 153.600 94.800 154.400 ;
        RECT 97.200 153.600 98.000 159.800 ;
        RECT 98.800 157.000 99.600 159.800 ;
        RECT 100.400 157.000 101.200 159.800 ;
        RECT 102.000 157.000 102.800 159.800 ;
        RECT 100.400 154.400 104.600 155.200 ;
        RECT 105.200 154.400 106.000 159.800 ;
        RECT 108.400 155.200 109.200 159.800 ;
        RECT 108.400 154.600 111.000 155.200 ;
        RECT 105.200 153.600 107.800 154.400 ;
        RECT 98.800 153.000 99.600 153.200 ;
        RECT 91.000 152.400 99.600 153.000 ;
        RECT 102.000 153.000 102.800 153.200 ;
        RECT 110.400 153.000 111.000 154.600 ;
        RECT 102.000 152.400 111.000 153.000 ;
        RECT 82.800 151.800 83.600 152.400 ;
        RECT 86.000 151.800 87.000 152.000 ;
        RECT 82.800 151.200 109.800 151.800 ;
        RECT 109.000 151.000 109.800 151.200 ;
        RECT 110.400 150.600 111.000 152.400 ;
        RECT 111.600 152.000 112.400 159.800 ;
        RECT 111.600 151.200 112.600 152.000 ;
        RECT 110.400 150.000 111.200 150.600 ;
        RECT 79.600 148.200 88.400 149.000 ;
        RECT 89.000 148.600 91.000 149.400 ;
        RECT 94.800 148.600 98.000 149.400 ;
        RECT 71.600 142.200 72.400 146.000 ;
        RECT 79.600 142.200 80.400 148.200 ;
        RECT 82.000 146.800 85.000 147.600 ;
        RECT 84.200 146.200 85.000 146.800 ;
        RECT 90.200 146.200 91.000 148.600 ;
        RECT 92.400 146.800 93.200 148.400 ;
        RECT 97.600 147.800 98.400 148.000 ;
        RECT 94.000 147.200 98.400 147.800 ;
        RECT 94.000 147.000 94.800 147.200 ;
        RECT 100.400 146.400 101.200 149.200 ;
        RECT 106.200 148.600 110.000 149.400 ;
        RECT 106.200 147.400 107.000 148.600 ;
        RECT 110.600 148.000 111.200 150.000 ;
        RECT 94.000 146.200 94.800 146.400 ;
        RECT 84.200 145.400 86.800 146.200 ;
        RECT 90.200 145.600 94.800 146.200 ;
        RECT 95.600 145.600 97.200 146.400 ;
        RECT 100.200 145.600 101.200 146.400 ;
        RECT 105.200 146.800 107.000 147.400 ;
        RECT 110.000 147.400 111.200 148.000 ;
        RECT 105.200 146.200 106.000 146.800 ;
        RECT 86.000 142.200 86.800 145.400 ;
        RECT 103.600 145.400 106.000 146.200 ;
        RECT 87.600 142.200 88.400 145.000 ;
        RECT 89.200 142.200 90.000 145.000 ;
        RECT 90.800 142.200 91.600 145.000 ;
        RECT 94.000 142.200 94.800 145.000 ;
        RECT 97.200 142.200 98.000 145.000 ;
        RECT 98.800 142.200 99.600 145.000 ;
        RECT 100.400 142.200 101.200 145.000 ;
        RECT 102.000 142.200 102.800 145.000 ;
        RECT 103.600 142.200 104.400 145.400 ;
        RECT 110.000 142.200 110.800 147.400 ;
        RECT 111.800 146.800 112.600 151.200 ;
        RECT 116.400 151.200 117.200 159.800 ;
        RECT 119.600 151.200 120.400 159.800 ;
        RECT 122.800 151.200 123.600 159.800 ;
        RECT 126.000 151.200 126.800 159.800 ;
        RECT 130.800 156.400 131.600 159.800 ;
        RECT 130.600 155.800 131.600 156.400 ;
        RECT 130.600 155.200 131.200 155.800 ;
        RECT 134.000 155.200 134.800 159.800 ;
        RECT 137.200 157.000 138.000 159.800 ;
        RECT 138.800 157.000 139.600 159.800 ;
        RECT 129.200 154.600 131.200 155.200 ;
        RECT 116.400 150.400 118.200 151.200 ;
        RECT 119.600 150.400 121.800 151.200 ;
        RECT 122.800 150.400 125.000 151.200 ;
        RECT 126.000 150.400 128.400 151.200 ;
        RECT 117.400 149.000 118.200 150.400 ;
        RECT 121.000 149.000 121.800 150.400 ;
        RECT 124.200 149.000 125.000 150.400 ;
        RECT 117.400 148.200 120.000 149.000 ;
        RECT 121.000 148.200 123.400 149.000 ;
        RECT 124.200 148.200 126.800 149.000 ;
        RECT 117.400 147.600 118.200 148.200 ;
        RECT 121.000 147.600 121.800 148.200 ;
        RECT 124.200 147.600 125.000 148.200 ;
        RECT 127.600 147.600 128.400 150.400 ;
        RECT 111.600 146.000 112.600 146.800 ;
        RECT 116.400 146.800 118.200 147.600 ;
        RECT 119.600 146.800 121.800 147.600 ;
        RECT 122.800 146.800 125.000 147.600 ;
        RECT 126.000 146.800 128.400 147.600 ;
        RECT 129.200 149.000 130.000 154.600 ;
        RECT 131.800 154.400 136.000 155.200 ;
        RECT 140.400 155.000 141.200 159.800 ;
        RECT 143.600 155.000 144.400 159.800 ;
        RECT 131.800 154.000 132.400 154.400 ;
        RECT 130.800 153.200 132.400 154.000 ;
        RECT 135.400 153.800 141.200 154.400 ;
        RECT 133.400 153.200 134.800 153.800 ;
        RECT 133.400 153.000 139.600 153.200 ;
        RECT 134.200 152.600 139.600 153.000 ;
        RECT 138.800 152.400 139.600 152.600 ;
        RECT 140.600 153.000 141.200 153.800 ;
        RECT 141.800 153.600 144.400 154.400 ;
        RECT 146.800 153.600 147.600 159.800 ;
        RECT 148.400 157.000 149.200 159.800 ;
        RECT 150.000 157.000 150.800 159.800 ;
        RECT 151.600 157.000 152.400 159.800 ;
        RECT 150.000 154.400 154.200 155.200 ;
        RECT 154.800 154.400 155.600 159.800 ;
        RECT 158.000 155.200 158.800 159.800 ;
        RECT 158.000 154.600 160.600 155.200 ;
        RECT 154.800 153.600 157.400 154.400 ;
        RECT 148.400 153.000 149.200 153.200 ;
        RECT 140.600 152.400 149.200 153.000 ;
        RECT 151.600 153.000 152.400 153.200 ;
        RECT 160.000 153.000 160.600 154.600 ;
        RECT 151.600 152.400 160.600 153.000 ;
        RECT 160.000 150.600 160.600 152.400 ;
        RECT 161.200 152.000 162.000 159.800 ;
        RECT 162.800 154.300 163.600 154.400 ;
        RECT 162.800 153.700 170.000 154.300 ;
        RECT 162.800 153.600 163.600 153.700 ;
        RECT 161.200 151.200 162.200 152.000 ;
        RECT 169.200 151.600 170.000 153.700 ;
        RECT 130.600 150.000 154.000 150.600 ;
        RECT 160.000 150.000 160.800 150.600 ;
        RECT 130.600 149.800 131.400 150.000 ;
        RECT 132.400 149.600 133.200 150.000 ;
        RECT 135.600 149.600 136.400 150.000 ;
        RECT 153.200 149.400 154.000 150.000 ;
        RECT 129.200 148.200 138.000 149.000 ;
        RECT 138.600 148.600 140.600 149.400 ;
        RECT 144.400 148.600 147.600 149.400 ;
        RECT 111.600 142.200 112.400 146.000 ;
        RECT 116.400 142.200 117.200 146.800 ;
        RECT 119.600 142.200 120.400 146.800 ;
        RECT 122.800 142.200 123.600 146.800 ;
        RECT 126.000 142.200 126.800 146.800 ;
        RECT 129.200 142.200 130.000 148.200 ;
        RECT 131.600 146.800 134.600 147.600 ;
        RECT 133.800 146.200 134.600 146.800 ;
        RECT 139.800 146.200 140.600 148.600 ;
        RECT 142.000 146.800 142.800 148.400 ;
        RECT 147.200 147.800 148.000 148.000 ;
        RECT 143.600 147.200 148.000 147.800 ;
        RECT 143.600 147.000 144.400 147.200 ;
        RECT 150.000 146.400 150.800 149.200 ;
        RECT 155.800 148.600 159.600 149.400 ;
        RECT 155.800 147.400 156.600 148.600 ;
        RECT 160.200 148.000 160.800 150.000 ;
        RECT 143.600 146.200 144.400 146.400 ;
        RECT 133.800 145.400 136.400 146.200 ;
        RECT 139.800 145.600 144.400 146.200 ;
        RECT 145.200 145.600 146.800 146.400 ;
        RECT 149.800 145.600 150.800 146.400 ;
        RECT 154.800 146.800 156.600 147.400 ;
        RECT 159.600 147.400 160.800 148.000 ;
        RECT 154.800 146.200 155.600 146.800 ;
        RECT 135.600 142.200 136.400 145.400 ;
        RECT 153.200 145.400 155.600 146.200 ;
        RECT 137.200 142.200 138.000 145.000 ;
        RECT 138.800 142.200 139.600 145.000 ;
        RECT 140.400 142.200 141.200 145.000 ;
        RECT 143.600 142.200 144.400 145.000 ;
        RECT 146.800 142.200 147.600 145.000 ;
        RECT 148.400 142.200 149.200 145.000 ;
        RECT 150.000 142.200 150.800 145.000 ;
        RECT 151.600 142.200 152.400 145.000 ;
        RECT 153.200 142.200 154.000 145.400 ;
        RECT 159.600 142.200 160.400 147.400 ;
        RECT 161.400 146.800 162.200 151.200 ;
        RECT 161.200 146.000 162.200 146.800 ;
        RECT 170.800 146.200 171.600 159.800 ;
        RECT 175.600 156.400 176.400 159.800 ;
        RECT 175.400 155.800 176.400 156.400 ;
        RECT 175.400 155.200 176.000 155.800 ;
        RECT 178.800 155.200 179.600 159.800 ;
        RECT 182.000 157.000 182.800 159.800 ;
        RECT 183.600 157.000 184.400 159.800 ;
        RECT 174.000 154.600 176.000 155.200 ;
        RECT 174.000 149.000 174.800 154.600 ;
        RECT 176.600 154.400 180.800 155.200 ;
        RECT 185.200 155.000 186.000 159.800 ;
        RECT 188.400 155.000 189.200 159.800 ;
        RECT 176.600 154.000 177.200 154.400 ;
        RECT 175.600 153.200 177.200 154.000 ;
        RECT 180.200 153.800 186.000 154.400 ;
        RECT 178.200 153.200 179.600 153.800 ;
        RECT 178.200 153.000 184.400 153.200 ;
        RECT 179.000 152.600 184.400 153.000 ;
        RECT 183.600 152.400 184.400 152.600 ;
        RECT 185.400 153.000 186.000 153.800 ;
        RECT 186.600 153.600 189.200 154.400 ;
        RECT 191.600 153.600 192.400 159.800 ;
        RECT 193.200 157.000 194.000 159.800 ;
        RECT 194.800 157.000 195.600 159.800 ;
        RECT 196.400 157.000 197.200 159.800 ;
        RECT 194.800 154.400 199.000 155.200 ;
        RECT 199.600 154.400 200.400 159.800 ;
        RECT 202.800 155.200 203.600 159.800 ;
        RECT 202.800 154.600 205.400 155.200 ;
        RECT 199.600 153.600 202.200 154.400 ;
        RECT 193.200 153.000 194.000 153.200 ;
        RECT 185.400 152.400 194.000 153.000 ;
        RECT 196.400 153.000 197.200 153.200 ;
        RECT 204.800 153.000 205.400 154.600 ;
        RECT 196.400 152.400 205.400 153.000 ;
        RECT 204.800 150.600 205.400 152.400 ;
        RECT 206.000 152.000 206.800 159.800 ;
        RECT 209.200 152.400 210.000 159.800 ;
        RECT 214.000 152.400 214.800 159.800 ;
        RECT 206.000 151.200 207.000 152.000 ;
        RECT 209.200 151.800 211.400 152.400 ;
        RECT 214.000 151.800 216.200 152.400 ;
        RECT 175.400 150.000 198.800 150.600 ;
        RECT 204.800 150.000 205.600 150.600 ;
        RECT 175.400 149.800 176.200 150.000 ;
        RECT 177.200 149.600 178.000 150.000 ;
        RECT 180.400 149.600 181.200 150.000 ;
        RECT 198.000 149.400 198.800 150.000 ;
        RECT 172.400 146.800 173.200 148.400 ;
        RECT 174.000 148.200 182.800 149.000 ;
        RECT 183.400 148.600 185.400 149.400 ;
        RECT 189.200 148.600 192.400 149.400 ;
        RECT 161.200 142.200 162.000 146.000 ;
        RECT 169.800 145.600 171.600 146.200 ;
        RECT 169.800 144.400 170.600 145.600 ;
        RECT 169.800 143.600 171.600 144.400 ;
        RECT 169.800 142.200 170.600 143.600 ;
        RECT 174.000 142.200 174.800 148.200 ;
        RECT 176.400 146.800 179.400 147.600 ;
        RECT 178.600 146.200 179.400 146.800 ;
        RECT 184.600 146.200 185.400 148.600 ;
        RECT 186.800 146.800 187.600 148.400 ;
        RECT 192.000 147.800 192.800 148.000 ;
        RECT 188.400 147.200 192.800 147.800 ;
        RECT 188.400 147.000 189.200 147.200 ;
        RECT 194.800 146.400 195.600 149.200 ;
        RECT 200.600 148.600 204.400 149.400 ;
        RECT 200.600 147.400 201.400 148.600 ;
        RECT 205.000 148.000 205.600 150.000 ;
        RECT 188.400 146.200 189.200 146.400 ;
        RECT 178.600 145.400 181.200 146.200 ;
        RECT 184.600 145.600 189.200 146.200 ;
        RECT 190.000 145.600 191.600 146.400 ;
        RECT 194.600 145.600 195.600 146.400 ;
        RECT 199.600 146.800 201.400 147.400 ;
        RECT 204.400 147.400 205.600 148.000 ;
        RECT 206.200 150.300 207.000 151.200 ;
        RECT 210.800 151.200 211.400 151.800 ;
        RECT 215.600 151.200 216.200 151.800 ;
        RECT 210.800 150.400 212.000 151.200 ;
        RECT 215.600 150.400 216.800 151.200 ;
        RECT 209.200 150.300 210.000 150.400 ;
        RECT 206.200 149.700 210.000 150.300 ;
        RECT 199.600 146.200 200.400 146.800 ;
        RECT 180.400 142.200 181.200 145.400 ;
        RECT 198.000 145.400 200.400 146.200 ;
        RECT 182.000 142.200 182.800 145.000 ;
        RECT 183.600 142.200 184.400 145.000 ;
        RECT 185.200 142.200 186.000 145.000 ;
        RECT 188.400 142.200 189.200 145.000 ;
        RECT 191.600 142.200 192.400 145.000 ;
        RECT 193.200 142.200 194.000 145.000 ;
        RECT 194.800 142.200 195.600 145.000 ;
        RECT 196.400 142.200 197.200 145.000 ;
        RECT 198.000 142.200 198.800 145.400 ;
        RECT 204.400 142.200 205.200 147.400 ;
        RECT 206.200 146.800 207.000 149.700 ;
        RECT 209.200 148.800 210.000 149.700 ;
        RECT 210.800 147.400 211.400 150.400 ;
        RECT 214.000 148.800 214.800 150.400 ;
        RECT 215.600 147.400 216.200 150.400 ;
        RECT 206.000 146.000 207.000 146.800 ;
        RECT 209.200 146.800 211.400 147.400 ;
        RECT 214.000 146.800 216.200 147.400 ;
        RECT 206.000 142.200 206.800 146.000 ;
        RECT 209.200 142.200 210.000 146.800 ;
        RECT 214.000 142.200 214.800 146.800 ;
        RECT 2.800 136.000 3.600 139.800 ;
        RECT 2.600 135.200 3.600 136.000 ;
        RECT 2.600 130.800 3.400 135.200 ;
        RECT 4.400 134.600 5.200 139.800 ;
        RECT 10.800 136.600 11.600 139.800 ;
        RECT 12.400 137.000 13.200 139.800 ;
        RECT 14.000 137.000 14.800 139.800 ;
        RECT 15.600 137.000 16.400 139.800 ;
        RECT 17.200 137.000 18.000 139.800 ;
        RECT 20.400 137.000 21.200 139.800 ;
        RECT 23.600 137.000 24.400 139.800 ;
        RECT 25.200 137.000 26.000 139.800 ;
        RECT 26.800 137.000 27.600 139.800 ;
        RECT 9.200 135.800 11.600 136.600 ;
        RECT 28.400 136.600 29.200 139.800 ;
        RECT 9.200 135.200 10.000 135.800 ;
        RECT 4.000 134.000 5.200 134.600 ;
        RECT 8.200 134.600 10.000 135.200 ;
        RECT 14.000 135.600 15.000 136.400 ;
        RECT 18.000 135.600 19.600 136.400 ;
        RECT 20.400 135.800 25.000 136.400 ;
        RECT 28.400 135.800 31.000 136.600 ;
        RECT 20.400 135.600 21.200 135.800 ;
        RECT 4.000 132.000 4.600 134.000 ;
        RECT 8.200 133.400 9.000 134.600 ;
        RECT 5.200 132.600 9.000 133.400 ;
        RECT 14.000 132.800 14.800 135.600 ;
        RECT 20.400 134.800 21.200 135.000 ;
        RECT 16.800 134.200 21.200 134.800 ;
        RECT 16.800 134.000 17.600 134.200 ;
        RECT 22.000 133.600 22.800 135.200 ;
        RECT 24.200 133.400 25.000 135.800 ;
        RECT 30.200 135.200 31.000 135.800 ;
        RECT 30.200 134.400 33.200 135.200 ;
        RECT 34.800 133.800 35.600 139.800 ;
        RECT 39.600 138.400 40.400 139.800 ;
        RECT 39.600 137.800 40.600 138.400 ;
        RECT 40.000 137.600 40.600 137.800 ;
        RECT 42.800 137.800 43.600 139.800 ;
        RECT 42.800 137.600 44.000 137.800 ;
        RECT 40.000 137.000 44.000 137.600 ;
        RECT 36.400 136.300 37.200 136.400 ;
        RECT 38.000 136.300 39.800 136.400 ;
        RECT 36.400 135.700 39.800 136.300 ;
        RECT 36.400 135.600 37.200 135.700 ;
        RECT 38.000 135.600 39.800 135.700 ;
        RECT 17.200 132.600 20.400 133.400 ;
        RECT 24.200 132.600 26.200 133.400 ;
        RECT 26.800 133.000 35.600 133.800 ;
        RECT 38.000 134.300 38.800 134.400 ;
        RECT 39.600 134.300 41.200 134.400 ;
        RECT 38.000 133.700 41.200 134.300 ;
        RECT 38.000 133.600 38.800 133.700 ;
        RECT 39.600 133.600 41.200 133.700 ;
        RECT 10.800 132.000 11.600 132.600 ;
        RECT 28.400 132.000 29.200 132.400 ;
        RECT 31.600 132.000 32.400 132.400 ;
        RECT 33.400 132.000 34.200 132.200 ;
        RECT 4.000 131.400 4.800 132.000 ;
        RECT 10.800 131.400 34.200 132.000 ;
        RECT 2.600 130.000 3.600 130.800 ;
        RECT 2.800 122.200 3.600 130.000 ;
        RECT 4.200 129.600 4.800 131.400 ;
        RECT 4.200 129.000 13.200 129.600 ;
        RECT 4.200 127.400 4.800 129.000 ;
        RECT 12.400 128.800 13.200 129.000 ;
        RECT 15.600 129.000 24.200 129.600 ;
        RECT 15.600 128.800 16.400 129.000 ;
        RECT 7.400 127.600 10.000 128.400 ;
        RECT 4.200 126.800 6.800 127.400 ;
        RECT 6.000 122.200 6.800 126.800 ;
        RECT 9.200 122.200 10.000 127.600 ;
        RECT 10.600 126.800 14.800 127.600 ;
        RECT 12.400 122.200 13.200 125.000 ;
        RECT 14.000 122.200 14.800 125.000 ;
        RECT 15.600 122.200 16.400 125.000 ;
        RECT 17.200 122.200 18.000 128.400 ;
        RECT 20.400 127.600 23.000 128.400 ;
        RECT 23.600 128.200 24.200 129.000 ;
        RECT 25.200 129.400 26.000 129.600 ;
        RECT 25.200 129.000 30.600 129.400 ;
        RECT 25.200 128.800 31.400 129.000 ;
        RECT 30.000 128.200 31.400 128.800 ;
        RECT 23.600 127.600 29.400 128.200 ;
        RECT 32.400 128.000 34.000 128.800 ;
        RECT 32.400 127.600 33.000 128.000 ;
        RECT 20.400 122.200 21.200 127.000 ;
        RECT 23.600 122.200 24.400 127.000 ;
        RECT 28.800 126.800 33.000 127.600 ;
        RECT 34.800 127.400 35.600 133.000 ;
        RECT 41.200 131.600 42.800 132.400 ;
        RECT 43.400 130.600 44.000 137.000 ;
        RECT 49.200 135.800 50.000 139.800 ;
        RECT 53.600 136.200 55.200 139.800 ;
        RECT 49.200 135.200 51.400 135.800 ;
        RECT 52.400 135.400 54.000 135.600 ;
        RECT 50.600 135.000 51.400 135.200 ;
        RECT 52.000 134.800 54.000 135.400 ;
        RECT 52.000 134.400 52.600 134.800 ;
        RECT 49.200 133.800 52.600 134.400 ;
        RECT 49.200 133.600 50.800 133.800 ;
        RECT 53.200 133.400 54.000 134.200 ;
        RECT 53.200 132.800 53.800 133.400 ;
        RECT 51.200 132.200 53.800 132.800 ;
        RECT 54.600 132.800 55.200 136.200 ;
        RECT 58.800 135.800 59.600 139.800 ;
        RECT 66.800 136.000 67.600 139.800 ;
        RECT 55.800 134.800 56.600 135.600 ;
        RECT 57.200 135.200 59.600 135.800 ;
        RECT 66.600 135.200 67.600 136.000 ;
        RECT 57.200 135.000 58.000 135.200 ;
        RECT 56.000 134.400 56.600 134.800 ;
        RECT 56.000 133.600 56.800 134.400 ;
        RECT 58.000 134.300 59.600 134.400 ;
        RECT 66.600 134.300 67.400 135.200 ;
        RECT 68.400 134.600 69.200 139.800 ;
        RECT 74.800 136.600 75.600 139.800 ;
        RECT 76.400 137.000 77.200 139.800 ;
        RECT 78.000 137.000 78.800 139.800 ;
        RECT 79.600 137.000 80.400 139.800 ;
        RECT 81.200 137.000 82.000 139.800 ;
        RECT 84.400 137.000 85.200 139.800 ;
        RECT 87.600 137.000 88.400 139.800 ;
        RECT 89.200 137.000 90.000 139.800 ;
        RECT 90.800 137.000 91.600 139.800 ;
        RECT 73.200 135.800 75.600 136.600 ;
        RECT 92.400 136.600 93.200 139.800 ;
        RECT 73.200 135.200 74.000 135.800 ;
        RECT 58.000 133.700 67.400 134.300 ;
        RECT 58.000 133.600 59.600 133.700 ;
        RECT 54.600 132.400 55.600 132.800 ;
        RECT 54.600 132.200 56.400 132.400 ;
        RECT 51.200 132.000 52.000 132.200 ;
        RECT 55.000 131.600 56.400 132.200 ;
        RECT 53.400 131.400 54.200 131.600 ;
        RECT 50.800 130.800 54.200 131.400 ;
        RECT 43.400 130.400 45.200 130.600 ;
        RECT 43.400 129.800 46.800 130.400 ;
        RECT 50.800 130.200 51.400 130.800 ;
        RECT 55.000 130.200 55.600 131.600 ;
        RECT 66.600 130.800 67.400 133.700 ;
        RECT 68.000 134.000 69.200 134.600 ;
        RECT 72.200 134.600 74.000 135.200 ;
        RECT 78.000 135.600 79.000 136.400 ;
        RECT 82.000 135.600 83.600 136.400 ;
        RECT 84.400 135.800 89.000 136.400 ;
        RECT 92.400 135.800 95.000 136.600 ;
        RECT 84.400 135.600 85.200 135.800 ;
        RECT 68.000 132.000 68.600 134.000 ;
        RECT 72.200 133.400 73.000 134.600 ;
        RECT 69.200 132.600 73.000 133.400 ;
        RECT 78.000 132.800 78.800 135.600 ;
        RECT 84.400 134.800 85.200 135.000 ;
        RECT 80.800 134.200 85.200 134.800 ;
        RECT 80.800 134.000 81.600 134.200 ;
        RECT 86.000 133.600 86.800 135.200 ;
        RECT 88.200 133.400 89.000 135.800 ;
        RECT 94.200 135.200 95.000 135.800 ;
        RECT 94.200 134.400 97.200 135.200 ;
        RECT 98.800 133.800 99.600 139.800 ;
        RECT 100.400 135.800 101.200 139.800 ;
        RECT 104.800 136.200 106.400 139.800 ;
        RECT 100.400 135.200 102.800 135.800 ;
        RECT 102.000 135.000 102.800 135.200 ;
        RECT 103.400 134.800 104.200 135.600 ;
        RECT 103.400 134.400 104.000 134.800 ;
        RECT 81.200 132.600 84.400 133.400 ;
        RECT 88.200 132.600 90.200 133.400 ;
        RECT 90.800 133.000 99.600 133.800 ;
        RECT 100.400 133.600 102.000 134.400 ;
        RECT 103.200 133.600 104.000 134.400 ;
        RECT 68.000 131.400 68.800 132.000 ;
        RECT 46.000 129.600 46.800 129.800 ;
        RECT 49.200 129.600 51.400 130.200 ;
        RECT 36.600 128.800 40.200 129.400 ;
        RECT 36.600 128.200 37.200 128.800 ;
        RECT 33.600 126.800 35.600 127.400 ;
        RECT 25.200 122.200 26.000 125.000 ;
        RECT 26.800 122.200 27.600 125.000 ;
        RECT 30.000 122.200 30.800 126.800 ;
        RECT 33.600 126.200 34.200 126.800 ;
        RECT 33.200 125.600 34.200 126.200 ;
        RECT 33.200 122.200 34.000 125.600 ;
        RECT 36.400 122.200 37.200 128.200 ;
        RECT 39.600 128.200 40.200 128.800 ;
        RECT 41.400 129.000 45.000 129.200 ;
        RECT 46.000 129.000 46.600 129.600 ;
        RECT 41.400 128.600 45.200 129.000 ;
        RECT 41.400 128.200 42.000 128.600 ;
        RECT 39.600 122.800 40.400 128.200 ;
        RECT 41.200 123.400 42.000 128.200 ;
        RECT 42.800 122.800 43.600 128.000 ;
        RECT 44.400 123.000 45.200 128.600 ;
        RECT 46.000 123.400 46.800 129.000 ;
        RECT 39.600 122.200 43.600 122.800 ;
        RECT 44.600 122.800 45.200 123.000 ;
        RECT 47.600 123.000 48.400 129.000 ;
        RECT 47.600 122.800 48.200 123.000 ;
        RECT 44.600 122.200 48.200 122.800 ;
        RECT 49.200 122.200 50.000 129.600 ;
        RECT 50.600 129.400 51.400 129.600 ;
        RECT 53.600 129.600 55.600 130.200 ;
        RECT 57.200 129.600 59.600 130.200 ;
        RECT 66.600 130.000 67.600 130.800 ;
        RECT 53.600 122.200 55.200 129.600 ;
        RECT 57.200 129.400 58.000 129.600 ;
        RECT 58.800 122.200 59.600 129.600 ;
        RECT 66.800 122.200 67.600 130.000 ;
        RECT 68.200 129.600 68.800 131.400 ;
        RECT 69.400 130.800 70.200 131.000 ;
        RECT 69.400 130.200 96.400 130.800 ;
        RECT 92.200 130.000 93.200 130.200 ;
        RECT 95.600 129.600 96.400 130.200 ;
        RECT 68.200 129.000 77.200 129.600 ;
        RECT 68.200 127.400 68.800 129.000 ;
        RECT 76.400 128.800 77.200 129.000 ;
        RECT 79.600 129.000 88.200 129.600 ;
        RECT 79.600 128.800 80.400 129.000 ;
        RECT 71.400 127.600 74.000 128.400 ;
        RECT 68.200 126.800 70.800 127.400 ;
        RECT 70.000 122.200 70.800 126.800 ;
        RECT 73.200 122.200 74.000 127.600 ;
        RECT 74.600 126.800 78.800 127.600 ;
        RECT 76.400 122.200 77.200 125.000 ;
        RECT 78.000 122.200 78.800 125.000 ;
        RECT 79.600 122.200 80.400 125.000 ;
        RECT 81.200 122.200 82.000 128.400 ;
        RECT 84.400 127.600 87.000 128.400 ;
        RECT 87.600 128.200 88.200 129.000 ;
        RECT 89.200 129.400 90.000 129.600 ;
        RECT 89.200 129.000 94.600 129.400 ;
        RECT 89.200 128.800 95.400 129.000 ;
        RECT 94.000 128.200 95.400 128.800 ;
        RECT 87.600 127.600 93.400 128.200 ;
        RECT 96.400 128.000 98.000 128.800 ;
        RECT 96.400 127.600 97.000 128.000 ;
        RECT 84.400 122.200 85.200 127.000 ;
        RECT 87.600 122.200 88.400 127.000 ;
        RECT 92.800 126.800 97.000 127.600 ;
        RECT 98.800 127.400 99.600 133.000 ;
        RECT 104.800 132.800 105.400 136.200 ;
        RECT 110.000 135.800 110.800 139.800 ;
        RECT 113.200 136.400 114.000 139.800 ;
        RECT 106.000 135.400 107.600 135.600 ;
        RECT 106.000 134.800 108.000 135.400 ;
        RECT 108.600 135.200 110.800 135.800 ;
        RECT 113.000 135.800 114.000 136.400 ;
        RECT 108.600 135.000 109.400 135.200 ;
        RECT 107.400 134.400 108.000 134.800 ;
        RECT 113.000 134.400 113.600 135.800 ;
        RECT 116.400 135.200 117.200 139.800 ;
        RECT 118.600 136.400 119.400 139.800 ;
        RECT 118.600 135.800 120.400 136.400 ;
        RECT 114.600 134.600 117.200 135.200 ;
        RECT 106.000 133.400 106.800 134.200 ;
        RECT 107.400 133.800 110.800 134.400 ;
        RECT 109.200 133.600 110.800 133.800 ;
        RECT 113.000 133.600 114.000 134.400 ;
        RECT 104.400 132.400 105.400 132.800 ;
        RECT 103.600 132.200 105.400 132.400 ;
        RECT 106.200 132.800 106.800 133.400 ;
        RECT 106.200 132.200 108.800 132.800 ;
        RECT 103.600 131.600 105.000 132.200 ;
        RECT 108.000 132.000 108.800 132.200 ;
        RECT 104.400 130.200 105.000 131.600 ;
        RECT 105.800 131.400 106.600 131.600 ;
        RECT 105.800 130.800 109.200 131.400 ;
        RECT 108.600 130.200 109.200 130.800 ;
        RECT 113.000 130.200 113.600 133.600 ;
        RECT 114.600 133.000 115.200 134.600 ;
        RECT 118.000 134.300 118.800 134.400 ;
        RECT 119.600 134.300 120.400 135.800 ;
        RECT 122.800 135.800 123.600 139.800 ;
        RECT 127.200 136.200 128.800 139.800 ;
        RECT 122.800 135.200 125.200 135.800 ;
        RECT 118.000 133.700 120.400 134.300 ;
        RECT 118.000 133.600 118.800 133.700 ;
        RECT 114.200 132.200 115.200 133.000 ;
        RECT 114.600 130.200 115.200 132.200 ;
        RECT 116.200 132.400 117.000 133.200 ;
        RECT 116.200 131.600 117.200 132.400 ;
        RECT 97.600 126.800 99.600 127.400 ;
        RECT 100.400 129.600 102.800 130.200 ;
        RECT 104.400 129.600 106.400 130.200 ;
        RECT 89.200 122.200 90.000 125.000 ;
        RECT 90.800 122.200 91.600 125.000 ;
        RECT 94.000 122.200 94.800 126.800 ;
        RECT 97.600 126.200 98.200 126.800 ;
        RECT 97.200 125.600 98.200 126.200 ;
        RECT 97.200 122.200 98.000 125.600 ;
        RECT 100.400 122.200 101.200 129.600 ;
        RECT 102.000 129.400 102.800 129.600 ;
        RECT 104.800 124.400 106.400 129.600 ;
        RECT 108.600 129.600 110.800 130.200 ;
        RECT 108.600 129.400 109.400 129.600 ;
        RECT 103.600 123.600 106.400 124.400 ;
        RECT 104.800 122.200 106.400 123.600 ;
        RECT 110.000 122.200 110.800 129.600 ;
        RECT 113.000 129.200 114.000 130.200 ;
        RECT 114.600 129.600 117.200 130.200 ;
        RECT 113.200 122.200 114.000 129.200 ;
        RECT 116.400 122.200 117.200 129.600 ;
        RECT 118.000 128.800 118.800 130.400 ;
        RECT 119.600 122.200 120.400 133.700 ;
        RECT 121.200 134.300 122.000 135.200 ;
        RECT 124.400 135.000 125.200 135.200 ;
        RECT 125.800 134.800 126.600 135.600 ;
        RECT 125.800 134.400 126.400 134.800 ;
        RECT 122.800 134.300 124.400 134.400 ;
        RECT 121.200 133.700 124.400 134.300 ;
        RECT 121.200 133.600 122.000 133.700 ;
        RECT 122.800 133.600 124.400 133.700 ;
        RECT 125.600 133.600 126.400 134.400 ;
        RECT 127.200 134.200 127.800 136.200 ;
        RECT 132.400 135.800 133.200 139.800 ;
        RECT 128.400 134.800 130.000 135.600 ;
        RECT 130.600 135.200 133.200 135.800 ;
        RECT 130.600 135.000 131.400 135.200 ;
        RECT 131.600 134.200 133.200 134.400 ;
        RECT 127.200 133.600 128.200 134.200 ;
        RECT 131.000 134.000 133.200 134.200 ;
        RECT 127.600 132.400 128.200 133.600 ;
        RECT 128.800 133.600 133.200 134.000 ;
        RECT 134.000 133.800 134.800 139.800 ;
        RECT 140.400 136.600 141.200 139.800 ;
        RECT 142.000 137.000 142.800 139.800 ;
        RECT 143.600 137.000 144.400 139.800 ;
        RECT 145.200 137.000 146.000 139.800 ;
        RECT 148.400 137.000 149.200 139.800 ;
        RECT 151.600 137.000 152.400 139.800 ;
        RECT 153.200 137.000 154.000 139.800 ;
        RECT 154.800 137.000 155.600 139.800 ;
        RECT 156.400 137.000 157.200 139.800 ;
        RECT 138.600 135.800 141.200 136.600 ;
        RECT 158.000 136.600 158.800 139.800 ;
        RECT 144.600 135.800 149.200 136.400 ;
        RECT 138.600 135.200 139.400 135.800 ;
        RECT 136.400 134.400 139.400 135.200 ;
        RECT 128.800 133.400 131.600 133.600 ;
        RECT 128.800 133.200 129.600 133.400 ;
        RECT 134.000 133.000 142.800 133.800 ;
        RECT 144.600 133.400 145.400 135.800 ;
        RECT 148.400 135.600 149.200 135.800 ;
        RECT 150.000 135.600 151.600 136.400 ;
        RECT 154.600 135.600 155.600 136.400 ;
        RECT 158.000 135.800 160.400 136.600 ;
        RECT 146.800 133.600 147.600 135.200 ;
        RECT 148.400 134.800 149.200 135.000 ;
        RECT 148.400 134.200 152.800 134.800 ;
        RECT 152.000 134.000 152.800 134.200 ;
        RECT 127.600 131.600 128.400 132.400 ;
        RECT 130.200 132.200 131.000 132.400 ;
        RECT 129.400 131.600 131.000 132.200 ;
        RECT 127.600 130.200 128.200 131.600 ;
        RECT 129.400 131.400 130.200 131.600 ;
        RECT 122.800 129.600 125.200 130.200 ;
        RECT 122.800 122.200 123.600 129.600 ;
        RECT 124.400 129.400 125.200 129.600 ;
        RECT 127.200 122.200 128.800 130.200 ;
        RECT 130.600 129.600 133.200 130.200 ;
        RECT 130.600 129.400 131.400 129.600 ;
        RECT 132.400 122.200 133.200 129.600 ;
        RECT 134.000 127.400 134.800 133.000 ;
        RECT 143.400 132.600 145.400 133.400 ;
        RECT 149.200 132.600 152.400 133.400 ;
        RECT 154.800 132.800 155.600 135.600 ;
        RECT 159.600 135.200 160.400 135.800 ;
        RECT 159.600 134.600 161.400 135.200 ;
        RECT 160.600 133.400 161.400 134.600 ;
        RECT 164.400 134.600 165.200 139.800 ;
        RECT 166.000 136.000 166.800 139.800 ;
        RECT 166.000 135.200 167.000 136.000 ;
        RECT 174.000 135.800 174.800 139.800 ;
        RECT 178.400 136.200 180.000 139.800 ;
        RECT 174.000 135.200 176.400 135.800 ;
        RECT 164.400 134.000 165.600 134.600 ;
        RECT 160.600 132.600 164.400 133.400 ;
        RECT 135.400 132.000 136.200 132.200 ;
        RECT 137.200 132.000 138.000 132.400 ;
        RECT 140.400 132.000 141.200 132.400 ;
        RECT 158.000 132.000 158.800 132.600 ;
        RECT 165.000 132.000 165.600 134.000 ;
        RECT 135.400 131.400 158.800 132.000 ;
        RECT 164.800 131.400 165.600 132.000 ;
        RECT 164.800 129.600 165.400 131.400 ;
        RECT 166.200 130.800 167.000 135.200 ;
        RECT 175.600 135.000 176.400 135.200 ;
        RECT 177.000 134.800 177.800 135.600 ;
        RECT 177.000 134.400 177.600 134.800 ;
        RECT 174.000 134.300 175.600 134.400 ;
        RECT 169.300 133.700 175.600 134.300 ;
        RECT 167.600 132.300 168.400 132.400 ;
        RECT 169.300 132.300 169.900 133.700 ;
        RECT 174.000 133.600 175.600 133.700 ;
        RECT 176.800 133.600 177.600 134.400 ;
        RECT 178.400 132.800 179.000 136.200 ;
        RECT 183.600 135.800 184.400 139.800 ;
        RECT 179.600 135.400 181.200 135.600 ;
        RECT 179.600 134.800 181.600 135.400 ;
        RECT 182.200 135.200 184.400 135.800 ;
        RECT 186.800 137.800 187.600 139.800 ;
        RECT 182.200 135.000 183.000 135.200 ;
        RECT 181.000 134.400 181.600 134.800 ;
        RECT 186.800 134.400 187.400 137.800 ;
        RECT 188.400 135.600 189.200 137.200 ;
        RECT 191.200 136.300 192.000 139.800 ;
        RECT 193.200 136.300 194.000 136.400 ;
        RECT 191.200 135.700 194.000 136.300 ;
        RECT 179.600 133.400 180.400 134.200 ;
        RECT 181.000 133.800 184.400 134.400 ;
        RECT 182.800 133.600 184.400 133.800 ;
        RECT 186.800 133.600 187.600 134.400 ;
        RECT 191.200 134.200 192.000 135.700 ;
        RECT 193.200 135.600 194.000 135.700 ;
        RECT 196.400 135.800 197.200 139.800 ;
        RECT 200.800 138.400 202.400 139.800 ;
        RECT 199.600 137.600 202.400 138.400 ;
        RECT 200.800 136.200 202.400 137.600 ;
        RECT 196.400 135.200 198.600 135.800 ;
        RECT 199.600 135.400 201.200 135.600 ;
        RECT 197.800 135.000 198.600 135.200 ;
        RECT 199.200 134.800 201.200 135.400 ;
        RECT 199.200 134.400 199.800 134.800 ;
        RECT 190.200 133.800 192.000 134.200 ;
        RECT 196.400 133.800 199.800 134.400 ;
        RECT 190.200 133.600 191.800 133.800 ;
        RECT 196.400 133.600 198.000 133.800 ;
        RECT 178.000 132.400 179.000 132.800 ;
        RECT 167.600 131.700 169.900 132.300 ;
        RECT 177.200 132.200 179.000 132.400 ;
        RECT 179.800 132.800 180.400 133.400 ;
        RECT 179.800 132.200 182.400 132.800 ;
        RECT 167.600 131.600 168.400 131.700 ;
        RECT 177.200 131.600 178.600 132.200 ;
        RECT 181.600 132.000 182.400 132.200 ;
        RECT 183.700 132.300 184.300 133.600 ;
        RECT 185.200 132.300 186.000 132.400 ;
        RECT 183.700 131.700 186.000 132.300 ;
        RECT 143.600 129.400 144.400 129.600 ;
        RECT 139.000 129.000 144.400 129.400 ;
        RECT 138.200 128.800 144.400 129.000 ;
        RECT 145.400 129.000 154.000 129.600 ;
        RECT 135.600 128.000 137.200 128.800 ;
        RECT 138.200 128.200 139.600 128.800 ;
        RECT 145.400 128.200 146.000 129.000 ;
        RECT 153.200 128.800 154.000 129.000 ;
        RECT 156.400 129.000 165.400 129.600 ;
        RECT 156.400 128.800 157.200 129.000 ;
        RECT 136.600 127.600 137.200 128.000 ;
        RECT 140.200 127.600 146.000 128.200 ;
        RECT 146.600 127.600 149.200 128.400 ;
        RECT 134.000 126.800 136.000 127.400 ;
        RECT 136.600 126.800 140.800 127.600 ;
        RECT 135.400 126.200 136.000 126.800 ;
        RECT 135.400 125.600 136.400 126.200 ;
        RECT 135.600 122.200 136.400 125.600 ;
        RECT 138.800 122.200 139.600 126.800 ;
        RECT 142.000 122.200 142.800 125.000 ;
        RECT 143.600 122.200 144.400 125.000 ;
        RECT 145.200 122.200 146.000 127.000 ;
        RECT 148.400 122.200 149.200 127.000 ;
        RECT 151.600 122.200 152.400 128.400 ;
        RECT 159.600 127.600 162.200 128.400 ;
        RECT 154.800 126.800 159.000 127.600 ;
        RECT 153.200 122.200 154.000 125.000 ;
        RECT 154.800 122.200 155.600 125.000 ;
        RECT 156.400 122.200 157.200 125.000 ;
        RECT 159.600 122.200 160.400 127.600 ;
        RECT 164.800 127.400 165.400 129.000 ;
        RECT 162.800 126.800 165.400 127.400 ;
        RECT 166.000 130.000 167.000 130.800 ;
        RECT 178.000 130.200 178.600 131.600 ;
        RECT 179.400 131.400 180.200 131.600 ;
        RECT 179.400 130.800 182.800 131.400 ;
        RECT 185.200 130.800 186.000 131.700 ;
        RECT 182.200 130.200 182.800 130.800 ;
        RECT 186.800 130.200 187.400 133.600 ;
        RECT 190.200 130.400 190.800 133.600 ;
        RECT 200.400 133.400 201.200 134.200 ;
        RECT 200.400 132.800 201.000 133.400 ;
        RECT 192.400 131.600 194.000 132.400 ;
        RECT 198.400 132.200 201.000 132.800 ;
        RECT 201.800 132.800 202.400 136.200 ;
        RECT 206.000 135.800 206.800 139.800 ;
        RECT 208.200 138.400 209.000 139.800 ;
        RECT 207.600 137.600 209.000 138.400 ;
        RECT 208.200 136.400 209.000 137.600 ;
        RECT 208.200 135.800 210.000 136.400 ;
        RECT 203.000 134.800 203.800 135.600 ;
        RECT 204.400 135.200 206.800 135.800 ;
        RECT 204.400 135.000 205.200 135.200 ;
        RECT 203.200 134.400 203.800 134.800 ;
        RECT 203.200 133.600 204.000 134.400 ;
        RECT 205.200 133.600 206.800 134.400 ;
        RECT 201.800 132.400 202.800 132.800 ;
        RECT 201.800 132.200 203.600 132.400 ;
        RECT 198.400 132.000 199.200 132.200 ;
        RECT 202.200 131.600 203.600 132.200 ;
        RECT 200.600 131.400 201.400 131.600 ;
        RECT 162.800 122.200 163.600 126.800 ;
        RECT 166.000 122.200 166.800 130.000 ;
        RECT 174.000 129.600 176.400 130.200 ;
        RECT 178.000 129.600 180.000 130.200 ;
        RECT 174.000 122.200 174.800 129.600 ;
        RECT 175.600 129.400 176.400 129.600 ;
        RECT 178.400 124.400 180.000 129.600 ;
        RECT 182.200 129.600 184.400 130.200 ;
        RECT 182.200 129.400 183.000 129.600 ;
        RECT 177.200 123.600 180.000 124.400 ;
        RECT 178.400 122.200 180.000 123.600 ;
        RECT 183.600 122.200 184.400 129.600 ;
        RECT 185.800 129.400 187.600 130.200 ;
        RECT 190.000 129.600 190.800 130.400 ;
        RECT 194.800 129.600 195.600 131.200 ;
        RECT 198.000 130.800 201.400 131.400 ;
        RECT 198.000 130.200 198.600 130.800 ;
        RECT 202.200 130.200 202.800 131.600 ;
        RECT 196.400 129.600 198.600 130.200 ;
        RECT 185.800 128.400 186.600 129.400 ;
        RECT 185.200 127.600 186.600 128.400 ;
        RECT 185.800 122.200 186.600 127.600 ;
        RECT 190.200 127.000 190.800 129.600 ;
        RECT 191.600 127.600 192.400 129.200 ;
        RECT 190.200 126.400 193.800 127.000 ;
        RECT 190.200 126.200 190.800 126.400 ;
        RECT 190.000 122.200 190.800 126.200 ;
        RECT 193.200 126.200 193.800 126.400 ;
        RECT 193.200 122.200 194.000 126.200 ;
        RECT 196.400 122.200 197.200 129.600 ;
        RECT 197.800 129.400 198.600 129.600 ;
        RECT 200.800 129.600 202.800 130.200 ;
        RECT 204.400 129.600 206.800 130.200 ;
        RECT 200.800 122.200 202.400 129.600 ;
        RECT 204.400 129.400 205.200 129.600 ;
        RECT 206.000 122.200 206.800 129.600 ;
        RECT 207.600 128.800 208.400 130.400 ;
        RECT 209.200 122.200 210.000 135.800 ;
        RECT 212.400 135.200 213.200 139.800 ;
        RECT 210.800 133.600 211.600 135.200 ;
        RECT 212.400 134.600 214.600 135.200 ;
        RECT 210.800 132.300 211.600 132.400 ;
        RECT 212.400 132.300 213.200 133.200 ;
        RECT 210.800 131.700 213.200 132.300 ;
        RECT 210.800 131.600 211.600 131.700 ;
        RECT 212.400 131.600 213.200 131.700 ;
        RECT 214.000 131.600 214.600 134.600 ;
        RECT 214.000 130.800 215.200 131.600 ;
        RECT 214.000 130.200 214.600 130.800 ;
        RECT 212.400 129.600 214.600 130.200 ;
        RECT 212.400 122.200 213.200 129.600 ;
        RECT 4.400 112.400 5.200 119.800 ;
        RECT 9.200 112.400 10.000 119.800 ;
        RECT 3.000 111.800 5.200 112.400 ;
        RECT 7.800 111.800 10.000 112.400 ;
        RECT 10.800 112.400 11.600 119.800 ;
        RECT 12.400 112.400 13.200 112.600 ;
        RECT 15.200 112.400 16.800 119.800 ;
        RECT 10.800 111.800 13.200 112.400 ;
        RECT 14.800 111.800 16.800 112.400 ;
        RECT 19.000 112.400 19.800 112.600 ;
        RECT 20.400 112.400 21.200 119.800 ;
        RECT 19.000 111.800 21.200 112.400 ;
        RECT 3.000 111.200 3.600 111.800 ;
        RECT 7.800 111.200 8.400 111.800 ;
        RECT 2.400 110.400 3.600 111.200 ;
        RECT 7.200 110.400 8.400 111.200 ;
        RECT 14.800 110.400 15.400 111.800 ;
        RECT 19.000 111.200 19.600 111.800 ;
        RECT 16.200 110.600 19.600 111.200 ;
        RECT 16.200 110.400 17.000 110.600 ;
        RECT 3.000 107.400 3.600 110.400 ;
        RECT 4.400 108.800 5.200 110.400 ;
        RECT 7.800 107.400 8.400 110.400 ;
        RECT 9.200 108.800 10.000 110.400 ;
        RECT 14.000 109.800 15.400 110.400 ;
        RECT 18.400 109.800 19.200 110.000 ;
        RECT 14.000 109.600 15.800 109.800 ;
        RECT 14.800 109.200 15.800 109.600 ;
        RECT 10.800 107.600 12.400 108.400 ;
        RECT 13.600 107.600 14.400 108.400 ;
        RECT 3.000 106.800 5.200 107.400 ;
        RECT 7.800 106.800 10.000 107.400 ;
        RECT 13.800 107.200 14.400 107.600 ;
        RECT 12.400 106.800 13.200 107.000 ;
        RECT 4.400 102.200 5.200 106.800 ;
        RECT 9.200 102.200 10.000 106.800 ;
        RECT 10.800 106.200 13.200 106.800 ;
        RECT 13.800 106.400 14.600 107.200 ;
        RECT 10.800 102.200 11.600 106.200 ;
        RECT 15.200 105.800 15.800 109.200 ;
        RECT 16.600 109.200 19.200 109.800 ;
        RECT 16.600 108.600 17.200 109.200 ;
        RECT 16.400 107.800 17.200 108.600 ;
        RECT 19.600 108.200 21.200 108.400 ;
        RECT 17.800 107.600 21.200 108.200 ;
        RECT 17.800 107.200 18.400 107.600 ;
        RECT 16.400 106.600 18.400 107.200 ;
        RECT 19.000 106.800 19.800 107.000 ;
        RECT 16.400 106.400 18.000 106.600 ;
        RECT 19.000 106.200 21.200 106.800 ;
        RECT 15.200 102.200 16.800 105.800 ;
        RECT 20.400 102.200 21.200 106.200 ;
        RECT 22.000 104.800 22.800 106.400 ;
        RECT 23.600 102.200 24.400 119.800 ;
        RECT 25.200 104.800 26.000 106.400 ;
        RECT 26.800 102.200 27.600 119.800 ;
        RECT 30.000 115.800 30.800 119.800 ;
        RECT 30.200 115.600 30.800 115.800 ;
        RECT 33.200 115.800 34.000 119.800 ;
        RECT 33.200 115.600 33.800 115.800 ;
        RECT 30.200 115.000 33.800 115.600 ;
        RECT 31.600 112.800 32.400 114.400 ;
        RECT 33.200 112.400 33.800 115.000 ;
        RECT 38.000 112.400 38.800 119.800 ;
        RECT 28.400 110.800 29.200 112.400 ;
        RECT 33.200 111.600 34.000 112.400 ;
        RECT 36.600 111.800 38.800 112.400 ;
        RECT 30.000 109.600 31.600 110.400 ;
        RECT 33.200 108.400 33.800 111.600 ;
        RECT 36.600 111.200 37.200 111.800 ;
        RECT 36.000 110.400 37.200 111.200 ;
        RECT 41.200 111.200 42.000 119.800 ;
        RECT 44.400 111.200 45.200 119.800 ;
        RECT 47.600 112.400 48.400 119.800 ;
        RECT 50.800 112.800 51.600 119.800 ;
        RECT 47.600 111.800 50.200 112.400 ;
        RECT 50.800 111.800 51.800 112.800 ;
        RECT 60.400 112.000 61.200 119.800 ;
        RECT 63.600 115.200 64.400 119.800 ;
        RECT 41.200 110.400 45.200 111.200 ;
        RECT 32.200 108.200 33.800 108.400 ;
        RECT 32.000 107.800 33.800 108.200 ;
        RECT 32.000 104.400 32.800 107.800 ;
        RECT 36.600 107.400 37.200 110.400 ;
        RECT 38.000 110.300 38.800 110.400 ;
        RECT 39.600 110.300 40.400 110.400 ;
        RECT 38.000 109.700 40.400 110.300 ;
        RECT 38.000 108.800 38.800 109.700 ;
        RECT 39.600 109.600 40.400 109.700 ;
        RECT 41.200 107.600 42.000 110.400 ;
        RECT 44.400 110.300 45.200 110.400 ;
        RECT 47.600 110.300 48.600 110.400 ;
        RECT 44.400 109.700 48.600 110.300 ;
        RECT 47.600 109.600 48.600 109.700 ;
        RECT 47.800 108.800 48.600 109.600 ;
        RECT 49.600 109.800 50.200 111.800 ;
        RECT 49.600 109.000 50.600 109.800 ;
        RECT 36.600 106.800 38.800 107.400 ;
        RECT 32.000 103.600 34.000 104.400 ;
        RECT 32.000 102.200 32.800 103.600 ;
        RECT 38.000 102.200 38.800 106.800 ;
        RECT 41.200 106.800 45.200 107.600 ;
        RECT 49.600 107.400 50.200 109.000 ;
        RECT 51.200 108.400 51.800 111.800 ;
        RECT 60.200 111.200 61.200 112.000 ;
        RECT 61.800 114.600 64.400 115.200 ;
        RECT 61.800 113.000 62.400 114.600 ;
        RECT 66.800 114.400 67.600 119.800 ;
        RECT 70.000 117.000 70.800 119.800 ;
        RECT 71.600 117.000 72.400 119.800 ;
        RECT 73.200 117.000 74.000 119.800 ;
        RECT 68.200 114.400 72.400 115.200 ;
        RECT 65.000 113.600 67.600 114.400 ;
        RECT 74.800 113.600 75.600 119.800 ;
        RECT 78.000 115.000 78.800 119.800 ;
        RECT 81.200 115.000 82.000 119.800 ;
        RECT 82.800 117.000 83.600 119.800 ;
        RECT 84.400 117.000 85.200 119.800 ;
        RECT 87.600 115.200 88.400 119.800 ;
        RECT 90.800 116.400 91.600 119.800 ;
        RECT 90.800 115.800 91.800 116.400 ;
        RECT 91.200 115.200 91.800 115.800 ;
        RECT 86.400 114.400 90.600 115.200 ;
        RECT 91.200 114.600 93.200 115.200 ;
        RECT 78.000 113.600 80.600 114.400 ;
        RECT 81.200 113.800 87.000 114.400 ;
        RECT 90.000 114.000 90.600 114.400 ;
        RECT 70.000 113.000 70.800 113.200 ;
        RECT 61.800 112.400 70.800 113.000 ;
        RECT 73.200 113.000 74.000 113.200 ;
        RECT 81.200 113.000 81.800 113.800 ;
        RECT 87.600 113.200 89.000 113.800 ;
        RECT 90.000 113.200 91.600 114.000 ;
        RECT 73.200 112.400 81.800 113.000 ;
        RECT 82.800 113.000 89.000 113.200 ;
        RECT 82.800 112.600 88.200 113.000 ;
        RECT 82.800 112.400 83.600 112.600 ;
        RECT 50.800 108.300 51.800 108.400 ;
        RECT 58.800 108.300 59.600 108.400 ;
        RECT 50.800 107.700 59.600 108.300 ;
        RECT 50.800 107.600 51.800 107.700 ;
        RECT 58.800 107.600 59.600 107.700 ;
        RECT 41.200 102.200 42.000 106.800 ;
        RECT 44.400 102.200 45.200 106.800 ;
        RECT 47.600 106.800 50.200 107.400 ;
        RECT 47.600 102.200 48.400 106.800 ;
        RECT 51.200 106.200 51.800 107.600 ;
        RECT 50.800 105.600 51.800 106.200 ;
        RECT 60.200 106.800 61.000 111.200 ;
        RECT 61.800 110.600 62.400 112.400 ;
        RECT 61.600 110.000 62.400 110.600 ;
        RECT 68.400 110.000 91.800 110.600 ;
        RECT 61.600 108.000 62.200 110.000 ;
        RECT 68.400 109.400 69.200 110.000 ;
        RECT 86.000 109.600 86.800 110.000 ;
        RECT 90.800 109.800 91.800 110.000 ;
        RECT 90.800 109.600 91.600 109.800 ;
        RECT 62.800 108.600 66.600 109.400 ;
        RECT 61.600 107.400 62.800 108.000 ;
        RECT 60.200 106.000 61.200 106.800 ;
        RECT 50.800 102.200 51.600 105.600 ;
        RECT 60.400 102.200 61.200 106.000 ;
        RECT 62.000 102.200 62.800 107.400 ;
        RECT 65.800 107.400 66.600 108.600 ;
        RECT 65.800 106.800 67.600 107.400 ;
        RECT 66.800 106.200 67.600 106.800 ;
        RECT 71.600 106.400 72.400 109.200 ;
        RECT 74.800 108.600 78.000 109.400 ;
        RECT 81.800 108.600 83.800 109.400 ;
        RECT 92.400 109.000 93.200 114.600 ;
        RECT 95.600 112.000 96.400 119.800 ;
        RECT 98.800 115.200 99.600 119.800 ;
        RECT 74.400 107.800 75.200 108.000 ;
        RECT 74.400 107.200 78.800 107.800 ;
        RECT 78.000 107.000 78.800 107.200 ;
        RECT 79.600 106.800 80.400 108.400 ;
        RECT 66.800 105.400 69.200 106.200 ;
        RECT 71.600 105.600 72.600 106.400 ;
        RECT 75.600 105.600 77.200 106.400 ;
        RECT 78.000 106.200 78.800 106.400 ;
        RECT 81.800 106.200 82.600 108.600 ;
        RECT 84.400 108.200 93.200 109.000 ;
        RECT 87.800 106.800 90.800 107.600 ;
        RECT 87.800 106.200 88.600 106.800 ;
        RECT 78.000 105.600 82.600 106.200 ;
        RECT 68.400 102.200 69.200 105.400 ;
        RECT 86.000 105.400 88.600 106.200 ;
        RECT 70.000 102.200 70.800 105.000 ;
        RECT 71.600 102.200 72.400 105.000 ;
        RECT 73.200 102.200 74.000 105.000 ;
        RECT 74.800 102.200 75.600 105.000 ;
        RECT 78.000 102.200 78.800 105.000 ;
        RECT 81.200 102.200 82.000 105.000 ;
        RECT 82.800 102.200 83.600 105.000 ;
        RECT 84.400 102.200 85.200 105.000 ;
        RECT 86.000 102.200 86.800 105.400 ;
        RECT 92.400 102.200 93.200 108.200 ;
        RECT 95.400 111.200 96.400 112.000 ;
        RECT 97.000 114.600 99.600 115.200 ;
        RECT 97.000 113.000 97.600 114.600 ;
        RECT 102.000 114.400 102.800 119.800 ;
        RECT 105.200 117.000 106.000 119.800 ;
        RECT 106.800 117.000 107.600 119.800 ;
        RECT 108.400 117.000 109.200 119.800 ;
        RECT 103.400 114.400 107.600 115.200 ;
        RECT 100.200 113.600 102.800 114.400 ;
        RECT 110.000 113.600 110.800 119.800 ;
        RECT 113.200 115.000 114.000 119.800 ;
        RECT 116.400 115.000 117.200 119.800 ;
        RECT 118.000 117.000 118.800 119.800 ;
        RECT 119.600 117.000 120.400 119.800 ;
        RECT 122.800 115.200 123.600 119.800 ;
        RECT 126.000 116.400 126.800 119.800 ;
        RECT 126.000 115.800 127.000 116.400 ;
        RECT 126.400 115.200 127.000 115.800 ;
        RECT 121.600 114.400 125.800 115.200 ;
        RECT 126.400 114.600 128.400 115.200 ;
        RECT 113.200 113.600 115.800 114.400 ;
        RECT 116.400 113.800 122.200 114.400 ;
        RECT 125.200 114.000 125.800 114.400 ;
        RECT 105.200 113.000 106.000 113.200 ;
        RECT 97.000 112.400 106.000 113.000 ;
        RECT 108.400 113.000 109.200 113.200 ;
        RECT 116.400 113.000 117.000 113.800 ;
        RECT 122.800 113.200 124.200 113.800 ;
        RECT 125.200 113.200 126.800 114.000 ;
        RECT 108.400 112.400 117.000 113.000 ;
        RECT 118.000 113.000 124.200 113.200 ;
        RECT 118.000 112.600 123.400 113.000 ;
        RECT 118.000 112.400 118.800 112.600 ;
        RECT 95.400 106.800 96.200 111.200 ;
        RECT 97.000 110.600 97.600 112.400 ;
        RECT 96.800 110.000 97.600 110.600 ;
        RECT 103.600 110.000 127.000 110.600 ;
        RECT 96.800 108.000 97.400 110.000 ;
        RECT 103.600 109.400 104.400 110.000 ;
        RECT 121.200 109.600 122.000 110.000 ;
        RECT 124.400 109.600 125.200 110.000 ;
        RECT 126.200 109.800 127.000 110.000 ;
        RECT 98.000 108.600 101.800 109.400 ;
        RECT 96.800 107.400 98.000 108.000 ;
        RECT 94.000 106.300 94.800 106.400 ;
        RECT 95.400 106.300 96.400 106.800 ;
        RECT 94.000 105.700 96.400 106.300 ;
        RECT 94.000 105.600 94.800 105.700 ;
        RECT 95.600 102.200 96.400 105.700 ;
        RECT 97.200 102.200 98.000 107.400 ;
        RECT 101.000 107.400 101.800 108.600 ;
        RECT 101.000 106.800 102.800 107.400 ;
        RECT 102.000 106.200 102.800 106.800 ;
        RECT 106.800 106.400 107.600 109.200 ;
        RECT 110.000 108.600 113.200 109.400 ;
        RECT 117.000 108.600 119.000 109.400 ;
        RECT 127.600 109.000 128.400 114.600 ;
        RECT 129.200 112.400 130.000 119.800 ;
        RECT 132.400 112.800 133.200 119.800 ;
        RECT 137.200 116.400 138.000 119.800 ;
        RECT 137.000 115.800 138.000 116.400 ;
        RECT 137.000 115.200 137.600 115.800 ;
        RECT 140.400 115.200 141.200 119.800 ;
        RECT 143.600 117.000 144.400 119.800 ;
        RECT 145.200 117.000 146.000 119.800 ;
        RECT 135.600 114.600 137.600 115.200 ;
        RECT 129.200 111.800 131.800 112.400 ;
        RECT 132.400 111.800 133.400 112.800 ;
        RECT 129.200 109.600 130.200 110.400 ;
        RECT 109.600 107.800 110.400 108.000 ;
        RECT 109.600 107.200 114.000 107.800 ;
        RECT 113.200 107.000 114.000 107.200 ;
        RECT 114.800 106.800 115.600 108.400 ;
        RECT 102.000 105.400 104.400 106.200 ;
        RECT 106.800 105.600 107.800 106.400 ;
        RECT 110.800 105.600 112.400 106.400 ;
        RECT 113.200 106.200 114.000 106.400 ;
        RECT 117.000 106.200 117.800 108.600 ;
        RECT 119.600 108.200 128.400 109.000 ;
        RECT 129.400 108.800 130.200 109.600 ;
        RECT 131.200 109.800 131.800 111.800 ;
        RECT 131.200 109.000 132.200 109.800 ;
        RECT 123.000 106.800 126.000 107.600 ;
        RECT 123.000 106.200 123.800 106.800 ;
        RECT 113.200 105.600 117.800 106.200 ;
        RECT 103.600 102.200 104.400 105.400 ;
        RECT 121.200 105.400 123.800 106.200 ;
        RECT 105.200 102.200 106.000 105.000 ;
        RECT 106.800 102.200 107.600 105.000 ;
        RECT 108.400 102.200 109.200 105.000 ;
        RECT 110.000 102.200 110.800 105.000 ;
        RECT 113.200 102.200 114.000 105.000 ;
        RECT 116.400 102.200 117.200 105.000 ;
        RECT 118.000 102.200 118.800 105.000 ;
        RECT 119.600 102.200 120.400 105.000 ;
        RECT 121.200 102.200 122.000 105.400 ;
        RECT 127.600 102.200 128.400 108.200 ;
        RECT 131.200 107.400 131.800 109.000 ;
        RECT 132.800 108.400 133.400 111.800 ;
        RECT 135.600 109.000 136.400 114.600 ;
        RECT 138.200 114.400 142.400 115.200 ;
        RECT 146.800 115.000 147.600 119.800 ;
        RECT 150.000 115.000 150.800 119.800 ;
        RECT 138.200 114.000 138.800 114.400 ;
        RECT 137.200 113.200 138.800 114.000 ;
        RECT 141.800 113.800 147.600 114.400 ;
        RECT 139.800 113.200 141.200 113.800 ;
        RECT 139.800 113.000 146.000 113.200 ;
        RECT 140.600 112.600 146.000 113.000 ;
        RECT 145.200 112.400 146.000 112.600 ;
        RECT 147.000 113.000 147.600 113.800 ;
        RECT 148.200 113.600 150.800 114.400 ;
        RECT 153.200 113.600 154.000 119.800 ;
        RECT 154.800 117.000 155.600 119.800 ;
        RECT 156.400 117.000 157.200 119.800 ;
        RECT 158.000 117.000 158.800 119.800 ;
        RECT 156.400 114.400 160.600 115.200 ;
        RECT 161.200 114.400 162.000 119.800 ;
        RECT 164.400 115.200 165.200 119.800 ;
        RECT 164.400 114.600 167.000 115.200 ;
        RECT 161.200 113.600 163.800 114.400 ;
        RECT 154.800 113.000 155.600 113.200 ;
        RECT 147.000 112.400 155.600 113.000 ;
        RECT 158.000 113.000 158.800 113.200 ;
        RECT 166.400 113.000 167.000 114.600 ;
        RECT 158.000 112.400 167.000 113.000 ;
        RECT 166.400 110.600 167.000 112.400 ;
        RECT 167.600 112.000 168.400 119.800 ;
        RECT 177.200 116.400 178.000 119.800 ;
        RECT 177.000 115.800 178.000 116.400 ;
        RECT 177.000 115.200 177.600 115.800 ;
        RECT 180.400 115.200 181.200 119.800 ;
        RECT 183.600 117.000 184.400 119.800 ;
        RECT 185.200 117.000 186.000 119.800 ;
        RECT 175.600 114.600 177.600 115.200 ;
        RECT 167.600 111.200 168.600 112.000 ;
        RECT 137.000 110.000 160.400 110.600 ;
        RECT 166.400 110.000 167.200 110.600 ;
        RECT 137.000 109.800 137.800 110.000 ;
        RECT 138.800 109.600 139.600 110.000 ;
        RECT 142.000 109.600 142.800 110.000 ;
        RECT 159.600 109.400 160.400 110.000 ;
        RECT 132.400 108.300 133.400 108.400 ;
        RECT 134.000 108.300 134.800 108.400 ;
        RECT 132.400 107.700 134.800 108.300 ;
        RECT 132.400 107.600 133.400 107.700 ;
        RECT 134.000 107.600 134.800 107.700 ;
        RECT 135.600 108.200 144.400 109.000 ;
        RECT 145.000 108.600 147.000 109.400 ;
        RECT 150.800 108.600 154.000 109.400 ;
        RECT 129.200 106.800 131.800 107.400 ;
        RECT 129.200 102.200 130.000 106.800 ;
        RECT 132.800 106.200 133.400 107.600 ;
        RECT 132.400 105.600 133.400 106.200 ;
        RECT 132.400 102.200 133.200 105.600 ;
        RECT 135.600 102.200 136.400 108.200 ;
        RECT 138.000 106.800 141.000 107.600 ;
        RECT 140.200 106.200 141.000 106.800 ;
        RECT 146.200 106.200 147.000 108.600 ;
        RECT 148.400 106.800 149.200 108.400 ;
        RECT 153.600 107.800 154.400 108.000 ;
        RECT 150.000 107.200 154.400 107.800 ;
        RECT 150.000 107.000 150.800 107.200 ;
        RECT 156.400 106.400 157.200 109.200 ;
        RECT 162.200 108.600 166.000 109.400 ;
        RECT 162.200 107.400 163.000 108.600 ;
        RECT 166.600 108.000 167.200 110.000 ;
        RECT 150.000 106.200 150.800 106.400 ;
        RECT 140.200 105.400 142.800 106.200 ;
        RECT 146.200 105.600 150.800 106.200 ;
        RECT 151.600 105.600 153.200 106.400 ;
        RECT 156.200 105.600 157.200 106.400 ;
        RECT 161.200 106.800 163.000 107.400 ;
        RECT 166.000 107.400 167.200 108.000 ;
        RECT 161.200 106.200 162.000 106.800 ;
        RECT 142.000 102.200 142.800 105.400 ;
        RECT 159.600 105.400 162.000 106.200 ;
        RECT 143.600 102.200 144.400 105.000 ;
        RECT 145.200 102.200 146.000 105.000 ;
        RECT 146.800 102.200 147.600 105.000 ;
        RECT 150.000 102.200 150.800 105.000 ;
        RECT 153.200 102.200 154.000 105.000 ;
        RECT 154.800 102.200 155.600 105.000 ;
        RECT 156.400 102.200 157.200 105.000 ;
        RECT 158.000 102.200 158.800 105.000 ;
        RECT 159.600 102.200 160.400 105.400 ;
        RECT 166.000 102.200 166.800 107.400 ;
        RECT 167.800 106.800 168.600 111.200 ;
        RECT 167.600 106.000 168.600 106.800 ;
        RECT 175.600 109.000 176.400 114.600 ;
        RECT 178.200 114.400 182.400 115.200 ;
        RECT 186.800 115.000 187.600 119.800 ;
        RECT 190.000 115.000 190.800 119.800 ;
        RECT 178.200 114.000 178.800 114.400 ;
        RECT 177.200 113.200 178.800 114.000 ;
        RECT 181.800 113.800 187.600 114.400 ;
        RECT 179.800 113.200 181.200 113.800 ;
        RECT 179.800 113.000 186.000 113.200 ;
        RECT 180.600 112.600 186.000 113.000 ;
        RECT 185.200 112.400 186.000 112.600 ;
        RECT 187.000 113.000 187.600 113.800 ;
        RECT 188.200 113.600 190.800 114.400 ;
        RECT 193.200 113.600 194.000 119.800 ;
        RECT 194.800 117.000 195.600 119.800 ;
        RECT 196.400 117.000 197.200 119.800 ;
        RECT 198.000 117.000 198.800 119.800 ;
        RECT 196.400 114.400 200.600 115.200 ;
        RECT 201.200 114.400 202.000 119.800 ;
        RECT 204.400 115.200 205.200 119.800 ;
        RECT 204.400 114.600 207.000 115.200 ;
        RECT 201.200 113.600 203.800 114.400 ;
        RECT 194.800 113.000 195.600 113.200 ;
        RECT 187.000 112.400 195.600 113.000 ;
        RECT 198.000 113.000 198.800 113.200 ;
        RECT 206.400 113.000 207.000 114.600 ;
        RECT 198.000 112.400 207.000 113.000 ;
        RECT 206.400 110.600 207.000 112.400 ;
        RECT 207.600 112.000 208.400 119.800 ;
        RECT 210.800 112.400 211.600 119.800 ;
        RECT 207.600 111.200 208.600 112.000 ;
        RECT 210.800 111.800 213.000 112.400 ;
        RECT 177.000 110.000 200.400 110.600 ;
        RECT 206.400 110.000 207.200 110.600 ;
        RECT 177.000 109.800 177.800 110.000 ;
        RECT 178.800 109.600 179.600 110.000 ;
        RECT 182.000 109.600 182.800 110.000 ;
        RECT 199.600 109.400 200.400 110.000 ;
        RECT 175.600 108.200 184.400 109.000 ;
        RECT 185.000 108.600 187.000 109.400 ;
        RECT 190.800 108.600 194.000 109.400 ;
        RECT 167.600 102.200 168.400 106.000 ;
        RECT 175.600 102.200 176.400 108.200 ;
        RECT 178.000 106.800 181.000 107.600 ;
        RECT 180.200 106.200 181.000 106.800 ;
        RECT 186.200 106.200 187.000 108.600 ;
        RECT 188.400 106.800 189.200 108.400 ;
        RECT 193.600 107.800 194.400 108.000 ;
        RECT 190.000 107.200 194.400 107.800 ;
        RECT 190.000 107.000 190.800 107.200 ;
        RECT 196.400 106.400 197.200 109.200 ;
        RECT 202.200 108.600 206.000 109.400 ;
        RECT 202.200 107.400 203.000 108.600 ;
        RECT 206.600 108.000 207.200 110.000 ;
        RECT 190.000 106.200 190.800 106.400 ;
        RECT 180.200 105.400 182.800 106.200 ;
        RECT 186.200 105.600 190.800 106.200 ;
        RECT 191.600 105.600 193.200 106.400 ;
        RECT 196.200 105.600 197.200 106.400 ;
        RECT 201.200 106.800 203.000 107.400 ;
        RECT 206.000 107.400 207.200 108.000 ;
        RECT 207.800 110.300 208.600 111.200 ;
        RECT 212.400 111.200 213.000 111.800 ;
        RECT 212.400 110.400 213.600 111.200 ;
        RECT 210.800 110.300 211.600 110.400 ;
        RECT 207.800 109.700 211.600 110.300 ;
        RECT 201.200 106.200 202.000 106.800 ;
        RECT 182.000 102.200 182.800 105.400 ;
        RECT 199.600 105.400 202.000 106.200 ;
        RECT 183.600 102.200 184.400 105.000 ;
        RECT 185.200 102.200 186.000 105.000 ;
        RECT 186.800 102.200 187.600 105.000 ;
        RECT 190.000 102.200 190.800 105.000 ;
        RECT 193.200 102.200 194.000 105.000 ;
        RECT 194.800 102.200 195.600 105.000 ;
        RECT 196.400 102.200 197.200 105.000 ;
        RECT 198.000 102.200 198.800 105.000 ;
        RECT 199.600 102.200 200.400 105.400 ;
        RECT 206.000 102.200 206.800 107.400 ;
        RECT 207.800 106.800 208.600 109.700 ;
        RECT 210.800 108.800 211.600 109.700 ;
        RECT 212.400 107.400 213.000 110.400 ;
        RECT 207.600 106.000 208.600 106.800 ;
        RECT 210.800 106.800 213.000 107.400 ;
        RECT 207.600 102.200 208.400 106.000 ;
        RECT 210.800 102.200 211.600 106.800 ;
        RECT 2.800 96.000 3.600 99.800 ;
        RECT 2.600 95.200 3.600 96.000 ;
        RECT 2.600 90.800 3.400 95.200 ;
        RECT 4.400 94.600 5.200 99.800 ;
        RECT 10.800 96.600 11.600 99.800 ;
        RECT 12.400 97.000 13.200 99.800 ;
        RECT 14.000 97.000 14.800 99.800 ;
        RECT 15.600 97.000 16.400 99.800 ;
        RECT 17.200 97.000 18.000 99.800 ;
        RECT 20.400 97.000 21.200 99.800 ;
        RECT 23.600 97.000 24.400 99.800 ;
        RECT 25.200 97.000 26.000 99.800 ;
        RECT 26.800 97.000 27.600 99.800 ;
        RECT 9.200 95.800 11.600 96.600 ;
        RECT 28.400 96.600 29.200 99.800 ;
        RECT 9.200 95.200 10.000 95.800 ;
        RECT 4.000 94.000 5.200 94.600 ;
        RECT 8.200 94.600 10.000 95.200 ;
        RECT 14.000 95.600 15.000 96.400 ;
        RECT 18.000 95.600 19.600 96.400 ;
        RECT 20.400 95.800 25.000 96.400 ;
        RECT 28.400 95.800 31.000 96.600 ;
        RECT 20.400 95.600 21.200 95.800 ;
        RECT 4.000 92.000 4.600 94.000 ;
        RECT 8.200 93.400 9.000 94.600 ;
        RECT 5.200 92.600 9.000 93.400 ;
        RECT 14.000 92.800 14.800 95.600 ;
        RECT 20.400 94.800 21.200 95.000 ;
        RECT 16.800 94.200 21.200 94.800 ;
        RECT 16.800 94.000 17.600 94.200 ;
        RECT 22.000 93.600 22.800 95.200 ;
        RECT 24.200 93.400 25.000 95.800 ;
        RECT 30.200 95.200 31.000 95.800 ;
        RECT 30.200 94.400 33.200 95.200 ;
        RECT 34.800 93.800 35.600 99.800 ;
        RECT 38.000 96.000 38.800 99.800 ;
        RECT 17.200 92.600 20.400 93.400 ;
        RECT 24.200 92.600 26.200 93.400 ;
        RECT 26.800 93.000 35.600 93.800 ;
        RECT 4.000 91.400 4.800 92.000 ;
        RECT 2.600 90.000 3.600 90.800 ;
        RECT 2.800 82.200 3.600 90.000 ;
        RECT 4.200 89.600 4.800 91.400 ;
        RECT 5.400 90.800 6.200 91.000 ;
        RECT 5.400 90.200 32.400 90.800 ;
        RECT 28.200 90.000 29.000 90.200 ;
        RECT 31.600 89.600 32.400 90.200 ;
        RECT 4.200 89.000 13.200 89.600 ;
        RECT 4.200 87.400 4.800 89.000 ;
        RECT 12.400 88.800 13.200 89.000 ;
        RECT 15.600 89.000 24.200 89.600 ;
        RECT 15.600 88.800 16.400 89.000 ;
        RECT 7.400 87.600 10.000 88.400 ;
        RECT 4.200 86.800 6.800 87.400 ;
        RECT 6.000 82.200 6.800 86.800 ;
        RECT 9.200 82.200 10.000 87.600 ;
        RECT 10.600 86.800 14.800 87.600 ;
        RECT 12.400 82.200 13.200 85.000 ;
        RECT 14.000 82.200 14.800 85.000 ;
        RECT 15.600 82.200 16.400 85.000 ;
        RECT 17.200 82.200 18.000 88.400 ;
        RECT 20.400 87.600 23.000 88.400 ;
        RECT 23.600 88.200 24.200 89.000 ;
        RECT 25.200 89.400 26.000 89.600 ;
        RECT 25.200 89.000 30.600 89.400 ;
        RECT 25.200 88.800 31.400 89.000 ;
        RECT 30.000 88.200 31.400 88.800 ;
        RECT 23.600 87.600 29.400 88.200 ;
        RECT 32.400 88.000 34.000 88.800 ;
        RECT 32.400 87.600 33.000 88.000 ;
        RECT 20.400 82.200 21.200 87.000 ;
        RECT 23.600 82.200 24.400 87.000 ;
        RECT 28.800 86.800 33.000 87.600 ;
        RECT 34.800 87.400 35.600 93.000 ;
        RECT 37.800 95.200 38.800 96.000 ;
        RECT 37.800 90.800 38.600 95.200 ;
        RECT 39.600 94.600 40.400 99.800 ;
        RECT 46.000 96.600 46.800 99.800 ;
        RECT 47.600 97.000 48.400 99.800 ;
        RECT 49.200 97.000 50.000 99.800 ;
        RECT 50.800 97.000 51.600 99.800 ;
        RECT 52.400 97.000 53.200 99.800 ;
        RECT 55.600 97.000 56.400 99.800 ;
        RECT 58.800 97.000 59.600 99.800 ;
        RECT 60.400 97.000 61.200 99.800 ;
        RECT 62.000 97.000 62.800 99.800 ;
        RECT 44.400 95.800 46.800 96.600 ;
        RECT 63.600 96.600 64.400 99.800 ;
        RECT 44.400 95.200 45.200 95.800 ;
        RECT 39.200 94.000 40.400 94.600 ;
        RECT 43.400 94.600 45.200 95.200 ;
        RECT 49.200 95.600 50.200 96.400 ;
        RECT 53.200 95.600 54.800 96.400 ;
        RECT 55.600 95.800 60.200 96.400 ;
        RECT 63.600 95.800 66.200 96.600 ;
        RECT 55.600 95.600 56.400 95.800 ;
        RECT 39.200 92.000 39.800 94.000 ;
        RECT 43.400 93.400 44.200 94.600 ;
        RECT 40.400 92.600 44.200 93.400 ;
        RECT 49.200 92.800 50.000 95.600 ;
        RECT 55.600 94.800 56.400 95.000 ;
        RECT 52.000 94.200 56.400 94.800 ;
        RECT 52.000 94.000 52.800 94.200 ;
        RECT 57.200 93.600 58.000 95.200 ;
        RECT 59.400 93.400 60.200 95.800 ;
        RECT 65.400 95.200 66.200 95.800 ;
        RECT 65.400 94.400 68.400 95.200 ;
        RECT 70.000 93.800 70.800 99.800 ;
        RECT 78.000 96.400 78.800 99.800 ;
        RECT 52.400 92.600 55.600 93.400 ;
        RECT 59.400 92.600 61.400 93.400 ;
        RECT 62.000 93.000 70.800 93.800 ;
        RECT 39.200 91.400 40.000 92.000 ;
        RECT 37.800 90.000 38.800 90.800 ;
        RECT 33.600 86.800 35.600 87.400 ;
        RECT 25.200 82.200 26.000 85.000 ;
        RECT 26.800 82.200 27.600 85.000 ;
        RECT 30.000 82.200 30.800 86.800 ;
        RECT 33.600 86.200 34.200 86.800 ;
        RECT 33.200 85.600 34.200 86.200 ;
        RECT 33.200 82.200 34.000 85.600 ;
        RECT 38.000 82.200 38.800 90.000 ;
        RECT 39.400 89.600 40.000 91.400 ;
        RECT 40.600 90.800 41.400 91.000 ;
        RECT 40.600 90.200 67.600 90.800 ;
        RECT 63.400 90.000 64.200 90.200 ;
        RECT 66.800 89.600 67.600 90.200 ;
        RECT 39.400 89.000 48.400 89.600 ;
        RECT 39.400 87.400 40.000 89.000 ;
        RECT 47.600 88.800 48.400 89.000 ;
        RECT 50.800 89.000 59.400 89.600 ;
        RECT 50.800 88.800 51.600 89.000 ;
        RECT 42.600 87.600 45.200 88.400 ;
        RECT 39.400 86.800 42.000 87.400 ;
        RECT 41.200 82.200 42.000 86.800 ;
        RECT 44.400 82.200 45.200 87.600 ;
        RECT 45.800 86.800 50.000 87.600 ;
        RECT 47.600 82.200 48.400 85.000 ;
        RECT 49.200 82.200 50.000 85.000 ;
        RECT 50.800 82.200 51.600 85.000 ;
        RECT 52.400 82.200 53.200 88.400 ;
        RECT 55.600 87.600 58.200 88.400 ;
        RECT 58.800 88.200 59.400 89.000 ;
        RECT 60.400 89.400 61.200 89.600 ;
        RECT 60.400 89.000 65.800 89.400 ;
        RECT 60.400 88.800 66.600 89.000 ;
        RECT 65.200 88.200 66.600 88.800 ;
        RECT 58.800 87.600 64.600 88.200 ;
        RECT 67.600 88.000 69.200 88.800 ;
        RECT 67.600 87.600 68.200 88.000 ;
        RECT 55.600 82.200 56.400 87.000 ;
        RECT 58.800 82.200 59.600 87.000 ;
        RECT 64.000 86.800 68.200 87.600 ;
        RECT 70.000 87.400 70.800 93.000 ;
        RECT 77.800 95.800 78.800 96.400 ;
        RECT 77.800 94.400 78.400 95.800 ;
        RECT 81.200 95.200 82.000 99.800 ;
        RECT 82.800 95.800 83.600 99.800 ;
        RECT 87.200 98.400 88.800 99.800 ;
        RECT 87.200 97.600 90.000 98.400 ;
        RECT 87.200 96.200 88.800 97.600 ;
        RECT 82.800 95.200 85.000 95.800 ;
        RECT 86.000 95.400 87.600 95.600 ;
        RECT 79.400 94.600 82.000 95.200 ;
        RECT 84.200 95.000 85.000 95.200 ;
        RECT 85.600 94.800 87.600 95.400 ;
        RECT 77.800 93.600 78.800 94.400 ;
        RECT 77.800 90.200 78.400 93.600 ;
        RECT 79.400 93.000 80.000 94.600 ;
        RECT 85.600 94.400 86.200 94.800 ;
        RECT 82.800 93.800 86.200 94.400 ;
        RECT 82.800 93.600 84.400 93.800 ;
        RECT 86.800 93.400 87.600 94.200 ;
        RECT 79.000 92.200 80.000 93.000 ;
        RECT 79.400 90.200 80.000 92.200 ;
        RECT 81.000 92.400 81.800 93.200 ;
        RECT 86.800 92.800 87.400 93.400 ;
        RECT 81.000 91.600 82.000 92.400 ;
        RECT 84.800 92.200 87.400 92.800 ;
        RECT 88.200 92.800 88.800 96.200 ;
        RECT 92.400 95.800 93.200 99.800 ;
        RECT 94.000 96.000 94.800 99.800 ;
        RECT 97.200 96.000 98.000 99.800 ;
        RECT 94.000 95.800 98.000 96.000 ;
        RECT 98.800 95.800 99.600 99.800 ;
        RECT 89.400 94.800 90.200 95.600 ;
        RECT 90.800 95.200 93.200 95.800 ;
        RECT 94.200 95.400 97.800 95.800 ;
        RECT 90.800 95.000 91.600 95.200 ;
        RECT 89.600 94.400 90.200 94.800 ;
        RECT 94.800 94.400 95.600 94.800 ;
        RECT 98.800 94.400 99.400 95.800 ;
        RECT 100.400 95.600 101.200 97.200 ;
        RECT 89.600 93.600 90.400 94.400 ;
        RECT 91.600 94.300 93.200 94.400 ;
        RECT 94.000 94.300 95.600 94.400 ;
        RECT 91.600 93.800 95.600 94.300 ;
        RECT 97.000 94.300 99.600 94.400 ;
        RECT 100.400 94.300 101.200 94.400 ;
        RECT 91.600 93.700 94.800 93.800 ;
        RECT 91.600 93.600 93.200 93.700 ;
        RECT 94.000 93.600 94.800 93.700 ;
        RECT 97.000 93.700 101.200 94.300 ;
        RECT 97.000 93.600 99.600 93.700 ;
        RECT 100.400 93.600 101.200 93.700 ;
        RECT 88.200 92.400 89.200 92.800 ;
        RECT 88.200 92.200 90.000 92.400 ;
        RECT 84.800 92.000 85.600 92.200 ;
        RECT 88.600 91.600 90.000 92.200 ;
        RECT 95.600 91.600 96.400 93.200 ;
        RECT 87.000 91.400 87.800 91.600 ;
        RECT 84.400 90.800 87.800 91.400 ;
        RECT 84.400 90.200 85.000 90.800 ;
        RECT 88.600 90.200 89.200 91.600 ;
        RECT 97.000 90.200 97.600 93.600 ;
        RECT 98.800 90.300 99.600 90.400 ;
        RECT 100.400 90.300 101.200 90.400 ;
        RECT 98.800 90.200 101.200 90.300 ;
        RECT 77.800 89.200 78.800 90.200 ;
        RECT 79.400 89.600 82.000 90.200 ;
        RECT 68.800 86.800 70.800 87.400 ;
        RECT 60.400 82.200 61.200 85.000 ;
        RECT 62.000 82.200 62.800 85.000 ;
        RECT 65.200 82.200 66.000 86.800 ;
        RECT 68.800 86.200 69.400 86.800 ;
        RECT 68.400 85.600 69.400 86.200 ;
        RECT 68.400 82.200 69.200 85.600 ;
        RECT 78.000 82.200 78.800 89.200 ;
        RECT 81.200 82.200 82.000 89.600 ;
        RECT 82.800 89.600 85.000 90.200 ;
        RECT 82.800 82.200 83.600 89.600 ;
        RECT 84.200 89.400 85.000 89.600 ;
        RECT 87.200 89.600 89.200 90.200 ;
        RECT 90.800 89.600 93.200 90.200 ;
        RECT 87.200 82.200 88.800 89.600 ;
        RECT 90.800 89.400 91.600 89.600 ;
        RECT 92.400 82.200 93.200 89.600 ;
        RECT 96.600 89.600 97.600 90.200 ;
        RECT 98.200 89.700 101.200 90.200 ;
        RECT 98.200 89.600 99.600 89.700 ;
        RECT 100.400 89.600 101.200 89.700 ;
        RECT 96.600 82.200 97.400 89.600 ;
        RECT 98.200 88.400 98.800 89.600 ;
        RECT 98.000 87.600 98.800 88.400 ;
        RECT 102.000 88.300 102.800 99.800 ;
        RECT 106.200 96.400 107.000 99.800 ;
        RECT 105.200 95.800 107.000 96.400 ;
        RECT 110.000 96.000 110.800 99.800 ;
        RECT 103.600 93.600 104.400 95.200 ;
        RECT 105.200 94.300 106.000 95.800 ;
        RECT 109.800 95.200 110.800 96.000 ;
        RECT 108.400 94.300 109.200 94.400 ;
        RECT 105.200 93.700 109.200 94.300 ;
        RECT 103.600 88.300 104.400 88.400 ;
        RECT 102.000 87.700 104.400 88.300 ;
        RECT 102.000 82.200 102.800 87.700 ;
        RECT 103.600 87.600 104.400 87.700 ;
        RECT 105.200 82.200 106.000 93.700 ;
        RECT 108.400 93.600 109.200 93.700 ;
        RECT 109.800 90.800 110.600 95.200 ;
        RECT 111.600 94.600 112.400 99.800 ;
        RECT 118.000 96.600 118.800 99.800 ;
        RECT 119.600 97.000 120.400 99.800 ;
        RECT 121.200 97.000 122.000 99.800 ;
        RECT 122.800 97.000 123.600 99.800 ;
        RECT 124.400 97.000 125.200 99.800 ;
        RECT 127.600 97.000 128.400 99.800 ;
        RECT 130.800 97.000 131.600 99.800 ;
        RECT 132.400 97.000 133.200 99.800 ;
        RECT 134.000 97.000 134.800 99.800 ;
        RECT 116.400 95.800 118.800 96.600 ;
        RECT 135.600 96.600 136.400 99.800 ;
        RECT 116.400 95.200 117.200 95.800 ;
        RECT 111.200 94.000 112.400 94.600 ;
        RECT 115.400 94.600 117.200 95.200 ;
        RECT 121.200 95.600 122.200 96.400 ;
        RECT 125.200 95.600 126.800 96.400 ;
        RECT 127.600 95.800 132.200 96.400 ;
        RECT 135.600 95.800 138.200 96.600 ;
        RECT 127.600 95.600 128.400 95.800 ;
        RECT 111.200 92.000 111.800 94.000 ;
        RECT 115.400 93.400 116.200 94.600 ;
        RECT 112.400 92.600 116.200 93.400 ;
        RECT 121.200 92.800 122.000 95.600 ;
        RECT 127.600 94.800 128.400 95.000 ;
        RECT 124.000 94.200 128.400 94.800 ;
        RECT 124.000 94.000 124.800 94.200 ;
        RECT 129.200 93.600 130.000 95.200 ;
        RECT 131.400 93.400 132.200 95.800 ;
        RECT 137.400 95.200 138.200 95.800 ;
        RECT 137.400 94.400 140.400 95.200 ;
        RECT 142.000 93.800 142.800 99.800 ;
        RECT 124.400 92.600 127.600 93.400 ;
        RECT 131.400 92.600 133.400 93.400 ;
        RECT 134.000 93.000 142.800 93.800 ;
        RECT 118.000 92.000 118.800 92.600 ;
        RECT 135.600 92.000 136.400 92.400 ;
        RECT 138.800 92.000 139.600 92.400 ;
        RECT 140.600 92.000 141.400 92.200 ;
        RECT 111.200 91.400 112.000 92.000 ;
        RECT 118.000 91.400 141.400 92.000 ;
        RECT 106.800 90.300 107.600 90.400 ;
        RECT 108.400 90.300 109.200 90.400 ;
        RECT 106.800 89.700 109.200 90.300 ;
        RECT 109.800 90.000 110.800 90.800 ;
        RECT 106.800 88.800 107.600 89.700 ;
        RECT 108.400 89.600 109.200 89.700 ;
        RECT 110.000 82.200 110.800 90.000 ;
        RECT 111.400 89.600 112.000 91.400 ;
        RECT 111.400 89.000 120.400 89.600 ;
        RECT 111.400 87.400 112.000 89.000 ;
        RECT 119.600 88.800 120.400 89.000 ;
        RECT 122.800 89.000 131.400 89.600 ;
        RECT 122.800 88.800 123.600 89.000 ;
        RECT 114.600 87.600 117.200 88.400 ;
        RECT 111.400 86.800 114.000 87.400 ;
        RECT 113.200 82.200 114.000 86.800 ;
        RECT 116.400 82.200 117.200 87.600 ;
        RECT 117.800 86.800 122.000 87.600 ;
        RECT 119.600 82.200 120.400 85.000 ;
        RECT 121.200 82.200 122.000 85.000 ;
        RECT 122.800 82.200 123.600 85.000 ;
        RECT 124.400 82.200 125.200 88.400 ;
        RECT 127.600 87.600 130.200 88.400 ;
        RECT 130.800 88.200 131.400 89.000 ;
        RECT 132.400 89.400 133.200 89.600 ;
        RECT 132.400 89.000 137.800 89.400 ;
        RECT 132.400 88.800 138.600 89.000 ;
        RECT 137.200 88.200 138.600 88.800 ;
        RECT 130.800 87.600 136.600 88.200 ;
        RECT 139.600 88.000 141.200 88.800 ;
        RECT 139.600 87.600 140.200 88.000 ;
        RECT 127.600 82.200 128.400 87.000 ;
        RECT 130.800 82.200 131.600 87.000 ;
        RECT 136.000 86.800 140.200 87.600 ;
        RECT 142.000 87.400 142.800 93.000 ;
        RECT 140.800 86.800 142.800 87.400 ;
        RECT 148.400 93.800 149.200 99.800 ;
        RECT 154.800 96.600 155.600 99.800 ;
        RECT 156.400 97.000 157.200 99.800 ;
        RECT 158.000 97.000 158.800 99.800 ;
        RECT 159.600 97.000 160.400 99.800 ;
        RECT 162.800 97.000 163.600 99.800 ;
        RECT 166.000 97.000 166.800 99.800 ;
        RECT 167.600 97.000 168.400 99.800 ;
        RECT 169.200 97.000 170.000 99.800 ;
        RECT 170.800 97.000 171.600 99.800 ;
        RECT 153.000 95.800 155.600 96.600 ;
        RECT 172.400 96.600 173.200 99.800 ;
        RECT 159.000 95.800 163.600 96.400 ;
        RECT 153.000 95.200 153.800 95.800 ;
        RECT 150.800 94.400 153.800 95.200 ;
        RECT 148.400 93.000 157.200 93.800 ;
        RECT 159.000 93.400 159.800 95.800 ;
        RECT 162.800 95.600 163.600 95.800 ;
        RECT 164.400 95.600 166.000 96.400 ;
        RECT 169.000 95.600 170.000 96.400 ;
        RECT 172.400 95.800 174.800 96.600 ;
        RECT 161.200 93.600 162.000 95.200 ;
        RECT 162.800 94.800 163.600 95.000 ;
        RECT 162.800 94.200 167.200 94.800 ;
        RECT 166.400 94.000 167.200 94.200 ;
        RECT 148.400 87.400 149.200 93.000 ;
        RECT 157.800 92.600 159.800 93.400 ;
        RECT 163.600 92.600 166.800 93.400 ;
        RECT 169.200 92.800 170.000 95.600 ;
        RECT 174.000 95.200 174.800 95.800 ;
        RECT 174.000 94.600 175.800 95.200 ;
        RECT 175.000 93.400 175.800 94.600 ;
        RECT 178.800 94.600 179.600 99.800 ;
        RECT 180.400 96.000 181.200 99.800 ;
        RECT 180.400 95.200 181.400 96.000 ;
        RECT 183.600 95.800 184.400 99.800 ;
        RECT 188.000 96.200 189.600 99.800 ;
        RECT 183.600 95.200 186.000 95.800 ;
        RECT 178.800 94.000 180.000 94.600 ;
        RECT 175.000 92.600 178.800 93.400 ;
        RECT 149.800 92.000 150.600 92.200 ;
        RECT 151.600 92.000 152.400 92.400 ;
        RECT 154.800 92.000 155.600 92.400 ;
        RECT 172.400 92.000 173.200 92.600 ;
        RECT 179.400 92.000 180.000 94.000 ;
        RECT 149.800 91.400 173.200 92.000 ;
        RECT 179.200 91.400 180.000 92.000 ;
        RECT 180.600 94.300 181.400 95.200 ;
        RECT 185.200 95.000 186.000 95.200 ;
        RECT 186.600 94.800 187.400 95.600 ;
        RECT 186.600 94.400 187.200 94.800 ;
        RECT 183.600 94.300 185.200 94.400 ;
        RECT 180.600 93.700 185.200 94.300 ;
        RECT 179.200 89.600 179.800 91.400 ;
        RECT 180.600 90.800 181.400 93.700 ;
        RECT 183.600 93.600 185.200 93.700 ;
        RECT 186.400 93.600 187.200 94.400 ;
        RECT 188.000 92.800 188.600 96.200 ;
        RECT 193.200 95.800 194.000 99.800 ;
        RECT 195.400 96.400 196.200 99.800 ;
        RECT 200.200 96.400 201.000 99.800 ;
        RECT 195.400 95.800 197.200 96.400 ;
        RECT 200.200 95.800 202.000 96.400 ;
        RECT 189.200 95.400 190.800 95.600 ;
        RECT 189.200 94.800 191.200 95.400 ;
        RECT 191.800 95.200 194.000 95.800 ;
        RECT 191.800 95.000 192.600 95.200 ;
        RECT 190.600 94.400 191.200 94.800 ;
        RECT 190.600 94.300 194.000 94.400 ;
        RECT 196.400 94.300 197.200 95.800 ;
        RECT 189.200 93.400 190.000 94.200 ;
        RECT 190.600 93.800 197.200 94.300 ;
        RECT 192.400 93.700 197.200 93.800 ;
        RECT 192.400 93.600 194.000 93.700 ;
        RECT 187.600 92.400 188.600 92.800 ;
        RECT 182.000 92.300 182.800 92.400 ;
        RECT 186.800 92.300 188.600 92.400 ;
        RECT 182.000 92.200 188.600 92.300 ;
        RECT 189.400 92.800 190.000 93.400 ;
        RECT 189.400 92.200 192.000 92.800 ;
        RECT 182.000 91.700 188.200 92.200 ;
        RECT 191.200 92.000 192.000 92.200 ;
        RECT 182.000 91.600 182.800 91.700 ;
        RECT 186.800 91.600 188.200 91.700 ;
        RECT 158.000 89.400 158.800 89.600 ;
        RECT 153.400 89.000 158.800 89.400 ;
        RECT 152.600 88.800 158.800 89.000 ;
        RECT 159.800 89.000 168.400 89.600 ;
        RECT 150.000 88.000 151.600 88.800 ;
        RECT 152.600 88.200 154.000 88.800 ;
        RECT 159.800 88.200 160.400 89.000 ;
        RECT 167.600 88.800 168.400 89.000 ;
        RECT 170.800 89.000 179.800 89.600 ;
        RECT 170.800 88.800 171.600 89.000 ;
        RECT 151.000 87.600 151.600 88.000 ;
        RECT 154.600 87.600 160.400 88.200 ;
        RECT 161.000 87.600 163.600 88.400 ;
        RECT 148.400 86.800 150.400 87.400 ;
        RECT 151.000 86.800 155.200 87.600 ;
        RECT 132.400 82.200 133.200 85.000 ;
        RECT 134.000 82.200 134.800 85.000 ;
        RECT 137.200 82.200 138.000 86.800 ;
        RECT 140.800 86.200 141.400 86.800 ;
        RECT 140.400 85.600 141.400 86.200 ;
        RECT 149.800 86.200 150.400 86.800 ;
        RECT 149.800 85.600 150.800 86.200 ;
        RECT 140.400 82.200 141.200 85.600 ;
        RECT 150.000 82.200 150.800 85.600 ;
        RECT 153.200 82.200 154.000 86.800 ;
        RECT 156.400 82.200 157.200 85.000 ;
        RECT 158.000 82.200 158.800 85.000 ;
        RECT 159.600 82.200 160.400 87.000 ;
        RECT 162.800 82.200 163.600 87.000 ;
        RECT 166.000 82.200 166.800 88.400 ;
        RECT 174.000 87.600 176.600 88.400 ;
        RECT 169.200 86.800 173.400 87.600 ;
        RECT 167.600 82.200 168.400 85.000 ;
        RECT 169.200 82.200 170.000 85.000 ;
        RECT 170.800 82.200 171.600 85.000 ;
        RECT 174.000 82.200 174.800 87.600 ;
        RECT 179.200 87.400 179.800 89.000 ;
        RECT 177.200 86.800 179.800 87.400 ;
        RECT 180.400 90.000 181.400 90.800 ;
        RECT 187.600 90.200 188.200 91.600 ;
        RECT 189.000 91.400 189.800 91.600 ;
        RECT 189.000 90.800 192.400 91.400 ;
        RECT 191.800 90.200 192.400 90.800 ;
        RECT 177.200 82.200 178.000 86.800 ;
        RECT 180.400 82.200 181.200 90.000 ;
        RECT 183.600 89.600 186.000 90.200 ;
        RECT 187.600 89.600 189.600 90.200 ;
        RECT 183.600 82.200 184.400 89.600 ;
        RECT 185.200 89.400 186.000 89.600 ;
        RECT 188.000 82.200 189.600 89.600 ;
        RECT 191.800 89.600 194.000 90.200 ;
        RECT 191.800 89.400 192.600 89.600 ;
        RECT 193.200 82.200 194.000 89.600 ;
        RECT 194.800 88.800 195.600 90.400 ;
        RECT 196.400 82.200 197.200 93.700 ;
        RECT 198.000 93.600 198.800 95.200 ;
        RECT 199.600 88.800 200.400 90.400 ;
        RECT 201.200 82.200 202.000 95.800 ;
        RECT 204.400 95.800 205.200 99.800 ;
        RECT 208.800 98.400 210.400 99.800 ;
        RECT 207.600 97.600 210.400 98.400 ;
        RECT 208.800 96.200 210.400 97.600 ;
        RECT 204.400 95.200 207.000 95.800 ;
        RECT 202.800 93.600 203.600 95.200 ;
        RECT 206.200 95.000 207.000 95.200 ;
        RECT 207.600 94.800 209.200 95.600 ;
        RECT 204.400 94.200 206.000 94.400 ;
        RECT 209.800 94.200 210.400 96.200 ;
        RECT 214.000 95.800 214.800 99.800 ;
        RECT 211.000 94.800 211.800 95.600 ;
        RECT 212.400 95.200 214.800 95.800 ;
        RECT 215.600 95.200 216.400 99.800 ;
        RECT 212.400 95.000 213.200 95.200 ;
        RECT 204.400 94.000 206.600 94.200 ;
        RECT 204.400 93.600 208.800 94.000 ;
        RECT 206.000 93.400 208.800 93.600 ;
        RECT 208.000 93.200 208.800 93.400 ;
        RECT 209.400 93.600 210.400 94.200 ;
        RECT 211.200 94.400 211.800 94.800 ;
        RECT 215.600 94.600 217.800 95.200 ;
        RECT 211.200 93.600 212.000 94.400 ;
        RECT 213.200 93.600 214.800 94.400 ;
        RECT 209.400 92.400 210.000 93.600 ;
        RECT 206.600 92.200 207.400 92.400 ;
        RECT 206.600 91.600 208.200 92.200 ;
        RECT 209.200 91.600 210.000 92.400 ;
        RECT 215.600 91.600 216.400 93.200 ;
        RECT 217.200 91.600 217.800 94.600 ;
        RECT 207.400 91.400 208.200 91.600 ;
        RECT 209.400 90.200 210.000 91.600 ;
        RECT 217.200 90.800 218.400 91.600 ;
        RECT 217.200 90.200 217.800 90.800 ;
        RECT 204.400 89.600 207.000 90.200 ;
        RECT 204.400 82.200 205.200 89.600 ;
        RECT 206.200 89.400 207.000 89.600 ;
        RECT 208.800 82.200 210.400 90.200 ;
        RECT 212.400 89.600 214.800 90.200 ;
        RECT 212.400 89.400 213.200 89.600 ;
        RECT 214.000 82.200 214.800 89.600 ;
        RECT 215.600 89.600 217.800 90.200 ;
        RECT 215.600 82.200 216.400 89.600 ;
        RECT 4.400 72.400 5.200 79.800 ;
        RECT 9.200 72.400 10.000 79.800 ;
        RECT 10.800 73.800 11.600 79.800 ;
        RECT 11.000 73.200 11.600 73.800 ;
        RECT 14.000 79.200 18.000 79.800 ;
        RECT 14.000 73.800 14.800 79.200 ;
        RECT 15.600 73.800 16.400 78.600 ;
        RECT 17.200 74.000 18.000 79.200 ;
        RECT 19.000 79.200 22.600 79.800 ;
        RECT 19.000 79.000 19.600 79.200 ;
        RECT 14.000 73.200 14.600 73.800 ;
        RECT 11.000 72.600 14.600 73.200 ;
        RECT 15.800 73.400 16.400 73.800 ;
        RECT 18.800 73.400 19.600 79.000 ;
        RECT 22.000 79.000 22.600 79.200 ;
        RECT 15.800 73.000 19.600 73.400 ;
        RECT 20.400 73.000 21.200 78.600 ;
        RECT 22.000 73.000 22.800 79.000 ;
        RECT 15.800 72.800 19.400 73.000 ;
        RECT 3.000 71.800 5.200 72.400 ;
        RECT 7.800 71.800 10.000 72.400 ;
        RECT 20.400 72.400 21.000 73.000 ;
        RECT 26.200 72.400 27.000 79.800 ;
        RECT 27.600 73.600 28.400 74.400 ;
        RECT 30.000 74.300 30.800 74.400 ;
        RECT 31.600 74.300 32.400 79.800 ;
        RECT 30.000 73.700 32.400 74.300 ;
        RECT 30.000 73.600 30.800 73.700 ;
        RECT 27.800 72.400 28.400 73.600 ;
        RECT 20.400 72.200 21.200 72.400 ;
        RECT 3.000 71.200 3.600 71.800 ;
        RECT 7.800 71.200 8.400 71.800 ;
        RECT 2.400 70.400 3.600 71.200 ;
        RECT 7.200 70.400 8.400 71.200 ;
        RECT 17.800 71.600 21.200 72.200 ;
        RECT 26.200 71.800 27.200 72.400 ;
        RECT 27.800 71.800 29.200 72.400 ;
        RECT 3.000 67.400 3.600 70.400 ;
        RECT 4.400 68.800 5.200 70.400 ;
        RECT 7.800 67.400 8.400 70.400 ;
        RECT 9.200 68.800 10.000 70.400 ;
        RECT 15.600 69.600 17.200 70.400 ;
        RECT 10.800 68.300 11.600 68.400 ;
        RECT 14.000 68.300 15.600 68.400 ;
        RECT 10.800 67.700 15.600 68.300 ;
        RECT 10.800 67.600 11.600 67.700 ;
        RECT 14.000 67.600 15.600 67.700 ;
        RECT 3.000 66.800 5.200 67.400 ;
        RECT 7.800 66.800 10.000 67.400 ;
        RECT 4.400 62.200 5.200 66.800 ;
        RECT 9.200 62.200 10.000 66.800 ;
        RECT 12.400 66.300 14.200 66.400 ;
        RECT 15.600 66.300 16.400 66.400 ;
        RECT 12.400 65.700 16.400 66.300 ;
        RECT 12.400 65.600 14.200 65.700 ;
        RECT 15.600 65.600 16.400 65.700 ;
        RECT 17.800 65.000 18.400 71.600 ;
        RECT 25.200 68.800 26.000 70.400 ;
        RECT 26.600 68.400 27.200 71.800 ;
        RECT 28.400 71.600 29.200 71.800 ;
        RECT 23.600 68.200 24.400 68.400 ;
        RECT 26.600 68.300 29.200 68.400 ;
        RECT 30.000 68.300 30.800 68.400 ;
        RECT 23.600 67.600 25.200 68.200 ;
        RECT 26.600 67.700 30.800 68.300 ;
        RECT 26.600 67.600 29.200 67.700 ;
        RECT 24.400 67.200 25.200 67.600 ;
        RECT 23.800 66.200 27.400 66.600 ;
        RECT 28.400 66.200 29.000 67.600 ;
        RECT 30.000 66.800 30.800 67.700 ;
        RECT 31.600 66.200 32.400 73.700 ;
        RECT 33.200 71.600 34.000 73.200 ;
        RECT 34.800 72.400 35.600 79.800 ;
        RECT 36.200 72.400 37.000 72.600 ;
        RECT 34.800 71.800 37.000 72.400 ;
        RECT 39.200 72.400 40.800 79.800 ;
        RECT 42.800 72.400 43.600 72.600 ;
        RECT 44.400 72.400 45.200 79.800 ;
        RECT 39.200 71.800 41.200 72.400 ;
        RECT 42.800 71.800 45.200 72.400 ;
        RECT 52.400 72.000 53.200 79.800 ;
        RECT 55.600 75.200 56.400 79.800 ;
        RECT 36.400 71.200 37.000 71.800 ;
        RECT 36.400 70.600 39.800 71.200 ;
        RECT 39.000 70.400 39.800 70.600 ;
        RECT 40.600 70.400 41.200 71.800 ;
        RECT 52.200 71.200 53.200 72.000 ;
        RECT 53.800 74.600 56.400 75.200 ;
        RECT 53.800 73.000 54.400 74.600 ;
        RECT 58.800 74.400 59.600 79.800 ;
        RECT 62.000 77.000 62.800 79.800 ;
        RECT 63.600 77.000 64.400 79.800 ;
        RECT 65.200 77.000 66.000 79.800 ;
        RECT 60.200 74.400 64.400 75.200 ;
        RECT 57.000 73.600 59.600 74.400 ;
        RECT 66.800 73.600 67.600 79.800 ;
        RECT 70.000 75.000 70.800 79.800 ;
        RECT 73.200 75.000 74.000 79.800 ;
        RECT 74.800 77.000 75.600 79.800 ;
        RECT 76.400 77.000 77.200 79.800 ;
        RECT 79.600 75.200 80.400 79.800 ;
        RECT 82.800 76.400 83.600 79.800 ;
        RECT 82.800 75.800 83.800 76.400 ;
        RECT 83.200 75.200 83.800 75.800 ;
        RECT 78.400 74.400 82.600 75.200 ;
        RECT 83.200 74.600 85.200 75.200 ;
        RECT 70.000 73.600 72.600 74.400 ;
        RECT 73.200 73.800 79.000 74.400 ;
        RECT 82.000 74.000 82.600 74.400 ;
        RECT 62.000 73.000 62.800 73.200 ;
        RECT 53.800 72.400 62.800 73.000 ;
        RECT 65.200 73.000 66.000 73.200 ;
        RECT 73.200 73.000 73.800 73.800 ;
        RECT 79.600 73.200 81.000 73.800 ;
        RECT 82.000 73.200 83.600 74.000 ;
        RECT 65.200 72.400 73.800 73.000 ;
        RECT 74.800 73.000 81.000 73.200 ;
        RECT 74.800 72.600 80.200 73.000 ;
        RECT 74.800 72.400 75.600 72.600 ;
        RECT 40.600 70.300 42.000 70.400 ;
        RECT 50.800 70.300 51.600 70.400 ;
        RECT 36.800 69.800 37.600 70.000 ;
        RECT 40.600 69.800 51.600 70.300 ;
        RECT 36.800 69.200 39.400 69.800 ;
        RECT 38.800 68.600 39.400 69.200 ;
        RECT 40.200 69.700 51.600 69.800 ;
        RECT 40.200 69.600 42.000 69.700 ;
        RECT 50.800 69.600 51.600 69.700 ;
        RECT 40.200 69.200 41.200 69.600 ;
        RECT 34.800 68.200 36.400 68.400 ;
        RECT 34.800 67.600 38.200 68.200 ;
        RECT 38.800 67.800 39.600 68.600 ;
        RECT 37.600 67.200 38.200 67.600 ;
        RECT 36.200 66.800 37.000 67.000 ;
        RECT 34.800 66.200 37.000 66.800 ;
        RECT 37.600 66.600 39.600 67.200 ;
        RECT 38.000 66.400 39.600 66.600 ;
        RECT 14.400 64.400 18.400 65.000 ;
        RECT 14.000 63.600 15.000 64.400 ;
        RECT 17.200 64.200 18.400 64.400 ;
        RECT 23.600 66.000 27.600 66.200 ;
        RECT 14.000 62.200 14.800 63.600 ;
        RECT 17.200 62.200 18.000 64.200 ;
        RECT 23.600 62.200 24.400 66.000 ;
        RECT 26.800 62.200 27.600 66.000 ;
        RECT 28.400 62.200 29.200 66.200 ;
        RECT 31.600 65.600 33.400 66.200 ;
        RECT 32.600 62.200 33.400 65.600 ;
        RECT 34.800 62.200 35.600 66.200 ;
        RECT 40.200 65.800 40.800 69.200 ;
        RECT 41.600 67.600 42.400 68.400 ;
        RECT 43.600 68.300 45.200 68.400 ;
        RECT 52.200 68.300 53.000 71.200 ;
        RECT 53.800 70.600 54.400 72.400 ;
        RECT 77.800 71.800 78.800 72.000 ;
        RECT 81.200 71.800 82.000 72.400 ;
        RECT 55.000 71.200 82.000 71.800 ;
        RECT 55.000 71.000 55.800 71.200 ;
        RECT 43.600 67.700 53.000 68.300 ;
        RECT 43.600 67.600 45.200 67.700 ;
        RECT 41.600 67.200 42.200 67.600 ;
        RECT 41.400 66.400 42.200 67.200 ;
        RECT 42.800 66.800 43.600 67.000 ;
        RECT 52.200 66.800 53.000 67.700 ;
        RECT 53.600 70.000 54.400 70.600 ;
        RECT 53.600 68.000 54.200 70.000 ;
        RECT 54.800 68.600 58.600 69.400 ;
        RECT 53.600 67.400 54.800 68.000 ;
        RECT 42.800 66.200 45.200 66.800 ;
        RECT 39.200 62.200 40.800 65.800 ;
        RECT 44.400 62.200 45.200 66.200 ;
        RECT 52.200 66.000 53.200 66.800 ;
        RECT 52.400 62.200 53.200 66.000 ;
        RECT 54.000 62.200 54.800 67.400 ;
        RECT 57.800 67.400 58.600 68.600 ;
        RECT 57.800 66.800 59.600 67.400 ;
        RECT 58.800 66.200 59.600 66.800 ;
        RECT 63.600 66.400 64.400 69.200 ;
        RECT 66.800 68.600 70.000 69.400 ;
        RECT 73.800 68.600 75.800 69.400 ;
        RECT 84.400 69.000 85.200 74.600 ;
        RECT 66.400 67.800 67.200 68.000 ;
        RECT 66.400 67.200 70.800 67.800 ;
        RECT 70.000 67.000 70.800 67.200 ;
        RECT 71.600 66.800 72.400 68.400 ;
        RECT 58.800 65.400 61.200 66.200 ;
        RECT 63.600 65.600 64.600 66.400 ;
        RECT 67.600 65.600 69.200 66.400 ;
        RECT 70.000 66.200 70.800 66.400 ;
        RECT 73.800 66.200 74.600 68.600 ;
        RECT 76.400 68.200 85.200 69.000 ;
        RECT 79.800 66.800 82.800 67.600 ;
        RECT 79.800 66.200 80.600 66.800 ;
        RECT 70.000 65.600 74.600 66.200 ;
        RECT 60.400 62.200 61.200 65.400 ;
        RECT 78.000 65.400 80.600 66.200 ;
        RECT 62.000 62.200 62.800 65.000 ;
        RECT 63.600 62.200 64.400 65.000 ;
        RECT 65.200 62.200 66.000 65.000 ;
        RECT 66.800 62.200 67.600 65.000 ;
        RECT 70.000 62.200 70.800 65.000 ;
        RECT 73.200 62.200 74.000 65.000 ;
        RECT 74.800 62.200 75.600 65.000 ;
        RECT 76.400 62.200 77.200 65.000 ;
        RECT 78.000 62.200 78.800 65.400 ;
        RECT 84.400 62.200 85.200 68.200 ;
        RECT 86.000 62.200 86.800 79.800 ;
        RECT 90.800 71.200 91.600 79.800 ;
        RECT 94.000 71.200 94.800 79.800 ;
        RECT 97.200 71.200 98.000 79.800 ;
        RECT 100.400 71.200 101.200 79.800 ;
        RECT 105.200 75.800 106.000 79.800 ;
        RECT 105.400 75.600 106.000 75.800 ;
        RECT 108.400 75.800 109.200 79.800 ;
        RECT 108.400 75.600 109.000 75.800 ;
        RECT 105.400 75.000 109.000 75.600 ;
        RECT 105.200 74.300 106.000 74.400 ;
        RECT 106.800 74.300 107.600 74.400 ;
        RECT 105.200 73.700 107.600 74.300 ;
        RECT 105.200 73.600 106.000 73.700 ;
        RECT 106.800 72.800 107.600 73.700 ;
        RECT 108.400 72.400 109.000 75.000 ;
        RECT 89.200 70.400 91.600 71.200 ;
        RECT 92.600 70.400 94.800 71.200 ;
        RECT 95.800 70.400 98.000 71.200 ;
        RECT 99.400 70.400 101.200 71.200 ;
        RECT 103.600 70.800 104.400 72.400 ;
        RECT 108.400 71.600 109.200 72.400 ;
        RECT 89.200 67.600 90.000 70.400 ;
        RECT 92.600 69.000 93.400 70.400 ;
        RECT 95.800 69.000 96.600 70.400 ;
        RECT 99.400 69.000 100.200 70.400 ;
        RECT 105.200 69.600 106.800 70.400 ;
        RECT 90.800 68.200 93.400 69.000 ;
        RECT 94.200 68.200 96.600 69.000 ;
        RECT 97.600 68.200 100.200 69.000 ;
        RECT 108.400 68.400 109.000 71.600 ;
        RECT 110.000 70.300 110.800 70.400 ;
        RECT 111.600 70.300 112.400 79.800 ;
        RECT 114.800 71.200 115.600 79.800 ;
        RECT 118.000 71.200 118.800 79.800 ;
        RECT 121.200 71.200 122.000 79.800 ;
        RECT 124.400 71.200 125.200 79.800 ;
        RECT 127.600 72.400 128.400 79.800 ;
        RECT 130.800 72.800 131.600 79.800 ;
        RECT 127.600 71.800 130.200 72.400 ;
        RECT 130.800 71.800 131.800 72.800 ;
        RECT 110.000 69.700 112.400 70.300 ;
        RECT 110.000 69.600 110.800 69.700 ;
        RECT 107.400 68.200 109.000 68.400 ;
        RECT 92.600 67.600 93.400 68.200 ;
        RECT 95.800 67.600 96.600 68.200 ;
        RECT 99.400 67.600 100.200 68.200 ;
        RECT 107.200 67.800 109.000 68.200 ;
        RECT 89.200 66.800 91.600 67.600 ;
        RECT 92.600 66.800 94.800 67.600 ;
        RECT 95.800 66.800 98.000 67.600 ;
        RECT 99.400 66.800 101.200 67.600 ;
        RECT 87.600 64.800 88.400 66.400 ;
        RECT 90.800 62.200 91.600 66.800 ;
        RECT 94.000 62.200 94.800 66.800 ;
        RECT 97.200 62.200 98.000 66.800 ;
        RECT 100.400 62.200 101.200 66.800 ;
        RECT 107.200 62.200 108.000 67.800 ;
        RECT 110.000 64.800 110.800 66.400 ;
        RECT 111.600 62.200 112.400 69.700 ;
        RECT 113.200 70.400 115.600 71.200 ;
        RECT 116.600 70.400 118.800 71.200 ;
        RECT 119.800 70.400 122.000 71.200 ;
        RECT 123.400 70.400 125.200 71.200 ;
        RECT 113.200 67.600 114.000 70.400 ;
        RECT 116.600 69.000 117.400 70.400 ;
        RECT 119.800 69.000 120.600 70.400 ;
        RECT 123.400 69.000 124.200 70.400 ;
        RECT 127.600 69.600 128.600 70.400 ;
        RECT 114.800 68.200 117.400 69.000 ;
        RECT 118.200 68.200 120.600 69.000 ;
        RECT 121.600 68.200 124.200 69.000 ;
        RECT 127.800 68.800 128.600 69.600 ;
        RECT 129.600 69.800 130.200 71.800 ;
        RECT 129.600 69.000 130.600 69.800 ;
        RECT 116.600 67.600 117.400 68.200 ;
        RECT 119.800 67.600 120.600 68.200 ;
        RECT 123.400 67.600 124.200 68.200 ;
        RECT 113.200 66.800 115.600 67.600 ;
        RECT 116.600 66.800 118.800 67.600 ;
        RECT 119.800 66.800 122.000 67.600 ;
        RECT 123.400 66.800 125.200 67.600 ;
        RECT 129.600 67.400 130.200 69.000 ;
        RECT 131.200 68.400 131.800 71.800 ;
        RECT 135.600 71.200 136.400 79.800 ;
        RECT 138.800 71.200 139.600 79.800 ;
        RECT 142.000 71.200 142.800 79.800 ;
        RECT 145.200 71.200 146.000 79.800 ;
        RECT 151.000 72.600 151.800 79.800 ;
        RECT 150.000 71.800 151.800 72.600 ;
        RECT 158.600 72.600 159.400 79.800 ;
        RECT 164.400 75.800 165.200 79.800 ;
        RECT 158.600 71.800 160.400 72.600 ;
        RECT 135.600 70.400 137.400 71.200 ;
        RECT 138.800 70.400 141.000 71.200 ;
        RECT 142.000 70.400 144.200 71.200 ;
        RECT 145.200 70.400 147.600 71.200 ;
        RECT 130.800 67.600 131.800 68.400 ;
        RECT 136.600 69.000 137.400 70.400 ;
        RECT 140.200 69.000 141.000 70.400 ;
        RECT 143.400 69.000 144.200 70.400 ;
        RECT 136.600 68.200 139.200 69.000 ;
        RECT 140.200 68.200 142.600 69.000 ;
        RECT 143.400 68.200 146.000 69.000 ;
        RECT 136.600 67.600 137.400 68.200 ;
        RECT 140.200 67.600 141.000 68.200 ;
        RECT 143.400 67.600 144.200 68.200 ;
        RECT 146.800 67.600 147.600 70.400 ;
        RECT 150.200 68.400 150.800 71.800 ;
        RECT 151.600 69.600 152.400 71.200 ;
        RECT 158.000 69.600 158.800 71.200 ;
        RECT 150.000 67.600 150.800 68.400 ;
        RECT 114.800 62.200 115.600 66.800 ;
        RECT 118.000 62.200 118.800 66.800 ;
        RECT 121.200 62.200 122.000 66.800 ;
        RECT 124.400 62.200 125.200 66.800 ;
        RECT 127.600 66.800 130.200 67.400 ;
        RECT 127.600 62.200 128.400 66.800 ;
        RECT 131.200 66.200 131.800 67.600 ;
        RECT 130.800 65.600 131.800 66.200 ;
        RECT 135.600 66.800 137.400 67.600 ;
        RECT 138.800 66.800 141.000 67.600 ;
        RECT 142.000 66.800 144.200 67.600 ;
        RECT 145.200 66.800 147.600 67.600 ;
        RECT 130.800 62.200 131.600 65.600 ;
        RECT 135.600 62.200 136.400 66.800 ;
        RECT 138.800 62.200 139.600 66.800 ;
        RECT 142.000 62.200 142.800 66.800 ;
        RECT 145.200 62.200 146.000 66.800 ;
        RECT 148.400 64.800 149.200 66.400 ;
        RECT 150.200 64.400 150.800 67.600 ;
        RECT 159.600 68.400 160.200 71.800 ;
        RECT 164.600 71.600 165.200 75.800 ;
        RECT 167.600 71.800 168.400 79.800 ;
        RECT 169.200 72.400 170.000 79.800 ;
        RECT 174.000 72.400 174.800 79.800 ;
        RECT 175.800 72.400 176.600 72.600 ;
        RECT 169.200 71.800 171.400 72.400 ;
        RECT 174.000 71.800 176.600 72.400 ;
        RECT 178.400 71.800 180.000 79.800 ;
        RECT 182.000 72.400 182.800 72.600 ;
        RECT 183.600 72.400 184.400 79.800 ;
        RECT 186.800 75.800 187.600 79.800 ;
        RECT 182.000 71.800 184.400 72.400 ;
        RECT 164.600 71.000 167.000 71.600 ;
        RECT 164.400 69.600 165.200 70.400 ;
        RECT 159.600 67.600 160.400 68.400 ;
        RECT 162.800 67.600 163.600 69.200 ;
        RECT 164.600 68.800 165.200 69.600 ;
        RECT 164.600 68.200 165.600 68.800 ;
        RECT 164.800 68.000 165.600 68.200 ;
        RECT 166.400 67.600 167.000 71.000 ;
        RECT 167.800 70.400 168.400 71.800 ;
        RECT 170.800 71.200 171.400 71.800 ;
        RECT 170.800 70.400 172.000 71.200 ;
        RECT 177.000 70.400 177.800 70.600 ;
        RECT 179.000 70.400 179.600 71.800 ;
        RECT 187.000 71.600 187.600 75.800 ;
        RECT 190.000 71.800 190.800 79.800 ;
        RECT 187.000 71.000 189.400 71.600 ;
        RECT 167.600 69.600 168.400 70.400 ;
        RECT 151.600 66.300 152.400 66.400 ;
        RECT 159.600 66.300 160.200 67.600 ;
        RECT 166.400 67.400 167.200 67.600 ;
        RECT 164.200 67.000 167.200 67.400 ;
        RECT 163.000 66.800 167.200 67.000 ;
        RECT 163.000 66.400 164.800 66.800 ;
        RECT 151.600 65.700 160.300 66.300 ;
        RECT 151.600 65.600 152.400 65.700 ;
        RECT 150.000 62.200 150.800 64.400 ;
        RECT 159.600 64.200 160.200 65.700 ;
        RECT 161.200 64.800 162.000 66.400 ;
        RECT 163.000 66.200 163.600 66.400 ;
        RECT 167.800 66.200 168.400 69.600 ;
        RECT 169.200 68.800 170.000 70.400 ;
        RECT 170.800 67.400 171.400 70.400 ;
        RECT 176.200 69.800 177.800 70.400 ;
        RECT 176.200 69.600 177.000 69.800 ;
        RECT 178.800 69.600 179.600 70.400 ;
        RECT 186.800 69.600 187.600 70.400 ;
        RECT 177.600 68.600 178.400 68.800 ;
        RECT 175.600 68.400 178.400 68.600 ;
        RECT 174.000 68.000 178.400 68.400 ;
        RECT 179.000 68.400 179.600 69.600 ;
        RECT 174.000 67.800 176.200 68.000 ;
        RECT 179.000 67.800 180.000 68.400 ;
        RECT 174.000 67.600 175.600 67.800 ;
        RECT 159.600 62.200 160.400 64.200 ;
        RECT 162.800 62.200 163.600 66.200 ;
        RECT 167.000 65.200 168.400 66.200 ;
        RECT 169.200 66.800 171.400 67.400 ;
        RECT 175.800 66.800 176.600 67.000 ;
        RECT 167.000 62.200 167.800 65.200 ;
        RECT 169.200 62.200 170.000 66.800 ;
        RECT 174.000 66.200 176.600 66.800 ;
        RECT 177.200 66.400 178.800 67.200 ;
        RECT 174.000 62.200 174.800 66.200 ;
        RECT 179.400 65.800 180.000 67.800 ;
        RECT 180.800 67.600 181.600 68.400 ;
        RECT 182.800 67.600 184.400 68.400 ;
        RECT 185.200 67.600 186.000 69.200 ;
        RECT 187.000 68.800 187.600 69.600 ;
        RECT 187.000 68.200 188.000 68.800 ;
        RECT 187.200 68.000 188.000 68.200 ;
        RECT 188.800 67.600 189.400 71.000 ;
        RECT 190.200 70.400 190.800 71.800 ;
        RECT 190.000 69.600 190.800 70.400 ;
        RECT 180.800 67.200 181.400 67.600 ;
        RECT 188.800 67.400 189.600 67.600 ;
        RECT 180.600 66.400 181.400 67.200 ;
        RECT 186.600 67.000 189.600 67.400 ;
        RECT 182.000 66.800 182.800 67.000 ;
        RECT 185.400 66.800 189.600 67.000 ;
        RECT 182.000 66.200 184.400 66.800 ;
        RECT 185.400 66.400 187.200 66.800 ;
        RECT 185.400 66.200 186.000 66.400 ;
        RECT 190.200 66.200 190.800 69.600 ;
        RECT 178.400 64.400 180.000 65.800 ;
        RECT 177.200 63.600 180.000 64.400 ;
        RECT 178.400 62.200 180.000 63.600 ;
        RECT 183.600 62.200 184.400 66.200 ;
        RECT 185.200 62.200 186.000 66.200 ;
        RECT 189.400 65.200 190.800 66.200 ;
        RECT 191.600 71.800 192.400 79.800 ;
        RECT 194.800 75.800 195.600 79.800 ;
        RECT 191.600 70.400 192.200 71.800 ;
        RECT 194.800 71.600 195.400 75.800 ;
        RECT 198.600 72.600 199.400 79.800 ;
        RECT 205.400 78.400 206.200 79.800 ;
        RECT 204.400 77.600 206.200 78.400 ;
        RECT 205.400 72.600 206.200 77.600 ;
        RECT 198.600 71.800 200.400 72.600 ;
        RECT 204.400 71.800 206.200 72.600 ;
        RECT 193.000 71.000 195.400 71.600 ;
        RECT 199.600 71.600 200.400 71.800 ;
        RECT 191.600 69.600 192.400 70.400 ;
        RECT 191.600 66.200 192.200 69.600 ;
        RECT 193.000 67.600 193.600 71.000 ;
        RECT 194.800 69.600 195.600 70.400 ;
        RECT 198.000 69.600 198.800 71.200 ;
        RECT 194.800 68.800 195.400 69.600 ;
        RECT 194.400 68.200 195.400 68.800 ;
        RECT 194.400 68.000 195.200 68.200 ;
        RECT 196.400 67.600 197.200 69.200 ;
        RECT 199.600 68.400 200.200 71.600 ;
        RECT 204.600 68.400 205.200 71.800 ;
        RECT 206.000 70.300 206.800 71.200 ;
        RECT 207.600 70.300 208.400 79.800 ;
        RECT 210.800 72.400 211.600 79.800 ;
        RECT 210.800 71.800 213.000 72.400 ;
        RECT 212.400 71.200 213.000 71.800 ;
        RECT 212.400 70.400 213.600 71.200 ;
        RECT 206.000 69.700 208.400 70.300 ;
        RECT 206.000 69.600 206.800 69.700 ;
        RECT 199.600 67.600 200.400 68.400 ;
        RECT 204.400 67.600 205.200 68.400 ;
        RECT 192.800 67.400 193.600 67.600 ;
        RECT 192.800 67.000 195.800 67.400 ;
        RECT 192.800 66.800 197.000 67.000 ;
        RECT 195.200 66.400 197.000 66.800 ;
        RECT 196.400 66.200 197.000 66.400 ;
        RECT 191.600 65.200 193.000 66.200 ;
        RECT 189.400 62.200 190.200 65.200 ;
        RECT 192.200 62.200 193.000 65.200 ;
        RECT 196.400 62.200 197.200 66.200 ;
        RECT 199.600 64.200 200.200 67.600 ;
        RECT 201.200 66.300 202.000 66.400 ;
        RECT 202.800 66.300 203.600 66.400 ;
        RECT 201.200 65.700 203.600 66.300 ;
        RECT 201.200 64.800 202.000 65.700 ;
        RECT 202.800 64.800 203.600 65.700 ;
        RECT 204.600 64.400 205.200 67.600 ;
        RECT 199.600 62.200 200.400 64.200 ;
        RECT 204.400 62.200 205.200 64.400 ;
        RECT 207.600 62.200 208.400 69.700 ;
        RECT 210.800 68.800 211.600 70.400 ;
        RECT 212.400 67.400 213.000 70.400 ;
        RECT 210.800 66.800 213.000 67.400 ;
        RECT 209.200 64.800 210.000 66.400 ;
        RECT 210.800 62.200 211.600 66.800 ;
        RECT 2.800 56.000 3.600 59.800 ;
        RECT 2.600 55.200 3.600 56.000 ;
        RECT 2.600 50.800 3.400 55.200 ;
        RECT 4.400 54.600 5.200 59.800 ;
        RECT 10.800 56.600 11.600 59.800 ;
        RECT 12.400 57.000 13.200 59.800 ;
        RECT 14.000 57.000 14.800 59.800 ;
        RECT 15.600 57.000 16.400 59.800 ;
        RECT 17.200 57.000 18.000 59.800 ;
        RECT 20.400 57.000 21.200 59.800 ;
        RECT 23.600 57.000 24.400 59.800 ;
        RECT 25.200 57.000 26.000 59.800 ;
        RECT 26.800 57.000 27.600 59.800 ;
        RECT 9.200 55.800 11.600 56.600 ;
        RECT 28.400 56.600 29.200 59.800 ;
        RECT 9.200 55.200 10.000 55.800 ;
        RECT 4.000 54.000 5.200 54.600 ;
        RECT 8.200 54.600 10.000 55.200 ;
        RECT 14.000 55.600 15.000 56.400 ;
        RECT 18.000 55.600 19.600 56.400 ;
        RECT 20.400 55.800 25.000 56.400 ;
        RECT 28.400 55.800 31.000 56.600 ;
        RECT 20.400 55.600 21.200 55.800 ;
        RECT 4.000 52.000 4.600 54.000 ;
        RECT 8.200 53.400 9.000 54.600 ;
        RECT 5.200 52.600 9.000 53.400 ;
        RECT 14.000 52.800 14.800 55.600 ;
        RECT 20.400 54.800 21.200 55.000 ;
        RECT 16.800 54.200 21.200 54.800 ;
        RECT 16.800 54.000 17.600 54.200 ;
        RECT 22.000 53.600 22.800 55.200 ;
        RECT 24.200 53.400 25.000 55.800 ;
        RECT 30.200 55.200 31.000 55.800 ;
        RECT 30.200 54.400 33.200 55.200 ;
        RECT 34.800 53.800 35.600 59.800 ;
        RECT 37.000 56.400 37.800 59.800 ;
        RECT 37.000 55.800 38.800 56.400 ;
        RECT 17.200 52.600 20.400 53.400 ;
        RECT 24.200 52.600 26.200 53.400 ;
        RECT 26.800 53.000 35.600 53.800 ;
        RECT 36.400 54.300 37.200 54.400 ;
        RECT 38.000 54.300 38.800 55.800 ;
        RECT 41.200 55.600 42.000 57.200 ;
        RECT 36.400 53.700 38.800 54.300 ;
        RECT 36.400 53.600 37.200 53.700 ;
        RECT 4.000 51.400 4.800 52.000 ;
        RECT 2.600 50.000 3.600 50.800 ;
        RECT 2.800 42.200 3.600 50.000 ;
        RECT 4.200 49.600 4.800 51.400 ;
        RECT 5.400 50.800 6.200 51.000 ;
        RECT 5.400 50.200 32.400 50.800 ;
        RECT 28.200 50.000 29.000 50.200 ;
        RECT 31.600 49.600 32.400 50.200 ;
        RECT 4.200 49.000 13.200 49.600 ;
        RECT 4.200 47.400 4.800 49.000 ;
        RECT 12.400 48.800 13.200 49.000 ;
        RECT 15.600 49.000 24.200 49.600 ;
        RECT 15.600 48.800 16.400 49.000 ;
        RECT 7.400 47.600 10.000 48.400 ;
        RECT 4.200 46.800 6.800 47.400 ;
        RECT 6.000 42.200 6.800 46.800 ;
        RECT 9.200 42.200 10.000 47.600 ;
        RECT 10.600 46.800 14.800 47.600 ;
        RECT 12.400 42.200 13.200 45.000 ;
        RECT 14.000 42.200 14.800 45.000 ;
        RECT 15.600 42.200 16.400 45.000 ;
        RECT 17.200 42.200 18.000 48.400 ;
        RECT 20.400 47.600 23.000 48.400 ;
        RECT 23.600 48.200 24.200 49.000 ;
        RECT 25.200 49.400 26.000 49.600 ;
        RECT 25.200 49.000 30.600 49.400 ;
        RECT 25.200 48.800 31.400 49.000 ;
        RECT 30.000 48.200 31.400 48.800 ;
        RECT 23.600 47.600 29.400 48.200 ;
        RECT 32.400 48.000 34.000 48.800 ;
        RECT 32.400 47.600 33.000 48.000 ;
        RECT 20.400 42.200 21.200 47.000 ;
        RECT 23.600 42.200 24.400 47.000 ;
        RECT 28.800 46.800 33.000 47.600 ;
        RECT 34.800 47.400 35.600 53.000 ;
        RECT 36.400 48.800 37.200 50.400 ;
        RECT 33.600 46.800 35.600 47.400 ;
        RECT 25.200 42.200 26.000 45.000 ;
        RECT 26.800 42.200 27.600 45.000 ;
        RECT 30.000 42.200 30.800 46.800 ;
        RECT 33.600 46.200 34.200 46.800 ;
        RECT 33.200 45.600 34.200 46.200 ;
        RECT 33.200 42.200 34.000 45.600 ;
        RECT 38.000 42.200 38.800 53.700 ;
        RECT 39.600 53.600 40.400 55.200 ;
        RECT 42.800 50.300 43.600 59.800 ;
        RECT 48.000 54.200 48.800 59.800 ;
        RECT 50.800 55.800 51.600 59.800 ;
        RECT 52.400 56.000 53.200 59.800 ;
        RECT 55.600 56.000 56.400 59.800 ;
        RECT 65.200 58.400 66.000 59.800 ;
        RECT 65.200 57.800 66.200 58.400 ;
        RECT 65.600 57.600 66.200 57.800 ;
        RECT 68.400 57.800 69.200 59.800 ;
        RECT 68.400 57.600 69.600 57.800 ;
        RECT 65.600 57.000 69.600 57.600 ;
        RECT 52.400 55.800 56.400 56.000 ;
        RECT 51.000 54.400 51.600 55.800 ;
        RECT 52.600 55.400 56.200 55.800 ;
        RECT 63.600 55.600 65.400 56.400 ;
        RECT 54.800 54.400 55.600 54.800 ;
        RECT 48.000 53.800 49.800 54.200 ;
        RECT 48.200 53.600 49.800 53.800 ;
        RECT 50.800 53.600 53.400 54.400 ;
        RECT 54.800 54.300 56.400 54.400 ;
        RECT 63.700 54.300 64.300 55.600 ;
        RECT 54.800 53.800 64.300 54.300 ;
        RECT 55.600 53.700 64.300 53.800 ;
        RECT 55.600 53.600 56.400 53.700 ;
        RECT 65.200 53.600 66.800 54.400 ;
        RECT 46.000 51.600 47.600 52.400 ;
        RECT 44.400 50.300 45.200 51.200 ;
        RECT 42.800 49.700 45.200 50.300 ;
        RECT 42.800 42.200 43.600 49.700 ;
        RECT 44.400 49.600 45.200 49.700 ;
        RECT 49.200 50.400 49.800 53.600 ;
        RECT 52.800 52.400 53.400 53.600 ;
        RECT 52.400 51.600 53.400 52.400 ;
        RECT 54.000 52.300 54.800 53.200 ;
        RECT 66.800 52.300 68.400 52.400 ;
        RECT 54.000 51.700 68.400 52.300 ;
        RECT 54.000 51.600 54.800 51.700 ;
        RECT 66.800 51.600 68.400 51.700 ;
        RECT 49.200 49.600 50.000 50.400 ;
        RECT 50.800 50.200 51.600 50.400 ;
        RECT 52.800 50.200 53.400 51.600 ;
        RECT 69.000 50.400 69.600 57.000 ;
        RECT 73.200 56.300 74.000 56.400 ;
        RECT 74.800 56.300 75.600 57.200 ;
        RECT 73.200 55.700 75.600 56.300 ;
        RECT 73.200 55.600 74.000 55.700 ;
        RECT 74.800 55.600 75.600 55.700 ;
        RECT 50.800 49.600 52.200 50.200 ;
        RECT 52.800 49.600 53.800 50.200 ;
        RECT 69.000 49.800 72.400 50.400 ;
        RECT 47.600 47.600 48.400 49.200 ;
        RECT 49.200 47.000 49.800 49.600 ;
        RECT 51.600 48.400 52.200 49.600 ;
        RECT 50.800 47.600 52.400 48.400 ;
        RECT 46.200 46.400 49.800 47.000 ;
        RECT 46.200 46.200 46.800 46.400 ;
        RECT 46.000 42.200 46.800 46.200 ;
        RECT 49.200 46.200 49.800 46.400 ;
        RECT 49.200 42.200 50.000 46.200 ;
        RECT 53.000 42.200 53.800 49.600 ;
        RECT 71.600 49.600 72.400 49.800 ;
        RECT 76.400 50.300 77.200 59.800 ;
        RECT 81.600 58.400 82.400 59.800 ;
        RECT 81.600 57.600 83.600 58.400 ;
        RECT 89.200 57.800 90.000 59.800 ;
        RECT 92.400 58.400 93.200 59.800 ;
        RECT 88.800 57.600 90.000 57.800 ;
        RECT 92.200 57.600 93.200 58.400 ;
        RECT 81.600 54.200 82.400 57.600 ;
        RECT 88.800 57.000 92.800 57.600 ;
        RECT 81.600 53.800 83.400 54.200 ;
        RECT 81.800 53.600 83.400 53.800 ;
        RECT 79.600 51.600 81.200 52.400 ;
        RECT 78.000 50.300 78.800 51.200 ;
        RECT 76.400 49.700 78.800 50.300 ;
        RECT 62.200 48.800 65.800 49.400 ;
        RECT 62.200 48.200 62.800 48.800 ;
        RECT 62.000 42.200 62.800 48.200 ;
        RECT 65.200 48.200 65.800 48.800 ;
        RECT 67.000 49.000 70.600 49.200 ;
        RECT 71.600 49.000 72.200 49.600 ;
        RECT 67.000 48.600 70.800 49.000 ;
        RECT 67.000 48.200 67.600 48.600 ;
        RECT 65.200 42.800 66.000 48.200 ;
        RECT 66.800 43.400 67.600 48.200 ;
        RECT 68.400 42.800 69.200 48.000 ;
        RECT 70.000 43.000 70.800 48.600 ;
        RECT 71.600 43.400 72.400 49.000 ;
        RECT 65.200 42.200 69.200 42.800 ;
        RECT 70.200 42.800 70.800 43.000 ;
        RECT 73.200 43.000 74.000 49.000 ;
        RECT 73.200 42.800 73.800 43.000 ;
        RECT 70.200 42.200 73.800 42.800 ;
        RECT 76.400 42.200 77.200 49.700 ;
        RECT 78.000 49.600 78.800 49.700 ;
        RECT 82.800 50.400 83.400 53.600 ;
        RECT 88.800 50.400 89.400 57.000 ;
        RECT 92.400 56.300 94.800 56.400 ;
        RECT 92.400 55.700 96.300 56.300 ;
        RECT 97.200 56.000 98.000 59.800 ;
        RECT 100.400 56.000 101.200 59.800 ;
        RECT 97.200 55.800 101.200 56.000 ;
        RECT 102.000 55.800 102.800 59.800 ;
        RECT 106.200 56.400 107.000 59.800 ;
        RECT 110.000 57.800 110.800 59.800 ;
        RECT 105.200 55.800 107.000 56.400 ;
        RECT 92.400 55.600 94.800 55.700 ;
        RECT 91.600 53.600 93.200 54.400 ;
        RECT 95.700 54.300 96.300 55.700 ;
        RECT 97.400 55.400 101.000 55.800 ;
        RECT 98.000 54.400 98.800 54.800 ;
        RECT 102.000 54.400 102.600 55.800 ;
        RECT 97.200 54.300 98.800 54.400 ;
        RECT 95.700 53.800 98.800 54.300 ;
        RECT 95.700 53.700 98.000 53.800 ;
        RECT 97.200 53.600 98.000 53.700 ;
        RECT 100.200 53.600 102.800 54.400 ;
        RECT 103.600 53.600 104.400 55.200 ;
        RECT 90.000 52.300 91.600 52.400 ;
        RECT 98.800 52.300 99.600 53.200 ;
        RECT 90.000 51.700 99.600 52.300 ;
        RECT 90.000 51.600 91.600 51.700 ;
        RECT 98.800 51.600 99.600 51.700 ;
        RECT 100.200 52.300 100.800 53.600 ;
        RECT 103.600 52.300 104.400 52.400 ;
        RECT 100.200 51.700 104.400 52.300 ;
        RECT 82.800 49.600 83.600 50.400 ;
        RECT 86.000 49.800 89.400 50.400 ;
        RECT 100.200 50.200 100.800 51.700 ;
        RECT 103.600 51.600 104.400 51.700 ;
        RECT 102.000 50.200 102.800 50.400 ;
        RECT 86.000 49.600 86.800 49.800 ;
        RECT 81.200 47.600 82.000 49.200 ;
        RECT 82.800 47.000 83.400 49.600 ;
        RECT 86.200 49.000 86.800 49.600 ;
        RECT 99.800 49.600 100.800 50.200 ;
        RECT 101.400 49.600 102.800 50.200 ;
        RECT 87.800 49.000 91.400 49.200 ;
        RECT 79.800 46.400 83.400 47.000 ;
        RECT 79.800 46.200 80.400 46.400 ;
        RECT 79.600 42.200 80.400 46.200 ;
        RECT 82.800 46.200 83.400 46.400 ;
        RECT 82.800 42.200 83.600 46.200 ;
        RECT 84.400 43.000 85.200 49.000 ;
        RECT 86.000 43.400 86.800 49.000 ;
        RECT 87.600 48.600 91.400 49.000 ;
        RECT 84.600 42.800 85.200 43.000 ;
        RECT 87.600 43.000 88.400 48.600 ;
        RECT 90.800 48.200 91.400 48.600 ;
        RECT 92.600 48.800 96.200 49.400 ;
        RECT 92.600 48.200 93.200 48.800 ;
        RECT 87.600 42.800 88.200 43.000 ;
        RECT 84.600 42.200 88.200 42.800 ;
        RECT 89.200 42.800 90.000 48.000 ;
        RECT 90.800 43.400 91.600 48.200 ;
        RECT 92.400 42.800 93.200 48.200 ;
        RECT 89.200 42.200 93.200 42.800 ;
        RECT 95.600 48.200 96.200 48.800 ;
        RECT 95.600 42.200 96.400 48.200 ;
        RECT 99.800 42.200 100.600 49.600 ;
        RECT 101.400 48.400 102.000 49.600 ;
        RECT 101.200 47.600 102.000 48.400 ;
        RECT 103.600 48.300 104.400 48.400 ;
        RECT 105.200 48.300 106.000 55.800 ;
        RECT 108.400 55.600 109.200 57.200 ;
        RECT 110.200 56.300 110.800 57.800 ;
        RECT 111.600 56.300 112.400 56.400 ;
        RECT 110.100 55.700 112.400 56.300 ;
        RECT 113.200 55.800 114.000 59.800 ;
        RECT 117.400 56.800 118.200 59.800 ;
        RECT 121.200 57.800 122.000 59.800 ;
        RECT 117.400 55.800 118.800 56.800 ;
        RECT 110.200 54.400 110.800 55.700 ;
        RECT 111.600 55.600 112.400 55.700 ;
        RECT 113.400 55.600 114.000 55.800 ;
        RECT 113.400 55.200 115.200 55.600 ;
        RECT 113.400 55.000 117.600 55.200 ;
        RECT 114.600 54.600 117.600 55.000 ;
        RECT 116.800 54.400 117.600 54.600 ;
        RECT 110.000 53.600 110.800 54.400 ;
        RECT 106.800 48.800 107.600 50.400 ;
        RECT 110.200 50.200 110.800 53.600 ;
        RECT 113.200 52.800 114.000 54.400 ;
        RECT 115.200 53.800 116.000 54.000 ;
        RECT 115.000 53.200 116.000 53.800 ;
        RECT 115.000 52.400 115.600 53.200 ;
        RECT 111.600 50.800 112.400 52.400 ;
        RECT 114.800 51.600 115.600 52.400 ;
        RECT 116.800 51.000 117.400 54.400 ;
        RECT 118.200 52.400 118.800 55.800 ;
        RECT 119.600 55.600 120.400 57.200 ;
        RECT 121.400 54.400 122.000 57.800 ;
        RECT 121.200 53.600 122.000 54.400 ;
        RECT 118.000 52.300 118.800 52.400 ;
        RECT 119.600 52.300 120.400 52.400 ;
        RECT 118.000 51.700 120.400 52.300 ;
        RECT 118.000 51.600 118.800 51.700 ;
        RECT 119.600 51.600 120.400 51.700 ;
        RECT 115.000 50.400 117.400 51.000 ;
        RECT 110.000 49.400 111.800 50.200 ;
        RECT 103.600 47.700 106.000 48.300 ;
        RECT 103.600 47.600 104.400 47.700 ;
        RECT 105.200 42.200 106.000 47.700 ;
        RECT 111.000 42.200 111.800 49.400 ;
        RECT 115.000 46.200 115.600 50.400 ;
        RECT 118.200 50.200 118.800 51.600 ;
        RECT 121.400 50.200 122.000 53.600 ;
        RECT 124.400 53.800 125.200 59.800 ;
        RECT 130.800 56.600 131.600 59.800 ;
        RECT 132.400 57.000 133.200 59.800 ;
        RECT 134.000 57.000 134.800 59.800 ;
        RECT 135.600 57.000 136.400 59.800 ;
        RECT 138.800 57.000 139.600 59.800 ;
        RECT 142.000 57.000 142.800 59.800 ;
        RECT 143.600 57.000 144.400 59.800 ;
        RECT 145.200 57.000 146.000 59.800 ;
        RECT 146.800 57.000 147.600 59.800 ;
        RECT 129.000 55.800 131.600 56.600 ;
        RECT 148.400 56.600 149.200 59.800 ;
        RECT 135.000 55.800 139.600 56.400 ;
        RECT 129.000 55.200 129.800 55.800 ;
        RECT 126.800 54.400 129.800 55.200 ;
        RECT 124.400 53.000 133.200 53.800 ;
        RECT 135.000 53.400 135.800 55.800 ;
        RECT 138.800 55.600 139.600 55.800 ;
        RECT 140.400 55.600 142.000 56.400 ;
        RECT 145.000 55.600 146.000 56.400 ;
        RECT 148.400 55.800 150.800 56.600 ;
        RECT 137.200 53.600 138.000 55.200 ;
        RECT 138.800 54.800 139.600 55.000 ;
        RECT 138.800 54.200 143.200 54.800 ;
        RECT 142.400 54.000 143.200 54.200 ;
        RECT 122.800 50.800 123.600 52.400 ;
        RECT 114.800 42.200 115.600 46.200 ;
        RECT 118.000 42.200 118.800 50.200 ;
        RECT 121.200 49.400 123.000 50.200 ;
        RECT 122.200 44.400 123.000 49.400 ;
        RECT 124.400 47.400 125.200 53.000 ;
        RECT 133.800 52.600 135.800 53.400 ;
        RECT 139.600 52.600 142.800 53.400 ;
        RECT 145.200 52.800 146.000 55.600 ;
        RECT 150.000 55.200 150.800 55.800 ;
        RECT 150.000 54.600 151.800 55.200 ;
        RECT 151.000 53.400 151.800 54.600 ;
        RECT 154.800 54.600 155.600 59.800 ;
        RECT 156.400 56.300 157.200 59.800 ;
        RECT 159.600 58.300 160.400 58.400 ;
        RECT 162.800 58.300 163.600 58.400 ;
        RECT 159.600 57.700 163.600 58.300 ;
        RECT 159.600 57.600 160.400 57.700 ;
        RECT 162.800 57.600 163.600 57.700 ;
        RECT 162.800 56.300 163.600 56.400 ;
        RECT 156.400 55.700 163.600 56.300 ;
        RECT 156.400 55.200 157.400 55.700 ;
        RECT 162.800 55.600 163.600 55.700 ;
        RECT 154.800 54.000 156.000 54.600 ;
        RECT 151.000 52.600 154.800 53.400 ;
        RECT 125.800 52.000 126.600 52.200 ;
        RECT 130.800 52.000 131.600 52.400 ;
        RECT 148.400 52.000 149.200 52.600 ;
        RECT 155.400 52.000 156.000 54.000 ;
        RECT 125.800 51.400 149.200 52.000 ;
        RECT 155.200 51.400 156.000 52.000 ;
        RECT 155.200 49.600 155.800 51.400 ;
        RECT 156.600 50.800 157.400 55.200 ;
        RECT 134.000 49.400 134.800 49.600 ;
        RECT 129.400 49.000 134.800 49.400 ;
        RECT 128.600 48.800 134.800 49.000 ;
        RECT 135.800 49.000 144.400 49.600 ;
        RECT 126.000 48.000 127.600 48.800 ;
        RECT 128.600 48.200 130.000 48.800 ;
        RECT 135.800 48.200 136.400 49.000 ;
        RECT 143.600 48.800 144.400 49.000 ;
        RECT 146.800 49.000 155.800 49.600 ;
        RECT 146.800 48.800 147.600 49.000 ;
        RECT 127.000 47.600 127.600 48.000 ;
        RECT 130.600 47.600 136.400 48.200 ;
        RECT 137.000 47.600 139.600 48.400 ;
        RECT 124.400 46.800 126.400 47.400 ;
        RECT 127.000 46.800 131.200 47.600 ;
        RECT 125.800 46.200 126.400 46.800 ;
        RECT 125.800 45.600 126.800 46.200 ;
        RECT 122.200 43.600 123.600 44.400 ;
        RECT 122.200 42.200 123.000 43.600 ;
        RECT 126.000 42.200 126.800 45.600 ;
        RECT 129.200 42.200 130.000 46.800 ;
        RECT 132.400 42.200 133.200 45.000 ;
        RECT 134.000 42.200 134.800 45.000 ;
        RECT 135.600 42.200 136.400 47.000 ;
        RECT 138.800 42.200 139.600 47.000 ;
        RECT 142.000 42.200 142.800 48.400 ;
        RECT 150.000 47.600 152.600 48.400 ;
        RECT 145.200 46.800 149.400 47.600 ;
        RECT 143.600 42.200 144.400 45.000 ;
        RECT 145.200 42.200 146.000 45.000 ;
        RECT 146.800 42.200 147.600 45.000 ;
        RECT 150.000 42.200 150.800 47.600 ;
        RECT 155.200 47.400 155.800 49.000 ;
        RECT 153.200 46.800 155.800 47.400 ;
        RECT 156.400 50.000 157.400 50.800 ;
        RECT 164.400 53.800 165.200 59.800 ;
        RECT 170.800 56.600 171.600 59.800 ;
        RECT 172.400 57.000 173.200 59.800 ;
        RECT 174.000 57.000 174.800 59.800 ;
        RECT 175.600 57.000 176.400 59.800 ;
        RECT 178.800 57.000 179.600 59.800 ;
        RECT 182.000 57.000 182.800 59.800 ;
        RECT 183.600 57.000 184.400 59.800 ;
        RECT 185.200 57.000 186.000 59.800 ;
        RECT 186.800 57.000 187.600 59.800 ;
        RECT 169.000 55.800 171.600 56.600 ;
        RECT 188.400 56.600 189.200 59.800 ;
        RECT 175.000 55.800 179.600 56.400 ;
        RECT 169.000 55.200 169.800 55.800 ;
        RECT 166.800 54.400 169.800 55.200 ;
        RECT 164.400 53.000 173.200 53.800 ;
        RECT 175.000 53.400 175.800 55.800 ;
        RECT 178.800 55.600 179.600 55.800 ;
        RECT 180.400 55.600 182.000 56.400 ;
        RECT 185.000 55.600 186.000 56.400 ;
        RECT 188.400 55.800 190.800 56.600 ;
        RECT 177.200 53.600 178.000 55.200 ;
        RECT 178.800 54.800 179.600 55.000 ;
        RECT 178.800 54.200 183.200 54.800 ;
        RECT 182.400 54.000 183.200 54.200 ;
        RECT 153.200 42.200 154.000 46.800 ;
        RECT 156.400 42.200 157.200 50.000 ;
        RECT 164.400 47.400 165.200 53.000 ;
        RECT 173.800 52.600 175.800 53.400 ;
        RECT 179.600 52.600 182.800 53.400 ;
        RECT 185.200 52.800 186.000 55.600 ;
        RECT 190.000 55.200 190.800 55.800 ;
        RECT 190.000 54.600 191.800 55.200 ;
        RECT 191.000 53.400 191.800 54.600 ;
        RECT 194.800 54.600 195.600 59.800 ;
        RECT 196.400 56.000 197.200 59.800 ;
        RECT 201.200 57.800 202.000 59.800 ;
        RECT 205.000 58.400 205.800 59.800 ;
        RECT 196.400 55.200 197.400 56.000 ;
        RECT 194.800 54.000 196.000 54.600 ;
        RECT 191.000 52.600 194.800 53.400 ;
        RECT 165.800 52.000 166.600 52.200 ;
        RECT 167.600 52.000 168.400 52.400 ;
        RECT 170.800 52.000 171.600 52.400 ;
        RECT 188.400 52.000 189.200 52.600 ;
        RECT 195.400 52.000 196.000 54.000 ;
        RECT 165.800 51.400 189.200 52.000 ;
        RECT 195.200 51.400 196.000 52.000 ;
        RECT 195.200 49.600 195.800 51.400 ;
        RECT 196.600 50.800 197.400 55.200 ;
        RECT 201.200 54.400 201.800 57.800 ;
        RECT 204.400 57.600 205.800 58.400 ;
        RECT 202.800 55.600 203.600 57.200 ;
        RECT 205.000 56.400 205.800 57.600 ;
        RECT 205.000 55.800 206.800 56.400 ;
        RECT 201.200 53.600 202.000 54.400 ;
        RECT 199.600 50.800 200.400 52.400 ;
        RECT 174.000 49.400 174.800 49.600 ;
        RECT 169.400 49.000 174.800 49.400 ;
        RECT 168.600 48.800 174.800 49.000 ;
        RECT 175.800 49.000 184.400 49.600 ;
        RECT 166.000 48.000 167.600 48.800 ;
        RECT 168.600 48.200 170.000 48.800 ;
        RECT 175.800 48.200 176.400 49.000 ;
        RECT 183.600 48.800 184.400 49.000 ;
        RECT 186.800 49.000 195.800 49.600 ;
        RECT 186.800 48.800 187.600 49.000 ;
        RECT 167.000 47.600 167.600 48.000 ;
        RECT 170.600 47.600 176.400 48.200 ;
        RECT 177.000 47.600 179.600 48.400 ;
        RECT 164.400 46.800 166.400 47.400 ;
        RECT 167.000 46.800 171.200 47.600 ;
        RECT 165.800 46.200 166.400 46.800 ;
        RECT 165.800 45.600 166.800 46.200 ;
        RECT 166.000 42.200 166.800 45.600 ;
        RECT 169.200 42.200 170.000 46.800 ;
        RECT 172.400 42.200 173.200 45.000 ;
        RECT 174.000 42.200 174.800 45.000 ;
        RECT 175.600 42.200 176.400 47.000 ;
        RECT 178.800 42.200 179.600 47.000 ;
        RECT 182.000 42.200 182.800 48.400 ;
        RECT 190.000 47.600 192.600 48.400 ;
        RECT 185.200 46.800 189.400 47.600 ;
        RECT 183.600 42.200 184.400 45.000 ;
        RECT 185.200 42.200 186.000 45.000 ;
        RECT 186.800 42.200 187.600 45.000 ;
        RECT 190.000 42.200 190.800 47.600 ;
        RECT 195.200 47.400 195.800 49.000 ;
        RECT 193.200 46.800 195.800 47.400 ;
        RECT 196.400 50.000 197.400 50.800 ;
        RECT 201.200 50.200 201.800 53.600 ;
        RECT 193.200 42.200 194.000 46.800 ;
        RECT 196.400 42.200 197.200 50.000 ;
        RECT 200.200 49.400 202.000 50.200 ;
        RECT 200.200 42.200 201.000 49.400 ;
        RECT 204.400 47.600 205.200 50.400 ;
        RECT 206.000 42.200 206.800 55.800 ;
        RECT 212.400 55.600 213.200 59.800 ;
        RECT 213.800 56.400 214.600 57.200 ;
        RECT 214.000 55.600 214.800 56.400 ;
        RECT 207.600 54.300 208.400 55.200 ;
        RECT 210.800 54.300 211.600 54.400 ;
        RECT 207.600 53.700 211.600 54.300 ;
        RECT 207.600 53.600 208.400 53.700 ;
        RECT 210.800 52.800 211.600 53.700 ;
        RECT 209.200 52.200 210.000 52.400 ;
        RECT 212.400 52.200 213.000 55.600 ;
        RECT 215.600 55.200 216.400 59.800 ;
        RECT 215.600 54.600 217.800 55.200 ;
        RECT 214.000 52.200 214.800 52.400 ;
        RECT 209.200 51.600 210.800 52.200 ;
        RECT 212.400 51.600 214.800 52.200 ;
        RECT 215.600 51.600 216.400 53.200 ;
        RECT 217.200 51.600 217.800 54.600 ;
        RECT 210.000 51.200 210.800 51.600 ;
        RECT 214.000 50.200 214.600 51.600 ;
        RECT 217.200 50.800 218.400 51.600 ;
        RECT 217.200 50.200 217.800 50.800 ;
        RECT 209.200 49.600 213.200 50.200 ;
        RECT 209.200 42.200 210.000 49.600 ;
        RECT 212.400 42.200 213.200 49.600 ;
        RECT 214.000 42.200 214.800 50.200 ;
        RECT 215.600 49.600 217.800 50.200 ;
        RECT 215.600 42.200 216.400 49.600 ;
        RECT 4.400 32.400 5.200 39.800 ;
        RECT 3.000 31.800 5.200 32.400 ;
        RECT 3.000 31.200 3.600 31.800 ;
        RECT 2.400 30.400 3.600 31.200 ;
        RECT 3.000 27.400 3.600 30.400 ;
        RECT 4.400 28.800 5.200 30.400 ;
        RECT 3.000 26.800 5.200 27.400 ;
        RECT 4.400 22.200 5.200 26.800 ;
        RECT 6.000 24.800 6.800 26.400 ;
        RECT 7.600 22.200 8.400 39.800 ;
        RECT 9.200 35.800 10.000 39.800 ;
        RECT 9.400 35.600 10.000 35.800 ;
        RECT 12.400 35.800 13.200 39.800 ;
        RECT 12.400 35.600 13.000 35.800 ;
        RECT 9.400 35.000 13.000 35.600 ;
        RECT 9.400 32.400 10.000 35.000 ;
        RECT 10.800 32.800 11.600 34.400 ;
        RECT 9.200 31.600 10.000 32.400 ;
        RECT 9.400 28.400 10.000 31.600 ;
        RECT 14.000 32.300 14.800 32.400 ;
        RECT 15.600 32.300 16.400 39.800 ;
        RECT 14.000 31.700 16.400 32.300 ;
        RECT 18.800 32.400 19.600 39.800 ;
        RECT 20.400 32.400 21.200 32.600 ;
        RECT 23.200 32.400 24.800 39.800 ;
        RECT 18.800 31.800 21.200 32.400 ;
        RECT 22.800 31.800 24.800 32.400 ;
        RECT 27.000 32.400 27.800 32.600 ;
        RECT 28.400 32.400 29.200 39.800 ;
        RECT 32.600 38.400 33.400 39.800 ;
        RECT 31.600 37.600 33.400 38.400 ;
        RECT 27.000 31.800 29.200 32.400 ;
        RECT 32.600 32.400 33.400 37.600 ;
        RECT 34.000 33.600 34.800 34.400 ;
        RECT 36.400 33.800 37.200 39.800 ;
        RECT 34.200 32.400 34.800 33.600 ;
        RECT 36.600 33.200 37.200 33.800 ;
        RECT 39.600 39.200 43.600 39.800 ;
        RECT 39.600 33.800 40.400 39.200 ;
        RECT 41.200 33.800 42.000 38.600 ;
        RECT 42.800 34.000 43.600 39.200 ;
        RECT 44.600 39.200 48.200 39.800 ;
        RECT 44.600 39.000 45.200 39.200 ;
        RECT 39.600 33.200 40.200 33.800 ;
        RECT 36.600 32.600 40.200 33.200 ;
        RECT 41.400 33.400 42.000 33.800 ;
        RECT 44.400 33.400 45.200 39.000 ;
        RECT 47.600 39.000 48.200 39.200 ;
        RECT 41.400 33.000 45.200 33.400 ;
        RECT 46.000 33.000 46.800 38.600 ;
        RECT 47.600 33.000 48.400 39.000 ;
        RECT 41.400 32.800 45.000 33.000 ;
        RECT 46.000 32.400 46.600 33.000 ;
        RECT 32.600 31.800 33.600 32.400 ;
        RECT 34.200 31.800 35.600 32.400 ;
        RECT 46.000 32.200 46.800 32.400 ;
        RECT 14.000 30.800 14.800 31.700 ;
        RECT 11.600 29.600 13.200 30.400 ;
        RECT 9.400 28.200 11.000 28.400 ;
        RECT 9.400 27.800 11.200 28.200 ;
        RECT 10.400 22.200 11.200 27.800 ;
        RECT 15.600 22.200 16.400 31.700 ;
        RECT 22.800 30.400 23.400 31.800 ;
        RECT 27.000 31.200 27.600 31.800 ;
        RECT 24.200 30.600 27.600 31.200 ;
        RECT 24.200 30.400 25.000 30.600 ;
        RECT 22.000 29.800 23.400 30.400 ;
        RECT 30.000 30.300 30.800 30.400 ;
        RECT 31.600 30.300 32.400 30.400 ;
        RECT 26.400 29.800 27.200 30.000 ;
        RECT 22.000 29.600 23.800 29.800 ;
        RECT 22.800 29.200 23.800 29.600 ;
        RECT 18.800 28.300 20.400 28.400 ;
        RECT 17.300 27.700 20.400 28.300 ;
        RECT 17.300 26.400 17.900 27.700 ;
        RECT 18.800 27.600 20.400 27.700 ;
        RECT 21.600 27.600 22.400 28.400 ;
        RECT 21.800 27.200 22.400 27.600 ;
        RECT 20.400 26.800 21.200 27.000 ;
        RECT 17.200 24.800 18.000 26.400 ;
        RECT 18.800 26.200 21.200 26.800 ;
        RECT 21.800 26.400 22.600 27.200 ;
        RECT 18.800 22.200 19.600 26.200 ;
        RECT 23.200 25.800 23.800 29.200 ;
        RECT 24.600 29.200 27.200 29.800 ;
        RECT 28.500 29.700 32.400 30.300 ;
        RECT 24.600 28.600 25.200 29.200 ;
        RECT 24.400 27.800 25.200 28.600 ;
        RECT 28.500 28.400 29.100 29.700 ;
        RECT 30.000 29.600 30.800 29.700 ;
        RECT 31.600 28.800 32.400 29.700 ;
        RECT 33.000 28.400 33.600 31.800 ;
        RECT 34.800 31.600 35.600 31.800 ;
        RECT 43.400 31.600 46.800 32.200 ;
        RECT 34.900 30.300 35.500 31.600 ;
        RECT 34.900 29.700 38.700 30.300 ;
        RECT 27.600 28.200 29.200 28.400 ;
        RECT 25.800 27.600 29.200 28.200 ;
        RECT 30.000 28.200 30.800 28.400 ;
        RECT 30.000 27.600 31.600 28.200 ;
        RECT 33.000 27.600 35.600 28.400 ;
        RECT 38.100 28.300 38.700 29.700 ;
        RECT 41.200 29.600 42.800 30.400 ;
        RECT 39.600 28.300 41.200 28.400 ;
        RECT 38.100 27.700 41.200 28.300 ;
        RECT 39.600 27.600 41.200 27.700 ;
        RECT 25.800 27.200 26.400 27.600 ;
        RECT 30.800 27.200 31.600 27.600 ;
        RECT 24.400 26.600 26.400 27.200 ;
        RECT 27.000 26.800 27.800 27.000 ;
        RECT 24.400 26.400 26.000 26.600 ;
        RECT 27.000 26.200 29.200 26.800 ;
        RECT 30.200 26.200 33.800 26.600 ;
        RECT 34.800 26.200 35.400 27.600 ;
        RECT 23.200 24.400 24.800 25.800 ;
        RECT 23.200 23.600 26.000 24.400 ;
        RECT 23.200 22.200 24.800 23.600 ;
        RECT 28.400 22.200 29.200 26.200 ;
        RECT 30.000 26.000 34.000 26.200 ;
        RECT 30.000 22.200 30.800 26.000 ;
        RECT 33.200 22.200 34.000 26.000 ;
        RECT 34.800 22.200 35.600 26.200 ;
        RECT 38.000 25.600 39.800 26.400 ;
        RECT 43.400 25.000 44.000 31.600 ;
        RECT 40.000 24.400 44.000 25.000 ;
        RECT 40.000 24.200 40.600 24.400 ;
        RECT 39.600 23.600 40.600 24.200 ;
        RECT 42.800 24.200 44.000 24.400 ;
        RECT 39.600 22.200 40.400 23.600 ;
        RECT 42.800 22.200 43.600 24.200 ;
        RECT 49.200 22.200 50.000 39.800 ;
        RECT 52.400 26.800 53.200 28.400 ;
        RECT 50.800 24.800 51.600 26.400 ;
        RECT 54.000 26.200 54.800 39.800 ;
        RECT 55.600 31.600 56.400 33.200 ;
        RECT 62.000 32.400 62.800 39.800 ;
        RECT 63.400 32.400 64.200 32.600 ;
        RECT 62.000 31.800 64.200 32.400 ;
        RECT 66.400 32.400 68.000 39.800 ;
        RECT 70.000 32.400 70.800 32.600 ;
        RECT 71.600 32.400 72.400 39.800 ;
        RECT 74.800 36.400 75.600 39.800 ;
        RECT 74.600 35.800 75.600 36.400 ;
        RECT 74.600 35.200 75.200 35.800 ;
        RECT 78.000 35.200 78.800 39.800 ;
        RECT 81.200 37.000 82.000 39.800 ;
        RECT 82.800 37.000 83.600 39.800 ;
        RECT 66.400 31.800 68.400 32.400 ;
        RECT 70.000 31.800 72.400 32.400 ;
        RECT 73.200 34.600 75.200 35.200 ;
        RECT 63.600 31.200 64.200 31.800 ;
        RECT 63.600 30.600 67.000 31.200 ;
        RECT 66.200 30.400 67.000 30.600 ;
        RECT 67.800 30.400 68.400 31.800 ;
        RECT 67.800 30.300 69.200 30.400 ;
        RECT 71.600 30.300 72.400 30.400 ;
        RECT 64.000 29.800 64.800 30.000 ;
        RECT 67.800 29.800 72.400 30.300 ;
        RECT 64.000 29.200 66.600 29.800 ;
        RECT 66.000 28.600 66.600 29.200 ;
        RECT 67.400 29.700 72.400 29.800 ;
        RECT 67.400 29.600 69.200 29.700 ;
        RECT 71.600 29.600 72.400 29.700 ;
        RECT 67.400 29.200 68.400 29.600 ;
        RECT 55.600 28.300 56.400 28.400 ;
        RECT 62.000 28.300 63.600 28.400 ;
        RECT 55.600 28.200 63.600 28.300 ;
        RECT 55.600 27.700 65.400 28.200 ;
        RECT 66.000 27.800 66.800 28.600 ;
        RECT 55.600 27.600 56.400 27.700 ;
        RECT 62.000 27.600 65.400 27.700 ;
        RECT 64.800 27.200 65.400 27.600 ;
        RECT 63.400 26.800 64.200 27.000 ;
        RECT 62.000 26.200 64.200 26.800 ;
        RECT 64.800 26.600 66.800 27.200 ;
        RECT 65.200 26.400 66.800 26.600 ;
        RECT 54.000 25.600 55.800 26.200 ;
        RECT 55.000 24.300 55.800 25.600 ;
        RECT 60.400 24.300 61.200 24.400 ;
        RECT 55.000 23.700 61.200 24.300 ;
        RECT 55.000 22.200 55.800 23.700 ;
        RECT 60.400 23.600 61.200 23.700 ;
        RECT 62.000 22.200 62.800 26.200 ;
        RECT 67.400 25.800 68.000 29.200 ;
        RECT 73.200 29.000 74.000 34.600 ;
        RECT 75.800 34.400 80.000 35.200 ;
        RECT 84.400 35.000 85.200 39.800 ;
        RECT 87.600 35.000 88.400 39.800 ;
        RECT 75.800 34.000 76.400 34.400 ;
        RECT 74.800 33.200 76.400 34.000 ;
        RECT 79.400 33.800 85.200 34.400 ;
        RECT 77.400 33.200 78.800 33.800 ;
        RECT 77.400 33.000 83.600 33.200 ;
        RECT 78.200 32.600 83.600 33.000 ;
        RECT 82.800 32.400 83.600 32.600 ;
        RECT 84.600 33.000 85.200 33.800 ;
        RECT 85.800 33.600 88.400 34.400 ;
        RECT 90.800 33.600 91.600 39.800 ;
        RECT 92.400 37.000 93.200 39.800 ;
        RECT 94.000 37.000 94.800 39.800 ;
        RECT 95.600 37.000 96.400 39.800 ;
        RECT 94.000 34.400 98.200 35.200 ;
        RECT 98.800 34.400 99.600 39.800 ;
        RECT 102.000 35.200 102.800 39.800 ;
        RECT 102.000 34.600 104.600 35.200 ;
        RECT 98.800 33.600 101.400 34.400 ;
        RECT 92.400 33.000 93.200 33.200 ;
        RECT 84.600 32.400 93.200 33.000 ;
        RECT 95.600 33.000 96.400 33.200 ;
        RECT 104.000 33.000 104.600 34.600 ;
        RECT 95.600 32.400 104.600 33.000 ;
        RECT 104.000 30.600 104.600 32.400 ;
        RECT 105.200 32.000 106.000 39.800 ;
        RECT 110.000 32.000 110.800 39.800 ;
        RECT 113.200 35.200 114.000 39.800 ;
        RECT 105.200 31.200 106.200 32.000 ;
        RECT 74.600 30.000 98.000 30.600 ;
        RECT 104.000 30.000 104.800 30.600 ;
        RECT 74.600 29.800 75.400 30.000 ;
        RECT 78.000 29.600 78.800 30.000 ;
        RECT 79.600 29.600 80.400 30.000 ;
        RECT 97.200 29.400 98.000 30.000 ;
        RECT 68.800 27.600 69.600 28.400 ;
        RECT 70.800 27.600 72.400 28.400 ;
        RECT 73.200 28.200 82.000 29.000 ;
        RECT 82.600 28.600 84.600 29.400 ;
        RECT 88.400 28.600 91.600 29.400 ;
        RECT 68.800 27.200 69.400 27.600 ;
        RECT 68.600 26.400 69.400 27.200 ;
        RECT 70.000 26.800 70.800 27.000 ;
        RECT 70.000 26.200 72.400 26.800 ;
        RECT 66.400 22.200 68.000 25.800 ;
        RECT 71.600 22.200 72.400 26.200 ;
        RECT 73.200 22.200 74.000 28.200 ;
        RECT 75.600 26.800 78.600 27.600 ;
        RECT 77.800 26.200 78.600 26.800 ;
        RECT 83.800 26.200 84.600 28.600 ;
        RECT 86.000 26.800 86.800 28.400 ;
        RECT 91.200 27.800 92.000 28.000 ;
        RECT 87.600 27.200 92.000 27.800 ;
        RECT 87.600 27.000 88.400 27.200 ;
        RECT 94.000 26.400 94.800 29.200 ;
        RECT 99.800 28.600 103.600 29.400 ;
        RECT 99.800 27.400 100.600 28.600 ;
        RECT 104.200 28.000 104.800 30.000 ;
        RECT 87.600 26.200 88.400 26.400 ;
        RECT 77.800 25.400 80.400 26.200 ;
        RECT 83.800 25.600 88.400 26.200 ;
        RECT 89.200 25.600 90.800 26.400 ;
        RECT 93.800 25.600 94.800 26.400 ;
        RECT 98.800 26.800 100.600 27.400 ;
        RECT 103.600 27.400 104.800 28.000 ;
        RECT 98.800 26.200 99.600 26.800 ;
        RECT 79.600 22.200 80.400 25.400 ;
        RECT 97.200 25.400 99.600 26.200 ;
        RECT 81.200 22.200 82.000 25.000 ;
        RECT 82.800 22.200 83.600 25.000 ;
        RECT 84.400 22.200 85.200 25.000 ;
        RECT 87.600 22.200 88.400 25.000 ;
        RECT 90.800 22.200 91.600 25.000 ;
        RECT 92.400 22.200 93.200 25.000 ;
        RECT 94.000 22.200 94.800 25.000 ;
        RECT 95.600 22.200 96.400 25.000 ;
        RECT 97.200 22.200 98.000 25.400 ;
        RECT 103.600 22.200 104.400 27.400 ;
        RECT 105.400 26.800 106.200 31.200 ;
        RECT 105.200 26.000 106.200 26.800 ;
        RECT 109.800 31.200 110.800 32.000 ;
        RECT 111.400 34.600 114.000 35.200 ;
        RECT 111.400 33.000 112.000 34.600 ;
        RECT 116.400 34.400 117.200 39.800 ;
        RECT 119.600 37.000 120.400 39.800 ;
        RECT 121.200 37.000 122.000 39.800 ;
        RECT 122.800 37.000 123.600 39.800 ;
        RECT 117.800 34.400 122.000 35.200 ;
        RECT 114.600 33.600 117.200 34.400 ;
        RECT 124.400 33.600 125.200 39.800 ;
        RECT 127.600 35.000 128.400 39.800 ;
        RECT 130.800 35.000 131.600 39.800 ;
        RECT 132.400 37.000 133.200 39.800 ;
        RECT 134.000 37.000 134.800 39.800 ;
        RECT 137.200 35.200 138.000 39.800 ;
        RECT 140.400 36.400 141.200 39.800 ;
        RECT 140.400 35.800 141.400 36.400 ;
        RECT 140.800 35.200 141.400 35.800 ;
        RECT 136.000 34.400 140.200 35.200 ;
        RECT 140.800 34.600 142.800 35.200 ;
        RECT 127.600 33.600 130.200 34.400 ;
        RECT 130.800 33.800 136.600 34.400 ;
        RECT 139.600 34.000 140.200 34.400 ;
        RECT 119.600 33.000 120.400 33.200 ;
        RECT 111.400 32.400 120.400 33.000 ;
        RECT 122.800 33.000 123.600 33.200 ;
        RECT 130.800 33.000 131.400 33.800 ;
        RECT 137.200 33.200 138.600 33.800 ;
        RECT 139.600 33.200 141.200 34.000 ;
        RECT 122.800 32.400 131.400 33.000 ;
        RECT 132.400 33.000 138.600 33.200 ;
        RECT 132.400 32.600 137.800 33.000 ;
        RECT 132.400 32.400 133.200 32.600 ;
        RECT 109.800 26.800 110.600 31.200 ;
        RECT 111.400 30.600 112.000 32.400 ;
        RECT 135.400 31.800 136.400 32.000 ;
        RECT 138.800 31.800 139.600 32.400 ;
        RECT 112.600 31.200 139.600 31.800 ;
        RECT 112.600 31.000 113.400 31.200 ;
        RECT 111.200 30.000 112.000 30.600 ;
        RECT 111.200 28.000 111.800 30.000 ;
        RECT 112.400 28.600 116.200 29.400 ;
        RECT 111.200 27.400 112.400 28.000 ;
        RECT 109.800 26.000 110.800 26.800 ;
        RECT 105.200 22.200 106.000 26.000 ;
        RECT 110.000 22.200 110.800 26.000 ;
        RECT 111.600 22.200 112.400 27.400 ;
        RECT 115.400 27.400 116.200 28.600 ;
        RECT 115.400 26.800 117.200 27.400 ;
        RECT 116.400 26.200 117.200 26.800 ;
        RECT 121.200 26.400 122.000 29.200 ;
        RECT 124.400 28.600 127.600 29.400 ;
        RECT 131.400 28.600 133.400 29.400 ;
        RECT 142.000 29.000 142.800 34.600 ;
        RECT 124.000 27.800 124.800 28.000 ;
        RECT 124.000 27.200 128.400 27.800 ;
        RECT 127.600 27.000 128.400 27.200 ;
        RECT 129.200 26.800 130.000 28.400 ;
        RECT 116.400 25.400 118.800 26.200 ;
        RECT 121.200 25.600 122.200 26.400 ;
        RECT 125.200 25.600 126.800 26.400 ;
        RECT 127.600 26.200 128.400 26.400 ;
        RECT 131.400 26.200 132.200 28.600 ;
        RECT 134.000 28.200 142.800 29.000 ;
        RECT 137.400 26.800 140.400 27.600 ;
        RECT 137.400 26.200 138.200 26.800 ;
        RECT 127.600 25.600 132.200 26.200 ;
        RECT 118.000 22.200 118.800 25.400 ;
        RECT 135.600 25.400 138.200 26.200 ;
        RECT 119.600 22.200 120.400 25.000 ;
        RECT 121.200 22.200 122.000 25.000 ;
        RECT 122.800 22.200 123.600 25.000 ;
        RECT 124.400 22.200 125.200 25.000 ;
        RECT 127.600 22.200 128.400 25.000 ;
        RECT 130.800 22.200 131.600 25.000 ;
        RECT 132.400 22.200 133.200 25.000 ;
        RECT 134.000 22.200 134.800 25.000 ;
        RECT 135.600 22.200 136.400 25.400 ;
        RECT 142.000 22.200 142.800 28.200 ;
        RECT 143.600 26.800 144.400 28.400 ;
        RECT 145.200 26.200 146.000 39.800 ;
        RECT 146.800 31.600 147.600 33.200 ;
        RECT 149.000 32.600 149.800 39.800 ;
        RECT 149.000 31.800 150.800 32.600 ;
        RECT 146.900 30.300 147.500 31.600 ;
        RECT 148.400 30.300 149.200 31.200 ;
        RECT 146.900 29.700 149.200 30.300 ;
        RECT 148.400 29.600 149.200 29.700 ;
        RECT 150.000 28.400 150.600 31.800 ;
        RECT 159.600 30.300 160.400 39.800 ;
        RECT 161.800 32.600 162.600 39.800 ;
        RECT 167.600 36.400 168.400 39.800 ;
        RECT 167.400 35.800 168.400 36.400 ;
        RECT 167.400 35.200 168.000 35.800 ;
        RECT 170.800 35.200 171.600 39.800 ;
        RECT 174.000 37.000 174.800 39.800 ;
        RECT 175.600 37.000 176.400 39.800 ;
        RECT 166.000 34.600 168.000 35.200 ;
        RECT 161.800 31.800 163.600 32.600 ;
        RECT 161.200 30.300 162.000 31.200 ;
        RECT 159.600 29.700 162.000 30.300 ;
        RECT 150.000 28.300 150.800 28.400 ;
        RECT 156.400 28.300 157.200 28.400 ;
        RECT 150.000 27.700 157.200 28.300 ;
        RECT 150.000 27.600 150.800 27.700 ;
        RECT 156.400 27.600 157.200 27.700 ;
        RECT 145.200 25.600 147.000 26.200 ;
        RECT 146.200 24.400 147.000 25.600 ;
        RECT 146.200 23.600 147.600 24.400 ;
        RECT 150.000 24.200 150.600 27.600 ;
        RECT 151.600 24.800 152.400 26.400 ;
        RECT 158.000 24.800 158.800 26.400 ;
        RECT 146.200 22.200 147.000 23.600 ;
        RECT 150.000 22.200 150.800 24.200 ;
        RECT 159.600 22.200 160.400 29.700 ;
        RECT 161.200 29.600 162.000 29.700 ;
        RECT 162.800 28.400 163.400 31.800 ;
        RECT 166.000 29.000 166.800 34.600 ;
        RECT 168.600 34.400 172.800 35.200 ;
        RECT 177.200 35.000 178.000 39.800 ;
        RECT 180.400 35.000 181.200 39.800 ;
        RECT 168.600 34.000 169.200 34.400 ;
        RECT 167.600 33.200 169.200 34.000 ;
        RECT 172.200 33.800 178.000 34.400 ;
        RECT 170.200 33.200 171.600 33.800 ;
        RECT 170.200 33.000 176.400 33.200 ;
        RECT 171.000 32.600 176.400 33.000 ;
        RECT 175.600 32.400 176.400 32.600 ;
        RECT 177.400 33.000 178.000 33.800 ;
        RECT 178.600 33.600 181.200 34.400 ;
        RECT 183.600 33.600 184.400 39.800 ;
        RECT 185.200 37.000 186.000 39.800 ;
        RECT 186.800 37.000 187.600 39.800 ;
        RECT 188.400 37.000 189.200 39.800 ;
        RECT 186.800 34.400 191.000 35.200 ;
        RECT 191.600 34.400 192.400 39.800 ;
        RECT 194.800 35.200 195.600 39.800 ;
        RECT 194.800 34.600 197.400 35.200 ;
        RECT 191.600 33.600 194.200 34.400 ;
        RECT 185.200 33.000 186.000 33.200 ;
        RECT 177.400 32.400 186.000 33.000 ;
        RECT 188.400 33.000 189.200 33.200 ;
        RECT 196.800 33.000 197.400 34.600 ;
        RECT 188.400 32.400 197.400 33.000 ;
        RECT 196.800 30.600 197.400 32.400 ;
        RECT 198.000 32.000 198.800 39.800 ;
        RECT 201.200 32.400 202.000 39.800 ;
        RECT 203.000 32.400 203.800 32.600 ;
        RECT 198.000 31.200 199.000 32.000 ;
        RECT 201.200 31.800 203.800 32.400 ;
        RECT 205.600 31.800 207.200 39.800 ;
        RECT 209.200 32.400 210.000 32.600 ;
        RECT 210.800 32.400 211.600 39.800 ;
        RECT 209.200 31.800 211.600 32.400 ;
        RECT 212.400 32.400 213.200 39.800 ;
        RECT 212.400 31.800 214.600 32.400 ;
        RECT 167.400 30.000 190.800 30.600 ;
        RECT 196.800 30.000 197.600 30.600 ;
        RECT 167.400 29.800 168.200 30.000 ;
        RECT 170.800 29.600 171.600 30.000 ;
        RECT 172.400 29.600 173.200 30.000 ;
        RECT 190.000 29.400 190.800 30.000 ;
        RECT 162.800 27.600 163.600 28.400 ;
        RECT 166.000 28.200 174.800 29.000 ;
        RECT 175.400 28.600 177.400 29.400 ;
        RECT 181.200 28.600 184.400 29.400 ;
        RECT 162.800 24.400 163.400 27.600 ;
        RECT 164.400 24.800 165.200 26.400 ;
        RECT 162.800 22.200 163.600 24.400 ;
        RECT 166.000 22.200 166.800 28.200 ;
        RECT 168.400 26.800 171.400 27.600 ;
        RECT 170.600 26.200 171.400 26.800 ;
        RECT 176.600 26.200 177.400 28.600 ;
        RECT 178.800 26.800 179.600 28.400 ;
        RECT 184.000 27.800 184.800 28.000 ;
        RECT 180.400 27.200 184.800 27.800 ;
        RECT 180.400 27.000 181.200 27.200 ;
        RECT 186.800 26.400 187.600 29.200 ;
        RECT 192.600 28.600 196.400 29.400 ;
        RECT 192.600 27.400 193.400 28.600 ;
        RECT 197.000 28.000 197.600 30.000 ;
        RECT 180.400 26.200 181.200 26.400 ;
        RECT 170.600 25.400 173.200 26.200 ;
        RECT 176.600 25.600 181.200 26.200 ;
        RECT 182.000 25.600 183.600 26.400 ;
        RECT 186.600 25.600 187.600 26.400 ;
        RECT 191.600 26.800 193.400 27.400 ;
        RECT 196.400 27.400 197.600 28.000 ;
        RECT 191.600 26.200 192.400 26.800 ;
        RECT 172.400 22.200 173.200 25.400 ;
        RECT 190.000 25.400 192.400 26.200 ;
        RECT 174.000 22.200 174.800 25.000 ;
        RECT 175.600 22.200 176.400 25.000 ;
        RECT 177.200 22.200 178.000 25.000 ;
        RECT 180.400 22.200 181.200 25.000 ;
        RECT 183.600 22.200 184.400 25.000 ;
        RECT 185.200 22.200 186.000 25.000 ;
        RECT 186.800 22.200 187.600 25.000 ;
        RECT 188.400 22.200 189.200 25.000 ;
        RECT 190.000 22.200 190.800 25.400 ;
        RECT 196.400 22.200 197.200 27.400 ;
        RECT 198.200 26.800 199.000 31.200 ;
        RECT 204.200 30.400 205.000 30.600 ;
        RECT 206.200 30.400 206.800 31.800 ;
        RECT 214.000 31.200 214.600 31.800 ;
        RECT 214.000 30.400 215.200 31.200 ;
        RECT 203.400 29.800 205.000 30.400 ;
        RECT 203.400 29.600 204.200 29.800 ;
        RECT 206.000 29.600 206.800 30.400 ;
        RECT 210.800 30.300 211.600 30.400 ;
        RECT 212.400 30.300 213.200 30.400 ;
        RECT 210.800 29.700 213.200 30.300 ;
        RECT 210.800 29.600 211.600 29.700 ;
        RECT 204.800 28.600 205.600 28.800 ;
        RECT 202.800 28.400 205.600 28.600 ;
        RECT 201.200 28.000 205.600 28.400 ;
        RECT 206.200 28.400 206.800 29.600 ;
        RECT 210.900 28.400 211.500 29.600 ;
        RECT 212.400 28.800 213.200 29.700 ;
        RECT 201.200 27.800 203.400 28.000 ;
        RECT 206.200 27.800 207.200 28.400 ;
        RECT 201.200 27.600 202.800 27.800 ;
        RECT 203.000 26.800 203.800 27.000 ;
        RECT 198.000 26.000 199.000 26.800 ;
        RECT 201.200 26.200 203.800 26.800 ;
        RECT 204.400 26.400 206.000 27.200 ;
        RECT 198.000 22.200 198.800 26.000 ;
        RECT 201.200 22.200 202.000 26.200 ;
        RECT 206.600 25.800 207.200 27.800 ;
        RECT 208.000 27.600 208.800 28.400 ;
        RECT 210.000 27.600 211.600 28.400 ;
        RECT 208.000 27.200 208.600 27.600 ;
        RECT 214.000 27.400 214.600 30.400 ;
        RECT 207.800 26.400 208.600 27.200 ;
        RECT 209.200 26.800 210.000 27.000 ;
        RECT 212.400 26.800 214.600 27.400 ;
        RECT 209.200 26.200 211.600 26.800 ;
        RECT 205.600 24.400 207.200 25.800 ;
        RECT 204.400 23.600 207.200 24.400 ;
        RECT 205.600 22.200 207.200 23.600 ;
        RECT 210.800 22.200 211.600 26.200 ;
        RECT 212.400 22.200 213.200 26.800 ;
        RECT 4.400 15.200 5.200 19.800 ;
        RECT 7.600 16.000 8.400 19.800 ;
        RECT 3.000 14.600 5.200 15.200 ;
        RECT 7.400 15.200 8.400 16.000 ;
        RECT 3.000 11.600 3.600 14.600 ;
        RECT 4.400 12.300 5.200 13.200 ;
        RECT 7.400 12.300 8.200 15.200 ;
        RECT 9.200 14.600 10.000 19.800 ;
        RECT 15.600 16.600 16.400 19.800 ;
        RECT 17.200 17.000 18.000 19.800 ;
        RECT 18.800 17.000 19.600 19.800 ;
        RECT 20.400 17.000 21.200 19.800 ;
        RECT 22.000 17.000 22.800 19.800 ;
        RECT 25.200 17.000 26.000 19.800 ;
        RECT 28.400 17.000 29.200 19.800 ;
        RECT 30.000 17.000 30.800 19.800 ;
        RECT 31.600 17.000 32.400 19.800 ;
        RECT 14.000 15.800 16.400 16.600 ;
        RECT 33.200 16.600 34.000 19.800 ;
        RECT 14.000 15.200 14.800 15.800 ;
        RECT 4.400 11.700 8.200 12.300 ;
        RECT 4.400 11.600 5.200 11.700 ;
        RECT 2.400 10.800 3.600 11.600 ;
        RECT 3.000 10.200 3.600 10.800 ;
        RECT 7.400 10.800 8.200 11.700 ;
        RECT 8.800 14.000 10.000 14.600 ;
        RECT 13.000 14.600 14.800 15.200 ;
        RECT 18.800 15.600 19.800 16.400 ;
        RECT 22.800 15.600 24.400 16.400 ;
        RECT 25.200 15.800 29.800 16.400 ;
        RECT 33.200 15.800 35.800 16.600 ;
        RECT 25.200 15.600 26.000 15.800 ;
        RECT 8.800 12.000 9.400 14.000 ;
        RECT 13.000 13.400 13.800 14.600 ;
        RECT 10.000 12.600 13.800 13.400 ;
        RECT 18.800 12.800 19.600 15.600 ;
        RECT 25.200 14.800 26.000 15.000 ;
        RECT 21.600 14.200 26.000 14.800 ;
        RECT 21.600 14.000 22.400 14.200 ;
        RECT 26.800 13.600 27.600 15.200 ;
        RECT 29.000 13.400 29.800 15.800 ;
        RECT 35.000 15.200 35.800 15.800 ;
        RECT 35.000 14.400 38.000 15.200 ;
        RECT 39.600 13.800 40.400 19.800 ;
        RECT 44.400 15.200 45.200 19.800 ;
        RECT 50.800 16.300 51.600 16.400 ;
        RECT 52.400 16.300 53.200 19.800 ;
        RECT 50.800 15.700 53.200 16.300 ;
        RECT 50.800 15.600 51.600 15.700 ;
        RECT 22.000 12.600 25.200 13.400 ;
        RECT 29.000 12.600 31.000 13.400 ;
        RECT 31.600 13.000 40.400 13.800 ;
        RECT 15.600 12.000 16.400 12.600 ;
        RECT 33.200 12.000 34.000 12.400 ;
        RECT 38.200 12.000 39.000 12.200 ;
        RECT 8.800 11.400 9.600 12.000 ;
        RECT 15.600 11.400 39.000 12.000 ;
        RECT 3.000 9.600 5.200 10.200 ;
        RECT 7.400 10.000 8.400 10.800 ;
        RECT 4.400 2.200 5.200 9.600 ;
        RECT 7.600 2.200 8.400 10.000 ;
        RECT 9.000 9.600 9.600 11.400 ;
        RECT 9.000 9.000 18.000 9.600 ;
        RECT 9.000 7.400 9.600 9.000 ;
        RECT 17.200 8.800 18.000 9.000 ;
        RECT 20.400 9.000 29.000 9.600 ;
        RECT 20.400 8.800 21.200 9.000 ;
        RECT 12.200 7.600 14.800 8.400 ;
        RECT 9.000 6.800 11.600 7.400 ;
        RECT 10.800 2.200 11.600 6.800 ;
        RECT 14.000 2.200 14.800 7.600 ;
        RECT 15.400 6.800 19.600 7.600 ;
        RECT 17.200 2.200 18.000 5.000 ;
        RECT 18.800 2.200 19.600 5.000 ;
        RECT 20.400 2.200 21.200 5.000 ;
        RECT 22.000 2.200 22.800 8.400 ;
        RECT 25.200 7.600 27.800 8.400 ;
        RECT 28.400 8.200 29.000 9.000 ;
        RECT 30.000 9.400 30.800 9.600 ;
        RECT 30.000 9.000 35.400 9.400 ;
        RECT 30.000 8.800 36.200 9.000 ;
        RECT 34.800 8.200 36.200 8.800 ;
        RECT 28.400 7.600 34.200 8.200 ;
        RECT 37.200 8.000 38.800 8.800 ;
        RECT 37.200 7.600 37.800 8.000 ;
        RECT 25.200 2.200 26.000 7.000 ;
        RECT 28.400 2.200 29.200 7.000 ;
        RECT 33.600 6.800 37.800 7.600 ;
        RECT 39.600 7.400 40.400 13.000 ;
        RECT 43.000 14.600 45.200 15.200 ;
        RECT 52.200 15.200 53.200 15.700 ;
        RECT 43.000 11.600 43.600 14.600 ;
        RECT 44.400 12.300 45.200 13.200 ;
        RECT 52.200 12.300 53.000 15.200 ;
        RECT 54.000 14.600 54.800 19.800 ;
        RECT 60.400 16.600 61.200 19.800 ;
        RECT 62.000 17.000 62.800 19.800 ;
        RECT 63.600 17.000 64.400 19.800 ;
        RECT 65.200 17.000 66.000 19.800 ;
        RECT 66.800 17.000 67.600 19.800 ;
        RECT 70.000 17.000 70.800 19.800 ;
        RECT 73.200 17.000 74.000 19.800 ;
        RECT 74.800 17.000 75.600 19.800 ;
        RECT 76.400 17.000 77.200 19.800 ;
        RECT 58.800 15.800 61.200 16.600 ;
        RECT 78.000 16.600 78.800 19.800 ;
        RECT 58.800 15.200 59.600 15.800 ;
        RECT 44.400 11.700 53.000 12.300 ;
        RECT 44.400 11.600 45.200 11.700 ;
        RECT 42.400 10.800 43.600 11.600 ;
        RECT 43.000 10.200 43.600 10.800 ;
        RECT 52.200 10.800 53.000 11.700 ;
        RECT 53.600 14.000 54.800 14.600 ;
        RECT 57.800 14.600 59.600 15.200 ;
        RECT 63.600 15.600 64.600 16.400 ;
        RECT 67.600 15.600 69.200 16.400 ;
        RECT 70.000 15.800 74.600 16.400 ;
        RECT 78.000 15.800 80.600 16.600 ;
        RECT 70.000 15.600 70.800 15.800 ;
        RECT 53.600 12.000 54.200 14.000 ;
        RECT 57.800 13.400 58.600 14.600 ;
        RECT 54.800 12.600 58.600 13.400 ;
        RECT 63.600 12.800 64.400 15.600 ;
        RECT 70.000 14.800 70.800 15.000 ;
        RECT 66.400 14.200 70.800 14.800 ;
        RECT 66.400 14.000 67.200 14.200 ;
        RECT 71.600 13.600 72.400 15.200 ;
        RECT 73.800 13.400 74.600 15.800 ;
        RECT 79.800 15.200 80.600 15.800 ;
        RECT 79.800 14.400 82.800 15.200 ;
        RECT 84.400 13.800 85.200 19.800 ;
        RECT 89.200 15.200 90.000 19.800 ;
        RECT 66.800 12.600 70.000 13.400 ;
        RECT 73.800 12.600 75.800 13.400 ;
        RECT 76.400 13.000 85.200 13.800 ;
        RECT 60.400 12.000 61.200 12.600 ;
        RECT 78.000 12.000 78.800 12.400 ;
        RECT 83.000 12.000 83.800 12.200 ;
        RECT 53.600 11.400 54.400 12.000 ;
        RECT 60.400 11.400 83.800 12.000 ;
        RECT 43.000 9.600 45.200 10.200 ;
        RECT 52.200 10.000 53.200 10.800 ;
        RECT 38.400 6.800 40.400 7.400 ;
        RECT 30.000 2.200 30.800 5.000 ;
        RECT 31.600 2.200 32.400 5.000 ;
        RECT 34.800 2.200 35.600 6.800 ;
        RECT 38.400 6.200 39.000 6.800 ;
        RECT 38.000 5.600 39.000 6.200 ;
        RECT 38.000 2.200 38.800 5.600 ;
        RECT 44.400 2.200 45.200 9.600 ;
        RECT 52.400 2.200 53.200 10.000 ;
        RECT 53.800 9.600 54.400 11.400 ;
        RECT 53.800 9.000 62.800 9.600 ;
        RECT 53.800 7.400 54.400 9.000 ;
        RECT 62.000 8.800 62.800 9.000 ;
        RECT 65.200 9.000 73.800 9.600 ;
        RECT 65.200 8.800 66.000 9.000 ;
        RECT 57.000 7.600 59.600 8.400 ;
        RECT 53.800 6.800 56.400 7.400 ;
        RECT 55.600 2.200 56.400 6.800 ;
        RECT 58.800 2.200 59.600 7.600 ;
        RECT 60.200 6.800 64.400 7.600 ;
        RECT 62.000 2.200 62.800 5.000 ;
        RECT 63.600 2.200 64.400 5.000 ;
        RECT 65.200 2.200 66.000 5.000 ;
        RECT 66.800 2.200 67.600 8.400 ;
        RECT 70.000 7.600 72.600 8.400 ;
        RECT 73.200 8.200 73.800 9.000 ;
        RECT 74.800 9.400 75.600 9.600 ;
        RECT 74.800 9.000 80.200 9.400 ;
        RECT 74.800 8.800 81.000 9.000 ;
        RECT 79.600 8.200 81.000 8.800 ;
        RECT 73.200 7.600 79.000 8.200 ;
        RECT 82.000 8.000 83.600 8.800 ;
        RECT 82.000 7.600 82.600 8.000 ;
        RECT 70.000 2.200 70.800 7.000 ;
        RECT 73.200 2.200 74.000 7.000 ;
        RECT 78.400 6.800 82.600 7.600 ;
        RECT 84.400 7.400 85.200 13.000 ;
        RECT 87.800 14.600 90.000 15.200 ;
        RECT 90.800 15.200 91.600 19.800 ;
        RECT 95.600 15.200 96.400 19.800 ;
        RECT 100.400 15.200 101.200 19.800 ;
        RECT 106.800 16.000 107.600 19.800 ;
        RECT 106.600 15.200 107.600 16.000 ;
        RECT 90.800 14.600 93.000 15.200 ;
        RECT 95.600 14.600 97.800 15.200 ;
        RECT 100.400 14.600 102.600 15.200 ;
        RECT 87.800 11.600 88.400 14.600 ;
        RECT 89.200 11.600 90.000 13.200 ;
        RECT 90.800 11.600 91.600 13.200 ;
        RECT 92.400 11.600 93.000 14.600 ;
        RECT 95.600 11.600 96.400 13.200 ;
        RECT 97.200 11.600 97.800 14.600 ;
        RECT 100.400 11.600 101.200 13.200 ;
        RECT 102.000 11.600 102.600 14.600 ;
        RECT 87.200 10.800 88.400 11.600 ;
        RECT 87.800 10.200 88.400 10.800 ;
        RECT 92.400 10.800 93.600 11.600 ;
        RECT 97.200 10.800 98.400 11.600 ;
        RECT 102.000 10.800 103.200 11.600 ;
        RECT 106.600 10.800 107.400 15.200 ;
        RECT 108.400 14.600 109.200 19.800 ;
        RECT 114.800 16.600 115.600 19.800 ;
        RECT 116.400 17.000 117.200 19.800 ;
        RECT 118.000 17.000 118.800 19.800 ;
        RECT 119.600 17.000 120.400 19.800 ;
        RECT 121.200 17.000 122.000 19.800 ;
        RECT 124.400 17.000 125.200 19.800 ;
        RECT 127.600 17.000 128.400 19.800 ;
        RECT 129.200 17.000 130.000 19.800 ;
        RECT 130.800 17.000 131.600 19.800 ;
        RECT 113.200 15.800 115.600 16.600 ;
        RECT 132.400 16.600 133.200 19.800 ;
        RECT 113.200 15.200 114.000 15.800 ;
        RECT 108.000 14.000 109.200 14.600 ;
        RECT 112.200 14.600 114.000 15.200 ;
        RECT 118.000 15.600 119.000 16.400 ;
        RECT 122.000 15.600 123.600 16.400 ;
        RECT 124.400 15.800 129.000 16.400 ;
        RECT 132.400 15.800 135.000 16.600 ;
        RECT 124.400 15.600 125.200 15.800 ;
        RECT 108.000 12.000 108.600 14.000 ;
        RECT 112.200 13.400 113.000 14.600 ;
        RECT 109.200 12.600 113.000 13.400 ;
        RECT 118.000 12.800 118.800 15.600 ;
        RECT 124.400 14.800 125.200 15.000 ;
        RECT 120.800 14.200 125.200 14.800 ;
        RECT 120.800 14.000 121.600 14.200 ;
        RECT 126.000 13.600 126.800 15.200 ;
        RECT 128.200 13.400 129.000 15.800 ;
        RECT 134.200 15.200 135.000 15.800 ;
        RECT 134.200 14.400 137.200 15.200 ;
        RECT 138.800 13.800 139.600 19.800 ;
        RECT 143.600 16.300 144.400 16.400 ;
        RECT 146.800 16.300 147.600 19.800 ;
        RECT 143.600 15.700 147.600 16.300 ;
        RECT 143.600 15.600 144.400 15.700 ;
        RECT 121.200 12.600 124.400 13.400 ;
        RECT 128.200 12.600 130.200 13.400 ;
        RECT 130.800 13.000 139.600 13.800 ;
        RECT 114.800 12.000 115.600 12.600 ;
        RECT 132.400 12.000 133.200 12.400 ;
        RECT 135.600 12.000 136.400 12.400 ;
        RECT 137.400 12.000 138.200 12.200 ;
        RECT 108.000 11.400 108.800 12.000 ;
        RECT 114.800 11.400 138.200 12.000 ;
        RECT 92.400 10.200 93.000 10.800 ;
        RECT 97.200 10.200 97.800 10.800 ;
        RECT 102.000 10.200 102.600 10.800 ;
        RECT 87.800 9.600 90.000 10.200 ;
        RECT 83.200 6.800 85.200 7.400 ;
        RECT 74.800 2.200 75.600 5.000 ;
        RECT 76.400 2.200 77.200 5.000 ;
        RECT 79.600 2.200 80.400 6.800 ;
        RECT 83.200 6.200 83.800 6.800 ;
        RECT 82.800 5.600 83.800 6.200 ;
        RECT 82.800 2.200 83.600 5.600 ;
        RECT 89.200 2.200 90.000 9.600 ;
        RECT 90.800 9.600 93.000 10.200 ;
        RECT 95.600 9.600 97.800 10.200 ;
        RECT 100.400 9.600 102.600 10.200 ;
        RECT 106.600 10.000 107.600 10.800 ;
        RECT 90.800 2.200 91.600 9.600 ;
        RECT 95.600 2.200 96.400 9.600 ;
        RECT 100.400 2.200 101.200 9.600 ;
        RECT 106.800 2.200 107.600 10.000 ;
        RECT 108.200 9.600 108.800 11.400 ;
        RECT 108.200 9.000 117.200 9.600 ;
        RECT 108.200 7.400 108.800 9.000 ;
        RECT 116.400 8.800 117.200 9.000 ;
        RECT 119.600 9.000 128.200 9.600 ;
        RECT 119.600 8.800 120.400 9.000 ;
        RECT 111.400 7.600 114.000 8.400 ;
        RECT 108.200 6.800 110.800 7.400 ;
        RECT 110.000 2.200 110.800 6.800 ;
        RECT 113.200 2.200 114.000 7.600 ;
        RECT 114.600 6.800 118.800 7.600 ;
        RECT 116.400 2.200 117.200 5.000 ;
        RECT 118.000 2.200 118.800 5.000 ;
        RECT 119.600 2.200 120.400 5.000 ;
        RECT 121.200 2.200 122.000 8.400 ;
        RECT 124.400 7.600 127.000 8.400 ;
        RECT 127.600 8.200 128.200 9.000 ;
        RECT 129.200 9.400 130.000 9.600 ;
        RECT 129.200 9.000 134.600 9.400 ;
        RECT 129.200 8.800 135.400 9.000 ;
        RECT 134.000 8.200 135.400 8.800 ;
        RECT 127.600 7.600 133.400 8.200 ;
        RECT 136.400 8.000 138.000 8.800 ;
        RECT 136.400 7.600 137.000 8.000 ;
        RECT 124.400 2.200 125.200 7.000 ;
        RECT 127.600 2.200 128.400 7.000 ;
        RECT 132.800 6.800 137.000 7.600 ;
        RECT 138.800 7.400 139.600 13.000 ;
        RECT 146.600 15.200 147.600 15.700 ;
        RECT 146.600 10.800 147.400 15.200 ;
        RECT 148.400 14.600 149.200 19.800 ;
        RECT 154.800 16.600 155.600 19.800 ;
        RECT 156.400 17.000 157.200 19.800 ;
        RECT 158.000 17.000 158.800 19.800 ;
        RECT 159.600 17.000 160.400 19.800 ;
        RECT 161.200 17.000 162.000 19.800 ;
        RECT 164.400 17.000 165.200 19.800 ;
        RECT 167.600 17.000 168.400 19.800 ;
        RECT 169.200 17.000 170.000 19.800 ;
        RECT 170.800 17.000 171.600 19.800 ;
        RECT 153.200 15.800 155.600 16.600 ;
        RECT 172.400 16.600 173.200 19.800 ;
        RECT 153.200 15.200 154.000 15.800 ;
        RECT 148.000 14.000 149.200 14.600 ;
        RECT 152.200 14.600 154.000 15.200 ;
        RECT 158.000 15.600 159.000 16.400 ;
        RECT 162.000 15.600 163.600 16.400 ;
        RECT 164.400 15.800 169.000 16.400 ;
        RECT 172.400 15.800 175.000 16.600 ;
        RECT 164.400 15.600 165.200 15.800 ;
        RECT 148.000 12.000 148.600 14.000 ;
        RECT 152.200 13.400 153.000 14.600 ;
        RECT 149.200 12.600 153.000 13.400 ;
        RECT 158.000 12.800 158.800 15.600 ;
        RECT 164.400 14.800 165.200 15.000 ;
        RECT 160.800 14.200 165.200 14.800 ;
        RECT 160.800 14.000 161.600 14.200 ;
        RECT 166.000 13.600 166.800 15.200 ;
        RECT 168.200 13.400 169.000 15.800 ;
        RECT 174.200 15.200 175.000 15.800 ;
        RECT 174.200 14.400 177.200 15.200 ;
        RECT 178.800 13.800 179.600 19.800 ;
        RECT 161.200 12.600 164.400 13.400 ;
        RECT 168.200 12.600 170.200 13.400 ;
        RECT 170.800 13.000 179.600 13.800 ;
        RECT 154.800 12.000 155.600 12.600 ;
        RECT 172.400 12.000 173.200 12.400 ;
        RECT 174.000 12.000 174.800 12.400 ;
        RECT 177.400 12.000 178.200 12.200 ;
        RECT 148.000 11.400 148.800 12.000 ;
        RECT 154.800 11.400 178.200 12.000 ;
        RECT 146.600 10.000 147.600 10.800 ;
        RECT 137.600 6.800 139.600 7.400 ;
        RECT 129.200 2.200 130.000 5.000 ;
        RECT 130.800 2.200 131.600 5.000 ;
        RECT 134.000 2.200 134.800 6.800 ;
        RECT 137.600 6.200 138.200 6.800 ;
        RECT 137.200 5.600 138.200 6.200 ;
        RECT 137.200 2.200 138.000 5.600 ;
        RECT 146.800 2.200 147.600 10.000 ;
        RECT 148.200 9.600 148.800 11.400 ;
        RECT 148.200 9.000 157.200 9.600 ;
        RECT 148.200 7.400 148.800 9.000 ;
        RECT 156.400 8.800 157.200 9.000 ;
        RECT 159.600 9.000 168.200 9.600 ;
        RECT 159.600 8.800 160.400 9.000 ;
        RECT 151.400 7.600 154.000 8.400 ;
        RECT 148.200 6.800 150.800 7.400 ;
        RECT 150.000 2.200 150.800 6.800 ;
        RECT 153.200 2.200 154.000 7.600 ;
        RECT 154.600 6.800 158.800 7.600 ;
        RECT 156.400 2.200 157.200 5.000 ;
        RECT 158.000 2.200 158.800 5.000 ;
        RECT 159.600 2.200 160.400 5.000 ;
        RECT 161.200 2.200 162.000 8.400 ;
        RECT 164.400 7.600 167.000 8.400 ;
        RECT 167.600 8.200 168.200 9.000 ;
        RECT 169.200 9.400 170.000 9.600 ;
        RECT 169.200 9.000 174.600 9.400 ;
        RECT 169.200 8.800 175.400 9.000 ;
        RECT 174.000 8.200 175.400 8.800 ;
        RECT 167.600 7.600 173.400 8.200 ;
        RECT 176.400 8.000 178.000 8.800 ;
        RECT 176.400 7.600 177.000 8.000 ;
        RECT 164.400 2.200 165.200 7.000 ;
        RECT 167.600 2.200 168.400 7.000 ;
        RECT 172.800 6.800 177.000 7.600 ;
        RECT 178.800 7.400 179.600 13.000 ;
        RECT 177.600 6.800 179.600 7.400 ;
        RECT 180.400 13.800 181.200 19.800 ;
        RECT 186.800 16.600 187.600 19.800 ;
        RECT 188.400 17.000 189.200 19.800 ;
        RECT 190.000 17.000 190.800 19.800 ;
        RECT 191.600 17.000 192.400 19.800 ;
        RECT 194.800 17.000 195.600 19.800 ;
        RECT 198.000 17.000 198.800 19.800 ;
        RECT 199.600 17.000 200.400 19.800 ;
        RECT 201.200 17.000 202.000 19.800 ;
        RECT 202.800 17.000 203.600 19.800 ;
        RECT 185.000 15.800 187.600 16.600 ;
        RECT 204.400 16.600 205.200 19.800 ;
        RECT 191.000 15.800 195.600 16.400 ;
        RECT 185.000 15.200 185.800 15.800 ;
        RECT 182.800 14.400 185.800 15.200 ;
        RECT 180.400 13.000 189.200 13.800 ;
        RECT 191.000 13.400 191.800 15.800 ;
        RECT 194.800 15.600 195.600 15.800 ;
        RECT 196.400 15.600 198.000 16.400 ;
        RECT 201.000 15.600 202.000 16.400 ;
        RECT 204.400 15.800 206.800 16.600 ;
        RECT 193.200 13.600 194.000 15.200 ;
        RECT 194.800 14.800 195.600 15.000 ;
        RECT 194.800 14.200 199.200 14.800 ;
        RECT 198.400 14.000 199.200 14.200 ;
        RECT 180.400 7.400 181.200 13.000 ;
        RECT 189.800 12.600 191.800 13.400 ;
        RECT 195.600 12.600 198.800 13.400 ;
        RECT 201.200 12.800 202.000 15.600 ;
        RECT 206.000 15.200 206.800 15.800 ;
        RECT 206.000 14.600 207.800 15.200 ;
        RECT 207.000 13.400 207.800 14.600 ;
        RECT 210.800 14.600 211.600 19.800 ;
        RECT 212.400 16.000 213.200 19.800 ;
        RECT 212.400 15.200 213.400 16.000 ;
        RECT 210.800 14.000 212.000 14.600 ;
        RECT 207.000 12.600 210.800 13.400 ;
        RECT 181.800 12.000 182.600 12.200 ;
        RECT 183.600 12.000 184.400 12.400 ;
        RECT 186.800 12.000 187.600 12.400 ;
        RECT 204.400 12.000 205.200 12.600 ;
        RECT 211.400 12.000 212.000 14.000 ;
        RECT 181.800 11.400 205.200 12.000 ;
        RECT 211.200 11.400 212.000 12.000 ;
        RECT 211.200 9.600 211.800 11.400 ;
        RECT 212.600 10.800 213.400 15.200 ;
        RECT 190.000 9.400 190.800 9.600 ;
        RECT 185.400 9.000 190.800 9.400 ;
        RECT 184.600 8.800 190.800 9.000 ;
        RECT 191.800 9.000 200.400 9.600 ;
        RECT 182.000 8.000 183.600 8.800 ;
        RECT 184.600 8.200 186.000 8.800 ;
        RECT 191.800 8.200 192.400 9.000 ;
        RECT 199.600 8.800 200.400 9.000 ;
        RECT 202.800 9.000 211.800 9.600 ;
        RECT 202.800 8.800 203.600 9.000 ;
        RECT 183.000 7.600 183.600 8.000 ;
        RECT 186.600 7.600 192.400 8.200 ;
        RECT 193.000 7.600 195.600 8.400 ;
        RECT 180.400 6.800 182.400 7.400 ;
        RECT 183.000 6.800 187.200 7.600 ;
        RECT 169.200 2.200 170.000 5.000 ;
        RECT 170.800 2.200 171.600 5.000 ;
        RECT 174.000 2.200 174.800 6.800 ;
        RECT 177.600 6.200 178.200 6.800 ;
        RECT 177.200 5.600 178.200 6.200 ;
        RECT 181.800 6.200 182.400 6.800 ;
        RECT 181.800 5.600 182.800 6.200 ;
        RECT 177.200 2.200 178.000 5.600 ;
        RECT 182.000 2.200 182.800 5.600 ;
        RECT 185.200 2.200 186.000 6.800 ;
        RECT 188.400 2.200 189.200 5.000 ;
        RECT 190.000 2.200 190.800 5.000 ;
        RECT 191.600 2.200 192.400 7.000 ;
        RECT 194.800 2.200 195.600 7.000 ;
        RECT 198.000 2.200 198.800 8.400 ;
        RECT 206.000 7.600 208.600 8.400 ;
        RECT 201.200 6.800 205.400 7.600 ;
        RECT 199.600 2.200 200.400 5.000 ;
        RECT 201.200 2.200 202.000 5.000 ;
        RECT 202.800 2.200 203.600 5.000 ;
        RECT 206.000 2.200 206.800 7.600 ;
        RECT 211.200 7.400 211.800 9.000 ;
        RECT 209.200 6.800 211.800 7.400 ;
        RECT 212.400 10.000 213.400 10.800 ;
        RECT 209.200 2.200 210.000 6.800 ;
        RECT 212.400 2.200 213.200 10.000 ;
      LAYER via1 ;
        RECT 7.800 191.800 8.600 192.600 ;
        RECT 4.400 189.600 5.200 190.400 ;
        RECT 9.000 189.800 9.800 190.600 ;
        RECT 7.800 186.200 8.600 187.000 ;
        RECT 10.800 183.600 11.600 184.400 ;
        RECT 17.200 185.600 18.000 186.400 ;
        RECT 26.800 189.600 27.600 190.400 ;
        RECT 28.400 187.600 29.200 188.400 ;
        RECT 50.800 193.600 51.600 194.400 ;
        RECT 54.000 193.600 54.800 194.400 ;
        RECT 47.600 191.600 48.400 192.400 ;
        RECT 46.000 187.600 46.800 188.400 ;
        RECT 28.400 183.600 29.200 184.400 ;
        RECT 44.400 185.600 45.200 186.400 ;
        RECT 52.400 187.600 53.200 188.400 ;
        RECT 57.200 187.600 58.000 188.400 ;
        RECT 58.800 187.600 59.600 188.400 ;
        RECT 55.600 185.600 56.400 186.400 ;
        RECT 79.600 194.400 80.400 195.200 ;
        RECT 82.800 195.000 83.600 195.800 ;
        RECT 78.000 192.400 78.800 193.200 ;
        RECT 68.200 189.600 69.000 190.400 ;
        RECT 87.600 187.600 88.400 188.400 ;
        RECT 84.400 185.600 85.200 186.400 ;
        RECT 102.000 189.600 102.800 190.400 ;
        RECT 78.000 184.200 78.800 185.000 ;
        RECT 79.600 184.200 80.400 185.000 ;
        RECT 81.200 184.200 82.000 185.000 ;
        RECT 82.800 184.200 83.600 185.000 ;
        RECT 86.000 184.200 86.800 185.000 ;
        RECT 89.200 184.200 90.000 185.000 ;
        RECT 90.800 184.200 91.600 185.000 ;
        RECT 92.400 184.200 93.200 185.000 ;
        RECT 124.400 195.000 125.200 195.800 ;
        RECT 121.200 193.600 122.000 194.400 ;
        RECT 126.000 192.400 126.800 193.200 ;
        RECT 148.400 191.800 149.200 192.600 ;
        RECT 114.800 188.200 115.600 189.000 ;
        RECT 124.400 188.600 125.200 189.400 ;
        RECT 119.600 187.600 120.400 188.400 ;
        RECT 139.000 189.600 139.800 190.400 ;
        RECT 114.800 184.200 115.600 185.000 ;
        RECT 116.400 184.200 117.200 185.000 ;
        RECT 118.000 184.200 118.800 185.000 ;
        RECT 121.200 184.200 122.000 185.000 ;
        RECT 124.400 184.200 125.200 185.000 ;
        RECT 126.000 184.200 126.800 185.000 ;
        RECT 127.600 184.200 128.400 185.000 ;
        RECT 129.200 184.200 130.000 185.000 ;
        RECT 145.200 189.600 146.000 190.400 ;
        RECT 148.400 186.200 149.200 187.000 ;
        RECT 162.800 189.600 163.600 190.400 ;
        RECT 156.400 187.600 157.200 188.400 ;
        RECT 153.200 186.400 154.000 187.200 ;
        RECT 167.600 185.600 168.400 186.400 ;
        RECT 170.800 185.600 171.600 186.400 ;
        RECT 172.400 183.600 173.200 184.400 ;
        RECT 199.600 195.000 200.400 195.800 ;
        RECT 196.400 193.600 197.200 194.400 ;
        RECT 201.200 192.400 202.000 193.200 ;
        RECT 190.000 188.200 190.800 189.000 ;
        RECT 199.600 188.600 200.400 189.400 ;
        RECT 180.400 183.600 181.200 184.400 ;
        RECT 194.800 187.600 195.600 188.400 ;
        RECT 190.000 184.200 190.800 185.000 ;
        RECT 191.600 184.200 192.400 185.000 ;
        RECT 193.200 184.200 194.000 185.000 ;
        RECT 196.400 184.200 197.200 185.000 ;
        RECT 199.600 184.200 200.400 185.000 ;
        RECT 201.200 184.200 202.000 185.000 ;
        RECT 202.800 184.200 203.600 185.000 ;
        RECT 204.400 184.200 205.200 185.000 ;
        RECT 214.000 183.600 214.800 184.400 ;
        RECT 2.800 177.600 3.600 178.400 ;
        RECT 18.800 175.600 19.600 176.400 ;
        RECT 20.400 174.200 21.200 175.000 ;
        RECT 14.000 166.800 14.800 167.600 ;
        RECT 17.200 166.200 18.000 167.000 ;
        RECT 12.400 164.200 13.200 165.000 ;
        RECT 14.000 164.200 14.800 165.000 ;
        RECT 15.600 164.200 16.400 165.000 ;
        RECT 20.400 166.200 21.200 167.000 ;
        RECT 23.600 166.200 24.400 167.000 ;
        RECT 44.400 171.600 45.200 172.400 ;
        RECT 47.600 171.600 48.400 172.400 ;
        RECT 25.200 164.200 26.000 165.000 ;
        RECT 26.800 164.200 27.600 165.000 ;
        RECT 41.200 163.600 42.000 164.400 ;
        RECT 68.400 175.600 69.200 176.400 ;
        RECT 81.200 174.800 82.000 175.600 ;
        RECT 90.800 177.600 91.600 178.400 ;
        RECT 87.600 173.600 88.400 174.400 ;
        RECT 111.600 173.000 112.400 173.800 ;
        RECT 82.800 163.600 83.600 164.400 ;
        RECT 121.200 172.600 122.000 173.400 ;
        RECT 135.600 175.600 136.400 176.400 ;
        RECT 110.000 171.600 110.800 172.400 ;
        RECT 146.800 174.800 147.600 175.600 ;
        RECT 161.200 177.600 162.000 178.400 ;
        RECT 164.400 177.600 165.200 178.400 ;
        RECT 113.200 168.800 114.000 169.600 ;
        RECT 118.000 167.600 118.800 168.400 ;
        RECT 114.800 166.200 115.600 167.000 ;
        RECT 111.600 164.200 112.400 165.000 ;
        RECT 113.200 164.200 114.000 165.000 ;
        RECT 118.000 166.200 118.800 167.000 ;
        RECT 121.200 166.200 122.000 167.000 ;
        RECT 122.800 164.200 123.600 165.000 ;
        RECT 124.400 164.200 125.200 165.000 ;
        RECT 126.000 164.200 126.800 165.000 ;
        RECT 162.800 169.600 163.600 170.400 ;
        RECT 174.000 174.800 174.800 175.600 ;
        RECT 182.000 169.600 182.800 170.400 ;
        RECT 201.200 173.600 202.000 174.400 ;
        RECT 207.600 173.600 208.400 174.400 ;
        RECT 4.400 149.600 5.200 150.400 ;
        RECT 9.200 149.600 10.000 150.400 ;
        RECT 20.400 153.600 21.200 154.400 ;
        RECT 10.800 145.600 11.600 146.400 ;
        RECT 14.000 145.600 14.800 146.400 ;
        RECT 57.200 155.000 58.000 155.800 ;
        RECT 54.000 153.600 54.800 154.400 ;
        RECT 71.600 157.600 72.400 158.400 ;
        RECT 58.800 152.400 59.600 153.200 ;
        RECT 46.000 151.200 46.800 152.000 ;
        RECT 36.400 147.600 37.200 148.400 ;
        RECT 38.000 147.600 38.800 148.400 ;
        RECT 47.600 148.200 48.400 149.000 ;
        RECT 57.200 148.600 58.000 149.400 ;
        RECT 52.400 147.600 53.200 148.400 ;
        RECT 47.600 144.200 48.400 145.000 ;
        RECT 49.200 144.200 50.000 145.000 ;
        RECT 50.800 144.200 51.600 145.000 ;
        RECT 54.000 144.200 54.800 145.000 ;
        RECT 57.200 144.200 58.000 145.000 ;
        RECT 58.800 144.200 59.600 145.000 ;
        RECT 60.400 144.200 61.200 145.000 ;
        RECT 62.000 144.200 62.800 145.000 ;
        RECT 97.200 155.000 98.000 155.800 ;
        RECT 94.000 153.600 94.800 154.400 ;
        RECT 111.600 157.600 112.400 158.400 ;
        RECT 98.800 152.400 99.600 153.200 ;
        RECT 86.000 151.200 86.800 152.000 ;
        RECT 87.600 148.200 88.400 149.000 ;
        RECT 97.200 148.600 98.000 149.400 ;
        RECT 92.400 147.600 93.200 148.400 ;
        RECT 87.600 144.200 88.400 145.000 ;
        RECT 89.200 144.200 90.000 145.000 ;
        RECT 90.800 144.200 91.600 145.000 ;
        RECT 94.000 144.200 94.800 145.000 ;
        RECT 97.200 144.200 98.000 145.000 ;
        RECT 98.800 144.200 99.600 145.000 ;
        RECT 100.400 144.200 101.200 145.000 ;
        RECT 102.000 144.200 102.800 145.000 ;
        RECT 146.800 155.000 147.600 155.800 ;
        RECT 143.600 153.600 144.400 154.400 ;
        RECT 161.200 157.600 162.000 158.400 ;
        RECT 148.400 152.400 149.200 153.200 ;
        RECT 153.200 149.600 154.000 150.400 ;
        RECT 137.200 148.200 138.000 149.000 ;
        RECT 146.800 148.600 147.600 149.400 ;
        RECT 142.000 147.600 142.800 148.400 ;
        RECT 137.200 144.200 138.000 145.000 ;
        RECT 138.800 144.200 139.600 145.000 ;
        RECT 140.400 144.200 141.200 145.000 ;
        RECT 143.600 144.200 144.400 145.000 ;
        RECT 146.800 144.200 147.600 145.000 ;
        RECT 148.400 144.200 149.200 145.000 ;
        RECT 150.000 144.200 150.800 145.000 ;
        RECT 151.600 144.200 152.400 145.000 ;
        RECT 191.600 155.000 192.400 155.800 ;
        RECT 188.400 153.600 189.200 154.400 ;
        RECT 193.200 152.400 194.000 153.200 ;
        RECT 172.400 147.600 173.200 148.400 ;
        RECT 182.000 148.200 182.800 149.000 ;
        RECT 191.600 148.600 192.400 149.400 ;
        RECT 170.800 143.600 171.600 144.400 ;
        RECT 186.800 147.600 187.600 148.400 ;
        RECT 182.000 144.200 182.800 145.000 ;
        RECT 183.600 144.200 184.400 145.000 ;
        RECT 185.200 144.200 186.000 145.000 ;
        RECT 188.400 144.200 189.200 145.000 ;
        RECT 191.600 144.200 192.400 145.000 ;
        RECT 193.200 144.200 194.000 145.000 ;
        RECT 194.800 144.200 195.600 145.000 ;
        RECT 196.400 144.200 197.200 145.000 ;
        RECT 214.000 149.600 214.800 150.400 ;
        RECT 206.000 143.600 206.800 144.400 ;
        RECT 2.800 137.600 3.600 138.400 ;
        RECT 18.800 135.600 19.600 136.400 ;
        RECT 20.400 134.200 21.200 135.000 ;
        RECT 31.600 131.600 32.400 132.400 ;
        RECT 14.000 126.800 14.800 127.600 ;
        RECT 17.200 126.200 18.000 127.000 ;
        RECT 12.400 124.200 13.200 125.000 ;
        RECT 14.000 124.200 14.800 125.000 ;
        RECT 15.600 124.200 16.400 125.000 ;
        RECT 20.400 126.200 21.200 127.000 ;
        RECT 23.600 126.200 24.400 127.000 ;
        RECT 52.400 134.800 53.200 135.600 ;
        RECT 58.800 133.600 59.600 134.400 ;
        RECT 44.400 129.800 45.200 130.600 ;
        RECT 82.800 135.600 83.600 136.400 ;
        RECT 84.400 134.200 85.200 135.000 ;
        RECT 25.200 124.200 26.000 125.000 ;
        RECT 26.800 124.200 27.600 125.000 ;
        RECT 54.000 127.600 54.800 128.400 ;
        RECT 92.400 130.000 93.200 130.800 ;
        RECT 78.000 126.800 78.800 127.600 ;
        RECT 81.200 126.200 82.000 127.000 ;
        RECT 76.400 124.200 77.200 125.000 ;
        RECT 78.000 124.200 78.800 125.000 ;
        RECT 79.600 124.200 80.400 125.000 ;
        RECT 84.400 126.200 85.200 127.000 ;
        RECT 87.600 126.200 88.400 127.000 ;
        RECT 113.200 137.600 114.000 138.400 ;
        RECT 106.800 134.800 107.600 135.600 ;
        RECT 110.000 133.600 110.800 134.400 ;
        RECT 116.400 131.600 117.200 132.400 ;
        RECT 89.200 124.200 90.000 125.000 ;
        RECT 90.800 124.200 91.600 125.000 ;
        RECT 118.000 129.600 118.800 130.400 ;
        RECT 129.200 134.800 130.000 135.600 ;
        RECT 132.400 133.600 133.200 134.400 ;
        RECT 142.000 133.000 142.800 133.800 ;
        RECT 151.600 132.600 152.400 133.400 ;
        RECT 137.200 131.600 138.000 132.400 ;
        RECT 166.200 133.600 167.000 134.400 ;
        RECT 180.400 134.800 181.200 135.600 ;
        RECT 183.600 133.600 184.400 134.400 ;
        RECT 199.600 134.800 200.400 135.600 ;
        RECT 143.600 128.800 144.400 129.600 ;
        RECT 148.400 127.600 149.200 128.400 ;
        RECT 145.200 126.200 146.000 127.000 ;
        RECT 142.000 124.200 142.800 125.000 ;
        RECT 143.600 124.200 144.400 125.000 ;
        RECT 148.400 126.200 149.200 127.000 ;
        RECT 151.600 126.200 152.400 127.000 ;
        RECT 153.200 124.200 154.000 125.000 ;
        RECT 154.800 124.200 155.600 125.000 ;
        RECT 156.400 124.200 157.200 125.000 ;
        RECT 193.200 131.600 194.000 132.400 ;
        RECT 206.000 133.600 206.800 134.400 ;
        RECT 207.600 129.600 208.400 130.400 ;
        RECT 12.400 111.800 13.200 112.600 ;
        RECT 23.600 111.600 24.400 112.400 ;
        RECT 4.400 109.600 5.200 110.400 ;
        RECT 9.200 109.600 10.000 110.400 ;
        RECT 12.400 106.200 13.200 107.000 ;
        RECT 20.400 107.600 21.200 108.400 ;
        RECT 17.200 106.400 18.000 107.200 ;
        RECT 15.600 103.600 16.400 104.400 ;
        RECT 22.000 105.600 22.800 106.400 ;
        RECT 31.600 113.600 32.400 114.400 ;
        RECT 28.400 111.600 29.200 112.400 ;
        RECT 26.800 109.600 27.600 110.400 ;
        RECT 25.200 105.600 26.000 106.400 ;
        RECT 60.400 117.600 61.200 118.400 ;
        RECT 33.200 103.600 34.000 104.400 ;
        RECT 71.600 114.400 72.400 115.200 ;
        RECT 74.800 115.000 75.600 115.800 ;
        RECT 70.000 112.400 70.800 113.200 ;
        RECT 44.400 103.600 45.200 104.400 ;
        RECT 68.400 109.600 69.200 110.400 ;
        RECT 79.600 107.600 80.400 108.400 ;
        RECT 76.400 105.600 77.200 106.400 ;
        RECT 70.000 104.200 70.800 105.000 ;
        RECT 71.600 104.200 72.400 105.000 ;
        RECT 73.200 104.200 74.000 105.000 ;
        RECT 74.800 104.200 75.600 105.000 ;
        RECT 78.000 104.200 78.800 105.000 ;
        RECT 81.200 104.200 82.000 105.000 ;
        RECT 82.800 104.200 83.600 105.000 ;
        RECT 84.400 104.200 85.200 105.000 ;
        RECT 106.800 114.400 107.600 115.200 ;
        RECT 110.000 115.000 110.800 115.800 ;
        RECT 105.200 112.400 106.000 113.200 ;
        RECT 114.800 107.600 115.600 108.400 ;
        RECT 111.600 105.600 112.400 106.400 ;
        RECT 105.200 104.200 106.000 105.000 ;
        RECT 106.800 104.200 107.600 105.000 ;
        RECT 108.400 104.200 109.200 105.000 ;
        RECT 110.000 104.200 110.800 105.000 ;
        RECT 113.200 104.200 114.000 105.000 ;
        RECT 116.400 104.200 117.200 105.000 ;
        RECT 118.000 104.200 118.800 105.000 ;
        RECT 119.600 104.200 120.400 105.000 ;
        RECT 153.200 115.000 154.000 115.800 ;
        RECT 150.000 113.600 150.800 114.400 ;
        RECT 167.600 117.600 168.400 118.400 ;
        RECT 154.800 112.400 155.600 113.200 ;
        RECT 159.600 109.600 160.400 110.400 ;
        RECT 143.600 108.200 144.400 109.000 ;
        RECT 153.200 108.600 154.000 109.400 ;
        RECT 148.400 107.600 149.200 108.400 ;
        RECT 143.600 104.200 144.400 105.000 ;
        RECT 145.200 104.200 146.000 105.000 ;
        RECT 146.800 104.200 147.600 105.000 ;
        RECT 150.000 104.200 150.800 105.000 ;
        RECT 153.200 104.200 154.000 105.000 ;
        RECT 154.800 104.200 155.600 105.000 ;
        RECT 156.400 104.200 157.200 105.000 ;
        RECT 158.000 104.200 158.800 105.000 ;
        RECT 193.200 115.000 194.000 115.800 ;
        RECT 190.000 113.600 190.800 114.400 ;
        RECT 194.800 112.400 195.600 113.200 ;
        RECT 183.600 108.200 184.400 109.000 ;
        RECT 193.200 108.600 194.000 109.400 ;
        RECT 188.400 107.600 189.200 108.400 ;
        RECT 183.600 104.200 184.400 105.000 ;
        RECT 185.200 104.200 186.000 105.000 ;
        RECT 186.800 104.200 187.600 105.000 ;
        RECT 190.000 104.200 190.800 105.000 ;
        RECT 193.200 104.200 194.000 105.000 ;
        RECT 194.800 104.200 195.600 105.000 ;
        RECT 196.400 104.200 197.200 105.000 ;
        RECT 198.000 104.200 198.800 105.000 ;
        RECT 207.600 103.600 208.400 104.400 ;
        RECT 2.800 97.600 3.600 98.400 ;
        RECT 18.800 95.600 19.600 96.400 ;
        RECT 20.400 94.200 21.200 95.000 ;
        RECT 38.000 97.600 38.800 98.400 ;
        RECT 2.800 83.600 3.600 84.400 ;
        RECT 14.000 86.800 14.800 87.600 ;
        RECT 17.200 86.200 18.000 87.000 ;
        RECT 12.400 84.200 13.200 85.000 ;
        RECT 14.000 84.200 14.800 85.000 ;
        RECT 15.600 84.200 16.400 85.000 ;
        RECT 20.400 86.200 21.200 87.000 ;
        RECT 23.600 86.200 24.400 87.000 ;
        RECT 54.000 95.600 54.800 96.400 ;
        RECT 55.600 94.200 56.400 95.000 ;
        RECT 25.200 84.200 26.000 85.000 ;
        RECT 26.800 84.200 27.600 85.000 ;
        RECT 38.000 83.600 38.800 84.400 ;
        RECT 49.200 86.800 50.000 87.600 ;
        RECT 52.400 86.200 53.200 87.000 ;
        RECT 47.600 84.200 48.400 85.000 ;
        RECT 49.200 84.200 50.000 85.000 ;
        RECT 50.800 84.200 51.600 85.000 ;
        RECT 55.600 86.200 56.400 87.000 ;
        RECT 58.800 86.200 59.600 87.000 ;
        RECT 89.200 97.600 90.000 98.400 ;
        RECT 86.000 94.800 86.800 95.600 ;
        RECT 81.200 91.600 82.000 92.400 ;
        RECT 60.400 84.200 61.200 85.000 ;
        RECT 62.000 84.200 62.800 85.000 ;
        RECT 78.000 83.600 78.800 84.400 ;
        RECT 126.000 95.600 126.800 96.400 ;
        RECT 127.600 94.200 128.400 95.000 ;
        RECT 138.800 91.600 139.600 92.400 ;
        RECT 110.000 89.600 110.800 90.400 ;
        RECT 121.200 86.800 122.000 87.600 ;
        RECT 124.400 86.200 125.200 87.000 ;
        RECT 119.600 84.200 120.400 85.000 ;
        RECT 121.200 84.200 122.000 85.000 ;
        RECT 122.800 84.200 123.600 85.000 ;
        RECT 127.600 86.200 128.400 87.000 ;
        RECT 130.800 86.200 131.600 87.000 ;
        RECT 156.400 93.000 157.200 93.800 ;
        RECT 166.000 92.600 166.800 93.400 ;
        RECT 151.600 91.600 152.400 92.400 ;
        RECT 190.000 94.800 190.800 95.600 ;
        RECT 158.000 88.800 158.800 89.600 ;
        RECT 162.800 87.600 163.600 88.400 ;
        RECT 132.400 84.200 133.200 85.000 ;
        RECT 134.000 84.200 134.800 85.000 ;
        RECT 159.600 86.200 160.400 87.000 ;
        RECT 156.400 84.200 157.200 85.000 ;
        RECT 158.000 84.200 158.800 85.000 ;
        RECT 162.800 86.200 163.600 87.000 ;
        RECT 166.000 86.200 166.800 87.000 ;
        RECT 167.600 84.200 168.400 85.000 ;
        RECT 169.200 84.200 170.000 85.000 ;
        RECT 170.800 84.200 171.600 85.000 ;
        RECT 194.800 89.600 195.600 90.400 ;
        RECT 199.600 89.600 200.400 90.400 ;
        RECT 214.000 93.600 214.800 94.400 ;
        RECT 201.200 83.600 202.000 84.400 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 9.200 69.600 10.000 70.400 ;
        RECT 25.200 69.600 26.000 70.400 ;
        RECT 36.200 71.800 37.000 72.600 ;
        RECT 63.600 74.400 64.400 75.200 ;
        RECT 66.800 75.000 67.600 75.800 ;
        RECT 62.000 72.400 62.800 73.200 ;
        RECT 36.200 66.200 37.000 67.000 ;
        RECT 78.000 71.200 78.800 72.000 ;
        RECT 52.400 63.600 53.200 64.400 ;
        RECT 71.600 67.600 72.400 68.400 ;
        RECT 68.400 65.600 69.200 66.400 ;
        RECT 62.000 64.200 62.800 65.000 ;
        RECT 63.600 64.200 64.400 65.000 ;
        RECT 65.200 64.200 66.000 65.000 ;
        RECT 66.800 64.200 67.600 65.000 ;
        RECT 70.000 64.200 70.800 65.000 ;
        RECT 73.200 64.200 74.000 65.000 ;
        RECT 74.800 64.200 75.600 65.000 ;
        RECT 76.400 64.200 77.200 65.000 ;
        RECT 108.400 77.600 109.200 78.400 ;
        RECT 103.600 71.600 104.400 72.400 ;
        RECT 114.800 77.600 115.600 78.400 ;
        RECT 87.600 65.600 88.400 66.400 ;
        RECT 86.000 63.600 86.800 64.400 ;
        RECT 110.000 65.600 110.800 66.400 ;
        RECT 145.200 77.600 146.000 78.400 ;
        RECT 130.800 63.600 131.600 64.400 ;
        RECT 148.400 65.600 149.200 66.400 ;
        RECT 175.800 71.800 176.600 72.600 ;
        RECT 150.000 63.600 150.800 64.400 ;
        RECT 161.200 65.600 162.000 66.400 ;
        RECT 169.200 69.600 170.000 70.400 ;
        RECT 177.000 69.800 177.800 70.600 ;
        RECT 175.800 66.200 176.600 67.000 ;
        RECT 183.600 67.600 184.400 68.400 ;
        RECT 191.600 77.600 192.400 78.400 ;
        RECT 202.800 65.600 203.600 66.400 ;
        RECT 204.400 63.600 205.200 64.400 ;
        RECT 210.800 69.600 211.600 70.400 ;
        RECT 209.200 65.600 210.000 66.400 ;
        RECT 18.800 55.600 19.600 56.400 ;
        RECT 20.400 54.200 21.200 55.000 ;
        RECT 2.800 43.600 3.600 44.400 ;
        RECT 14.000 46.800 14.800 47.600 ;
        RECT 17.200 46.200 18.000 47.000 ;
        RECT 12.400 44.200 13.200 45.000 ;
        RECT 14.000 44.200 14.800 45.000 ;
        RECT 15.600 44.200 16.400 45.000 ;
        RECT 20.400 46.200 21.200 47.000 ;
        RECT 23.600 46.200 24.400 47.000 ;
        RECT 36.400 49.600 37.200 50.400 ;
        RECT 25.200 44.200 26.000 45.000 ;
        RECT 26.800 44.200 27.600 45.000 ;
        RECT 49.200 43.600 50.000 44.400 ;
        RECT 82.800 57.600 83.600 58.400 ;
        RECT 92.400 57.600 93.200 58.400 ;
        RECT 71.600 47.600 72.400 48.400 ;
        RECT 92.400 53.600 93.200 54.400 ;
        RECT 90.800 51.600 91.600 52.400 ;
        RECT 102.000 49.600 102.800 50.400 ;
        RECT 106.800 49.600 107.600 50.400 ;
        RECT 113.200 53.600 114.000 54.400 ;
        RECT 111.600 51.600 112.400 52.400 ;
        RECT 132.400 53.000 133.200 53.800 ;
        RECT 122.800 51.600 123.600 52.400 ;
        RECT 142.000 52.600 142.800 53.400 ;
        RECT 130.800 51.600 131.600 52.400 ;
        RECT 148.400 51.600 149.200 52.400 ;
        RECT 134.000 48.800 134.800 49.600 ;
        RECT 138.800 47.600 139.600 48.400 ;
        RECT 122.800 43.600 123.600 44.400 ;
        RECT 135.600 46.200 136.400 47.000 ;
        RECT 132.400 44.200 133.200 45.000 ;
        RECT 134.000 44.200 134.800 45.000 ;
        RECT 138.800 46.200 139.600 47.000 ;
        RECT 142.000 46.200 142.800 47.000 ;
        RECT 143.600 44.200 144.400 45.000 ;
        RECT 145.200 44.200 146.000 45.000 ;
        RECT 146.800 44.200 147.600 45.000 ;
        RECT 172.400 53.000 173.200 53.800 ;
        RECT 182.000 52.600 182.800 53.400 ;
        RECT 167.600 51.600 168.400 52.400 ;
        RECT 170.800 51.600 171.600 52.400 ;
        RECT 199.600 51.600 200.400 52.400 ;
        RECT 174.000 48.800 174.800 49.600 ;
        RECT 178.800 47.600 179.600 48.400 ;
        RECT 175.600 46.200 176.400 47.000 ;
        RECT 172.400 44.200 173.200 45.000 ;
        RECT 174.000 44.200 174.800 45.000 ;
        RECT 178.800 46.200 179.600 47.000 ;
        RECT 182.000 46.200 182.800 47.000 ;
        RECT 183.600 44.200 184.400 45.000 ;
        RECT 185.200 44.200 186.000 45.000 ;
        RECT 186.800 44.200 187.600 45.000 ;
        RECT 196.400 47.600 197.200 48.400 ;
        RECT 210.800 53.600 211.600 54.400 ;
        RECT 12.400 37.600 13.200 38.400 ;
        RECT 10.800 33.600 11.600 34.400 ;
        RECT 4.400 29.600 5.200 30.400 ;
        RECT 7.600 29.600 8.400 30.400 ;
        RECT 6.000 25.600 6.800 26.400 ;
        RECT 20.400 31.800 21.200 32.600 ;
        RECT 46.000 37.600 46.800 38.400 ;
        RECT 49.200 37.600 50.000 38.400 ;
        RECT 12.400 29.600 13.200 30.400 ;
        RECT 20.400 26.200 21.200 27.000 ;
        RECT 25.200 26.400 26.000 27.200 ;
        RECT 25.200 23.600 26.000 24.400 ;
        RECT 52.400 27.600 53.200 28.400 ;
        RECT 50.800 25.600 51.600 26.400 ;
        RECT 63.400 31.800 64.200 32.600 ;
        RECT 63.400 26.200 64.200 27.000 ;
        RECT 90.800 35.000 91.600 35.800 ;
        RECT 87.600 33.600 88.400 34.400 ;
        RECT 105.200 37.600 106.000 38.400 ;
        RECT 92.400 32.400 93.200 33.200 ;
        RECT 110.000 37.600 110.800 38.400 ;
        RECT 71.600 27.600 72.400 28.400 ;
        RECT 81.200 28.200 82.000 29.000 ;
        RECT 90.800 28.600 91.600 29.400 ;
        RECT 86.000 27.600 86.800 28.400 ;
        RECT 81.200 24.200 82.000 25.000 ;
        RECT 82.800 24.200 83.600 25.000 ;
        RECT 84.400 24.200 85.200 25.000 ;
        RECT 87.600 24.200 88.400 25.000 ;
        RECT 90.800 24.200 91.600 25.000 ;
        RECT 92.400 24.200 93.200 25.000 ;
        RECT 94.000 24.200 94.800 25.000 ;
        RECT 95.600 24.200 96.400 25.000 ;
        RECT 121.200 34.400 122.000 35.200 ;
        RECT 124.400 35.000 125.200 35.800 ;
        RECT 119.600 32.400 120.400 33.200 ;
        RECT 135.600 31.200 136.400 32.000 ;
        RECT 138.800 31.600 139.600 32.400 ;
        RECT 110.000 23.600 110.800 24.400 ;
        RECT 129.200 27.600 130.000 28.400 ;
        RECT 126.000 25.600 126.800 26.400 ;
        RECT 119.600 24.200 120.400 25.000 ;
        RECT 121.200 24.200 122.000 25.000 ;
        RECT 122.800 24.200 123.600 25.000 ;
        RECT 124.400 24.200 125.200 25.000 ;
        RECT 127.600 24.200 128.400 25.000 ;
        RECT 130.800 24.200 131.600 25.000 ;
        RECT 132.400 24.200 133.200 25.000 ;
        RECT 134.000 24.200 134.800 25.000 ;
        RECT 143.600 27.600 144.400 28.400 ;
        RECT 159.600 37.600 160.400 38.400 ;
        RECT 146.800 23.600 147.600 24.400 ;
        RECT 151.600 25.600 152.400 26.400 ;
        RECT 158.000 25.600 158.800 26.400 ;
        RECT 183.600 35.000 184.400 35.800 ;
        RECT 180.400 33.600 181.200 34.400 ;
        RECT 198.000 37.600 198.800 38.400 ;
        RECT 185.200 32.400 186.000 33.200 ;
        RECT 203.000 31.800 203.800 32.600 ;
        RECT 174.000 28.200 174.800 29.000 ;
        RECT 183.600 28.600 184.400 29.400 ;
        RECT 164.400 25.600 165.200 26.400 ;
        RECT 162.800 23.600 163.600 24.400 ;
        RECT 178.800 27.600 179.600 28.400 ;
        RECT 174.000 24.200 174.800 25.000 ;
        RECT 175.600 24.200 176.400 25.000 ;
        RECT 177.200 24.200 178.000 25.000 ;
        RECT 180.400 24.200 181.200 25.000 ;
        RECT 183.600 24.200 184.400 25.000 ;
        RECT 185.200 24.200 186.000 25.000 ;
        RECT 186.800 24.200 187.600 25.000 ;
        RECT 188.400 24.200 189.200 25.000 ;
        RECT 204.200 29.800 205.000 30.600 ;
        RECT 212.400 29.600 213.200 30.400 ;
        RECT 203.000 26.200 203.800 27.000 ;
        RECT 7.600 17.600 8.400 18.400 ;
        RECT 23.600 15.600 24.400 16.400 ;
        RECT 25.200 14.200 26.000 15.000 ;
        RECT 33.200 11.600 34.000 12.400 ;
        RECT 18.800 6.800 19.600 7.600 ;
        RECT 22.000 6.200 22.800 7.000 ;
        RECT 17.200 4.200 18.000 5.000 ;
        RECT 18.800 4.200 19.600 5.000 ;
        RECT 20.400 4.200 21.200 5.000 ;
        RECT 25.200 6.200 26.000 7.000 ;
        RECT 28.400 6.200 29.200 7.000 ;
        RECT 68.400 15.600 69.200 16.400 ;
        RECT 70.000 14.200 70.800 15.000 ;
        RECT 60.400 11.600 61.200 12.400 ;
        RECT 78.000 11.600 78.800 12.400 ;
        RECT 30.000 4.200 30.800 5.000 ;
        RECT 31.600 4.200 32.400 5.000 ;
        RECT 63.600 6.800 64.400 7.600 ;
        RECT 66.800 6.200 67.600 7.000 ;
        RECT 62.000 4.200 62.800 5.000 ;
        RECT 63.600 4.200 64.400 5.000 ;
        RECT 65.200 4.200 66.000 5.000 ;
        RECT 70.000 6.200 70.800 7.000 ;
        RECT 73.200 6.200 74.000 7.000 ;
        RECT 106.800 17.600 107.600 18.400 ;
        RECT 122.800 15.600 123.600 16.400 ;
        RECT 124.400 14.200 125.200 15.000 ;
        RECT 135.600 11.600 136.400 12.400 ;
        RECT 74.800 4.200 75.600 5.000 ;
        RECT 76.400 4.200 77.200 5.000 ;
        RECT 118.000 6.800 118.800 7.600 ;
        RECT 121.200 6.200 122.000 7.000 ;
        RECT 116.400 4.200 117.200 5.000 ;
        RECT 118.000 4.200 118.800 5.000 ;
        RECT 119.600 4.200 120.400 5.000 ;
        RECT 124.400 6.200 125.200 7.000 ;
        RECT 127.600 6.200 128.400 7.000 ;
        RECT 162.800 15.600 163.600 16.400 ;
        RECT 164.400 14.200 165.200 15.000 ;
        RECT 174.000 11.600 174.800 12.400 ;
        RECT 129.200 4.200 130.000 5.000 ;
        RECT 130.800 4.200 131.600 5.000 ;
        RECT 158.000 6.800 158.800 7.600 ;
        RECT 161.200 6.200 162.000 7.000 ;
        RECT 156.400 4.200 157.200 5.000 ;
        RECT 158.000 4.200 158.800 5.000 ;
        RECT 159.600 4.200 160.400 5.000 ;
        RECT 164.400 6.200 165.200 7.000 ;
        RECT 167.600 6.200 168.400 7.000 ;
        RECT 188.400 13.000 189.200 13.800 ;
        RECT 198.000 12.600 198.800 13.400 ;
        RECT 212.400 17.600 213.200 18.400 ;
        RECT 183.600 11.600 184.400 12.400 ;
        RECT 190.000 8.800 190.800 9.600 ;
        RECT 194.800 7.600 195.600 8.400 ;
        RECT 169.200 4.200 170.000 5.000 ;
        RECT 170.800 4.200 171.600 5.000 ;
        RECT 191.600 6.200 192.400 7.000 ;
        RECT 188.400 4.200 189.200 5.000 ;
        RECT 190.000 4.200 190.800 5.000 ;
        RECT 194.800 6.200 195.600 7.000 ;
        RECT 198.000 6.200 198.800 7.000 ;
        RECT 199.600 4.200 200.400 5.000 ;
        RECT 201.200 4.200 202.000 5.000 ;
        RECT 202.800 4.200 203.600 5.000 ;
      LAYER metal2 ;
        RECT 50.800 193.600 51.600 194.400 ;
        RECT 54.000 193.600 54.800 194.400 ;
        RECT 7.800 191.800 8.600 192.600 ;
        RECT 14.000 191.800 14.800 192.600 ;
        RECT 4.400 189.600 5.200 190.400 ;
        RECT 4.500 186.400 5.100 189.600 ;
        RECT 7.800 187.000 8.400 191.800 ;
        RECT 9.000 189.800 9.800 190.600 ;
        RECT 9.200 188.400 9.800 189.800 ;
        RECT 14.200 188.400 14.800 191.800 ;
        RECT 34.800 191.600 35.600 192.400 ;
        RECT 47.600 191.600 48.400 192.400 ;
        RECT 60.400 191.600 61.200 192.400 ;
        RECT 22.000 189.600 22.800 190.400 ;
        RECT 26.800 189.600 27.600 190.400 ;
        RECT 38.000 189.600 38.800 190.400 ;
        RECT 38.100 188.400 38.700 189.600 ;
        RECT 9.200 187.800 14.800 188.400 ;
        RECT 9.200 187.000 10.000 187.200 ;
        RECT 12.600 187.000 13.400 187.200 ;
        RECT 14.200 187.000 14.800 187.800 ;
        RECT 28.400 187.600 29.200 188.400 ;
        RECT 38.000 187.600 38.800 188.400 ;
        RECT 46.000 187.600 46.800 188.400 ;
        RECT 7.800 186.400 13.400 187.000 ;
        RECT 4.400 185.600 5.200 186.400 ;
        RECT 7.800 186.200 8.600 186.400 ;
        RECT 14.000 186.200 14.800 187.000 ;
        RECT 47.700 186.400 48.300 191.600 ;
        RECT 49.200 189.600 50.000 190.400 ;
        RECT 55.600 189.600 56.400 190.400 ;
        RECT 68.200 189.600 69.200 190.400 ;
        RECT 49.300 188.400 49.900 189.600 ;
        RECT 49.200 187.600 50.000 188.400 ;
        RECT 52.400 187.600 53.200 188.400 ;
        RECT 55.700 186.400 56.300 189.600 ;
        RECT 57.200 187.600 58.000 188.400 ;
        RECT 58.800 187.600 59.600 188.400 ;
        RECT 17.200 185.600 18.000 186.400 ;
        RECT 28.400 185.600 29.200 186.400 ;
        RECT 44.400 185.600 45.200 186.400 ;
        RECT 47.600 185.600 48.400 186.400 ;
        RECT 55.600 185.600 56.400 186.400 ;
        RECT 4.500 180.300 5.100 185.600 ;
        RECT 10.800 183.600 11.600 184.400 ;
        RECT 17.300 182.400 17.900 185.600 ;
        RECT 22.000 183.600 22.800 184.400 ;
        RECT 28.400 183.600 29.200 184.400 ;
        RECT 17.200 181.600 18.000 182.400 ;
        RECT 2.900 179.700 5.100 180.300 ;
        RECT 2.900 178.400 3.500 179.700 ;
        RECT 2.800 177.600 3.600 178.400 ;
        RECT 12.400 164.200 13.200 177.800 ;
        RECT 14.000 164.200 14.800 177.800 ;
        RECT 15.600 164.200 16.400 177.800 ;
        RECT 17.200 166.200 18.000 177.800 ;
        RECT 18.800 175.600 19.600 176.400 ;
        RECT 18.900 152.300 19.500 175.600 ;
        RECT 20.400 166.200 21.200 177.800 ;
        RECT 22.100 174.400 22.700 183.600 ;
        RECT 22.000 173.600 22.800 174.400 ;
        RECT 23.600 166.200 24.400 177.800 ;
        RECT 25.200 164.200 26.000 177.800 ;
        RECT 26.800 164.200 27.600 177.800 ;
        RECT 28.500 168.400 29.100 183.600 ;
        RECT 39.600 175.600 40.400 176.400 ;
        RECT 49.200 175.600 50.000 176.400 ;
        RECT 52.400 175.600 53.200 176.400 ;
        RECT 39.700 172.400 40.300 175.600 ;
        RECT 39.600 171.600 40.400 172.400 ;
        RECT 44.400 171.600 45.200 172.400 ;
        RECT 47.600 171.600 48.400 172.400 ;
        RECT 49.300 170.400 49.900 175.600 ;
        RECT 57.300 172.400 57.900 187.600 ;
        RECT 78.000 184.200 78.800 197.800 ;
        RECT 79.600 184.200 80.400 197.800 ;
        RECT 81.200 184.200 82.000 197.800 ;
        RECT 82.800 184.200 83.600 195.800 ;
        RECT 84.400 185.600 85.200 186.400 ;
        RECT 84.500 182.400 85.100 185.600 ;
        RECT 86.000 184.200 86.800 195.800 ;
        RECT 87.600 187.600 88.400 188.400 ;
        RECT 89.200 184.200 90.000 195.800 ;
        RECT 90.800 184.200 91.600 197.800 ;
        RECT 92.400 184.200 93.200 197.800 ;
        RECT 97.200 189.600 98.000 190.400 ;
        RECT 102.000 189.600 102.800 190.400 ;
        RECT 110.000 189.600 110.800 190.400 ;
        RECT 84.400 181.600 85.200 182.400 ;
        RECT 90.800 181.600 91.600 182.400 ;
        RECT 95.600 181.600 96.400 182.400 ;
        RECT 90.900 178.400 91.500 181.600 ;
        RECT 68.400 178.300 69.200 178.400 ;
        RECT 66.900 177.700 69.200 178.300 ;
        RECT 55.600 171.600 56.400 172.400 ;
        RECT 57.200 171.600 58.000 172.400 ;
        RECT 31.600 169.600 32.400 170.400 ;
        RECT 46.000 169.600 46.800 170.400 ;
        RECT 49.200 169.600 50.000 170.400 ;
        RECT 54.000 169.600 54.800 170.400 ;
        RECT 28.400 167.600 29.200 168.400 ;
        RECT 20.400 153.600 21.200 154.400 ;
        RECT 18.900 151.700 21.100 152.300 ;
        RECT 4.400 149.600 5.200 150.400 ;
        RECT 9.200 149.600 10.000 150.400 ;
        RECT 14.000 149.600 14.800 150.400 ;
        RECT 18.800 149.600 19.600 150.400 ;
        RECT 4.500 146.400 5.100 149.600 ;
        RECT 9.300 148.400 9.900 149.600 ;
        RECT 9.200 147.600 10.000 148.400 ;
        RECT 14.000 147.600 14.800 148.400 ;
        RECT 20.500 148.300 21.100 151.700 ;
        RECT 28.400 151.600 29.200 152.400 ;
        RECT 18.900 147.700 21.100 148.300 ;
        RECT 14.100 146.400 14.700 147.600 ;
        RECT 4.400 146.300 5.200 146.400 ;
        RECT 2.900 145.700 5.200 146.300 ;
        RECT 2.900 138.400 3.500 145.700 ;
        RECT 4.400 145.600 5.200 145.700 ;
        RECT 10.800 145.600 11.600 146.400 ;
        RECT 14.000 145.600 14.800 146.400 ;
        RECT 18.900 138.400 19.500 147.700 ;
        RECT 28.500 146.400 29.100 151.600 ;
        RECT 25.200 145.600 26.000 146.400 ;
        RECT 28.400 145.600 29.200 146.400 ;
        RECT 25.300 144.400 25.900 145.600 ;
        RECT 20.400 143.600 21.200 144.400 ;
        RECT 22.000 143.600 22.800 144.400 ;
        RECT 25.200 143.600 26.000 144.400 ;
        RECT 2.800 137.600 3.600 138.400 ;
        RECT 12.400 124.200 13.200 137.800 ;
        RECT 14.000 124.200 14.800 137.800 ;
        RECT 15.600 124.200 16.400 137.800 ;
        RECT 17.200 126.200 18.000 137.800 ;
        RECT 18.800 137.600 19.600 138.400 ;
        RECT 18.900 136.400 19.500 137.600 ;
        RECT 18.800 135.600 19.600 136.400 ;
        RECT 20.400 126.200 21.200 137.800 ;
        RECT 22.100 134.400 22.700 143.600 ;
        RECT 22.000 133.600 22.800 134.400 ;
        RECT 23.600 126.200 24.400 137.800 ;
        RECT 25.200 124.200 26.000 137.800 ;
        RECT 26.800 124.200 27.600 137.800 ;
        RECT 31.700 132.400 32.300 169.600 ;
        RECT 46.100 168.400 46.700 169.600 ;
        RECT 42.800 167.600 43.600 168.400 ;
        RECT 46.000 167.600 46.800 168.400 ;
        RECT 49.200 167.600 50.000 168.400 ;
        RECT 41.200 163.600 42.000 164.400 ;
        RECT 41.300 152.400 41.900 163.600 ;
        RECT 34.800 151.600 35.600 152.400 ;
        RECT 41.200 151.600 42.000 152.400 ;
        RECT 38.000 149.600 38.800 150.400 ;
        RECT 38.100 148.400 38.700 149.600 ;
        RECT 34.800 147.600 35.600 148.400 ;
        RECT 36.400 147.600 37.200 148.400 ;
        RECT 38.000 147.600 38.800 148.400 ;
        RECT 34.900 146.300 35.500 147.600 ;
        RECT 34.900 145.700 37.100 146.300 ;
        RECT 36.500 136.400 37.100 145.700 ;
        RECT 38.000 145.600 38.800 146.400 ;
        RECT 36.400 135.600 37.200 136.400 ;
        RECT 38.100 134.400 38.700 145.600 ;
        RECT 41.300 134.400 41.900 151.600 ;
        RECT 46.000 151.200 46.800 152.000 ;
        RECT 38.000 133.600 38.800 134.400 ;
        RECT 41.200 133.600 42.000 134.400 ;
        RECT 41.300 132.400 41.900 133.600 ;
        RECT 46.100 132.400 46.700 151.200 ;
        RECT 47.600 144.200 48.400 157.800 ;
        RECT 49.200 144.200 50.000 157.800 ;
        RECT 50.800 144.200 51.600 155.800 ;
        RECT 52.400 147.600 53.200 148.400 ;
        RECT 54.000 144.200 54.800 155.800 ;
        RECT 55.700 150.400 56.300 171.600 ;
        RECT 55.600 149.600 56.400 150.400 ;
        RECT 55.600 145.600 56.400 146.400 ;
        RECT 55.700 138.400 56.300 145.600 ;
        RECT 57.200 144.200 58.000 155.800 ;
        RECT 58.800 144.200 59.600 157.800 ;
        RECT 60.400 144.200 61.200 157.800 ;
        RECT 62.000 144.200 62.800 157.800 ;
        RECT 66.900 154.400 67.500 177.700 ;
        RECT 68.400 177.600 69.200 177.700 ;
        RECT 90.800 177.600 91.600 178.400 ;
        RECT 68.400 175.600 69.200 176.400 ;
        RECT 79.400 175.000 80.200 175.800 ;
        RECT 81.200 175.000 85.400 175.600 ;
        RECT 86.000 175.000 86.800 175.800 ;
        RECT 87.600 175.600 88.400 176.400 ;
        RECT 68.400 173.600 69.200 174.400 ;
        RECT 70.000 173.600 70.800 174.400 ;
        RECT 78.000 173.600 78.800 174.400 ;
        RECT 68.500 170.400 69.100 173.600 ;
        RECT 70.100 172.400 70.700 173.600 ;
        RECT 70.000 171.600 70.800 172.400 ;
        RECT 68.400 169.600 69.200 170.400 ;
        RECT 71.600 169.600 72.400 170.400 ;
        RECT 79.400 170.200 80.000 175.000 ;
        RECT 81.200 174.800 82.000 175.000 ;
        RECT 84.600 174.800 85.400 175.000 ;
        RECT 86.200 174.200 86.800 175.000 ;
        RECT 87.700 174.400 88.300 175.600 ;
        RECT 82.000 173.600 86.800 174.200 ;
        RECT 87.600 173.600 88.400 174.400 ;
        RECT 82.000 173.400 82.800 173.600 ;
        RECT 86.200 170.200 86.800 173.600 ;
        RECT 71.700 158.400 72.300 169.600 ;
        RECT 79.400 169.400 80.200 170.200 ;
        RECT 86.000 169.400 86.800 170.200 ;
        RECT 82.800 163.600 83.600 164.400 ;
        RECT 71.600 157.600 72.400 158.400 ;
        RECT 66.800 153.600 67.600 154.400 ;
        RECT 82.900 148.400 83.500 163.600 ;
        RECT 86.000 151.200 86.800 152.000 ;
        RECT 82.800 147.600 83.600 148.400 ;
        RECT 82.800 145.600 83.600 146.400 ;
        RECT 55.600 137.600 56.400 138.400 ;
        RECT 50.600 135.000 51.400 135.800 ;
        RECT 52.400 135.000 56.600 135.600 ;
        RECT 57.200 135.000 58.000 135.800 ;
        RECT 58.800 135.600 59.600 136.400 ;
        RECT 49.200 133.600 50.000 134.400 ;
        RECT 31.600 131.600 32.400 132.400 ;
        RECT 41.200 131.600 42.000 132.400 ;
        RECT 46.000 131.600 46.800 132.400 ;
        RECT 44.400 129.800 45.200 130.600 ;
        RECT 9.200 117.600 10.000 118.400 ;
        RECT 9.300 110.400 9.900 117.600 ;
        RECT 44.500 114.400 45.100 129.800 ;
        RECT 31.600 113.600 32.400 114.400 ;
        RECT 44.400 113.600 45.200 114.400 ;
        RECT 12.400 111.800 13.200 112.600 ;
        RECT 19.000 111.800 19.800 112.600 ;
        RECT 4.400 110.300 5.200 110.400 ;
        RECT 2.900 109.700 5.200 110.300 ;
        RECT 2.900 98.400 3.500 109.700 ;
        RECT 4.400 109.600 5.200 109.700 ;
        RECT 9.200 109.600 10.000 110.400 ;
        RECT 4.500 108.400 5.100 109.600 ;
        RECT 12.400 108.400 13.000 111.800 ;
        RECT 16.400 108.400 17.200 108.600 ;
        RECT 4.400 107.600 5.200 108.400 ;
        RECT 10.800 107.600 11.600 108.400 ;
        RECT 12.400 107.800 17.200 108.400 ;
        RECT 12.400 107.000 13.000 107.800 ;
        RECT 13.800 107.000 14.600 107.200 ;
        RECT 17.200 107.000 18.000 107.200 ;
        RECT 19.200 107.000 19.800 111.800 ;
        RECT 23.600 111.600 24.400 112.400 ;
        RECT 28.400 111.600 29.200 112.400 ;
        RECT 46.100 110.400 46.700 131.600 ;
        RECT 50.600 130.200 51.200 135.000 ;
        RECT 52.400 134.800 53.200 135.000 ;
        RECT 55.800 134.800 56.600 135.000 ;
        RECT 57.400 134.200 58.000 135.000 ;
        RECT 58.900 134.400 59.500 135.600 ;
        RECT 53.200 133.600 58.000 134.200 ;
        RECT 58.800 133.600 59.600 134.400 ;
        RECT 53.200 133.400 54.000 133.600 ;
        RECT 57.400 130.200 58.000 133.600 ;
        RECT 50.600 129.400 51.400 130.200 ;
        RECT 57.200 129.400 58.000 130.200 ;
        RECT 54.000 127.600 54.800 128.400 ;
        RECT 76.400 124.200 77.200 137.800 ;
        RECT 78.000 124.200 78.800 137.800 ;
        RECT 79.600 124.200 80.400 137.800 ;
        RECT 81.200 126.200 82.000 137.800 ;
        RECT 82.900 136.400 83.500 145.600 ;
        RECT 86.100 142.400 86.700 151.200 ;
        RECT 87.600 144.200 88.400 157.800 ;
        RECT 89.200 144.200 90.000 157.800 ;
        RECT 90.800 144.200 91.600 155.800 ;
        RECT 92.400 147.600 93.200 148.400 ;
        RECT 94.000 144.200 94.800 155.800 ;
        RECT 95.700 146.400 96.300 181.600 ;
        RECT 102.100 176.400 102.700 189.600 ;
        RECT 102.000 175.600 102.800 176.400 ;
        RECT 108.400 175.600 109.200 176.400 ;
        RECT 108.500 158.400 109.100 175.600 ;
        RECT 110.100 172.400 110.700 189.600 ;
        RECT 114.800 184.200 115.600 197.800 ;
        RECT 116.400 184.200 117.200 197.800 ;
        RECT 118.000 184.200 118.800 195.800 ;
        RECT 119.600 191.600 120.400 192.400 ;
        RECT 119.700 188.400 120.300 191.600 ;
        RECT 119.600 187.600 120.400 188.400 ;
        RECT 119.600 185.600 120.400 186.400 ;
        RECT 110.000 171.600 110.800 172.400 ;
        RECT 95.600 145.600 96.400 146.400 ;
        RECT 86.000 141.600 86.800 142.400 ;
        RECT 92.400 141.600 93.200 142.400 ;
        RECT 82.800 135.600 83.600 136.400 ;
        RECT 84.400 126.200 85.200 137.800 ;
        RECT 86.000 133.600 86.800 134.400 ;
        RECT 86.100 128.400 86.700 133.600 ;
        RECT 86.000 127.600 86.800 128.400 ;
        RECT 87.600 126.200 88.400 137.800 ;
        RECT 89.200 124.200 90.000 137.800 ;
        RECT 90.800 124.200 91.600 137.800 ;
        RECT 92.500 130.800 93.100 141.600 ;
        RECT 95.700 136.400 96.300 145.600 ;
        RECT 97.200 144.200 98.000 155.800 ;
        RECT 98.800 144.200 99.600 157.800 ;
        RECT 100.400 144.200 101.200 157.800 ;
        RECT 102.000 144.200 102.800 157.800 ;
        RECT 108.400 157.600 109.200 158.400 ;
        RECT 110.100 148.400 110.700 171.600 ;
        RECT 111.600 164.200 112.400 177.800 ;
        RECT 113.200 164.200 114.000 177.800 ;
        RECT 114.800 166.200 115.600 177.800 ;
        RECT 116.400 173.600 117.200 174.400 ;
        RECT 116.500 170.400 117.100 173.600 ;
        RECT 116.400 169.600 117.200 170.400 ;
        RECT 118.000 166.200 118.800 177.800 ;
        RECT 119.700 176.400 120.300 185.600 ;
        RECT 121.200 184.200 122.000 195.800 ;
        RECT 122.800 185.600 123.600 186.400 ;
        RECT 124.400 184.200 125.200 195.800 ;
        RECT 126.000 184.200 126.800 197.800 ;
        RECT 127.600 184.200 128.400 197.800 ;
        RECT 129.200 184.200 130.000 197.800 ;
        RECT 148.400 191.800 149.200 192.600 ;
        RECT 138.800 189.600 139.800 190.400 ;
        RECT 145.200 189.600 146.000 190.400 ;
        RECT 148.400 188.400 149.000 191.800 ;
        RECT 150.000 191.600 150.800 192.400 ;
        RECT 155.000 191.800 155.800 192.600 ;
        RECT 152.400 188.400 153.200 188.600 ;
        RECT 148.400 187.800 153.200 188.400 ;
        RECT 148.400 187.000 149.000 187.800 ;
        RECT 149.800 187.000 150.600 187.200 ;
        RECT 153.200 187.000 154.000 187.200 ;
        RECT 155.200 187.000 155.800 191.800 ;
        RECT 162.800 189.600 163.600 190.400 ;
        RECT 167.600 189.600 168.400 190.400 ;
        RECT 170.800 189.600 171.600 190.400 ;
        RECT 174.000 189.600 174.800 190.400 ;
        RECT 185.200 189.600 186.000 190.400 ;
        RECT 156.400 187.600 157.200 188.400 ;
        RECT 148.400 186.200 149.200 187.000 ;
        RECT 149.800 186.400 154.000 187.000 ;
        RECT 155.000 186.200 155.800 187.000 ;
        RECT 119.600 175.600 120.400 176.400 ;
        RECT 111.600 157.600 112.400 158.400 ;
        RECT 110.000 147.600 110.800 148.400 ;
        RECT 113.200 147.600 114.000 148.400 ;
        RECT 113.300 138.400 113.900 147.600 ;
        RECT 119.700 146.400 120.300 175.600 ;
        RECT 121.200 166.200 122.000 177.800 ;
        RECT 122.800 164.200 123.600 177.800 ;
        RECT 124.400 164.200 125.200 177.800 ;
        RECT 126.000 164.200 126.800 177.800 ;
        RECT 161.200 177.600 162.000 178.400 ;
        RECT 162.900 176.400 163.500 189.600 ;
        RECT 164.400 187.600 165.200 188.400 ;
        RECT 164.500 178.400 165.100 187.600 ;
        RECT 167.700 186.400 168.300 189.600 ;
        RECT 177.200 188.000 178.000 188.800 ;
        RECT 167.600 185.600 168.400 186.400 ;
        RECT 170.800 185.600 171.600 186.400 ;
        RECT 170.900 178.400 171.500 185.600 ;
        RECT 172.400 183.600 173.200 184.400 ;
        RECT 172.500 180.400 173.100 183.600 ;
        RECT 177.300 182.400 177.900 188.000 ;
        RECT 180.400 183.600 181.200 184.400 ;
        RECT 177.200 181.600 178.000 182.400 ;
        RECT 172.400 179.600 173.200 180.400 ;
        RECT 178.800 179.600 179.600 180.400 ;
        RECT 164.400 177.600 165.200 178.400 ;
        RECT 170.800 177.600 171.600 178.400 ;
        RECT 135.600 175.600 136.400 176.400 ;
        RECT 145.000 175.000 145.800 175.800 ;
        RECT 146.800 175.000 151.000 175.600 ;
        RECT 151.600 175.000 152.400 175.800 ;
        RECT 159.600 175.600 160.400 176.400 ;
        RECT 162.800 175.600 163.600 176.400 ;
        RECT 166.000 175.600 166.800 176.400 ;
        RECT 167.600 175.600 168.400 176.400 ;
        RECT 143.600 173.600 144.400 174.400 ;
        RECT 142.000 171.600 142.800 172.400 ;
        RECT 145.000 170.200 145.600 175.000 ;
        RECT 146.800 174.800 147.600 175.000 ;
        RECT 150.200 174.800 151.000 175.000 ;
        RECT 151.800 174.200 152.400 175.000 ;
        RECT 166.100 174.400 166.700 175.600 ;
        RECT 167.700 174.400 168.300 175.600 ;
        RECT 169.200 175.000 170.000 175.800 ;
        RECT 170.600 175.000 174.800 175.600 ;
        RECT 175.800 175.000 176.600 175.800 ;
        RECT 147.600 173.600 152.400 174.200 ;
        RECT 162.800 173.600 163.600 174.400 ;
        RECT 166.000 173.600 166.800 174.400 ;
        RECT 167.600 173.600 168.400 174.400 ;
        RECT 169.200 174.200 169.800 175.000 ;
        RECT 170.600 174.800 171.400 175.000 ;
        RECT 174.000 174.800 174.800 175.000 ;
        RECT 169.200 173.600 174.000 174.200 ;
        RECT 147.600 173.400 148.400 173.600 ;
        RECT 145.000 169.400 145.800 170.200 ;
        RECT 146.800 169.600 147.600 170.400 ;
        RECT 151.800 170.200 152.400 173.600 ;
        RECT 162.900 170.400 163.500 173.600 ;
        RECT 146.900 168.400 147.500 169.600 ;
        RECT 151.600 169.400 152.400 170.200 ;
        RECT 162.800 169.600 163.600 170.400 ;
        RECT 146.800 167.600 147.600 168.400 ;
        RECT 132.400 149.600 133.200 150.400 ;
        RECT 132.500 148.400 133.100 149.600 ;
        RECT 127.600 147.600 128.400 148.400 ;
        RECT 132.400 147.600 133.200 148.400 ;
        RECT 127.700 146.400 128.300 147.600 ;
        RECT 119.600 145.600 120.400 146.400 ;
        RECT 127.600 145.600 128.400 146.400 ;
        RECT 137.200 144.200 138.000 157.800 ;
        RECT 138.800 144.200 139.600 157.800 ;
        RECT 140.400 144.200 141.200 155.800 ;
        RECT 142.000 147.600 142.800 148.400 ;
        RECT 143.600 144.200 144.400 155.800 ;
        RECT 145.200 145.600 146.000 146.400 ;
        RECT 145.300 140.400 145.900 145.600 ;
        RECT 146.800 144.200 147.600 155.800 ;
        RECT 148.400 144.200 149.200 157.800 ;
        RECT 150.000 144.200 150.800 157.800 ;
        RECT 151.600 144.200 152.400 157.800 ;
        RECT 161.200 157.600 162.000 158.400 ;
        RECT 162.900 154.400 163.500 169.600 ;
        RECT 167.700 158.400 168.300 173.600 ;
        RECT 169.200 170.200 169.800 173.600 ;
        RECT 173.200 173.400 174.000 173.600 ;
        RECT 176.000 170.200 176.600 175.000 ;
        RECT 178.900 174.400 179.500 179.600 ;
        RECT 178.800 173.600 179.600 174.400 ;
        RECT 177.200 171.600 178.000 172.400 ;
        RECT 169.200 169.400 170.000 170.200 ;
        RECT 175.800 169.400 176.600 170.200 ;
        RECT 170.800 163.600 171.600 164.400 ;
        RECT 167.600 157.600 168.400 158.400 ;
        RECT 162.800 153.600 163.600 154.400 ;
        RECT 169.200 151.600 170.000 152.400 ;
        RECT 153.200 149.600 154.000 150.400 ;
        RECT 145.200 139.600 146.000 140.400 ;
        RECT 150.000 139.600 150.800 140.400 ;
        RECT 113.200 137.600 114.000 138.400 ;
        RECT 95.600 135.600 96.400 136.400 ;
        RECT 102.000 135.000 102.800 135.800 ;
        RECT 103.400 135.000 107.600 135.600 ;
        RECT 108.600 135.000 109.400 135.800 ;
        RECT 100.400 133.600 101.200 134.400 ;
        RECT 102.000 134.200 102.600 135.000 ;
        RECT 103.400 134.800 104.200 135.000 ;
        RECT 106.800 134.800 107.600 135.000 ;
        RECT 102.000 133.600 106.800 134.200 ;
        RECT 92.400 130.000 93.200 130.800 ;
        RECT 92.500 122.300 93.100 130.000 ;
        RECT 90.900 121.700 93.100 122.300 ;
        RECT 60.400 117.600 61.200 118.400 ;
        RECT 26.800 109.600 27.600 110.400 ;
        RECT 30.000 109.600 30.800 110.400 ;
        RECT 39.600 109.600 40.400 110.400 ;
        RECT 46.000 109.600 46.800 110.400 ;
        RECT 58.800 109.600 59.600 110.400 ;
        RECT 68.400 109.600 69.200 110.400 ;
        RECT 20.400 107.600 21.200 108.400 ;
        RECT 22.000 107.600 22.800 108.400 ;
        RECT 12.400 106.200 13.200 107.000 ;
        RECT 13.800 106.400 18.000 107.000 ;
        RECT 19.000 106.200 19.800 107.000 ;
        RECT 15.600 103.600 16.400 104.400 ;
        RECT 20.500 102.400 21.100 107.600 ;
        RECT 22.100 106.400 22.700 107.600 ;
        RECT 22.000 105.600 22.800 106.400 ;
        RECT 25.200 105.600 26.000 106.400 ;
        RECT 22.000 103.600 22.800 104.400 ;
        RECT 20.400 101.600 21.200 102.400 ;
        RECT 2.800 97.600 3.600 98.400 ;
        RECT 2.800 83.600 3.600 84.400 ;
        RECT 12.400 84.200 13.200 97.800 ;
        RECT 14.000 84.200 14.800 97.800 ;
        RECT 15.600 84.200 16.400 97.800 ;
        RECT 17.200 86.200 18.000 97.800 ;
        RECT 18.800 95.600 19.600 96.400 ;
        RECT 2.900 68.400 3.500 83.600 ;
        RECT 4.400 71.600 5.200 72.400 ;
        RECT 10.800 71.600 11.600 72.400 ;
        RECT 4.500 70.400 5.100 71.600 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 9.200 69.600 10.000 70.400 ;
        RECT 2.800 67.600 3.600 68.400 ;
        RECT 9.300 56.400 9.900 69.600 ;
        RECT 10.900 68.400 11.500 71.600 ;
        RECT 15.600 69.600 16.400 70.400 ;
        RECT 10.800 67.600 11.600 68.400 ;
        RECT 15.600 67.600 16.400 68.400 ;
        RECT 15.700 66.400 16.300 67.600 ;
        RECT 18.900 66.400 19.500 95.600 ;
        RECT 20.400 86.200 21.200 97.800 ;
        RECT 22.100 94.400 22.700 103.600 ;
        RECT 25.300 102.400 25.900 105.600 ;
        RECT 33.200 103.600 34.000 104.400 ;
        RECT 25.200 101.600 26.000 102.400 ;
        RECT 22.000 93.600 22.800 94.400 ;
        RECT 23.600 86.200 24.400 97.800 ;
        RECT 25.200 84.200 26.000 97.800 ;
        RECT 26.800 84.200 27.600 97.800 ;
        RECT 30.000 93.600 30.800 94.400 ;
        RECT 30.100 74.400 30.700 93.600 ;
        RECT 31.600 89.600 32.400 90.400 ;
        RECT 30.000 73.600 30.800 74.400 ;
        RECT 28.400 71.600 29.200 72.400 ;
        RECT 25.200 69.600 26.000 70.400 ;
        RECT 23.600 67.600 24.400 68.400 ;
        RECT 15.600 65.600 16.400 66.400 ;
        RECT 18.800 65.600 19.600 66.400 ;
        RECT 14.000 63.600 14.800 64.400 ;
        RECT 14.100 60.400 14.700 63.600 ;
        RECT 14.000 59.600 14.800 60.400 ;
        RECT 9.200 55.600 10.000 56.400 ;
        RECT 2.800 43.600 3.600 44.400 ;
        RECT 12.400 44.200 13.200 57.800 ;
        RECT 14.000 44.200 14.800 57.800 ;
        RECT 15.600 44.200 16.400 57.800 ;
        RECT 17.200 46.200 18.000 57.800 ;
        RECT 18.900 56.400 19.500 65.600 ;
        RECT 18.800 55.600 19.600 56.400 ;
        RECT 20.400 46.200 21.200 57.800 ;
        RECT 22.000 53.600 22.800 54.400 ;
        RECT 23.600 46.200 24.400 57.800 ;
        RECT 25.200 44.200 26.000 57.800 ;
        RECT 26.800 44.200 27.600 57.800 ;
        RECT 30.000 51.600 30.800 52.400 ;
        RECT 2.900 32.300 3.500 43.600 ;
        RECT 12.400 41.600 13.200 42.400 ;
        RECT 12.500 38.400 13.100 41.600 ;
        RECT 12.400 37.600 13.200 38.400 ;
        RECT 10.800 33.600 11.600 34.400 ;
        RECT 4.400 32.300 5.200 32.400 ;
        RECT 2.900 31.700 5.200 32.300 ;
        RECT 4.400 31.600 5.200 31.700 ;
        RECT 20.400 31.800 21.200 32.600 ;
        RECT 27.000 31.800 27.800 32.600 ;
        RECT 4.500 30.400 5.100 31.600 ;
        RECT 4.400 30.300 5.200 30.400 ;
        RECT 4.400 29.700 6.700 30.300 ;
        RECT 4.400 29.600 5.200 29.700 ;
        RECT 6.100 26.400 6.700 29.700 ;
        RECT 7.600 29.600 8.400 30.400 ;
        RECT 12.400 29.600 13.200 30.400 ;
        RECT 20.400 28.400 21.000 31.800 ;
        RECT 24.400 28.400 25.200 28.600 ;
        RECT 7.600 27.600 8.400 28.400 ;
        RECT 18.800 27.600 19.600 28.400 ;
        RECT 20.400 27.800 25.200 28.400 ;
        RECT 6.000 25.600 6.800 26.400 ;
        RECT 7.700 18.400 8.300 27.600 ;
        RECT 20.400 27.000 21.000 27.800 ;
        RECT 21.800 27.000 22.600 27.200 ;
        RECT 25.200 27.000 26.000 27.200 ;
        RECT 27.200 27.000 27.800 31.800 ;
        RECT 30.100 30.400 30.700 51.600 ;
        RECT 31.700 50.400 32.300 89.600 ;
        RECT 33.300 72.400 33.900 103.600 ;
        RECT 38.000 101.600 38.800 102.400 ;
        RECT 38.100 98.400 38.700 101.600 ;
        RECT 38.000 97.600 38.800 98.400 ;
        RECT 39.700 96.400 40.300 109.600 ;
        RECT 58.900 108.400 59.500 109.600 ;
        RECT 58.800 107.600 59.600 108.400 ;
        RECT 54.000 105.600 54.800 106.400 ;
        RECT 44.400 103.600 45.200 104.400 ;
        RECT 39.600 95.600 40.400 96.400 ;
        RECT 44.500 84.400 45.100 103.600 ;
        RECT 38.000 83.600 38.800 84.400 ;
        RECT 44.400 83.600 45.200 84.400 ;
        RECT 47.600 84.200 48.400 97.800 ;
        RECT 49.200 84.200 50.000 97.800 ;
        RECT 50.800 84.200 51.600 97.800 ;
        RECT 52.400 86.200 53.200 97.800 ;
        RECT 54.100 96.400 54.700 105.600 ;
        RECT 70.000 104.200 70.800 117.800 ;
        RECT 71.600 104.200 72.400 117.800 ;
        RECT 73.200 104.200 74.000 117.800 ;
        RECT 74.800 104.200 75.600 115.800 ;
        RECT 76.400 105.600 77.200 106.400 ;
        RECT 78.000 104.200 78.800 115.800 ;
        RECT 79.600 109.600 80.400 110.400 ;
        RECT 79.700 108.400 80.300 109.600 ;
        RECT 79.600 107.600 80.400 108.400 ;
        RECT 81.200 104.200 82.000 115.800 ;
        RECT 82.800 104.200 83.600 117.800 ;
        RECT 84.400 104.200 85.200 117.800 ;
        RECT 90.900 110.400 91.500 121.700 ;
        RECT 100.500 118.400 101.100 133.600 ;
        RECT 102.000 130.200 102.600 133.600 ;
        RECT 106.000 133.400 106.800 133.600 ;
        RECT 108.800 130.200 109.400 135.000 ;
        RECT 124.400 135.000 125.200 135.800 ;
        RECT 130.600 135.600 131.400 135.800 ;
        RECT 125.800 135.000 131.400 135.600 ;
        RECT 110.000 133.600 110.800 134.400 ;
        RECT 118.000 133.600 118.800 134.400 ;
        RECT 122.800 133.600 123.600 134.400 ;
        RECT 124.400 134.200 125.000 135.000 ;
        RECT 125.800 134.800 126.600 135.000 ;
        RECT 129.200 134.800 130.000 135.000 ;
        RECT 124.400 133.600 130.000 134.200 ;
        RECT 116.400 131.600 117.200 132.400 ;
        RECT 102.000 129.400 102.800 130.200 ;
        RECT 108.600 129.400 109.400 130.200 ;
        RECT 116.500 128.400 117.100 131.600 ;
        RECT 118.000 129.600 118.800 130.400 ;
        RECT 124.400 130.200 125.000 133.600 ;
        RECT 127.600 131.600 128.400 132.400 ;
        RECT 129.400 132.200 130.000 133.600 ;
        RECT 129.400 131.400 130.200 132.200 ;
        RECT 130.800 130.200 131.400 135.000 ;
        RECT 132.400 133.600 133.200 134.400 ;
        RECT 132.500 130.400 133.100 133.600 ;
        RECT 137.200 131.600 138.000 132.400 ;
        RECT 124.400 129.400 125.200 130.200 ;
        RECT 130.600 129.400 131.400 130.200 ;
        RECT 132.400 129.600 133.200 130.400 ;
        RECT 116.400 127.600 117.200 128.400 ;
        RECT 129.200 127.600 130.000 128.400 ;
        RECT 103.600 123.600 104.400 124.400 ;
        RECT 100.400 117.600 101.200 118.400 ;
        RECT 103.700 110.400 104.300 123.600 ;
        RECT 90.800 109.600 91.600 110.400 ;
        RECT 103.600 109.600 104.400 110.400 ;
        RECT 89.200 107.600 90.000 108.400 ;
        RECT 89.300 98.400 89.900 107.600 ;
        RECT 94.000 105.600 94.800 106.400 ;
        RECT 54.000 95.600 54.800 96.400 ;
        RECT 33.200 71.600 34.000 72.400 ;
        RECT 36.200 71.800 37.000 72.600 ;
        RECT 38.100 72.400 38.700 83.600 ;
        RECT 33.300 52.400 33.900 71.600 ;
        RECT 34.800 67.600 35.600 68.400 ;
        RECT 33.200 51.600 34.000 52.400 ;
        RECT 31.600 50.300 32.400 50.400 ;
        RECT 31.600 49.700 33.900 50.300 ;
        RECT 31.600 49.600 32.400 49.700 ;
        RECT 31.600 47.600 32.400 48.400 ;
        RECT 31.700 38.400 32.300 47.600 ;
        RECT 31.600 37.600 32.400 38.400 ;
        RECT 30.000 29.600 30.800 30.400 ;
        RECT 30.000 27.600 30.800 28.400 ;
        RECT 20.400 26.200 21.200 27.000 ;
        RECT 21.800 26.400 26.000 27.000 ;
        RECT 27.000 26.200 27.800 27.000 ;
        RECT 25.200 23.600 26.000 24.400 ;
        RECT 23.600 21.600 24.400 22.400 ;
        RECT 7.600 17.600 8.400 18.400 ;
        RECT 17.200 4.200 18.000 17.800 ;
        RECT 18.800 4.200 19.600 17.800 ;
        RECT 20.400 4.200 21.200 17.800 ;
        RECT 22.000 6.200 22.800 17.800 ;
        RECT 23.700 16.400 24.300 21.600 ;
        RECT 25.300 20.300 25.900 23.600 ;
        RECT 25.300 19.700 27.500 20.300 ;
        RECT 23.600 15.600 24.400 16.400 ;
        RECT 25.200 6.200 26.000 17.800 ;
        RECT 26.900 14.400 27.500 19.700 ;
        RECT 26.800 13.600 27.600 14.400 ;
        RECT 28.400 6.200 29.200 17.800 ;
        RECT 30.000 4.200 30.800 17.800 ;
        RECT 31.600 4.200 32.400 17.800 ;
        RECT 33.300 12.400 33.900 49.700 ;
        RECT 34.900 42.400 35.500 67.600 ;
        RECT 36.200 67.000 36.800 71.800 ;
        RECT 38.000 71.600 38.800 72.400 ;
        RECT 42.800 71.800 43.600 72.600 ;
        RECT 38.800 68.400 39.600 68.600 ;
        RECT 43.000 68.400 43.600 71.800 ;
        RECT 50.800 69.600 51.600 70.400 ;
        RECT 50.900 68.400 51.500 69.600 ;
        RECT 38.800 67.800 43.600 68.400 ;
        RECT 38.000 67.000 38.800 67.200 ;
        RECT 41.400 67.000 42.200 67.200 ;
        RECT 43.000 67.000 43.600 67.800 ;
        RECT 50.800 67.600 51.600 68.400 ;
        RECT 36.200 66.200 37.000 67.000 ;
        RECT 38.000 66.400 42.200 67.000 ;
        RECT 42.800 66.200 43.600 67.000 ;
        RECT 54.100 66.400 54.700 95.600 ;
        RECT 55.600 86.200 56.400 97.800 ;
        RECT 57.200 93.600 58.000 94.400 ;
        RECT 58.800 86.200 59.600 97.800 ;
        RECT 60.400 84.200 61.200 97.800 ;
        RECT 62.000 84.200 62.800 97.800 ;
        RECT 89.200 97.600 90.000 98.400 ;
        RECT 94.100 96.400 94.700 105.600 ;
        RECT 105.200 104.200 106.000 117.800 ;
        RECT 106.800 104.200 107.600 117.800 ;
        RECT 108.400 104.200 109.200 117.800 ;
        RECT 110.000 104.200 110.800 115.800 ;
        RECT 111.600 105.600 112.400 106.400 ;
        RECT 111.700 96.400 112.300 105.600 ;
        RECT 113.200 104.200 114.000 115.800 ;
        RECT 114.800 107.600 115.600 108.400 ;
        RECT 116.400 104.200 117.200 115.800 ;
        RECT 118.000 104.200 118.800 117.800 ;
        RECT 119.600 104.200 120.400 117.800 ;
        RECT 129.300 110.400 129.900 127.600 ;
        RECT 137.300 110.400 137.900 131.600 ;
        RECT 142.000 124.200 142.800 137.800 ;
        RECT 143.600 124.200 144.400 137.800 ;
        RECT 145.200 126.200 146.000 137.800 ;
        RECT 146.800 133.600 147.600 134.400 ;
        RECT 146.900 132.400 147.500 133.600 ;
        RECT 146.800 131.600 147.600 132.400 ;
        RECT 148.400 126.200 149.200 137.800 ;
        RECT 150.100 136.400 150.700 139.600 ;
        RECT 150.000 135.600 150.800 136.400 ;
        RECT 151.600 126.200 152.400 137.800 ;
        RECT 153.200 124.200 154.000 137.800 ;
        RECT 154.800 124.200 155.600 137.800 ;
        RECT 156.400 124.200 157.200 137.800 ;
        RECT 166.000 133.600 167.000 134.400 ;
        RECT 167.600 131.600 168.400 132.400 ;
        RECT 167.700 128.400 168.300 131.600 ;
        RECT 167.600 127.600 168.400 128.400 ;
        RECT 167.700 118.400 168.300 127.600 ;
        RECT 169.300 120.400 169.900 151.600 ;
        RECT 170.900 148.400 171.500 163.600 ;
        RECT 172.400 159.600 173.200 160.400 ;
        RECT 172.500 148.400 173.100 159.600 ;
        RECT 177.300 150.400 177.900 171.600 ;
        RECT 180.500 160.400 181.100 183.600 ;
        RECT 185.300 172.400 185.900 189.600 ;
        RECT 190.000 184.200 190.800 197.800 ;
        RECT 191.600 184.200 192.400 197.800 ;
        RECT 193.200 184.200 194.000 195.800 ;
        RECT 194.800 187.600 195.600 188.400 ;
        RECT 194.900 178.400 195.500 187.600 ;
        RECT 196.400 184.200 197.200 195.800 ;
        RECT 198.000 185.600 198.800 186.400 ;
        RECT 198.100 184.400 198.700 185.600 ;
        RECT 198.000 183.600 198.800 184.400 ;
        RECT 199.600 184.200 200.400 195.800 ;
        RECT 201.200 184.200 202.000 197.800 ;
        RECT 202.800 184.200 203.600 197.800 ;
        RECT 204.400 184.200 205.200 197.800 ;
        RECT 214.000 183.600 214.800 184.400 ;
        RECT 202.800 181.600 203.600 182.400 ;
        RECT 202.900 178.400 203.500 181.600 ;
        RECT 194.800 177.600 195.600 178.400 ;
        RECT 202.800 177.600 203.600 178.400 ;
        RECT 190.000 175.600 190.800 176.400 ;
        RECT 193.400 175.600 194.200 175.800 ;
        RECT 193.400 175.000 199.000 175.600 ;
        RECT 199.600 175.000 200.400 175.800 ;
        RECT 207.600 175.600 208.400 176.400 ;
        RECT 186.800 173.600 187.600 174.400 ;
        RECT 191.600 173.600 192.400 174.400 ;
        RECT 185.200 171.600 186.000 172.400 ;
        RECT 182.000 169.600 182.800 170.400 ;
        RECT 193.400 170.200 194.000 175.000 ;
        RECT 194.800 174.800 195.600 175.000 ;
        RECT 198.200 174.800 199.000 175.000 ;
        RECT 199.800 174.200 200.400 175.000 ;
        RECT 207.700 174.400 208.300 175.600 ;
        RECT 194.800 173.600 200.400 174.200 ;
        RECT 201.200 173.600 202.000 174.400 ;
        RECT 207.600 173.600 208.400 174.400 ;
        RECT 194.800 172.200 195.400 173.600 ;
        RECT 194.600 171.400 195.400 172.200 ;
        RECT 199.800 170.200 200.400 173.600 ;
        RECT 201.300 172.400 201.900 173.600 ;
        RECT 214.100 172.400 214.700 183.600 ;
        RECT 201.200 171.600 202.000 172.400 ;
        RECT 206.000 171.600 206.800 172.400 ;
        RECT 214.000 171.600 214.800 172.400 ;
        RECT 193.400 169.400 194.200 170.200 ;
        RECT 199.600 169.400 200.400 170.200 ;
        RECT 180.400 159.600 181.200 160.400 ;
        RECT 177.200 149.600 178.000 150.400 ;
        RECT 170.800 147.600 171.600 148.400 ;
        RECT 172.400 147.600 173.200 148.400 ;
        RECT 170.800 143.600 171.600 144.400 ;
        RECT 170.900 136.400 171.500 143.600 ;
        RECT 170.800 135.600 171.600 136.400 ;
        RECT 172.500 132.400 173.100 147.600 ;
        RECT 182.000 144.200 182.800 157.800 ;
        RECT 183.600 144.200 184.400 157.800 ;
        RECT 185.200 144.200 186.000 155.800 ;
        RECT 186.800 147.600 187.600 148.400 ;
        RECT 188.400 144.200 189.200 155.800 ;
        RECT 190.000 145.600 190.800 146.400 ;
        RECT 191.600 144.200 192.400 155.800 ;
        RECT 193.200 144.200 194.000 157.800 ;
        RECT 194.800 144.200 195.600 157.800 ;
        RECT 196.400 144.200 197.200 157.800 ;
        RECT 214.000 149.600 214.800 150.400 ;
        RECT 199.600 147.600 200.400 148.400 ;
        RECT 199.700 138.400 200.300 147.600 ;
        RECT 206.000 143.600 206.800 144.400 ;
        RECT 188.400 137.600 189.200 138.400 ;
        RECT 199.600 137.600 200.400 138.400 ;
        RECT 188.500 136.400 189.100 137.600 ;
        RECT 175.600 135.000 176.400 135.800 ;
        RECT 177.000 135.000 181.200 135.600 ;
        RECT 182.200 135.000 183.000 135.800 ;
        RECT 183.600 135.600 184.400 136.400 ;
        RECT 188.400 135.600 189.200 136.400 ;
        RECT 193.200 135.600 194.000 136.400 ;
        RECT 196.400 135.600 197.200 136.400 ;
        RECT 175.600 134.200 176.200 135.000 ;
        RECT 177.000 134.800 177.800 135.000 ;
        RECT 180.400 134.800 181.200 135.000 ;
        RECT 175.600 133.600 180.400 134.200 ;
        RECT 172.400 131.600 173.200 132.400 ;
        RECT 175.600 130.200 176.200 133.600 ;
        RECT 179.600 133.400 180.400 133.600 ;
        RECT 182.400 130.200 183.000 135.000 ;
        RECT 183.700 134.400 184.300 135.600 ;
        RECT 196.500 134.400 197.100 135.600 ;
        RECT 197.800 135.000 198.600 135.800 ;
        RECT 199.600 135.000 203.800 135.600 ;
        RECT 204.400 135.000 205.200 135.800 ;
        RECT 183.600 133.600 184.400 134.400 ;
        RECT 196.400 133.600 197.200 134.400 ;
        RECT 193.200 131.600 194.000 132.400 ;
        RECT 175.600 129.400 176.400 130.200 ;
        RECT 182.200 129.400 183.000 130.200 ;
        RECT 185.200 129.600 186.000 130.400 ;
        RECT 194.800 129.600 195.600 130.400 ;
        RECT 197.800 130.200 198.400 135.000 ;
        RECT 199.600 134.800 200.400 135.000 ;
        RECT 203.000 134.800 203.800 135.000 ;
        RECT 204.600 134.200 205.200 135.000 ;
        RECT 206.100 134.400 206.700 143.600 ;
        RECT 207.600 137.600 208.400 138.400 ;
        RECT 214.100 134.400 214.700 149.600 ;
        RECT 200.400 133.600 205.200 134.200 ;
        RECT 206.000 134.300 206.800 134.400 ;
        RECT 206.000 133.700 208.300 134.300 ;
        RECT 206.000 133.600 206.800 133.700 ;
        RECT 200.400 133.400 201.200 133.600 ;
        RECT 204.600 130.200 205.200 133.600 ;
        RECT 207.700 130.400 208.300 133.700 ;
        RECT 210.800 133.600 211.600 134.400 ;
        RECT 214.000 133.600 214.800 134.400 ;
        RECT 210.900 132.400 211.500 133.600 ;
        RECT 210.800 131.600 211.600 132.400 ;
        RECT 185.300 128.400 185.900 129.600 ;
        RECT 194.900 128.400 195.500 129.600 ;
        RECT 197.800 129.400 198.600 130.200 ;
        RECT 204.400 129.400 205.200 130.200 ;
        RECT 207.600 129.600 208.400 130.400 ;
        RECT 210.900 128.400 211.500 131.600 ;
        RECT 185.200 127.600 186.000 128.400 ;
        RECT 191.600 127.600 192.400 128.400 ;
        RECT 194.800 127.600 195.600 128.400 ;
        RECT 210.800 127.600 211.600 128.400 ;
        RECT 177.200 123.600 178.000 124.400 ;
        RECT 169.200 119.600 170.000 120.400 ;
        RECT 124.400 109.600 125.200 110.400 ;
        RECT 129.200 109.600 130.000 110.400 ;
        RECT 134.000 109.600 134.800 110.400 ;
        RECT 137.200 109.600 138.000 110.400 ;
        RECT 138.800 109.600 139.600 110.400 ;
        RECT 124.500 108.400 125.100 109.600 ;
        RECT 134.100 108.400 134.700 109.600 ;
        RECT 124.400 107.600 125.200 108.400 ;
        RECT 134.000 107.600 134.800 108.400 ;
        RECT 84.200 95.000 85.000 95.800 ;
        RECT 86.000 95.000 90.200 95.600 ;
        RECT 90.800 95.000 91.600 95.800 ;
        RECT 94.000 95.600 94.800 96.400 ;
        RECT 100.400 95.600 101.200 96.400 ;
        RECT 111.600 95.600 112.400 96.400 ;
        RECT 82.800 93.600 83.600 94.400 ;
        RECT 82.900 92.400 83.500 93.600 ;
        RECT 81.200 91.600 82.000 92.400 ;
        RECT 82.800 91.600 83.600 92.400 ;
        RECT 66.800 89.600 67.600 90.400 ;
        RECT 78.000 89.600 78.800 90.400 ;
        RECT 78.100 84.400 78.700 89.600 ;
        RECT 81.300 84.400 81.900 91.600 ;
        RECT 78.000 83.600 78.800 84.400 ;
        RECT 81.200 83.600 82.000 84.400 ;
        RECT 54.000 65.600 54.800 66.400 ;
        RECT 52.400 63.600 53.200 64.400 ;
        RECT 62.000 64.200 62.800 77.800 ;
        RECT 63.600 64.200 64.400 77.800 ;
        RECT 65.200 64.200 66.000 77.800 ;
        RECT 66.800 64.200 67.600 75.800 ;
        RECT 68.400 65.600 69.200 66.400 ;
        RECT 70.000 64.200 70.800 75.800 ;
        RECT 71.600 67.600 72.400 68.400 ;
        RECT 73.200 64.200 74.000 75.800 ;
        RECT 74.800 64.200 75.600 77.800 ;
        RECT 76.400 64.200 77.200 77.800 ;
        RECT 78.100 72.000 78.700 83.600 ;
        RECT 78.000 71.200 78.800 72.000 ;
        RECT 52.500 56.400 53.100 63.600 ;
        RECT 82.900 58.400 83.500 91.600 ;
        RECT 84.200 90.200 84.800 95.000 ;
        RECT 86.000 94.800 86.800 95.000 ;
        RECT 89.400 94.800 90.200 95.000 ;
        RECT 91.000 94.200 91.600 95.000 ;
        RECT 94.100 94.400 94.700 95.600 ;
        RECT 86.800 93.600 91.600 94.200 ;
        RECT 94.000 93.600 94.800 94.400 ;
        RECT 100.400 93.600 101.200 94.400 ;
        RECT 103.600 93.600 104.400 94.400 ;
        RECT 108.400 93.600 109.200 94.400 ;
        RECT 86.800 93.400 87.600 93.600 ;
        RECT 91.000 90.200 91.600 93.600 ;
        RECT 95.600 91.600 96.400 92.400 ;
        RECT 84.200 89.400 85.000 90.200 ;
        RECT 90.800 89.400 91.600 90.200 ;
        RECT 100.400 89.600 101.200 90.400 ;
        RECT 108.400 89.600 109.200 90.400 ;
        RECT 110.000 89.600 110.800 90.400 ;
        RECT 103.600 87.600 104.400 88.400 ;
        RECT 92.400 73.600 93.200 74.400 ;
        RECT 89.200 67.600 90.000 68.400 ;
        RECT 89.300 66.400 89.900 67.600 ;
        RECT 87.600 65.600 88.400 66.400 ;
        RECT 89.200 65.600 90.000 66.400 ;
        RECT 86.000 63.600 86.800 64.400 ;
        RECT 82.800 57.600 83.600 58.400 ;
        RECT 41.200 55.600 42.000 56.400 ;
        RECT 52.400 55.600 53.200 56.400 ;
        RECT 55.600 55.600 56.400 56.400 ;
        RECT 73.200 55.600 74.000 56.400 ;
        RECT 55.700 54.400 56.300 55.600 ;
        RECT 36.400 53.600 37.200 54.400 ;
        RECT 39.600 53.600 40.400 54.400 ;
        RECT 50.800 53.600 51.600 54.400 ;
        RECT 55.600 53.600 56.400 54.400 ;
        RECT 65.200 53.600 66.000 54.400 ;
        RECT 39.700 52.400 40.300 53.600 ;
        RECT 39.600 51.600 40.400 52.400 ;
        RECT 46.000 51.600 46.800 52.400 ;
        RECT 36.400 49.600 37.200 50.400 ;
        RECT 36.500 48.400 37.100 49.600 ;
        RECT 36.400 47.600 37.200 48.400 ;
        RECT 39.700 42.400 40.300 51.600 ;
        RECT 34.800 41.600 35.600 42.400 ;
        RECT 39.600 41.600 40.400 42.400 ;
        RECT 46.100 40.400 46.700 51.600 ;
        RECT 50.900 48.400 51.500 53.600 ;
        RECT 52.400 51.600 53.200 52.400 ;
        RECT 54.000 51.600 54.800 52.400 ;
        RECT 47.600 47.600 48.400 48.400 ;
        RECT 50.800 47.600 51.600 48.400 ;
        RECT 46.000 39.600 46.800 40.400 ;
        RECT 46.000 38.300 46.800 38.400 ;
        RECT 47.700 38.300 48.300 47.600 ;
        RECT 49.200 43.600 50.000 44.400 ;
        RECT 49.300 42.400 49.900 43.600 ;
        RECT 49.200 41.600 50.000 42.400 ;
        RECT 49.200 39.600 50.000 40.400 ;
        RECT 49.300 38.400 49.900 39.600 ;
        RECT 46.000 37.700 48.300 38.300 ;
        RECT 46.000 37.600 46.800 37.700 ;
        RECT 49.200 37.600 50.000 38.400 ;
        RECT 34.800 31.600 35.600 32.400 ;
        RECT 41.200 29.600 42.000 30.400 ;
        RECT 38.000 27.600 38.800 28.400 ;
        RECT 38.100 26.400 38.700 27.600 ;
        RECT 50.900 26.400 51.500 47.600 ;
        RECT 52.500 28.400 53.100 51.600 ;
        RECT 55.600 49.600 56.400 50.400 ;
        RECT 55.700 42.400 56.300 49.600 ;
        RECT 71.600 47.600 72.400 48.400 ;
        RECT 55.600 41.600 56.400 42.400 ;
        RECT 55.700 32.400 56.300 41.600 ;
        RECT 55.600 31.600 56.400 32.400 ;
        RECT 63.400 31.800 64.200 32.600 ;
        RECT 70.000 31.800 70.800 32.600 ;
        RECT 55.700 28.400 56.300 31.600 ;
        RECT 52.400 27.600 53.200 28.400 ;
        RECT 55.600 27.600 56.400 28.400 ;
        RECT 63.400 27.000 64.000 31.800 ;
        RECT 66.000 28.400 66.800 28.600 ;
        RECT 70.200 28.400 70.800 31.800 ;
        RECT 71.600 29.600 72.400 30.400 ;
        RECT 66.000 27.800 70.800 28.400 ;
        RECT 65.200 27.000 66.000 27.200 ;
        RECT 68.600 27.000 69.400 27.200 ;
        RECT 70.200 27.000 70.800 27.800 ;
        RECT 71.600 28.300 72.400 28.400 ;
        RECT 73.300 28.300 73.900 55.600 ;
        RECT 82.900 54.400 83.500 57.600 ;
        RECT 82.800 53.600 83.600 54.400 ;
        RECT 86.100 52.400 86.700 63.600 ;
        RECT 87.700 52.400 88.300 65.600 ;
        RECT 92.500 58.400 93.100 73.600 ;
        RECT 103.700 72.400 104.300 87.600 ;
        RECT 108.500 78.400 109.100 89.600 ;
        RECT 111.700 82.400 112.300 95.600 ;
        RECT 113.200 89.600 114.000 90.400 ;
        RECT 111.600 81.600 112.400 82.400 ;
        RECT 108.400 77.600 109.200 78.400 ;
        RECT 105.200 73.600 106.000 74.400 ;
        RECT 103.600 71.600 104.400 72.400 ;
        RECT 105.200 69.600 106.000 70.400 ;
        RECT 110.000 69.600 110.800 70.400 ;
        RECT 113.300 66.400 113.900 89.600 ;
        RECT 119.600 84.200 120.400 97.800 ;
        RECT 121.200 84.200 122.000 97.800 ;
        RECT 122.800 84.200 123.600 97.800 ;
        RECT 124.400 86.200 125.200 97.800 ;
        RECT 126.000 95.600 126.800 96.400 ;
        RECT 127.600 86.200 128.400 97.800 ;
        RECT 129.200 93.600 130.000 94.400 ;
        RECT 130.800 86.200 131.600 97.800 ;
        RECT 127.600 83.600 128.400 84.400 ;
        RECT 132.400 84.200 133.200 97.800 ;
        RECT 134.000 84.200 134.800 97.800 ;
        RECT 138.900 92.400 139.500 109.600 ;
        RECT 143.600 104.200 144.400 117.800 ;
        RECT 145.200 104.200 146.000 117.800 ;
        RECT 146.800 104.200 147.600 115.800 ;
        RECT 148.400 107.600 149.200 108.400 ;
        RECT 150.000 104.200 150.800 115.800 ;
        RECT 151.600 105.600 152.400 106.400 ;
        RECT 151.700 102.400 152.300 105.600 ;
        RECT 153.200 104.200 154.000 115.800 ;
        RECT 154.800 104.200 155.600 117.800 ;
        RECT 156.400 104.200 157.200 117.800 ;
        RECT 158.000 104.200 158.800 117.800 ;
        RECT 167.600 117.600 168.400 118.400 ;
        RECT 159.600 109.600 160.400 110.400 ;
        RECT 177.300 108.400 177.900 123.600 ;
        RECT 191.700 120.400 192.300 127.600 ;
        RECT 191.600 119.600 192.400 120.400 ;
        RECT 178.800 109.600 179.600 110.400 ;
        RECT 177.200 107.600 178.000 108.400 ;
        RECT 164.400 103.600 165.200 104.400 ;
        RECT 183.600 104.200 184.400 117.800 ;
        RECT 185.200 104.200 186.000 117.800 ;
        RECT 186.800 104.200 187.600 115.800 ;
        RECT 188.400 107.600 189.200 108.400 ;
        RECT 145.200 101.600 146.000 102.400 ;
        RECT 151.600 101.600 152.400 102.400 ;
        RECT 138.800 91.600 139.600 92.400 ;
        RECT 114.800 81.600 115.600 82.400 ;
        RECT 114.900 78.400 115.500 81.600 ;
        RECT 114.800 77.600 115.600 78.400 ;
        RECT 127.700 70.400 128.300 83.600 ;
        RECT 140.400 81.600 141.200 82.400 ;
        RECT 127.600 69.600 128.400 70.400 ;
        RECT 110.000 66.300 110.800 66.400 ;
        RECT 108.500 65.700 110.800 66.300 ;
        RECT 92.400 57.600 93.200 58.400 ;
        RECT 108.500 56.400 109.100 65.700 ;
        RECT 110.000 65.600 110.800 65.700 ;
        RECT 113.200 65.600 114.000 66.400 ;
        RECT 92.400 55.600 93.200 56.400 ;
        RECT 105.200 55.600 106.000 56.400 ;
        RECT 108.400 55.600 109.200 56.400 ;
        RECT 111.600 55.600 112.400 56.400 ;
        RECT 92.400 53.600 93.200 54.400 ;
        RECT 103.600 53.600 104.400 54.400 ;
        RECT 92.500 52.400 93.100 53.600 ;
        RECT 79.600 51.600 80.400 52.400 ;
        RECT 86.000 51.600 86.800 52.400 ;
        RECT 87.600 51.600 88.400 52.400 ;
        RECT 90.800 51.600 91.600 52.400 ;
        RECT 92.400 51.600 93.200 52.400 ;
        RECT 102.000 51.600 102.800 52.400 ;
        RECT 103.600 51.600 104.400 52.400 ;
        RECT 90.900 50.400 91.500 51.600 ;
        RECT 102.100 50.400 102.700 51.600 ;
        RECT 103.700 50.400 104.300 51.600 ;
        RECT 90.800 49.600 91.600 50.400 ;
        RECT 102.000 49.600 102.800 50.400 ;
        RECT 103.600 49.600 104.400 50.400 ;
        RECT 81.200 47.600 82.000 48.400 ;
        RECT 103.600 47.600 104.400 48.400 ;
        RECT 78.000 29.600 78.800 30.400 ;
        RECT 71.600 27.700 73.900 28.300 ;
        RECT 71.600 27.600 72.400 27.700 ;
        RECT 38.000 25.600 38.800 26.400 ;
        RECT 50.800 25.600 51.600 26.400 ;
        RECT 63.400 26.200 64.200 27.000 ;
        RECT 65.200 26.400 69.400 27.000 ;
        RECT 70.000 26.200 70.800 27.000 ;
        RECT 50.900 16.400 51.500 25.600 ;
        RECT 60.400 23.600 61.200 24.400 ;
        RECT 50.800 15.600 51.600 16.400 ;
        RECT 60.500 14.400 61.100 23.600 ;
        RECT 68.400 21.600 69.200 22.400 ;
        RECT 60.400 13.600 61.200 14.400 ;
        RECT 33.200 11.600 34.000 12.400 ;
        RECT 60.400 11.600 61.200 12.400 ;
        RECT 62.000 4.200 62.800 17.800 ;
        RECT 63.600 4.200 64.400 17.800 ;
        RECT 65.200 4.200 66.000 17.800 ;
        RECT 66.800 6.200 67.600 17.800 ;
        RECT 68.500 16.400 69.100 21.600 ;
        RECT 73.300 20.400 73.900 27.700 ;
        RECT 73.200 19.600 74.000 20.400 ;
        RECT 68.400 15.600 69.200 16.400 ;
        RECT 70.000 6.200 70.800 17.800 ;
        RECT 71.600 13.600 72.400 14.400 ;
        RECT 73.200 6.200 74.000 17.800 ;
        RECT 74.800 4.200 75.600 17.800 ;
        RECT 76.400 4.200 77.200 17.800 ;
        RECT 78.100 12.400 78.700 29.600 ;
        RECT 81.200 24.200 82.000 37.800 ;
        RECT 82.800 24.200 83.600 37.800 ;
        RECT 84.400 24.200 85.200 35.800 ;
        RECT 86.000 29.600 86.800 30.400 ;
        RECT 86.100 28.400 86.700 29.600 ;
        RECT 86.000 27.600 86.800 28.400 ;
        RECT 87.600 24.200 88.400 35.800 ;
        RECT 89.200 25.600 90.000 26.400 ;
        RECT 90.800 24.200 91.600 35.800 ;
        RECT 92.400 24.200 93.200 37.800 ;
        RECT 94.000 24.200 94.800 37.800 ;
        RECT 95.600 24.200 96.400 37.800 ;
        RECT 103.700 28.400 104.300 47.600 ;
        RECT 105.300 38.400 105.900 55.600 ;
        RECT 106.800 49.600 107.600 50.400 ;
        RECT 105.200 37.600 106.000 38.400 ;
        RECT 103.600 27.600 104.400 28.400 ;
        RECT 89.200 19.600 90.000 20.400 ;
        RECT 89.300 12.400 89.900 19.600 ;
        RECT 100.400 17.600 101.200 18.400 ;
        RECT 106.800 17.600 107.600 18.400 ;
        RECT 90.800 13.600 91.600 14.400 ;
        RECT 90.900 12.400 91.500 13.600 ;
        RECT 100.500 12.400 101.100 17.600 ;
        RECT 108.500 12.400 109.100 55.600 ;
        RECT 113.300 54.400 113.900 65.600 ;
        RECT 130.800 63.600 131.600 64.400 ;
        RECT 119.600 55.600 120.400 56.400 ;
        RECT 113.200 53.600 114.000 54.400 ;
        RECT 130.900 52.400 131.500 63.600 ;
        RECT 110.000 51.600 110.800 52.400 ;
        RECT 111.600 51.600 112.400 52.400 ;
        RECT 114.800 51.600 115.600 52.400 ;
        RECT 119.600 51.600 120.400 52.400 ;
        RECT 122.800 51.600 123.600 52.400 ;
        RECT 130.800 51.600 131.600 52.400 ;
        RECT 110.100 38.400 110.700 51.600 ;
        RECT 110.000 37.600 110.800 38.400 ;
        RECT 110.000 23.600 110.800 24.400 ;
        RECT 110.100 14.400 110.700 23.600 ;
        RECT 111.700 18.400 112.300 51.600 ;
        RECT 119.700 40.400 120.300 51.600 ;
        RECT 122.800 43.600 123.600 44.400 ;
        RECT 122.900 42.400 123.500 43.600 ;
        RECT 122.800 41.600 123.600 42.400 ;
        RECT 119.600 39.600 120.400 40.400 ;
        RECT 130.900 38.400 131.500 51.600 ;
        RECT 132.400 44.200 133.200 57.800 ;
        RECT 134.000 44.200 134.800 57.800 ;
        RECT 135.600 46.200 136.400 57.800 ;
        RECT 137.200 53.600 138.000 54.400 ;
        RECT 138.800 46.200 139.600 57.800 ;
        RECT 140.500 56.400 141.100 81.600 ;
        RECT 145.300 78.400 145.900 101.600 ;
        RECT 151.700 96.400 152.300 101.600 ;
        RECT 151.600 95.600 152.400 96.400 ;
        RECT 151.600 91.600 152.400 92.400 ;
        RECT 156.400 84.200 157.200 97.800 ;
        RECT 158.000 84.200 158.800 97.800 ;
        RECT 159.600 86.200 160.400 97.800 ;
        RECT 161.200 93.600 162.000 94.400 ;
        RECT 162.800 86.200 163.600 97.800 ;
        RECT 164.500 96.400 165.100 103.600 ;
        RECT 188.500 102.400 189.100 107.600 ;
        RECT 190.000 104.200 190.800 115.800 ;
        RECT 191.600 105.600 192.400 106.400 ;
        RECT 191.700 104.400 192.300 105.600 ;
        RECT 191.600 103.600 192.400 104.400 ;
        RECT 193.200 104.200 194.000 115.800 ;
        RECT 194.800 104.200 195.600 117.800 ;
        RECT 196.400 104.200 197.200 117.800 ;
        RECT 198.000 104.200 198.800 117.800 ;
        RECT 202.800 103.600 203.600 104.400 ;
        RECT 207.600 103.600 208.400 104.400 ;
        RECT 188.400 101.600 189.200 102.400 ;
        RECT 164.400 95.600 165.200 96.400 ;
        RECT 166.000 86.200 166.800 97.800 ;
        RECT 167.600 84.200 168.400 97.800 ;
        RECT 169.200 84.200 170.000 97.800 ;
        RECT 170.800 84.200 171.600 97.800 ;
        RECT 185.200 95.000 186.000 95.800 ;
        RECT 186.600 95.000 190.800 95.600 ;
        RECT 191.800 95.000 192.600 95.800 ;
        RECT 182.000 93.600 182.800 94.400 ;
        RECT 183.600 93.600 184.400 94.400 ;
        RECT 185.200 94.200 185.800 95.000 ;
        RECT 186.600 94.800 187.400 95.000 ;
        RECT 190.000 94.800 190.800 95.000 ;
        RECT 185.200 93.600 190.000 94.200 ;
        RECT 182.100 92.400 182.700 93.600 ;
        RECT 183.700 92.400 184.300 93.600 ;
        RECT 182.000 91.600 182.800 92.400 ;
        RECT 183.600 91.600 184.400 92.400 ;
        RECT 185.200 90.200 185.800 93.600 ;
        RECT 189.200 93.400 190.000 93.600 ;
        RECT 192.000 90.200 192.600 95.000 ;
        RECT 202.900 94.400 203.500 103.600 ;
        RECT 207.600 101.600 208.400 102.400 ;
        RECT 207.700 98.400 208.300 101.600 ;
        RECT 207.600 97.600 208.400 98.400 ;
        RECT 206.200 95.600 207.000 95.800 ;
        RECT 206.200 95.000 211.800 95.600 ;
        RECT 212.400 95.000 213.200 95.800 ;
        RECT 198.000 93.600 198.800 94.400 ;
        RECT 202.800 93.600 203.600 94.400 ;
        RECT 204.400 93.600 205.200 94.400 ;
        RECT 199.600 91.600 200.400 92.400 ;
        RECT 199.700 90.400 200.300 91.600 ;
        RECT 204.500 90.400 205.100 93.600 ;
        RECT 185.200 89.400 186.000 90.200 ;
        RECT 191.800 89.400 192.600 90.200 ;
        RECT 194.800 89.600 195.600 90.400 ;
        RECT 199.600 89.600 200.400 90.400 ;
        RECT 204.400 89.600 205.200 90.400 ;
        RECT 206.200 90.200 206.800 95.000 ;
        RECT 207.600 94.800 208.400 95.000 ;
        RECT 211.000 94.800 211.800 95.000 ;
        RECT 212.600 94.200 213.200 95.000 ;
        RECT 207.600 93.600 213.200 94.200 ;
        RECT 214.000 93.600 214.800 94.400 ;
        RECT 207.600 92.200 208.200 93.600 ;
        RECT 207.400 91.400 208.200 92.200 ;
        RECT 212.600 90.200 213.200 93.600 ;
        RECT 215.600 91.600 216.400 92.400 ;
        RECT 191.600 87.600 192.400 88.400 ;
        RECT 191.700 78.400 192.300 87.600 ;
        RECT 201.200 83.600 202.000 84.400 ;
        RECT 145.200 77.600 146.000 78.400 ;
        RECT 191.600 77.600 192.400 78.400 ;
        RECT 175.800 71.800 176.600 72.600 ;
        RECT 182.000 71.800 182.800 72.600 ;
        RECT 151.600 69.600 152.400 70.400 ;
        RECT 158.000 69.600 158.800 70.400 ;
        RECT 162.800 69.600 163.600 70.400 ;
        RECT 164.400 69.600 165.200 70.400 ;
        RECT 167.600 69.600 168.400 70.400 ;
        RECT 169.200 69.600 170.000 70.400 ;
        RECT 151.700 68.400 152.300 69.600 ;
        RECT 162.900 68.400 163.500 69.600 ;
        RECT 151.600 67.600 152.400 68.400 ;
        RECT 162.800 67.600 163.600 68.400 ;
        RECT 148.400 65.600 149.200 66.400 ;
        RECT 151.600 65.600 152.400 66.400 ;
        RECT 161.200 65.600 162.000 66.400 ;
        RECT 150.000 63.600 150.800 64.400 ;
        RECT 140.400 55.600 141.200 56.400 ;
        RECT 119.600 24.200 120.400 37.800 ;
        RECT 121.200 24.200 122.000 37.800 ;
        RECT 122.800 24.200 123.600 37.800 ;
        RECT 130.800 37.600 131.600 38.400 ;
        RECT 124.400 24.200 125.200 35.800 ;
        RECT 126.000 25.600 126.800 26.400 ;
        RECT 111.600 17.600 112.400 18.400 ;
        RECT 110.000 13.600 110.800 14.400 ;
        RECT 78.000 11.600 78.800 12.400 ;
        RECT 89.200 11.600 90.000 12.400 ;
        RECT 90.800 11.600 91.600 12.400 ;
        RECT 95.600 11.600 96.400 12.400 ;
        RECT 100.400 11.600 101.200 12.400 ;
        RECT 108.400 11.600 109.200 12.400 ;
        RECT 116.400 4.200 117.200 17.800 ;
        RECT 118.000 4.200 118.800 17.800 ;
        RECT 119.600 4.200 120.400 17.800 ;
        RECT 121.200 6.200 122.000 17.800 ;
        RECT 122.800 15.600 123.600 16.400 ;
        RECT 124.400 6.200 125.200 17.800 ;
        RECT 126.100 16.400 126.700 25.600 ;
        RECT 127.600 24.200 128.400 35.800 ;
        RECT 129.200 27.600 130.000 28.400 ;
        RECT 130.800 24.200 131.600 35.800 ;
        RECT 132.400 24.200 133.200 37.800 ;
        RECT 134.000 24.200 134.800 37.800 ;
        RECT 135.600 37.600 136.400 38.400 ;
        RECT 135.700 32.000 136.300 37.600 ;
        RECT 135.600 31.200 136.400 32.000 ;
        RECT 138.800 31.600 139.600 32.400 ;
        RECT 126.000 15.600 126.800 16.400 ;
        RECT 126.000 13.600 126.800 14.400 ;
        RECT 127.600 6.200 128.400 17.800 ;
        RECT 129.200 4.200 130.000 17.800 ;
        RECT 130.800 4.200 131.600 17.800 ;
        RECT 138.900 12.400 139.500 31.600 ;
        RECT 140.500 26.400 141.100 55.600 ;
        RECT 142.000 46.200 142.800 57.800 ;
        RECT 143.600 44.200 144.400 57.800 ;
        RECT 145.200 44.200 146.000 57.800 ;
        RECT 146.800 44.200 147.600 57.800 ;
        RECT 150.100 54.400 150.700 63.600 ;
        RECT 162.900 58.400 163.500 67.600 ;
        RECT 164.500 66.400 165.100 69.600 ;
        RECT 167.700 68.400 168.300 69.600 ;
        RECT 167.600 67.600 168.400 68.400 ;
        RECT 174.000 67.600 174.800 68.400 ;
        RECT 175.800 67.000 176.400 71.800 ;
        RECT 177.000 69.800 177.800 70.600 ;
        RECT 177.200 68.400 177.800 69.800 ;
        RECT 182.200 68.400 182.800 71.800 ;
        RECT 194.800 71.600 195.600 72.400 ;
        RECT 199.600 71.600 200.400 72.400 ;
        RECT 194.900 70.400 195.500 71.600 ;
        RECT 201.300 70.400 201.900 83.600 ;
        RECT 204.500 78.400 205.100 89.600 ;
        RECT 206.200 89.400 207.000 90.200 ;
        RECT 212.400 89.400 213.200 90.200 ;
        RECT 204.400 77.600 205.200 78.400 ;
        RECT 183.600 69.600 184.400 70.400 ;
        RECT 186.800 69.600 187.600 70.400 ;
        RECT 190.000 69.600 190.800 70.400 ;
        RECT 194.800 69.600 195.600 70.400 ;
        RECT 198.000 69.600 198.800 70.400 ;
        RECT 201.200 69.600 202.000 70.400 ;
        RECT 210.800 69.600 211.600 70.400 ;
        RECT 183.700 68.400 184.300 69.600 ;
        RECT 177.200 67.800 182.800 68.400 ;
        RECT 177.200 67.000 178.000 67.200 ;
        RECT 180.600 67.000 181.400 67.200 ;
        RECT 182.200 67.000 182.800 67.800 ;
        RECT 183.600 67.600 184.400 68.400 ;
        RECT 185.200 67.600 186.000 68.400 ;
        RECT 175.800 66.400 181.400 67.000 ;
        RECT 164.400 65.600 165.200 66.400 ;
        RECT 175.800 66.200 176.600 66.400 ;
        RECT 182.000 66.200 182.800 67.000 ;
        RECT 186.900 66.400 187.500 69.600 ;
        RECT 190.100 68.400 190.700 69.600 ;
        RECT 190.000 67.600 190.800 68.400 ;
        RECT 196.400 67.600 197.200 68.400 ;
        RECT 209.200 67.600 210.000 68.400 ;
        RECT 209.300 66.400 209.900 67.600 ;
        RECT 210.900 66.400 211.500 69.600 ;
        RECT 186.800 65.600 187.600 66.400 ;
        RECT 198.000 65.600 198.800 66.400 ;
        RECT 202.800 65.600 203.600 66.400 ;
        RECT 209.200 65.600 210.000 66.400 ;
        RECT 210.800 65.600 211.600 66.400 ;
        RECT 159.600 57.600 160.400 58.400 ;
        RECT 162.800 57.600 163.600 58.400 ;
        RECT 150.000 53.600 150.800 54.400 ;
        RECT 148.400 51.600 149.200 52.400 ;
        RECT 146.800 39.600 147.600 40.400 ;
        RECT 146.900 32.400 147.500 39.600 ;
        RECT 159.700 38.400 160.300 57.600 ;
        RECT 162.800 56.300 163.600 56.400 ;
        RECT 164.500 56.300 165.100 65.600 ;
        RECT 177.200 63.600 178.000 64.400 ;
        RECT 162.800 55.700 165.100 56.300 ;
        RECT 162.800 55.600 163.600 55.700 ;
        RECT 167.600 51.600 168.400 52.400 ;
        RECT 170.800 51.600 171.600 52.400 ;
        RECT 159.600 37.600 160.400 38.400 ;
        RECT 146.800 31.600 147.600 32.400 ;
        RECT 170.900 30.400 171.500 51.600 ;
        RECT 172.400 44.200 173.200 57.800 ;
        RECT 174.000 44.200 174.800 57.800 ;
        RECT 175.600 46.200 176.400 57.800 ;
        RECT 177.200 53.600 178.000 54.400 ;
        RECT 178.800 46.200 179.600 57.800 ;
        RECT 180.400 55.600 181.200 56.400 ;
        RECT 170.800 29.600 171.600 30.400 ;
        RECT 143.600 27.600 144.400 28.400 ;
        RECT 156.400 27.600 157.200 28.400 ;
        RECT 143.700 26.400 144.300 27.600 ;
        RECT 156.500 26.400 157.100 27.600 ;
        RECT 140.400 25.600 141.200 26.400 ;
        RECT 143.600 25.600 144.400 26.400 ;
        RECT 151.600 25.600 152.400 26.400 ;
        RECT 156.400 25.600 157.200 26.400 ;
        RECT 158.000 25.600 158.800 26.400 ;
        RECT 164.400 25.600 165.200 26.400 ;
        RECT 143.700 16.400 144.300 25.600 ;
        RECT 158.100 24.400 158.700 25.600 ;
        RECT 146.800 23.600 147.600 24.400 ;
        RECT 158.000 23.600 158.800 24.400 ;
        RECT 162.800 23.600 163.600 24.400 ;
        RECT 162.900 18.400 163.500 23.600 ;
        RECT 170.900 20.400 171.500 29.600 ;
        RECT 174.000 24.200 174.800 37.800 ;
        RECT 175.600 24.200 176.400 37.800 ;
        RECT 178.800 37.600 179.600 38.400 ;
        RECT 180.500 38.300 181.100 55.600 ;
        RECT 182.000 46.200 182.800 57.800 ;
        RECT 183.600 44.200 184.400 57.800 ;
        RECT 185.200 44.200 186.000 57.800 ;
        RECT 186.800 44.200 187.600 57.800 ;
        RECT 196.400 47.600 197.200 48.400 ;
        RECT 198.100 38.400 198.700 65.600 ;
        RECT 199.600 63.600 200.400 64.400 ;
        RECT 199.700 52.400 200.300 63.600 ;
        RECT 202.900 62.300 203.500 65.600 ;
        RECT 204.400 63.600 205.200 64.400 ;
        RECT 202.900 61.700 205.100 62.300 ;
        RECT 204.500 58.400 205.100 61.700 ;
        RECT 204.400 57.600 205.200 58.400 ;
        RECT 202.800 55.600 203.600 56.400 ;
        RECT 201.200 53.600 202.000 54.400 ;
        RECT 209.300 52.400 209.900 65.600 ;
        RECT 212.400 55.600 213.200 56.400 ;
        RECT 214.000 55.600 214.800 56.400 ;
        RECT 210.800 53.600 211.600 54.400 ;
        RECT 199.600 51.600 200.400 52.400 ;
        RECT 209.200 51.600 210.000 52.400 ;
        RECT 204.400 47.600 205.200 48.400 ;
        RECT 180.500 37.700 182.700 38.300 ;
        RECT 177.200 24.200 178.000 35.800 ;
        RECT 178.900 28.400 179.500 37.600 ;
        RECT 178.800 27.600 179.600 28.400 ;
        RECT 180.400 24.200 181.200 35.800 ;
        RECT 182.100 26.400 182.700 37.700 ;
        RECT 182.000 25.600 182.800 26.400 ;
        RECT 170.800 19.600 171.600 20.400 ;
        RECT 174.000 19.600 174.800 20.400 ;
        RECT 143.600 15.600 144.400 16.400 ;
        RECT 135.600 11.600 136.400 12.400 ;
        RECT 138.800 11.600 139.600 12.400 ;
        RECT 156.400 4.200 157.200 17.800 ;
        RECT 158.000 4.200 158.800 17.800 ;
        RECT 159.600 4.200 160.400 17.800 ;
        RECT 161.200 6.200 162.000 17.800 ;
        RECT 162.800 17.600 163.600 18.400 ;
        RECT 162.800 15.600 163.600 16.400 ;
        RECT 164.400 6.200 165.200 17.800 ;
        RECT 166.000 17.600 166.800 18.400 ;
        RECT 166.100 14.400 166.700 17.600 ;
        RECT 166.000 13.600 166.800 14.400 ;
        RECT 167.600 6.200 168.400 17.800 ;
        RECT 169.200 4.200 170.000 17.800 ;
        RECT 170.800 4.200 171.600 17.800 ;
        RECT 174.100 12.400 174.700 19.600 ;
        RECT 182.100 16.400 182.700 25.600 ;
        RECT 183.600 24.200 184.400 35.800 ;
        RECT 185.200 24.200 186.000 37.800 ;
        RECT 186.800 24.200 187.600 37.800 ;
        RECT 188.400 24.200 189.200 37.800 ;
        RECT 198.000 37.600 198.800 38.400 ;
        RECT 209.300 36.400 209.900 51.600 ;
        RECT 201.200 35.600 202.000 36.400 ;
        RECT 209.200 35.600 210.000 36.400 ;
        RECT 201.300 28.400 201.900 35.600 ;
        RECT 203.000 31.800 203.800 32.600 ;
        RECT 209.200 31.800 210.000 32.600 ;
        RECT 201.200 27.600 202.000 28.400 ;
        RECT 203.000 27.000 203.600 31.800 ;
        RECT 204.200 29.800 205.000 30.600 ;
        RECT 204.400 28.400 205.000 29.800 ;
        RECT 209.400 28.400 210.000 31.800 ;
        RECT 210.900 30.400 211.500 53.600 ;
        RECT 214.100 48.400 214.700 55.600 ;
        RECT 215.600 51.600 216.400 52.400 ;
        RECT 215.700 48.400 216.300 51.600 ;
        RECT 214.000 47.600 214.800 48.400 ;
        RECT 215.600 47.600 216.400 48.400 ;
        RECT 210.800 29.600 211.600 30.400 ;
        RECT 212.400 29.600 213.200 30.400 ;
        RECT 204.400 27.800 210.000 28.400 ;
        RECT 204.400 27.000 205.200 27.200 ;
        RECT 207.800 27.000 208.600 27.200 ;
        RECT 209.400 27.000 210.000 27.800 ;
        RECT 203.000 26.400 208.600 27.000 ;
        RECT 203.000 26.200 203.800 26.400 ;
        RECT 209.200 26.200 210.000 27.000 ;
        RECT 204.400 23.600 205.200 24.400 ;
        RECT 183.600 19.600 184.400 20.400 ;
        RECT 182.000 15.600 182.800 16.400 ;
        RECT 183.700 12.400 184.300 19.600 ;
        RECT 174.000 11.600 174.800 12.400 ;
        RECT 183.600 11.600 184.400 12.400 ;
        RECT 188.400 4.200 189.200 17.800 ;
        RECT 190.000 4.200 190.800 17.800 ;
        RECT 191.600 6.200 192.400 17.800 ;
        RECT 193.200 13.600 194.000 14.400 ;
        RECT 194.800 6.200 195.600 17.800 ;
        RECT 196.400 15.600 197.200 16.400 ;
        RECT 198.000 6.200 198.800 17.800 ;
        RECT 199.600 4.200 200.400 17.800 ;
        RECT 201.200 4.200 202.000 17.800 ;
        RECT 202.800 4.200 203.600 17.800 ;
        RECT 204.500 14.400 205.100 23.600 ;
        RECT 212.500 18.400 213.100 29.600 ;
        RECT 212.400 17.600 213.200 18.400 ;
        RECT 204.400 13.600 205.200 14.400 ;
      LAYER via2 ;
        RECT 68.400 189.600 69.200 190.400 ;
        RECT 138.800 189.600 139.600 190.400 ;
        RECT 166.000 133.600 166.800 134.400 ;
      LAYER metal3 ;
        RECT 50.800 194.300 51.600 194.400 ;
        RECT 54.000 194.300 54.800 194.400 ;
        RECT 50.800 193.700 54.800 194.300 ;
        RECT 50.800 193.600 51.600 193.700 ;
        RECT 54.000 193.600 54.800 193.700 ;
        RECT 34.800 192.300 35.600 192.400 ;
        RECT 60.400 192.300 61.200 192.400 ;
        RECT 34.800 191.700 61.200 192.300 ;
        RECT 34.800 191.600 35.600 191.700 ;
        RECT 60.400 191.600 61.200 191.700 ;
        RECT 119.600 192.300 120.400 192.400 ;
        RECT 150.000 192.300 150.800 192.400 ;
        RECT 119.600 191.700 150.800 192.300 ;
        RECT 119.600 191.600 120.400 191.700 ;
        RECT 150.000 191.600 150.800 191.700 ;
        RECT 22.000 190.300 22.800 190.400 ;
        RECT 26.800 190.300 27.600 190.400 ;
        RECT 22.000 189.700 27.600 190.300 ;
        RECT 22.000 189.600 22.800 189.700 ;
        RECT 26.800 189.600 27.600 189.700 ;
        RECT 38.000 190.300 38.800 190.400 ;
        RECT 55.600 190.300 56.400 190.400 ;
        RECT 68.400 190.300 69.200 190.400 ;
        RECT 38.000 189.700 69.200 190.300 ;
        RECT 38.000 189.600 38.800 189.700 ;
        RECT 55.600 189.600 56.400 189.700 ;
        RECT 68.400 189.600 69.200 189.700 ;
        RECT 97.200 190.300 98.000 190.400 ;
        RECT 110.000 190.300 110.800 190.400 ;
        RECT 97.200 189.700 110.800 190.300 ;
        RECT 97.200 189.600 98.000 189.700 ;
        RECT 110.000 189.600 110.800 189.700 ;
        RECT 138.800 190.300 139.600 190.400 ;
        RECT 145.200 190.300 146.000 190.400 ;
        RECT 167.600 190.300 168.400 190.400 ;
        RECT 138.800 189.700 168.400 190.300 ;
        RECT 138.800 189.600 139.600 189.700 ;
        RECT 145.200 189.600 146.000 189.700 ;
        RECT 167.600 189.600 168.400 189.700 ;
        RECT 170.800 190.300 171.600 190.400 ;
        RECT 174.000 190.300 174.800 190.400 ;
        RECT 170.800 189.700 174.800 190.300 ;
        RECT 170.800 189.600 171.600 189.700 ;
        RECT 174.000 189.600 174.800 189.700 ;
        RECT 28.400 188.300 29.200 188.400 ;
        RECT 38.000 188.300 38.800 188.400 ;
        RECT 28.400 187.700 38.800 188.300 ;
        RECT 28.400 187.600 29.200 187.700 ;
        RECT 38.000 187.600 38.800 187.700 ;
        RECT 46.000 188.300 46.800 188.400 ;
        RECT 49.200 188.300 50.000 188.400 ;
        RECT 46.000 187.700 50.000 188.300 ;
        RECT 46.000 187.600 46.800 187.700 ;
        RECT 49.200 187.600 50.000 187.700 ;
        RECT 52.400 188.300 53.200 188.400 ;
        RECT 57.200 188.300 58.000 188.400 ;
        RECT 52.400 187.700 58.000 188.300 ;
        RECT 52.400 187.600 53.200 187.700 ;
        RECT 57.200 187.600 58.000 187.700 ;
        RECT 58.800 188.300 59.600 188.400 ;
        RECT 87.600 188.300 88.400 188.400 ;
        RECT 58.800 187.700 88.400 188.300 ;
        RECT 58.800 187.600 59.600 187.700 ;
        RECT 87.600 187.600 88.400 187.700 ;
        RECT 156.400 188.300 157.200 188.400 ;
        RECT 164.400 188.300 165.200 188.400 ;
        RECT 156.400 187.700 165.200 188.300 ;
        RECT 156.400 187.600 157.200 187.700 ;
        RECT 164.400 187.600 165.200 187.700 ;
        RECT 4.400 186.300 5.200 186.400 ;
        RECT 28.400 186.300 29.200 186.400 ;
        RECT 44.400 186.300 45.200 186.400 ;
        RECT 4.400 185.700 45.200 186.300 ;
        RECT 4.400 185.600 5.200 185.700 ;
        RECT 28.400 185.600 29.200 185.700 ;
        RECT 44.400 185.600 45.200 185.700 ;
        RECT 46.000 186.300 46.800 186.400 ;
        RECT 47.600 186.300 48.400 186.400 ;
        RECT 46.000 185.700 48.400 186.300 ;
        RECT 46.000 185.600 46.800 185.700 ;
        RECT 47.600 185.600 48.400 185.700 ;
        RECT 119.600 186.300 120.400 186.400 ;
        RECT 122.800 186.300 123.600 186.400 ;
        RECT 119.600 185.700 123.600 186.300 ;
        RECT 119.600 185.600 120.400 185.700 ;
        RECT 122.800 185.600 123.600 185.700 ;
        RECT 10.800 184.300 11.600 184.400 ;
        RECT 22.000 184.300 22.800 184.400 ;
        RECT 10.800 183.700 22.800 184.300 ;
        RECT 10.800 183.600 11.600 183.700 ;
        RECT 22.000 183.600 22.800 183.700 ;
        RECT 193.200 184.300 194.000 184.400 ;
        RECT 198.000 184.300 198.800 184.400 ;
        RECT 193.200 183.700 198.800 184.300 ;
        RECT 193.200 183.600 194.000 183.700 ;
        RECT 198.000 183.600 198.800 183.700 ;
        RECT 17.200 182.300 18.000 182.400 ;
        RECT 46.000 182.300 46.800 182.400 ;
        RECT 17.200 181.700 46.800 182.300 ;
        RECT 17.200 181.600 18.000 181.700 ;
        RECT 46.000 181.600 46.800 181.700 ;
        RECT 84.400 182.300 85.200 182.400 ;
        RECT 90.800 182.300 91.600 182.400 ;
        RECT 95.600 182.300 96.400 182.400 ;
        RECT 84.400 181.700 96.400 182.300 ;
        RECT 84.400 181.600 85.200 181.700 ;
        RECT 90.800 181.600 91.600 181.700 ;
        RECT 95.600 181.600 96.400 181.700 ;
        RECT 177.200 182.300 178.000 182.400 ;
        RECT 202.800 182.300 203.600 182.400 ;
        RECT 177.200 181.700 203.600 182.300 ;
        RECT 177.200 181.600 178.000 181.700 ;
        RECT 202.800 181.600 203.600 181.700 ;
        RECT 172.400 180.300 173.200 180.400 ;
        RECT 178.800 180.300 179.600 180.400 ;
        RECT 172.400 179.700 179.600 180.300 ;
        RECT 172.400 179.600 173.200 179.700 ;
        RECT 178.800 179.600 179.600 179.700 ;
        RECT 161.200 178.300 162.000 178.400 ;
        RECT 170.800 178.300 171.600 178.400 ;
        RECT 161.200 177.700 171.600 178.300 ;
        RECT 161.200 177.600 162.000 177.700 ;
        RECT 170.800 177.600 171.600 177.700 ;
        RECT 39.600 176.300 40.400 176.400 ;
        RECT 49.200 176.300 50.000 176.400 ;
        RECT 39.600 175.700 50.000 176.300 ;
        RECT 39.600 175.600 40.400 175.700 ;
        RECT 49.200 175.600 50.000 175.700 ;
        RECT 52.400 176.300 53.200 176.400 ;
        RECT 68.400 176.300 69.200 176.400 ;
        RECT 87.600 176.300 88.400 176.400 ;
        RECT 102.000 176.300 102.800 176.400 ;
        RECT 108.400 176.300 109.200 176.400 ;
        RECT 52.400 175.700 109.200 176.300 ;
        RECT 52.400 175.600 53.200 175.700 ;
        RECT 68.400 175.600 69.200 175.700 ;
        RECT 87.600 175.600 88.400 175.700 ;
        RECT 102.000 175.600 102.800 175.700 ;
        RECT 108.400 175.600 109.200 175.700 ;
        RECT 135.600 176.300 136.400 176.400 ;
        RECT 159.600 176.300 160.400 176.400 ;
        RECT 162.800 176.300 163.600 176.400 ;
        RECT 166.000 176.300 166.800 176.400 ;
        RECT 135.600 175.700 166.800 176.300 ;
        RECT 135.600 175.600 136.400 175.700 ;
        RECT 159.600 175.600 160.400 175.700 ;
        RECT 162.800 175.600 163.600 175.700 ;
        RECT 166.000 175.600 166.800 175.700 ;
        RECT 167.600 176.300 168.400 176.400 ;
        RECT 190.000 176.300 190.800 176.400 ;
        RECT 207.600 176.300 208.400 176.400 ;
        RECT 167.600 175.700 208.400 176.300 ;
        RECT 167.600 175.600 168.400 175.700 ;
        RECT 190.000 175.600 190.800 175.700 ;
        RECT 207.600 175.600 208.400 175.700 ;
        RECT 70.000 174.300 70.800 174.400 ;
        RECT 78.000 174.300 78.800 174.400 ;
        RECT 70.000 173.700 78.800 174.300 ;
        RECT 70.000 173.600 70.800 173.700 ;
        RECT 78.000 173.600 78.800 173.700 ;
        RECT 143.600 174.300 144.400 174.400 ;
        RECT 162.800 174.300 163.600 174.400 ;
        RECT 143.600 173.700 163.600 174.300 ;
        RECT 143.600 173.600 144.400 173.700 ;
        RECT 162.800 173.600 163.600 173.700 ;
        RECT 186.800 174.300 187.600 174.400 ;
        RECT 191.600 174.300 192.400 174.400 ;
        RECT 186.800 173.700 192.400 174.300 ;
        RECT 186.800 173.600 187.600 173.700 ;
        RECT 191.600 173.600 192.400 173.700 ;
        RECT 44.400 172.300 45.200 172.400 ;
        RECT 47.600 172.300 48.400 172.400 ;
        RECT 44.400 171.700 48.400 172.300 ;
        RECT 44.400 171.600 45.200 171.700 ;
        RECT 47.600 171.600 48.400 171.700 ;
        RECT 142.000 171.600 142.800 172.400 ;
        RECT 177.200 172.300 178.000 172.400 ;
        RECT 185.200 172.300 186.000 172.400 ;
        RECT 177.200 171.700 186.000 172.300 ;
        RECT 177.200 171.600 178.000 171.700 ;
        RECT 185.200 171.600 186.000 171.700 ;
        RECT 201.200 172.300 202.000 172.400 ;
        RECT 206.000 172.300 206.800 172.400 ;
        RECT 214.000 172.300 214.800 172.400 ;
        RECT 201.200 171.700 214.800 172.300 ;
        RECT 201.200 171.600 202.000 171.700 ;
        RECT 206.000 171.600 206.800 171.700 ;
        RECT 214.000 171.600 214.800 171.700 ;
        RECT 49.200 170.300 50.000 170.400 ;
        RECT 54.000 170.300 54.800 170.400 ;
        RECT 68.400 170.300 69.200 170.400 ;
        RECT 71.600 170.300 72.400 170.400 ;
        RECT 49.200 169.700 72.400 170.300 ;
        RECT 49.200 169.600 50.000 169.700 ;
        RECT 54.000 169.600 54.800 169.700 ;
        RECT 68.400 169.600 69.200 169.700 ;
        RECT 71.600 169.600 72.400 169.700 ;
        RECT 116.400 170.300 117.200 170.400 ;
        RECT 146.800 170.300 147.600 170.400 ;
        RECT 116.400 169.700 147.600 170.300 ;
        RECT 116.400 169.600 117.200 169.700 ;
        RECT 146.800 169.600 147.600 169.700 ;
        RECT 162.800 170.300 163.600 170.400 ;
        RECT 182.000 170.300 182.800 170.400 ;
        RECT 162.800 169.700 182.800 170.300 ;
        RECT 162.800 169.600 163.600 169.700 ;
        RECT 182.000 169.600 182.800 169.700 ;
        RECT 28.400 168.300 29.200 168.400 ;
        RECT 42.800 168.300 43.600 168.400 ;
        RECT 28.400 167.700 43.600 168.300 ;
        RECT 28.400 167.600 29.200 167.700 ;
        RECT 42.800 167.600 43.600 167.700 ;
        RECT 46.000 168.300 46.800 168.400 ;
        RECT 49.200 168.300 50.000 168.400 ;
        RECT 46.000 167.700 50.000 168.300 ;
        RECT 46.000 167.600 46.800 167.700 ;
        RECT 49.200 167.600 50.000 167.700 ;
        RECT 172.400 160.300 173.200 160.400 ;
        RECT 180.400 160.300 181.200 160.400 ;
        RECT 172.400 159.700 181.200 160.300 ;
        RECT 172.400 159.600 173.200 159.700 ;
        RECT 180.400 159.600 181.200 159.700 ;
        RECT 108.400 158.300 109.200 158.400 ;
        RECT 111.600 158.300 112.400 158.400 ;
        RECT 108.400 157.700 112.400 158.300 ;
        RECT 108.400 157.600 109.200 157.700 ;
        RECT 111.600 157.600 112.400 157.700 ;
        RECT 161.200 158.300 162.000 158.400 ;
        RECT 167.600 158.300 168.400 158.400 ;
        RECT 161.200 157.700 168.400 158.300 ;
        RECT 161.200 157.600 162.000 157.700 ;
        RECT 167.600 157.600 168.400 157.700 ;
        RECT 20.400 154.300 21.200 154.400 ;
        RECT 66.800 154.300 67.600 154.400 ;
        RECT 20.400 153.700 67.600 154.300 ;
        RECT 20.400 153.600 21.200 153.700 ;
        RECT 66.800 153.600 67.600 153.700 ;
        RECT 34.800 152.300 35.600 152.400 ;
        RECT 41.200 152.300 42.000 152.400 ;
        RECT 34.800 151.700 42.000 152.300 ;
        RECT 34.800 151.600 35.600 151.700 ;
        RECT 41.200 151.600 42.000 151.700 ;
        RECT 14.000 150.300 14.800 150.400 ;
        RECT 18.800 150.300 19.600 150.400 ;
        RECT 14.000 149.700 19.600 150.300 ;
        RECT 14.000 149.600 14.800 149.700 ;
        RECT 18.800 149.600 19.600 149.700 ;
        RECT 38.000 150.300 38.800 150.400 ;
        RECT 55.600 150.300 56.400 150.400 ;
        RECT 38.000 149.700 56.400 150.300 ;
        RECT 38.000 149.600 38.800 149.700 ;
        RECT 55.600 149.600 56.400 149.700 ;
        RECT 153.200 150.300 154.000 150.400 ;
        RECT 177.200 150.300 178.000 150.400 ;
        RECT 153.200 149.700 178.000 150.300 ;
        RECT 153.200 149.600 154.000 149.700 ;
        RECT 177.200 149.600 178.000 149.700 ;
        RECT 9.200 148.300 10.000 148.400 ;
        RECT 14.000 148.300 14.800 148.400 ;
        RECT 34.800 148.300 35.600 148.400 ;
        RECT 9.200 147.700 35.600 148.300 ;
        RECT 9.200 147.600 10.000 147.700 ;
        RECT 14.000 147.600 14.800 147.700 ;
        RECT 34.800 147.600 35.600 147.700 ;
        RECT 36.400 148.300 37.200 148.400 ;
        RECT 52.400 148.300 53.200 148.400 ;
        RECT 36.400 147.700 53.200 148.300 ;
        RECT 36.400 147.600 37.200 147.700 ;
        RECT 52.400 147.600 53.200 147.700 ;
        RECT 82.800 148.300 83.600 148.400 ;
        RECT 92.400 148.300 93.200 148.400 ;
        RECT 82.800 147.700 93.200 148.300 ;
        RECT 82.800 147.600 83.600 147.700 ;
        RECT 92.400 147.600 93.200 147.700 ;
        RECT 110.000 148.300 110.800 148.400 ;
        RECT 113.200 148.300 114.000 148.400 ;
        RECT 132.400 148.300 133.200 148.400 ;
        RECT 110.000 147.700 133.200 148.300 ;
        RECT 110.000 147.600 110.800 147.700 ;
        RECT 113.200 147.600 114.000 147.700 ;
        RECT 132.400 147.600 133.200 147.700 ;
        RECT 142.000 148.300 142.800 148.400 ;
        RECT 170.800 148.300 171.600 148.400 ;
        RECT 142.000 147.700 171.600 148.300 ;
        RECT 142.000 147.600 142.800 147.700 ;
        RECT 170.800 147.600 171.600 147.700 ;
        RECT 186.800 148.300 187.600 148.400 ;
        RECT 199.600 148.300 200.400 148.400 ;
        RECT 186.800 147.700 200.400 148.300 ;
        RECT 186.800 147.600 187.600 147.700 ;
        RECT 199.600 147.600 200.400 147.700 ;
        RECT 4.400 146.300 5.200 146.400 ;
        RECT 10.800 146.300 11.600 146.400 ;
        RECT 28.400 146.300 29.200 146.400 ;
        RECT 38.000 146.300 38.800 146.400 ;
        RECT 4.400 145.700 38.800 146.300 ;
        RECT 4.400 145.600 5.200 145.700 ;
        RECT 10.800 145.600 11.600 145.700 ;
        RECT 28.400 145.600 29.200 145.700 ;
        RECT 38.000 145.600 38.800 145.700 ;
        RECT 55.600 146.300 56.400 146.400 ;
        RECT 82.800 146.300 83.600 146.400 ;
        RECT 55.600 145.700 83.600 146.300 ;
        RECT 55.600 145.600 56.400 145.700 ;
        RECT 82.800 145.600 83.600 145.700 ;
        RECT 119.600 146.300 120.400 146.400 ;
        RECT 127.600 146.300 128.400 146.400 ;
        RECT 145.200 146.300 146.000 146.400 ;
        RECT 190.000 146.300 190.800 146.400 ;
        RECT 193.200 146.300 194.000 146.400 ;
        RECT 119.600 145.700 194.000 146.300 ;
        RECT 119.600 145.600 120.400 145.700 ;
        RECT 127.600 145.600 128.400 145.700 ;
        RECT 145.200 145.600 146.000 145.700 ;
        RECT 190.000 145.600 190.800 145.700 ;
        RECT 193.200 145.600 194.000 145.700 ;
        RECT 14.000 144.300 14.800 144.400 ;
        RECT 20.400 144.300 21.200 144.400 ;
        RECT 14.000 143.700 21.200 144.300 ;
        RECT 14.000 143.600 14.800 143.700 ;
        RECT 20.400 143.600 21.200 143.700 ;
        RECT 22.000 144.300 22.800 144.400 ;
        RECT 25.200 144.300 26.000 144.400 ;
        RECT 22.000 143.700 26.000 144.300 ;
        RECT 22.000 143.600 22.800 143.700 ;
        RECT 25.200 143.600 26.000 143.700 ;
        RECT 86.000 142.300 86.800 142.400 ;
        RECT 92.400 142.300 93.200 142.400 ;
        RECT 86.000 141.700 93.200 142.300 ;
        RECT 86.000 141.600 86.800 141.700 ;
        RECT 92.400 141.600 93.200 141.700 ;
        RECT 145.200 140.300 146.000 140.400 ;
        RECT 150.000 140.300 150.800 140.400 ;
        RECT 145.200 139.700 150.800 140.300 ;
        RECT 145.200 139.600 146.000 139.700 ;
        RECT 150.000 139.600 150.800 139.700 ;
        RECT 18.800 138.300 19.600 138.400 ;
        RECT 55.600 138.300 56.400 138.400 ;
        RECT 18.800 137.700 56.400 138.300 ;
        RECT 18.800 137.600 19.600 137.700 ;
        RECT 55.600 137.600 56.400 137.700 ;
        RECT 188.400 138.300 189.200 138.400 ;
        RECT 207.600 138.300 208.400 138.400 ;
        RECT 188.400 137.700 208.400 138.300 ;
        RECT 188.400 137.600 189.200 137.700 ;
        RECT 207.600 137.600 208.400 137.700 ;
        RECT 36.400 136.300 37.200 136.400 ;
        RECT 58.800 136.300 59.600 136.400 ;
        RECT 36.400 135.700 59.600 136.300 ;
        RECT 36.400 135.600 37.200 135.700 ;
        RECT 58.800 135.600 59.600 135.700 ;
        RECT 82.800 136.300 83.600 136.400 ;
        RECT 95.600 136.300 96.400 136.400 ;
        RECT 82.800 135.700 96.400 136.300 ;
        RECT 82.800 135.600 83.600 135.700 ;
        RECT 95.600 135.600 96.400 135.700 ;
        RECT 170.800 136.300 171.600 136.400 ;
        RECT 183.600 136.300 184.400 136.400 ;
        RECT 170.800 135.700 184.400 136.300 ;
        RECT 170.800 135.600 171.600 135.700 ;
        RECT 183.600 135.600 184.400 135.700 ;
        RECT 193.200 136.300 194.000 136.400 ;
        RECT 196.400 136.300 197.200 136.400 ;
        RECT 193.200 135.700 197.200 136.300 ;
        RECT 193.200 135.600 194.000 135.700 ;
        RECT 196.400 135.600 197.200 135.700 ;
        RECT 41.200 134.300 42.000 134.400 ;
        RECT 49.200 134.300 50.000 134.400 ;
        RECT 41.200 133.700 50.000 134.300 ;
        RECT 41.200 133.600 42.000 133.700 ;
        RECT 49.200 133.600 50.000 133.700 ;
        RECT 110.000 134.300 110.800 134.400 ;
        RECT 118.000 134.300 118.800 134.400 ;
        RECT 110.000 133.700 118.800 134.300 ;
        RECT 110.000 133.600 110.800 133.700 ;
        RECT 118.000 133.600 118.800 133.700 ;
        RECT 122.800 134.300 123.600 134.400 ;
        RECT 166.000 134.300 166.800 134.400 ;
        RECT 214.000 134.300 214.800 134.400 ;
        RECT 122.800 133.700 214.800 134.300 ;
        RECT 122.800 133.600 123.600 133.700 ;
        RECT 166.000 133.600 166.800 133.700 ;
        RECT 214.000 133.600 214.800 133.700 ;
        RECT 31.600 132.300 32.400 132.400 ;
        RECT 46.000 132.300 46.800 132.400 ;
        RECT 31.600 131.700 46.800 132.300 ;
        RECT 31.600 131.600 32.400 131.700 ;
        RECT 46.000 131.600 46.800 131.700 ;
        RECT 127.600 132.300 128.400 132.400 ;
        RECT 146.800 132.300 147.600 132.400 ;
        RECT 127.600 131.700 147.600 132.300 ;
        RECT 127.600 131.600 128.400 131.700 ;
        RECT 146.800 131.600 147.600 131.700 ;
        RECT 172.400 132.300 173.200 132.400 ;
        RECT 193.200 132.300 194.000 132.400 ;
        RECT 172.400 131.700 194.000 132.300 ;
        RECT 172.400 131.600 173.200 131.700 ;
        RECT 193.200 131.600 194.000 131.700 ;
        RECT 118.000 130.300 118.800 130.400 ;
        RECT 132.400 130.300 133.200 130.400 ;
        RECT 185.200 130.300 186.000 130.400 ;
        RECT 118.000 129.700 186.000 130.300 ;
        RECT 118.000 129.600 118.800 129.700 ;
        RECT 132.400 129.600 133.200 129.700 ;
        RECT 185.200 129.600 186.000 129.700 ;
        RECT 54.000 128.300 54.800 128.400 ;
        RECT 86.000 128.300 86.800 128.400 ;
        RECT 54.000 127.700 86.800 128.300 ;
        RECT 54.000 127.600 54.800 127.700 ;
        RECT 86.000 127.600 86.800 127.700 ;
        RECT 116.400 128.300 117.200 128.400 ;
        RECT 129.200 128.300 130.000 128.400 ;
        RECT 116.400 127.700 130.000 128.300 ;
        RECT 116.400 127.600 117.200 127.700 ;
        RECT 129.200 127.600 130.000 127.700 ;
        RECT 167.600 128.300 168.400 128.400 ;
        RECT 194.800 128.300 195.600 128.400 ;
        RECT 210.800 128.300 211.600 128.400 ;
        RECT 167.600 127.700 211.600 128.300 ;
        RECT 167.600 127.600 168.400 127.700 ;
        RECT 194.800 127.600 195.600 127.700 ;
        RECT 210.800 127.600 211.600 127.700 ;
        RECT 169.200 120.300 170.000 120.400 ;
        RECT 190.000 120.300 190.800 120.400 ;
        RECT 191.600 120.300 192.400 120.400 ;
        RECT 169.200 119.700 192.400 120.300 ;
        RECT 169.200 119.600 170.000 119.700 ;
        RECT 190.000 119.600 190.800 119.700 ;
        RECT 191.600 119.600 192.400 119.700 ;
        RECT 9.200 118.300 10.000 118.400 ;
        RECT 46.000 118.300 46.800 118.400 ;
        RECT 60.400 118.300 61.200 118.400 ;
        RECT 100.400 118.300 101.200 118.400 ;
        RECT 9.200 117.700 101.200 118.300 ;
        RECT 9.200 117.600 10.000 117.700 ;
        RECT 46.000 117.600 46.800 117.700 ;
        RECT 60.400 117.600 61.200 117.700 ;
        RECT 100.400 117.600 101.200 117.700 ;
        RECT 31.600 114.300 32.400 114.400 ;
        RECT 44.400 114.300 45.200 114.400 ;
        RECT 31.600 113.700 45.200 114.300 ;
        RECT 31.600 113.600 32.400 113.700 ;
        RECT 44.400 113.600 45.200 113.700 ;
        RECT 23.600 112.300 24.400 112.400 ;
        RECT 28.400 112.300 29.200 112.400 ;
        RECT 23.600 111.700 29.200 112.300 ;
        RECT 23.600 111.600 24.400 111.700 ;
        RECT 28.400 111.600 29.200 111.700 ;
        RECT 26.800 110.300 27.600 110.400 ;
        RECT 30.000 110.300 30.800 110.400 ;
        RECT 26.800 109.700 30.800 110.300 ;
        RECT 26.800 109.600 27.600 109.700 ;
        RECT 30.000 109.600 30.800 109.700 ;
        RECT 46.000 110.300 46.800 110.400 ;
        RECT 58.800 110.300 59.600 110.400 ;
        RECT 68.400 110.300 69.200 110.400 ;
        RECT 46.000 109.700 69.200 110.300 ;
        RECT 46.000 109.600 46.800 109.700 ;
        RECT 58.800 109.600 59.600 109.700 ;
        RECT 68.400 109.600 69.200 109.700 ;
        RECT 79.600 110.300 80.400 110.400 ;
        RECT 103.600 110.300 104.400 110.400 ;
        RECT 79.600 109.700 104.400 110.300 ;
        RECT 79.600 109.600 80.400 109.700 ;
        RECT 103.600 109.600 104.400 109.700 ;
        RECT 129.200 109.600 130.000 110.400 ;
        RECT 134.000 110.300 134.800 110.400 ;
        RECT 137.200 110.300 138.000 110.400 ;
        RECT 138.800 110.300 139.600 110.400 ;
        RECT 134.000 109.700 139.600 110.300 ;
        RECT 134.000 109.600 134.800 109.700 ;
        RECT 137.200 109.600 138.000 109.700 ;
        RECT 138.800 109.600 139.600 109.700 ;
        RECT 159.600 110.300 160.400 110.400 ;
        RECT 178.800 110.300 179.600 110.400 ;
        RECT 159.600 109.700 179.600 110.300 ;
        RECT 159.600 109.600 160.400 109.700 ;
        RECT 178.800 109.600 179.600 109.700 ;
        RECT 4.400 108.300 5.200 108.400 ;
        RECT 10.800 108.300 11.600 108.400 ;
        RECT 22.000 108.300 22.800 108.400 ;
        RECT 4.400 107.700 22.800 108.300 ;
        RECT 4.400 107.600 5.200 107.700 ;
        RECT 10.800 107.600 11.600 107.700 ;
        RECT 22.000 107.600 22.800 107.700 ;
        RECT 89.200 108.300 90.000 108.400 ;
        RECT 114.800 108.300 115.600 108.400 ;
        RECT 89.200 107.700 115.600 108.300 ;
        RECT 89.200 107.600 90.000 107.700 ;
        RECT 114.800 107.600 115.600 107.700 ;
        RECT 124.400 108.300 125.200 108.400 ;
        RECT 134.000 108.300 134.800 108.400 ;
        RECT 124.400 107.700 134.800 108.300 ;
        RECT 124.400 107.600 125.200 107.700 ;
        RECT 134.000 107.600 134.800 107.700 ;
        RECT 148.400 108.300 149.200 108.400 ;
        RECT 177.200 108.300 178.000 108.400 ;
        RECT 148.400 107.700 178.000 108.300 ;
        RECT 148.400 107.600 149.200 107.700 ;
        RECT 177.200 107.600 178.000 107.700 ;
        RECT 54.000 106.300 54.800 106.400 ;
        RECT 76.400 106.300 77.200 106.400 ;
        RECT 54.000 105.700 77.200 106.300 ;
        RECT 54.000 105.600 54.800 105.700 ;
        RECT 76.400 105.600 77.200 105.700 ;
        RECT 15.600 104.300 16.400 104.400 ;
        RECT 22.000 104.300 22.800 104.400 ;
        RECT 15.600 103.700 22.800 104.300 ;
        RECT 15.600 103.600 16.400 103.700 ;
        RECT 22.000 103.600 22.800 103.700 ;
        RECT 164.400 104.300 165.200 104.400 ;
        RECT 183.600 104.300 184.400 104.400 ;
        RECT 191.600 104.300 192.400 104.400 ;
        RECT 164.400 103.700 192.400 104.300 ;
        RECT 164.400 103.600 165.200 103.700 ;
        RECT 183.600 103.600 184.400 103.700 ;
        RECT 191.600 103.600 192.400 103.700 ;
        RECT 202.800 104.300 203.600 104.400 ;
        RECT 207.600 104.300 208.400 104.400 ;
        RECT 202.800 103.700 208.400 104.300 ;
        RECT 202.800 103.600 203.600 103.700 ;
        RECT 207.600 103.600 208.400 103.700 ;
        RECT 14.000 102.300 14.800 102.400 ;
        RECT 20.400 102.300 21.200 102.400 ;
        RECT 14.000 101.700 21.200 102.300 ;
        RECT 14.000 101.600 14.800 101.700 ;
        RECT 20.400 101.600 21.200 101.700 ;
        RECT 25.200 102.300 26.000 102.400 ;
        RECT 38.000 102.300 38.800 102.400 ;
        RECT 25.200 101.700 38.800 102.300 ;
        RECT 25.200 101.600 26.000 101.700 ;
        RECT 38.000 101.600 38.800 101.700 ;
        RECT 145.200 102.300 146.000 102.400 ;
        RECT 151.600 102.300 152.400 102.400 ;
        RECT 145.200 101.700 152.400 102.300 ;
        RECT 145.200 101.600 146.000 101.700 ;
        RECT 151.600 101.600 152.400 101.700 ;
        RECT 188.400 102.300 189.200 102.400 ;
        RECT 207.600 102.300 208.400 102.400 ;
        RECT 188.400 101.700 208.400 102.300 ;
        RECT 188.400 101.600 189.200 101.700 ;
        RECT 207.600 101.600 208.400 101.700 ;
        RECT 39.600 96.300 40.400 96.400 ;
        RECT 94.000 96.300 94.800 96.400 ;
        RECT 100.400 96.300 101.200 96.400 ;
        RECT 39.600 95.700 101.200 96.300 ;
        RECT 39.600 95.600 40.400 95.700 ;
        RECT 94.000 95.600 94.800 95.700 ;
        RECT 100.400 95.600 101.200 95.700 ;
        RECT 111.600 96.300 112.400 96.400 ;
        RECT 126.000 96.300 126.800 96.400 ;
        RECT 111.600 95.700 126.800 96.300 ;
        RECT 111.600 95.600 112.400 95.700 ;
        RECT 126.000 95.600 126.800 95.700 ;
        RECT 151.600 96.300 152.400 96.400 ;
        RECT 164.400 96.300 165.200 96.400 ;
        RECT 151.600 95.700 165.200 96.300 ;
        RECT 151.600 95.600 152.400 95.700 ;
        RECT 164.400 95.600 165.200 95.700 ;
        RECT 30.000 94.300 30.800 94.400 ;
        RECT 57.200 94.300 58.000 94.400 ;
        RECT 30.000 93.700 58.000 94.300 ;
        RECT 30.000 93.600 30.800 93.700 ;
        RECT 57.200 93.600 58.000 93.700 ;
        RECT 100.400 94.300 101.200 94.400 ;
        RECT 103.600 94.300 104.400 94.400 ;
        RECT 100.400 93.700 104.400 94.300 ;
        RECT 100.400 93.600 101.200 93.700 ;
        RECT 103.600 93.600 104.400 93.700 ;
        RECT 108.400 94.300 109.200 94.400 ;
        RECT 129.200 94.300 130.000 94.400 ;
        RECT 108.400 93.700 130.000 94.300 ;
        RECT 108.400 93.600 109.200 93.700 ;
        RECT 129.200 93.600 130.000 93.700 ;
        RECT 161.200 94.300 162.000 94.400 ;
        RECT 182.000 94.300 182.800 94.400 ;
        RECT 161.200 93.700 182.800 94.300 ;
        RECT 161.200 93.600 162.000 93.700 ;
        RECT 182.000 93.600 182.800 93.700 ;
        RECT 198.000 94.300 198.800 94.400 ;
        RECT 202.800 94.300 203.600 94.400 ;
        RECT 214.000 94.300 214.800 94.400 ;
        RECT 198.000 93.700 214.800 94.300 ;
        RECT 198.000 93.600 198.800 93.700 ;
        RECT 202.800 93.600 203.600 93.700 ;
        RECT 214.000 93.600 214.800 93.700 ;
        RECT 82.800 92.300 83.600 92.400 ;
        RECT 95.600 92.300 96.400 92.400 ;
        RECT 82.800 91.700 96.400 92.300 ;
        RECT 82.800 91.600 83.600 91.700 ;
        RECT 95.600 91.600 96.400 91.700 ;
        RECT 138.800 92.300 139.600 92.400 ;
        RECT 151.600 92.300 152.400 92.400 ;
        RECT 138.800 91.700 152.400 92.300 ;
        RECT 138.800 91.600 139.600 91.700 ;
        RECT 151.600 91.600 152.400 91.700 ;
        RECT 183.600 92.300 184.400 92.400 ;
        RECT 199.600 92.300 200.400 92.400 ;
        RECT 215.600 92.300 216.400 92.400 ;
        RECT 183.600 91.700 216.400 92.300 ;
        RECT 183.600 91.600 184.400 91.700 ;
        RECT 199.600 91.600 200.400 91.700 ;
        RECT 215.600 91.600 216.400 91.700 ;
        RECT 31.600 90.300 32.400 90.400 ;
        RECT 66.800 90.300 67.600 90.400 ;
        RECT 78.000 90.300 78.800 90.400 ;
        RECT 31.600 89.700 78.800 90.300 ;
        RECT 31.600 89.600 32.400 89.700 ;
        RECT 66.800 89.600 67.600 89.700 ;
        RECT 78.000 89.600 78.800 89.700 ;
        RECT 100.400 90.300 101.200 90.400 ;
        RECT 110.000 90.300 110.800 90.400 ;
        RECT 113.200 90.300 114.000 90.400 ;
        RECT 100.400 89.700 114.000 90.300 ;
        RECT 100.400 89.600 101.200 89.700 ;
        RECT 110.000 89.600 110.800 89.700 ;
        RECT 113.200 89.600 114.000 89.700 ;
        RECT 194.800 90.300 195.600 90.400 ;
        RECT 204.400 90.300 205.200 90.400 ;
        RECT 194.800 89.700 205.200 90.300 ;
        RECT 194.800 89.600 195.600 89.700 ;
        RECT 204.400 89.600 205.200 89.700 ;
        RECT 190.000 88.300 190.800 88.400 ;
        RECT 191.600 88.300 192.400 88.400 ;
        RECT 190.000 87.700 192.400 88.300 ;
        RECT 190.000 87.600 190.800 87.700 ;
        RECT 191.600 87.600 192.400 87.700 ;
        RECT 44.400 84.300 45.200 84.400 ;
        RECT 81.200 84.300 82.000 84.400 ;
        RECT 127.600 84.300 128.400 84.400 ;
        RECT 129.200 84.300 130.000 84.400 ;
        RECT 44.400 83.700 130.000 84.300 ;
        RECT 44.400 83.600 45.200 83.700 ;
        RECT 81.200 83.600 82.000 83.700 ;
        RECT 127.600 83.600 128.400 83.700 ;
        RECT 129.200 83.600 130.000 83.700 ;
        RECT 111.600 82.300 112.400 82.400 ;
        RECT 114.800 82.300 115.600 82.400 ;
        RECT 140.400 82.300 141.200 82.400 ;
        RECT 111.600 81.700 141.200 82.300 ;
        RECT 111.600 81.600 112.400 81.700 ;
        RECT 114.800 81.600 115.600 81.700 ;
        RECT 140.400 81.600 141.200 81.700 ;
        RECT 92.400 74.300 93.200 74.400 ;
        RECT 105.200 74.300 106.000 74.400 ;
        RECT 92.400 73.700 106.000 74.300 ;
        RECT 92.400 73.600 93.200 73.700 ;
        RECT 105.200 73.600 106.000 73.700 ;
        RECT 4.400 72.300 5.200 72.400 ;
        RECT 10.800 72.300 11.600 72.400 ;
        RECT 28.400 72.300 29.200 72.400 ;
        RECT 38.000 72.300 38.800 72.400 ;
        RECT 4.400 71.700 38.800 72.300 ;
        RECT 4.400 71.600 5.200 71.700 ;
        RECT 10.800 71.600 11.600 71.700 ;
        RECT 28.400 71.600 29.200 71.700 ;
        RECT 38.000 71.600 38.800 71.700 ;
        RECT 194.800 72.300 195.600 72.400 ;
        RECT 199.600 72.300 200.400 72.400 ;
        RECT 194.800 71.700 200.400 72.300 ;
        RECT 194.800 71.600 195.600 71.700 ;
        RECT 199.600 71.600 200.400 71.700 ;
        RECT 14.000 70.300 14.800 70.400 ;
        RECT 15.600 70.300 16.400 70.400 ;
        RECT 25.200 70.300 26.000 70.400 ;
        RECT 14.000 69.700 26.000 70.300 ;
        RECT 14.000 69.600 14.800 69.700 ;
        RECT 15.600 69.600 16.400 69.700 ;
        RECT 25.200 69.600 26.000 69.700 ;
        RECT 105.200 70.300 106.000 70.400 ;
        RECT 110.000 70.300 110.800 70.400 ;
        RECT 105.200 69.700 110.800 70.300 ;
        RECT 105.200 69.600 106.000 69.700 ;
        RECT 110.000 69.600 110.800 69.700 ;
        RECT 158.000 70.300 158.800 70.400 ;
        RECT 162.800 70.300 163.600 70.400 ;
        RECT 158.000 69.700 163.600 70.300 ;
        RECT 158.000 69.600 158.800 69.700 ;
        RECT 162.800 69.600 163.600 69.700 ;
        RECT 164.400 70.300 165.200 70.400 ;
        RECT 169.200 70.300 170.000 70.400 ;
        RECT 164.400 69.700 170.000 70.300 ;
        RECT 164.400 69.600 165.200 69.700 ;
        RECT 169.200 69.600 170.000 69.700 ;
        RECT 183.600 70.300 184.400 70.400 ;
        RECT 186.800 70.300 187.600 70.400 ;
        RECT 183.600 69.700 187.600 70.300 ;
        RECT 183.600 69.600 184.400 69.700 ;
        RECT 186.800 69.600 187.600 69.700 ;
        RECT 198.000 70.300 198.800 70.400 ;
        RECT 201.200 70.300 202.000 70.400 ;
        RECT 198.000 69.700 202.000 70.300 ;
        RECT 198.000 69.600 198.800 69.700 ;
        RECT 201.200 69.600 202.000 69.700 ;
        RECT 2.800 68.300 3.600 68.400 ;
        RECT 15.600 68.300 16.400 68.400 ;
        RECT 23.600 68.300 24.400 68.400 ;
        RECT 2.800 67.700 24.400 68.300 ;
        RECT 2.800 67.600 3.600 67.700 ;
        RECT 15.600 67.600 16.400 67.700 ;
        RECT 23.600 67.600 24.400 67.700 ;
        RECT 50.800 68.300 51.600 68.400 ;
        RECT 71.600 68.300 72.400 68.400 ;
        RECT 50.800 67.700 72.400 68.300 ;
        RECT 50.800 67.600 51.600 67.700 ;
        RECT 71.600 67.600 72.400 67.700 ;
        RECT 151.600 68.300 152.400 68.400 ;
        RECT 167.600 68.300 168.400 68.400 ;
        RECT 174.000 68.300 174.800 68.400 ;
        RECT 185.200 68.300 186.000 68.400 ;
        RECT 151.600 67.700 186.000 68.300 ;
        RECT 151.600 67.600 152.400 67.700 ;
        RECT 167.600 67.600 168.400 67.700 ;
        RECT 174.000 67.600 174.800 67.700 ;
        RECT 185.200 67.600 186.000 67.700 ;
        RECT 190.000 68.300 190.800 68.400 ;
        RECT 196.400 68.300 197.200 68.400 ;
        RECT 209.200 68.300 210.000 68.400 ;
        RECT 190.000 67.700 210.000 68.300 ;
        RECT 190.000 67.600 190.800 67.700 ;
        RECT 196.400 67.600 197.200 67.700 ;
        RECT 209.200 67.600 210.000 67.700 ;
        RECT 18.800 66.300 19.600 66.400 ;
        RECT 23.600 66.300 24.400 66.400 ;
        RECT 54.000 66.300 54.800 66.400 ;
        RECT 68.400 66.300 69.200 66.400 ;
        RECT 89.200 66.300 90.000 66.400 ;
        RECT 18.800 65.700 90.000 66.300 ;
        RECT 18.800 65.600 19.600 65.700 ;
        RECT 23.600 65.600 24.400 65.700 ;
        RECT 54.000 65.600 54.800 65.700 ;
        RECT 68.400 65.600 69.200 65.700 ;
        RECT 89.200 65.600 90.000 65.700 ;
        RECT 110.000 66.300 110.800 66.400 ;
        RECT 113.200 66.300 114.000 66.400 ;
        RECT 110.000 65.700 114.000 66.300 ;
        RECT 110.000 65.600 110.800 65.700 ;
        RECT 113.200 65.600 114.000 65.700 ;
        RECT 148.400 66.300 149.200 66.400 ;
        RECT 151.600 66.300 152.400 66.400 ;
        RECT 148.400 65.700 152.400 66.300 ;
        RECT 148.400 65.600 149.200 65.700 ;
        RECT 151.600 65.600 152.400 65.700 ;
        RECT 161.200 66.300 162.000 66.400 ;
        RECT 164.400 66.300 165.200 66.400 ;
        RECT 161.200 65.700 165.200 66.300 ;
        RECT 161.200 65.600 162.000 65.700 ;
        RECT 164.400 65.600 165.200 65.700 ;
        RECT 186.800 66.300 187.600 66.400 ;
        RECT 198.000 66.300 198.800 66.400 ;
        RECT 210.800 66.300 211.600 66.400 ;
        RECT 186.800 65.700 211.600 66.300 ;
        RECT 186.800 65.600 187.600 65.700 ;
        RECT 198.000 65.600 198.800 65.700 ;
        RECT 210.800 65.600 211.600 65.700 ;
        RECT 177.200 63.600 178.000 64.400 ;
        RECT 199.600 64.300 200.400 64.400 ;
        RECT 204.400 64.300 205.200 64.400 ;
        RECT 199.600 63.700 205.200 64.300 ;
        RECT 199.600 63.600 200.400 63.700 ;
        RECT 204.400 63.600 205.200 63.700 ;
        RECT 10.800 60.300 11.600 60.400 ;
        RECT 14.000 60.300 14.800 60.400 ;
        RECT 10.800 59.700 14.800 60.300 ;
        RECT 10.800 59.600 11.600 59.700 ;
        RECT 14.000 59.600 14.800 59.700 ;
        RECT 9.200 56.300 10.000 56.400 ;
        RECT 41.200 56.300 42.000 56.400 ;
        RECT 52.400 56.300 53.200 56.400 ;
        RECT 55.600 56.300 56.400 56.400 ;
        RECT 9.200 55.700 56.400 56.300 ;
        RECT 9.200 55.600 10.000 55.700 ;
        RECT 41.200 55.600 42.000 55.700 ;
        RECT 52.400 55.600 53.200 55.700 ;
        RECT 55.600 55.600 56.400 55.700 ;
        RECT 73.200 56.300 74.000 56.400 ;
        RECT 92.400 56.300 93.200 56.400 ;
        RECT 105.200 56.300 106.000 56.400 ;
        RECT 73.200 55.700 106.000 56.300 ;
        RECT 73.200 55.600 74.000 55.700 ;
        RECT 92.400 55.600 93.200 55.700 ;
        RECT 105.200 55.600 106.000 55.700 ;
        RECT 111.600 56.300 112.400 56.400 ;
        RECT 119.600 56.300 120.400 56.400 ;
        RECT 111.600 55.700 120.400 56.300 ;
        RECT 111.600 55.600 112.400 55.700 ;
        RECT 119.600 55.600 120.400 55.700 ;
        RECT 180.400 56.300 181.200 56.400 ;
        RECT 183.600 56.300 184.400 56.400 ;
        RECT 180.400 55.700 184.400 56.300 ;
        RECT 180.400 55.600 181.200 55.700 ;
        RECT 183.600 55.600 184.400 55.700 ;
        RECT 202.800 56.300 203.600 56.400 ;
        RECT 212.400 56.300 213.200 56.400 ;
        RECT 202.800 55.700 213.200 56.300 ;
        RECT 202.800 55.600 203.600 55.700 ;
        RECT 212.400 55.600 213.200 55.700 ;
        RECT 22.000 54.300 22.800 54.400 ;
        RECT 36.400 54.300 37.200 54.400 ;
        RECT 22.000 53.700 37.200 54.300 ;
        RECT 22.000 53.600 22.800 53.700 ;
        RECT 36.400 53.600 37.200 53.700 ;
        RECT 50.800 54.300 51.600 54.400 ;
        RECT 65.200 54.300 66.000 54.400 ;
        RECT 50.800 53.700 66.000 54.300 ;
        RECT 50.800 53.600 51.600 53.700 ;
        RECT 65.200 53.600 66.000 53.700 ;
        RECT 82.800 54.300 83.600 54.400 ;
        RECT 103.600 54.300 104.400 54.400 ;
        RECT 82.800 53.700 104.400 54.300 ;
        RECT 82.800 53.600 83.600 53.700 ;
        RECT 103.600 53.600 104.400 53.700 ;
        RECT 137.200 54.300 138.000 54.400 ;
        RECT 150.000 54.300 150.800 54.400 ;
        RECT 137.200 53.700 150.800 54.300 ;
        RECT 137.200 53.600 138.000 53.700 ;
        RECT 150.000 53.600 150.800 53.700 ;
        RECT 177.200 54.300 178.000 54.400 ;
        RECT 201.200 54.300 202.000 54.400 ;
        RECT 177.200 53.700 202.000 54.300 ;
        RECT 177.200 53.600 178.000 53.700 ;
        RECT 201.200 53.600 202.000 53.700 ;
        RECT 30.000 52.300 30.800 52.400 ;
        RECT 33.200 52.300 34.000 52.400 ;
        RECT 30.000 51.700 34.000 52.300 ;
        RECT 30.000 51.600 30.800 51.700 ;
        RECT 33.200 51.600 34.000 51.700 ;
        RECT 39.600 52.300 40.400 52.400 ;
        RECT 54.000 52.300 54.800 52.400 ;
        RECT 39.600 51.700 54.800 52.300 ;
        RECT 39.600 51.600 40.400 51.700 ;
        RECT 54.000 51.600 54.800 51.700 ;
        RECT 79.600 52.300 80.400 52.400 ;
        RECT 86.000 52.300 86.800 52.400 ;
        RECT 79.600 51.700 86.800 52.300 ;
        RECT 79.600 51.600 80.400 51.700 ;
        RECT 86.000 51.600 86.800 51.700 ;
        RECT 87.600 52.300 88.400 52.400 ;
        RECT 92.400 52.300 93.200 52.400 ;
        RECT 102.000 52.300 102.800 52.400 ;
        RECT 110.000 52.300 110.800 52.400 ;
        RECT 87.600 51.700 110.800 52.300 ;
        RECT 87.600 51.600 88.400 51.700 ;
        RECT 92.400 51.600 93.200 51.700 ;
        RECT 102.000 51.600 102.800 51.700 ;
        RECT 110.000 51.600 110.800 51.700 ;
        RECT 111.600 52.300 112.400 52.400 ;
        RECT 114.800 52.300 115.600 52.400 ;
        RECT 111.600 51.700 115.600 52.300 ;
        RECT 111.600 51.600 112.400 51.700 ;
        RECT 114.800 51.600 115.600 51.700 ;
        RECT 119.600 52.300 120.400 52.400 ;
        RECT 122.800 52.300 123.600 52.400 ;
        RECT 119.600 51.700 123.600 52.300 ;
        RECT 119.600 51.600 120.400 51.700 ;
        RECT 122.800 51.600 123.600 51.700 ;
        RECT 148.400 52.300 149.200 52.400 ;
        RECT 167.600 52.300 168.400 52.400 ;
        RECT 148.400 51.700 168.400 52.300 ;
        RECT 148.400 51.600 149.200 51.700 ;
        RECT 167.600 51.600 168.400 51.700 ;
        RECT 55.600 50.300 56.400 50.400 ;
        RECT 90.800 50.300 91.600 50.400 ;
        RECT 55.600 49.700 91.600 50.300 ;
        RECT 55.600 49.600 56.400 49.700 ;
        RECT 90.800 49.600 91.600 49.700 ;
        RECT 103.600 50.300 104.400 50.400 ;
        RECT 106.800 50.300 107.600 50.400 ;
        RECT 103.600 49.700 107.600 50.300 ;
        RECT 103.600 49.600 104.400 49.700 ;
        RECT 106.800 49.600 107.600 49.700 ;
        RECT 31.600 48.300 32.400 48.400 ;
        RECT 36.400 48.300 37.200 48.400 ;
        RECT 31.600 47.700 37.200 48.300 ;
        RECT 31.600 47.600 32.400 47.700 ;
        RECT 36.400 47.600 37.200 47.700 ;
        RECT 71.600 48.300 72.400 48.400 ;
        RECT 81.200 48.300 82.000 48.400 ;
        RECT 71.600 47.700 82.000 48.300 ;
        RECT 71.600 47.600 72.400 47.700 ;
        RECT 81.200 47.600 82.000 47.700 ;
        RECT 196.400 48.300 197.200 48.400 ;
        RECT 204.400 48.300 205.200 48.400 ;
        RECT 214.000 48.300 214.800 48.400 ;
        RECT 215.600 48.300 216.400 48.400 ;
        RECT 196.400 47.700 216.400 48.300 ;
        RECT 196.400 47.600 197.200 47.700 ;
        RECT 204.400 47.600 205.200 47.700 ;
        RECT 214.000 47.600 214.800 47.700 ;
        RECT 215.600 47.600 216.400 47.700 ;
        RECT 12.400 42.300 13.200 42.400 ;
        RECT 34.800 42.300 35.600 42.400 ;
        RECT 39.600 42.300 40.400 42.400 ;
        RECT 12.400 41.700 40.400 42.300 ;
        RECT 12.400 41.600 13.200 41.700 ;
        RECT 34.800 41.600 35.600 41.700 ;
        RECT 39.600 41.600 40.400 41.700 ;
        RECT 49.200 42.300 50.000 42.400 ;
        RECT 55.600 42.300 56.400 42.400 ;
        RECT 49.200 41.700 56.400 42.300 ;
        RECT 49.200 41.600 50.000 41.700 ;
        RECT 55.600 41.600 56.400 41.700 ;
        RECT 122.800 42.300 123.600 42.400 ;
        RECT 126.000 42.300 126.800 42.400 ;
        RECT 122.800 41.700 126.800 42.300 ;
        RECT 122.800 41.600 123.600 41.700 ;
        RECT 126.000 41.600 126.800 41.700 ;
        RECT 46.000 40.300 46.800 40.400 ;
        RECT 49.200 40.300 50.000 40.400 ;
        RECT 46.000 39.700 50.000 40.300 ;
        RECT 46.000 39.600 46.800 39.700 ;
        RECT 49.200 39.600 50.000 39.700 ;
        RECT 119.600 40.300 120.400 40.400 ;
        RECT 146.800 40.300 147.600 40.400 ;
        RECT 119.600 39.700 147.600 40.300 ;
        RECT 119.600 39.600 120.400 39.700 ;
        RECT 146.800 39.600 147.600 39.700 ;
        RECT 130.800 38.300 131.600 38.400 ;
        RECT 135.600 38.300 136.400 38.400 ;
        RECT 130.800 37.700 136.400 38.300 ;
        RECT 130.800 37.600 131.600 37.700 ;
        RECT 135.600 37.600 136.400 37.700 ;
        RECT 177.200 38.300 178.000 38.400 ;
        RECT 178.800 38.300 179.600 38.400 ;
        RECT 177.200 37.700 179.600 38.300 ;
        RECT 177.200 37.600 178.000 37.700 ;
        RECT 178.800 37.600 179.600 37.700 ;
        RECT 201.200 36.300 202.000 36.400 ;
        RECT 209.200 36.300 210.000 36.400 ;
        RECT 201.200 35.700 210.000 36.300 ;
        RECT 201.200 35.600 202.000 35.700 ;
        RECT 209.200 35.600 210.000 35.700 ;
        RECT 10.800 33.600 11.600 34.400 ;
        RECT 4.400 32.300 5.200 32.400 ;
        RECT 34.800 32.300 35.600 32.400 ;
        RECT 4.400 31.700 35.600 32.300 ;
        RECT 4.400 31.600 5.200 31.700 ;
        RECT 34.800 31.600 35.600 31.700 ;
        RECT 7.600 30.300 8.400 30.400 ;
        RECT 12.400 30.300 13.200 30.400 ;
        RECT 7.600 29.700 13.200 30.300 ;
        RECT 7.600 29.600 8.400 29.700 ;
        RECT 12.400 29.600 13.200 29.700 ;
        RECT 30.000 30.300 30.800 30.400 ;
        RECT 41.200 30.300 42.000 30.400 ;
        RECT 30.000 29.700 42.000 30.300 ;
        RECT 30.000 29.600 30.800 29.700 ;
        RECT 41.200 29.600 42.000 29.700 ;
        RECT 71.600 30.300 72.400 30.400 ;
        RECT 86.000 30.300 86.800 30.400 ;
        RECT 71.600 29.700 86.800 30.300 ;
        RECT 71.600 29.600 72.400 29.700 ;
        RECT 86.000 29.600 86.800 29.700 ;
        RECT 7.600 28.300 8.400 28.400 ;
        RECT 18.800 28.300 19.600 28.400 ;
        RECT 30.000 28.300 30.800 28.400 ;
        RECT 38.000 28.300 38.800 28.400 ;
        RECT 7.600 27.700 38.800 28.300 ;
        RECT 7.600 27.600 8.400 27.700 ;
        RECT 18.800 27.600 19.600 27.700 ;
        RECT 30.000 27.600 30.800 27.700 ;
        RECT 38.000 27.600 38.800 27.700 ;
        RECT 103.600 28.300 104.400 28.400 ;
        RECT 129.200 28.300 130.000 28.400 ;
        RECT 103.600 27.700 130.000 28.300 ;
        RECT 103.600 27.600 104.400 27.700 ;
        RECT 129.200 27.600 130.000 27.700 ;
        RECT 89.200 26.300 90.000 26.400 ;
        RECT 126.000 26.300 126.800 26.400 ;
        RECT 140.400 26.300 141.200 26.400 ;
        RECT 89.200 25.700 141.200 26.300 ;
        RECT 89.200 25.600 90.000 25.700 ;
        RECT 126.000 25.600 126.800 25.700 ;
        RECT 140.400 25.600 141.200 25.700 ;
        RECT 142.000 26.300 142.800 26.400 ;
        RECT 143.600 26.300 144.400 26.400 ;
        RECT 151.600 26.300 152.400 26.400 ;
        RECT 142.000 25.700 152.400 26.300 ;
        RECT 142.000 25.600 142.800 25.700 ;
        RECT 143.600 25.600 144.400 25.700 ;
        RECT 151.600 25.600 152.400 25.700 ;
        RECT 156.400 26.300 157.200 26.400 ;
        RECT 164.400 26.300 165.200 26.400 ;
        RECT 156.400 25.700 165.200 26.300 ;
        RECT 156.400 25.600 157.200 25.700 ;
        RECT 164.400 25.600 165.200 25.700 ;
        RECT 146.800 24.300 147.600 24.400 ;
        RECT 158.000 24.300 158.800 24.400 ;
        RECT 146.800 23.700 158.800 24.300 ;
        RECT 146.800 23.600 147.600 23.700 ;
        RECT 158.000 23.600 158.800 23.700 ;
        RECT 23.600 22.300 24.400 22.400 ;
        RECT 68.400 22.300 69.200 22.400 ;
        RECT 23.600 21.700 69.200 22.300 ;
        RECT 23.600 21.600 24.400 21.700 ;
        RECT 68.400 21.600 69.200 21.700 ;
        RECT 73.200 20.300 74.000 20.400 ;
        RECT 89.200 20.300 90.000 20.400 ;
        RECT 73.200 19.700 90.000 20.300 ;
        RECT 73.200 19.600 74.000 19.700 ;
        RECT 89.200 19.600 90.000 19.700 ;
        RECT 170.800 20.300 171.600 20.400 ;
        RECT 174.000 20.300 174.800 20.400 ;
        RECT 183.600 20.300 184.400 20.400 ;
        RECT 170.800 19.700 184.400 20.300 ;
        RECT 170.800 19.600 171.600 19.700 ;
        RECT 174.000 19.600 174.800 19.700 ;
        RECT 183.600 19.600 184.400 19.700 ;
        RECT 100.400 18.300 101.200 18.400 ;
        RECT 106.800 18.300 107.600 18.400 ;
        RECT 111.600 18.300 112.400 18.400 ;
        RECT 100.400 17.700 112.400 18.300 ;
        RECT 100.400 17.600 101.200 17.700 ;
        RECT 106.800 17.600 107.600 17.700 ;
        RECT 111.600 17.600 112.400 17.700 ;
        RECT 162.800 18.300 163.600 18.400 ;
        RECT 166.000 18.300 166.800 18.400 ;
        RECT 162.800 17.700 166.800 18.300 ;
        RECT 162.800 17.600 163.600 17.700 ;
        RECT 166.000 17.600 166.800 17.700 ;
        RECT 122.800 16.300 123.600 16.400 ;
        RECT 126.000 16.300 126.800 16.400 ;
        RECT 122.800 15.700 126.800 16.300 ;
        RECT 122.800 15.600 123.600 15.700 ;
        RECT 126.000 15.600 126.800 15.700 ;
        RECT 162.800 16.300 163.600 16.400 ;
        RECT 182.000 16.300 182.800 16.400 ;
        RECT 196.400 16.300 197.200 16.400 ;
        RECT 162.800 15.700 197.200 16.300 ;
        RECT 162.800 15.600 163.600 15.700 ;
        RECT 182.000 15.600 182.800 15.700 ;
        RECT 196.400 15.600 197.200 15.700 ;
        RECT 60.400 14.300 61.200 14.400 ;
        RECT 71.600 14.300 72.400 14.400 ;
        RECT 60.400 13.700 72.400 14.300 ;
        RECT 60.400 13.600 61.200 13.700 ;
        RECT 71.600 13.600 72.400 13.700 ;
        RECT 90.800 14.300 91.600 14.400 ;
        RECT 110.000 14.300 110.800 14.400 ;
        RECT 90.800 13.700 110.800 14.300 ;
        RECT 90.800 13.600 91.600 13.700 ;
        RECT 110.000 13.600 110.800 13.700 ;
        RECT 126.000 13.600 126.800 14.400 ;
        RECT 193.200 14.300 194.000 14.400 ;
        RECT 204.400 14.300 205.200 14.400 ;
        RECT 193.200 13.700 205.200 14.300 ;
        RECT 193.200 13.600 194.000 13.700 ;
        RECT 204.400 13.600 205.200 13.700 ;
        RECT 33.200 12.300 34.000 12.400 ;
        RECT 60.400 12.300 61.200 12.400 ;
        RECT 33.200 11.700 61.200 12.300 ;
        RECT 33.200 11.600 34.000 11.700 ;
        RECT 60.400 11.600 61.200 11.700 ;
        RECT 95.600 12.300 96.400 12.400 ;
        RECT 108.400 12.300 109.200 12.400 ;
        RECT 95.600 11.700 109.200 12.300 ;
        RECT 95.600 11.600 96.400 11.700 ;
        RECT 108.400 11.600 109.200 11.700 ;
        RECT 135.600 12.300 136.400 12.400 ;
        RECT 138.800 12.300 139.600 12.400 ;
        RECT 135.600 11.700 139.600 12.300 ;
        RECT 135.600 11.600 136.400 11.700 ;
        RECT 138.800 11.600 139.600 11.700 ;
      LAYER metal4 ;
        RECT 13.800 69.400 15.000 144.600 ;
        RECT 45.800 117.400 47.000 186.600 ;
        RECT 129.000 83.400 130.200 110.600 ;
        RECT 10.600 33.400 11.800 60.600 ;
        RECT 23.400 21.400 24.600 66.600 ;
        RECT 125.800 13.400 127.000 42.600 ;
        RECT 141.800 25.400 143.000 172.600 ;
        RECT 193.000 145.400 194.200 184.600 ;
        RECT 177.000 37.400 178.200 64.600 ;
        RECT 183.400 55.400 184.600 104.600 ;
        RECT 189.800 87.400 191.000 120.600 ;
  END
END cordic
END LIBRARY


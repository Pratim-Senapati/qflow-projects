* NGSPICE file created from noc_top.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

.subckt noc_top vdd gnd clk rst ext_data_in[0] ext_data_in[1] ext_data_in[2] ext_data_in[3]
+ ext_data_in[4] ext_data_in[5] ext_data_in[6] ext_data_in[7] ext_data_in[8] ext_data_in[9]
+ ext_data_in[10] ext_data_in[11] ext_data_in[12] ext_data_in[13] ext_data_in[14]
+ ext_data_in[15] ext_data_out[0] ext_data_out[1] ext_data_out[2] ext_data_out[3]
+ ext_data_out[4] ext_data_out[5] ext_data_out[6] ext_data_out[7] ext_data_out[8]
+ ext_data_out[9] ext_data_out[10] ext_data_out[11] ext_data_out[12] ext_data_out[13]
+ ext_data_out[14] ext_data_out[15] pe_busy[0] pe_busy[1] pe_busy[2] pe_busy[3]
XFILL_22_0_2 gnd vdd FILL
XFILL_5_1_2 gnd vdd FILL
XAND2X2_5 INVX2_6/A INVX4_1/A gnd AND2X2_5/Y vdd AND2X2
XOAI21X1_382 BUFX4_31/Y OR2X2_10/B INVX1_114/A gnd OAI21X1_383/C vdd OAI21X1
XOAI21X1_360 INVX1_99/Y OR2X2_9/Y OAI21X1_360/C gnd DFFSR_84/D vdd OAI21X1
XOAI21X1_371 DFFSR_90/Q INVX1_105/Y OAI21X1_371/C gnd DFFSR_78/D vdd OAI21X1
XFILL_13_0_2 gnd vdd FILL
XOAI21X1_393 BUFX4_61/Y BUFX2_24/A DFFSR_112/Q gnd OAI21X1_394/C vdd OAI21X1
XFILL_23_3_0 gnd vdd FILL
XMUX2X1_28 MUX2X1_42/A MUX2X1_28/B NOR2X1_13/Y gnd MUX2X1_28/Y vdd MUX2X1
XMUX2X1_17 MUX2X1_3/A INVX1_18/A NOR2X1_7/Y gnd MUX2X1_17/Y vdd MUX2X1
XMUX2X1_39 INVX1_45/A MUX2X1_39/B MUX2X1_39/S gnd MUX2X1_39/Y vdd MUX2X1
XFILL_14_3_0 gnd vdd FILL
XOAI21X1_190 BUFX4_62/Y BUFX4_16/Y MUX2X1_56/B gnd OAI21X1_191/C vdd OAI21X1
XDFFSR_9 DFFSR_9/Q DFFSR_9/CLK DFFSR_6/R vdd DFFSR_9/D gnd vdd DFFSR
XNAND2X1_43 MUX2X1_48/B NOR2X1_19/Y gnd NAND2X1_43/Y vdd NAND2X1
XNAND2X1_32 DFFSR_95/Q DFFSR_100/Q gnd NAND2X1_32/Y vdd NAND2X1
XNAND2X1_10 INVX1_4/A INVX1_5/Y gnd MUX2X1_9/S vdd NAND2X1
XNAND2X1_21 MUX2X1_25/B NOR2X1_9/Y gnd NAND2X1_21/Y vdd NAND2X1
XNAND2X1_98 NAND2X1_98/A NAND2X1_98/B gnd DFFSR_64/D vdd NAND2X1
XNAND2X1_65 NAND2X1_65/A NAND2X1_65/B gnd DFFSR_57/D vdd NAND2X1
XNAND2X1_87 DFFSR_123/Q DFFSR_127/Q gnd NAND2X1_87/Y vdd NAND2X1
XNAND2X1_54 NAND2X1_54/A NAND2X1_44/B gnd DFFSR_23/D vdd NAND2X1
XNAND2X1_76 NAND2X1_76/A NAND2X1_76/B gnd DFFSR_48/D vdd NAND2X1
XOAI22X1_3 OAI22X1_3/A OAI22X1_4/B INVX1_146/Y OAI22X1_4/D gnd OAI22X1_3/Y vdd OAI22X1
XFILL_20_1_0 gnd vdd FILL
XINVX2_12 INVX2_12/A gnd INVX2_12/Y vdd INVX2
XFILL_3_2_0 gnd vdd FILL
XOAI21X1_19 BUFX4_10/Y MUX2X1_6/Y OAI21X1_19/C gnd OAI21X1_19/Y vdd OAI21X1
XFILL_11_1_0 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XBUFX4_85 INVX8_4/Y gnd DFFSR_71/R vdd BUFX4
XBUFX4_74 DFFSR_1/Q gnd BUFX4_74/Y vdd BUFX4
XBUFX4_52 INVX8_1/Y gnd DFFSR_2/S vdd BUFX4
XBUFX4_41 NOR2X1_4/Y gnd BUFX4_41/Y vdd BUFX4
XBUFX4_30 INVX8_3/Y gnd DFFSR_43/R vdd BUFX4
XBUFX4_63 BUFX4_63/A gnd BUFX4_63/Y vdd BUFX4
XBUFX4_96 BUFX4_93/A gnd BUFX4_96/Y vdd BUFX4
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XOR2X2_11 BUFX4_63/Y BUFX2_24/A gnd OR2X2_11/Y vdd OR2X2
XXNOR2X1_6 NOR2X1_16/Y INVX2_2/Y gnd DFFSR_32/D vdd XNOR2X1
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XFILL_8_1_0 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XOAI21X1_383 INVX1_114/Y OR2X2_10/Y OAI21X1_383/C gnd DFFSR_101/D vdd OAI21X1
XOAI21X1_372 DFFSR_90/Q INVX1_106/Y OAI21X1_372/C gnd DFFSR_79/D vdd OAI21X1
XOAI21X1_361 OR2X2_9/A OR2X2_9/B DFFSR_85/Q gnd OAI21X1_362/C vdd OAI21X1
XOAI21X1_394 INVX1_123/Y OR2X2_11/Y OAI21X1_394/C gnd DFFSR_112/D vdd OAI21X1
XOAI21X1_350 OAI21X1_350/A OAI21X1_349/Y NOR2X1_36/Y gnd NAND2X1_108/B vdd OAI21X1
XFILL_23_3_1 gnd vdd FILL
XMUX2X1_18 MUX2X1_4/A INVX1_20/A NOR2X1_7/Y gnd MUX2X1_18/Y vdd MUX2X1
XMUX2X1_29 MUX2X1_49/A MUX2X1_29/B NOR2X1_13/Y gnd MUX2X1_29/Y vdd MUX2X1
XFILL_14_3_1 gnd vdd FILL
XOAI21X1_191 BUFX4_92/Y MUX2X1_56/Y OAI21X1_191/C gnd OAI21X1_191/Y vdd OAI21X1
XAOI22X1_1 INVX2_5/A AND2X2_5/Y BUFX2_4/Y NOR2X1_49/Y gnd AOI22X1_1/Y vdd AOI22X1
XOAI21X1_180 DFFSR_109/Q INVX1_51/Y NAND2X1_57/Y gnd MUX2X1_53/A vdd OAI21X1
XNAND2X1_66 DFFSR_54/Q INVX1_53/Y gnd MUX2X1_66/S vdd NAND2X1
XNAND2X1_33 DFFSR_95/Q INVX1_114/A gnd NAND2X1_33/Y vdd NAND2X1
XNAND2X1_44 NAND2X1_44/A NAND2X1_44/B gnd DFFSR_27/D vdd NAND2X1
XNAND2X1_11 DFFSR_14/Q INVX2_1/Y gnd OAI21X1_69/B vdd NAND2X1
XNAND2X1_55 NAND2X1_55/A NAND2X1_46/B gnd DFFSR_24/D vdd NAND2X1
XNAND2X1_22 NAND2X1_22/A OAI21X1_79/Y gnd DFFSR_11/D vdd NAND2X1
XNAND2X1_77 MUX2X1_77/B NOR2X1_29/Y gnd NAND2X1_77/Y vdd NAND2X1
XNAND2X1_99 NAND2X1_99/A NOR2X1_39/Y gnd NAND2X1_99/Y vdd NAND2X1
XNAND2X1_88 DFFSR_123/Q DFFSR_128/Q gnd NAND2X1_88/Y vdd NAND2X1
XOAI22X1_4 OAI22X1_4/A OAI22X1_4/B OAI22X1_3/A OAI22X1_4/D gnd OAI22X1_4/Y vdd OAI22X1
XFILL_20_1_1 gnd vdd FILL
XINVX2_13 INVX2_13/A gnd INVX2_13/Y vdd INVX2
XFILL_3_2_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_19_2_1 gnd vdd FILL
XBUFX4_20 DFFSR_58/Q gnd BUFX4_20/Y vdd BUFX4
XBUFX4_64 BUFX4_63/A gnd BUFX4_64/Y vdd BUFX4
XBUFX4_86 INVX8_4/Y gnd DFFSR_69/R vdd BUFX4
XBUFX4_42 NOR2X1_4/Y gnd BUFX4_42/Y vdd BUFX4
XBUFX4_53 INVX8_1/Y gnd DFFSR_5/R vdd BUFX4
XBUFX4_97 DFFSR_2/Q gnd BUFX4_97/Y vdd BUFX4
XBUFX4_75 DFFSR_1/Q gnd INVX1_2/A vdd BUFX4
XBUFX4_31 DFFSR_20/Q gnd BUFX4_31/Y vdd BUFX4
XOR2X2_12 OR2X2_12/A BUFX2_25/A gnd OR2X2_12/Y vdd OR2X2
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XXNOR2X1_7 BUFX4_93/Y DFFSR_53/Q gnd DFFSR_53/D vdd XNOR2X1
XFILL_0_0_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XFILL_8_1_1 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XOAI21X1_395 BUFX4_62/Y BUFX2_24/A DFFSR_113/Q gnd OAI21X1_395/Y vdd OAI21X1
XOAI21X1_351 INVX2_4/Y OR2X2_8/Y DFFSR_71/Q gnd OAI21X1_352/C vdd OAI21X1
XOAI21X1_384 BUFX4_31/Y OR2X2_10/B DFFSR_102/Q gnd OAI21X1_385/C vdd OAI21X1
XOAI21X1_373 DFFSR_90/Q INVX1_107/Y OAI21X1_373/C gnd DFFSR_80/D vdd OAI21X1
XOAI21X1_362 INVX1_100/Y OR2X2_9/Y OAI21X1_362/C gnd DFFSR_85/D vdd OAI21X1
XOAI21X1_340 INVX1_91/Y NAND2X1_95/Y NAND3X1_26/Y gnd OAI21X1_342/A vdd OAI21X1
XFILL_23_3_2 gnd vdd FILL
XMUX2X1_19 MUX2X1_5/A INVX1_22/A NOR2X1_7/Y gnd MUX2X1_19/Y vdd MUX2X1
XFILL_14_3_2 gnd vdd FILL
XAOI22X1_2 DFFSR_68/Q AND2X2_5/Y DFFSR_30/Q NOR2X1_48/Y gnd AOI22X1_2/Y vdd AOI22X1
XOAI21X1_181 BUFX4_62/Y BUFX4_15/Y MUX2X1_53/B gnd OAI21X1_181/Y vdd OAI21X1
XOAI21X1_170 INVX1_47/Y NAND2X1_39/Y NAND3X1_14/Y gnd OAI21X1_170/Y vdd OAI21X1
XOAI21X1_192 DFFSR_109/Q INVX1_57/Y NAND2X1_61/Y gnd MUX2X1_71/A vdd OAI21X1
XNAND2X1_89 DFFSR_123/Q INVX1_138/A gnd NAND2X1_89/Y vdd NAND2X1
XNAND2X1_34 DFFSR_95/Q DFFSR_102/Q gnd NAND2X1_34/Y vdd NAND2X1
XNAND2X1_56 NAND2X1_56/A NAND2X1_56/B gnd DFFSR_25/D vdd NAND2X1
XNAND2X1_12 MUX2X1_21/B NOR2X1_9/Y gnd NAND2X1_12/Y vdd NAND2X1
XNAND2X1_23 MUX2X1_26/B NOR2X1_9/Y gnd NAND2X1_23/Y vdd NAND2X1
XNAND2X1_45 MUX2X1_49/B NOR2X1_19/Y gnd NAND2X1_45/Y vdd NAND2X1
XNAND2X1_67 DFFSR_52/Q INVX2_3/Y gnd NAND2X1_67/Y vdd NAND2X1
XNAND2X1_78 NAND2X1_78/A NAND2X1_78/B gnd DFFSR_49/D vdd NAND2X1
XAOI22X1_10 DFFSR_49/Q AND2X2_5/Y DFFSR_30/Q NOR2X1_49/Y gnd AOI22X1_10/Y vdd AOI22X1
XOAI22X1_5 OAI22X1_1/Y NOR2X1_42/B OAI22X1_3/Y NOR2X1_45/B gnd NOR2X1_52/A vdd OAI22X1
XFILL_20_1_2 gnd vdd FILL
XFILL_3_2_2 gnd vdd FILL
XFILL_11_1_2 gnd vdd FILL
XFILL_19_2_2 gnd vdd FILL
XINVX8_1 rst gnd INVX8_1/Y vdd INVX8
XBUFX4_21 DFFSR_58/Q gnd BUFX4_21/Y vdd BUFX4
XBUFX4_32 DFFSR_20/Q gnd BUFX4_32/Y vdd BUFX4
XBUFX4_43 NOR2X1_4/Y gnd BUFX4_43/Y vdd BUFX4
XBUFX4_10 BUFX4_13/A gnd BUFX4_10/Y vdd BUFX4
XBUFX4_87 INVX8_4/Y gnd DFFSR_74/R vdd BUFX4
XBUFX4_65 BUFX4_63/A gnd BUFX4_65/Y vdd BUFX4
XBUFX4_76 DFFSR_1/Q gnd BUFX4_76/Y vdd BUFX4
XBUFX4_54 BUFX4_57/A gnd BUFX4_54/Y vdd BUFX4
XBUFX4_98 DFFSR_2/Q gnd INVX2_5/A vdd BUFX4
XXNOR2X1_8 NOR2X1_30/Y INVX1_52/Y gnd DFFSR_54/D vdd XNOR2X1
XOR2X2_13 BUFX2_26/A gnd gnd OR2X2_13/Y vdd OR2X2
XOR2X2_6 OR2X2_6/A OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XFILL_0_0_2 gnd vdd FILL
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_8_1_2 gnd vdd FILL
XFILL_16_0_2 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XOAI21X1_330 OAI21X1_328/Y OAI21X1_329/Y NOR2X1_36/Y gnd NAND2X1_98/B vdd OAI21X1
XOAI21X1_341 INVX1_92/Y NAND2X1_97/Y OAI21X1_341/C gnd OAI21X1_341/Y vdd OAI21X1
XOAI21X1_396 INVX1_124/Y OR2X2_11/Y OAI21X1_395/Y gnd DFFSR_113/D vdd OAI21X1
XOAI21X1_385 INVX1_115/Y OR2X2_10/Y OAI21X1_385/C gnd DFFSR_102/D vdd OAI21X1
XOAI21X1_374 BUFX4_35/Y OR2X2_10/B DFFSR_97/Q gnd OAI21X1_375/C vdd OAI21X1
XOAI21X1_352 OR2X2_8/Y NAND2X1_97/Y OAI21X1_352/C gnd DFFSR_71/D vdd OAI21X1
XOAI21X1_363 BUFX4_74/Y OR2X2_9/B DFFSR_86/Q gnd OAI21X1_363/Y vdd OAI21X1
XFILL_17_3_0 gnd vdd FILL
XOAI21X1_182 BUFX4_92/Y MUX2X1_53/Y OAI21X1_181/Y gnd OAI21X1_182/Y vdd OAI21X1
XOAI21X1_160 OAI21X1_158/Y OAI21X1_160/B NOR2X1_16/Y gnd NAND2X1_46/B vdd OAI21X1
XOAI21X1_171 INVX1_48/Y NAND2X1_41/Y NAND2X1_51/Y gnd OAI21X1_172/B vdd OAI21X1
XAOI22X1_3 DFFSR_11/Q AOI21X1_9/A DFFSR_49/Q NOR2X1_49/Y gnd AOI22X1_3/Y vdd AOI22X1
XOAI21X1_193 BUFX4_61/Y BUFX4_15/Y MUX2X1_57/B gnd OAI21X1_193/Y vdd OAI21X1
XNAND2X1_57 DFFSR_109/Q DFFSR_111/Q gnd NAND2X1_57/Y vdd NAND2X1
XNAND2X1_13 INVX2_1/A INVX1_14/Y gnd OAI21X1_78/B vdd NAND2X1
XNAND2X1_24 NAND2X1_24/A OAI21X1_83/Y gnd DFFSR_12/D vdd NAND2X1
XNAND2X1_46 NAND2X1_46/A NAND2X1_46/B gnd DFFSR_28/D vdd NAND2X1
XNAND2X1_35 OR2X2_3/A OR2X2_3/B gnd NAND2X1_36/B vdd NAND2X1
XNAND2X1_68 MUX2X1_73/B NOR2X1_29/Y gnd NAND2X1_68/Y vdd NAND2X1
XNAND2X1_79 MUX2X1_78/B NOR2X1_29/Y gnd NAND2X1_79/Y vdd NAND2X1
XAOI22X1_11 AOI21X1_9/A DFFSR_12/Q DFFSR_69/Q AND2X2_5/Y gnd NAND3X1_45/A vdd AOI22X1
XFILL_23_1_0 gnd vdd FILL
XOAI22X1_6 OAI22X1_6/A OAI22X1_6/B INVX4_3/Y OAI22X1_6/D gnd OAI22X1_6/Y vdd OAI22X1
XFILL_6_2_0 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XFILL_3_0_0 gnd vdd FILL
XINVX8_2 rst gnd INVX8_2/Y vdd INVX8
XBUFX4_55 BUFX4_57/A gnd BUFX4_55/Y vdd BUFX4
XBUFX4_11 BUFX4_13/A gnd BUFX4_11/Y vdd BUFX4
XBUFX4_44 NOR2X1_4/Y gnd BUFX4_44/Y vdd BUFX4
XBUFX4_33 DFFSR_20/Q gnd BUFX4_33/Y vdd BUFX4
XBUFX4_77 INVX8_2/Y gnd DFFSR_38/R vdd BUFX4
XBUFX4_66 INVX8_9/Y gnd BUFX4_66/Y vdd BUFX4
XBUFX4_22 DFFSR_58/Q gnd BUFX4_22/Y vdd BUFX4
XBUFX4_88 INVX8_4/Y gnd BUFX4_88/Y vdd BUFX4
XBUFX4_99 DFFSR_2/Q gnd OR2X2_2/B vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XOR2X2_14 BUFX2_1/Y gnd gnd OR2X2_14/Y vdd OR2X2
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XXNOR2X1_9 NOR2X1_26/Y INVX2_3/Y gnd DFFSR_51/D vdd XNOR2X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XFILL_1_3_1 gnd vdd FILL
XOAI21X1_353 BUFX4_89/Y OR2X2_8/A DFFSR_60/Q gnd NAND2X1_109/A vdd OAI21X1
XOAI21X1_364 INVX1_101/Y OR2X2_9/Y OAI21X1_363/Y gnd DFFSR_86/D vdd OAI21X1
XOAI21X1_320 BUFX4_47/Y MUX2X1_101/Y OAI21X1_319/Y gnd DFFPOSX1_75/D vdd OAI21X1
XOAI21X1_342 OAI21X1_342/A OAI21X1_341/Y NOR2X1_36/Y gnd NAND2X1_112/B vdd OAI21X1
XOAI21X1_331 BUFX4_91/Y OR2X2_8/A DFFSR_65/Q gnd OAI21X1_331/Y vdd OAI21X1
XOAI21X1_397 BUFX4_65/Y BUFX2_24/A DFFSR_114/Q gnd OAI21X1_397/Y vdd OAI21X1
XOAI21X1_386 BUFX4_35/Y DFFSR_95/Q OAI21X1_386/C gnd DFFSR_103/D vdd OAI21X1
XOAI21X1_375 INVX1_110/Y OR2X2_10/Y OAI21X1_375/C gnd DFFSR_97/D vdd OAI21X1
XFILL_17_3_1 gnd vdd FILL
XOAI21X1_194 BUFX4_92/Y MUX2X1_57/Y OAI21X1_193/Y gnd DFFPOSX1_71/D vdd OAI21X1
XOAI21X1_150 INVX1_36/Y NAND2X1_39/Y NAND3X1_9/Y gnd OAI21X1_150/Y vdd OAI21X1
XOAI21X1_161 BUFX2_3/Y OR2X2_4/A DFFSR_29/Q gnd NAND2X1_48/A vdd OAI21X1
XOAI21X1_172 OAI21X1_170/Y OAI21X1_172/B NOR2X1_16/Y gnd NAND2X1_52/B vdd OAI21X1
XOAI21X1_183 DFFSR_109/Q INVX1_54/Y NAND2X1_58/Y gnd MUX2X1_68/A vdd OAI21X1
XAOI22X1_4 DFFSR_11/Q AND2X2_5/Y DFFSR_68/Q NOR2X1_49/Y gnd AOI22X1_4/Y vdd AOI22X1
XNAND2X1_25 OAI21X1_86/Y NAND2X1_14/B gnd DFFSR_3/D vdd NAND2X1
XNAND2X1_14 OAI21X1_60/Y NAND2X1_14/B gnd DFFSR_7/D vdd NAND2X1
XNAND2X1_47 MUX2X1_50/B NOR2X1_19/Y gnd NAND2X1_47/Y vdd NAND2X1
XNAND2X1_36 INVX1_25/A NAND2X1_36/B gnd AOI21X1_2/A vdd NAND2X1
XNAND2X1_58 DFFSR_109/Q DFFSR_112/Q gnd NAND2X1_58/Y vdd NAND2X1
XNAND2X1_69 INVX2_3/A INVX1_62/Y gnd NAND2X1_69/Y vdd NAND2X1
XAOI22X1_12 DFFSR_12/Q AND2X2_5/Y DFFSR_50/Q NOR2X1_48/Y gnd AOI22X1_12/Y vdd AOI22X1
XFILL_23_1_1 gnd vdd FILL
XOAI22X1_7 OAI22X1_6/A OAI22X1_7/B INVX4_3/Y OAI22X1_7/D gnd DFFSR_140/D vdd OAI22X1
XFILL_6_2_1 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XCLKBUF1_1 BUFX4_4/Y gnd DFFSR_9/CLK vdd CLKBUF1
XFILL_3_0_1 gnd vdd FILL
XINVX8_3 rst gnd INVX8_3/Y vdd INVX8
XBUFX4_23 DFFSR_58/Q gnd OR2X2_12/A vdd BUFX4
XBUFX4_89 BUFX2_4/A gnd BUFX4_89/Y vdd BUFX4
XBUFX4_12 BUFX4_13/A gnd AND2X2_1/A vdd BUFX4
XBUFX4_78 INVX8_2/Y gnd BUFX4_78/Y vdd BUFX4
XBUFX4_56 BUFX4_57/A gnd BUFX4_56/Y vdd BUFX4
XBUFX4_34 DFFSR_20/Q gnd BUFX4_34/Y vdd BUFX4
XBUFX4_67 INVX8_9/Y gnd BUFX4_67/Y vdd BUFX4
XBUFX4_45 BUFX4_48/A gnd BUFX4_45/Y vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XFILL_1_3_2 gnd vdd FILL
XOAI21X1_398 INVX1_125/Y OR2X2_11/Y OAI21X1_397/Y gnd DFFSR_114/D vdd OAI21X1
XOAI21X1_354 BUFX4_89/Y OR2X2_8/A DFFSR_61/Q gnd NAND2X1_110/A vdd OAI21X1
XOAI21X1_310 BUFX4_47/Y MUX2X1_96/Y OAI21X1_309/Y gnd DFFPOSX1_82/D vdd OAI21X1
XOAI21X1_376 BUFX4_35/Y OR2X2_10/B DFFSR_98/Q gnd OAI21X1_377/C vdd OAI21X1
XOAI21X1_387 DFFSR_104/Q INVX1_116/Y OAI21X1_387/C gnd DFFSR_91/D vdd OAI21X1
XOAI21X1_365 OR2X2_9/A OR2X2_9/B DFFSR_87/Q gnd OAI21X1_365/Y vdd OAI21X1
XOAI21X1_321 BUFX4_22/Y BUFX4_84/Y MUX2X1_102/B gnd OAI21X1_321/Y vdd OAI21X1
XOAI21X1_332 INVX1_87/Y NAND2X1_95/Y NAND3X1_24/Y gnd OAI21X1_332/Y vdd OAI21X1
XOAI21X1_343 BUFX4_91/Y OR2X2_8/A DFFSR_68/Q gnd NAND2X1_106/A vdd OAI21X1
XFILL_17_3_2 gnd vdd FILL
XOAI21X1_162 INVX1_43/Y NAND2X1_39/Y NAND3X1_12/Y gnd OAI21X1_162/Y vdd OAI21X1
XOAI21X1_140 BUFX4_40/Y MUX2X1_48/Y OAI21X1_139/Y gnd OAI21X1_140/Y vdd OAI21X1
XOAI21X1_151 INVX1_37/Y NAND2X1_41/Y NAND2X1_40/Y gnd OAI21X1_152/B vdd OAI21X1
XOAI21X1_173 INVX2_2/Y OR2X2_4/Y DFFSR_33/Q gnd OAI21X1_174/C vdd OAI21X1
XOAI21X1_195 DFFSR_109/Q INVX1_58/Y NAND2X1_62/Y gnd MUX2X1_66/B vdd OAI21X1
XOAI21X1_184 BUFX4_61/Y BUFX4_15/Y MUX2X1_54/B gnd OAI21X1_185/C vdd OAI21X1
XAOI22X1_5 AOI22X1_5/A AOI22X1_5/B AOI22X1_5/C AOI21X1_7/C gnd AOI22X1_5/Y vdd AOI22X1
XNAND2X1_59 DFFSR_109/Q DFFSR_113/Q gnd NAND2X1_59/Y vdd NAND2X1
XNAND2X1_48 NAND2X1_48/A NAND2X1_56/B gnd DFFSR_29/D vdd NAND2X1
XNAND2X1_15 MUX2X1_22/B NOR2X1_9/Y gnd NAND2X1_15/Y vdd NAND2X1
XNAND2X1_26 OAI21X1_87/Y NAND2X1_16/B gnd DFFSR_4/D vdd NAND2X1
XNAND2X1_37 NAND2X1_37/A NAND2X1_37/B gnd DFFSR_38/D vdd NAND2X1
XAOI22X1_13 AOI22X1_5/A AOI22X1_5/B NAND3X1_48/Y AOI21X1_7/C gnd NAND3X1_49/C vdd
+ AOI22X1
XFILL_23_1_2 gnd vdd FILL
XOAI22X1_8 INVX4_3/Y OAI22X1_8/B OR2X2_14/Y OAI22X1_6/A gnd DFFSR_178/D vdd OAI22X1
XFILL_6_2_2 gnd vdd FILL
XFILL_14_1_2 gnd vdd FILL
XFILL_19_1 gnd vdd FILL
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B MUX2X1_5/S gnd MUX2X1_1/Y vdd MUX2X1
XCLKBUF1_2 BUFX4_4/Y gnd DFFSR_8/CLK vdd CLKBUF1
XFILL_3_0_2 gnd vdd FILL
XINVX8_4 rst gnd INVX8_4/Y vdd INVX8
XDFFPOSX1_90 INVX1_95/A CLKBUF1_7/Y OAI21X1_302/Y gnd vdd DFFPOSX1
XBUFX4_35 DFFSR_20/Q gnd BUFX4_35/Y vdd BUFX4
XBUFX4_79 INVX8_2/Y gnd DFFSR_29/R vdd BUFX4
XBUFX4_13 BUFX4_13/A gnd MUX2X1_7/S vdd BUFX4
XBUFX4_57 BUFX4_57/A gnd BUFX4_57/Y vdd BUFX4
XBUFX4_68 INVX8_9/Y gnd BUFX4_68/Y vdd BUFX4
XBUFX4_46 BUFX4_48/A gnd BUFX4_46/Y vdd BUFX4
XBUFX4_24 BUFX2_2/A gnd OR2X2_6/B vdd BUFX4
XFILL_19_0_2 gnd vdd FILL
XOR2X2_9 OR2X2_9/A OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XFILL_21_2_0 gnd vdd FILL
XFILL_4_3_0 gnd vdd FILL
XFILL_12_2_0 gnd vdd FILL
XOAI21X1_355 OR2X2_8/B OR2X2_8/A DFFSR_62/Q gnd NAND2X1_111/A vdd OAI21X1
XOAI21X1_377 INVX1_111/Y OR2X2_10/Y OAI21X1_377/C gnd DFFSR_98/D vdd OAI21X1
XOAI21X1_388 DFFSR_104/Q INVX1_117/Y OAI21X1_388/C gnd DFFSR_92/D vdd OAI21X1
XOAI21X1_366 INVX1_102/Y OR2X2_9/Y OAI21X1_365/Y gnd DFFSR_87/D vdd OAI21X1
XOAI21X1_322 BUFX4_47/Y MUX2X1_102/Y OAI21X1_321/Y gnd OAI21X1_322/Y vdd OAI21X1
XOAI21X1_399 BUFX4_61/Y BUFX2_24/A INVX1_126/A gnd OAI21X1_399/Y vdd OAI21X1
XOAI21X1_333 INVX1_88/Y NAND2X1_97/Y NAND2X1_99/Y gnd OAI21X1_333/Y vdd OAI21X1
XOAI21X1_300 BUFX4_46/Y MUX2X1_91/Y OAI21X1_300/C gnd OAI21X1_300/Y vdd OAI21X1
XOAI21X1_344 INVX1_93/Y NAND2X1_95/Y NAND3X1_27/Y gnd OAI21X1_344/Y vdd OAI21X1
XOAI21X1_311 OR2X2_12/A BUFX4_82/Y INVX1_94/A gnd OAI21X1_311/Y vdd OAI21X1
XNAND3X1_1 OR2X2_1/A OR2X2_1/B INVX1_1/Y gnd AOI21X1_1/B vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XOAI21X1_130 BUFX4_37/Y MUX2X1_43/Y OAI21X1_130/C gnd DFFPOSX1_33/D vdd OAI21X1
XOAI21X1_196 BUFX4_62/Y BUFX4_15/Y MUX2X1_58/B gnd OAI21X1_197/C vdd OAI21X1
XOAI21X1_163 INVX1_44/Y NAND2X1_41/Y NAND2X1_47/Y gnd OAI21X1_164/B vdd OAI21X1
XOAI21X1_152 OAI21X1_150/Y OAI21X1_152/B NOR2X1_16/Y gnd NAND2X1_42/B vdd OAI21X1
XOAI21X1_141 BUFX4_34/Y BUFX4_57/Y MUX2X1_49/B gnd OAI21X1_142/C vdd OAI21X1
XOAI21X1_174 OR2X2_4/Y NAND2X1_41/Y OAI21X1_174/C gnd DFFSR_33/D vdd OAI21X1
XOAI21X1_185 BUFX4_94/Y MUX2X1_54/Y OAI21X1_185/C gnd DFFPOSX1_68/D vdd OAI21X1
XAOI22X1_6 DFFSR_49/Q AOI21X1_9/A DFFSR_11/Q NOR2X1_49/Y gnd AOI22X1_6/Y vdd AOI22X1
XNAND2X1_27 OAI21X1_88/Y NAND2X1_18/B gnd DFFSR_5/D vdd NAND2X1
XNAND2X1_16 NAND2X1_16/A NAND2X1_16/B gnd DFFSR_8/D vdd NAND2X1
XNAND2X1_49 MUX2X1_51/B NOR2X1_19/Y gnd NAND2X1_49/Y vdd NAND2X1
XNAND2X1_38 INVX1_28/A INVX1_29/Y gnd MUX2X1_39/S vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XNAND2X1_180 NAND2X1_179/Y NAND2X1_180/B gnd DFFSR_176/D vdd NAND2X1
XFILL_17_1_0 gnd vdd FILL
XAOI22X1_14 AOI21X1_9/A DFFSR_50/Q DFFSR_31/Q AND2X2_5/Y gnd NAND3X1_50/A vdd AOI22X1
XOAI22X1_9 OAI22X1_6/A OAI22X1_9/B INVX4_3/Y OAI22X1_9/D gnd DFFSR_141/D vdd OAI22X1
XXOR2X1_1 XOR2X1_1/A OR2X2_1/B gnd DFFSR_17/D vdd XOR2X1
XFILL_6_0_0 gnd vdd FILL
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B MUX2X1_5/S gnd MUX2X1_2/Y vdd MUX2X1
XCLKBUF1_3 BUFX4_1/Y gnd CLKBUF1_3/Y vdd CLKBUF1
XINVX8_5 rst gnd INVX8_5/Y vdd INVX8
XDFFPOSX1_91 MUX2X1_79/B CLKBUF1_7/Y OAI21X1_271/Y gnd vdd DFFPOSX1
XBUFX4_14 BUFX4_13/A gnd BUFX4_14/Y vdd BUFX4
XDFFPOSX1_80 INVX1_88/A CLKBUF1_7/Y OAI21X1_306/Y gnd vdd DFFPOSX1
XBUFX4_25 BUFX2_2/A gnd BUFX4_25/Y vdd BUFX4
XBUFX4_36 BUFX4_36/A gnd BUFX4_36/Y vdd BUFX4
XBUFX4_58 BUFX2_3/A gnd BUFX4_58/Y vdd BUFX4
XBUFX4_69 INVX8_9/Y gnd BUFX4_69/Y vdd BUFX4
XBUFX4_47 BUFX4_48/A gnd BUFX4_47/Y vdd BUFX4
XFILL_21_2_1 gnd vdd FILL
XFILL_4_3_1 gnd vdd FILL
XFILL_12_2_1 gnd vdd FILL
XOAI21X1_323 BUFX4_20/Y BUFX4_82/Y MUX2X1_103/B gnd OAI21X1_324/C vdd OAI21X1
XOAI21X1_301 BUFX4_20/Y BUFX4_82/Y INVX1_95/A gnd OAI21X1_301/Y vdd OAI21X1
XOAI21X1_312 BUFX4_45/Y MUX2X1_97/Y OAI21X1_311/Y gnd DFFPOSX1_83/D vdd OAI21X1
XOAI21X1_356 OR2X2_8/B OR2X2_8/A DFFSR_63/Q gnd NAND2X1_112/A vdd OAI21X1
XOAI21X1_389 DFFSR_104/Q INVX1_118/Y OAI21X1_389/C gnd DFFSR_93/D vdd OAI21X1
XOAI21X1_378 BUFX4_31/Y OR2X2_10/B DFFSR_99/Q gnd OAI21X1_379/C vdd OAI21X1
XOAI21X1_367 OR2X2_9/A OR2X2_9/B DFFSR_88/Q gnd OAI21X1_368/C vdd OAI21X1
XOAI21X1_334 OAI21X1_332/Y OAI21X1_333/Y NOR2X1_36/Y gnd NAND2X1_110/B vdd OAI21X1
XOAI21X1_345 INVX1_94/Y NAND2X1_97/Y OAI21X1_345/C gnd OAI21X1_345/Y vdd OAI21X1
XNAND3X1_2 MUX2X1_1/B DFFSR_14/Q INVX2_1/A gnd NAND3X1_2/Y vdd NAND3X1
XFILL_1_1_1 gnd vdd FILL
XOAI21X1_131 BUFX4_34/Y BUFX4_57/Y INVX1_44/A gnd OAI21X1_132/C vdd OAI21X1
XOAI21X1_164 OAI21X1_162/Y OAI21X1_164/B NOR2X1_16/Y gnd NAND2X1_56/B vdd OAI21X1
XOAI21X1_153 BUFX4_59/Y OR2X2_4/A DFFSR_27/Q gnd NAND2X1_44/A vdd OAI21X1
XOAI21X1_120 BUFX4_40/Y MUX2X1_38/Y OAI21X1_119/Y gnd DFFPOSX1_40/D vdd OAI21X1
XOAI21X1_142 BUFX4_40/Y MUX2X1_49/Y OAI21X1_142/C gnd OAI21X1_142/Y vdd OAI21X1
XAOI22X1_7 DFFSR_30/Q AND2X2_5/Y DFFSR_68/Q NOR2X1_48/Y gnd AOI22X1_7/Y vdd AOI22X1
XOAI21X1_197 BUFX4_92/Y MUX2X1_58/Y OAI21X1_197/C gnd OAI21X1_197/Y vdd OAI21X1
XOAI21X1_175 BUFX2_3/Y OR2X2_4/A DFFSR_22/Q gnd NAND2X1_53/A vdd OAI21X1
XFILL_9_2_1 gnd vdd FILL
XOAI21X1_186 DFFSR_109/Q INVX1_55/Y NAND2X1_59/Y gnd MUX2X1_55/A vdd OAI21X1
XNAND2X1_28 NAND2X1_28/A NAND2X1_20/B gnd DFFSR_6/D vdd NAND2X1
XNAND2X1_17 MUX2X1_23/B NOR2X1_9/Y gnd NAND2X1_17/Y vdd NAND2X1
XNAND2X1_39 DFFSR_33/Q INVX2_2/Y gnd NAND2X1_39/Y vdd NAND2X1
XNAND2X1_170 INVX2_9/A INVX4_3/Y gnd NAND2X1_171/A vdd NAND2X1
XNAND2X1_181 NAND3X1_71/Y NAND3X1_70/Y gnd OAI21X1_463/A vdd NAND2X1
XFILL_17_1_1 gnd vdd FILL
XAOI22X1_15 NOR2X1_48/Y DFFSR_69/Q DFFSR_12/Q NOR2X1_49/Y gnd NAND3X1_50/B vdd AOI22X1
XFILL_6_0_1 gnd vdd FILL
XXOR2X1_2 OR2X2_1/A OR2X2_1/B gnd XOR2X1_2/Y vdd XOR2X1
XMUX2X1_3 MUX2X1_3/A MUX2X1_3/B MUX2X1_5/S gnd MUX2X1_3/Y vdd MUX2X1
XCLKBUF1_4 BUFX4_4/Y gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_24_1 gnd vdd FILL
XINVX8_6 rst gnd INVX8_6/Y vdd INVX8
XDFFPOSX1_70 MUX2X1_56/B CLKBUF1_21/Y OAI21X1_191/Y gnd vdd DFFPOSX1
XDFFPOSX1_81 INVX1_90/A CLKBUF1_25/Y OAI21X1_308/Y gnd vdd DFFPOSX1
XBUFX4_37 BUFX4_36/A gnd BUFX4_37/Y vdd BUFX4
XBUFX4_59 BUFX2_3/A gnd BUFX4_59/Y vdd BUFX4
XDFFPOSX1_92 MUX2X1_80/B CLKBUF1_25/Y OAI21X1_274/Y gnd vdd DFFPOSX1
XBUFX4_26 BUFX2_2/A gnd BUFX4_26/Y vdd BUFX4
XBUFX4_15 BUFX4_18/A gnd BUFX4_15/Y vdd BUFX4
XBUFX4_48 BUFX4_48/A gnd AND2X2_4/A vdd BUFX4
XFILL_21_2_2 gnd vdd FILL
XFILL_4_3_2 gnd vdd FILL
XFILL_12_2_2 gnd vdd FILL
XOAI21X1_313 BUFX4_22/Y BUFX4_84/Y INVX1_96/A gnd OAI21X1_313/Y vdd OAI21X1
XOAI21X1_335 BUFX4_91/Y OR2X2_8/A DFFSR_66/Q gnd OAI21X1_335/Y vdd OAI21X1
XOAI21X1_324 BUFX4_45/Y MUX2X1_103/Y OAI21X1_324/C gnd DFFPOSX1_77/D vdd OAI21X1
XOAI21X1_302 BUFX4_49/Y MUX2X1_92/Y OAI21X1_301/Y gnd OAI21X1_302/Y vdd OAI21X1
XOAI21X1_346 OAI21X1_344/Y OAI21X1_345/Y NOR2X1_36/Y gnd NAND2X1_106/B vdd OAI21X1
XOAI21X1_379 INVX1_112/Y OR2X2_10/Y OAI21X1_379/C gnd DFFSR_99/D vdd OAI21X1
XOAI21X1_368 INVX1_103/Y OR2X2_9/Y OAI21X1_368/C gnd DFFSR_88/D vdd OAI21X1
XOAI21X1_357 OR2X2_9/A OR2X2_9/B DFFSR_83/Q gnd OAI21X1_357/Y vdd OAI21X1
XDFFSR_170 INVX1_82/A DFFSR_21/CLK BUFX4_70/Y vdd DFFSR_170/D gnd vdd DFFSR
XNAND3X1_3 MUX2X1_2/B DFFSR_14/Q INVX2_1/A gnd NAND3X1_3/Y vdd NAND3X1
XFILL_1_1_2 gnd vdd FILL
XOAI21X1_187 BUFX4_64/Y BUFX4_18/Y MUX2X1_55/B gnd OAI21X1_187/Y vdd OAI21X1
XOAI21X1_132 BUFX4_37/Y MUX2X1_44/Y OAI21X1_132/C gnd DFFPOSX1_34/D vdd OAI21X1
XOAI21X1_176 BUFX4_59/Y OR2X2_4/A DFFSR_23/Q gnd NAND2X1_54/A vdd OAI21X1
XOAI21X1_154 INVX1_39/Y NAND2X1_39/Y NAND3X1_10/Y gnd OAI21X1_154/Y vdd OAI21X1
XOAI21X1_143 BUFX4_35/Y BUFX4_56/Y MUX2X1_50/B gnd OAI21X1_143/Y vdd OAI21X1
XOAI21X1_165 BUFX4_59/Y OR2X2_4/A DFFSR_30/Q gnd NAND2X1_50/A vdd OAI21X1
XOAI21X1_121 BUFX4_33/Y BUFX4_54/Y INVX1_45/A gnd OAI21X1_121/Y vdd OAI21X1
XOAI21X1_110 AND2X2_2/Y AOI21X1_2/Y OR2X2_4/Y gnd NAND2X1_37/B vdd OAI21X1
XOAI21X1_198 OR2X2_6/B OR2X2_6/A AND2X2_3/A gnd XOR2X1_5/A vdd OAI21X1
XAOI22X1_8 AOI22X1_8/A INVX1_152/Y AOI22X1_8/C AOI22X1_8/D gnd AOI22X1_8/Y vdd AOI22X1
XFILL_9_2_2 gnd vdd FILL
XNAND2X1_18 NAND2X1_18/A NAND2X1_18/B gnd DFFSR_9/D vdd NAND2X1
XNAND2X1_29 DFFSR_95/Q DFFSR_97/Q gnd NAND2X1_29/Y vdd NAND2X1
XNAND2X1_171 NAND2X1_171/A NAND2X1_171/B gnd DFFSR_173/D vdd NAND2X1
XNAND2X1_182 INVX2_13/A INVX4_3/Y gnd NAND2X1_182/Y vdd NAND2X1
XNAND2X1_160 INVX2_7/A INVX4_3/Y gnd OAI22X1_6/A vdd NAND2X1
XFILL_17_1_2 gnd vdd FILL
XAOI22X1_16 AOI22X1_8/A INVX1_152/Y NAND3X1_50/Y AOI22X1_16/D gnd AOI22X1_16/Y vdd
+ AOI22X1
XFILL_10_3_0 gnd vdd FILL
XFILL_6_0_2 gnd vdd FILL
XXOR2X1_3 XOR2X1_3/A OR2X2_3/B gnd XOR2X1_3/Y vdd XOR2X1
XMUX2X1_4 MUX2X1_4/A MUX2X1_4/B MUX2X1_5/S gnd MUX2X1_4/Y vdd MUX2X1
XCLKBUF1_5 BUFX4_5/Y gnd CLKBUF1_5/Y vdd CLKBUF1
XFILL_24_2 gnd vdd FILL
XFILL_24_2_0 gnd vdd FILL
XINVX8_7 rst gnd INVX8_7/Y vdd INVX8
XDFFPOSX1_60 INVX1_72/A CLKBUF1_21/Y OAI21X1_225/Y gnd vdd DFFPOSX1
XDFFPOSX1_71 MUX2X1_57/B CLKBUF1_41/Y DFFPOSX1_71/D gnd vdd DFFPOSX1
XDFFPOSX1_93 MUX2X1_81/B CLKBUF1_25/Y DFFPOSX1_93/D gnd vdd DFFPOSX1
XDFFPOSX1_82 INVX1_92/A CLKBUF1_7/Y DFFPOSX1_82/D gnd vdd DFFPOSX1
XBUFX4_16 BUFX4_18/A gnd BUFX4_16/Y vdd BUFX4
XBUFX4_38 BUFX4_36/A gnd BUFX4_38/Y vdd BUFX4
XFILL_7_3_0 gnd vdd FILL
XBUFX4_49 BUFX4_48/A gnd BUFX4_49/Y vdd BUFX4
XBUFX4_27 INVX8_3/Y gnd DFFSR_54/R vdd BUFX4
XFILL_15_2_0 gnd vdd FILL
XFILL_21_0_0 gnd vdd FILL
XOAI21X1_369 BUFX4_76/Y NOR2X1_4/B OAI21X1_369/C gnd DFFSR_89/D vdd OAI21X1
XOAI21X1_358 INVX1_98/Y OR2X2_9/Y OAI21X1_357/Y gnd DFFSR_83/D vdd OAI21X1
XOAI21X1_314 BUFX4_47/Y MUX2X1_98/Y OAI21X1_313/Y gnd DFFPOSX1_84/D vdd OAI21X1
XOAI21X1_325 BUFX4_22/Y BUFX4_84/Y MUX2X1_104/B gnd OAI21X1_326/C vdd OAI21X1
XOAI21X1_336 INVX1_89/Y NAND2X1_95/Y NAND3X1_25/Y gnd OAI21X1_336/Y vdd OAI21X1
XOAI21X1_347 BUFX4_91/Y OR2X2_8/A DFFSR_69/Q gnd OAI21X1_347/Y vdd OAI21X1
XOAI21X1_303 BUFX4_20/Y BUFX4_82/Y INVX1_85/A gnd OAI21X1_304/C vdd OAI21X1
XDFFSR_171 INVX4_3/A CLKBUF1_12/Y BUFX4_66/Y vdd DFFSR_171/D gnd vdd DFFSR
XDFFSR_160 INVX1_54/A DFFSR_87/CLK BUFX4_68/Y vdd DFFSR_160/D gnd vdd DFFSR
XBUFX4_1 clk gnd BUFX4_1/Y vdd BUFX4
XFILL_4_1_0 gnd vdd FILL
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XFILL_12_0_0 gnd vdd FILL
XNAND3X1_4 MUX2X1_3/B DFFSR_14/Q INVX2_1/A gnd NAND3X1_4/Y vdd NAND3X1
XOAI21X1_199 AND2X2_3/Y AOI21X1_3/Y OR2X2_6/Y gnd NAND2X1_65/B vdd OAI21X1
XOAI21X1_188 AND2X2_3/A MUX2X1_55/Y OAI21X1_187/Y gnd OAI21X1_188/Y vdd OAI21X1
XOAI21X1_155 INVX1_40/Y NAND2X1_41/Y NAND2X1_43/Y gnd OAI21X1_156/B vdd OAI21X1
XOAI21X1_177 BUFX2_3/Y OR2X2_4/A DFFSR_24/Q gnd NAND2X1_55/A vdd OAI21X1
XOAI21X1_100 DFFSR_95/Q INVX1_32/Y NAND2X1_32/Y gnd MUX2X1_44/A vdd OAI21X1
XOAI21X1_144 BUFX4_36/Y MUX2X1_50/Y OAI21X1_143/Y gnd DFFPOSX1_28/D vdd OAI21X1
XOAI21X1_166 INVX1_45/Y NAND2X1_39/Y NAND3X1_13/Y gnd OAI21X1_168/A vdd OAI21X1
XOAI21X1_122 BUFX4_38/Y MUX2X1_39/Y OAI21X1_121/Y gnd OAI21X1_122/Y vdd OAI21X1
XOAI21X1_133 BUFX4_34/Y BUFX4_57/Y INVX1_46/A gnd OAI21X1_134/C vdd OAI21X1
XOAI21X1_111 OR2X2_3/A OR2X2_3/B INVX1_25/A gnd INVX1_35/A vdd OAI21X1
XAOI22X1_9 DFFSR_68/Q AOI21X1_9/A DFFSR_11/Q NOR2X1_48/Y gnd AOI22X1_9/Y vdd AOI22X1
XNAND2X1_19 MUX2X1_24/B NOR2X1_9/Y gnd NAND2X1_19/Y vdd NAND2X1
XNAND2X1_161 NOR2X1_4/A DFFSR_171/D gnd NAND2X1_161/Y vdd NAND2X1
XNAND2X1_150 DFFSR_49/Q NOR2X1_48/Y gnd NAND3X1_42/B vdd NAND2X1
XNAND2X1_183 NAND2X1_182/Y NAND2X1_183/B gnd DFFSR_177/D vdd NAND2X1
XNAND2X1_172 NAND3X1_62/Y NAND3X1_61/Y gnd OAI21X1_457/A vdd NAND2X1
XAOI22X1_17 DFFSR_69/Q AOI21X1_9/A DFFSR_31/Q NOR2X1_49/Y gnd AOI22X1_17/Y vdd AOI22X1
XFILL_10_3_1 gnd vdd FILL
XOAI21X1_1 NOR2X1_4/A NOR2X1_4/B INVX1_2/Y gnd BUFX4_13/A vdd OAI21X1
XFILL_9_0_0 gnd vdd FILL
XXOR2X1_4 OR2X2_3/A OR2X2_3/B gnd XOR2X1_4/Y vdd XOR2X1
XMUX2X1_5 MUX2X1_5/A MUX2X1_5/B MUX2X1_5/S gnd MUX2X1_5/Y vdd MUX2X1
XCLKBUF1_6 BUFX4_4/Y gnd DFFSR_2/CLK vdd CLKBUF1
XFILL_24_3 gnd vdd FILL
XFILL_24_2_1 gnd vdd FILL
XINVX8_8 rst gnd INVX8_8/Y vdd INVX8
XDFFPOSX1_72 MUX2X1_58/B CLKBUF1_41/Y OAI21X1_197/Y gnd vdd DFFPOSX1
XDFFPOSX1_61 INVX1_60/A CLKBUF1_9/Y DFFPOSX1_61/D gnd vdd DFFPOSX1
XDFFPOSX1_94 MUX2X1_82/B CLKBUF1_25/Y DFFPOSX1_94/D gnd vdd DFFPOSX1
XDFFPOSX1_50 MUX2X1_74/B CLKBUF1_9/Y DFFPOSX1_50/D gnd vdd DFFPOSX1
XDFFPOSX1_83 INVX1_94/A CLKBUF1_14/Y DFFPOSX1_83/D gnd vdd DFFPOSX1
XBUFX4_39 BUFX4_36/A gnd AND2X2_2/A vdd BUFX4
XFILL_7_3_1 gnd vdd FILL
XBUFX4_28 INVX8_3/Y gnd BUFX4_28/Y vdd BUFX4
XBUFX4_17 BUFX4_18/A gnd BUFX4_17/Y vdd BUFX4
XFILL_15_2_1 gnd vdd FILL
XFILL_21_0_1 gnd vdd FILL
XOAI21X1_315 BUFX4_21/Y BUFX4_83/Y MUX2X1_99/B gnd OAI21X1_315/Y vdd OAI21X1
XOAI21X1_359 BUFX4_74/Y OR2X2_9/B DFFSR_84/Q gnd OAI21X1_360/C vdd OAI21X1
XDFFSR_150 INVX1_8/A CLKBUF1_38/Y BUFX4_66/Y vdd DFFSR_150/D gnd vdd DFFSR
XDFFSR_161 INVX1_55/A CLKBUF1_38/Y BUFX4_68/Y vdd DFFSR_161/D gnd vdd DFFSR
XOAI21X1_326 BUFX4_47/Y MUX2X1_104/Y OAI21X1_326/C gnd OAI21X1_326/Y vdd OAI21X1
XOAI21X1_337 INVX1_90/Y NAND2X1_97/Y NAND2X1_101/Y gnd OAI21X1_337/Y vdd OAI21X1
XOAI21X1_348 INVX1_95/Y NAND2X1_95/Y NAND3X1_28/Y gnd OAI21X1_350/A vdd OAI21X1
XOAI21X1_304 BUFX4_45/Y MUX2X1_93/Y OAI21X1_304/C gnd DFFPOSX1_79/D vdd OAI21X1
XDFFSR_172 INVX2_8/A CLKBUF1_35/Y BUFX4_69/Y vdd DFFSR_172/D gnd vdd DFFSR
XBUFX4_2 clk gnd BUFX4_2/Y vdd BUFX4
XFILL_4_1_1 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XINVX4_2 rst gnd INVX4_2/Y vdd INVX4
XNAND3X1_5 MUX2X1_4/B DFFSR_14/Q INVX2_1/A gnd NAND3X1_5/Y vdd NAND3X1
XOAI21X1_101 BUFX4_34/Y BUFX4_55/Y MUX2X1_30/B gnd OAI21X1_102/C vdd OAI21X1
XOAI21X1_112 INVX1_35/Y DFFSR_21/D NOR2X1_16/Y gnd NAND2X1_37/A vdd OAI21X1
XOAI21X1_189 DFFSR_109/Q INVX1_56/Y NAND2X1_60/Y gnd MUX2X1_56/A vdd OAI21X1
XOAI21X1_123 BUFX4_34/Y BUFX4_55/Y INVX1_47/A gnd OAI21X1_124/C vdd OAI21X1
XOAI21X1_156 OAI21X1_154/Y OAI21X1_156/B NOR2X1_16/Y gnd NAND2X1_44/B vdd OAI21X1
XOAI21X1_178 BUFX2_3/Y OR2X2_4/A DFFSR_25/Q gnd NAND2X1_56/A vdd OAI21X1
XOAI21X1_134 BUFX4_38/Y MUX2X1_45/Y OAI21X1_134/C gnd OAI21X1_134/Y vdd OAI21X1
XOAI21X1_167 INVX1_46/Y NAND2X1_41/Y NAND2X1_49/Y gnd OAI21X1_168/B vdd OAI21X1
XOAI21X1_145 BUFX4_33/Y BUFX4_54/Y MUX2X1_51/B gnd OAI21X1_146/C vdd OAI21X1
XNAND2X1_140 BUFX2_26/A MUX2X1_105/Y gnd AOI21X1_6/A vdd NAND2X1
XNAND2X1_173 INVX2_10/A INVX4_3/Y gnd NAND2X1_173/Y vdd NAND2X1
XNAND2X1_162 BUFX4_8/Y gnd gnd OAI22X1_6/B vdd NAND2X1
XNAND2X1_151 AOI22X1_9/Y AOI22X1_10/Y gnd OAI21X1_436/A vdd NAND2X1
XAOI22X1_18 DFFSR_50/Q AND2X2_5/Y DFFSR_12/Q NOR2X1_48/Y gnd AOI22X1_18/Y vdd AOI22X1
XFILL_10_3_2 gnd vdd FILL
XOAI21X1_2 NOR2X1_4/B INVX1_3/Y NAND2X1_1/Y gnd MUX2X1_1/A vdd OAI21X1
XFILL_9_0_1 gnd vdd FILL
XXOR2X1_5 XOR2X1_5/A OR2X2_5/B gnd DFFSR_55/D vdd XOR2X1
XMUX2X1_6 MUX2X1_6/A MUX2X1_6/B MUX2X1_5/S gnd MUX2X1_6/Y vdd MUX2X1
XCLKBUF1_7 BUFX4_2/Y gnd CLKBUF1_7/Y vdd CLKBUF1
XFILL_24_4 gnd vdd FILL
XFILL_24_2_2 gnd vdd FILL
XINVX8_9 rst gnd INVX8_9/Y vdd INVX8
XDFFPOSX1_73 MUX2X1_99/B CLKBUF1_14/Y OAI21X1_316/Y gnd vdd DFFPOSX1
XDFFPOSX1_40 INVX1_43/A CLKBUF1_20/Y DFFPOSX1_40/D gnd vdd DFFPOSX1
XFILL_7_3_2 gnd vdd FILL
XDFFPOSX1_84 INVX1_96/A DFFSR_36/CLK DFFPOSX1_84/D gnd vdd DFFPOSX1
XDFFPOSX1_51 MUX2X1_75/B CLKBUF1_24/Y DFFPOSX1_51/D gnd vdd DFFPOSX1
XDFFPOSX1_95 MUX2X1_83/B CLKBUF1_14/Y DFFPOSX1_95/D gnd vdd DFFPOSX1
XDFFPOSX1_62 INVX1_63/A CLKBUF1_9/Y DFFPOSX1_62/D gnd vdd DFFPOSX1
XBUFX4_18 BUFX4_18/A gnd BUFX4_18/Y vdd BUFX4
XBUFX4_29 INVX8_3/Y gnd DFFSR_41/R vdd BUFX4
XFILL_15_2_2 gnd vdd FILL
XFILL_22_1 gnd vdd FILL
XFILL_21_0_2 gnd vdd FILL
XOAI21X1_305 BUFX4_20/Y BUFX4_84/Y INVX1_88/A gnd OAI21X1_305/Y vdd OAI21X1
XOAI21X1_327 BUFX4_89/Y OR2X2_8/A DFFSR_64/Q gnd NAND2X1_98/A vdd OAI21X1
XOAI21X1_316 BUFX4_45/Y MUX2X1_99/Y OAI21X1_315/Y gnd OAI21X1_316/Y vdd OAI21X1
XDFFSR_140 NOR2X1_15/A CLKBUF1_35/Y BUFX4_67/Y vdd DFFSR_140/D gnd vdd DFFSR
XDFFSR_173 INVX2_9/A CLKBUF1_12/Y BUFX4_66/Y vdd DFFSR_173/D gnd vdd DFFSR
XBUFX4_3 clk gnd BUFX4_3/Y vdd BUFX4
XDFFSR_162 INVX1_56/A CLKBUF1_38/Y BUFX4_66/Y vdd DFFSR_162/D gnd vdd DFFSR
XDFFSR_151 INVX1_9/A CLKBUF1_12/Y BUFX4_66/Y vdd DFFSR_151/D gnd vdd DFFSR
XOAI21X1_349 INVX1_96/Y NAND2X1_97/Y NAND2X1_107/Y gnd OAI21X1_349/Y vdd OAI21X1
XOAI21X1_338 OAI21X1_336/Y OAI21X1_337/Y NOR2X1_36/Y gnd NAND2X1_111/B vdd OAI21X1
XFILL_4_1_2 gnd vdd FILL
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XFILL_12_0_2 gnd vdd FILL
XNAND3X1_6 MUX2X1_5/B DFFSR_14/Q INVX2_1/A gnd NAND3X1_6/Y vdd NAND3X1
XFILL_22_3_0 gnd vdd FILL
XOAI21X1_124 BUFX4_40/Y MUX2X1_40/Y OAI21X1_124/C gnd OAI21X1_124/Y vdd OAI21X1
XOAI21X1_102 BUFX4_37/Y MUX2X1_30/Y OAI21X1_102/C gnd OAI21X1_102/Y vdd OAI21X1
XOAI21X1_113 BUFX4_35/Y BUFX4_56/Y INVX1_36/A gnd OAI21X1_113/Y vdd OAI21X1
XOAI21X1_135 BUFX4_33/Y BUFX4_54/Y INVX1_48/A gnd OAI21X1_135/Y vdd OAI21X1
XOAI21X1_146 AND2X2_2/A MUX2X1_51/Y OAI21X1_146/C gnd DFFPOSX1_29/D vdd OAI21X1
XOAI21X1_168 OAI21X1_168/A OAI21X1_168/B NOR2X1_16/Y gnd NAND2X1_50/B vdd OAI21X1
XOAI21X1_157 BUFX4_58/Y OR2X2_4/A DFFSR_28/Q gnd NAND2X1_46/A vdd OAI21X1
XOAI21X1_179 INVX1_161/A DFFSR_109/Q INVX1_50/Y gnd BUFX4_93/A vdd OAI21X1
XNAND2X1_130 DFFSR_132/Q DFFSR_61/Q gnd OAI21X1_422/C vdd NAND2X1
XNAND2X1_141 INVX1_148/Y MUX2X1_106/Y gnd AOI21X1_6/B vdd NAND2X1
XNAND2X1_152 DFFSR_135/Q DFFSR_137/D gnd OAI21X1_439/C vdd NAND2X1
XNAND2X1_163 BUFX4_9/Y INVX4_5/Y gnd OAI22X1_7/B vdd NAND2X1
XNAND2X1_174 NAND2X1_173/Y NAND2X1_174/B gnd DFFSR_174/D vdd NAND2X1
XFILL_13_3_0 gnd vdd FILL
XOAI21X1_3 BUFX4_74/Y BUFX4_42/Y MUX2X1_1/B gnd OAI21X1_3/Y vdd OAI21X1
XFILL_9_0_2 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XXOR2X1_6 OR2X2_5/A OR2X2_5/B gnd XOR2X1_6/Y vdd XOR2X1
XMUX2X1_7 OR2X2_1/A XOR2X1_2/Y MUX2X1_7/S gnd MUX2X1_8/A vdd MUX2X1
XCLKBUF1_8 BUFX4_4/Y gnd DFFSR_1/CLK vdd CLKBUF1
XFILL_10_1_0 gnd vdd FILL
XFILL_18_2_0 gnd vdd FILL
XDFFPOSX1_30 MUX2X1_52/B CLKBUF1_27/Y OAI21X1_148/Y gnd vdd DFFPOSX1
XDFFPOSX1_41 INVX1_45/A CLKBUF1_42/Y OAI21X1_122/Y gnd vdd DFFPOSX1
XDFFPOSX1_52 MUX2X1_76/B CLKBUF1_9/Y DFFPOSX1_52/D gnd vdd DFFPOSX1
XDFFPOSX1_63 INVX1_65/A DFFSR_54/CLK OAI21X1_207/Y gnd vdd DFFPOSX1
XDFFPOSX1_85 INVX1_84/A CLKBUF1_14/Y OAI21X1_292/Y gnd vdd DFFPOSX1
XDFFPOSX1_74 NAND2X1_99/A CLKBUF1_25/Y DFFPOSX1_74/D gnd vdd DFFPOSX1
XBUFX4_19 DFFSR_58/Q gnd BUFX4_19/Y vdd BUFX4
XDFFPOSX1_96 MUX2X1_84/B CLKBUF1_7/Y OAI21X1_286/Y gnd vdd DFFPOSX1
XFILL_22_2 gnd vdd FILL
XFILL_15_1 gnd vdd FILL
XFILL_24_0_0 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XOAI21X1_328 INVX1_84/Y NAND2X1_95/Y NAND3X1_23/Y gnd OAI21X1_328/Y vdd OAI21X1
XOAI21X1_317 BUFX4_20/Y BUFX4_84/Y NAND2X1_99/A gnd OAI21X1_318/C vdd OAI21X1
XOAI21X1_306 BUFX4_49/Y MUX2X1_94/Y OAI21X1_305/Y gnd OAI21X1_306/Y vdd OAI21X1
XDFFSR_130 DFFSR_130/Q CLKBUF1_32/Y INVX8_8/Y vdd DFFSR_130/D gnd vdd DFFSR
XOAI21X1_339 BUFX4_91/Y OR2X2_8/A DFFSR_67/Q gnd OAI21X1_339/Y vdd OAI21X1
XBUFX4_4 clk gnd BUFX4_4/Y vdd BUFX4
XDFFSR_152 INVX1_10/A CLKBUF1_38/Y BUFX4_66/Y vdd DFFSR_152/D gnd vdd DFFSR
XDFFSR_174 INVX2_10/A CLKBUF1_34/Y BUFX4_71/Y vdd DFFSR_174/D gnd vdd DFFSR
XDFFSR_163 INVX1_57/A CLKBUF1_12/Y BUFX4_68/Y vdd DFFSR_163/D gnd vdd DFFSR
XDFFSR_141 NOR2X1_25/A CLKBUF1_12/Y BUFX4_69/Y vdd DFFSR_141/D gnd vdd DFFSR
XINVX4_4 INVX4_4/A gnd INVX4_4/Y vdd INVX4
XNAND3X1_7 MUX2X1_6/B DFFSR_14/Q INVX2_1/A gnd NAND3X1_7/Y vdd NAND3X1
XFILL_22_3_1 gnd vdd FILL
XOAI21X1_158 INVX1_41/Y NAND2X1_39/Y NAND3X1_11/Y gnd OAI21X1_158/Y vdd OAI21X1
XOAI21X1_114 BUFX4_36/Y MUX2X1_35/Y OAI21X1_113/Y gnd OAI21X1_114/Y vdd OAI21X1
XOAI21X1_147 BUFX4_33/Y BUFX4_57/Y MUX2X1_52/B gnd OAI21X1_148/C vdd OAI21X1
XOAI21X1_103 DFFSR_95/Q INVX1_33/Y NAND2X1_33/Y gnd MUX2X1_39/B vdd OAI21X1
XOAI21X1_136 BUFX4_38/Y MUX2X1_46/Y OAI21X1_135/Y gnd DFFPOSX1_36/D vdd OAI21X1
XOAI21X1_169 OR2X2_4/B OR2X2_4/A DFFSR_31/Q gnd NAND2X1_52/A vdd OAI21X1
XOAI21X1_125 BUFX4_33/Y BUFX4_54/Y INVX1_37/A gnd OAI21X1_126/C vdd OAI21X1
XBUFX2_1 BUFX4_8/A gnd BUFX2_1/Y vdd BUFX2
XNAND2X1_131 DFFSR_132/Q DFFSR_62/Q gnd NAND2X1_131/Y vdd NAND2X1
XNAND2X1_142 AOI21X1_6/A AOI21X1_6/B gnd NOR2X1_50/B vdd NAND2X1
XNAND2X1_120 DFFSR_104/Q DFFSR_23/Q gnd OAI21X1_388/C vdd NAND2X1
XNAND2X1_164 INVX4_3/A NOR2X1_54/Y gnd MUX2X1_118/S vdd NAND2X1
XNAND2X1_175 NAND3X1_65/Y NAND3X1_64/Y gnd NAND2X1_175/Y vdd NAND2X1
XNAND2X1_153 DFFSR_31/Q NOR2X1_48/Y gnd NAND3X1_45/B vdd NAND2X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XFILL_13_3_1 gnd vdd FILL
XAOI21X1_1 NAND2X1_8/Y AOI21X1_1/B AND2X2_1/A gnd AOI21X1_1/Y vdd AOI21X1
XOAI21X1_4 BUFX4_14/Y MUX2X1_1/Y OAI21X1_3/Y gnd OAI21X1_4/Y vdd OAI21X1
XXOR2X1_7 XOR2X1_7/A OR2X2_7/B gnd XOR2X1_7/Y vdd XOR2X1
XFILL_2_2_1 gnd vdd FILL
XMUX2X1_8 MUX2X1_8/A XOR2X1_2/Y OR2X2_2/Y gnd MUX2X1_8/Y vdd MUX2X1
XFILL_10_1_1 gnd vdd FILL
XCLKBUF1_9 BUFX4_1/Y gnd CLKBUF1_9/Y vdd CLKBUF1
XFILL_18_2_1 gnd vdd FILL
XDFFPOSX1_53 MUX2X1_77/B CLKBUF1_26/Y DFFPOSX1_53/D gnd vdd DFFPOSX1
XDFFPOSX1_64 INVX1_67/A CLKBUF1_41/Y OAI21X1_209/Y gnd vdd DFFPOSX1
XDFFPOSX1_42 INVX1_47/A CLKBUF1_36/Y OAI21X1_124/Y gnd vdd DFFPOSX1
XDFFPOSX1_20 MUX2X1_2/B CLKBUF1_40/Y OAI21X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_31 INVX1_37/A CLKBUF1_42/Y OAI21X1_126/Y gnd vdd DFFPOSX1
XDFFPOSX1_75 MUX2X1_101/B DFFSR_36/CLK DFFPOSX1_75/D gnd vdd DFFPOSX1
XDFFPOSX1_86 INVX1_87/A CLKBUF1_25/Y OAI21X1_294/Y gnd vdd DFFPOSX1
XFILL_22_3 gnd vdd FILL
XFILL_15_2 gnd vdd FILL
XINVX1_180 DFFSR_7/Q gnd INVX1_180/Y vdd INVX1
XFILL_24_0_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XOAI21X1_329 INVX1_85/Y NAND2X1_97/Y NAND2X1_96/Y gnd OAI21X1_329/Y vdd OAI21X1
XOAI21X1_307 BUFX4_22/Y BUFX4_81/Y INVX1_90/A gnd OAI21X1_308/C vdd OAI21X1
XOAI21X1_318 BUFX4_49/Y MUX2X1_100/Y OAI21X1_318/C gnd DFFPOSX1_74/D vdd OAI21X1
XDFFSR_120 BUFX2_19/A CLKBUF1_5/Y INVX8_8/Y vdd DFFSR_120/D gnd vdd DFFSR
XDFFSR_131 BUFX2_25/A CLKBUF1_32/Y INVX8_8/Y vdd DFFSR_131/D gnd vdd DFFSR
XDFFSR_164 INVX1_58/A CLKBUF1_38/Y BUFX4_68/Y vdd DFFSR_164/D gnd vdd DFFSR
XDFFSR_153 INVX1_27/A DFFSR_33/CLK BUFX4_71/Y vdd DFFSR_153/D gnd vdd DFFSR
XDFFSR_175 INVX2_11/A DFFSR_45/CLK BUFX4_69/Y vdd DFFSR_175/D gnd vdd DFFSR
XDFFSR_142 DFFSR_142/Q CLKBUF1_30/Y BUFX4_70/Y vdd OAI22X1_6/Y gnd vdd DFFSR
XBUFX4_5 clk gnd BUFX4_5/Y vdd BUFX4
XINVX4_5 gnd gnd INVX4_5/Y vdd INVX4
XNAND3X1_8 OR2X2_3/A OR2X2_3/B INVX1_25/Y gnd AOI21X1_2/B vdd NAND3X1
XFILL_22_3_2 gnd vdd FILL
XOAI21X1_104 BUFX4_34/Y BUFX4_57/Y MUX2X1_31/B gnd OAI21X1_105/C vdd OAI21X1
XOAI21X1_115 BUFX4_32/Y BUFX4_56/Y INVX1_39/A gnd OAI21X1_116/C vdd OAI21X1
XOAI21X1_159 INVX1_42/Y NAND2X1_41/Y NAND2X1_45/Y gnd OAI21X1_160/B vdd OAI21X1
XOAI21X1_137 BUFX4_33/Y BUFX4_54/Y MUX2X1_47/B gnd OAI21X1_138/C vdd OAI21X1
XOAI21X1_148 BUFX4_36/Y MUX2X1_52/Y OAI21X1_148/C gnd OAI21X1_148/Y vdd OAI21X1
XOAI21X1_126 AND2X2_2/A MUX2X1_41/Y OAI21X1_126/C gnd OAI21X1_126/Y vdd OAI21X1
XNAND2X1_132 DFFSR_132/Q DFFSR_63/Q gnd OAI21X1_424/C vdd NAND2X1
XNAND2X1_110 NAND2X1_110/A NAND2X1_110/B gnd DFFSR_61/D vdd NAND2X1
XNAND2X1_143 DFFSR_137/Q NOR2X1_50/B gnd NOR2X1_53/A vdd NAND2X1
XNAND2X1_121 DFFSR_104/Q DFFSR_24/Q gnd OAI21X1_389/C vdd NAND2X1
XBUFX2_2 BUFX2_2/A gnd BUFX2_2/Y vdd BUFX2
XNAND2X1_165 gnd INVX4_4/Y gnd OAI22X1_9/B vdd NAND2X1
XNAND2X1_176 INVX2_11/A INVX4_3/Y gnd NAND2X1_176/Y vdd NAND2X1
XNAND2X1_154 DFFSR_50/Q NOR2X1_49/Y gnd NAND3X1_45/C vdd NAND2X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XFILL_13_3_2 gnd vdd FILL
XAOI21X1_2 AOI21X1_2/A AOI21X1_2/B AND2X2_2/A gnd AOI21X1_2/Y vdd AOI21X1
XXNOR2X1_10 AND2X2_4/A DFFSR_72/Q gnd DFFSR_72/D vdd XNOR2X1
XBUFX2_20 BUFX2_20/A gnd ext_data_out[14] vdd BUFX2
XAOI21X1_10 NAND3X1_51/Y AOI21X1_10/B NOR2X1_52/A gnd AOI21X1_10/Y vdd AOI21X1
XOAI21X1_5 NOR2X1_4/B INVX1_6/Y NAND2X1_2/Y gnd MUX2X1_2/A vdd OAI21X1
XXOR2X1_8 OR2X2_7/A OR2X2_7/B gnd XOR2X1_8/Y vdd XOR2X1
XFILL_2_2_2 gnd vdd FILL
XMUX2X1_9 INVX1_12/A MUX2X1_1/A MUX2X1_9/S gnd MUX2X1_9/Y vdd MUX2X1
XFILL_10_1_2 gnd vdd FILL
XFILL_18_2_2 gnd vdd FILL
XDFFPOSX1_65 INVX1_69/A CLKBUF1_26/Y OAI21X1_211/Y gnd vdd DFFPOSX1
XDFFPOSX1_54 MUX2X1_78/B CLKBUF1_41/Y OAI21X1_237/Y gnd vdd DFFPOSX1
XDFFPOSX1_32 INVX1_40/A CLKBUF1_27/Y OAI21X1_128/Y gnd vdd DFFPOSX1
XDFFPOSX1_10 INVX1_20/A CLKBUF1_4/Y OAI21X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_43 NAND3X1_9/A CLKBUF1_20/Y OAI21X1_93/Y gnd vdd DFFPOSX1
XDFFPOSX1_21 MUX2X1_3/B DFFSR_1/CLK OAI21X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_76 MUX2X1_102/B CLKBUF1_7/Y OAI21X1_322/Y gnd vdd DFFPOSX1
XDFFPOSX1_87 INVX1_89/A CLKBUF1_30/Y DFFPOSX1_87/D gnd vdd DFFPOSX1
XFILL_15_3 gnd vdd FILL
XINVX1_170 INVX1_55/A gnd INVX1_170/Y vdd INVX1
XINVX1_181 DFFSR_8/Q gnd INVX1_181/Y vdd INVX1
XFILL_24_0_2 gnd vdd FILL
XFILL_7_1_2 gnd vdd FILL
XFILL_15_0_2 gnd vdd FILL
XFILL_20_1 gnd vdd FILL
XDFFSR_121 BUFX2_20/A DFFSR_74/CLK INVX8_8/Y vdd DFFSR_121/D gnd vdd DFFSR
XDFFSR_132 DFFSR_132/Q DFFSR_60/CLK INVX8_8/Y vdd NOR2X1_35/B gnd vdd DFFSR
XDFFSR_143 NOR2X1_4/A CLKBUF1_12/Y BUFX4_69/Y vdd DFFSR_143/D gnd vdd DFFSR
XDFFSR_110 NOR2X1_25/B CLKBUF1_38/Y INVX8_7/Y vdd INVX1_132/Y gnd vdd DFFSR
XOAI21X1_308 BUFX4_46/Y MUX2X1_95/Y OAI21X1_308/C gnd OAI21X1_308/Y vdd OAI21X1
XOAI21X1_319 BUFX4_22/Y BUFX4_81/Y MUX2X1_101/B gnd OAI21X1_319/Y vdd OAI21X1
XDFFSR_154 INVX1_30/A CLKBUF1_16/Y BUFX4_67/Y vdd DFFSR_154/D gnd vdd DFFSR
XBUFX4_6 clk gnd BUFX4_6/Y vdd BUFX4
XDFFSR_165 INVX1_75/A DFFSR_21/CLK BUFX4_71/Y vdd DFFSR_165/D gnd vdd DFFSR
XDFFSR_176 INVX2_12/A DFFSR_45/CLK BUFX4_69/Y vdd DFFSR_176/D gnd vdd DFFSR
XFILL_0_3_0 gnd vdd FILL
XFILL_16_3_0 gnd vdd FILL
XNAND3X1_9 NAND3X1_9/A DFFSR_33/Q INVX2_2/A gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_127 BUFX4_35/Y BUFX4_56/Y INVX1_40/A gnd OAI21X1_127/Y vdd OAI21X1
XOAI21X1_116 BUFX4_37/Y MUX2X1_36/Y OAI21X1_116/C gnd DFFPOSX1_38/D vdd OAI21X1
XOAI21X1_149 BUFX4_59/Y OR2X2_4/A DFFSR_26/Q gnd NAND2X1_42/A vdd OAI21X1
XBUFX2_3 BUFX2_3/A gnd BUFX2_3/Y vdd BUFX2
XOAI21X1_138 BUFX4_36/Y MUX2X1_47/Y OAI21X1_138/C gnd DFFPOSX1_25/D vdd OAI21X1
XOAI21X1_105 BUFX4_38/Y MUX2X1_31/Y OAI21X1_105/C gnd OAI21X1_105/Y vdd OAI21X1
XNAND2X1_133 INVX4_1/A INVX2_6/Y gnd OAI22X1_4/D vdd NAND2X1
XNAND2X1_111 NAND2X1_111/A NAND2X1_111/B gnd DFFSR_62/D vdd NAND2X1
XNAND2X1_144 INVX2_6/A INVX4_1/Y gnd OAI21X1_427/B vdd NAND2X1
XNAND2X1_122 DFFSR_104/Q DFFSR_25/Q gnd OAI21X1_390/C vdd NAND2X1
XNAND2X1_166 NAND3X1_56/Y NAND3X1_55/Y gnd OAI21X1_453/A vdd NAND2X1
XNAND2X1_177 NAND2X1_176/Y OAI21X1_459/Y gnd DFFSR_175/D vdd NAND2X1
XNAND2X1_100 OAI21X1_331/Y NAND2X1_110/B gnd DFFSR_65/D vdd NAND2X1
XNAND2X1_155 DFFSR_31/Q AOI21X1_9/A gnd NAND3X1_48/A vdd NAND2X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XAOI21X1_3 AOI21X1_3/A AOI21X1_3/B BUFX4_93/Y gnd AOI21X1_3/Y vdd AOI21X1
XXNOR2X1_11 NOR2X1_40/Y INVX1_76/Y gnd DFFSR_73/D vdd XNOR2X1
XBUFX2_10 BUFX2_10/A gnd ext_data_out[4] vdd BUFX2
XINVX1_90 INVX1_90/A gnd INVX1_90/Y vdd INVX1
XBUFX2_21 BUFX2_21/A gnd ext_data_out[15] vdd BUFX2
XNOR2X1_1 INVX1_1/A OR2X2_1/Y gnd DFFSR_2/D vdd NOR2X1
XFILL_22_1_0 gnd vdd FILL
XAOI21X1_11 NOR2X1_47/Y NAND3X1_39/Y AOI21X1_8/C gnd AOI21X1_11/Y vdd AOI21X1
XOAI21X1_6 OR2X2_9/A BUFX4_44/Y MUX2X1_2/B gnd OAI21X1_6/Y vdd OAI21X1
XFILL_5_2_0 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XDFFPOSX1_11 INVX1_22/A CLKBUF1_31/Y OAI21X1_45/Y gnd vdd DFFPOSX1
XDFFPOSX1_66 INVX1_71/A CLKBUF1_41/Y OAI21X1_213/Y gnd vdd DFFPOSX1
XDFFPOSX1_22 MUX2X1_4/B CLKBUF1_40/Y OAI21X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_44 MUX2X1_28/B CLKBUF1_36/Y OAI21X1_96/Y gnd vdd DFFPOSX1
XDFFPOSX1_33 INVX1_42/A CLKBUF1_27/Y DFFPOSX1_33/D gnd vdd DFFPOSX1
XDFFPOSX1_88 INVX1_91/A DFFSR_36/CLK DFFPOSX1_88/D gnd vdd DFFPOSX1
XDFFPOSX1_77 MUX2X1_103/B CLKBUF1_14/Y DFFPOSX1_77/D gnd vdd DFFPOSX1
XDFFPOSX1_55 INVX1_61/A CLKBUF1_9/Y DFFPOSX1_55/D gnd vdd DFFPOSX1
XFILL_2_0_0 gnd vdd FILL
XFILL_18_0_0 gnd vdd FILL
XINVX1_182 DFFSR_9/Q gnd INVX1_182/Y vdd INVX1
XINVX1_171 INVX1_56/A gnd INVX1_171/Y vdd INVX1
XINVX1_160 gnd gnd INVX1_160/Y vdd INVX1
XFILL_20_2 gnd vdd FILL
XDFFSR_122 BUFX2_21/A DFFSR_61/CLK INVX8_8/Y vdd DFFSR_122/D gnd vdd DFFSR
XDFFSR_111 DFFSR_111/Q CLKBUF1_21/Y INVX8_7/Y vdd DFFSR_111/D gnd vdd DFFSR
XDFFSR_100 DFFSR_100/Q CLKBUF1_13/Y INVX8_6/Y vdd DFFSR_100/D gnd vdd DFFSR
XDFFSR_144 INVX1_159/A CLKBUF1_16/Y BUFX4_67/Y vdd DFFSR_144/D gnd vdd DFFSR
XDFFSR_155 INVX1_31/A DFFSR_21/CLK BUFX4_71/Y vdd DFFSR_155/D gnd vdd DFFSR
XDFFSR_133 BUFX4_8/A DFFSR_45/CLK INVX4_2/Y vdd DFFSR_133/D gnd vdd DFFSR
XOAI21X1_309 BUFX4_22/Y BUFX4_84/Y INVX1_92/A gnd OAI21X1_309/Y vdd OAI21X1
XBUFX4_7 BUFX4_8/A gnd INVX4_4/A vdd BUFX4
XDFFSR_166 INVX1_78/A CLKBUF1_30/Y BUFX4_70/Y vdd DFFSR_166/D gnd vdd DFFSR
XDFFSR_177 INVX2_13/A CLKBUF1_35/Y BUFX4_67/Y vdd DFFSR_177/D gnd vdd DFFSR
XFILL_0_3_1 gnd vdd FILL
XFILL_16_3_1 gnd vdd FILL
XOAI21X1_128 BUFX4_36/Y MUX2X1_42/Y OAI21X1_127/Y gnd OAI21X1_128/Y vdd OAI21X1
XOAI21X1_117 BUFX4_32/Y BUFX4_55/Y INVX1_41/A gnd OAI21X1_117/Y vdd OAI21X1
XOAI21X1_106 DFFSR_95/Q INVX1_34/Y NAND2X1_34/Y gnd MUX2X1_46/A vdd OAI21X1
XBUFX2_4 BUFX2_4/A gnd BUFX2_4/Y vdd BUFX2
XOAI21X1_139 BUFX4_32/Y BUFX4_55/Y MUX2X1_48/B gnd OAI21X1_139/Y vdd OAI21X1
XNAND2X1_134 INVX2_6/A INVX4_1/A gnd OAI22X1_4/B vdd NAND2X1
XNAND2X1_112 NAND2X1_112/A NAND2X1_112/B gnd DFFSR_63/D vdd NAND2X1
XNAND2X1_123 BUFX4_65/Y BUFX2_24/A gnd OAI21X1_403/C vdd NAND2X1
XNAND2X1_145 OAI21X1_427/B OAI22X1_4/D gnd NAND2X1_145/Y vdd NAND2X1
XNAND2X1_167 INVX2_8/A INVX4_3/Y gnd NAND2X1_168/A vdd NAND2X1
XNAND2X1_101 MUX2X1_101/B NOR2X1_39/Y gnd NAND2X1_101/Y vdd NAND2X1
XNAND2X1_178 NAND3X1_68/Y NAND3X1_67/Y gnd OAI21X1_461/A vdd NAND2X1
XNAND2X1_156 DFFSR_69/Q NOR2X1_49/Y gnd NAND3X1_48/B vdd NAND2X1
XAOI21X1_4 AOI21X1_4/A AOI21X1_4/B AND2X2_4/A gnd AOI21X1_4/Y vdd AOI21X1
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XXNOR2X1_12 NOR2X1_36/Y INVX2_4/Y gnd DFFSR_70/D vdd XNOR2X1
XBUFX2_22 OR2X2_9/B gnd pe_busy[0] vdd BUFX2
XBUFX2_11 DFFSR_92/Q gnd ext_data_out[5] vdd BUFX2
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XNOR2X1_2 INVX1_1/Y OR2X2_1/Y gnd DFFSR_1/D vdd NOR2X1
XFILL_22_1_1 gnd vdd FILL
XAOI21X1_12 INVX2_8/Y NOR2X1_58/B NOR2X1_56/Y gnd DFFSR_147/D vdd AOI21X1
XOAI21X1_7 BUFX4_10/Y MUX2X1_2/Y OAI21X1_6/Y gnd OAI21X1_7/Y vdd OAI21X1
XFILL_5_2_1 gnd vdd FILL
XFILL_13_1_1 gnd vdd FILL
XFILL_1_1 gnd vdd FILL
XDFFPOSX1_34 INVX1_44/A CLKBUF1_36/Y DFFPOSX1_34/D gnd vdd DFFPOSX1
XDFFPOSX1_45 MUX2X1_29/B CLKBUF1_20/Y OAI21X1_99/Y gnd vdd DFFPOSX1
XDFFPOSX1_12 INVX1_24/A CLKBUF1_40/Y OAI21X1_47/Y gnd vdd DFFPOSX1
XDFFPOSX1_23 MUX2X1_5/B CLKBUF1_31/Y OAI21X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_67 MUX2X1_53/B CLKBUF1_41/Y OAI21X1_182/Y gnd vdd DFFPOSX1
XDFFPOSX1_56 INVX1_64/A CLKBUF1_21/Y DFFPOSX1_56/D gnd vdd DFFPOSX1
XDFFPOSX1_78 MUX2X1_104/B DFFSR_36/CLK OAI21X1_326/Y gnd vdd DFFPOSX1
XDFFPOSX1_89 INVX1_93/A CLKBUF1_14/Y OAI21X1_300/Y gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XFILL_18_0_1 gnd vdd FILL
XINVX1_150 AOI21X1_8/C gnd INVX1_150/Y vdd INVX1
XINVX1_183 DFFSR_10/Q gnd INVX1_183/Y vdd INVX1
XINVX1_172 INVX1_57/A gnd INVX1_172/Y vdd INVX1
XINVX1_161 INVX1_161/A gnd INVX1_161/Y vdd INVX1
XFILL_20_3 gnd vdd FILL
XDFFSR_123 DFFSR_123/Q DFFSR_60/CLK INVX8_8/Y vdd DFFSR_123/D gnd vdd DFFSR
XDFFSR_101 INVX1_114/A CLKBUF1_13/Y INVX8_6/Y vdd DFFSR_101/D gnd vdd DFFSR
XDFFSR_156 INVX1_32/A CLKBUF1_34/Y BUFX4_67/Y vdd DFFSR_156/D gnd vdd DFFSR
XDFFSR_178 NOR2X1_5/A CLKBUF1_35/Y BUFX4_67/Y vdd DFFSR_178/D gnd vdd DFFSR
XDFFSR_112 DFFSR_112/Q CLKBUF1_9/Y INVX8_7/Y vdd DFFSR_112/D gnd vdd DFFSR
XDFFSR_145 INVX1_161/A CLKBUF1_12/Y BUFX4_69/Y vdd DFFSR_145/D gnd vdd DFFSR
XDFFSR_167 INVX1_79/A DFFSR_21/CLK BUFX4_70/Y vdd DFFSR_167/D gnd vdd DFFSR
XBUFX4_8 BUFX4_8/A gnd BUFX4_8/Y vdd BUFX4
XDFFSR_134 BUFX2_26/A DFFSR_45/CLK INVX4_2/Y vdd DFFSR_134/D gnd vdd DFFSR
XFILL_0_3_2 gnd vdd FILL
XFILL_16_3_2 gnd vdd FILL
XOAI21X1_118 BUFX4_40/Y MUX2X1_37/Y OAI21X1_117/Y gnd OAI21X1_118/Y vdd OAI21X1
XOAI21X1_129 BUFX4_34/Y BUFX4_57/Y INVX1_42/A gnd OAI21X1_130/C vdd OAI21X1
XOAI21X1_107 BUFX4_33/Y BUFX4_54/Y MUX2X1_32/B gnd OAI21X1_107/Y vdd OAI21X1
XBUFX2_5 DFFSR_2/Q gnd BUFX2_5/Y vdd BUFX2
XNAND2X1_146 INVX4_1/Y AOI21X1_7/Y gnd AOI21X1_8/A vdd NAND2X1
XNAND2X1_124 DFFSR_41/Q DFFSR_118/Q gnd NAND2X1_124/Y vdd NAND2X1
XNAND2X1_135 BUFX4_25/Y AOI21X1_9/A gnd NAND3X1_30/C vdd NAND2X1
XNAND2X1_113 BUFX4_76/Y OR2X2_9/B gnd OAI21X1_369/C vdd NAND2X1
XNAND2X1_168 NAND2X1_168/A NAND2X1_168/B gnd DFFSR_172/D vdd NAND2X1
XNAND2X1_179 INVX2_12/A INVX4_3/Y gnd NAND2X1_179/Y vdd NAND2X1
XNAND2X1_157 AOI22X1_17/Y AOI22X1_18/Y gnd NAND2X1_157/Y vdd NAND2X1
XNAND2X1_102 OAI21X1_335/Y NAND2X1_111/B gnd DFFSR_66/D vdd NAND2X1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XAOI21X1_5 AOI21X1_9/A BUFX2_4/Y INVX2_7/A gnd AOI21X1_5/Y vdd AOI21X1
XXNOR2X1_13 XNOR2X1_13/A INVX2_6/A gnd DFFSR_138/D vdd XNOR2X1
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XBUFX2_23 OR2X2_10/B gnd pe_busy[1] vdd BUFX2
XBUFX2_12 BUFX2_12/A gnd ext_data_out[6] vdd BUFX2
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XNOR2X1_3 INVX1_4/Y INVX1_5/Y gnd MUX2X1_5/S vdd NOR2X1
XFILL_22_1_2 gnd vdd FILL
XAOI21X1_13 INVX2_9/Y NOR2X1_58/B NOR2X1_57/Y gnd DFFSR_148/D vdd AOI21X1
XOAI21X1_8 NOR2X1_4/B INVX1_7/Y NAND2X1_3/Y gnd MUX2X1_3/A vdd OAI21X1
XFILL_5_2_2 gnd vdd FILL
XFILL_13_1_2 gnd vdd FILL
XOAI21X1_460 INVX1_184/Y OR2X2_14/Y NAND3X1_66/Y gnd OAI21X1_461/B vdd OAI21X1
XOAI21X1_290 INVX1_83/Y DFFSR_59/D NOR2X1_36/Y gnd NAND2X1_93/A vdd OAI21X1
XDFFPOSX1_46 MUX2X1_30/B CLKBUF1_36/Y OAI21X1_102/Y gnd vdd DFFPOSX1
XDFFPOSX1_13 INVX1_12/A DFFSR_89/CLK OAI21X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_35 INVX1_46/A CLKBUF1_42/Y OAI21X1_134/Y gnd vdd DFFPOSX1
XDFFPOSX1_24 MUX2X1_6/B CLKBUF1_31/Y OAI21X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_68 MUX2X1_54/B CLKBUF1_24/Y DFFPOSX1_68/D gnd vdd DFFPOSX1
XDFFPOSX1_57 INVX1_66/A DFFSR_50/CLK DFFPOSX1_57/D gnd vdd DFFPOSX1
XDFFPOSX1_79 INVX1_85/A CLKBUF1_14/Y DFFPOSX1_79/D gnd vdd DFFPOSX1
XFILL_2_0_2 gnd vdd FILL
XDFFSR_90 DFFSR_90/Q DFFSR_23/CLK INVX8_5/Y vdd NOR2X1_5/B gnd vdd DFFSR
XFILL_18_0_2 gnd vdd FILL
XINVX1_140 BUFX2_18/A gnd INVX1_140/Y vdd INVX1
XINVX1_173 INVX1_58/A gnd INVX1_173/Y vdd INVX1
XINVX1_162 INVX1_75/A gnd INVX1_162/Y vdd INVX1
XINVX1_184 DFFSR_11/Q gnd INVX1_184/Y vdd INVX1
XINVX1_151 OAI22X1_3/Y gnd AOI22X1_8/A vdd INVX1
XFILL_20_2_0 gnd vdd FILL
XFILL_3_3_0 gnd vdd FILL
XFILL_11_2_0 gnd vdd FILL
XFILL_19_3_0 gnd vdd FILL
XDFFSR_113 DFFSR_113/Q CLKBUF1_26/Y INVX8_7/Y vdd DFFSR_113/D gnd vdd DFFSR
XDFFSR_124 NOR2X1_35/B DFFSR_60/CLK INVX8_8/Y vdd DFFSR_124/D gnd vdd DFFSR
XDFFSR_135 DFFSR_135/Q DFFSR_67/CLK INVX4_2/Y vdd DFFSR_135/D gnd vdd DFFSR
XDFFSR_102 DFFSR_102/Q CLKBUF1_13/Y INVX8_6/Y vdd DFFSR_102/D gnd vdd DFFSR
XDFFSR_157 INVX1_33/A CLKBUF1_16/Y BUFX4_67/Y vdd DFFSR_157/D gnd vdd DFFSR
XBUFX4_9 BUFX4_8/A gnd BUFX4_9/Y vdd BUFX4
XDFFSR_168 INVX1_80/A CLKBUF1_30/Y BUFX4_70/Y vdd DFFSR_168/D gnd vdd DFFSR
XDFFSR_146 NOR2X1_34/A CLKBUF1_30/Y BUFX4_70/Y vdd DFFSR_146/D gnd vdd DFFSR
XOAI21X1_119 BUFX4_32/Y BUFX4_55/Y INVX1_43/A gnd OAI21X1_119/Y vdd OAI21X1
XOAI21X1_108 BUFX4_36/Y MUX2X1_32/Y OAI21X1_107/Y gnd DFFPOSX1_48/D vdd OAI21X1
XNAND2X1_114 DFFSR_3/Q DFFSR_90/Q gnd OAI21X1_370/C vdd NAND2X1
XBUFX2_6 BUFX2_6/A gnd ext_data_out[0] vdd BUFX2
XNAND2X1_103 MUX2X1_102/B NOR2X1_39/Y gnd OAI21X1_341/C vdd NAND2X1
XNAND2X1_125 DFFSR_118/Q DFFSR_42/Q gnd NAND2X1_125/Y vdd NAND2X1
XNAND2X1_136 BUFX4_25/Y INVX4_1/A gnd OAI21X1_425/C vdd NAND2X1
XNAND2X1_158 INVX2_6/Y AOI21X1_7/C gnd AOI21X1_10/B vdd NAND2X1
XNAND2X1_1 NOR2X1_4/B DFFSR_83/Q gnd NAND2X1_1/Y vdd NAND2X1
XNAND2X1_169 NAND3X1_59/Y NAND3X1_58/Y gnd OAI21X1_455/A vdd NAND2X1
XNAND2X1_147 BUFX2_26/A DFFSR_137/D gnd OAI21X1_437/C vdd NAND2X1
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XFILL_0_1_0 gnd vdd FILL
XAOI21X1_6 AOI21X1_6/A AOI21X1_6/B INVX4_1/Y gnd AOI21X1_6/Y vdd AOI21X1
XMUX2X1_120 INVX1_175/Y INVX2_9/Y MUX2X1_122/S gnd DFFSR_154/D vdd MUX2X1
XFILL_8_2_0 gnd vdd FILL
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XINVX1_71 INVX1_71/A gnd INVX1_71/Y vdd INVX1
XDFFPOSX1_1 MUX2X1_21/B CLKBUF1_4/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XBUFX2_13 BUFX2_13/A gnd ext_data_out[7] vdd BUFX2
XINVX1_82 INVX1_82/A gnd INVX1_82/Y vdd INVX1
XFILL_16_1_0 gnd vdd FILL
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XBUFX2_24 BUFX2_24/A gnd pe_busy[2] vdd BUFX2
XNOR2X1_4 NOR2X1_4/A NOR2X1_4/B gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_14 INVX2_10/Y NOR2X1_58/B NOR2X1_58/Y gnd DFFSR_149/D vdd AOI21X1
XOAI21X1_9 BUFX4_76/Y BUFX4_43/Y MUX2X1_3/B gnd OAI21X1_9/Y vdd OAI21X1
XOAI21X1_450 INVX1_161/Y OAI22X1_6/A MUX2X1_118/S gnd DFFSR_145/D vdd OAI21X1
XOAI21X1_461 OAI21X1_461/A OAI21X1_461/B INVX4_3/A gnd NAND2X1_180/B vdd OAI21X1
XFILL_5_0_0 gnd vdd FILL
XOAI21X1_280 BUFX4_49/Y MUX2X1_82/Y OAI21X1_279/Y gnd DFFPOSX1_94/D vdd OAI21X1
XOAI21X1_291 OR2X2_12/A BUFX4_83/Y INVX1_84/A gnd OAI21X1_291/Y vdd OAI21X1
XDFFPOSX1_58 INVX1_68/A CLKBUF1_21/Y DFFPOSX1_58/D gnd vdd DFFPOSX1
XDFFPOSX1_69 MUX2X1_55/B CLKBUF1_26/Y OAI21X1_188/Y gnd vdd DFFPOSX1
XDFFPOSX1_14 INVX1_15/A CLKBUF1_40/Y OAI21X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_25 MUX2X1_47/B CLKBUF1_27/Y DFFPOSX1_25/D gnd vdd DFFPOSX1
XDFFPOSX1_47 MUX2X1_31/B CLKBUF1_42/Y OAI21X1_105/Y gnd vdd DFFPOSX1
XDFFPOSX1_36 INVX1_48/A CLKBUF1_42/Y DFFPOSX1_36/D gnd vdd DFFPOSX1
XDFFSR_80 BUFX2_9/A DFFSR_9/CLK INVX8_5/Y vdd DFFSR_80/D gnd vdd DFFSR
XDFFSR_91 BUFX2_10/A DFFSR_23/CLK INVX8_6/Y vdd DFFSR_91/D gnd vdd DFFSR
XINVX1_141 BUFX2_19/A gnd INVX1_141/Y vdd INVX1
XINVX1_130 BUFX2_16/A gnd INVX1_130/Y vdd INVX1
XINVX1_152 NOR2X1_45/B gnd INVX1_152/Y vdd INVX1
XINVX1_174 INVX1_27/A gnd INVX1_174/Y vdd INVX1
XINVX1_185 DFFSR_12/Q gnd INVX1_185/Y vdd INVX1
XINVX1_163 INVX1_78/A gnd INVX1_163/Y vdd INVX1
XFILL_20_2_1 gnd vdd FILL
XFILL_3_3_1 gnd vdd FILL
XFILL_11_2_1 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XDFFSR_114 DFFSR_114/Q CLKBUF1_21/Y INVX8_7/Y vdd DFFSR_114/D gnd vdd DFFSR
XDFFSR_103 OR2X2_10/B CLKBUF1_20/Y INVX8_6/Y vdd DFFSR_103/D gnd vdd DFFSR
XDFFSR_125 DFFSR_125/Q DFFSR_67/CLK INVX8_8/Y vdd DFFSR_125/D gnd vdd DFFSR
XDFFSR_136 INVX2_7/A CLKBUF1_5/Y INVX4_2/Y vdd NOR2X1_53/Y gnd vdd DFFSR
XDFFSR_147 INVX1_3/A DFFSR_87/CLK BUFX4_68/Y vdd DFFSR_147/D gnd vdd DFFSR
XDFFSR_158 INVX1_34/A DFFSR_21/CLK BUFX4_71/Y vdd DFFSR_158/D gnd vdd DFFSR
XDFFSR_169 INVX1_81/A CLKBUF1_30/Y BUFX4_71/Y vdd DFFSR_169/D gnd vdd DFFSR
XBUFX2_7 BUFX2_7/A gnd ext_data_out[1] vdd BUFX2
XOAI21X1_109 OR2X2_4/B OR2X2_4/A AND2X2_2/A gnd XOR2X1_3/A vdd OAI21X1
XFILL_11_1 gnd vdd FILL
XNAND2X1_137 INVX2_6/Y OAI21X1_425/Y gnd NAND3X1_34/B vdd NAND2X1
XNAND2X1_104 OAI21X1_339/Y NAND2X1_112/B gnd DFFSR_67/D vdd NAND2X1
XNAND2X1_159 INVX2_6/Y NOR2X1_46/A gnd NAND2X1_159/Y vdd NAND2X1
XNAND2X1_115 DFFSR_90/Q DFFSR_4/Q gnd OAI21X1_371/C vdd NAND2X1
XNAND2X1_126 DFFSR_118/Q DFFSR_43/Q gnd OAI21X1_406/C vdd NAND2X1
XNAND2X1_148 AOI22X1_2/Y AOI22X1_3/Y gnd NAND3X1_40/A vdd NAND2X1
XNAND2X1_2 NOR2X1_4/B DFFSR_84/Q gnd NAND2X1_2/Y vdd NAND2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XFILL_0_1_1 gnd vdd FILL
XAOI21X1_7 NOR2X1_47/Y INVX2_6/A AOI21X1_7/C gnd AOI21X1_7/Y vdd AOI21X1
XMUX2X1_121 INVX1_176/Y INVX2_10/Y MUX2X1_122/S gnd DFFSR_155/D vdd MUX2X1
XMUX2X1_110 INVX1_165/Y INVX2_11/Y MUX2X1_108/S gnd DFFSR_168/D vdd MUX2X1
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XFILL_8_2_1 gnd vdd FILL
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XINVX1_50 BUFX4_61/Y gnd INVX1_50/Y vdd INVX1
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XBUFX2_14 BUFX2_14/A gnd ext_data_out[8] vdd BUFX2
XBUFX2_25 BUFX2_25/A gnd pe_busy[3] vdd BUFX2
XDFFPOSX1_2 MUX2X1_22/B DFFSR_1/CLK OAI21X1_51/Y gnd vdd DFFPOSX1
XFILL_16_1_1 gnd vdd FILL
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd OR2X2_2/A vdd NOR2X1
XAOI21X1_15 INVX2_11/Y NOR2X1_58/B NOR2X1_59/Y gnd DFFSR_150/D vdd AOI21X1
XOAI21X1_440 OAI22X1_3/Y NOR2X1_45/B INVX2_6/A gnd OAI21X1_440/Y vdd OAI21X1
XOAI21X1_451 BUFX4_9/Y INVX4_5/Y NOR2X1_25/A gnd OAI22X1_9/D vdd OAI21X1
XOAI21X1_462 INVX1_185/Y OR2X2_14/Y NAND3X1_69/Y gnd OAI21X1_463/B vdd OAI21X1
XFILL_5_0_1 gnd vdd FILL
XOAI21X1_281 DFFSR_123/Q INVX1_81/Y NAND2X1_89/Y gnd MUX2X1_97/A vdd OAI21X1
XOAI21X1_292 BUFX4_45/Y MUX2X1_87/Y OAI21X1_291/Y gnd OAI21X1_292/Y vdd OAI21X1
XOAI21X1_270 OR2X2_12/A BUFX4_82/Y MUX2X1_79/B gnd OAI21X1_270/Y vdd OAI21X1
XDFFPOSX1_59 INVX1_70/A CLKBUF1_26/Y OAI21X1_223/Y gnd vdd DFFPOSX1
XDFFPOSX1_37 INVX1_36/A CLKBUF1_27/Y OAI21X1_114/Y gnd vdd DFFPOSX1
XDFFPOSX1_15 INVX1_17/A DFFSR_89/CLK OAI21X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_48 MUX2X1_32/B CLKBUF1_27/Y DFFPOSX1_48/D gnd vdd DFFPOSX1
XDFFPOSX1_26 MUX2X1_48/B CLKBUF1_20/Y OAI21X1_140/Y gnd vdd DFFPOSX1
XDFFSR_70 INVX2_4/A CLKBUF1_32/Y DFFSR_71/R vdd DFFSR_70/D gnd vdd DFFSR
XDFFSR_81 NOR2X1_4/B CLKBUF1_4/Y INVX8_5/Y vdd INVX1_97/Y gnd vdd DFFSR
XDFFSR_92 DFFSR_92/Q DFFSR_23/CLK INVX8_6/Y vdd DFFSR_92/D gnd vdd DFFSR
XINVX1_142 BUFX2_20/A gnd INVX1_142/Y vdd INVX1
XINVX1_120 BUFX4_59/Y gnd DFFSR_96/D vdd INVX1
XINVX1_175 INVX1_30/A gnd INVX1_175/Y vdd INVX1
XINVX1_164 INVX1_79/A gnd INVX1_164/Y vdd INVX1
XINVX1_131 BUFX2_17/A gnd INVX1_131/Y vdd INVX1
XINVX1_153 OAI22X1_1/Y gnd AOI22X1_5/A vdd INVX1
XFILL_20_2_2 gnd vdd FILL
XFILL_3_3_2 gnd vdd FILL
XFILL_11_2_2 gnd vdd FILL
XFILL_19_3_2 gnd vdd FILL
XDFFSR_126 DFFSR_126/Q DFFSR_61/CLK INVX8_8/Y vdd DFFSR_126/D gnd vdd DFFSR
XDFFSR_137 DFFSR_137/Q DFFSR_50/CLK INVX4_2/Y vdd DFFSR_137/D gnd vdd DFFSR
XDFFSR_104 DFFSR_104/Q DFFSR_8/CLK INVX8_6/Y vdd DFFSR_96/Q gnd vdd DFFSR
XDFFSR_148 INVX1_6/A DFFSR_2/CLK BUFX4_66/Y vdd DFFSR_148/D gnd vdd DFFSR
XDFFSR_115 INVX1_126/A CLKBUF1_24/Y INVX8_7/Y vdd DFFSR_115/D gnd vdd DFFSR
XDFFSR_159 INVX1_51/A CLKBUF1_31/Y BUFX4_68/Y vdd DFFSR_159/D gnd vdd DFFSR
XNAND3X1_70 BUFX4_8/Y DFFSR_31/Q INVX4_5/Y gnd NAND3X1_70/Y vdd NAND3X1
XFILL_11_2 gnd vdd FILL
XBUFX2_8 BUFX2_8/A gnd ext_data_out[2] vdd BUFX2
XNAND2X1_138 INVX4_1/A BUFX4_89/Y gnd OAI21X1_426/C vdd NAND2X1
XNAND2X1_116 DFFSR_90/Q DFFSR_5/Q gnd OAI21X1_372/C vdd NAND2X1
XNAND2X1_3 NOR2X1_4/B DFFSR_85/Q gnd NAND2X1_3/Y vdd NAND2X1
XNAND2X1_127 DFFSR_118/Q DFFSR_44/Q gnd OAI21X1_407/C vdd NAND2X1
XNAND2X1_149 DFFSR_30/Q AOI21X1_9/A gnd NAND3X1_42/A vdd NAND2X1
XNAND2X1_105 MUX2X1_103/B NOR2X1_39/Y gnd OAI21X1_345/C vdd NAND2X1
XFILL_0_1_2 gnd vdd FILL
XAOI21X1_8 AOI21X1_8/A AOI21X1_8/B AOI21X1_8/C gnd AOI21X1_8/Y vdd AOI21X1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XMUX2X1_122 INVX1_177/Y INVX2_11/Y MUX2X1_122/S gnd DFFSR_156/D vdd MUX2X1
XMUX2X1_111 INVX1_166/Y INVX2_12/Y MUX2X1_108/S gnd DFFSR_169/D vdd MUX2X1
XMUX2X1_100 MUX2X1_94/A NAND2X1_99/A NOR2X1_38/Y gnd MUX2X1_100/Y vdd MUX2X1
XINVX1_73 DFFSR_76/Q gnd INVX1_73/Y vdd INVX1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XFILL_8_2_2 gnd vdd FILL
XBUFX2_26 BUFX2_26/A gnd BUFX2_26/Y vdd BUFX2
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XINVX1_62 DFFSR_52/Q gnd INVX1_62/Y vdd INVX1
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XBUFX2_15 BUFX2_15/A gnd ext_data_out[9] vdd BUFX2
XDFFPOSX1_3 MUX2X1_23/B DFFSR_87/CLK OAI21X1_53/Y gnd vdd DFFPOSX1
XFILL_16_1_2 gnd vdd FILL
XNOR2X1_6 OR2X2_2/B OR2X2_2/A gnd NOR2X1_6/Y vdd NOR2X1
XAOI21X1_16 INVX2_12/Y NOR2X1_58/B NOR2X1_60/Y gnd DFFSR_151/D vdd AOI21X1
XOAI21X1_430 OAI22X1_2/Y NOR2X1_43/B NOR2X1_44/A gnd NOR2X1_52/B vdd OAI21X1
XOAI21X1_441 OAI21X1_440/Y AOI21X1_11/Y NAND2X1_159/Y gnd OAI21X1_441/Y vdd OAI21X1
XOAI21X1_452 INVX1_180/Y OR2X2_14/Y NAND3X1_54/Y gnd OAI21X1_453/B vdd OAI21X1
XOAI21X1_463 OAI21X1_463/A OAI21X1_463/B INVX4_3/A gnd NAND2X1_183/B vdd OAI21X1
XOAI21X1_90 INVX1_159/A DFFSR_95/Q INVX1_26/Y gnd BUFX4_36/A vdd OAI21X1
XFILL_5_0_2 gnd vdd FILL
XOAI21X1_293 BUFX4_19/Y BUFX4_83/Y INVX1_87/A gnd OAI21X1_294/C vdd OAI21X1
XOAI21X1_282 BUFX4_19/Y BUFX4_83/Y MUX2X1_83/B gnd OAI21X1_282/Y vdd OAI21X1
XOAI21X1_271 AND2X2_4/A MUX2X1_79/Y OAI21X1_270/Y gnd OAI21X1_271/Y vdd OAI21X1
XOAI21X1_260 INVX1_72/Y NAND2X1_69/Y NAND2X1_79/Y gnd OAI21X1_261/B vdd OAI21X1
XDFFPOSX1_27 MUX2X1_49/B CLKBUF1_36/Y OAI21X1_142/Y gnd vdd DFFPOSX1
XDFFPOSX1_16 INVX1_19/A DFFSR_89/CLK OAI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_38 INVX1_39/A CLKBUF1_20/Y DFFPOSX1_38/D gnd vdd DFFPOSX1
XDFFPOSX1_49 MUX2X1_73/B CLKBUF1_24/Y DFFPOSX1_49/D gnd vdd DFFPOSX1
XFILL_23_2_0 gnd vdd FILL
XDFFSR_60 DFFSR_60/Q DFFSR_60/CLK BUFX4_88/Y vdd DFFSR_60/D gnd vdd DFFSR
XDFFSR_71 DFFSR_71/Q CLKBUF1_32/Y DFFSR_71/R vdd DFFSR_71/D gnd vdd DFFSR
XDFFSR_82 NOR2X1_5/B DFFSR_8/CLK INVX8_5/Y vdd DFFSR_82/D gnd vdd DFFSR
XDFFSR_93 BUFX2_12/A DFFSR_23/CLK INVX8_6/Y vdd DFFSR_93/D gnd vdd DFFSR
XFILL_6_3_0 gnd vdd FILL
XFILL_14_2_0 gnd vdd FILL
XINVX1_143 BUFX2_21/A gnd INVX1_143/Y vdd INVX1
XINVX1_121 OR2X2_11/Y gnd INVX1_121/Y vdd INVX1
XINVX1_110 ext_data_in[4] gnd INVX1_110/Y vdd INVX1
XINVX1_176 INVX1_31/A gnd INVX1_176/Y vdd INVX1
XINVX1_132 BUFX2_2/Y gnd INVX1_132/Y vdd INVX1
XINVX1_165 INVX1_80/A gnd INVX1_165/Y vdd INVX1
XINVX1_154 NOR2X1_42/B gnd AOI22X1_5/B vdd INVX1
XDFFSR_138 INVX2_6/A CLKBUF1_5/Y INVX4_2/Y vdd DFFSR_138/D gnd vdd DFFSR
XDFFSR_105 BUFX2_14/A CLKBUF1_5/Y INVX8_7/Y vdd DFFSR_105/D gnd vdd DFFSR
XDFFSR_127 DFFSR_127/Q DFFSR_61/CLK INVX8_8/Y vdd DFFSR_127/D gnd vdd DFFSR
XDFFSR_149 INVX1_7/A CLKBUF1_31/Y BUFX4_68/Y vdd DFFSR_149/D gnd vdd DFFSR
XDFFSR_116 INVX1_127/A CLKBUF1_9/Y INVX8_7/Y vdd DFFSR_116/D gnd vdd DFFSR
XFILL_20_0_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XNOR2X1_60 INVX1_9/A NOR2X1_58/B gnd NOR2X1_60/Y vdd NOR2X1
XNAND3X1_60 gnd DFFSR_47/Q INVX4_4/Y gnd NAND3X1_60/Y vdd NAND3X1
XNAND3X1_71 BUFX4_8/Y gnd DFFSR_69/Q gnd NAND3X1_71/Y vdd NAND3X1
XFILL_19_1_0 gnd vdd FILL
XBUFX2_9 BUFX2_9/A gnd ext_data_out[3] vdd BUFX2
XNAND2X1_139 INVX2_6/A NAND2X1_139/B gnd NAND3X1_34/C vdd NAND2X1
XNAND2X1_128 OR2X2_12/A BUFX2_25/A gnd OAI21X1_420/C vdd NAND2X1
XNAND2X1_4 NOR2X1_4/B DFFSR_86/Q gnd NAND2X1_4/Y vdd NAND2X1
XNAND2X1_117 DFFSR_90/Q DFFSR_6/Q gnd OAI21X1_373/C vdd NAND2X1
XNAND2X1_106 NAND2X1_106/A NAND2X1_106/B gnd DFFSR_68/D vdd NAND2X1
XAOI21X1_9 AOI21X1_9/A BUFX4_58/Y INVX2_7/A gnd AOI21X1_9/Y vdd AOI21X1
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XMUX2X1_123 INVX1_178/Y INVX2_12/Y MUX2X1_122/S gnd DFFSR_157/D vdd MUX2X1
XMUX2X1_112 INVX1_167/Y INVX2_13/Y MUX2X1_108/S gnd DFFSR_170/D vdd MUX2X1
XMUX2X1_101 MUX2X1_89/B MUX2X1_101/B NOR2X1_38/Y gnd MUX2X1_101/Y vdd MUX2X1
XINVX1_52 DFFSR_54/Q gnd INVX1_52/Y vdd INVX1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XBUFX2_16 BUFX2_16/A gnd ext_data_out[10] vdd BUFX2
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XINVX1_74 BUFX4_19/Y gnd INVX1_74/Y vdd INVX1
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XDFFPOSX1_4 MUX2X1_24/B CLKBUF1_4/Y OAI21X1_55/Y gnd vdd DFFPOSX1
XNOR2X1_7 INVX1_4/A INVX1_5/Y gnd NOR2X1_7/Y vdd NOR2X1
XAOI21X1_17 INVX2_13/Y NOR2X1_58/B NOR2X1_61/Y gnd DFFSR_152/D vdd AOI21X1
XOAI21X1_431 NOR2X1_48/Y NOR2X1_49/Y NOR2X1_50/B gnd OAI21X1_431/Y vdd OAI21X1
XOAI21X1_420 OR2X2_12/A DFFSR_123/Q OAI21X1_420/C gnd DFFSR_131/D vdd OAI21X1
XOAI21X1_442 AOI21X1_10/Y OAI21X1_441/Y DFFSR_137/Q gnd OAI21X1_443/C vdd OAI21X1
XOAI21X1_453 OAI21X1_453/A OAI21X1_453/B INVX4_3/A gnd NAND2X1_168/B vdd OAI21X1
XFILL_8_0_0 gnd vdd FILL
XOAI21X1_91 DFFSR_95/Q INVX1_27/Y NAND2X1_29/Y gnd MUX2X1_41/A vdd OAI21X1
XOAI21X1_80 INVX2_5/A OR2X2_2/A DFFSR_12/Q gnd NAND2X1_24/A vdd OAI21X1
XOAI21X1_250 BUFX4_26/Y OR2X2_6/A DFFSR_48/Q gnd NAND2X1_76/A vdd OAI21X1
XOAI21X1_294 BUFX4_46/Y MUX2X1_88/Y OAI21X1_294/C gnd OAI21X1_294/Y vdd OAI21X1
XOAI21X1_272 DFFSR_123/Q INVX1_78/Y NAND2X1_86/Y gnd MUX2X1_94/A vdd OAI21X1
XOAI21X1_261 OAI21X1_261/A OAI21X1_261/B NOR2X1_26/Y gnd NAND2X1_80/B vdd OAI21X1
XOAI21X1_283 BUFX4_45/Y MUX2X1_83/Y OAI21X1_282/Y gnd DFFPOSX1_95/D vdd OAI21X1
XDFFPOSX1_39 INVX1_41/A CLKBUF1_36/Y OAI21X1_118/Y gnd vdd DFFPOSX1
XDFFPOSX1_28 MUX2X1_50/B CLKBUF1_20/Y DFFPOSX1_28/D gnd vdd DFFPOSX1
XDFFPOSX1_17 INVX1_21/A CLKBUF1_31/Y OAI21X1_33/Y gnd vdd DFFPOSX1
XFILL_23_2_1 gnd vdd FILL
XDFFSR_61 DFFSR_61/Q DFFSR_61/CLK BUFX4_88/Y vdd DFFSR_61/D gnd vdd DFFSR
XDFFSR_72 DFFSR_72/Q CLKBUF1_32/Y DFFSR_71/R vdd DFFSR_72/D gnd vdd DFFSR
XDFFSR_94 BUFX2_13/A DFFSR_23/CLK INVX8_6/Y vdd DFFSR_94/D gnd vdd DFFSR
XDFFSR_83 DFFSR_83/Q DFFSR_87/CLK INVX8_5/Y vdd DFFSR_83/D gnd vdd DFFSR
XDFFSR_50 DFFSR_50/Q DFFSR_50/CLK DFFSR_41/R vdd DFFSR_50/D gnd vdd DFFSR
XFILL_6_3_1 gnd vdd FILL
XFILL_14_2_1 gnd vdd FILL
XINVX1_100 ext_data_in[2] gnd INVX1_100/Y vdd INVX1
XINVX1_122 ext_data_in[8] gnd INVX1_122/Y vdd INVX1
XINVX1_133 OR2X2_12/Y gnd DFFSR_123/D vdd INVX1
XINVX1_144 BUFX4_89/Y gnd DFFSR_124/D vdd INVX1
XINVX1_111 ext_data_in[5] gnd INVX1_111/Y vdd INVX1
XINVX1_177 INVX1_32/A gnd INVX1_177/Y vdd INVX1
XINVX1_166 INVX1_81/A gnd INVX1_166/Y vdd INVX1
XINVX1_155 NOR2X1_46/A gnd INVX1_155/Y vdd INVX1
XDFFSR_117 BUFX2_24/A CLKBUF1_21/Y INVX8_7/Y vdd DFFSR_117/D gnd vdd DFFSR
XDFFSR_139 INVX4_1/A CLKBUF1_5/Y INVX4_2/Y vdd DFFSR_139/D gnd vdd DFFSR
XDFFSR_128 DFFSR_128/Q DFFSR_61/CLK INVX8_8/Y vdd DFFSR_128/D gnd vdd DFFSR
XDFFSR_106 BUFX2_15/A DFFSR_45/CLK INVX8_7/Y vdd DFFSR_106/D gnd vdd DFFSR
XFILL_20_0_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XNAND3X1_50 NAND3X1_50/A NAND3X1_50/B AOI21X1_8/C gnd NAND3X1_50/Y vdd NAND3X1
XNOR2X1_50 INVX4_1/A NOR2X1_50/B gnd NOR2X1_50/Y vdd NOR2X1
XNOR2X1_61 INVX1_10/A NOR2X1_58/B gnd NOR2X1_61/Y vdd NOR2X1
XNAND3X1_61 BUFX2_1/Y DFFSR_28/Q INVX4_5/Y gnd NAND3X1_61/Y vdd NAND3X1
XFILL_19_1_1 gnd vdd FILL
XNAND2X1_107 MUX2X1_104/B NOR2X1_39/Y gnd NAND2X1_107/Y vdd NAND2X1
XNAND2X1_129 DFFSR_60/Q DFFSR_132/Q gnd OAI21X1_421/C vdd NAND2X1
XNAND2X1_118 BUFX4_35/Y OR2X2_10/B gnd OAI21X1_386/C vdd NAND2X1
XNAND2X1_5 NOR2X1_4/B DFFSR_87/Q gnd NAND2X1_5/Y vdd NAND2X1
XMUX2X1_90 INVX1_91/A MUX2X1_82/A MUX2X1_87/S gnd MUX2X1_90/Y vdd MUX2X1
XMUX2X1_113 INVX1_168/Y INVX2_8/Y MUX2X1_118/S gnd DFFSR_159/D vdd MUX2X1
XMUX2X1_102 MUX2X1_82/A MUX2X1_102/B NOR2X1_38/Y gnd MUX2X1_102/Y vdd MUX2X1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XMUX2X1_124 INVX1_179/Y INVX2_13/Y MUX2X1_122/S gnd DFFSR_158/D vdd MUX2X1
XINVX1_53 DFFSR_53/Q gnd INVX1_53/Y vdd INVX1
XINVX1_97 OR2X2_9/Y gnd INVX1_97/Y vdd INVX1
XDFFPOSX1_5 MUX2X1_25/B DFFSR_2/CLK OAI21X1_57/Y gnd vdd DFFPOSX1
XBUFX2_17 BUFX2_17/A gnd ext_data_out[11] vdd BUFX2
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XINVX1_64 INVX1_64/A gnd INVX1_64/Y vdd INVX1
XINVX1_86 DFFSR_71/Q gnd INVX1_86/Y vdd INVX1
XNOR2X1_8 INVX1_4/A INVX1_5/A gnd NOR2X1_8/Y vdd NOR2X1
XOAI21X1_421 DFFSR_132/Q INVX1_140/Y OAI21X1_421/C gnd DFFSR_119/D vdd OAI21X1
XOAI21X1_410 BUFX4_21/Y BUFX2_25/A DFFSR_126/Q gnd OAI21X1_410/Y vdd OAI21X1
XOAI21X1_432 OAI22X1_3/Y NOR2X1_45/B DFFSR_137/Q gnd NOR2X1_51/A vdd OAI21X1
XOAI21X1_454 INVX1_181/Y OR2X2_14/Y NAND3X1_57/Y gnd OAI21X1_455/B vdd OAI21X1
XOAI21X1_443 DFFSR_137/Q INVX1_156/Y OAI21X1_443/C gnd DFFSR_133/D vdd OAI21X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_81 INVX1_23/Y OAI21X1_69/B NAND3X1_7/Y gnd OAI21X1_81/Y vdd OAI21X1
XOAI21X1_70 INVX1_18/Y OAI21X1_78/B NAND2X1_17/Y gnd OAI21X1_71/B vdd OAI21X1
XOAI21X1_92 BUFX4_32/Y BUFX4_56/Y NAND3X1_9/A gnd OAI21X1_93/C vdd OAI21X1
XOAI21X1_273 BUFX4_19/Y BUFX4_81/Y MUX2X1_80/B gnd OAI21X1_274/C vdd OAI21X1
XOAI21X1_240 INVX1_61/Y NAND2X1_69/Y NAND2X1_68/Y gnd OAI21X1_240/Y vdd OAI21X1
XOAI21X1_262 INVX2_3/Y OR2X2_6/Y DFFSR_52/Q gnd OAI21X1_262/Y vdd OAI21X1
XOAI21X1_251 INVX1_67/Y NAND2X1_67/Y NAND3X1_19/Y gnd OAI21X1_253/A vdd OAI21X1
XOAI21X1_295 BUFX4_19/Y BUFX4_83/Y INVX1_89/A gnd OAI21X1_296/C vdd OAI21X1
XOAI21X1_284 DFFSR_123/Q INVX1_82/Y NAND2X1_90/Y gnd MUX2X1_92/B vdd OAI21X1
XDFFPOSX1_18 INVX1_23/A DFFSR_87/CLK OAI21X1_35/Y gnd vdd DFFPOSX1
XDFFPOSX1_29 MUX2X1_51/B DFFSR_33/CLK DFFPOSX1_29/D gnd vdd DFFPOSX1
XFILL_23_2_2 gnd vdd FILL
XDFFSR_62 DFFSR_62/Q DFFSR_74/CLK DFFSR_74/R vdd DFFSR_62/D gnd vdd DFFSR
XDFFSR_40 BUFX2_2/A DFFSR_54/CLK vdd DFFSR_54/R DFFSR_40/D gnd vdd DFFSR
XDFFSR_84 DFFSR_84/Q CLKBUF1_4/Y INVX8_5/Y vdd DFFSR_84/D gnd vdd DFFSR
XDFFSR_95 DFFSR_95/Q CLKBUF1_13/Y INVX8_6/Y vdd DFFSR_95/D gnd vdd DFFSR
XDFFSR_51 INVX2_3/A CLKBUF1_3/Y DFFSR_43/R vdd DFFSR_51/D gnd vdd DFFSR
XDFFSR_73 DFFSR_73/Q CLKBUF1_7/Y DFFSR_71/R vdd DFFSR_73/D gnd vdd DFFSR
XFILL_6_3_2 gnd vdd FILL
XFILL_14_2_2 gnd vdd FILL
XINVX1_134 ext_data_in[12] gnd INVX1_134/Y vdd INVX1
XINVX1_101 ext_data_in[3] gnd INVX1_101/Y vdd INVX1
XINVX1_112 ext_data_in[6] gnd INVX1_112/Y vdd INVX1
XINVX1_123 ext_data_in[9] gnd INVX1_123/Y vdd INVX1
XINVX1_178 INVX1_33/A gnd INVX1_178/Y vdd INVX1
XINVX1_167 INVX1_82/A gnd INVX1_167/Y vdd INVX1
XINVX1_156 INVX4_4/A gnd INVX1_156/Y vdd INVX1
XINVX1_145 DFFSR_137/Q gnd DFFSR_137/D vdd INVX1
XDFFSR_107 BUFX2_16/A CLKBUF1_24/Y INVX8_7/Y vdd DFFSR_107/D gnd vdd DFFSR
XDFFSR_129 INVX1_138/A DFFSR_60/CLK INVX8_8/Y vdd DFFSR_129/D gnd vdd DFFSR
XDFFSR_118 DFFSR_118/Q CLKBUF1_3/Y INVX8_7/Y vdd NOR2X1_25/B gnd vdd DFFSR
XFILL_20_0_2 gnd vdd FILL
XFILL_3_1_2 gnd vdd FILL
XFILL_11_0_2 gnd vdd FILL
XNAND3X1_62 BUFX4_8/Y gnd DFFSR_66/Q gnd NAND3X1_62/Y vdd NAND3X1
XNAND3X1_51 INVX4_4/A NOR2X1_44/A NAND3X1_39/Y gnd NAND3X1_51/Y vdd NAND3X1
XNAND3X1_40 NAND3X1_40/A NAND3X1_39/Y NOR2X1_47/Y gnd NAND3X1_43/B vdd NAND3X1
XNOR2X1_51 NOR2X1_51/A NOR2X1_50/Y gnd NOR2X1_51/Y vdd NOR2X1
XNOR2X1_40 INVX1_77/Y BUFX4_49/Y gnd NOR2X1_40/Y vdd NOR2X1
XFILL_19_1_2 gnd vdd FILL
XNAND2X1_119 DFFSR_22/Q DFFSR_104/Q gnd OAI21X1_387/C vdd NAND2X1
XNAND2X1_108 OAI21X1_347/Y NAND2X1_108/B gnd DFFSR_69/D vdd NAND2X1
XNAND2X1_6 NOR2X1_4/B DFFSR_88/Q gnd NAND2X1_6/Y vdd NAND2X1
XFILL_21_3_0 gnd vdd FILL
XMUX2X1_80 MUX2X1_94/A MUX2X1_80/B MUX2X1_79/S gnd MUX2X1_80/Y vdd MUX2X1
XMUX2X1_91 INVX1_93/A MUX2X1_97/A MUX2X1_87/S gnd MUX2X1_91/Y vdd MUX2X1
XMUX2X1_114 INVX1_169/Y INVX2_9/Y MUX2X1_118/S gnd DFFSR_160/D vdd MUX2X1
XMUX2X1_103 MUX2X1_97/A MUX2X1_103/B NOR2X1_38/Y gnd MUX2X1_103/Y vdd MUX2X1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XINVX1_76 DFFSR_73/Q gnd INVX1_76/Y vdd INVX1
XBUFX2_18 BUFX2_18/A gnd ext_data_out[12] vdd BUFX2
XDFFPOSX1_6 MUX2X1_26/B DFFSR_89/CLK DFFPOSX1_6/D gnd vdd DFFPOSX1
XINVX1_98 ext_data_in[0] gnd INVX1_98/Y vdd INVX1
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XFILL_12_3_0 gnd vdd FILL
XNOR2X1_9 DFFSR_14/Q INVX2_1/A gnd NOR2X1_9/Y vdd NOR2X1
XOAI21X1_422 DFFSR_132/Q INVX1_141/Y OAI21X1_422/C gnd DFFSR_120/D vdd OAI21X1
XOAI21X1_411 INVX1_135/Y OR2X2_12/Y OAI21X1_410/Y gnd DFFSR_126/D vdd OAI21X1
XOAI21X1_433 INVX1_150/Y OAI21X1_431/Y NOR2X1_51/Y gnd OAI21X1_433/Y vdd OAI21X1
XOAI21X1_455 OAI21X1_455/A OAI21X1_455/B INVX4_3/A gnd NAND2X1_171/B vdd OAI21X1
XOAI21X1_400 INVX1_126/Y OR2X2_11/Y OAI21X1_399/Y gnd DFFSR_115/D vdd OAI21X1
XOAI21X1_444 INVX1_158/Y OAI22X1_6/A MUX2X1_108/S gnd DFFSR_146/D vdd OAI21X1
XFILL_8_0_2 gnd vdd FILL
XOAI21X1_71 OAI21X1_69/Y OAI21X1_71/B NOR2X1_6/Y gnd NAND2X1_18/B vdd OAI21X1
XOAI21X1_93 BUFX4_37/Y MUX2X1_27/Y OAI21X1_93/C gnd OAI21X1_93/Y vdd OAI21X1
XOAI21X1_60 BUFX2_5/Y OR2X2_2/A DFFSR_7/Q gnd OAI21X1_60/Y vdd OAI21X1
XOAI21X1_82 INVX1_24/Y OAI21X1_78/B NAND2X1_23/Y gnd OAI21X1_82/Y vdd OAI21X1
XFILL_1_2_0 gnd vdd FILL
XOAI21X1_274 BUFX4_46/Y MUX2X1_80/Y OAI21X1_274/C gnd OAI21X1_274/Y vdd OAI21X1
XOAI21X1_296 BUFX4_46/Y MUX2X1_89/Y OAI21X1_296/C gnd DFFPOSX1_87/D vdd OAI21X1
XOAI21X1_252 INVX1_68/Y NAND2X1_69/Y NAND2X1_75/Y gnd OAI21X1_252/Y vdd OAI21X1
XOAI21X1_241 OAI21X1_241/A OAI21X1_240/Y NOR2X1_26/Y gnd NAND2X1_70/B vdd OAI21X1
XOAI21X1_230 BUFX4_61/Y BUFX4_15/Y MUX2X1_75/B gnd OAI21X1_231/C vdd OAI21X1
XOAI21X1_263 OR2X2_6/Y NAND2X1_69/Y OAI21X1_262/Y gnd DFFSR_52/D vdd OAI21X1
XOAI21X1_285 BUFX4_20/Y BUFX4_82/Y MUX2X1_84/B gnd OAI21X1_285/Y vdd OAI21X1
XFILL_9_3_0 gnd vdd FILL
XFILL_17_2_0 gnd vdd FILL
XDFFPOSX1_19 MUX2X1_1/B CLKBUF1_4/Y OAI21X1_4/Y gnd vdd DFFPOSX1
XDFFSR_30 DFFSR_30/Q CLKBUF1_34/Y DFFSR_29/R vdd DFFSR_30/D gnd vdd DFFSR
XDFFSR_74 OR2X2_7/B DFFSR_74/CLK DFFSR_74/R vdd XOR2X1_7/Y gnd vdd DFFSR
XDFFSR_63 DFFSR_63/Q DFFSR_61/CLK BUFX4_88/Y vdd DFFSR_63/D gnd vdd DFFSR
XDFFSR_96 DFFSR_96/Q DFFSR_8/CLK INVX8_6/Y vdd DFFSR_96/D gnd vdd DFFSR
XDFFSR_85 DFFSR_85/Q CLKBUF1_40/Y INVX8_5/Y vdd DFFSR_85/D gnd vdd DFFSR
XDFFSR_52 DFFSR_52/Q DFFSR_50/CLK BUFX4_28/Y vdd DFFSR_52/D gnd vdd DFFSR
XDFFSR_41 DFFSR_41/Q DFFSR_50/CLK DFFSR_41/R vdd DFFSR_41/D gnd vdd DFFSR
XINVX1_135 ext_data_in[13] gnd INVX1_135/Y vdd INVX1
XINVX1_124 ext_data_in[10] gnd INVX1_124/Y vdd INVX1
XINVX1_146 BUFX4_58/Y gnd INVX1_146/Y vdd INVX1
XINVX1_113 ext_data_in[7] gnd INVX1_113/Y vdd INVX1
XINVX1_102 DFFSR_87/Q gnd INVX1_102/Y vdd INVX1
XINVX1_157 OAI22X1_6/A gnd DFFSR_171/D vdd INVX1
XINVX1_168 INVX1_51/A gnd INVX1_168/Y vdd INVX1
XINVX1_179 INVX1_34/A gnd INVX1_179/Y vdd INVX1
XFILL_23_0_0 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XDFFSR_119 BUFX2_18/A DFFSR_60/CLK INVX8_8/Y vdd DFFSR_119/D gnd vdd DFFSR
XDFFSR_108 BUFX2_17/A CLKBUF1_24/Y INVX8_7/Y vdd DFFSR_108/D gnd vdd DFFSR
XFILL_14_0_0 gnd vdd FILL
XNOR2X1_30 INVX1_53/Y BUFX4_93/Y gnd NOR2X1_30/Y vdd NOR2X1
XNAND3X1_30 INVX2_7/Y NAND3X1_30/B NAND3X1_30/C gnd NOR2X1_42/B vdd NAND3X1
XNAND3X1_63 gnd DFFSR_48/Q INVX4_4/Y gnd NAND3X1_63/Y vdd NAND3X1
XNAND3X1_52 INVX4_3/A BUFX2_26/A gnd gnd MUX2X1_108/S vdd NAND3X1
XNAND3X1_41 BUFX2_26/A NOR2X1_44/A NAND3X1_39/Y gnd NAND3X1_43/A vdd NAND3X1
XNOR2X1_52 NOR2X1_52/A NOR2X1_52/B gnd NOR2X1_52/Y vdd NOR2X1
XNOR2X1_41 INVX2_6/A INVX4_1/A gnd AOI21X1_9/A vdd NOR2X1
XNAND2X1_109 NAND2X1_109/A NAND2X1_98/B gnd DFFSR_60/D vdd NAND2X1
XNAND2X1_7 OR2X2_1/A OR2X2_1/B gnd NAND2X1_7/Y vdd NAND2X1
XMUX2X1_70 MUX2X1_56/A INVX1_68/A NOR2X1_27/Y gnd MUX2X1_70/Y vdd MUX2X1
XMUX2X1_81 MUX2X1_89/B MUX2X1_81/B MUX2X1_79/S gnd MUX2X1_81/Y vdd MUX2X1
XFILL_21_3_1 gnd vdd FILL
XMUX2X1_92 INVX1_95/A MUX2X1_92/B MUX2X1_87/S gnd MUX2X1_92/Y vdd MUX2X1
XMUX2X1_115 INVX1_170/Y INVX2_10/Y MUX2X1_118/S gnd DFFSR_161/D vdd MUX2X1
XMUX2X1_104 MUX2X1_92/B MUX2X1_104/B NOR2X1_38/Y gnd MUX2X1_104/Y vdd MUX2X1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XINVX1_99 ext_data_in[1] gnd INVX1_99/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XINVX1_77 DFFSR_72/Q gnd INVX1_77/Y vdd INVX1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XBUFX2_19 BUFX2_19/A gnd ext_data_out[13] vdd BUFX2
XDFFPOSX1_7 INVX1_13/A DFFSR_89/CLK DFFPOSX1_7/D gnd vdd DFFPOSX1
XFILL_12_3_1 gnd vdd FILL
XOAI21X1_423 DFFSR_132/Q INVX1_142/Y NAND2X1_131/Y gnd DFFSR_121/D vdd OAI21X1
XOAI21X1_412 BUFX4_21/Y BUFX2_25/A DFFSR_127/Q gnd OAI21X1_412/Y vdd OAI21X1
XOAI21X1_434 DFFSR_137/D NOR2X1_46/A INVX4_1/A gnd OAI21X1_434/Y vdd OAI21X1
XOAI21X1_445 INVX1_159/Y OAI22X1_6/A MUX2X1_122/S gnd DFFSR_144/D vdd OAI21X1
XOAI21X1_456 INVX1_182/Y OR2X2_14/Y NAND3X1_60/Y gnd OAI21X1_456/Y vdd OAI21X1
XOAI21X1_401 BUFX4_61/Y BUFX2_24/A INVX1_127/A gnd OAI21X1_401/Y vdd OAI21X1
XOAI21X1_94 DFFSR_95/Q INVX1_30/Y NAND2X1_30/Y gnd MUX2X1_42/A vdd OAI21X1
XOAI21X1_50 BUFX4_76/Y BUFX4_43/Y MUX2X1_22/B gnd OAI21X1_50/Y vdd OAI21X1
XOAI21X1_61 INVX1_12/Y OAI21X1_69/B NAND3X1_2/Y gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_83 OAI21X1_81/Y OAI21X1_82/Y NOR2X1_6/Y gnd OAI21X1_83/Y vdd OAI21X1
XOAI21X1_72 OR2X2_2/B OR2X2_2/A DFFSR_10/Q gnd NAND2X1_20/A vdd OAI21X1
XFILL_1_2_1 gnd vdd FILL
XOAI21X1_220 BUFX4_65/Y BUFX4_16/Y INVX1_68/A gnd OAI21X1_221/C vdd OAI21X1
XOAI21X1_297 BUFX4_22/Y BUFX4_81/Y INVX1_91/A gnd OAI21X1_297/Y vdd OAI21X1
XOAI21X1_242 BUFX2_2/Y OR2X2_6/A DFFSR_46/Q gnd NAND2X1_72/A vdd OAI21X1
XOAI21X1_275 DFFSR_123/Q INVX1_79/Y NAND2X1_87/Y gnd MUX2X1_89/B vdd OAI21X1
XOAI21X1_253 OAI21X1_253/A OAI21X1_252/Y NOR2X1_26/Y gnd NAND2X1_76/B vdd OAI21X1
XOAI21X1_231 BUFX4_94/Y MUX2X1_75/Y OAI21X1_231/C gnd DFFPOSX1_51/D vdd OAI21X1
XOAI21X1_264 OR2X2_6/B OR2X2_6/A DFFSR_41/Q gnd NAND2X1_81/A vdd OAI21X1
XOAI21X1_286 BUFX4_49/Y MUX2X1_84/Y OAI21X1_285/Y gnd OAI21X1_286/Y vdd OAI21X1
XFILL_9_3_1 gnd vdd FILL
XFILL_17_2_1 gnd vdd FILL
XDFFSR_53 DFFSR_53/Q CLKBUF1_5/Y DFFSR_54/R vdd DFFSR_53/D gnd vdd DFFSR
XDFFSR_64 DFFSR_64/Q CLKBUF1_5/Y BUFX4_88/Y vdd DFFSR_64/D gnd vdd DFFSR
XDFFSR_31 DFFSR_31/Q CLKBUF1_34/Y DFFSR_29/R vdd DFFSR_31/D gnd vdd DFFSR
XDFFSR_20 DFFSR_20/Q DFFSR_33/CLK DFFSR_38/R vdd DFFSR_20/D gnd vdd DFFSR
XDFFSR_42 DFFSR_42/Q CLKBUF1_3/Y DFFSR_43/R vdd DFFSR_42/D gnd vdd DFFSR
XDFFSR_75 OR2X2_7/A DFFSR_74/CLK DFFSR_74/R vdd DFFSR_75/D gnd vdd DFFSR
XDFFSR_97 DFFSR_97/Q CLKBUF1_13/Y INVX8_6/Y vdd DFFSR_97/D gnd vdd DFFSR
XDFFSR_86 DFFSR_86/Q CLKBUF1_4/Y INVX8_5/Y vdd DFFSR_86/D gnd vdd DFFSR
XCLKBUF1_40 BUFX4_1/Y gnd CLKBUF1_40/Y vdd CLKBUF1
XINVX1_125 ext_data_in[11] gnd INVX1_125/Y vdd INVX1
XINVX1_136 ext_data_in[14] gnd INVX1_136/Y vdd INVX1
XINVX1_147 BUFX2_4/Y gnd OAI22X1_4/A vdd INVX1
XINVX1_114 INVX1_114/A gnd INVX1_114/Y vdd INVX1
XINVX1_103 DFFSR_88/Q gnd INVX1_103/Y vdd INVX1
XINVX1_169 INVX1_54/A gnd INVX1_169/Y vdd INVX1
XINVX1_158 NOR2X1_34/A gnd INVX1_158/Y vdd INVX1
XFILL_23_0_1 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XDFFSR_109 DFFSR_109/Q CLKBUF1_26/Y INVX8_7/Y vdd INVX1_121/Y gnd vdd DFFSR
XFILL_25_1 gnd vdd FILL
XNOR2X1_53 NOR2X1_53/A NOR2X1_52/Y gnd NOR2X1_53/Y vdd NOR2X1
XNOR2X1_31 DFFSR_76/Q OR2X2_7/Y gnd DFFSR_59/D vdd NOR2X1
XNAND3X1_31 INVX2_6/A BUFX4_25/Y INVX4_1/Y gnd NAND3X1_33/B vdd NAND3X1
XNOR2X1_42 OAI22X1_1/Y NOR2X1_42/B gnd AOI21X1_8/C vdd NOR2X1
XNOR2X1_20 INVX1_29/Y BUFX4_38/Y gnd NOR2X1_20/Y vdd NOR2X1
XNAND3X1_64 BUFX2_1/Y DFFSR_29/Q INVX4_5/Y gnd NAND3X1_64/Y vdd NAND3X1
XNAND3X1_53 INVX4_3/A BUFX2_26/A INVX1_160/Y gnd MUX2X1_122/S vdd NAND3X1
XNAND3X1_42 NAND3X1_42/A NAND3X1_42/B AOI22X1_4/Y gnd AOI22X1_5/C vdd NAND3X1
XNAND3X1_20 MUX2X1_57/B DFFSR_52/Q INVX2_3/A gnd NAND3X1_20/Y vdd NAND3X1
XNAND2X1_8 INVX1_1/A NAND2X1_7/Y gnd NAND2X1_8/Y vdd NAND2X1
XMUX2X1_71 MUX2X1_71/A INVX1_70/A NOR2X1_27/Y gnd MUX2X1_71/Y vdd MUX2X1
XMUX2X1_82 MUX2X1_82/A MUX2X1_82/B MUX2X1_79/S gnd MUX2X1_82/Y vdd MUX2X1
XMUX2X1_93 MUX2X1_79/A INVX1_85/A NOR2X1_37/Y gnd MUX2X1_93/Y vdd MUX2X1
XMUX2X1_60 MUX2X1_59/Y XOR2X1_6/Y OR2X2_6/Y gnd DFFSR_56/D vdd MUX2X1
XFILL_21_3_2 gnd vdd FILL
XMUX2X1_105 BUFX4_21/Y BUFX4_31/Y DFFSR_135/Q gnd MUX2X1_105/Y vdd MUX2X1
XMUX2X1_116 INVX1_171/Y INVX2_11/Y MUX2X1_118/S gnd DFFSR_162/D vdd MUX2X1
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XDFFPOSX1_8 INVX1_16/A DFFSR_89/CLK OAI21X1_39/Y gnd vdd DFFPOSX1
XFILL_12_3_2 gnd vdd FILL
XOAI21X1_424 DFFSR_132/Q INVX1_143/Y OAI21X1_424/C gnd DFFSR_122/D vdd OAI21X1
XOAI21X1_413 INVX1_136/Y OR2X2_12/Y OAI21X1_412/Y gnd DFFSR_127/D vdd OAI21X1
XOAI21X1_435 OAI21X1_433/Y AOI21X1_8/Y OAI21X1_434/Y gnd DFFSR_139/D vdd OAI21X1
XOAI21X1_446 INVX4_3/Y OR2X2_13/Y NAND2X1_161/Y gnd DFFSR_143/D vdd OAI21X1
XOAI21X1_457 OAI21X1_457/A OAI21X1_456/Y INVX4_3/A gnd NAND2X1_174/B vdd OAI21X1
XOAI21X1_402 INVX1_127/Y OR2X2_11/Y OAI21X1_401/Y gnd DFFSR_116/D vdd OAI21X1
XOAI21X1_51 AND2X2_1/A MUX2X1_22/Y OAI21X1_50/Y gnd OAI21X1_51/Y vdd OAI21X1
XOAI21X1_73 INVX1_19/Y OAI21X1_69/B NAND3X1_5/Y gnd OAI21X1_75/A vdd OAI21X1
XOAI21X1_62 INVX1_13/Y OAI21X1_78/B NAND2X1_12/Y gnd OAI21X1_62/Y vdd OAI21X1
XOAI21X1_95 BUFX4_32/Y BUFX4_55/Y MUX2X1_28/B gnd OAI21X1_95/Y vdd OAI21X1
XOAI21X1_84 INVX2_1/Y OR2X2_2/Y DFFSR_14/Q gnd OAI21X1_84/Y vdd OAI21X1
XOAI21X1_40 BUFX4_73/Y BUFX4_41/Y INVX1_18/A gnd OAI21X1_40/Y vdd OAI21X1
XFILL_1_2_2 gnd vdd FILL
XOAI21X1_221 BUFX4_96/Y MUX2X1_70/Y OAI21X1_221/C gnd DFFPOSX1_58/D vdd OAI21X1
XOAI21X1_210 BUFX4_64/Y BUFX4_18/Y INVX1_69/A gnd OAI21X1_210/Y vdd OAI21X1
XOAI21X1_287 OR2X2_8/B OR2X2_8/A AND2X2_4/A gnd XOR2X1_7/A vdd OAI21X1
XOAI21X1_298 BUFX4_47/Y MUX2X1_90/Y OAI21X1_297/Y gnd DFFPOSX1_88/D vdd OAI21X1
XOAI21X1_276 BUFX4_19/Y BUFX4_81/Y MUX2X1_81/B gnd OAI21X1_277/C vdd OAI21X1
XOAI21X1_265 BUFX2_2/Y OR2X2_6/A DFFSR_42/Q gnd NAND2X1_82/A vdd OAI21X1
XOAI21X1_243 INVX1_63/Y NAND2X1_67/Y NAND3X1_17/Y gnd OAI21X1_243/Y vdd OAI21X1
XOAI21X1_232 BUFX4_63/Y BUFX4_17/Y MUX2X1_76/B gnd OAI21X1_232/Y vdd OAI21X1
XOAI21X1_254 OR2X2_6/B OR2X2_6/A DFFSR_49/Q gnd NAND2X1_78/A vdd OAI21X1
XFILL_9_3_2 gnd vdd FILL
XFILL_17_2_2 gnd vdd FILL
XDFFSR_76 DFFSR_76/Q DFFSR_74/CLK DFFSR_74/R vdd DFFSR_76/D gnd vdd DFFSR
XDFFSR_54 DFFSR_54/Q DFFSR_54/CLK DFFSR_54/R vdd DFFSR_54/D gnd vdd DFFSR
XDFFSR_98 DFFSR_98/Q CLKBUF1_13/Y INVX8_6/Y vdd DFFSR_98/D gnd vdd DFFSR
XDFFSR_87 DFFSR_87/Q DFFSR_87/CLK INVX8_5/Y vdd DFFSR_87/D gnd vdd DFFSR
XDFFSR_10 DFFSR_10/Q DFFSR_2/CLK DFFSR_2/S vdd DFFSR_10/D gnd vdd DFFSR
XDFFSR_32 INVX2_2/A DFFSR_33/CLK DFFSR_38/R vdd DFFSR_32/D gnd vdd DFFSR
XDFFSR_21 BUFX2_3/A DFFSR_21/CLK vdd DFFSR_38/R DFFSR_21/D gnd vdd DFFSR
XDFFSR_43 DFFSR_43/Q CLKBUF1_3/Y DFFSR_43/R vdd DFFSR_43/D gnd vdd DFFSR
XDFFSR_65 DFFSR_65/Q DFFSR_67/CLK DFFSR_69/R vdd DFFSR_65/D gnd vdd DFFSR
XCLKBUF1_41 BUFX4_5/Y gnd CLKBUF1_41/Y vdd CLKBUF1
XCLKBUF1_30 BUFX4_6/Y gnd CLKBUF1_30/Y vdd CLKBUF1
XINVX1_137 ext_data_in[15] gnd INVX1_137/Y vdd INVX1
XINVX1_148 BUFX2_26/A gnd INVX1_148/Y vdd INVX1
XINVX1_115 DFFSR_102/Q gnd INVX1_115/Y vdd INVX1
XINVX1_104 BUFX2_6/A gnd INVX1_104/Y vdd INVX1
XINVX1_159 INVX1_159/A gnd INVX1_159/Y vdd INVX1
XINVX1_126 INVX1_126/A gnd INVX1_126/Y vdd INVX1
XFILL_23_0_2 gnd vdd FILL
XFILL_6_1_2 gnd vdd FILL
XFILL_14_0_2 gnd vdd FILL
XFILL_25_2 gnd vdd FILL
XFILL_18_1 gnd vdd FILL
XFILL_24_3_0 gnd vdd FILL
XNAND3X1_32 BUFX4_58/Y INVX2_6/Y INVX4_1/Y gnd NAND3X1_33/C vdd NAND3X1
XNAND3X1_21 MUX2X1_58/B DFFSR_52/Q INVX2_3/A gnd NAND3X1_21/Y vdd NAND3X1
XNAND3X1_10 MUX2X1_28/B DFFSR_33/Q INVX2_2/A gnd NAND3X1_10/Y vdd NAND3X1
XNOR2X1_32 INVX1_73/Y OR2X2_7/Y gnd DFFSR_58/D vdd NOR2X1
XNOR2X1_43 OAI22X1_2/Y NOR2X1_43/B gnd AOI21X1_7/C vdd NOR2X1
XNOR2X1_21 DFFSR_57/Q OR2X2_5/Y gnd DFFSR_40/D vdd NOR2X1
XNOR2X1_10 INVX1_5/Y BUFX4_11/Y gnd NOR2X1_10/Y vdd NOR2X1
XNOR2X1_54 BUFX2_26/A INVX1_160/Y gnd NOR2X1_54/Y vdd NOR2X1
XNAND3X1_65 BUFX2_1/Y gnd DFFSR_67/Q gnd NAND3X1_65/Y vdd NAND3X1
XNAND3X1_54 gnd DFFSR_45/Q INVX4_4/Y gnd NAND3X1_54/Y vdd NAND3X1
XNAND3X1_43 NAND3X1_43/A NAND3X1_43/B AOI22X1_5/Y gnd AOI22X1_8/D vdd NAND3X1
XFILL_15_3_0 gnd vdd FILL
XNAND2X1_9 NAND2X1_9/A NAND2X1_9/B gnd DFFSR_19/D vdd NAND2X1
XMUX2X1_72 MUX2X1_66/B INVX1_72/A NOR2X1_27/Y gnd MUX2X1_72/Y vdd MUX2X1
XMUX2X1_61 INVX1_60/A MUX2X1_53/A MUX2X1_66/S gnd MUX2X1_61/Y vdd MUX2X1
XMUX2X1_50 MUX2X1_44/A MUX2X1_50/B NOR2X1_18/Y gnd MUX2X1_50/Y vdd MUX2X1
XMUX2X1_94 MUX2X1_94/A INVX1_88/A NOR2X1_37/Y gnd MUX2X1_94/Y vdd MUX2X1
XMUX2X1_83 MUX2X1_97/A MUX2X1_83/B MUX2X1_79/S gnd MUX2X1_83/Y vdd MUX2X1
XMUX2X1_106 BUFX4_64/Y INVX1_2/A DFFSR_135/Q gnd MUX2X1_106/Y vdd MUX2X1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XMUX2X1_117 INVX1_172/Y INVX2_12/Y MUX2X1_118/S gnd DFFSR_163/D vdd MUX2X1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XDFFPOSX1_9 INVX1_18/A DFFSR_87/CLK OAI21X1_41/Y gnd vdd DFFPOSX1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XOAI21X1_403 BUFX4_65/Y DFFSR_109/Q OAI21X1_403/C gnd DFFSR_117/D vdd OAI21X1
XFILL_21_1_0 gnd vdd FILL
XOAI21X1_414 BUFX4_21/Y BUFX2_25/A DFFSR_128/Q gnd OAI21X1_414/Y vdd OAI21X1
XOAI21X1_425 INVX4_1/A INVX2_5/Y OAI21X1_425/C gnd OAI21X1_425/Y vdd OAI21X1
XOAI21X1_458 INVX1_183/Y OR2X2_14/Y NAND3X1_63/Y gnd OAI21X1_458/Y vdd OAI21X1
XOAI21X1_447 INVX4_4/Y INVX4_5/Y DFFSR_142/Q gnd OAI22X1_6/D vdd OAI21X1
XOAI21X1_436 OAI21X1_436/A INVX1_155/Y DFFSR_137/Q gnd OAI21X1_437/A vdd OAI21X1
XFILL_4_2_0 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XOAI21X1_30 BUFX4_73/Y BUFX4_42/Y INVX1_19/A gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_63 OAI21X1_61/Y OAI21X1_62/Y NOR2X1_6/Y gnd NAND2X1_14/B vdd OAI21X1
XOAI21X1_52 BUFX4_73/Y BUFX4_44/Y MUX2X1_23/B gnd OAI21X1_52/Y vdd OAI21X1
XOAI21X1_41 MUX2X1_7/S MUX2X1_17/Y OAI21X1_40/Y gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_74 INVX1_20/Y OAI21X1_78/B NAND2X1_19/Y gnd OAI21X1_74/Y vdd OAI21X1
XOAI21X1_96 BUFX4_40/Y MUX2X1_28/Y OAI21X1_95/Y gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_85 OR2X2_2/Y OAI21X1_78/B OAI21X1_84/Y gnd DFFSR_14/D vdd OAI21X1
XOAI21X1_200 OR2X2_5/A OR2X2_5/B DFFSR_57/Q gnd INVX1_59/A vdd OAI21X1
XOAI21X1_211 BUFX4_93/Y MUX2X1_65/Y OAI21X1_210/Y gnd OAI21X1_211/Y vdd OAI21X1
XOAI21X1_222 BUFX4_64/Y BUFX4_18/Y INVX1_70/A gnd OAI21X1_222/Y vdd OAI21X1
XOAI21X1_233 BUFX4_94/Y MUX2X1_76/Y OAI21X1_232/Y gnd DFFPOSX1_52/D vdd OAI21X1
XOAI21X1_244 INVX1_64/Y NAND2X1_69/Y NAND2X1_71/Y gnd OAI21X1_245/B vdd OAI21X1
XOAI21X1_255 INVX1_69/Y NAND2X1_67/Y NAND3X1_20/Y gnd OAI21X1_257/A vdd OAI21X1
XOAI21X1_288 AND2X2_4/Y AOI21X1_4/Y OR2X2_8/Y gnd NAND2X1_93/B vdd OAI21X1
XOAI21X1_266 BUFX2_2/Y OR2X2_6/A DFFSR_43/Q gnd NAND2X1_83/A vdd OAI21X1
XOAI21X1_277 BUFX4_46/Y MUX2X1_81/Y OAI21X1_277/C gnd DFFPOSX1_93/D vdd OAI21X1
XOAI21X1_299 BUFX4_19/Y BUFX4_83/Y INVX1_93/A gnd OAI21X1_300/C vdd OAI21X1
XDFFSR_77 BUFX2_6/A DFFSR_9/CLK INVX8_5/Y vdd DFFSR_77/D gnd vdd DFFSR
XDFFSR_99 DFFSR_99/Q CLKBUF1_13/Y INVX8_6/Y vdd DFFSR_99/D gnd vdd DFFSR
XDFFSR_22 DFFSR_22/Q CLKBUF1_16/Y BUFX4_78/Y vdd DFFSR_22/D gnd vdd DFFSR
XDFFSR_33 DFFSR_33/Q DFFSR_33/CLK DFFSR_38/R vdd DFFSR_33/D gnd vdd DFFSR
XDFFSR_11 DFFSR_11/Q CLKBUF1_35/Y DFFSR_8/R vdd DFFSR_11/D gnd vdd DFFSR
XDFFSR_88 DFFSR_88/Q CLKBUF1_40/Y INVX8_5/Y vdd DFFSR_88/D gnd vdd DFFSR
XDFFSR_44 DFFSR_44/Q CLKBUF1_3/Y BUFX4_28/Y vdd DFFSR_44/D gnd vdd DFFSR
XDFFSR_55 OR2X2_5/B DFFSR_50/CLK DFFSR_41/R vdd DFFSR_55/D gnd vdd DFFSR
XDFFSR_66 DFFSR_66/Q DFFSR_67/CLK DFFSR_69/R vdd DFFSR_66/D gnd vdd DFFSR
XCLKBUF1_20 BUFX4_3/Y gnd CLKBUF1_20/Y vdd CLKBUF1
XCLKBUF1_31 BUFX4_1/Y gnd CLKBUF1_31/Y vdd CLKBUF1
XCLKBUF1_42 BUFX4_3/Y gnd CLKBUF1_42/Y vdd CLKBUF1
XFILL_1_0_0 gnd vdd FILL
XINVX1_105 BUFX2_7/A gnd INVX1_105/Y vdd INVX1
XINVX1_116 BUFX2_10/A gnd INVX1_116/Y vdd INVX1
XINVX1_149 BUFX4_25/Y gnd OAI22X1_3/A vdd INVX1
XINVX1_138 INVX1_138/A gnd INVX1_138/Y vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XINVX1_127 INVX1_127/A gnd INVX1_127/Y vdd INVX1
XFILL_17_0_0 gnd vdd FILL
XFILL_18_2 gnd vdd FILL
XFILL_24_3_1 gnd vdd FILL
XNAND3X1_22 OR2X2_7/A OR2X2_7/B INVX1_73/Y gnd AOI21X1_4/B vdd NAND3X1
XNAND3X1_33 INVX2_7/Y NAND3X1_33/B NAND3X1_33/C gnd NOR2X1_43/B vdd NAND3X1
XNAND3X1_11 MUX2X1_29/B DFFSR_33/Q INVX2_2/A gnd NAND3X1_11/Y vdd NAND3X1
XNAND3X1_55 BUFX4_9/Y DFFSR_26/Q INVX4_5/Y gnd NAND3X1_55/Y vdd NAND3X1
XNAND3X1_66 gnd DFFSR_49/Q INVX4_4/Y gnd NAND3X1_66/Y vdd NAND3X1
XNAND3X1_44 AOI22X1_6/Y AOI22X1_7/Y AOI21X1_8/C gnd AOI22X1_8/C vdd NAND3X1
XNOR2X1_44 NOR2X1_44/A AOI21X1_7/C gnd NOR2X1_44/Y vdd NOR2X1
XNOR2X1_22 INVX1_49/Y OR2X2_5/Y gnd DFFSR_39/D vdd NOR2X1
XNOR2X1_55 INVX4_3/Y OR2X2_13/Y gnd NOR2X1_58/B vdd NOR2X1
XNOR2X1_11 INVX1_25/A OR2X2_3/Y gnd DFFSR_21/D vdd NOR2X1
XFILL_15_3_1 gnd vdd FILL
XNOR2X1_33 INVX1_76/Y INVX1_77/Y gnd MUX2X1_79/S vdd NOR2X1
XMUX2X1_40 INVX1_47/A MUX2X1_46/A MUX2X1_39/S gnd MUX2X1_40/Y vdd MUX2X1
XMUX2X1_51 MUX2X1_39/B MUX2X1_51/B NOR2X1_18/Y gnd MUX2X1_51/Y vdd MUX2X1
XMUX2X1_95 MUX2X1_89/B INVX1_90/A NOR2X1_37/Y gnd MUX2X1_95/Y vdd MUX2X1
XMUX2X1_84 MUX2X1_92/B MUX2X1_84/B MUX2X1_79/S gnd MUX2X1_84/Y vdd MUX2X1
XMUX2X1_73 MUX2X1_53/A MUX2X1_73/B NOR2X1_28/Y gnd MUX2X1_73/Y vdd MUX2X1
XMUX2X1_62 INVX1_63/A MUX2X1_68/A MUX2X1_66/S gnd MUX2X1_62/Y vdd MUX2X1
XMUX2X1_118 INVX1_173/Y INVX2_13/Y MUX2X1_118/S gnd DFFSR_164/D vdd MUX2X1
XMUX2X1_107 INVX1_162/Y INVX2_8/Y MUX2X1_108/S gnd DFFSR_165/D vdd MUX2X1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XINVX1_14 DFFSR_14/Q gnd INVX1_14/Y vdd INVX1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XOAI21X1_426 INVX4_1/A INVX1_146/Y OAI21X1_426/C gnd NAND2X1_139/B vdd OAI21X1
XOAI21X1_404 DFFSR_118/Q INVX1_128/Y NAND2X1_124/Y gnd DFFSR_105/D vdd OAI21X1
XFILL_21_1_1 gnd vdd FILL
XOAI21X1_415 INVX1_137/Y OR2X2_12/Y OAI21X1_414/Y gnd DFFSR_128/D vdd OAI21X1
XOAI21X1_448 gnd INVX4_4/Y NOR2X1_15/A gnd OAI22X1_7/D vdd OAI21X1
XOAI21X1_437 OAI21X1_437/A AOI22X1_8/Y OAI21X1_437/C gnd DFFSR_134/D vdd OAI21X1
XOAI21X1_459 NAND2X1_175/Y OAI21X1_458/Y INVX4_3/A gnd OAI21X1_459/Y vdd OAI21X1
XFILL_4_2_1 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XOAI21X1_86 BUFX2_5/Y OR2X2_2/A DFFSR_3/Q gnd OAI21X1_86/Y vdd OAI21X1
XOAI21X1_20 BUFX4_97/Y OR2X2_2/A AND2X2_1/A gnd XOR2X1_1/A vdd OAI21X1
XOAI21X1_31 BUFX4_14/Y MUX2X1_12/Y OAI21X1_30/Y gnd OAI21X1_31/Y vdd OAI21X1
XOAI21X1_75 OAI21X1_75/A OAI21X1_74/Y NOR2X1_6/Y gnd NAND2X1_20/B vdd OAI21X1
XOAI21X1_42 BUFX4_74/Y BUFX4_42/Y INVX1_20/A gnd OAI21X1_42/Y vdd OAI21X1
XOAI21X1_64 BUFX2_5/Y OR2X2_2/A DFFSR_8/Q gnd NAND2X1_16/A vdd OAI21X1
XOAI21X1_53 BUFX4_10/Y MUX2X1_23/Y OAI21X1_52/Y gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_97 DFFSR_95/Q INVX1_31/Y NAND2X1_31/Y gnd MUX2X1_49/A vdd OAI21X1
XOAI21X1_289 OR2X2_7/A OR2X2_7/B DFFSR_76/Q gnd INVX1_83/A vdd OAI21X1
XOAI21X1_212 BUFX4_62/Y BUFX4_15/Y INVX1_71/A gnd OAI21X1_212/Y vdd OAI21X1
XOAI21X1_223 BUFX4_93/Y MUX2X1_71/Y OAI21X1_222/Y gnd OAI21X1_223/Y vdd OAI21X1
XOAI21X1_201 INVX1_59/Y DFFSR_40/D NOR2X1_26/Y gnd NAND2X1_65/A vdd OAI21X1
XOAI21X1_234 BUFX4_64/Y BUFX4_18/Y MUX2X1_77/B gnd OAI21X1_234/Y vdd OAI21X1
XOAI21X1_267 BUFX4_26/Y OR2X2_6/A DFFSR_44/Q gnd NAND2X1_84/A vdd OAI21X1
XOAI21X1_278 DFFSR_123/Q INVX1_80/Y NAND2X1_88/Y gnd MUX2X1_82/A vdd OAI21X1
XOAI21X1_245 OAI21X1_243/Y OAI21X1_245/B NOR2X1_26/Y gnd NAND2X1_72/B vdd OAI21X1
XOAI21X1_256 INVX1_70/Y NAND2X1_69/Y NAND2X1_77/Y gnd OAI21X1_257/B vdd OAI21X1
XDFFSR_12 DFFSR_12/Q CLKBUF1_35/Y DFFSR_2/S vdd DFFSR_12/D gnd vdd DFFSR
XDFFSR_56 OR2X2_5/A DFFSR_54/CLK DFFSR_54/R vdd DFFSR_56/D gnd vdd DFFSR
XDFFSR_67 DFFSR_67/Q DFFSR_67/CLK DFFSR_69/R vdd DFFSR_67/D gnd vdd DFFSR
XDFFSR_23 DFFSR_23/Q DFFSR_23/CLK BUFX4_78/Y vdd DFFSR_23/D gnd vdd DFFSR
XDFFSR_89 OR2X2_9/B DFFSR_89/CLK INVX8_5/Y vdd DFFSR_89/D gnd vdd DFFSR
XDFFSR_78 BUFX2_7/A DFFSR_1/CLK INVX8_5/Y vdd DFFSR_78/D gnd vdd DFFSR
XDFFSR_34 DFFSR_34/Q DFFSR_36/CLK DFFSR_34/R vdd DFFSR_34/D gnd vdd DFFSR
XDFFSR_45 DFFSR_45/Q DFFSR_45/CLK BUFX4_28/Y vdd DFFSR_45/D gnd vdd DFFSR
XCLKBUF1_32 BUFX4_2/Y gnd CLKBUF1_32/Y vdd CLKBUF1
XCLKBUF1_21 BUFX4_5/Y gnd CLKBUF1_21/Y vdd CLKBUF1
XCLKBUF1_10 BUFX4_4/Y gnd DFFSR_89/CLK vdd CLKBUF1
XFILL_1_0_1 gnd vdd FILL
XINVX1_128 BUFX2_14/A gnd INVX1_128/Y vdd INVX1
XINVX1_139 DFFSR_130/Q gnd INVX1_139/Y vdd INVX1
XINVX1_106 BUFX2_8/A gnd INVX1_106/Y vdd INVX1
XINVX1_117 DFFSR_92/Q gnd INVX1_117/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XFILL_18_3 gnd vdd FILL
XFILL_24_3_2 gnd vdd FILL
XNAND3X1_34 INVX2_7/Y NAND3X1_34/B NAND3X1_34/C gnd NOR2X1_44/A vdd NAND3X1
XNAND3X1_23 MUX2X1_79/B DFFSR_71/Q INVX2_4/A gnd NAND3X1_23/Y vdd NAND3X1
XNAND3X1_12 MUX2X1_30/B DFFSR_33/Q INVX2_2/A gnd NAND3X1_12/Y vdd NAND3X1
XNOR2X1_12 INVX1_25/Y OR2X2_3/Y gnd DFFSR_20/D vdd NOR2X1
XNAND3X1_67 INVX4_4/A DFFSR_30/Q INVX4_5/Y gnd NAND3X1_67/Y vdd NAND3X1
XNAND3X1_56 BUFX4_8/Y gnd DFFSR_64/Q gnd NAND3X1_56/Y vdd NAND3X1
XNAND3X1_45 NAND3X1_45/A NAND3X1_45/B NAND3X1_45/C gnd NAND3X1_45/Y vdd NAND3X1
XNOR2X1_23 INVX1_52/Y INVX1_53/Y gnd NOR2X1_23/Y vdd NOR2X1
XNOR2X1_45 OAI22X1_3/Y NOR2X1_45/B gnd NOR2X1_46/A vdd NOR2X1
XNOR2X1_56 INVX1_3/A NOR2X1_58/B gnd NOR2X1_56/Y vdd NOR2X1
XNOR2X1_34 NOR2X1_34/A DFFSR_123/Q gnd BUFX4_82/A vdd NOR2X1
XFILL_15_3_2 gnd vdd FILL
XMUX2X1_30 MUX2X1_44/A MUX2X1_30/B NOR2X1_13/Y gnd MUX2X1_30/Y vdd MUX2X1
XMUX2X1_52 MUX2X1_46/A MUX2X1_52/B NOR2X1_18/Y gnd MUX2X1_52/Y vdd MUX2X1
XMUX2X1_41 MUX2X1_41/A INVX1_37/A MUX2X1_43/S gnd MUX2X1_41/Y vdd MUX2X1
XMUX2X1_63 INVX1_65/A MUX2X1_55/A MUX2X1_66/S gnd MUX2X1_63/Y vdd MUX2X1
XMUX2X1_85 OR2X2_7/A XOR2X1_8/Y AND2X2_4/A gnd MUX2X1_85/Y vdd MUX2X1
XFILL_23_1 gnd vdd FILL
XMUX2X1_96 MUX2X1_82/A INVX1_92/A NOR2X1_37/Y gnd MUX2X1_96/Y vdd MUX2X1
XMUX2X1_74 MUX2X1_68/A MUX2X1_74/B NOR2X1_28/Y gnd MUX2X1_74/Y vdd MUX2X1
XMUX2X1_119 INVX1_174/Y INVX2_8/Y MUX2X1_122/S gnd DFFSR_153/D vdd MUX2X1
XMUX2X1_108 INVX1_163/Y INVX2_9/Y MUX2X1_108/S gnd DFFSR_166/D vdd MUX2X1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XINVX1_26 BUFX4_31/Y gnd INVX1_26/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XOAI21X1_427 INVX2_5/Y OAI21X1_427/B AOI21X1_5/Y gnd NOR2X1_45/B vdd OAI21X1
XFILL_21_1_2 gnd vdd FILL
XOAI21X1_416 BUFX4_21/Y BUFX2_25/A INVX1_138/A gnd OAI21X1_416/Y vdd OAI21X1
XOAI21X1_449 BUFX4_9/Y gnd NOR2X1_5/A gnd OAI22X1_8/B vdd OAI21X1
XOAI21X1_405 DFFSR_118/Q INVX1_129/Y NAND2X1_125/Y gnd DFFSR_106/D vdd OAI21X1
XOAI21X1_438 NAND2X1_157/Y INVX1_155/Y DFFSR_137/Q gnd OAI21X1_438/Y vdd OAI21X1
XFILL_4_2_2 gnd vdd FILL
XFILL_12_1_2 gnd vdd FILL
XOAI21X1_54 BUFX4_74/Y BUFX4_42/Y MUX2X1_24/B gnd OAI21X1_55/C vdd OAI21X1
XOAI21X1_43 BUFX4_14/Y MUX2X1_18/Y OAI21X1_42/Y gnd OAI21X1_43/Y vdd OAI21X1
XOAI21X1_98 BUFX4_32/Y BUFX4_56/Y MUX2X1_29/B gnd OAI21X1_99/C vdd OAI21X1
XOAI21X1_10 BUFX4_11/Y MUX2X1_3/Y OAI21X1_9/Y gnd OAI21X1_10/Y vdd OAI21X1
XOAI21X1_65 INVX1_15/Y OAI21X1_69/B NAND3X1_3/Y gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_21 AND2X2_1/Y AOI21X1_1/Y OR2X2_2/Y gnd NAND2X1_9/B vdd OAI21X1
XOAI21X1_87 BUFX4_97/Y OR2X2_2/A DFFSR_4/Q gnd OAI21X1_87/Y vdd OAI21X1
XOAI21X1_32 INVX1_2/A BUFX4_41/Y INVX1_21/A gnd OAI21X1_33/C vdd OAI21X1
XOAI21X1_76 OR2X2_2/B OR2X2_2/A DFFSR_11/Q gnd NAND2X1_22/A vdd OAI21X1
XOAI21X1_213 BUFX4_92/Y MUX2X1_66/Y OAI21X1_212/Y gnd OAI21X1_213/Y vdd OAI21X1
XOAI21X1_224 BUFX4_65/Y BUFX4_16/Y INVX1_72/A gnd OAI21X1_224/Y vdd OAI21X1
XOAI21X1_235 BUFX4_93/Y MUX2X1_77/Y OAI21X1_234/Y gnd DFFPOSX1_53/D vdd OAI21X1
XOAI21X1_246 BUFX4_26/Y OR2X2_6/A DFFSR_47/Q gnd NAND2X1_74/A vdd OAI21X1
XOAI21X1_268 NOR2X1_34/A DFFSR_123/Q INVX1_74/Y gnd BUFX4_48/A vdd OAI21X1
XOAI21X1_279 BUFX4_20/Y BUFX4_81/Y MUX2X1_82/B gnd OAI21X1_279/Y vdd OAI21X1
XOAI21X1_257 OAI21X1_257/A OAI21X1_257/B NOR2X1_26/Y gnd NAND2X1_78/B vdd OAI21X1
XOAI21X1_202 BUFX4_63/Y BUFX4_17/Y INVX1_60/A gnd OAI21X1_202/Y vdd OAI21X1
XDFFSR_24 DFFSR_24/Q CLKBUF1_16/Y BUFX4_78/Y vdd DFFSR_24/D gnd vdd DFFSR
XDFFSR_13 INVX2_1/A DFFSR_1/CLK DFFSR_5/R vdd DFFSR_13/D gnd vdd DFFSR
XDFFSR_35 INVX1_28/A CLKBUF1_42/Y DFFSR_34/R vdd DFFSR_35/D gnd vdd DFFSR
XDFFSR_46 DFFSR_46/Q CLKBUF1_3/Y DFFSR_43/R vdd DFFSR_46/D gnd vdd DFFSR
XDFFSR_57 DFFSR_57/Q DFFSR_54/CLK DFFSR_54/R vdd DFFSR_57/D gnd vdd DFFSR
XCLKBUF1_33 BUFX4_2/Y gnd DFFSR_61/CLK vdd CLKBUF1
XDFFSR_79 BUFX2_8/A DFFSR_9/CLK INVX8_5/Y vdd DFFSR_79/D gnd vdd DFFSR
XCLKBUF1_11 BUFX4_1/Y gnd DFFSR_87/CLK vdd CLKBUF1
XCLKBUF1_22 BUFX4_5/Y gnd DFFSR_50/CLK vdd CLKBUF1
XDFFSR_68 DFFSR_68/Q DFFSR_67/CLK DFFSR_69/R vdd DFFSR_68/D gnd vdd DFFSR
XFILL_1_0_2 gnd vdd FILL
XINVX1_118 BUFX2_12/A gnd INVX1_118/Y vdd INVX1
XINVX1_107 BUFX2_9/A gnd INVX1_107/Y vdd INVX1
XINVX1_129 BUFX2_15/A gnd INVX1_129/Y vdd INVX1
XFILL_9_1_2 gnd vdd FILL
XFILL_17_0_2 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XFILL_18_3_0 gnd vdd FILL
XFILL_18_4 gnd vdd FILL
XNOR2X1_46 NOR2X1_46/A NOR2X1_53/A gnd NOR2X1_46/Y vdd NOR2X1
XNAND3X1_35 AOI21X1_6/Y NAND3X1_35/B NOR2X1_52/B gnd AOI21X1_8/B vdd NAND3X1
XNAND3X1_13 MUX2X1_31/B DFFSR_33/Q INVX2_2/A gnd NAND3X1_13/Y vdd NAND3X1
XNOR2X1_13 INVX1_28/Y INVX1_29/Y gnd NOR2X1_13/Y vdd NOR2X1
XNAND3X1_57 gnd DFFSR_46/Q INVX4_4/Y gnd NAND3X1_57/Y vdd NAND3X1
XNAND3X1_68 INVX4_4/A gnd DFFSR_68/Q gnd NAND3X1_68/Y vdd NAND3X1
XNAND3X1_24 MUX2X1_80/B DFFSR_71/Q INVX2_4/A gnd NAND3X1_24/Y vdd NAND3X1
XNOR2X1_24 INVX1_161/A DFFSR_109/Q gnd BUFX4_18/A vdd NOR2X1
XNAND3X1_46 NAND3X1_45/Y NAND3X1_39/Y NOR2X1_47/Y gnd NAND3X1_46/Y vdd NAND3X1
XNOR2X1_35 DFFSR_142/Q NOR2X1_35/B gnd OR2X2_8/A vdd NOR2X1
XNOR2X1_57 INVX1_6/A NOR2X1_58/B gnd NOR2X1_57/Y vdd NOR2X1
XMUX2X1_86 MUX2X1_85/Y XOR2X1_8/Y OR2X2_8/Y gnd DFFSR_75/D vdd MUX2X1
XMUX2X1_53 MUX2X1_53/A MUX2X1_53/B NOR2X1_23/Y gnd MUX2X1_53/Y vdd MUX2X1
XMUX2X1_64 INVX1_67/A MUX2X1_56/A MUX2X1_66/S gnd MUX2X1_64/Y vdd MUX2X1
XMUX2X1_42 MUX2X1_42/A INVX1_40/A MUX2X1_43/S gnd MUX2X1_42/Y vdd MUX2X1
XMUX2X1_20 MUX2X1_6/A INVX1_24/A NOR2X1_7/Y gnd MUX2X1_20/Y vdd MUX2X1
XMUX2X1_31 MUX2X1_39/B MUX2X1_31/B NOR2X1_13/Y gnd MUX2X1_31/Y vdd MUX2X1
XMUX2X1_75 MUX2X1_55/A MUX2X1_75/B NOR2X1_28/Y gnd MUX2X1_75/Y vdd MUX2X1
XMUX2X1_97 MUX2X1_97/A INVX1_94/A NOR2X1_37/Y gnd MUX2X1_97/Y vdd MUX2X1
XFILL_23_2 gnd vdd FILL
XFILL_16_1 gnd vdd FILL
XDFFSR_1 DFFSR_1/Q DFFSR_1/CLK DFFSR_6/R vdd DFFSR_1/D gnd vdd DFFSR
XMUX2X1_109 INVX1_164/Y INVX2_10/Y MUX2X1_108/S gnd DFFSR_167/D vdd MUX2X1
XINVX1_49 DFFSR_57/Q gnd INVX1_49/Y vdd INVX1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XINVX1_38 DFFSR_33/Q gnd INVX1_38/Y vdd INVX1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XFILL_24_1_0 gnd vdd FILL
XNAND2X1_90 DFFSR_123/Q DFFSR_130/Q gnd NAND2X1_90/Y vdd NAND2X1
XFILL_7_2_0 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XOAI21X1_428 AOI21X1_8/C NOR2X1_44/Y NOR2X1_46/Y gnd XNOR2X1_13/A vdd OAI21X1
XOAI21X1_417 INVX1_138/Y OR2X2_12/Y OAI21X1_416/Y gnd DFFSR_129/D vdd OAI21X1
XOAI21X1_406 DFFSR_118/Q INVX1_130/Y OAI21X1_406/C gnd DFFSR_107/D vdd OAI21X1
XOAI21X1_439 OAI21X1_438/Y AOI22X1_16/Y OAI21X1_439/C gnd DFFSR_135/D vdd OAI21X1
XOAI21X1_11 NOR2X1_4/B INVX1_8/Y NAND2X1_4/Y gnd MUX2X1_4/A vdd OAI21X1
XOAI21X1_22 OR2X2_1/A OR2X2_1/B INVX1_1/A gnd INVX1_11/A vdd OAI21X1
XOAI21X1_55 BUFX4_14/Y MUX2X1_24/Y OAI21X1_55/C gnd OAI21X1_55/Y vdd OAI21X1
XOAI21X1_88 BUFX4_97/Y OR2X2_2/A DFFSR_5/Q gnd OAI21X1_88/Y vdd OAI21X1
XOAI21X1_99 BUFX4_37/Y MUX2X1_29/Y OAI21X1_99/C gnd OAI21X1_99/Y vdd OAI21X1
XOAI21X1_66 INVX1_16/Y OAI21X1_78/B NAND2X1_15/Y gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_77 INVX1_21/Y OAI21X1_69/B NAND3X1_6/Y gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_33 MUX2X1_7/S MUX2X1_13/Y OAI21X1_33/C gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_44 INVX1_2/A BUFX4_41/Y INVX1_22/A gnd OAI21X1_45/C vdd OAI21X1
XOAI21X1_203 BUFX4_96/Y MUX2X1_61/Y OAI21X1_202/Y gnd DFFPOSX1_61/D vdd OAI21X1
XOAI21X1_225 BUFX4_96/Y MUX2X1_72/Y OAI21X1_224/Y gnd OAI21X1_225/Y vdd OAI21X1
XOAI21X1_236 BUFX4_65/Y BUFX4_16/Y MUX2X1_78/B gnd OAI21X1_236/Y vdd OAI21X1
XOAI21X1_214 BUFX4_63/Y BUFX4_17/Y INVX1_61/A gnd OAI21X1_214/Y vdd OAI21X1
XOAI21X1_247 INVX1_65/Y NAND2X1_67/Y NAND3X1_18/Y gnd OAI21X1_249/A vdd OAI21X1
XOAI21X1_258 BUFX4_25/Y OR2X2_6/A DFFSR_50/Q gnd NAND2X1_80/A vdd OAI21X1
XOAI21X1_269 DFFSR_123/Q INVX1_75/Y NAND2X1_85/Y gnd MUX2X1_79/A vdd OAI21X1
XFILL_4_0_0 gnd vdd FILL
XDFFSR_58 DFFSR_58/Q DFFSR_74/CLK DFFSR_74/R vdd DFFSR_58/D gnd vdd DFFSR
XDFFSR_25 DFFSR_25/Q DFFSR_23/CLK BUFX4_78/Y vdd DFFSR_25/D gnd vdd DFFSR
XDFFSR_14 DFFSR_14/Q DFFSR_2/CLK DFFSR_2/S vdd DFFSR_14/D gnd vdd DFFSR
XDFFSR_36 OR2X2_3/B DFFSR_36/CLK DFFSR_34/R vdd XOR2X1_3/Y gnd vdd DFFSR
XDFFSR_47 DFFSR_47/Q CLKBUF1_3/Y BUFX4_28/Y vdd DFFSR_47/D gnd vdd DFFSR
XDFFSR_69 DFFSR_69/Q DFFSR_67/CLK DFFSR_69/R vdd DFFSR_69/D gnd vdd DFFSR
XCLKBUF1_23 BUFX4_2/Y gnd DFFSR_60/CLK vdd CLKBUF1
XCLKBUF1_12 BUFX4_6/Y gnd CLKBUF1_12/Y vdd CLKBUF1
XCLKBUF1_34 BUFX4_6/Y gnd CLKBUF1_34/Y vdd CLKBUF1
XINVX1_108 BUFX2_5/Y gnd DFFSR_82/D vdd INVX1
XINVX1_119 BUFX2_13/A gnd INVX1_119/Y vdd INVX1
XFILL_4_1 gnd vdd FILL
XFILL_2_3_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XFILL_18_3_1 gnd vdd FILL
XNAND3X1_14 MUX2X1_32/B DFFSR_33/Q INVX2_2/A gnd NAND3X1_14/Y vdd NAND3X1
XNOR2X1_36 OR2X2_8/B OR2X2_8/A gnd NOR2X1_36/Y vdd NOR2X1
XNAND3X1_36 INVX2_6/A BUFX4_58/Y INVX4_1/Y gnd NAND3X1_38/B vdd NAND3X1
XNOR2X1_47 OAI22X1_4/Y NOR2X1_47/B gnd NOR2X1_47/Y vdd NOR2X1
XNAND3X1_47 DFFSR_135/Q NOR2X1_44/A NAND3X1_39/Y gnd NAND3X1_49/A vdd NAND3X1
XNOR2X1_14 INVX1_159/A DFFSR_95/Q gnd BUFX4_57/A vdd NOR2X1
XNAND3X1_58 BUFX4_9/Y DFFSR_27/Q INVX4_5/Y gnd NAND3X1_58/Y vdd NAND3X1
XNOR2X1_58 INVX1_7/A NOR2X1_58/B gnd NOR2X1_58/Y vdd NOR2X1
XNOR2X1_25 NOR2X1_25/A NOR2X1_25/B gnd OR2X2_6/A vdd NOR2X1
XNAND3X1_69 gnd DFFSR_50/Q INVX4_4/Y gnd NAND3X1_69/Y vdd NAND3X1
XNAND3X1_25 MUX2X1_81/B DFFSR_71/Q INVX2_4/A gnd NAND3X1_25/Y vdd NAND3X1
XMUX2X1_65 INVX1_69/A MUX2X1_71/A MUX2X1_66/S gnd MUX2X1_65/Y vdd MUX2X1
XMUX2X1_10 INVX1_15/A MUX2X1_2/A MUX2X1_9/S gnd MUX2X1_10/Y vdd MUX2X1
XMUX2X1_21 MUX2X1_1/A MUX2X1_21/B NOR2X1_8/Y gnd MUX2X1_21/Y vdd MUX2X1
XMUX2X1_43 MUX2X1_49/A INVX1_42/A MUX2X1_43/S gnd MUX2X1_43/Y vdd MUX2X1
XMUX2X1_32 MUX2X1_46/A MUX2X1_32/B NOR2X1_13/Y gnd MUX2X1_32/Y vdd MUX2X1
XMUX2X1_98 MUX2X1_92/B INVX1_96/A NOR2X1_37/Y gnd MUX2X1_98/Y vdd MUX2X1
XMUX2X1_76 MUX2X1_56/A MUX2X1_76/B NOR2X1_28/Y gnd MUX2X1_76/Y vdd MUX2X1
XMUX2X1_54 MUX2X1_68/A MUX2X1_54/B NOR2X1_23/Y gnd MUX2X1_54/Y vdd MUX2X1
XMUX2X1_87 INVX1_84/A MUX2X1_79/A MUX2X1_87/S gnd MUX2X1_87/Y vdd MUX2X1
XFILL_23_3 gnd vdd FILL
XDFFSR_2 DFFSR_2/Q DFFSR_2/CLK vdd DFFSR_2/S DFFSR_2/D gnd vdd DFFSR
XNAND2X1_91 OR2X2_7/A OR2X2_7/B gnd NAND2X1_92/B vdd NAND2X1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XNAND2X1_80 NAND2X1_80/A NAND2X1_80/B gnd DFFSR_50/D vdd NAND2X1
XFILL_24_1_1 gnd vdd FILL
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XOAI21X1_429 OAI22X1_2/Y NOR2X1_43/B NAND2X1_145/Y gnd NAND3X1_35/B vdd OAI21X1
XOAI21X1_418 OR2X2_12/A BUFX2_25/A DFFSR_130/Q gnd OAI21X1_419/C vdd OAI21X1
XOAI21X1_407 DFFSR_118/Q INVX1_131/Y OAI21X1_407/C gnd DFFSR_108/D vdd OAI21X1
XOAI21X1_12 BUFX4_74/Y BUFX4_42/Y MUX2X1_4/B gnd OAI21X1_13/C vdd OAI21X1
XOAI21X1_23 INVX1_11/Y DFFSR_2/D NOR2X1_6/Y gnd NAND2X1_9/A vdd OAI21X1
XOAI21X1_34 OR2X2_9/A BUFX4_44/Y INVX1_23/A gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_45 MUX2X1_7/S MUX2X1_19/Y OAI21X1_45/C gnd OAI21X1_45/Y vdd OAI21X1
XOAI21X1_89 BUFX4_97/Y OR2X2_2/A DFFSR_6/Q gnd NAND2X1_28/A vdd OAI21X1
XOAI21X1_67 OAI21X1_65/Y OAI21X1_66/Y NOR2X1_6/Y gnd NAND2X1_16/B vdd OAI21X1
XOAI21X1_78 INVX1_22/Y OAI21X1_78/B NAND2X1_21/Y gnd OAI21X1_78/Y vdd OAI21X1
XOAI21X1_56 INVX1_2/A BUFX4_41/Y MUX2X1_25/B gnd OAI21X1_56/Y vdd OAI21X1
XOAI21X1_237 BUFX4_96/Y MUX2X1_78/Y OAI21X1_236/Y gnd OAI21X1_237/Y vdd OAI21X1
XOAI21X1_215 BUFX4_94/Y MUX2X1_67/Y OAI21X1_214/Y gnd DFFPOSX1_55/D vdd OAI21X1
XOAI21X1_226 BUFX4_63/Y BUFX4_17/Y MUX2X1_73/B gnd OAI21X1_226/Y vdd OAI21X1
XOAI21X1_204 BUFX4_63/Y BUFX4_17/Y INVX1_63/A gnd OAI21X1_204/Y vdd OAI21X1
XOAI21X1_248 INVX1_66/Y NAND2X1_69/Y NAND2X1_73/Y gnd OAI21X1_249/B vdd OAI21X1
XOAI21X1_259 INVX1_71/Y NAND2X1_67/Y NAND3X1_21/Y gnd OAI21X1_261/A vdd OAI21X1
XFILL_4_0_1 gnd vdd FILL
XDFFSR_59 BUFX2_4/A CLKBUF1_32/Y vdd DFFSR_71/R DFFSR_59/D gnd vdd DFFSR
XDFFSR_15 INVX1_5/A DFFSR_1/CLK DFFSR_5/R vdd DFFSR_15/D gnd vdd DFFSR
XDFFSR_26 DFFSR_26/Q CLKBUF1_34/Y DFFSR_29/R vdd DFFSR_26/D gnd vdd DFFSR
XDFFSR_37 OR2X2_3/A DFFSR_36/CLK DFFSR_34/R vdd DFFSR_37/D gnd vdd DFFSR
XDFFSR_48 DFFSR_48/Q DFFSR_45/CLK BUFX4_28/Y vdd DFFSR_48/D gnd vdd DFFSR
XCLKBUF1_13 BUFX4_3/Y gnd CLKBUF1_13/Y vdd CLKBUF1
XCLKBUF1_35 BUFX4_6/Y gnd CLKBUF1_35/Y vdd CLKBUF1
XCLKBUF1_24 BUFX4_1/Y gnd CLKBUF1_24/Y vdd CLKBUF1
XINVX1_109 OR2X2_10/Y gnd DFFSR_95/D vdd INVX1
XFILL_2_3_2 gnd vdd FILL
XFILL_10_2_2 gnd vdd FILL
XFILL_18_3_2 gnd vdd FILL
XNAND3X1_15 OR2X2_5/A OR2X2_5/B INVX1_49/Y gnd AOI21X1_3/B vdd NAND3X1
XNAND3X1_37 INVX2_5/A INVX2_6/Y INVX4_1/Y gnd NAND3X1_37/Y vdd NAND3X1
XNAND3X1_26 MUX2X1_82/B DFFSR_71/Q INVX2_4/A gnd NAND3X1_26/Y vdd NAND3X1
XNAND3X1_48 NAND3X1_48/A NAND3X1_48/B AOI22X1_12/Y gnd NAND3X1_48/Y vdd NAND3X1
XNOR2X1_48 INVX4_1/A INVX2_6/Y gnd NOR2X1_48/Y vdd NOR2X1
XNOR2X1_15 NOR2X1_15/A DFFSR_96/Q gnd OR2X2_4/A vdd NOR2X1
XNOR2X1_59 INVX1_8/A NOR2X1_58/B gnd NOR2X1_59/Y vdd NOR2X1
XNAND3X1_59 BUFX2_1/Y gnd DFFSR_65/Q gnd NAND3X1_59/Y vdd NAND3X1
XNOR2X1_26 OR2X2_6/B OR2X2_6/A gnd NOR2X1_26/Y vdd NOR2X1
XNOR2X1_37 DFFSR_73/Q INVX1_77/Y gnd NOR2X1_37/Y vdd NOR2X1
XMUX2X1_11 INVX1_17/A MUX2X1_3/A MUX2X1_9/S gnd MUX2X1_11/Y vdd MUX2X1
XMUX2X1_66 INVX1_71/A MUX2X1_66/B MUX2X1_66/S gnd MUX2X1_66/Y vdd MUX2X1
XMUX2X1_77 MUX2X1_71/A MUX2X1_77/B NOR2X1_28/Y gnd MUX2X1_77/Y vdd MUX2X1
XMUX2X1_55 MUX2X1_55/A MUX2X1_55/B NOR2X1_23/Y gnd MUX2X1_55/Y vdd MUX2X1
XMUX2X1_44 MUX2X1_44/A INVX1_44/A MUX2X1_43/S gnd MUX2X1_44/Y vdd MUX2X1
XMUX2X1_22 MUX2X1_2/A MUX2X1_22/B NOR2X1_8/Y gnd MUX2X1_22/Y vdd MUX2X1
XMUX2X1_33 OR2X2_3/A XOR2X1_4/Y AND2X2_2/A gnd MUX2X1_33/Y vdd MUX2X1
XMUX2X1_88 INVX1_87/A MUX2X1_94/A MUX2X1_87/S gnd MUX2X1_88/Y vdd MUX2X1
XMUX2X1_99 MUX2X1_79/A MUX2X1_99/B NOR2X1_38/Y gnd MUX2X1_99/Y vdd MUX2X1
XDFFSR_3 DFFSR_3/Q DFFSR_8/CLK DFFSR_8/R vdd DFFSR_3/D gnd vdd DFFSR
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XINVX1_29 DFFSR_34/Q gnd INVX1_29/Y vdd INVX1
XNAND2X1_92 DFFSR_76/Q NAND2X1_92/B gnd AOI21X1_4/A vdd NAND2X1
XNAND2X1_70 NAND2X1_70/A NAND2X1_70/B gnd DFFSR_45/D vdd NAND2X1
XNAND2X1_81 NAND2X1_81/A NAND2X1_70/B gnd DFFSR_41/D vdd NAND2X1
XFILL_24_1_2 gnd vdd FILL
XFILL_7_2_2 gnd vdd FILL
XFILL_15_1_2 gnd vdd FILL
XFILL_21_1 gnd vdd FILL
XOAI21X1_419 INVX1_139/Y OR2X2_12/Y OAI21X1_419/C gnd DFFSR_130/D vdd OAI21X1
XOAI21X1_408 BUFX4_21/Y BUFX2_25/A DFFSR_125/Q gnd OAI21X1_408/Y vdd OAI21X1
XOAI21X1_13 BUFX4_14/Y MUX2X1_4/Y OAI21X1_13/C gnd OAI21X1_13/Y vdd OAI21X1
XOAI21X1_68 BUFX4_97/Y OR2X2_2/A DFFSR_9/Q gnd NAND2X1_18/A vdd OAI21X1
XOAI21X1_24 BUFX4_76/Y BUFX4_43/Y INVX1_12/A gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_46 BUFX4_73/Y BUFX4_44/Y INVX1_24/A gnd OAI21X1_46/Y vdd OAI21X1
XOAI21X1_35 BUFX4_10/Y MUX2X1_14/Y OAI21X1_34/Y gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_57 MUX2X1_7/S MUX2X1_25/Y OAI21X1_56/Y gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_79 OAI21X1_77/Y OAI21X1_78/Y NOR2X1_6/Y gnd OAI21X1_79/Y vdd OAI21X1
XOAI21X1_216 BUFX4_65/Y BUFX4_16/Y INVX1_64/A gnd OAI21X1_217/C vdd OAI21X1
XOAI21X1_238 BUFX4_26/Y OR2X2_6/A DFFSR_45/Q gnd NAND2X1_70/A vdd OAI21X1
XOAI21X1_249 OAI21X1_249/A OAI21X1_249/B NOR2X1_26/Y gnd NAND2X1_83/B vdd OAI21X1
XOAI21X1_227 BUFX4_94/Y MUX2X1_73/Y OAI21X1_226/Y gnd DFFPOSX1_49/D vdd OAI21X1
XOAI21X1_205 BUFX4_96/Y MUX2X1_62/Y OAI21X1_204/Y gnd DFFPOSX1_62/D vdd OAI21X1
XFILL_4_0_2 gnd vdd FILL
XDFFSR_27 DFFSR_27/Q CLKBUF1_16/Y BUFX4_78/Y vdd DFFSR_27/D gnd vdd DFFSR
XDFFSR_16 INVX1_4/A DFFSR_1/CLK DFFSR_5/R vdd DFFSR_16/D gnd vdd DFFSR
XDFFSR_38 INVX1_25/A DFFSR_33/CLK DFFSR_38/R vdd DFFSR_38/D gnd vdd DFFSR
XDFFSR_49 DFFSR_49/Q DFFSR_50/CLK DFFSR_41/R vdd DFFSR_49/D gnd vdd DFFSR
XCLKBUF1_36 BUFX4_3/Y gnd CLKBUF1_36/Y vdd CLKBUF1
XCLKBUF1_25 BUFX4_2/Y gnd CLKBUF1_25/Y vdd CLKBUF1
XCLKBUF1_14 BUFX4_2/Y gnd CLKBUF1_14/Y vdd CLKBUF1
XFILL_22_2_0 gnd vdd FILL
XBUFX4_90 BUFX2_4/A gnd OR2X2_8/B vdd BUFX4
XFILL_5_3_0 gnd vdd FILL
XFILL_13_2_0 gnd vdd FILL
XNAND3X1_38 INVX2_7/Y NAND3X1_38/B NAND3X1_37/Y gnd NOR2X1_47/B vdd NAND3X1
XNAND3X1_16 MUX2X1_53/B DFFSR_52/Q INVX2_3/A gnd NAND3X1_16/Y vdd NAND3X1
XNAND3X1_49 NAND3X1_49/A NAND3X1_46/Y NAND3X1_49/C gnd AOI22X1_16/D vdd NAND3X1
XNAND3X1_27 MUX2X1_83/B DFFSR_71/Q INVX2_4/A gnd NAND3X1_27/Y vdd NAND3X1
XNOR2X1_27 DFFSR_54/Q INVX1_53/Y gnd NOR2X1_27/Y vdd NOR2X1
XNOR2X1_49 INVX2_6/A INVX4_1/Y gnd NOR2X1_49/Y vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_16 OR2X2_4/B OR2X2_4/A gnd NOR2X1_16/Y vdd NOR2X1
XNOR2X1_38 DFFSR_73/Q DFFSR_72/Q gnd NOR2X1_38/Y vdd NOR2X1
XFILL_10_0_0 gnd vdd FILL
XMUX2X1_12 INVX1_19/A MUX2X1_4/A MUX2X1_9/S gnd MUX2X1_12/Y vdd MUX2X1
XMUX2X1_23 MUX2X1_3/A MUX2X1_23/B NOR2X1_8/Y gnd MUX2X1_23/Y vdd MUX2X1
XMUX2X1_45 MUX2X1_39/B INVX1_46/A MUX2X1_43/S gnd MUX2X1_45/Y vdd MUX2X1
XMUX2X1_34 MUX2X1_33/Y XOR2X1_4/Y OR2X2_4/Y gnd DFFSR_37/D vdd MUX2X1
XFILL_18_1_0 gnd vdd FILL
XMUX2X1_56 MUX2X1_56/A MUX2X1_56/B NOR2X1_23/Y gnd MUX2X1_56/Y vdd MUX2X1
XMUX2X1_78 MUX2X1_66/B MUX2X1_78/B NOR2X1_28/Y gnd MUX2X1_78/Y vdd MUX2X1
XMUX2X1_89 INVX1_89/A MUX2X1_89/B MUX2X1_87/S gnd MUX2X1_89/Y vdd MUX2X1
XMUX2X1_67 MUX2X1_53/A INVX1_61/A NOR2X1_27/Y gnd MUX2X1_67/Y vdd MUX2X1
XDFFSR_4 DFFSR_4/Q DFFSR_8/CLK DFFSR_8/R vdd DFFSR_4/D gnd vdd DFFSR
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XNAND2X1_93 NAND2X1_93/A NAND2X1_93/B gnd DFFSR_76/D vdd NAND2X1
XNAND2X1_60 DFFSR_109/Q DFFSR_114/Q gnd NAND2X1_60/Y vdd NAND2X1
XNAND2X1_82 NAND2X1_82/A NAND2X1_72/B gnd DFFSR_42/D vdd NAND2X1
XNAND2X1_71 MUX2X1_74/B NOR2X1_29/Y gnd NAND2X1_71/Y vdd NAND2X1
XFILL_21_2 gnd vdd FILL
XOAI21X1_409 INVX1_134/Y OR2X2_12/Y OAI21X1_408/Y gnd DFFSR_125/D vdd OAI21X1
XFILL_14_1 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_69 INVX1_17/Y OAI21X1_69/B NAND3X1_4/Y gnd OAI21X1_69/Y vdd OAI21X1
XOAI21X1_36 BUFX4_76/Y BUFX4_43/Y INVX1_13/A gnd OAI21X1_36/Y vdd OAI21X1
XOAI21X1_25 BUFX4_11/Y MUX2X1_9/Y OAI21X1_24/Y gnd OAI21X1_25/Y vdd OAI21X1
XOAI21X1_58 BUFX4_73/Y BUFX4_43/Y MUX2X1_26/B gnd OAI21X1_59/C vdd OAI21X1
XOAI21X1_47 BUFX4_10/Y MUX2X1_20/Y OAI21X1_46/Y gnd OAI21X1_47/Y vdd OAI21X1
XOAI21X1_14 NOR2X1_4/B INVX1_9/Y NAND2X1_5/Y gnd MUX2X1_5/A vdd OAI21X1
XOAI21X1_217 BUFX4_96/Y MUX2X1_68/Y OAI21X1_217/C gnd DFFPOSX1_56/D vdd OAI21X1
XOAI21X1_228 BUFX4_63/Y BUFX4_17/Y MUX2X1_74/B gnd OAI21X1_228/Y vdd OAI21X1
XOAI21X1_239 INVX1_60/Y NAND2X1_67/Y NAND3X1_16/Y gnd OAI21X1_241/A vdd OAI21X1
XOAI21X1_206 BUFX4_64/Y BUFX4_18/Y INVX1_65/A gnd OAI21X1_206/Y vdd OAI21X1
XDFFSR_17 OR2X2_1/B DFFSR_9/CLK DFFSR_6/R vdd DFFSR_17/D gnd vdd DFFSR
XDFFSR_28 DFFSR_28/Q CLKBUF1_34/Y DFFSR_29/R vdd DFFSR_28/D gnd vdd DFFSR
XDFFSR_39 BUFX4_63/A DFFSR_54/CLK DFFSR_41/R vdd DFFSR_39/D gnd vdd DFFSR
XCLKBUF1_15 BUFX4_3/Y gnd DFFSR_36/CLK vdd CLKBUF1
XCLKBUF1_26 BUFX4_5/Y gnd CLKBUF1_26/Y vdd CLKBUF1
XCLKBUF1_37 BUFX4_2/Y gnd DFFSR_74/CLK vdd CLKBUF1
XBUFX4_91 BUFX2_4/A gnd BUFX4_91/Y vdd BUFX4
XBUFX4_80 INVX8_2/Y gnd DFFSR_34/R vdd BUFX4
XFILL_22_2_1 gnd vdd FILL
XXNOR2X1_1 BUFX4_11/Y INVX1_5/A gnd DFFSR_15/D vdd XNOR2X1
XFILL_5_3_1 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XFILL_13_2_1 gnd vdd FILL
XAND2X2_1 AND2X2_1/A INVX1_1/A gnd AND2X2_1/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XNOR2X1_28 DFFSR_54/Q DFFSR_53/Q gnd NOR2X1_28/Y vdd NOR2X1
XNAND3X1_39 NAND3X1_33/B AOI21X1_9/Y AOI22X1_1/Y gnd NAND3X1_39/Y vdd NAND3X1
XNOR2X1_17 INVX1_28/A INVX1_29/Y gnd MUX2X1_43/S vdd NOR2X1
XNAND3X1_17 MUX2X1_54/B DFFSR_52/Q INVX2_3/A gnd NAND3X1_17/Y vdd NAND3X1
XNAND3X1_28 MUX2X1_84/B DFFSR_71/Q INVX2_4/A gnd NAND3X1_28/Y vdd NAND3X1
XFILL_2_1_1 gnd vdd FILL
XNOR2X1_39 DFFSR_71/Q INVX2_4/A gnd NOR2X1_39/Y vdd NOR2X1
XFILL_10_0_1 gnd vdd FILL
XMUX2X1_57 MUX2X1_71/A MUX2X1_57/B NOR2X1_23/Y gnd MUX2X1_57/Y vdd MUX2X1
XMUX2X1_24 MUX2X1_4/A MUX2X1_24/B NOR2X1_8/Y gnd MUX2X1_24/Y vdd MUX2X1
XMUX2X1_35 INVX1_36/A MUX2X1_41/A MUX2X1_39/S gnd MUX2X1_35/Y vdd MUX2X1
XMUX2X1_13 INVX1_21/A MUX2X1_5/A MUX2X1_9/S gnd MUX2X1_13/Y vdd MUX2X1
XMUX2X1_46 MUX2X1_46/A INVX1_48/A MUX2X1_43/S gnd MUX2X1_46/Y vdd MUX2X1
XFILL_18_1_1 gnd vdd FILL
XMUX2X1_79 MUX2X1_79/A MUX2X1_79/B MUX2X1_79/S gnd MUX2X1_79/Y vdd MUX2X1
XMUX2X1_68 MUX2X1_68/A INVX1_64/A NOR2X1_27/Y gnd MUX2X1_68/Y vdd MUX2X1
XDFFSR_5 DFFSR_5/Q DFFSR_9/CLK DFFSR_5/R vdd DFFSR_5/D gnd vdd DFFSR
XNAND2X1_50 NAND2X1_50/A NAND2X1_50/B gnd DFFSR_30/D vdd NAND2X1
XNAND2X1_61 DFFSR_109/Q INVX1_126/A gnd NAND2X1_61/Y vdd NAND2X1
XNAND2X1_83 NAND2X1_83/A NAND2X1_83/B gnd DFFSR_43/D vdd NAND2X1
XNAND2X1_72 NAND2X1_72/A NAND2X1_72/B gnd DFFSR_46/D vdd NAND2X1
XNAND2X1_94 DFFSR_73/Q INVX1_77/Y gnd MUX2X1_87/S vdd NAND2X1
XFILL_21_3 gnd vdd FILL
XFILL_14_2 gnd vdd FILL
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_37 BUFX4_11/Y MUX2X1_15/Y OAI21X1_36/Y gnd DFFPOSX1_7/D vdd OAI21X1
XOAI21X1_48 BUFX4_74/Y BUFX4_42/Y MUX2X1_21/B gnd OAI21X1_48/Y vdd OAI21X1
XOAI21X1_59 AND2X2_1/A MUX2X1_26/Y OAI21X1_59/C gnd DFFPOSX1_6/D vdd OAI21X1
XOAI21X1_26 BUFX4_73/Y BUFX4_44/Y INVX1_15/A gnd OAI21X1_27/C vdd OAI21X1
XOAI21X1_15 INVX1_2/A BUFX4_41/Y MUX2X1_5/B gnd OAI21X1_16/C vdd OAI21X1
XOAI21X1_229 BUFX4_94/Y MUX2X1_74/Y OAI21X1_228/Y gnd DFFPOSX1_50/D vdd OAI21X1
XOAI21X1_218 BUFX4_64/Y BUFX4_18/Y INVX1_66/A gnd OAI21X1_219/C vdd OAI21X1
XOAI21X1_207 AND2X2_3/A MUX2X1_63/Y OAI21X1_206/Y gnd OAI21X1_207/Y vdd OAI21X1
XDFFSR_29 DFFSR_29/Q CLKBUF1_16/Y DFFSR_29/R vdd DFFSR_29/D gnd vdd DFFSR
XDFFSR_18 OR2X2_1/A DFFSR_2/CLK DFFSR_2/S vdd MUX2X1_8/Y gnd vdd DFFSR
XCLKBUF1_16 BUFX4_3/Y gnd CLKBUF1_16/Y vdd CLKBUF1
XCLKBUF1_27 BUFX4_3/Y gnd CLKBUF1_27/Y vdd CLKBUF1
XCLKBUF1_38 BUFX4_1/Y gnd CLKBUF1_38/Y vdd CLKBUF1
XBUFX4_92 BUFX4_93/A gnd BUFX4_92/Y vdd BUFX4
XBUFX4_70 INVX8_9/Y gnd BUFX4_70/Y vdd BUFX4
XBUFX4_81 BUFX4_82/A gnd BUFX4_81/Y vdd BUFX4
XFILL_22_2_2 gnd vdd FILL
XXNOR2X1_2 NOR2X1_10/Y INVX1_4/Y gnd DFFSR_16/D vdd XNOR2X1
XFILL_5_3_2 gnd vdd FILL
XFILL_13_2_2 gnd vdd FILL
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XOAI21X1_390 DFFSR_104/Q INVX1_119/Y OAI21X1_390/C gnd DFFSR_94/D vdd OAI21X1
XAND2X2_2 AND2X2_2/A INVX1_25/A gnd AND2X2_2/Y vdd AND2X2
XFILL_2_2 gnd vdd FILL
XNAND3X1_29 INVX2_6/A BUFX2_4/Y INVX4_1/Y gnd NAND3X1_30/B vdd NAND3X1
XNAND3X1_18 MUX2X1_55/B DFFSR_52/Q INVX2_3/A gnd NAND3X1_18/Y vdd NAND3X1
XNOR2X1_18 INVX1_28/A DFFSR_34/Q gnd NOR2X1_18/Y vdd NOR2X1
XNOR2X1_29 DFFSR_52/Q INVX2_3/A gnd NOR2X1_29/Y vdd NOR2X1
XFILL_2_1_2 gnd vdd FILL
XFILL_10_0_2 gnd vdd FILL
XMUX2X1_58 MUX2X1_66/B MUX2X1_58/B NOR2X1_23/Y gnd MUX2X1_58/Y vdd MUX2X1
XMUX2X1_36 INVX1_39/A MUX2X1_42/A MUX2X1_39/S gnd MUX2X1_36/Y vdd MUX2X1
XMUX2X1_47 MUX2X1_41/A MUX2X1_47/B NOR2X1_18/Y gnd MUX2X1_47/Y vdd MUX2X1
XMUX2X1_14 INVX1_23/A MUX2X1_6/A MUX2X1_9/S gnd MUX2X1_14/Y vdd MUX2X1
XMUX2X1_25 MUX2X1_5/A MUX2X1_25/B NOR2X1_8/Y gnd MUX2X1_25/Y vdd MUX2X1
XFILL_18_1_2 gnd vdd FILL
XMUX2X1_69 MUX2X1_55/A INVX1_66/A NOR2X1_27/Y gnd MUX2X1_69/Y vdd MUX2X1
XDFFSR_6 DFFSR_6/Q DFFSR_9/CLK DFFSR_6/R vdd DFFSR_6/D gnd vdd DFFSR
XNAND2X1_95 DFFSR_71/Q INVX2_4/Y gnd NAND2X1_95/Y vdd NAND2X1
XNAND2X1_40 MUX2X1_47/B NOR2X1_19/Y gnd NAND2X1_40/Y vdd NAND2X1
XNAND2X1_51 MUX2X1_52/B NOR2X1_19/Y gnd NAND2X1_51/Y vdd NAND2X1
XNAND2X1_62 DFFSR_109/Q INVX1_127/A gnd NAND2X1_62/Y vdd NAND2X1
XNAND2X1_84 NAND2X1_84/A NAND2X1_76/B gnd DFFSR_44/D vdd NAND2X1
XNAND2X1_73 MUX2X1_75/B NOR2X1_29/Y gnd NAND2X1_73/Y vdd NAND2X1
XFILL_20_3_0 gnd vdd FILL
XFILL_11_3_0 gnd vdd FILL
XFILL_7_0_2 gnd vdd FILL
XOAI21X1_16 MUX2X1_7/S MUX2X1_5/Y OAI21X1_16/C gnd OAI21X1_16/Y vdd OAI21X1
XOAI21X1_49 BUFX4_14/Y MUX2X1_21/Y OAI21X1_48/Y gnd DFFPOSX1_1/D vdd OAI21X1
XOAI21X1_27 BUFX4_10/Y MUX2X1_10/Y OAI21X1_27/C gnd OAI21X1_27/Y vdd OAI21X1
XOAI21X1_38 INVX1_2/A BUFX4_41/Y INVX1_16/A gnd OAI21X1_39/C vdd OAI21X1
XOAI21X1_208 BUFX4_62/Y BUFX4_16/Y INVX1_67/A gnd OAI21X1_208/Y vdd OAI21X1
XOAI21X1_219 AND2X2_3/A MUX2X1_69/Y OAI21X1_219/C gnd DFFPOSX1_57/D vdd OAI21X1
XFILL_0_2_0 gnd vdd FILL
XFILL_8_3_0 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XDFFSR_19 INVX1_1/A DFFSR_2/CLK DFFSR_6/R vdd DFFSR_19/D gnd vdd DFFSR
XCLKBUF1_39 BUFX4_5/Y gnd DFFSR_54/CLK vdd CLKBUF1
XCLKBUF1_17 BUFX4_4/Y gnd DFFSR_23/CLK vdd CLKBUF1
XCLKBUF1_28 BUFX4_6/Y gnd DFFSR_33/CLK vdd CLKBUF1
XBUFX4_93 BUFX4_93/A gnd BUFX4_93/Y vdd BUFX4
XBUFX4_60 BUFX2_3/A gnd OR2X2_4/B vdd BUFX4
XBUFX4_71 INVX8_9/Y gnd BUFX4_71/Y vdd BUFX4
XBUFX4_82 BUFX4_82/A gnd BUFX4_82/Y vdd BUFX4
XXNOR2X1_3 NOR2X1_6/Y INVX2_1/Y gnd DFFSR_13/D vdd XNOR2X1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_22_0_0 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XOAI21X1_391 BUFX4_62/Y BUFX2_24/A DFFSR_111/Q gnd OAI21X1_392/C vdd OAI21X1
XAND2X2_3 AND2X2_3/A DFFSR_57/Q gnd AND2X2_3/Y vdd AND2X2
XOAI21X1_380 BUFX4_31/Y OR2X2_10/B DFFSR_100/Q gnd OAI21X1_380/Y vdd OAI21X1
XNAND3X1_19 MUX2X1_56/B DFFSR_52/Q INVX2_3/A gnd NAND3X1_19/Y vdd NAND3X1
XNOR2X1_19 DFFSR_33/Q INVX2_2/A gnd NOR2X1_19/Y vdd NOR2X1
XMUX2X1_37 INVX1_41/A MUX2X1_49/A MUX2X1_39/S gnd MUX2X1_37/Y vdd MUX2X1
XMUX2X1_48 MUX2X1_42/A MUX2X1_48/B NOR2X1_18/Y gnd MUX2X1_48/Y vdd MUX2X1
XMUX2X1_15 MUX2X1_1/A INVX1_13/A NOR2X1_7/Y gnd MUX2X1_15/Y vdd MUX2X1
XMUX2X1_26 MUX2X1_6/A MUX2X1_26/B NOR2X1_8/Y gnd MUX2X1_26/Y vdd MUX2X1
XMUX2X1_59 OR2X2_5/A XOR2X1_6/Y AND2X2_3/A gnd MUX2X1_59/Y vdd MUX2X1
XDFFSR_7 DFFSR_7/Q DFFSR_8/CLK DFFSR_8/R vdd DFFSR_7/D gnd vdd DFFSR
XNAND2X1_63 OR2X2_5/A OR2X2_5/B gnd NAND2X1_64/B vdd NAND2X1
XNAND2X1_30 DFFSR_95/Q DFFSR_98/Q gnd NAND2X1_30/Y vdd NAND2X1
XNAND2X1_41 INVX2_2/A INVX1_38/Y gnd NAND2X1_41/Y vdd NAND2X1
XNAND2X1_52 NAND2X1_52/A NAND2X1_52/B gnd DFFSR_31/D vdd NAND2X1
XNAND2X1_74 NAND2X1_74/A NAND2X1_83/B gnd DFFSR_47/D vdd NAND2X1
XNAND2X1_85 DFFSR_123/Q DFFSR_125/Q gnd NAND2X1_85/Y vdd NAND2X1
XNAND2X1_96 MUX2X1_99/B NOR2X1_39/Y gnd NAND2X1_96/Y vdd NAND2X1
XFILL_20_3_1 gnd vdd FILL
XFILL_11_3_1 gnd vdd FILL
XOAI22X1_1 INVX1_146/Y OAI22X1_4/B INVX2_5/Y OAI22X1_4/D gnd OAI22X1_1/Y vdd OAI22X1
XINVX2_10 INVX2_10/A gnd INVX2_10/Y vdd INVX2
XOAI21X1_28 BUFX4_76/Y BUFX4_43/Y INVX1_17/A gnd OAI21X1_29/C vdd OAI21X1
XOAI21X1_39 AND2X2_1/A MUX2X1_16/Y OAI21X1_39/C gnd OAI21X1_39/Y vdd OAI21X1
XOAI21X1_17 NOR2X1_4/B INVX1_10/Y NAND2X1_6/Y gnd MUX2X1_6/A vdd OAI21X1
XOAI21X1_209 BUFX4_92/Y MUX2X1_64/Y OAI21X1_208/Y gnd OAI21X1_209/Y vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XFILL_0_2_1 gnd vdd FILL
XFILL_8_3_1 gnd vdd FILL
XFILL_16_2_1 gnd vdd FILL
XBUFX4_50 INVX8_1/Y gnd DFFSR_6/R vdd BUFX4
XCLKBUF1_29 BUFX4_6/Y gnd DFFSR_21/CLK vdd CLKBUF1
XCLKBUF1_18 BUFX4_5/Y gnd DFFSR_67/CLK vdd CLKBUF1
XBUFX4_61 BUFX4_63/A gnd BUFX4_61/Y vdd BUFX4
XBUFX4_72 DFFSR_1/Q gnd OR2X2_9/A vdd BUFX4
XBUFX4_83 BUFX4_82/A gnd BUFX4_83/Y vdd BUFX4
XBUFX4_94 BUFX4_93/A gnd BUFX4_94/Y vdd BUFX4
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XXNOR2X1_4 BUFX4_38/Y DFFSR_34/Q gnd DFFSR_34/D vdd XNOR2X1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_22_0_1 gnd vdd FILL
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XOAI21X1_392 INVX1_122/Y OR2X2_11/Y OAI21X1_392/C gnd DFFSR_111/D vdd OAI21X1
XAND2X2_4 AND2X2_4/A DFFSR_76/Q gnd AND2X2_4/Y vdd AND2X2
XOAI21X1_381 INVX1_113/Y OR2X2_10/Y OAI21X1_380/Y gnd DFFSR_100/D vdd OAI21X1
XOAI21X1_370 DFFSR_90/Q INVX1_104/Y OAI21X1_370/C gnd DFFSR_77/D vdd OAI21X1
XMUX2X1_27 MUX2X1_41/A NAND3X1_9/A NOR2X1_13/Y gnd MUX2X1_27/Y vdd MUX2X1
XMUX2X1_16 MUX2X1_2/A INVX1_16/A NOR2X1_7/Y gnd MUX2X1_16/Y vdd MUX2X1
XMUX2X1_38 INVX1_43/A MUX2X1_44/A MUX2X1_39/S gnd MUX2X1_38/Y vdd MUX2X1
XMUX2X1_49 MUX2X1_49/A MUX2X1_49/B NOR2X1_18/Y gnd MUX2X1_49/Y vdd MUX2X1
XDFFSR_8 DFFSR_8/Q DFFSR_8/CLK DFFSR_8/R vdd DFFSR_8/D gnd vdd DFFSR
XNAND2X1_64 DFFSR_57/Q NAND2X1_64/B gnd AOI21X1_3/A vdd NAND2X1
XNAND2X1_86 DFFSR_123/Q DFFSR_126/Q gnd NAND2X1_86/Y vdd NAND2X1
XNAND2X1_31 DFFSR_95/Q DFFSR_99/Q gnd NAND2X1_31/Y vdd NAND2X1
XNAND2X1_42 NAND2X1_42/A NAND2X1_42/B gnd DFFSR_26/D vdd NAND2X1
XNAND2X1_53 NAND2X1_53/A NAND2X1_42/B gnd DFFSR_22/D vdd NAND2X1
XNAND2X1_20 NAND2X1_20/A NAND2X1_20/B gnd DFFSR_10/D vdd NAND2X1
XNAND2X1_75 MUX2X1_76/B NOR2X1_29/Y gnd NAND2X1_75/Y vdd NAND2X1
XNAND2X1_97 INVX2_4/A INVX1_86/Y gnd NAND2X1_97/Y vdd NAND2X1
XFILL_20_3_2 gnd vdd FILL
XFILL_11_3_2 gnd vdd FILL
XOAI22X1_2 INVX2_5/Y OAI22X1_4/B OAI22X1_4/A OAI22X1_4/D gnd OAI22X1_2/Y vdd OAI22X1
XINVX2_11 INVX2_11/A gnd INVX2_11/Y vdd INVX2
XOAI21X1_29 BUFX4_11/Y MUX2X1_11/Y OAI21X1_29/C gnd OAI21X1_29/Y vdd OAI21X1
XOAI21X1_18 BUFX4_73/Y BUFX4_44/Y MUX2X1_6/B gnd OAI21X1_19/C vdd OAI21X1
XFILL_0_2_2 gnd vdd FILL
XFILL_8_3_2 gnd vdd FILL
XFILL_16_2_2 gnd vdd FILL
XBUFX4_62 BUFX4_63/A gnd BUFX4_62/Y vdd BUFX4
XBUFX4_73 DFFSR_1/Q gnd BUFX4_73/Y vdd BUFX4
XBUFX4_51 INVX8_1/Y gnd DFFSR_8/R vdd BUFX4
XBUFX4_40 BUFX4_36/A gnd BUFX4_40/Y vdd BUFX4
XCLKBUF1_19 BUFX4_6/Y gnd DFFSR_45/CLK vdd CLKBUF1
XBUFX4_84 BUFX4_82/A gnd BUFX4_84/Y vdd BUFX4
XBUFX4_95 BUFX4_93/A gnd AND2X2_3/A vdd BUFX4
XOR2X2_10 BUFX4_31/Y OR2X2_10/B gnd OR2X2_10/Y vdd OR2X2
XXNOR2X1_5 NOR2X1_20/Y INVX1_28/Y gnd DFFSR_35/D vdd XNOR2X1
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
.ends


magic
tech scmos
magscale 1 2
timestamp 1742918108
<< metal1 >>
rect 1768 4806 1774 4814
rect 1782 4806 1788 4814
rect 1796 4806 1802 4814
rect 1810 4806 1816 4814
rect 4824 4806 4830 4814
rect 4838 4806 4844 4814
rect 4852 4806 4858 4814
rect 4866 4806 4872 4814
rect 445 4737 460 4743
rect 1597 4743 1603 4763
rect 4900 4756 4902 4764
rect 1597 4737 1628 4743
rect 5181 4743 5187 4763
rect 5181 4737 5212 4743
rect 5284 4736 5286 4744
rect 5469 4737 5484 4743
rect 6157 4737 6172 4743
rect 589 4717 611 4723
rect 804 4716 812 4724
rect 1044 4716 1052 4724
rect 2093 4717 2115 4723
rect 2237 4717 2259 4723
rect 157 4697 179 4703
rect 237 4697 275 4703
rect 717 4697 739 4703
rect 813 4697 828 4703
rect 877 4697 899 4703
rect 1053 4697 1091 4703
rect 1108 4697 1139 4703
rect 1293 4684 1299 4703
rect 1612 4703 1620 4708
rect 1612 4697 1628 4703
rect 1693 4697 1715 4703
rect 1780 4697 1836 4703
rect 2077 4697 2092 4703
rect 2180 4697 2195 4703
rect 2445 4703 2451 4723
rect 2468 4716 2476 4724
rect 2596 4717 2611 4723
rect 2372 4697 2403 4703
rect 2413 4697 2451 4703
rect 2557 4703 2563 4716
rect 2541 4697 2563 4703
rect 2701 4697 2723 4703
rect 2808 4697 2860 4703
rect 2893 4697 2908 4703
rect 2973 4697 3011 4703
rect 3101 4703 3107 4723
rect 3044 4697 3075 4703
rect 3101 4697 3139 4703
rect 3741 4697 3763 4703
rect 717 4677 732 4683
rect 836 4677 851 4683
rect 189 4657 204 4663
rect 740 4657 755 4663
rect 845 4657 851 4677
rect 1261 4677 1292 4683
rect 1348 4677 1363 4683
rect 1773 4677 1859 4683
rect 941 4657 956 4663
rect 980 4657 995 4663
rect 1645 4657 1667 4663
rect 1700 4657 1715 4663
rect 1773 4657 1779 4677
rect 1940 4677 1955 4683
rect 1965 4677 1987 4683
rect 2029 4677 2051 4683
rect 1949 4657 1955 4677
rect 2500 4677 2531 4683
rect 2637 4677 2675 4683
rect 2845 4677 2883 4683
rect 3101 4677 3116 4683
rect 3757 4677 3763 4697
rect 3805 4703 3811 4723
rect 5581 4717 5619 4723
rect 6180 4717 6195 4723
rect 3805 4697 3843 4703
rect 4429 4697 4460 4703
rect 4701 4697 4780 4703
rect 4797 4697 4876 4703
rect 5268 4697 5283 4703
rect 5645 4697 5676 4703
rect 3805 4677 3820 4683
rect 4269 4677 4316 4683
rect 4397 4677 4419 4683
rect 3340 4663 3348 4666
rect 4397 4664 4403 4677
rect 4516 4677 4547 4683
rect 4724 4677 4771 4683
rect 5021 4677 5036 4683
rect 5357 4677 5372 4683
rect 5405 4677 5436 4683
rect 5901 4683 5907 4703
rect 5876 4677 5907 4683
rect 6116 4677 6140 4683
rect 6237 4677 6275 4683
rect 3340 4657 3411 4663
rect 4605 4657 4636 4663
rect 5108 4657 5123 4663
rect 5700 4656 5708 4664
rect 72 4636 76 4644
rect 344 4636 348 4644
rect 2356 4636 2358 4644
rect 2618 4636 2620 4644
rect 5050 4636 5052 4644
rect 5549 4637 5564 4643
rect 5844 4636 5846 4644
rect 6516 4637 6531 4643
rect 6589 4637 6636 4643
rect 3304 4606 3310 4614
rect 3318 4606 3324 4614
rect 3332 4606 3338 4614
rect 3346 4606 3352 4614
rect 618 4576 620 4584
rect 788 4576 790 4584
rect 3544 4576 3548 4584
rect 5693 4577 5708 4583
rect 5853 4577 5868 4583
rect 5914 4576 5916 4584
rect 1348 4557 1363 4563
rect 1757 4557 1772 4563
rect 1869 4557 1900 4563
rect 109 4537 124 4543
rect 749 4537 764 4543
rect 909 4537 963 4543
rect 1101 4537 1123 4543
rect 1229 4537 1267 4543
rect 349 4517 380 4523
rect 413 4517 444 4523
rect 461 4517 499 4523
rect 1005 4517 1027 4523
rect 1165 4517 1196 4523
rect 1165 4497 1171 4517
rect 1380 4517 1395 4523
rect 1524 4517 1539 4523
rect 1645 4523 1651 4543
rect 2116 4537 2131 4543
rect 2173 4537 2188 4543
rect 2237 4543 2243 4563
rect 2541 4557 2579 4563
rect 2916 4557 2931 4563
rect 2948 4557 2963 4563
rect 4356 4556 4364 4564
rect 4504 4556 4508 4564
rect 5469 4557 5491 4563
rect 5565 4557 5580 4563
rect 2228 4537 2243 4543
rect 2605 4537 2643 4543
rect 1613 4517 1651 4523
rect 1940 4517 1964 4523
rect 1981 4517 2019 4523
rect 2013 4497 2019 4517
rect 2061 4523 2067 4536
rect 2061 4517 2083 4523
rect 2317 4517 2348 4523
rect 2381 4517 2396 4523
rect 2452 4517 2467 4523
rect 2509 4517 2524 4523
rect 2605 4517 2611 4537
rect 2781 4537 2796 4543
rect 3524 4537 3544 4543
rect 3613 4537 3628 4543
rect 4388 4537 4403 4543
rect 2660 4517 2675 4523
rect 2692 4517 2723 4523
rect 2829 4517 2860 4523
rect 2948 4517 2979 4523
rect 3421 4517 3436 4523
rect 3613 4517 3651 4523
rect 2397 4497 2412 4503
rect 3252 4496 3260 4504
rect 3613 4497 3619 4517
rect 3972 4517 3987 4523
rect 4404 4517 4419 4523
rect 4724 4517 4755 4523
rect 4868 4517 4915 4523
rect 4612 4497 4627 4503
rect 4909 4503 4915 4517
rect 4973 4517 4988 4523
rect 5037 4523 5043 4543
rect 5949 4543 5955 4563
rect 5940 4537 5955 4543
rect 5972 4537 5987 4543
rect 6212 4537 6227 4543
rect 5005 4517 5043 4523
rect 5181 4517 5219 4523
rect 5341 4523 5347 4536
rect 5341 4517 5363 4523
rect 4909 4497 4931 4503
rect 5357 4497 5363 4517
rect 5533 4517 5571 4523
rect 5597 4517 5635 4523
rect 6196 4517 6243 4523
rect 6148 4497 6163 4503
rect 6404 4497 6419 4503
rect 276 4476 278 4484
rect 1549 4477 1564 4483
rect 2205 4477 2220 4483
rect 3370 4476 3372 4484
rect 6500 4477 6515 4483
rect 6548 4477 6579 4483
rect 148 4436 150 4444
rect 410 4436 412 4444
rect 712 4436 716 4444
rect 852 4436 856 4444
rect 1450 4436 1452 4444
rect 1924 4436 1926 4444
rect 2042 4436 2044 4444
rect 2596 4436 2598 4444
rect 2868 4436 2870 4444
rect 3204 4436 3206 4444
rect 5812 4436 5814 4444
rect 6052 4436 6054 4444
rect 1768 4406 1774 4414
rect 1782 4406 1788 4414
rect 1796 4406 1802 4414
rect 1810 4406 1816 4414
rect 4824 4406 4830 4414
rect 4838 4406 4844 4414
rect 4852 4406 4858 4414
rect 4866 4406 4872 4414
rect 2964 4376 2966 4384
rect 3796 4376 3798 4384
rect 4698 4376 4700 4384
rect 5044 4376 5046 4384
rect 1252 4356 1254 4364
rect 3018 4356 3020 4364
rect 1165 4337 1180 4343
rect 2250 4336 2252 4344
rect 3396 4336 3398 4344
rect 4125 4337 4140 4343
rect 5322 4336 5324 4344
rect 5610 4336 5612 4344
rect 173 4317 195 4323
rect 1780 4317 1827 4323
rect 3085 4317 3107 4323
rect 29 4297 44 4303
rect 157 4297 172 4303
rect 189 4297 227 4303
rect 1053 4297 1068 4303
rect 1284 4297 1299 4303
rect 1668 4297 1731 4303
rect 2004 4297 2019 4303
rect 3181 4297 3196 4303
rect 3261 4297 3276 4303
rect 3821 4303 3827 4323
rect 4925 4317 4940 4323
rect 3821 4297 3859 4303
rect 3917 4297 3932 4303
rect 4589 4297 4604 4303
rect 4708 4297 4755 4303
rect 5133 4303 5139 4323
rect 5293 4304 5299 4323
rect 5789 4317 5804 4323
rect 5901 4317 5932 4323
rect 6420 4317 6435 4323
rect 5101 4297 5139 4303
rect 5261 4297 5292 4303
rect 5348 4297 5363 4303
rect 5373 4297 5388 4303
rect 5581 4303 5587 4316
rect 5581 4297 5603 4303
rect 5709 4297 5756 4303
rect 5773 4297 5788 4303
rect 5885 4297 5907 4303
rect 356 4277 371 4283
rect 365 4257 371 4277
rect 2276 4277 2291 4283
rect 2669 4277 2707 4283
rect 2717 4277 2755 4283
rect 893 4257 908 4263
rect 1149 4257 1164 4263
rect 1885 4257 1907 4263
rect 1981 4257 2003 4263
rect 2036 4257 2051 4263
rect 2061 4257 2076 4263
rect 2173 4257 2188 4263
rect 2269 4257 2275 4276
rect 2548 4257 2563 4263
rect 2637 4257 2652 4263
rect 2701 4257 2707 4277
rect 2788 4277 2835 4283
rect 2925 4277 2940 4283
rect 3117 4277 3132 4283
rect 3277 4277 3292 4283
rect 4637 4277 4652 4283
rect 4724 4277 4739 4283
rect 4781 4277 4796 4283
rect 5005 4283 5011 4296
rect 5005 4277 5027 4283
rect 5341 4277 5347 4296
rect 5452 4277 5468 4283
rect 5452 4276 5460 4277
rect 5565 4277 5596 4283
rect 5684 4277 5699 4283
rect 6020 4277 6035 4283
rect 6285 4277 6316 4283
rect 4220 4272 4228 4276
rect 2781 4257 2796 4263
rect 4813 4257 4860 4263
rect 4989 4257 5004 4263
rect 5220 4256 5228 4264
rect 5668 4256 5676 4264
rect 5821 4257 5843 4263
rect 6125 4257 6147 4263
rect 6509 4257 6524 4263
rect 282 4236 284 4244
rect 500 4236 504 4244
rect 1428 4236 1432 4244
rect 1636 4236 1640 4244
rect 2906 4236 2908 4244
rect 4410 4236 4412 4244
rect 6228 4236 6230 4244
rect 6330 4236 6332 4244
rect 3304 4206 3310 4214
rect 3318 4206 3324 4214
rect 3332 4206 3338 4214
rect 3346 4206 3352 4214
rect 2794 4176 2796 4184
rect 5668 4176 5670 4184
rect 333 4157 355 4163
rect 884 4156 892 4164
rect 1709 4157 1740 4163
rect 4797 4157 4812 4163
rect 4852 4157 4915 4163
rect 5924 4156 5932 4164
rect 6068 4157 6083 4163
rect 356 4137 371 4143
rect 381 4137 451 4143
rect 589 4137 643 4143
rect 1172 4137 1187 4143
rect 1229 4137 1244 4143
rect 1284 4137 1299 4143
rect 1332 4137 1347 4143
rect 2068 4137 2099 4143
rect 2372 4137 2387 4143
rect 116 4117 131 4123
rect 797 4117 835 4123
rect 868 4117 883 4123
rect 989 4117 1004 4123
rect 877 4097 883 4117
rect 2045 4117 2076 4123
rect 2253 4117 2268 4123
rect 2397 4123 2403 4143
rect 2493 4137 2531 4143
rect 2765 4137 2780 4143
rect 2813 4137 2828 4143
rect 3629 4137 3667 4143
rect 4253 4137 4268 4143
rect 5380 4137 5395 4143
rect 6020 4137 6035 4143
rect 6093 4137 6108 4143
rect 6452 4137 6467 4143
rect 6541 4137 6579 4143
rect 2397 4117 2420 4123
rect 2412 4112 2420 4117
rect 2845 4117 2876 4123
rect 2973 4117 3011 4123
rect 3229 4117 3283 4123
rect 3293 4117 3356 4123
rect 3949 4117 4003 4123
rect 4029 4117 4067 4123
rect 4189 4117 4227 4123
rect 4253 4117 4291 4123
rect 1325 4097 1347 4103
rect 2173 4097 2195 4103
rect 4029 4097 4035 4117
rect 4253 4097 4259 4117
rect 4589 4117 4620 4123
rect 5181 4117 5219 4123
rect 4564 4097 4579 4103
rect 5213 4097 5219 4117
rect 5485 4117 5516 4123
rect 5613 4117 5644 4123
rect 6381 4117 6396 4123
rect 1284 4077 1315 4083
rect 1364 4077 1379 4083
rect 5068 4083 5076 4088
rect 5044 4077 5076 4083
rect 6284 4077 6316 4083
rect 244 4036 248 4044
rect 484 4036 488 4044
rect 1956 4036 1960 4044
rect 2308 4036 2310 4044
rect 2900 4036 2902 4044
rect 4004 4036 4006 4044
rect 5140 4036 5142 4044
rect 5540 4036 5542 4044
rect 6484 4036 6486 4044
rect 1768 4006 1774 4014
rect 1782 4006 1788 4014
rect 1796 4006 1802 4014
rect 1810 4006 1816 4014
rect 4824 4006 4830 4014
rect 4838 4006 4844 4014
rect 4852 4006 4858 4014
rect 4866 4006 4872 4014
rect 4772 3976 4774 3984
rect 5338 3976 5340 3984
rect 26 3936 28 3944
rect 493 3937 508 3943
rect 5180 3937 5235 3943
rect 5805 3937 5820 3943
rect 5180 3932 5188 3937
rect 1245 3917 1260 3923
rect 100 3897 115 3903
rect 285 3897 300 3903
rect 836 3897 851 3903
rect 861 3897 876 3903
rect 996 3897 1011 3903
rect 1140 3897 1171 3903
rect 1501 3897 1532 3903
rect 1981 3903 1987 3923
rect 2404 3916 2412 3924
rect 3293 3917 3308 3923
rect 1981 3897 2019 3903
rect 2973 3897 3011 3903
rect 3021 3897 3036 3903
rect 3156 3897 3171 3903
rect 3277 3897 3340 3903
rect 3661 3897 3715 3903
rect 4349 3897 4364 3903
rect 4429 3897 4492 3903
rect 4557 3897 4572 3903
rect 77 3877 99 3883
rect 420 3876 422 3884
rect 605 3877 620 3883
rect 1229 3877 1251 3883
rect 2036 3877 2067 3883
rect 2525 3877 2540 3883
rect 2877 3877 2892 3883
rect 3741 3877 3763 3883
rect 3853 3877 3884 3883
rect 4333 3877 4348 3883
rect 4404 3877 4419 3883
rect 4557 3877 4563 3897
rect 4621 3903 4627 3923
rect 5053 3917 5075 3923
rect 4589 3897 4627 3903
rect 4685 3897 4700 3903
rect 4733 3897 4764 3903
rect 4973 3897 5027 3903
rect 5037 3897 5052 3903
rect 5268 3897 5283 3903
rect 5453 3903 5459 3916
rect 5453 3897 5491 3903
rect 5501 3897 5532 3903
rect 5565 3897 5596 3903
rect 5869 3903 5875 3923
rect 6173 3917 6211 3923
rect 5837 3897 5875 3903
rect 6397 3897 6419 3903
rect 4829 3877 4892 3883
rect 5357 3877 5411 3883
rect 5901 3877 5923 3883
rect 6557 3883 6563 3903
rect 6548 3877 6563 3883
rect 52 3857 67 3863
rect 636 3863 644 3866
rect 621 3857 644 3863
rect 5732 3856 5740 3864
rect 6205 3857 6227 3863
rect 554 3836 556 3844
rect 1210 3836 1212 3844
rect 4164 3836 4168 3844
rect 4330 3836 4332 3844
rect 4378 3836 4380 3844
rect 4520 3836 4524 3844
rect 6580 3836 6582 3844
rect 3304 3806 3310 3814
rect 3318 3806 3324 3814
rect 3332 3806 3338 3814
rect 3346 3806 3352 3814
rect 5066 3776 5068 3784
rect 5197 3777 5212 3783
rect 6004 3776 6008 3784
rect 6548 3776 6552 3784
rect 3293 3757 3356 3763
rect 253 3737 268 3743
rect 989 3737 1004 3743
rect 2068 3737 2099 3743
rect 3469 3743 3475 3763
rect 3444 3737 3475 3743
rect 4301 3737 4316 3743
rect 4909 3737 4924 3743
rect 4957 3737 4972 3743
rect 253 3717 291 3723
rect 253 3697 259 3717
rect 557 3717 595 3723
rect 669 3717 707 3723
rect 557 3697 563 3717
rect 701 3697 707 3717
rect 1069 3717 1107 3723
rect 1133 3717 1203 3723
rect 1101 3697 1107 3717
rect 1549 3717 1564 3723
rect 2573 3717 2611 3723
rect 1628 3704 1636 3714
rect 1725 3697 1740 3703
rect 2445 3697 2483 3703
rect 2605 3697 2611 3717
rect 2772 3717 2787 3723
rect 2900 3717 2915 3723
rect 3348 3717 3363 3723
rect 4804 3717 4883 3723
rect 4957 3717 4963 3737
rect 4980 3737 4995 3743
rect 5028 3737 5052 3743
rect 5140 3737 5155 3743
rect 5261 3737 5299 3743
rect 5773 3723 5779 3743
rect 5912 3736 5916 3744
rect 6168 3736 6172 3744
rect 6493 3743 6499 3763
rect 6429 3737 6467 3743
rect 6493 3737 6508 3743
rect 5773 3717 5811 3723
rect 6372 3717 6403 3723
rect 6461 3717 6467 3737
rect 2812 3704 2820 3714
rect 3540 3696 3548 3704
rect 4205 3697 4236 3703
rect 4434 3696 4444 3704
rect 5949 3697 5987 3703
rect 6109 3697 6124 3703
rect 6292 3697 6307 3703
rect 637 3677 652 3683
rect 1748 3677 1763 3683
rect 2244 3676 2250 3684
rect 2845 3677 2860 3683
rect 4660 3677 4691 3683
rect 5620 3677 5699 3683
rect 6013 3677 6044 3683
rect 6276 3677 6300 3683
rect 532 3636 534 3644
rect 1130 3636 1132 3644
rect 1306 3636 1308 3644
rect 1450 3636 1452 3644
rect 2634 3636 2636 3644
rect 4564 3636 4566 3644
rect 5352 3636 5356 3644
rect 5754 3636 5756 3644
rect 1768 3606 1774 3614
rect 1782 3606 1788 3614
rect 1796 3606 1802 3614
rect 1810 3606 1816 3614
rect 4824 3606 4830 3614
rect 4838 3606 4844 3614
rect 4852 3606 4858 3614
rect 4866 3606 4872 3614
rect 4356 3576 4358 3584
rect 3028 3536 3030 3544
rect 6045 3543 6051 3563
rect 6045 3537 6108 3543
rect 285 3503 291 3523
rect 365 3517 403 3523
rect 420 3516 428 3524
rect 797 3517 812 3523
rect 829 3517 844 3523
rect 253 3497 291 3503
rect 957 3503 963 3523
rect 1108 3516 1112 3524
rect 2228 3517 2243 3523
rect 3364 3516 3372 3524
rect 3428 3517 3443 3523
rect 4036 3517 4051 3523
rect 4589 3517 4604 3523
rect 948 3497 963 3503
rect 1332 3497 1363 3503
rect 1693 3497 1731 3503
rect 221 3477 243 3483
rect 221 3464 227 3477
rect 276 3477 291 3483
rect 333 3477 348 3483
rect 781 3477 796 3483
rect 996 3477 1011 3483
rect 1725 3477 1731 3497
rect 2148 3497 2179 3503
rect 2532 3497 2547 3503
rect 3268 3497 3283 3503
rect 3373 3497 3411 3503
rect 3709 3497 3747 3503
rect 4317 3497 4348 3503
rect 4525 3497 4540 3503
rect 4740 3497 4755 3503
rect 5309 3497 5324 3503
rect 5677 3497 5699 3503
rect 5789 3497 5804 3503
rect 6253 3497 6291 3503
rect 1876 3477 1891 3483
rect 2036 3477 2067 3483
rect 2141 3477 2156 3483
rect 2269 3477 2284 3483
rect 2925 3477 2940 3483
rect 2996 3477 3011 3483
rect 3588 3476 3590 3484
rect 4589 3477 4611 3483
rect 4660 3477 4675 3483
rect 4724 3477 4739 3483
rect 5053 3477 5091 3483
rect 5341 3483 5347 3496
rect 5325 3477 5347 3483
rect 5373 3477 5388 3483
rect 868 3456 876 3464
rect 4004 3456 4008 3464
rect 4692 3456 4700 3464
rect 5373 3457 5379 3477
rect 5700 3477 5715 3483
rect 5741 3477 5763 3483
rect 5741 3464 5747 3477
rect 6413 3477 6451 3483
rect 5405 3457 5420 3463
rect 6333 3457 6348 3463
rect 6445 3457 6451 3477
rect 666 3436 668 3444
rect 1748 3436 1750 3444
rect 1924 3436 1928 3444
rect 2020 3436 2022 3444
rect 2308 3436 2310 3444
rect 2804 3436 2806 3444
rect 4276 3436 4278 3444
rect 4628 3436 4630 3444
rect 4916 3436 4918 3444
rect 5000 3436 5004 3444
rect 5124 3436 5128 3444
rect 5236 3436 5240 3444
rect 6532 3436 6534 3444
rect 6600 3436 6604 3444
rect 3304 3406 3310 3414
rect 3318 3406 3324 3414
rect 3332 3406 3338 3414
rect 3346 3406 3352 3414
rect 660 3376 662 3384
rect 938 3376 940 3384
rect 2548 3376 2550 3384
rect 4989 3377 5004 3383
rect 5176 3376 5180 3384
rect 5405 3377 5420 3383
rect 332 3357 355 3363
rect 332 3354 340 3357
rect 5796 3356 5804 3364
rect 893 3337 924 3343
rect 1021 3337 1036 3343
rect 1260 3343 1268 3348
rect 1260 3337 1283 3343
rect 1652 3337 1683 3343
rect 1693 3337 1708 3343
rect 1780 3337 1827 3343
rect 2164 3337 2179 3343
rect 3172 3337 3188 3343
rect 3412 3337 3427 3343
rect 3965 3337 3980 3343
rect 4520 3336 4524 3344
rect 4920 3337 4940 3343
rect 5357 3337 5372 3343
rect 5884 3343 5892 3344
rect 5821 3337 5859 3343
rect 5884 3337 5900 3343
rect 5949 3337 5980 3343
rect 6013 3343 6019 3363
rect 6013 3337 6044 3343
rect 221 3317 236 3323
rect 365 3317 380 3323
rect 468 3317 499 3323
rect 509 3317 524 3323
rect 452 3296 460 3304
rect 493 3297 499 3317
rect 1021 3317 1059 3323
rect 1021 3297 1027 3317
rect 1293 3317 1331 3323
rect 1357 3317 1372 3323
rect 1325 3297 1331 3317
rect 1757 3317 1804 3323
rect 1860 3317 1891 3323
rect 1348 3296 1356 3304
rect 1885 3297 1891 3317
rect 2141 3317 2179 3323
rect 2173 3297 2179 3317
rect 2445 3317 2483 3323
rect 2589 3317 2627 3323
rect 2637 3317 2652 3323
rect 2772 3317 2787 3323
rect 2893 3317 2931 3323
rect 3908 3317 3939 3323
rect 3949 3317 3996 3323
rect 4221 3317 4236 3323
rect 5485 3317 5523 3323
rect 2884 3296 2892 3304
rect 4292 3297 4307 3303
rect 4429 3297 4444 3303
rect 5085 3297 5139 3303
rect 5517 3297 5523 3317
rect 5533 3297 5571 3303
rect 5917 3297 5932 3303
rect 6148 3296 6156 3304
rect 6237 3297 6252 3303
rect 413 3277 436 3283
rect 1924 3277 1939 3283
rect 2413 3277 2428 3283
rect 3812 3277 3827 3283
rect 3844 3277 3891 3283
rect 4004 3276 4006 3284
rect 4628 3277 4707 3283
rect 4989 3277 5004 3283
rect 1412 3236 1414 3244
rect 1626 3236 1628 3244
rect 4074 3236 4076 3244
rect 5736 3236 5740 3244
rect 1768 3206 1774 3214
rect 1782 3206 1788 3214
rect 1796 3206 1802 3214
rect 1810 3206 1816 3214
rect 4824 3206 4830 3214
rect 4838 3206 4844 3214
rect 4852 3206 4858 3214
rect 4866 3206 4872 3214
rect 570 3176 572 3184
rect 1208 3176 1212 3184
rect 3098 3176 3100 3184
rect 4845 3177 4892 3183
rect 4077 3137 4092 3143
rect 4804 3137 4835 3143
rect 5549 3137 5580 3143
rect 5677 3137 5708 3143
rect 5818 3136 5820 3144
rect 5962 3136 5964 3144
rect 1012 3116 1020 3124
rect 1277 3117 1292 3123
rect 1588 3117 1603 3123
rect 253 3097 300 3103
rect 525 3097 563 3103
rect 717 3097 732 3103
rect 1021 3097 1052 3103
rect 1309 3097 1340 3103
rect 1453 3097 1500 3103
rect 2301 3097 2316 3103
rect 2557 3103 2563 3123
rect 2525 3097 2563 3103
rect 2589 3097 2627 3103
rect 3069 3103 3075 3123
rect 4788 3117 4803 3123
rect 5581 3117 5596 3123
rect 6045 3117 6060 3123
rect 3037 3097 3075 3103
rect 3165 3097 3203 3103
rect 3533 3097 3548 3103
rect 4132 3097 4147 3103
rect 4180 3097 4211 3103
rect 4525 3097 4547 3103
rect 4957 3097 4972 3103
rect 5277 3097 5324 3103
rect 5501 3097 5516 3103
rect 5773 3097 5788 3103
rect 1332 3077 1347 3083
rect 1640 3077 1667 3083
rect 4173 3077 4195 3083
rect 4445 3077 4483 3083
rect 3213 3057 3260 3063
rect 3780 3056 3788 3064
rect 3860 3057 3884 3063
rect 4020 3056 4028 3064
rect 4253 3057 4291 3063
rect 4477 3057 4483 3077
rect 5197 3077 5228 3083
rect 5437 3077 5452 3083
rect 5469 3077 5491 3083
rect 6140 3077 6156 3083
rect 6140 3076 6148 3077
rect 680 3036 684 3044
rect 1066 3036 1068 3044
rect 3044 3036 3046 3044
rect 3956 3036 3958 3044
rect 5352 3036 5356 3044
rect 5640 3036 5644 3044
rect 5677 3037 5692 3043
rect 6564 3036 6568 3044
rect 3304 3006 3310 3014
rect 3318 3006 3324 3014
rect 3332 3006 3338 3014
rect 3346 3006 3352 3014
rect 228 2976 230 2984
rect 1172 2976 1176 2984
rect 4216 2976 4220 2984
rect 724 2956 728 2964
rect 1293 2957 1320 2963
rect 2868 2957 2883 2963
rect 5380 2956 5388 2964
rect 5764 2956 5772 2964
rect 5912 2957 5939 2963
rect 28 2943 36 2944
rect 28 2937 44 2943
rect 156 2943 164 2944
rect 156 2937 172 2943
rect 436 2937 451 2943
rect 573 2937 604 2943
rect 877 2937 899 2943
rect 956 2943 964 2944
rect 948 2937 964 2943
rect 1076 2937 1107 2943
rect 1556 2937 1571 2943
rect 1972 2937 1987 2943
rect 2797 2937 2828 2943
rect 4477 2937 4508 2943
rect 4840 2937 4876 2943
rect 5037 2937 5052 2943
rect 5736 2937 5756 2943
rect 5796 2937 5827 2943
rect 6013 2937 6028 2943
rect 6308 2936 6310 2944
rect 429 2917 444 2923
rect 836 2917 867 2923
rect 916 2917 932 2923
rect 924 2912 932 2917
rect 1108 2917 1123 2923
rect 1885 2917 1923 2923
rect 2276 2917 2291 2923
rect 2365 2917 2403 2923
rect 2493 2917 2508 2923
rect 3012 2917 3027 2923
rect 3117 2917 3155 2923
rect 3165 2917 3180 2923
rect 3396 2917 3443 2923
rect 3517 2917 3555 2923
rect 4068 2917 4099 2923
rect 4109 2917 4131 2923
rect 4605 2917 4620 2923
rect 4637 2917 4652 2923
rect 4957 2917 4972 2923
rect 4989 2917 5020 2923
rect 5325 2917 5356 2923
rect 5453 2917 5468 2923
rect 5629 2917 5644 2923
rect 5949 2917 5987 2923
rect 925 2897 940 2903
rect 1021 2897 1043 2903
rect 1149 2897 1171 2903
rect 1268 2897 1283 2903
rect 2029 2897 2051 2903
rect 2420 2897 2435 2903
rect 4322 2896 4332 2904
rect 4621 2897 4643 2903
rect 4900 2897 4915 2903
rect 5122 2896 5132 2904
rect 5645 2897 5660 2903
rect 5677 2897 5699 2903
rect 6141 2897 6163 2903
rect 1020 2884 1028 2888
rect 260 2877 275 2883
rect 269 2857 275 2877
rect 324 2877 355 2883
rect 509 2877 524 2883
rect 1228 2883 1236 2888
rect 1181 2877 1236 2883
rect 1325 2877 1356 2883
rect 4717 2877 4748 2883
rect 6100 2877 6131 2883
rect 3802 2856 3804 2864
rect 1124 2836 1126 2844
rect 4532 2836 4534 2844
rect 1768 2806 1774 2814
rect 1782 2806 1788 2814
rect 1796 2806 1802 2814
rect 1810 2806 1816 2814
rect 4824 2806 4830 2814
rect 4838 2806 4844 2814
rect 4852 2806 4858 2814
rect 4866 2806 4872 2814
rect 72 2776 76 2784
rect 500 2776 502 2784
rect 1124 2776 1126 2784
rect 1220 2776 1222 2784
rect 1322 2776 1324 2784
rect 1448 2776 1452 2784
rect 861 2743 867 2763
rect 2106 2756 2108 2764
rect 861 2737 892 2743
rect 2618 2736 2620 2744
rect 4077 2737 4092 2743
rect 653 2717 675 2723
rect 1149 2717 1180 2723
rect 1773 2717 1836 2723
rect 3028 2716 3036 2724
rect 253 2703 259 2716
rect 237 2697 259 2703
rect 461 2697 476 2703
rect 484 2697 492 2703
rect 532 2697 547 2703
rect 700 2703 708 2708
rect 692 2697 708 2703
rect 1709 2697 1747 2703
rect 1853 2697 1891 2703
rect 2013 2697 2051 2703
rect 2308 2697 2323 2703
rect 2621 2697 2636 2703
rect 2932 2697 2947 2703
rect 3060 2697 3091 2703
rect 3181 2697 3203 2703
rect 109 2677 147 2683
rect 157 2677 172 2683
rect 413 2677 451 2683
rect 1092 2677 1107 2683
rect 1676 2677 1692 2683
rect 2820 2677 2851 2683
rect 3197 2677 3203 2697
rect 3245 2703 3251 2723
rect 3437 2717 3460 2723
rect 3452 2712 3460 2717
rect 4333 2717 4348 2723
rect 4468 2716 4476 2724
rect 3245 2697 3260 2703
rect 3293 2697 3379 2703
rect 4164 2697 4195 2703
rect 4212 2697 4227 2703
rect 4397 2697 4419 2703
rect 4109 2677 4124 2683
rect 4253 2677 4268 2683
rect 260 2656 268 2664
rect 1796 2657 1843 2663
rect 2813 2657 2828 2663
rect 4253 2657 4259 2677
rect 4285 2677 4316 2683
rect 4333 2677 4355 2683
rect 4413 2677 4419 2697
rect 4525 2697 4563 2703
rect 4996 2697 5043 2703
rect 5053 2697 5068 2703
rect 4605 2677 4643 2683
rect 6292 2676 6294 2684
rect 5021 2657 5036 2663
rect 138 2636 140 2644
rect 6605 2637 6620 2643
rect 3304 2606 3310 2614
rect 3318 2606 3324 2614
rect 3332 2606 3338 2614
rect 3346 2606 3352 2614
rect 36 2576 38 2584
rect 618 2576 620 2584
rect 676 2576 678 2584
rect 714 2576 716 2584
rect 1114 2576 1116 2584
rect 116 2537 136 2543
rect 381 2543 387 2563
rect 1181 2557 1196 2563
rect 349 2537 387 2543
rect 413 2537 444 2543
rect 461 2537 476 2543
rect 212 2517 227 2523
rect 557 2523 563 2543
rect 637 2537 652 2543
rect 781 2537 812 2543
rect 1021 2537 1075 2543
rect 1133 2537 1171 2543
rect 1389 2543 1395 2563
rect 1660 2557 1692 2563
rect 1660 2548 1668 2557
rect 1380 2537 1395 2543
rect 1804 2537 1852 2543
rect 2093 2537 2108 2543
rect 2244 2537 2260 2543
rect 2605 2537 2620 2543
rect 2701 2543 2707 2563
rect 2692 2537 2707 2543
rect 2813 2537 2828 2543
rect 532 2517 563 2523
rect 740 2517 755 2523
rect 852 2517 915 2523
rect 1069 2517 1107 2523
rect 84 2497 99 2503
rect 141 2497 163 2503
rect 477 2497 492 2503
rect 1101 2497 1107 2517
rect 1140 2517 1155 2523
rect 1236 2517 1251 2523
rect 1693 2517 1708 2523
rect 2573 2517 2611 2523
rect 2765 2517 2796 2523
rect 3181 2523 3187 2543
rect 3229 2537 3244 2543
rect 3277 2537 3324 2543
rect 4061 2537 4076 2543
rect 4317 2537 4348 2543
rect 4381 2537 4396 2543
rect 4413 2543 4419 2563
rect 4429 2557 4444 2563
rect 5261 2557 5276 2563
rect 6061 2557 6083 2563
rect 4404 2537 4419 2543
rect 4452 2537 4467 2543
rect 3172 2517 3187 2523
rect 3229 2517 3267 2523
rect 3229 2497 3235 2517
rect 3613 2517 3651 2523
rect 4068 2517 4083 2523
rect 4125 2517 4147 2523
rect 4189 2517 4204 2523
rect 4244 2517 4259 2523
rect 4461 2517 4467 2537
rect 4909 2537 4924 2543
rect 4532 2517 4547 2523
rect 4685 2517 4716 2523
rect 4973 2523 4979 2543
rect 5069 2537 5107 2543
rect 5188 2537 5219 2543
rect 5956 2536 5958 2544
rect 6116 2536 6124 2544
rect 6189 2543 6195 2563
rect 6157 2537 6195 2543
rect 4813 2517 4899 2523
rect 4941 2517 4979 2523
rect 5181 2517 5196 2523
rect 4612 2496 4620 2504
rect 4813 2497 4819 2517
rect 5229 2517 5283 2523
rect 5428 2517 5443 2523
rect 6109 2517 6115 2536
rect 4916 2497 4931 2503
rect 6068 2497 6083 2503
rect 2733 2477 2748 2483
rect 4548 2456 4550 2464
rect 186 2436 188 2444
rect 522 2436 524 2444
rect 1258 2436 1260 2444
rect 2516 2436 2518 2444
rect 2938 2436 2940 2444
rect 3978 2436 3980 2444
rect 5012 2436 5016 2444
rect 1768 2406 1774 2414
rect 1782 2406 1788 2414
rect 1796 2406 1802 2414
rect 1810 2406 1816 2414
rect 4824 2406 4830 2414
rect 4838 2406 4844 2414
rect 4852 2406 4858 2414
rect 4866 2406 4872 2414
rect 4260 2376 4262 2384
rect 356 2337 380 2343
rect 442 2336 444 2344
rect 500 2336 502 2344
rect 1828 2336 1834 2344
rect 2900 2337 2915 2343
rect 3380 2336 3382 2344
rect 5300 2336 5302 2344
rect 5862 2336 5868 2344
rect 269 2317 284 2323
rect 532 2317 547 2323
rect 708 2317 739 2323
rect 156 2303 164 2308
rect 141 2297 164 2303
rect 445 2297 492 2303
rect 532 2297 563 2303
rect 1076 2297 1091 2303
rect 1229 2303 1235 2323
rect 1268 2317 1283 2323
rect 1604 2316 1612 2324
rect 1629 2317 1644 2323
rect 2036 2316 2044 2324
rect 1197 2297 1235 2303
rect 1309 2297 1340 2303
rect 1444 2297 1459 2303
rect 1565 2297 1603 2303
rect 1661 2297 1699 2303
rect 1997 2297 2035 2303
rect 2093 2297 2131 2303
rect 2237 2297 2252 2303
rect 2381 2297 2419 2303
rect 2509 2303 2515 2323
rect 2621 2303 2627 2323
rect 2509 2297 2547 2303
rect 2589 2297 2627 2303
rect 2724 2297 2755 2303
rect 2765 2297 2851 2303
rect 3364 2297 3379 2303
rect 3869 2297 3923 2303
rect 3933 2297 3964 2303
rect 52 2277 67 2283
rect 61 2257 67 2277
rect 468 2277 483 2283
rect 980 2277 995 2283
rect 1261 2277 1283 2283
rect 1373 2277 1395 2283
rect 1373 2264 1379 2277
rect 2669 2277 2707 2283
rect 2989 2277 3043 2283
rect 3165 2277 3212 2283
rect 3277 2277 3356 2283
rect 3469 2277 3484 2283
rect 4013 2283 4019 2303
rect 4420 2297 4435 2303
rect 4445 2297 4476 2303
rect 4621 2303 4627 2323
rect 4621 2297 4659 2303
rect 5325 2303 5331 2323
rect 6013 2317 6028 2323
rect 5261 2297 5299 2303
rect 5325 2297 5363 2303
rect 5468 2303 5476 2308
rect 5468 2297 5491 2303
rect 5485 2284 5491 2297
rect 5933 2297 5987 2303
rect 5997 2297 6012 2303
rect 6477 2297 6508 2303
rect 3981 2277 4019 2283
rect 4029 2277 4067 2283
rect 4125 2277 4163 2283
rect 4493 2277 4515 2283
rect 4557 2277 4579 2283
rect 4621 2277 4636 2283
rect 4884 2277 4932 2283
rect 5220 2277 5251 2283
rect 77 2257 99 2263
rect 1236 2256 1244 2264
rect 1348 2257 1363 2263
rect 3901 2257 3916 2263
rect 4084 2257 4108 2263
rect 4189 2257 4211 2263
rect 4468 2257 4483 2263
rect 5245 2257 5251 2277
rect 5956 2277 5971 2283
rect 6045 2277 6067 2283
rect 6100 2277 6131 2283
rect 6013 2257 6035 2263
rect 916 2236 918 2244
rect 1012 2236 1014 2244
rect 1725 2237 1772 2243
rect 2938 2236 2940 2244
rect 5188 2236 5190 2244
rect 6084 2236 6086 2244
rect 3304 2206 3310 2214
rect 3318 2206 3324 2214
rect 3332 2206 3338 2214
rect 3346 2206 3352 2214
rect 506 2176 508 2184
rect 1396 2176 1398 2184
rect 925 2157 947 2163
rect 1021 2157 1043 2163
rect 2820 2157 2835 2163
rect 2948 2157 2963 2163
rect 6125 2157 6147 2163
rect 6468 2157 6483 2163
rect 248 2136 252 2144
rect 509 2137 547 2143
rect 877 2137 915 2143
rect 612 2117 627 2123
rect 877 2117 883 2137
rect 1085 2137 1100 2143
rect 1352 2137 1379 2143
rect 2324 2137 2339 2143
rect 2788 2137 2803 2143
rect 3005 2137 3036 2143
rect 3053 2137 3100 2143
rect 3293 2137 3395 2143
rect 3964 2143 3972 2148
rect 3964 2137 3987 2143
rect 4077 2137 4099 2143
rect 4237 2137 4252 2143
rect 4324 2137 4339 2143
rect 4493 2137 4508 2143
rect 5428 2137 5443 2143
rect 5517 2137 5539 2143
rect 5636 2137 5651 2143
rect 5933 2137 5955 2143
rect 6493 2143 6499 2156
rect 6340 2137 6355 2143
rect 6493 2137 6515 2143
rect 941 2117 979 2123
rect 1092 2117 1123 2123
rect 1277 2117 1292 2123
rect 2301 2117 2339 2123
rect 189 2097 211 2103
rect 317 2097 332 2103
rect 701 2097 739 2103
rect 2333 2097 2339 2117
rect 2461 2117 2492 2123
rect 2820 2117 2851 2123
rect 3197 2117 3219 2123
rect 2540 2104 2548 2114
rect 3213 2104 3219 2117
rect 3629 2117 3667 2123
rect 3693 2117 3747 2123
rect 3661 2097 3667 2117
rect 3892 2117 3907 2123
rect 3997 2117 4028 2123
rect 4301 2123 4307 2136
rect 4285 2117 4307 2123
rect 4493 2117 4531 2123
rect 4493 2097 4499 2117
rect 5268 2117 5283 2123
rect 5565 2117 5596 2123
rect 5885 2117 5916 2123
rect 5956 2117 5971 2123
rect 6029 2117 6060 2123
rect 6077 2117 6099 2123
rect 4732 2103 4740 2108
rect 4732 2097 4755 2103
rect 5245 2097 5267 2103
rect 5380 2097 5395 2103
rect 1204 2076 1206 2084
rect 5357 2077 5372 2083
rect 6381 2077 6412 2083
rect 1156 2036 1158 2044
rect 2884 2036 2886 2044
rect 3060 2036 3062 2044
rect 4132 2036 4136 2044
rect 4964 2036 4968 2044
rect 5076 2036 5080 2044
rect 5172 2036 5174 2044
rect 5460 2036 5462 2044
rect 5972 2036 5974 2044
rect 6532 2036 6534 2044
rect 1768 2006 1774 2014
rect 1782 2006 1788 2014
rect 1796 2006 1802 2014
rect 1810 2006 1816 2014
rect 4824 2006 4830 2014
rect 4838 2006 4844 2014
rect 4852 2006 4858 2014
rect 4866 2006 4872 2014
rect 3066 1976 3068 1984
rect 3194 1976 3196 1984
rect 1117 1937 1140 1943
rect 1373 1937 1427 1943
rect 5028 1936 5030 1944
rect 5693 1937 5708 1943
rect 132 1917 147 1923
rect 317 1917 332 1923
rect 484 1916 492 1924
rect 1613 1917 1628 1923
rect 1908 1917 1923 1923
rect 564 1897 579 1903
rect 653 1883 659 1903
rect 845 1897 860 1903
rect 1460 1897 1475 1903
rect 1485 1897 1507 1903
rect 1981 1897 2019 1903
rect 628 1877 659 1883
rect 861 1877 876 1883
rect 1069 1877 1091 1883
rect 877 1857 883 1876
rect 1085 1864 1091 1877
rect 1236 1877 1244 1883
rect 1677 1883 1683 1896
rect 2797 1897 2812 1903
rect 2941 1897 2956 1903
rect 3021 1897 3052 1903
rect 3165 1903 3171 1923
rect 4692 1916 4700 1924
rect 5170 1916 5180 1924
rect 3133 1897 3171 1903
rect 3204 1897 3235 1903
rect 3268 1897 3283 1903
rect 3373 1897 3411 1903
rect 3556 1897 3571 1903
rect 3837 1897 3852 1903
rect 4004 1897 4019 1903
rect 4516 1897 4531 1903
rect 4797 1903 4803 1916
rect 4781 1897 4803 1903
rect 4996 1897 5027 1903
rect 5245 1897 5260 1903
rect 5277 1897 5292 1903
rect 5389 1903 5395 1923
rect 5620 1917 5635 1923
rect 5917 1917 5932 1923
rect 6132 1916 6140 1924
rect 6445 1917 6460 1923
rect 5389 1897 5427 1903
rect 5773 1897 5804 1903
rect 6020 1897 6035 1903
rect 6141 1897 6179 1903
rect 1661 1877 1683 1883
rect 3085 1877 3100 1883
rect 1229 1857 1235 1876
rect 2348 1872 2356 1876
rect 2964 1857 2979 1863
rect 3085 1857 3091 1877
rect 3268 1877 3299 1883
rect 3332 1877 3379 1883
rect 4036 1877 4051 1883
rect 4829 1877 4876 1883
rect 5213 1877 5235 1883
rect 5229 1864 5235 1877
rect 5389 1877 5404 1883
rect 5572 1877 5587 1883
rect 5661 1877 5699 1883
rect 5725 1877 5740 1883
rect 5917 1877 5955 1883
rect 3236 1857 3251 1863
rect 3261 1857 3276 1863
rect 3309 1857 3340 1863
rect 3389 1857 3404 1863
rect 4900 1857 4915 1863
rect 5917 1857 5923 1877
rect 6004 1877 6051 1883
rect 6173 1877 6211 1883
rect 6276 1877 6291 1883
rect 5949 1857 5971 1863
rect 248 1836 252 1844
rect 596 1836 598 1844
rect 788 1836 790 1844
rect 1604 1836 1606 1844
rect 1700 1836 1702 1844
rect 1828 1836 1830 1844
rect 2872 1836 2876 1844
rect 4084 1836 4088 1844
rect 4810 1836 4812 1844
rect 6468 1837 6483 1843
rect 3304 1806 3310 1814
rect 3318 1806 3324 1814
rect 3332 1806 3338 1814
rect 3346 1806 3352 1814
rect 666 1776 668 1784
rect 4516 1776 4518 1784
rect 5464 1776 5468 1784
rect 388 1757 419 1763
rect 1012 1757 1036 1763
rect 5764 1756 5772 1764
rect 52 1737 83 1743
rect 116 1737 131 1743
rect 196 1737 211 1743
rect 493 1737 508 1743
rect 29 1717 67 1723
rect 109 1717 124 1723
rect 685 1723 691 1743
rect 964 1737 995 1743
rect 1501 1737 1532 1743
rect 477 1717 531 1723
rect 589 1717 627 1723
rect 685 1717 708 1723
rect 356 1697 371 1703
rect 589 1697 595 1717
rect 700 1712 708 1717
rect 1501 1717 1507 1737
rect 1748 1737 1827 1743
rect 2028 1737 2052 1743
rect 2612 1737 2627 1743
rect 2925 1737 2940 1743
rect 3037 1737 3075 1743
rect 3108 1737 3155 1743
rect 3373 1737 3411 1743
rect 3421 1737 3475 1743
rect 3501 1737 3539 1743
rect 4589 1737 4604 1743
rect 5085 1737 5107 1743
rect 2109 1717 2124 1723
rect 2589 1717 2627 1723
rect 621 1697 659 1703
rect 1197 1697 1212 1703
rect 1389 1697 1404 1703
rect 1565 1697 1587 1703
rect 1796 1697 1811 1703
rect 2621 1697 2627 1717
rect 3229 1717 3260 1723
rect 3277 1717 3356 1723
rect 4340 1717 4387 1723
rect 4573 1717 4620 1723
rect 4660 1717 4675 1723
rect 4836 1717 4883 1723
rect 5085 1717 5091 1737
rect 5101 1712 5107 1737
rect 5332 1737 5347 1743
rect 6317 1737 6339 1743
rect 5869 1717 5884 1723
rect 5949 1717 5971 1723
rect 4692 1697 4707 1703
rect 5885 1697 5900 1703
rect 6557 1697 6579 1703
rect 788 1677 803 1683
rect 1357 1677 1436 1683
rect 4708 1677 4739 1683
rect 5140 1676 5142 1684
rect 6116 1677 6172 1683
rect 6356 1677 6387 1683
rect 6564 1677 6579 1683
rect 1092 1636 1094 1644
rect 1492 1636 1494 1644
rect 1684 1636 1688 1644
rect 3940 1636 3944 1644
rect 4052 1636 4056 1644
rect 4570 1636 4572 1644
rect 4628 1636 4630 1644
rect 4968 1636 4972 1644
rect 5194 1636 5196 1644
rect 5624 1636 5628 1644
rect 1768 1606 1774 1614
rect 1782 1606 1788 1614
rect 1796 1606 1802 1614
rect 1810 1606 1816 1614
rect 4824 1606 4830 1614
rect 4838 1606 4844 1614
rect 4852 1606 4858 1614
rect 4866 1606 4872 1614
rect 634 1576 636 1584
rect 692 1576 694 1584
rect 3290 1576 3292 1584
rect 5322 1576 5324 1584
rect 980 1536 982 1544
rect 4024 1536 4028 1544
rect 4493 1537 4524 1543
rect 4573 1537 4620 1543
rect 4492 1524 4500 1528
rect 164 1517 179 1523
rect 660 1497 684 1503
rect 724 1497 739 1503
rect 797 1497 851 1503
rect 989 1497 1027 1503
rect 1181 1497 1196 1503
rect 1357 1503 1363 1523
rect 1965 1517 1980 1523
rect 2020 1517 2035 1523
rect 3180 1517 3203 1523
rect 3389 1517 3404 1523
rect 3180 1512 3188 1517
rect 4125 1517 4140 1523
rect 4205 1517 4227 1523
rect 1348 1497 1363 1503
rect 1469 1497 1484 1503
rect 1492 1497 1523 1503
rect 1581 1497 1635 1503
rect 1972 1497 2003 1503
rect 2237 1497 2252 1503
rect 2308 1497 2323 1503
rect 2628 1497 2659 1503
rect 2845 1497 2867 1503
rect 3332 1497 3395 1503
rect 3421 1497 3436 1503
rect 3613 1497 3644 1503
rect 3757 1497 3795 1503
rect 4412 1503 4420 1508
rect 4412 1497 4435 1503
rect 365 1477 403 1483
rect 397 1457 403 1477
rect 1284 1477 1299 1483
rect 1485 1477 1500 1483
rect 2077 1477 2092 1483
rect 2932 1477 2947 1483
rect 3469 1477 3484 1483
rect 3629 1477 3644 1483
rect 900 1456 904 1464
rect 2461 1457 2492 1463
rect 2596 1456 2604 1464
rect 3309 1457 3324 1463
rect 3629 1457 3635 1477
rect 3661 1477 3676 1483
rect 4429 1477 4435 1497
rect 4573 1497 4579 1537
rect 4700 1537 4732 1543
rect 4700 1532 4708 1537
rect 5453 1537 5484 1543
rect 5652 1536 5654 1544
rect 6042 1536 6044 1544
rect 6260 1537 6284 1543
rect 6340 1537 6403 1543
rect 6396 1524 6404 1528
rect 4605 1517 4620 1523
rect 6196 1516 6204 1524
rect 5348 1497 5363 1503
rect 5421 1497 5443 1503
rect 5572 1497 5644 1503
rect 5780 1497 5804 1503
rect 6084 1497 6099 1503
rect 6205 1497 6220 1503
rect 5005 1477 5043 1483
rect 3924 1456 3932 1464
rect 4100 1456 4108 1464
rect 4285 1457 4307 1463
rect 4829 1457 4844 1463
rect 5005 1457 5011 1477
rect 5581 1477 5628 1483
rect 6148 1477 6163 1483
rect 6317 1457 6332 1463
rect 468 1436 470 1444
rect 1044 1436 1046 1444
rect 1220 1436 1224 1444
rect 1300 1436 1302 1444
rect 1588 1436 1590 1444
rect 1748 1436 1750 1444
rect 1860 1436 1864 1444
rect 1956 1436 1958 1444
rect 2724 1436 2726 1444
rect 3834 1436 3836 1444
rect 4168 1436 4172 1444
rect 4234 1436 4236 1444
rect 4692 1436 4694 1444
rect 4760 1436 4764 1444
rect 5402 1436 5404 1444
rect 6388 1437 6403 1443
rect 6580 1437 6595 1443
rect 3304 1406 3310 1414
rect 3318 1406 3324 1414
rect 3332 1406 3338 1414
rect 3346 1406 3352 1414
rect 154 1376 156 1384
rect 202 1376 204 1384
rect 260 1377 275 1383
rect 868 1377 883 1383
rect 2186 1376 2188 1384
rect 4090 1376 4092 1384
rect 4340 1376 4344 1384
rect 6404 1376 6408 1384
rect 2717 1357 2739 1363
rect 3316 1357 3379 1363
rect 3453 1357 3468 1363
rect 3533 1357 3548 1363
rect 28 1343 36 1344
rect 28 1337 44 1343
rect 733 1337 764 1343
rect 772 1337 787 1343
rect 669 1323 675 1336
rect 669 1317 691 1323
rect 717 1317 796 1323
rect 685 1297 691 1317
rect 909 1323 915 1343
rect 1133 1337 1148 1343
rect 1780 1337 1843 1343
rect 1853 1337 1868 1343
rect 2080 1343 2092 1344
rect 2045 1337 2092 1343
rect 2080 1336 2092 1337
rect 2429 1337 2444 1343
rect 2628 1337 2643 1343
rect 2717 1337 2732 1343
rect 3693 1337 3708 1343
rect 3757 1343 3763 1356
rect 3741 1337 3763 1343
rect 3965 1343 3971 1356
rect 3949 1337 3971 1343
rect 4004 1337 4019 1343
rect 4196 1337 4227 1343
rect 909 1317 932 1323
rect 924 1312 932 1317
rect 1069 1317 1084 1323
rect 1124 1317 1171 1323
rect 1668 1317 1699 1323
rect 1940 1317 1971 1323
rect 1981 1317 2019 1323
rect 2237 1317 2275 1323
rect 2372 1317 2403 1323
rect 2420 1317 2467 1323
rect 2500 1317 2531 1323
rect 2548 1317 2563 1323
rect 2765 1317 2796 1323
rect 2877 1317 2940 1323
rect 3060 1317 3091 1323
rect 3284 1317 3363 1323
rect 3373 1317 3404 1323
rect 3725 1317 3756 1323
rect 3997 1317 4012 1323
rect 4509 1317 4524 1323
rect 4797 1323 4803 1343
rect 4973 1337 4988 1343
rect 5028 1337 5059 1343
rect 5149 1343 5155 1363
rect 5293 1357 5308 1363
rect 5124 1337 5155 1343
rect 5549 1343 5555 1363
rect 5549 1337 5564 1343
rect 4685 1317 4723 1323
rect 4797 1317 4860 1323
rect 1373 1297 1395 1303
rect 1764 1297 1820 1303
rect 2493 1297 2499 1316
rect 4157 1297 4211 1303
rect 4244 1297 4259 1303
rect 4525 1297 4540 1303
rect 4717 1297 4723 1317
rect 5389 1317 5436 1323
rect 5613 1317 5644 1323
rect 4733 1297 4771 1303
rect 4884 1296 4892 1304
rect 5453 1297 5475 1303
rect 5613 1297 5619 1317
rect 5892 1317 5907 1323
rect 5917 1317 5932 1323
rect 5933 1297 5948 1303
rect 6029 1297 6051 1303
rect 6516 1297 6547 1303
rect 1388 1284 1396 1288
rect 1517 1277 1548 1283
rect 1917 1277 1932 1283
rect 2093 1277 2147 1283
rect 3146 1276 3148 1284
rect 3482 1276 3484 1284
rect 3820 1283 3828 1288
rect 3820 1277 3875 1283
rect 4564 1277 4579 1283
rect 4781 1277 4844 1283
rect 3988 1256 3990 1264
rect 1114 1236 1116 1244
rect 1172 1236 1174 1244
rect 1604 1236 1608 1244
rect 2276 1236 2278 1244
rect 2468 1236 2470 1244
rect 2874 1236 2876 1244
rect 3098 1236 3100 1244
rect 3274 1236 3276 1244
rect 3930 1236 3932 1244
rect 4436 1236 4438 1244
rect 5172 1236 5174 1244
rect 1768 1206 1774 1214
rect 1782 1206 1788 1214
rect 1796 1206 1802 1214
rect 1810 1206 1816 1214
rect 4824 1206 4830 1214
rect 4838 1206 4844 1214
rect 4852 1206 4858 1214
rect 4866 1206 4872 1214
rect 644 1136 646 1144
rect 2196 1137 2211 1143
rect 3028 1136 3030 1144
rect 4404 1137 4419 1143
rect 6621 1137 6643 1143
rect 5900 1132 5908 1136
rect 6637 1124 6643 1137
rect 84 1097 99 1103
rect 541 1103 547 1123
rect 2621 1117 2643 1123
rect 2749 1117 2764 1123
rect 2797 1117 2819 1123
rect 3076 1116 3084 1124
rect 3517 1117 3539 1123
rect 500 1097 515 1103
rect 541 1097 579 1103
rect 509 1077 515 1097
rect 596 1097 643 1103
rect 804 1097 835 1103
rect 1892 1097 1907 1103
rect 2340 1097 2355 1103
rect 2541 1097 2556 1103
rect 2564 1097 2595 1103
rect 2909 1097 2924 1103
rect 3197 1097 3219 1103
rect 3380 1097 3411 1103
rect 3580 1103 3588 1108
rect 3677 1103 3683 1123
rect 3917 1117 3932 1123
rect 3580 1097 3603 1103
rect 3677 1097 3715 1103
rect 605 1077 620 1083
rect 861 1083 867 1096
rect 845 1077 867 1083
rect 1197 1077 1235 1083
rect 772 1056 780 1064
rect 1197 1057 1203 1077
rect 1380 1077 1395 1083
rect 1476 1077 1507 1083
rect 1677 1083 1683 1096
rect 1613 1077 1651 1083
rect 1661 1077 1683 1083
rect 1837 1077 1852 1083
rect 1885 1077 1912 1083
rect 2045 1077 2060 1083
rect 2333 1077 2339 1096
rect 2436 1077 2451 1083
rect 2461 1077 2499 1083
rect 2557 1077 2572 1083
rect 2733 1077 2771 1083
rect 2884 1077 2899 1083
rect 3101 1077 3116 1083
rect 3204 1077 3219 1083
rect 3544 1076 3548 1084
rect 3597 1077 3603 1097
rect 3796 1097 3811 1103
rect 3965 1103 3971 1123
rect 4132 1117 4147 1123
rect 4196 1116 4204 1124
rect 5277 1117 5292 1123
rect 5997 1117 6012 1123
rect 3965 1097 4003 1103
rect 3748 1077 3763 1083
rect 1460 1056 1468 1064
rect 2356 1057 2371 1063
rect 2381 1057 2412 1063
rect 3284 1057 3363 1063
rect 3757 1057 3763 1077
rect 4029 1077 4083 1083
rect 4365 1083 4371 1103
rect 4381 1083 4387 1108
rect 4492 1103 4500 1108
rect 4492 1097 4515 1103
rect 4573 1097 4588 1103
rect 4749 1097 4771 1103
rect 5172 1097 5187 1103
rect 5380 1097 5411 1103
rect 5517 1097 5555 1103
rect 6109 1097 6124 1103
rect 6445 1097 6483 1103
rect 6493 1097 6508 1103
rect 4365 1077 4403 1083
rect 4781 1077 4812 1083
rect 4836 1077 4867 1083
rect 5140 1077 5155 1083
rect 5373 1077 5388 1083
rect 4317 1057 4344 1063
rect 4660 1057 4675 1063
rect 5012 1057 5027 1063
rect 5037 1057 5052 1063
rect 5069 1057 5084 1063
rect 5124 1057 5139 1063
rect 5373 1057 5379 1077
rect 5540 1077 5571 1083
rect 5597 1077 5635 1083
rect 5732 1077 5763 1083
rect 5837 1077 5859 1083
rect 5853 1064 5859 1077
rect 5964 1077 5980 1083
rect 5964 1076 5972 1077
rect 6212 1077 6227 1083
rect 6253 1077 6284 1083
rect 6452 1077 6467 1083
rect 5892 1057 5916 1063
rect 420 1036 422 1044
rect 532 1036 534 1044
rect 884 1036 886 1044
rect 954 1036 956 1044
rect 1412 1036 1414 1044
rect 1594 1036 1596 1044
rect 1748 1037 1795 1043
rect 2468 1036 2470 1044
rect 2682 1036 2684 1044
rect 2740 1036 2742 1044
rect 2788 1036 2790 1044
rect 2858 1036 2860 1044
rect 3130 1036 3132 1044
rect 3460 1036 3462 1044
rect 3508 1036 3510 1044
rect 3956 1036 3958 1044
rect 4900 1036 4904 1044
rect 5476 1036 5478 1044
rect 5594 1036 5596 1044
rect 6356 1037 6371 1043
rect 3304 1006 3310 1014
rect 3318 1006 3324 1014
rect 3332 1006 3338 1014
rect 3346 1006 3352 1014
rect 157 977 172 983
rect 420 977 435 983
rect 3704 976 3708 984
rect 4714 976 4716 984
rect 1108 957 1123 963
rect 2340 956 2348 964
rect 2621 957 2636 963
rect 2989 957 3011 963
rect 3092 956 3100 964
rect 125 917 147 923
rect 477 923 483 943
rect 685 937 700 943
rect 2308 937 2323 943
rect 2349 937 2364 943
rect 2461 937 2515 943
rect 2820 937 2835 943
rect 2948 936 2956 944
rect 3261 937 3283 943
rect 3581 937 3596 943
rect 477 917 508 923
rect 1140 917 1171 923
rect 1229 917 1267 923
rect 829 897 844 903
rect 1229 897 1235 917
rect 2253 917 2275 923
rect 2957 917 2963 936
rect 3261 917 3267 937
rect 3277 912 3283 937
rect 3613 937 3651 943
rect 3741 937 3756 943
rect 3956 937 3971 943
rect 4205 943 4211 963
rect 4285 943 4291 963
rect 4324 956 4332 964
rect 4173 937 4211 943
rect 4221 937 4259 943
rect 4285 937 4300 943
rect 4253 924 4259 937
rect 4429 943 4435 963
rect 4397 937 4435 943
rect 4924 943 4932 944
rect 4916 937 4932 943
rect 5085 937 5100 943
rect 5133 937 5155 943
rect 3405 917 3420 923
rect 3981 917 3996 923
rect 4381 917 4403 923
rect 4589 917 4611 923
rect 4605 904 4611 917
rect 5020 923 5028 928
rect 5133 924 5139 937
rect 5533 937 5571 943
rect 5597 937 5651 943
rect 6284 943 6292 944
rect 6284 937 6300 943
rect 4964 917 4979 923
rect 4989 917 5028 923
rect 5212 923 5220 928
rect 5181 917 5220 923
rect 5268 917 5315 923
rect 5325 917 5363 923
rect 5469 917 5500 923
rect 6380 917 6419 923
rect 6380 912 6388 917
rect 1588 897 1603 903
rect 1709 897 1724 903
rect 1828 897 1843 903
rect 797 877 828 883
rect 1549 877 1619 883
rect 1613 857 1619 877
rect 1796 877 1859 883
rect 1853 857 1859 877
rect 1997 883 2003 903
rect 2196 897 2211 903
rect 2404 896 2412 904
rect 2701 897 2723 903
rect 2765 897 2780 903
rect 3485 897 3507 903
rect 4740 897 4755 903
rect 4797 897 4812 903
rect 4829 897 4899 903
rect 5748 897 5763 903
rect 6141 897 6156 903
rect 3100 884 3108 888
rect 5804 884 5812 888
rect 1988 877 2003 883
rect 3194 876 3196 884
rect 3501 877 3516 883
rect 3562 876 3564 884
rect 5917 877 5996 883
rect 6388 877 6404 883
rect 298 836 300 844
rect 516 836 518 844
rect 3930 836 3932 844
rect 1768 806 1774 814
rect 1782 806 1788 814
rect 1796 806 1802 814
rect 1810 806 1816 814
rect 4824 806 4830 814
rect 4838 806 4844 814
rect 4852 806 4858 814
rect 4866 806 4872 814
rect 36 776 38 784
rect 164 776 166 784
rect 4612 776 4614 784
rect 6356 776 6358 784
rect 244 737 275 743
rect 612 737 627 743
rect 708 737 723 743
rect 1268 737 1283 743
rect 1428 737 1443 743
rect 1524 737 1555 743
rect 1924 737 1948 743
rect 4900 737 4947 743
rect 5356 737 5379 743
rect 5164 732 5172 736
rect 228 717 243 723
rect 621 717 643 723
rect 1677 717 1692 723
rect 3757 717 3772 723
rect 1764 697 1811 703
rect 1821 697 1859 703
rect 2381 697 2435 703
rect 2660 697 2691 703
rect 717 677 739 683
rect 836 677 851 683
rect 1069 677 1084 683
rect 2260 677 2291 683
rect 2301 677 2339 683
rect 2301 664 2307 677
rect 2493 677 2531 683
rect 2541 677 2556 683
rect 2372 656 2380 664
rect 2525 657 2531 677
rect 2612 677 2627 683
rect 2685 677 2691 697
rect 2909 697 2947 703
rect 3268 697 3395 703
rect 3821 703 3827 723
rect 3933 717 3948 723
rect 4468 717 4483 723
rect 5533 717 5548 723
rect 5709 717 5731 723
rect 6509 717 6524 723
rect 3789 697 3827 703
rect 4852 697 4892 703
rect 5149 697 5164 703
rect 5236 697 5251 703
rect 5293 697 5331 703
rect 5901 697 5923 703
rect 6388 697 6403 703
rect 2824 677 2844 683
rect 2957 677 2995 683
rect 2957 664 2963 677
rect 3080 676 3084 684
rect 3284 677 3379 683
rect 3853 677 3907 683
rect 3988 677 4003 683
rect 4189 677 4211 683
rect 4717 677 4732 683
rect 2733 657 2748 663
rect 4093 657 4108 663
rect 4285 657 4307 663
rect 4452 656 4460 664
rect 5229 657 5235 683
rect 5357 677 5372 683
rect 5412 677 5427 683
rect 5469 677 5491 683
rect 5565 677 5603 683
rect 5837 677 5875 683
rect 5828 657 5843 663
rect 5869 657 5875 677
rect 6196 677 6236 683
rect 772 636 776 644
rect 884 636 888 644
rect 1220 637 1235 643
rect 1364 636 1368 644
rect 1604 637 1619 643
rect 1668 636 1670 644
rect 2148 636 2152 644
rect 2244 636 2246 644
rect 3188 637 3203 643
rect 3796 636 3798 644
rect 4020 636 4022 644
rect 4554 636 4556 644
rect 5082 636 5084 644
rect 5572 636 5574 644
rect 5956 636 5960 644
rect 6093 637 6108 643
rect 6548 636 6550 644
rect 3304 606 3310 614
rect 3318 606 3324 614
rect 3332 606 3338 614
rect 3346 606 3352 614
rect 2052 576 2056 584
rect 3530 576 3532 584
rect 4180 576 4182 584
rect 4616 576 4620 584
rect 5604 577 5619 583
rect 157 537 179 543
rect 372 537 392 543
rect 596 537 611 543
rect 1965 537 1987 543
rect 2253 543 2259 563
rect 3204 557 3219 563
rect 2253 537 2268 543
rect 2308 537 2339 543
rect 2349 537 2371 543
rect 2436 537 2451 543
rect 2468 537 2483 543
rect 2797 537 2812 543
rect 3165 543 3171 556
rect 3133 537 3171 543
rect 3373 537 3420 543
rect 3476 537 3507 543
rect 3556 537 3587 543
rect 3613 537 3628 543
rect 4557 524 4563 543
rect 4669 543 4675 556
rect 4660 537 4675 543
rect 4989 537 5004 543
rect 612 517 643 523
rect 1005 517 1043 523
rect 1005 497 1011 517
rect 2612 517 2627 523
rect 3389 517 3404 523
rect 3805 517 3836 523
rect 3908 517 3923 523
rect 4845 517 4924 523
rect 4989 517 5011 523
rect 5101 523 5107 543
rect 5229 537 5267 543
rect 5277 537 5315 543
rect 5580 543 5588 544
rect 5580 537 5596 543
rect 5748 537 5763 543
rect 5805 537 5820 543
rect 5892 537 5907 543
rect 5933 537 5948 543
rect 6173 537 6188 543
rect 6221 537 6236 543
rect 5101 517 5132 523
rect 5789 517 5836 523
rect 6452 517 6483 523
rect 1357 497 1372 503
rect 2237 497 2268 503
rect 2900 497 2915 503
rect 3924 496 3932 504
rect 5140 496 5148 504
rect 5453 497 5475 503
rect 6013 497 6035 503
rect 6109 497 6124 503
rect 733 477 812 483
rect 1188 477 1219 483
rect 1348 477 1404 483
rect 1700 477 1731 483
rect 1908 476 1912 484
rect 2730 476 2732 484
rect 2781 477 2796 483
rect 5261 477 5276 483
rect 6045 477 6099 483
rect 3732 456 3734 464
rect 2164 436 2168 444
rect 2938 436 2940 444
rect 3674 436 3676 444
rect 3860 436 3862 444
rect 4522 436 4524 444
rect 4740 436 4742 444
rect 4836 436 4838 444
rect 4932 436 4934 444
rect 5844 436 5846 444
rect 6154 436 6156 444
rect 6589 437 6620 443
rect 1768 406 1774 414
rect 1782 406 1788 414
rect 1796 406 1802 414
rect 1810 406 1816 414
rect 4824 406 4830 414
rect 4838 406 4844 414
rect 4852 406 4858 414
rect 4866 406 4872 414
rect 333 343 339 363
rect 269 337 339 343
rect 461 337 515 343
rect 525 337 556 343
rect 717 343 723 363
rect 1066 356 1068 364
rect 676 337 723 343
rect 1348 337 1404 343
rect 1677 337 1708 343
rect 2372 336 2376 344
rect 2858 336 2860 344
rect 3085 337 3100 343
rect 3140 337 3171 343
rect 4228 337 4284 343
rect 5981 337 6012 343
rect 268 324 276 328
rect 460 324 468 328
rect 989 317 1011 323
rect 1357 317 1372 323
rect 2756 317 2771 323
rect 77 303 83 316
rect 61 297 83 303
rect 932 297 947 303
rect 1469 297 1484 303
rect 2557 297 2572 303
rect 2941 303 2947 323
rect 3124 317 3139 323
rect 3316 317 3379 323
rect 3492 317 3507 323
rect 4365 317 4387 323
rect 4605 317 4627 323
rect 2868 297 2915 303
rect 2941 297 2979 303
rect 3668 297 3683 303
rect 4317 297 4332 303
rect 4428 303 4436 308
rect 4428 297 4451 303
rect 4660 297 4675 303
rect 861 277 883 283
rect 1156 277 1171 283
rect 1181 277 1212 283
rect 1485 277 1500 283
rect 1768 277 1820 283
rect 2157 277 2172 283
rect 2269 277 2284 283
rect 2884 277 2899 283
rect 2964 277 2979 283
rect 3812 277 3843 283
rect 4220 277 4236 283
rect 4220 276 4228 277
rect 4733 283 4739 296
rect 5741 303 5747 323
rect 5732 297 5747 303
rect 5757 297 5772 303
rect 5949 297 5987 303
rect 4733 277 4755 283
rect 5668 277 5699 283
rect 788 257 803 263
rect 1108 256 1116 264
rect 1501 257 1507 276
rect 2173 257 2195 263
rect 3176 256 3180 264
rect 4013 257 4035 263
rect 4532 256 4540 264
rect 5693 257 5699 277
rect 5885 277 5923 283
rect 5832 256 5836 264
rect 5917 257 5923 277
rect 90 236 92 244
rect 644 236 648 244
rect 1316 236 1320 244
rect 1940 236 1944 244
rect 3268 236 3272 244
rect 3544 236 3548 244
rect 3796 236 3798 244
rect 3892 237 3907 243
rect 4692 236 4694 244
rect 3304 206 3310 214
rect 3318 206 3324 214
rect 3332 206 3338 214
rect 3346 206 3352 214
rect 152 176 156 184
rect 349 177 364 183
rect 4120 176 4124 184
rect 5002 176 5004 184
rect 6420 176 6424 184
rect 6490 176 6492 184
rect 6564 176 6568 184
rect 29 137 51 143
rect 253 143 259 163
rect 877 157 892 163
rect 1076 156 1084 164
rect 1277 157 1292 163
rect 1981 157 2003 163
rect 2285 157 2300 163
rect 253 137 291 143
rect 712 136 716 144
rect 1149 137 1196 143
rect 1492 137 1507 143
rect 1549 137 1564 143
rect 1597 137 1635 143
rect 2532 137 2547 143
rect 2605 143 2611 156
rect 2605 137 2627 143
rect 3181 137 3203 143
rect 3725 143 3731 163
rect 4829 157 4876 163
rect 3693 137 3731 143
rect 3757 137 3772 143
rect 3853 137 3868 143
rect 4029 137 4067 143
rect 4884 137 4899 143
rect 5060 137 5080 143
rect 877 117 892 123
rect 1053 117 1075 123
rect 788 77 812 83
rect 957 83 963 116
rect 1069 104 1075 117
rect 1412 117 1443 123
rect 1108 97 1123 103
rect 1348 98 1352 106
rect 1437 97 1443 117
rect 1476 117 1523 123
rect 2061 117 2076 123
rect 2573 117 2595 123
rect 3076 117 3091 123
rect 3124 117 3155 123
rect 4925 117 4963 123
rect 1460 96 1468 104
rect 2644 96 2652 104
rect 3293 97 3356 103
rect 4813 97 4892 103
rect 4925 97 4931 117
rect 5924 117 5960 123
rect 957 77 972 83
rect 1780 77 1843 83
rect 2365 77 2380 83
rect 1741 57 1788 63
rect 2196 56 2200 64
rect 2365 57 2371 77
rect 3261 77 3388 83
rect 3428 77 3443 83
rect 6285 77 6316 83
rect 3978 36 3980 44
rect 1768 6 1774 14
rect 1782 6 1788 14
rect 1796 6 1802 14
rect 1810 6 1816 14
rect 4824 6 4830 14
rect 4838 6 4844 14
rect 4852 6 4858 14
rect 4866 6 4872 14
<< m2contact >>
rect 1774 4806 1782 4814
rect 1788 4806 1796 4814
rect 1802 4806 1810 4814
rect 4830 4806 4838 4814
rect 4844 4806 4852 4814
rect 4858 4806 4866 4814
rect 460 4736 468 4744
rect 636 4736 644 4744
rect 892 4736 900 4744
rect 1580 4736 1588 4744
rect 4892 4756 4900 4764
rect 1628 4736 1636 4744
rect 3340 4736 3348 4744
rect 5116 4736 5124 4744
rect 5164 4736 5172 4744
rect 5212 4736 5220 4744
rect 5276 4736 5284 4744
rect 5484 4736 5492 4744
rect 5548 4736 5556 4744
rect 6172 4736 6180 4744
rect 6524 4736 6532 4744
rect 492 4716 500 4724
rect 780 4716 788 4724
rect 812 4716 820 4724
rect 1020 4716 1028 4724
rect 1052 4716 1060 4724
rect 1164 4716 1172 4724
rect 1180 4716 1188 4724
rect 1500 4716 1508 4724
rect 1612 4716 1620 4724
rect 2028 4716 2036 4724
rect 2204 4716 2212 4724
rect 2364 4716 2372 4724
rect 2428 4716 2436 4724
rect 508 4696 516 4704
rect 684 4696 692 4704
rect 828 4696 836 4704
rect 860 4696 868 4704
rect 956 4696 964 4704
rect 972 4696 980 4704
rect 1100 4696 1108 4704
rect 1212 4696 1220 4704
rect 1276 4696 1284 4704
rect 1324 4696 1332 4704
rect 1468 4696 1476 4704
rect 1548 4696 1556 4704
rect 1596 4696 1604 4704
rect 1628 4696 1636 4704
rect 1740 4696 1748 4704
rect 1772 4696 1780 4704
rect 1836 4696 1844 4704
rect 1868 4696 1876 4704
rect 1916 4696 1924 4704
rect 1996 4696 2004 4704
rect 2060 4696 2068 4704
rect 2092 4696 2100 4704
rect 2140 4696 2148 4704
rect 2172 4696 2180 4704
rect 2364 4696 2372 4704
rect 2476 4716 2484 4724
rect 2556 4716 2564 4724
rect 2588 4716 2596 4724
rect 3036 4716 3044 4724
rect 2476 4696 2484 4704
rect 2860 4696 2868 4704
rect 2908 4696 2916 4704
rect 2940 4696 2948 4704
rect 3036 4696 3044 4704
rect 3116 4716 3124 4724
rect 3628 4716 3636 4724
rect 3212 4694 3220 4702
rect 3484 4694 3492 4702
rect 3644 4696 3652 4704
rect 3660 4696 3668 4704
rect 12 4676 20 4684
rect 108 4676 116 4684
rect 380 4676 388 4684
rect 460 4676 468 4684
rect 556 4676 564 4684
rect 668 4676 676 4684
rect 732 4676 740 4684
rect 828 4676 836 4684
rect 124 4656 132 4664
rect 204 4656 212 4664
rect 252 4656 260 4664
rect 396 4656 404 4664
rect 428 4656 436 4664
rect 524 4656 532 4664
rect 540 4656 548 4664
rect 620 4656 628 4664
rect 636 4656 644 4664
rect 700 4656 708 4664
rect 732 4656 740 4664
rect 764 4656 772 4664
rect 1068 4676 1076 4684
rect 1116 4676 1124 4684
rect 1228 4676 1236 4684
rect 1292 4676 1300 4684
rect 1308 4676 1316 4684
rect 1340 4676 1348 4684
rect 1372 4680 1380 4688
rect 1420 4676 1428 4684
rect 1452 4676 1460 4684
rect 1484 4676 1492 4684
rect 908 4656 916 4664
rect 924 4656 932 4664
rect 956 4656 964 4664
rect 972 4656 980 4664
rect 1004 4656 1012 4664
rect 1100 4656 1108 4664
rect 1164 4656 1172 4664
rect 1244 4656 1252 4664
rect 1340 4656 1348 4664
rect 1436 4656 1444 4664
rect 1516 4656 1524 4664
rect 1628 4656 1636 4664
rect 1692 4656 1700 4664
rect 1724 4656 1732 4664
rect 1932 4676 1940 4684
rect 1836 4656 1844 4664
rect 2156 4676 2164 4684
rect 2172 4676 2180 4684
rect 2284 4676 2292 4684
rect 2332 4676 2340 4684
rect 2380 4676 2388 4684
rect 2492 4676 2500 4684
rect 2588 4676 2596 4684
rect 2684 4676 2692 4684
rect 2748 4676 2756 4684
rect 2988 4676 2996 4684
rect 3052 4676 3060 4684
rect 3116 4676 3124 4684
rect 3148 4676 3156 4684
rect 3244 4676 3252 4684
rect 3516 4676 3524 4684
rect 3676 4676 3684 4684
rect 3692 4676 3700 4684
rect 3708 4680 3716 4688
rect 3772 4696 3780 4704
rect 3820 4716 3828 4724
rect 4284 4716 4292 4724
rect 4444 4716 4452 4724
rect 4572 4716 4580 4724
rect 4812 4716 4820 4724
rect 4924 4716 4932 4724
rect 4988 4716 4996 4724
rect 5036 4716 5044 4724
rect 5084 4716 5092 4724
rect 5196 4716 5204 4724
rect 5244 4716 5252 4724
rect 5308 4716 5316 4724
rect 5324 4716 5332 4724
rect 5340 4716 5348 4724
rect 5372 4716 5380 4724
rect 5500 4716 5508 4724
rect 5516 4716 5524 4724
rect 5660 4716 5668 4724
rect 5708 4716 5716 4724
rect 6108 4716 6116 4724
rect 6140 4716 6148 4724
rect 6172 4716 6180 4724
rect 6252 4716 6260 4724
rect 6492 4716 6500 4724
rect 3916 4694 3924 4702
rect 4108 4694 4116 4702
rect 4364 4696 4372 4704
rect 4460 4696 4468 4704
rect 4524 4696 4532 4704
rect 4620 4696 4628 4704
rect 4780 4696 4788 4704
rect 4876 4696 4884 4704
rect 4892 4696 4900 4704
rect 4956 4696 4964 4704
rect 5100 4696 5108 4704
rect 5180 4696 5188 4704
rect 5260 4696 5268 4704
rect 5564 4696 5572 4704
rect 5676 4696 5684 4704
rect 5820 4696 5828 4704
rect 5884 4696 5892 4704
rect 3820 4676 3828 4684
rect 3852 4676 3860 4684
rect 3980 4676 3988 4684
rect 4076 4676 4084 4684
rect 4252 4676 4260 4684
rect 4316 4676 4324 4684
rect 2220 4656 2228 4664
rect 2316 4656 2324 4664
rect 2508 4656 2516 4664
rect 2652 4656 2660 4664
rect 2732 4656 2740 4664
rect 2860 4656 2868 4664
rect 2908 4656 2916 4664
rect 2956 4656 2964 4664
rect 3036 4656 3044 4664
rect 4476 4676 4484 4684
rect 4508 4676 4516 4684
rect 4684 4676 4692 4684
rect 4716 4676 4724 4684
rect 4876 4676 4884 4684
rect 4940 4676 4948 4684
rect 5036 4676 5044 4684
rect 5068 4676 5076 4684
rect 5212 4676 5220 4684
rect 5260 4676 5268 4684
rect 5372 4676 5380 4684
rect 5388 4676 5396 4684
rect 5436 4676 5444 4684
rect 5484 4676 5492 4684
rect 5612 4676 5620 4684
rect 5628 4676 5636 4684
rect 5676 4676 5684 4684
rect 5740 4676 5748 4684
rect 5772 4676 5780 4684
rect 5836 4676 5844 4684
rect 5868 4676 5876 4684
rect 5964 4696 5972 4704
rect 5980 4696 5988 4704
rect 6044 4696 6052 4704
rect 6060 4696 6068 4704
rect 6124 4696 6132 4704
rect 6220 4696 6228 4704
rect 6348 4694 6356 4702
rect 6508 4696 6516 4704
rect 6556 4696 6564 4704
rect 5916 4676 5924 4684
rect 5948 4676 5956 4684
rect 5996 4676 6004 4684
rect 6028 4676 6036 4684
rect 6076 4676 6084 4684
rect 6108 4676 6116 4684
rect 6140 4676 6148 4684
rect 6172 4676 6180 4684
rect 6284 4676 6292 4684
rect 6316 4676 6324 4684
rect 3916 4656 3924 4664
rect 4300 4656 4308 4664
rect 4396 4656 4404 4664
rect 4492 4656 4500 4664
rect 4588 4656 4596 4664
rect 4636 4656 4644 4664
rect 4732 4656 4740 4664
rect 4988 4656 4996 4664
rect 5004 4656 5012 4664
rect 5100 4656 5108 4664
rect 5420 4656 5428 4664
rect 5596 4656 5604 4664
rect 5708 4656 5716 4664
rect 5724 4656 5732 4664
rect 5804 4656 5812 4664
rect 6012 4656 6020 4664
rect 76 4636 84 4644
rect 140 4636 148 4644
rect 172 4636 180 4644
rect 220 4636 228 4644
rect 268 4636 276 4644
rect 348 4636 356 4644
rect 412 4636 420 4644
rect 492 4636 500 4644
rect 588 4636 596 4644
rect 1180 4636 1188 4644
rect 1404 4636 1412 4644
rect 1532 4636 1540 4644
rect 1676 4636 1684 4644
rect 1756 4636 1764 4644
rect 1884 4636 1892 4644
rect 2108 4636 2116 4644
rect 2236 4636 2244 4644
rect 2252 4636 2260 4644
rect 2300 4636 2308 4644
rect 2348 4636 2356 4644
rect 2556 4636 2564 4644
rect 2620 4636 2628 4644
rect 2876 4636 2884 4644
rect 2924 4636 2932 4644
rect 3420 4636 3428 4644
rect 3612 4636 3620 4644
rect 4044 4636 4052 4644
rect 4236 4636 4244 4644
rect 4348 4636 4356 4644
rect 4380 4636 4388 4644
rect 4572 4636 4580 4644
rect 4604 4636 4612 4644
rect 5052 4636 5060 4644
rect 5244 4636 5252 4644
rect 5564 4636 5572 4644
rect 5788 4636 5796 4644
rect 5836 4636 5844 4644
rect 5932 4636 5940 4644
rect 6188 4636 6196 4644
rect 6476 4636 6484 4644
rect 6508 4636 6516 4644
rect 6636 4636 6644 4644
rect 3310 4606 3318 4614
rect 3324 4606 3332 4614
rect 3338 4606 3346 4614
rect 620 4576 628 4584
rect 780 4576 788 4584
rect 1260 4576 1268 4584
rect 1292 4576 1300 4584
rect 1580 4576 1588 4584
rect 1836 4576 1844 4584
rect 2636 4576 2644 4584
rect 2748 4576 2756 4584
rect 2812 4576 2820 4584
rect 3436 4576 3444 4584
rect 3548 4576 3556 4584
rect 3852 4576 3860 4584
rect 4108 4576 4116 4584
rect 4300 4576 4308 4584
rect 4444 4576 4452 4584
rect 4684 4576 4692 4584
rect 4828 4576 4836 4584
rect 4988 4576 4996 4584
rect 5164 4576 5172 4584
rect 5292 4576 5300 4584
rect 5356 4576 5364 4584
rect 5500 4576 5508 4584
rect 5644 4576 5652 4584
rect 5708 4576 5716 4584
rect 5868 4576 5876 4584
rect 5916 4576 5924 4584
rect 6012 4576 6020 4584
rect 444 4556 452 4564
rect 940 4556 948 4564
rect 1052 4556 1060 4564
rect 1068 4556 1076 4564
rect 1084 4556 1092 4564
rect 1244 4556 1252 4564
rect 1340 4556 1348 4564
rect 1372 4556 1380 4564
rect 1404 4556 1412 4564
rect 1500 4556 1508 4564
rect 1516 4556 1524 4564
rect 1564 4556 1572 4564
rect 1772 4556 1780 4564
rect 1820 4556 1828 4564
rect 1852 4556 1860 4564
rect 1900 4556 1908 4564
rect 2108 4556 2116 4564
rect 2140 4556 2148 4564
rect 2156 4556 2164 4564
rect 92 4536 100 4544
rect 124 4536 132 4544
rect 252 4536 260 4544
rect 316 4536 324 4544
rect 428 4536 436 4544
rect 476 4536 484 4544
rect 636 4536 644 4544
rect 652 4536 660 4544
rect 764 4536 772 4544
rect 812 4536 820 4544
rect 972 4532 980 4540
rect 1036 4536 1044 4544
rect 1148 4536 1156 4544
rect 1324 4536 1332 4544
rect 1468 4536 1476 4544
rect 1628 4536 1636 4544
rect 44 4516 52 4524
rect 140 4516 148 4524
rect 220 4516 228 4524
rect 268 4516 276 4524
rect 332 4516 340 4524
rect 380 4516 388 4524
rect 444 4516 452 4524
rect 508 4516 516 4524
rect 572 4516 580 4524
rect 1132 4516 1140 4524
rect 60 4496 68 4504
rect 76 4496 84 4504
rect 172 4496 180 4504
rect 236 4496 244 4504
rect 300 4496 308 4504
rect 364 4496 372 4504
rect 380 4496 388 4504
rect 524 4496 532 4504
rect 588 4496 596 4504
rect 604 4496 612 4504
rect 796 4496 804 4504
rect 1196 4516 1204 4524
rect 1212 4516 1220 4524
rect 1276 4516 1284 4524
rect 1340 4516 1348 4524
rect 1372 4516 1380 4524
rect 1452 4516 1460 4524
rect 1516 4516 1524 4524
rect 1548 4516 1556 4524
rect 1724 4536 1732 4544
rect 1948 4536 1956 4544
rect 2060 4536 2068 4544
rect 2108 4536 2116 4544
rect 2188 4536 2196 4544
rect 2220 4536 2228 4544
rect 2412 4556 2420 4564
rect 2444 4556 2452 4564
rect 2524 4556 2532 4564
rect 2652 4556 2660 4564
rect 2684 4556 2692 4564
rect 2764 4556 2772 4564
rect 2796 4556 2804 4564
rect 2908 4556 2916 4564
rect 2940 4556 2948 4564
rect 3180 4556 3188 4564
rect 3404 4556 3412 4564
rect 3916 4556 3924 4564
rect 4364 4556 4372 4564
rect 4508 4556 4516 4564
rect 4604 4556 4612 4564
rect 5180 4556 5188 4564
rect 5276 4556 5284 4564
rect 5548 4556 5556 4564
rect 5580 4556 5588 4564
rect 5612 4556 5620 4564
rect 5660 4556 5668 4564
rect 5788 4556 5796 4564
rect 2284 4536 2292 4544
rect 2348 4536 2356 4544
rect 2492 4536 2500 4544
rect 1660 4516 1668 4524
rect 1676 4516 1684 4524
rect 1708 4516 1716 4524
rect 1884 4516 1892 4524
rect 1932 4516 1940 4524
rect 1964 4516 1972 4524
rect 1180 4496 1188 4504
rect 1292 4496 1300 4504
rect 1420 4496 1428 4504
rect 1484 4496 1492 4504
rect 1596 4496 1604 4504
rect 1692 4496 1700 4504
rect 1996 4496 2004 4504
rect 2044 4516 2052 4524
rect 2092 4516 2100 4524
rect 2268 4516 2276 4524
rect 2300 4516 2308 4524
rect 2348 4516 2356 4524
rect 2364 4516 2372 4524
rect 2396 4516 2404 4524
rect 2428 4516 2436 4524
rect 2444 4516 2452 4524
rect 2476 4516 2484 4524
rect 2524 4516 2532 4524
rect 2556 4516 2564 4524
rect 2700 4536 2708 4544
rect 2796 4536 2804 4544
rect 2844 4536 2852 4544
rect 3276 4536 3284 4544
rect 3388 4536 3396 4544
rect 3484 4536 3492 4544
rect 3516 4536 3524 4544
rect 3564 4536 3572 4544
rect 3628 4536 3636 4544
rect 3660 4536 3668 4544
rect 3692 4536 3700 4544
rect 3756 4536 3764 4544
rect 4060 4536 4068 4544
rect 4124 4536 4132 4544
rect 4268 4536 4276 4544
rect 4332 4536 4340 4544
rect 4364 4536 4372 4544
rect 4380 4536 4388 4544
rect 4716 4536 4724 4544
rect 4732 4536 4740 4544
rect 4812 4536 4820 4544
rect 4844 4536 4852 4544
rect 5020 4536 5028 4544
rect 2620 4516 2628 4524
rect 2652 4516 2660 4524
rect 2684 4516 2692 4524
rect 2860 4516 2868 4524
rect 2908 4516 2916 4524
rect 2940 4516 2948 4524
rect 3036 4518 3044 4526
rect 3100 4516 3108 4524
rect 3212 4516 3220 4524
rect 3260 4516 3268 4524
rect 3372 4516 3380 4524
rect 3436 4516 3444 4524
rect 3468 4516 3476 4524
rect 3516 4516 3524 4524
rect 3580 4516 3588 4524
rect 3724 4518 3732 4526
rect 3916 4518 3924 4526
rect 2188 4496 2196 4504
rect 2332 4496 2340 4504
rect 2412 4496 2420 4504
rect 2748 4496 2756 4504
rect 2892 4496 2900 4504
rect 3228 4496 3236 4504
rect 3260 4496 3268 4504
rect 3340 4496 3348 4504
rect 3436 4496 3444 4504
rect 3500 4496 3508 4504
rect 3964 4516 3972 4524
rect 4076 4516 4084 4524
rect 4316 4516 4324 4524
rect 4380 4516 4388 4524
rect 4396 4516 4404 4524
rect 4476 4516 4484 4524
rect 4540 4516 4548 4524
rect 4636 4516 4644 4524
rect 4716 4516 4724 4524
rect 4764 4516 4772 4524
rect 4796 4516 4804 4524
rect 4860 4516 4868 4524
rect 3628 4496 3636 4504
rect 4300 4496 4308 4504
rect 4444 4496 4452 4504
rect 4460 4496 4468 4504
rect 4524 4496 4532 4504
rect 4604 4496 4612 4504
rect 4668 4496 4676 4504
rect 4684 4496 4692 4504
rect 4780 4496 4788 4504
rect 4940 4516 4948 4524
rect 4988 4516 4996 4524
rect 5148 4536 5156 4544
rect 5196 4536 5204 4544
rect 5308 4536 5316 4544
rect 5340 4536 5348 4544
rect 5404 4536 5412 4544
rect 5420 4536 5428 4544
rect 5516 4536 5524 4544
rect 5740 4536 5748 4544
rect 5932 4536 5940 4544
rect 5964 4536 5972 4544
rect 6028 4536 6036 4544
rect 6092 4536 6100 4544
rect 6140 4536 6148 4544
rect 6204 4536 6212 4544
rect 5100 4516 5108 4524
rect 5132 4516 5140 4524
rect 5228 4516 5236 4524
rect 4988 4496 4996 4504
rect 5052 4496 5060 4504
rect 5116 4496 5124 4504
rect 5244 4496 5252 4504
rect 5388 4516 5396 4524
rect 5436 4516 5444 4524
rect 5580 4516 5588 4524
rect 5708 4516 5716 4524
rect 5820 4516 5828 4524
rect 5868 4516 5876 4524
rect 6044 4516 6052 4524
rect 6108 4516 6116 4524
rect 6172 4516 6180 4524
rect 6188 4516 6196 4524
rect 6252 4516 6260 4524
rect 6300 4516 6308 4524
rect 6380 4516 6388 4524
rect 6428 4516 6436 4524
rect 6492 4516 6500 4524
rect 6556 4516 6564 4524
rect 5468 4496 5476 4504
rect 5724 4496 5732 4504
rect 5756 4496 5764 4504
rect 5772 4496 5780 4504
rect 5884 4496 5892 4504
rect 5900 4496 5908 4504
rect 6012 4496 6020 4504
rect 6076 4496 6084 4504
rect 6140 4496 6148 4504
rect 6268 4496 6276 4504
rect 6284 4496 6292 4504
rect 6396 4496 6404 4504
rect 6476 4496 6484 4504
rect 6540 4496 6548 4504
rect 28 4476 36 4484
rect 204 4476 212 4484
rect 268 4476 276 4484
rect 556 4476 564 4484
rect 1100 4476 1108 4484
rect 1564 4476 1572 4484
rect 1756 4476 1764 4484
rect 2220 4476 2228 4484
rect 3372 4476 3380 4484
rect 3532 4476 3540 4484
rect 4492 4476 4500 4484
rect 4556 4476 4564 4484
rect 4588 4476 4596 4484
rect 4652 4476 4660 4484
rect 4956 4476 4964 4484
rect 5084 4476 5092 4484
rect 5692 4476 5700 4484
rect 5852 4476 5860 4484
rect 6316 4476 6324 4484
rect 6364 4476 6372 4484
rect 6444 4476 6452 4484
rect 6492 4476 6500 4484
rect 6540 4476 6548 4484
rect 220 4456 228 4464
rect 4540 4456 4548 4464
rect 5292 4456 5300 4464
rect 44 4436 52 4444
rect 140 4436 148 4444
rect 412 4436 420 4444
rect 572 4436 580 4444
rect 716 4436 724 4444
rect 844 4436 852 4444
rect 1452 4436 1460 4444
rect 1916 4436 1924 4444
rect 2044 4436 2052 4444
rect 2268 4436 2276 4444
rect 2588 4436 2596 4444
rect 2860 4436 2868 4444
rect 3164 4436 3172 4444
rect 3196 4436 3204 4444
rect 3420 4436 3428 4444
rect 4044 4436 4052 4444
rect 4236 4436 4244 4444
rect 4940 4436 4948 4444
rect 5100 4436 5108 4444
rect 5260 4436 5268 4444
rect 5324 4436 5332 4444
rect 5804 4436 5812 4444
rect 6044 4436 6052 4444
rect 6300 4436 6308 4444
rect 6380 4436 6388 4444
rect 6428 4436 6436 4444
rect 6492 4436 6500 4444
rect 6588 4436 6596 4444
rect 1774 4406 1782 4414
rect 1788 4406 1796 4414
rect 1802 4406 1810 4414
rect 4830 4406 4838 4414
rect 4844 4406 4852 4414
rect 4858 4406 4866 4414
rect 2956 4376 2964 4384
rect 3548 4376 3556 4384
rect 3788 4376 3796 4384
rect 4476 4376 4484 4384
rect 4540 4376 4548 4384
rect 4700 4376 4708 4384
rect 4956 4376 4964 4384
rect 5036 4376 5044 4384
rect 5532 4376 5540 4384
rect 5836 4376 5844 4384
rect 6092 4376 6100 4384
rect 6396 4376 6404 4384
rect 668 4356 676 4364
rect 812 4356 820 4364
rect 1244 4356 1252 4364
rect 2508 4356 2516 4364
rect 3020 4356 3028 4364
rect 572 4336 580 4344
rect 652 4336 660 4344
rect 1180 4336 1188 4344
rect 1980 4336 1988 4344
rect 2252 4336 2260 4344
rect 3068 4336 3076 4344
rect 3388 4336 3396 4344
rect 4140 4336 4148 4344
rect 4204 4336 4212 4344
rect 4460 4336 4468 4344
rect 4524 4336 4532 4344
rect 5324 4336 5332 4344
rect 5452 4336 5460 4344
rect 5612 4336 5620 4344
rect 6380 4336 6388 4344
rect 6460 4336 6468 4344
rect 6508 4336 6516 4344
rect 44 4316 52 4324
rect 124 4316 132 4324
rect 268 4316 276 4324
rect 316 4316 324 4324
rect 380 4316 388 4324
rect 396 4316 404 4324
rect 684 4316 692 4324
rect 860 4316 868 4324
rect 924 4316 932 4324
rect 956 4316 964 4324
rect 1116 4316 1124 4324
rect 1212 4316 1220 4324
rect 1276 4316 1284 4324
rect 1324 4316 1332 4324
rect 1708 4316 1716 4324
rect 1772 4316 1780 4324
rect 1900 4316 1908 4324
rect 2156 4316 2164 4324
rect 2332 4316 2340 4324
rect 2460 4316 2468 4324
rect 2636 4316 2644 4324
rect 2876 4316 2884 4324
rect 2892 4316 2900 4324
rect 2988 4316 2996 4324
rect 3420 4316 3428 4324
rect 3532 4316 3540 4324
rect 44 4296 52 4304
rect 76 4296 84 4304
rect 172 4296 180 4304
rect 428 4296 436 4304
rect 620 4296 628 4304
rect 668 4296 676 4304
rect 700 4296 708 4304
rect 780 4296 788 4304
rect 908 4296 916 4304
rect 1004 4296 1012 4304
rect 1068 4296 1076 4304
rect 1084 4296 1092 4304
rect 1164 4296 1172 4304
rect 1244 4296 1252 4304
rect 1276 4296 1284 4304
rect 1356 4296 1364 4304
rect 1580 4296 1588 4304
rect 1660 4296 1668 4304
rect 1740 4296 1748 4304
rect 1852 4296 1860 4304
rect 1932 4296 1940 4304
rect 1996 4296 2004 4304
rect 2028 4296 2036 4304
rect 2076 4296 2084 4304
rect 2092 4296 2100 4304
rect 2188 4296 2196 4304
rect 2236 4296 2244 4304
rect 2300 4296 2308 4304
rect 2540 4296 2548 4304
rect 2604 4296 2612 4304
rect 2652 4296 2660 4304
rect 2732 4296 2740 4304
rect 2844 4296 2852 4304
rect 2860 4296 2868 4304
rect 2956 4296 2964 4304
rect 3004 4296 3012 4304
rect 3196 4296 3204 4304
rect 3276 4296 3284 4304
rect 3388 4296 3396 4304
rect 3436 4296 3444 4304
rect 3628 4294 3636 4302
rect 3692 4296 3700 4304
rect 3788 4296 3796 4304
rect 3836 4316 3844 4324
rect 3932 4316 3940 4324
rect 4396 4316 4404 4324
rect 4492 4316 4500 4324
rect 4556 4316 4564 4324
rect 4668 4316 4676 4324
rect 4780 4316 4788 4324
rect 4940 4316 4948 4324
rect 5068 4316 5076 4324
rect 3900 4296 3908 4304
rect 3932 4296 3940 4304
rect 3996 4294 4004 4302
rect 4060 4296 4068 4304
rect 4156 4296 4164 4304
rect 4188 4296 4196 4304
rect 4268 4296 4276 4304
rect 4316 4296 4324 4304
rect 4476 4296 4484 4304
rect 4540 4296 4548 4304
rect 4604 4296 4612 4304
rect 4700 4296 4708 4304
rect 4892 4296 4900 4304
rect 5004 4296 5012 4304
rect 5036 4296 5044 4304
rect 5084 4296 5092 4304
rect 5228 4316 5236 4324
rect 5420 4316 5428 4324
rect 5484 4316 5492 4324
rect 5580 4316 5588 4324
rect 5676 4316 5684 4324
rect 5724 4316 5732 4324
rect 5804 4316 5812 4324
rect 5932 4316 5940 4324
rect 5964 4316 5972 4324
rect 6012 4316 6020 4324
rect 6060 4316 6068 4324
rect 6236 4316 6244 4324
rect 6316 4316 6324 4324
rect 6412 4316 6420 4324
rect 6540 4316 6548 4324
rect 6556 4316 6564 4324
rect 6604 4316 6612 4324
rect 5164 4296 5172 4304
rect 5244 4296 5252 4304
rect 5292 4296 5300 4304
rect 5324 4296 5332 4304
rect 5340 4296 5348 4304
rect 5388 4296 5396 4304
rect 5468 4296 5476 4304
rect 5532 4296 5540 4304
rect 5756 4296 5764 4304
rect 5788 4296 5796 4304
rect 6188 4296 6196 4304
rect 6300 4296 6308 4304
rect 6396 4296 6404 4304
rect 6444 4296 6452 4304
rect 6476 4296 6484 4304
rect 6524 4296 6532 4304
rect 92 4276 100 4284
rect 140 4276 148 4284
rect 300 4276 308 4284
rect 348 4276 356 4284
rect 12 4256 20 4264
rect 108 4256 116 4264
rect 204 4256 212 4264
rect 252 4256 260 4264
rect 444 4276 452 4284
rect 460 4276 468 4284
rect 556 4276 564 4284
rect 604 4276 612 4284
rect 716 4276 724 4284
rect 764 4276 772 4284
rect 828 4276 836 4284
rect 988 4276 996 4284
rect 1068 4276 1076 4284
rect 1180 4276 1188 4284
rect 1228 4276 1236 4284
rect 1340 4276 1348 4284
rect 1372 4276 1380 4284
rect 1388 4276 1396 4284
rect 1484 4276 1492 4284
rect 1596 4276 1604 4284
rect 1692 4276 1700 4284
rect 1756 4276 1764 4284
rect 1948 4276 1956 4284
rect 2108 4276 2116 4284
rect 2268 4276 2276 4284
rect 2348 4276 2356 4284
rect 2444 4276 2452 4284
rect 2492 4276 2500 4284
rect 2588 4276 2596 4284
rect 572 4256 580 4264
rect 748 4256 756 4264
rect 876 4256 884 4264
rect 908 4256 916 4264
rect 940 4256 948 4264
rect 1020 4256 1028 4264
rect 1036 4256 1044 4264
rect 1132 4256 1140 4264
rect 1164 4256 1172 4264
rect 1308 4256 1316 4264
rect 1516 4256 1524 4264
rect 1836 4256 1844 4264
rect 1964 4256 1972 4264
rect 2028 4256 2036 4264
rect 2076 4256 2084 4264
rect 2140 4256 2148 4264
rect 2188 4256 2196 4264
rect 2220 4256 2228 4264
rect 2524 4256 2532 4264
rect 2540 4256 2548 4264
rect 2572 4256 2580 4264
rect 2652 4256 2660 4264
rect 2684 4256 2692 4264
rect 2780 4276 2788 4284
rect 2940 4276 2948 4284
rect 3052 4276 3060 4284
rect 3100 4276 3108 4284
rect 3132 4276 3140 4284
rect 3164 4276 3172 4284
rect 3292 4276 3300 4284
rect 3372 4276 3380 4284
rect 3452 4276 3460 4284
rect 3500 4276 3508 4284
rect 3772 4276 3780 4284
rect 3868 4276 3876 4284
rect 3884 4276 3892 4284
rect 3964 4276 3972 4284
rect 4140 4276 4148 4284
rect 4220 4276 4228 4284
rect 4364 4276 4372 4284
rect 4428 4276 4436 4284
rect 4572 4276 4580 4284
rect 4620 4276 4628 4284
rect 4652 4276 4660 4284
rect 4716 4276 4724 4284
rect 4796 4276 4804 4284
rect 4876 4276 4884 4284
rect 5180 4276 5188 4284
rect 5196 4276 5204 4284
rect 5468 4276 5476 4284
rect 5548 4276 5556 4284
rect 5596 4276 5604 4284
rect 5644 4276 5652 4284
rect 5676 4276 5684 4284
rect 5740 4276 5748 4284
rect 5868 4276 5876 4284
rect 5932 4276 5940 4284
rect 5980 4276 5988 4284
rect 6012 4276 6020 4284
rect 6172 4276 6180 4284
rect 6204 4276 6212 4284
rect 6316 4276 6324 4284
rect 6348 4276 6356 4284
rect 6588 4276 6596 4284
rect 6636 4276 6644 4284
rect 2796 4256 2804 4264
rect 3036 4256 3044 4264
rect 3132 4256 3140 4264
rect 3276 4256 3284 4264
rect 3484 4256 3492 4264
rect 3564 4256 3572 4264
rect 4652 4256 4660 4264
rect 4796 4256 4804 4264
rect 4860 4256 4868 4264
rect 4940 4256 4948 4264
rect 4972 4256 4980 4264
rect 5004 4256 5012 4264
rect 5116 4256 5124 4264
rect 5132 4256 5140 4264
rect 5228 4256 5236 4264
rect 5276 4256 5284 4264
rect 5388 4256 5396 4264
rect 5404 4256 5412 4264
rect 5500 4256 5508 4264
rect 5628 4256 5636 4264
rect 5676 4256 5684 4264
rect 5804 4256 5812 4264
rect 5916 4256 5924 4264
rect 6076 4256 6084 4264
rect 6108 4256 6116 4264
rect 6252 4256 6260 4264
rect 6524 4256 6532 4264
rect 44 4236 52 4244
rect 236 4236 244 4244
rect 284 4236 292 4244
rect 316 4236 324 4244
rect 396 4236 404 4244
rect 492 4236 500 4244
rect 732 4236 740 4244
rect 860 4236 868 4244
rect 956 4236 964 4244
rect 1116 4236 1124 4244
rect 1212 4236 1220 4244
rect 1420 4236 1428 4244
rect 1500 4236 1508 4244
rect 1548 4236 1556 4244
rect 1628 4236 1636 4244
rect 1868 4236 1876 4244
rect 2124 4236 2132 4244
rect 2204 4236 2212 4244
rect 2332 4236 2340 4244
rect 2396 4236 2404 4244
rect 2460 4236 2468 4244
rect 2764 4236 2772 4244
rect 2908 4236 2916 4244
rect 3148 4236 3156 4244
rect 3244 4236 3252 4244
rect 3468 4236 3476 4244
rect 3532 4236 3540 4244
rect 3756 4236 3764 4244
rect 4124 4236 4132 4244
rect 4412 4236 4420 4244
rect 4924 4236 4932 4244
rect 5964 4236 5972 4244
rect 6012 4236 6020 4244
rect 6060 4236 6068 4244
rect 6156 4236 6164 4244
rect 6220 4236 6228 4244
rect 6268 4236 6276 4244
rect 6332 4236 6340 4244
rect 6556 4236 6564 4244
rect 6604 4236 6612 4244
rect 3310 4206 3318 4214
rect 3324 4206 3332 4214
rect 3338 4206 3346 4214
rect 12 4176 20 4184
rect 1100 4176 1108 4184
rect 1884 4176 1892 4184
rect 2796 4176 2804 4184
rect 3036 4176 3044 4184
rect 3228 4176 3236 4184
rect 3548 4176 3556 4184
rect 3564 4176 3572 4184
rect 3596 4176 3604 4184
rect 3804 4176 3812 4184
rect 3900 4176 3908 4184
rect 4092 4176 4100 4184
rect 4492 4176 4500 4184
rect 4508 4176 4516 4184
rect 4828 4176 4836 4184
rect 5068 4176 5076 4184
rect 5372 4176 5380 4184
rect 5660 4176 5668 4184
rect 5740 4176 5748 4184
rect 6284 4176 6292 4184
rect 6428 4176 6436 4184
rect 316 4156 324 4164
rect 428 4156 436 4164
rect 556 4156 564 4164
rect 652 4156 660 4164
rect 780 4156 788 4164
rect 876 4156 884 4164
rect 1164 4156 1172 4164
rect 1356 4156 1364 4164
rect 1900 4156 1908 4164
rect 2076 4156 2084 4164
rect 2204 4156 2212 4164
rect 2476 4156 2484 4164
rect 2508 4156 2516 4164
rect 2860 4156 2868 4164
rect 2876 4156 2884 4164
rect 3020 4156 3028 4164
rect 3244 4156 3252 4164
rect 3580 4156 3588 4164
rect 3644 4156 3652 4164
rect 3724 4156 3732 4164
rect 4140 4156 4148 4164
rect 4364 4156 4372 4164
rect 4620 4156 4628 4164
rect 4812 4156 4820 4164
rect 4844 4156 4852 4164
rect 5116 4156 5124 4164
rect 5692 4156 5700 4164
rect 5868 4156 5876 4164
rect 5932 4156 5940 4164
rect 6060 4156 6068 4164
rect 6156 4156 6164 4164
rect 6364 4156 6372 4164
rect 6444 4156 6452 4164
rect 6556 4156 6564 4164
rect 124 4136 132 4144
rect 204 4136 212 4144
rect 300 4136 308 4144
rect 348 4136 356 4144
rect 540 4136 548 4144
rect 668 4136 676 4144
rect 764 4136 772 4144
rect 812 4136 820 4144
rect 908 4136 916 4144
rect 988 4136 996 4144
rect 1148 4136 1156 4144
rect 1164 4136 1172 4144
rect 1244 4136 1252 4144
rect 1276 4136 1284 4144
rect 1324 4136 1332 4144
rect 1612 4136 1620 4144
rect 1676 4136 1684 4144
rect 1756 4136 1764 4144
rect 1868 4136 1876 4144
rect 1916 4136 1924 4144
rect 2012 4136 2020 4144
rect 2028 4136 2036 4144
rect 2060 4136 2068 4144
rect 2124 4136 2132 4144
rect 2156 4136 2164 4144
rect 2220 4136 2228 4144
rect 2284 4136 2292 4144
rect 2348 4136 2356 4144
rect 2364 4136 2372 4144
rect 108 4116 116 4124
rect 396 4116 404 4124
rect 572 4116 580 4124
rect 604 4116 612 4124
rect 620 4116 628 4124
rect 844 4116 852 4124
rect 860 4116 868 4124
rect 860 4096 868 4104
rect 1004 4116 1012 4124
rect 1212 4116 1220 4124
rect 1436 4116 1444 4124
rect 1484 4116 1492 4124
rect 1580 4116 1588 4124
rect 1596 4116 1604 4124
rect 1660 4116 1668 4124
rect 1836 4116 1844 4124
rect 1852 4116 1860 4124
rect 2076 4116 2084 4124
rect 2108 4116 2116 4124
rect 2140 4116 2148 4124
rect 2236 4116 2244 4124
rect 2268 4116 2276 4124
rect 2300 4116 2308 4124
rect 2332 4116 2340 4124
rect 2588 4136 2596 4144
rect 2636 4136 2644 4144
rect 2700 4136 2708 4144
rect 2716 4136 2724 4144
rect 2780 4136 2788 4144
rect 2828 4136 2836 4144
rect 2924 4136 2932 4144
rect 2988 4136 2996 4144
rect 3196 4136 3204 4144
rect 3260 4136 3268 4144
rect 3436 4136 3444 4144
rect 3740 4136 3748 4144
rect 3772 4136 3780 4144
rect 3852 4136 3860 4144
rect 3868 4136 3876 4144
rect 3916 4136 3924 4144
rect 3980 4136 3988 4144
rect 4076 4136 4084 4144
rect 4124 4136 4132 4144
rect 4156 4136 4164 4144
rect 4204 4136 4212 4144
rect 4268 4136 4276 4144
rect 4300 4136 4308 4144
rect 4556 4136 4564 4144
rect 4604 4136 4612 4144
rect 4668 4136 4676 4144
rect 4732 4136 4740 4144
rect 4748 4136 4756 4144
rect 5100 4136 5108 4144
rect 5164 4136 5172 4144
rect 5228 4136 5236 4144
rect 5260 4136 5268 4144
rect 5340 4136 5348 4144
rect 5372 4136 5380 4144
rect 5436 4136 5444 4144
rect 5500 4136 5508 4144
rect 5516 4136 5524 4144
rect 5580 4136 5588 4144
rect 5644 4136 5652 4144
rect 5708 4136 5716 4144
rect 5756 4136 5764 4144
rect 5852 4136 5860 4144
rect 5900 4136 5908 4144
rect 6012 4136 6020 4144
rect 6108 4136 6116 4144
rect 6124 4136 6132 4144
rect 6236 4136 6244 4144
rect 6412 4136 6420 4144
rect 6444 4136 6452 4144
rect 2428 4116 2436 4124
rect 2620 4116 2628 4124
rect 2652 4116 2660 4124
rect 2684 4116 2692 4124
rect 2748 4116 2756 4124
rect 2828 4116 2836 4124
rect 2876 4116 2884 4124
rect 2908 4116 2916 4124
rect 2940 4116 2948 4124
rect 2956 4116 2964 4124
rect 3148 4116 3156 4124
rect 3356 4116 3364 4124
rect 3420 4118 3428 4126
rect 3676 4116 3684 4124
rect 3692 4116 3700 4124
rect 3756 4116 3764 4124
rect 3836 4116 3844 4124
rect 3932 4116 3940 4124
rect 4364 4118 4372 4126
rect 1116 4096 1124 4104
rect 1180 4096 1188 4104
rect 1244 4096 1252 4104
rect 1260 4096 1268 4104
rect 1564 4096 1572 4104
rect 1724 4096 1732 4104
rect 1820 4096 1828 4104
rect 2060 4096 2068 4104
rect 2268 4096 2276 4104
rect 2364 4096 2372 4104
rect 2412 4096 2420 4104
rect 2716 4096 2724 4104
rect 2780 4096 2788 4104
rect 3308 4096 3316 4104
rect 3596 4096 3604 4104
rect 3788 4096 3796 4104
rect 3804 4096 3812 4104
rect 3900 4096 3908 4104
rect 3964 4096 3972 4104
rect 4044 4096 4052 4104
rect 4092 4096 4100 4104
rect 4540 4116 4548 4124
rect 4620 4116 4628 4124
rect 4652 4116 4660 4124
rect 4700 4116 4708 4124
rect 4716 4116 4724 4124
rect 4764 4116 4772 4124
rect 4812 4116 4820 4124
rect 4972 4116 4980 4124
rect 5036 4116 5044 4124
rect 5148 4116 5156 4124
rect 4268 4096 4276 4104
rect 4556 4096 4564 4104
rect 4620 4096 4628 4104
rect 4684 4096 4692 4104
rect 4796 4096 4804 4104
rect 4988 4096 4996 4104
rect 5052 4096 5060 4104
rect 5068 4096 5076 4104
rect 5196 4096 5204 4104
rect 5244 4116 5252 4124
rect 5292 4116 5300 4124
rect 5324 4116 5332 4124
rect 5516 4116 5524 4124
rect 5532 4116 5540 4124
rect 5596 4116 5604 4124
rect 5644 4116 5652 4124
rect 5804 4116 5812 4124
rect 5980 4116 5988 4124
rect 6012 4116 6020 4124
rect 6044 4116 6052 4124
rect 6108 4116 6116 4124
rect 6188 4116 6196 4124
rect 6252 4116 6260 4124
rect 6316 4116 6324 4124
rect 6396 4116 6404 4124
rect 6476 4116 6484 4124
rect 6524 4116 6532 4124
rect 6588 4116 6596 4124
rect 5276 4096 5284 4104
rect 5372 4096 5380 4104
rect 5420 4096 5428 4104
rect 5468 4096 5476 4104
rect 5564 4096 5572 4104
rect 5628 4096 5636 4104
rect 5676 4096 5684 4104
rect 5932 4096 5940 4104
rect 5996 4096 6004 4104
rect 6172 4096 6180 4104
rect 6284 4096 6292 4104
rect 6300 4096 6308 4104
rect 6508 4096 6516 4104
rect 1276 4076 1284 4084
rect 1356 4076 1364 4084
rect 2444 4076 2452 4084
rect 4924 4076 4932 4084
rect 4956 4076 4964 4084
rect 5020 4076 5028 4084
rect 5036 4076 5044 4084
rect 5308 4076 5316 4084
rect 5404 4076 5412 4084
rect 5964 4076 5972 4084
rect 6204 4076 6212 4084
rect 6220 4076 6228 4084
rect 6316 4076 6324 4084
rect 6332 4076 6340 4084
rect 4972 4056 4980 4064
rect 5980 4056 5988 4064
rect 12 4036 20 4044
rect 236 4036 244 4044
rect 476 4036 484 4044
rect 716 4036 724 4044
rect 1100 4036 1108 4044
rect 1628 4036 1636 4044
rect 1692 4036 1700 4044
rect 1948 4036 1956 4044
rect 2300 4036 2308 4044
rect 2428 4036 2436 4044
rect 2556 4036 2564 4044
rect 2668 4036 2676 4044
rect 2892 4036 2900 4044
rect 3692 4036 3700 4044
rect 3996 4036 4004 4044
rect 4188 4036 4196 4044
rect 5036 4036 5044 4044
rect 5132 4036 5140 4044
rect 5452 4036 5460 4044
rect 5532 4036 5540 4044
rect 5884 4036 5892 4044
rect 6156 4036 6164 4044
rect 6316 4036 6324 4044
rect 6444 4036 6452 4044
rect 6476 4036 6484 4044
rect 6620 4036 6628 4044
rect 1774 4006 1782 4014
rect 1788 4006 1796 4014
rect 1802 4006 1810 4014
rect 4830 4006 4838 4014
rect 4844 4006 4852 4014
rect 4858 4006 4866 4014
rect 636 3976 644 3984
rect 2092 3976 2100 3984
rect 2444 3976 2452 3984
rect 3660 3976 3668 3984
rect 4764 3976 4772 3984
rect 5244 3976 5252 3984
rect 5340 3976 5348 3984
rect 5612 3976 5620 3984
rect 6492 3976 6500 3984
rect 5068 3956 5076 3964
rect 6156 3956 6164 3964
rect 28 3936 36 3944
rect 508 3936 516 3944
rect 524 3936 532 3944
rect 1916 3936 1924 3944
rect 4108 3936 4116 3944
rect 5820 3936 5828 3944
rect 5980 3936 5988 3944
rect 5996 3936 6004 3944
rect 6140 3936 6148 3944
rect 140 3916 148 3924
rect 156 3916 164 3924
rect 204 3916 212 3924
rect 540 3916 548 3924
rect 876 3916 884 3924
rect 1132 3916 1140 3924
rect 1196 3916 1204 3924
rect 1260 3916 1268 3924
rect 1468 3916 1476 3924
rect 12 3896 20 3904
rect 92 3896 100 3904
rect 236 3896 244 3904
rect 268 3896 276 3904
rect 300 3896 308 3904
rect 364 3894 372 3902
rect 588 3896 596 3904
rect 700 3896 708 3904
rect 764 3894 772 3902
rect 828 3896 836 3904
rect 876 3896 884 3904
rect 940 3894 948 3902
rect 988 3896 996 3904
rect 1100 3896 1108 3904
rect 1132 3896 1140 3904
rect 1180 3896 1188 3904
rect 1404 3894 1412 3902
rect 1532 3896 1540 3904
rect 1548 3896 1556 3904
rect 1580 3896 1588 3904
rect 1628 3896 1636 3904
rect 1660 3896 1668 3904
rect 1804 3896 1812 3904
rect 1852 3896 1860 3904
rect 1948 3896 1956 3904
rect 1964 3896 1972 3904
rect 1996 3916 2004 3924
rect 2396 3916 2404 3924
rect 2428 3916 2436 3924
rect 3036 3916 3044 3924
rect 3308 3916 3316 3924
rect 3676 3916 3684 3924
rect 3740 3916 3748 3924
rect 3804 3916 3812 3924
rect 3884 3916 3892 3924
rect 4236 3916 4244 3924
rect 4364 3916 4372 3924
rect 4444 3916 4452 3924
rect 4604 3916 4612 3924
rect 2316 3894 2324 3902
rect 2396 3896 2404 3904
rect 2476 3896 2484 3904
rect 2540 3896 2548 3904
rect 2668 3896 2676 3904
rect 2940 3896 2948 3904
rect 3036 3896 3044 3904
rect 3116 3896 3124 3904
rect 3148 3896 3156 3904
rect 3260 3896 3268 3904
rect 3340 3896 3348 3904
rect 3404 3894 3412 3902
rect 3772 3896 3780 3904
rect 3788 3896 3796 3904
rect 3820 3896 3828 3904
rect 3980 3894 3988 3902
rect 4284 3896 4292 3904
rect 4364 3896 4372 3904
rect 4492 3896 4500 3904
rect 172 3876 180 3884
rect 188 3876 196 3884
rect 204 3876 212 3884
rect 252 3876 260 3884
rect 332 3876 340 3884
rect 412 3876 420 3884
rect 572 3876 580 3884
rect 620 3876 628 3884
rect 828 3876 836 3884
rect 908 3876 916 3884
rect 1084 3876 1092 3884
rect 1116 3876 1124 3884
rect 1436 3876 1444 3884
rect 1484 3876 1492 3884
rect 1516 3876 1524 3884
rect 1532 3876 1540 3884
rect 1596 3876 1604 3884
rect 1612 3876 1620 3884
rect 1676 3876 1684 3884
rect 1932 3876 1940 3884
rect 2028 3876 2036 3884
rect 2108 3876 2116 3884
rect 2348 3876 2356 3884
rect 2380 3876 2388 3884
rect 2492 3876 2500 3884
rect 2540 3876 2548 3884
rect 2620 3876 2628 3884
rect 2716 3876 2724 3884
rect 2892 3876 2900 3884
rect 2908 3876 2916 3884
rect 2988 3876 2996 3884
rect 3244 3876 3252 3884
rect 3436 3876 3444 3884
rect 3548 3876 3556 3884
rect 3564 3876 3572 3884
rect 3612 3880 3620 3888
rect 3628 3876 3636 3884
rect 3644 3876 3652 3884
rect 3692 3876 3700 3884
rect 3884 3876 3892 3884
rect 3900 3876 3908 3884
rect 3916 3876 3924 3884
rect 3948 3876 3956 3884
rect 4124 3876 4132 3884
rect 4220 3876 4228 3884
rect 4252 3876 4260 3884
rect 4268 3876 4276 3884
rect 4300 3876 4308 3884
rect 4348 3876 4356 3884
rect 4396 3876 4404 3884
rect 4460 3876 4468 3884
rect 4572 3896 4580 3904
rect 4668 3916 4676 3924
rect 4796 3916 4804 3924
rect 4940 3916 4948 3924
rect 5180 3916 5188 3924
rect 5196 3916 5204 3924
rect 5308 3916 5316 3924
rect 5452 3916 5460 3924
rect 5516 3916 5524 3924
rect 5580 3916 5588 3924
rect 5596 3916 5604 3924
rect 5692 3916 5700 3924
rect 5740 3916 5748 3924
rect 5852 3916 5860 3924
rect 4700 3896 4708 3904
rect 4764 3896 4772 3904
rect 4908 3896 4916 3904
rect 4924 3896 4932 3904
rect 4956 3896 4964 3904
rect 5052 3896 5060 3904
rect 5100 3896 5108 3904
rect 5164 3896 5172 3904
rect 5212 3896 5220 3904
rect 5260 3896 5268 3904
rect 5292 3896 5300 3904
rect 5340 3896 5348 3904
rect 5420 3896 5428 3904
rect 5532 3896 5540 3904
rect 5548 3896 5556 3904
rect 5596 3896 5604 3904
rect 5660 3896 5668 3904
rect 5948 3916 5956 3924
rect 6060 3916 6068 3924
rect 6444 3916 6452 3924
rect 5964 3896 5972 3904
rect 6028 3896 6036 3904
rect 6108 3896 6116 3904
rect 6156 3896 6164 3904
rect 6268 3896 6276 3904
rect 6284 3896 6292 3904
rect 6348 3896 6356 3904
rect 6540 3896 6548 3904
rect 4572 3876 4580 3884
rect 4652 3876 4660 3884
rect 4700 3876 4708 3884
rect 4748 3876 4756 3884
rect 4812 3876 4820 3884
rect 4892 3876 4900 3884
rect 5004 3876 5012 3884
rect 5148 3876 5156 3884
rect 5452 3876 5460 3884
rect 5468 3876 5476 3884
rect 5532 3876 5540 3884
rect 5628 3876 5636 3884
rect 5644 3876 5652 3884
rect 5708 3876 5716 3884
rect 5772 3876 5780 3884
rect 5820 3876 5828 3884
rect 6012 3876 6020 3884
rect 6252 3876 6260 3884
rect 6300 3876 6308 3884
rect 6332 3876 6340 3884
rect 6476 3876 6484 3884
rect 6524 3876 6532 3884
rect 6540 3876 6548 3884
rect 6620 3896 6628 3904
rect 6572 3876 6580 3884
rect 6604 3876 6612 3884
rect 44 3856 52 3864
rect 300 3856 308 3864
rect 508 3856 516 3864
rect 1148 3856 1156 3864
rect 1260 3856 1268 3864
rect 1580 3856 1588 3864
rect 2044 3856 2052 3864
rect 2316 3856 2324 3864
rect 2460 3856 2468 3864
rect 2956 3856 2964 3864
rect 4716 3856 4724 3864
rect 4988 3856 4996 3864
rect 5084 3856 5092 3864
rect 5132 3856 5140 3864
rect 5260 3856 5268 3864
rect 5372 3856 5380 3864
rect 5740 3856 5748 3864
rect 5756 3856 5764 3864
rect 5884 3856 5892 3864
rect 5932 3856 5940 3864
rect 6076 3856 6084 3864
rect 6188 3856 6196 3864
rect 6364 3856 6372 3864
rect 6428 3856 6436 3864
rect 6492 3856 6500 3864
rect 140 3836 148 3844
rect 556 3836 564 3844
rect 1068 3836 1076 3844
rect 1212 3836 1220 3844
rect 1276 3836 1284 3844
rect 1660 3836 1668 3844
rect 2156 3836 2164 3844
rect 2188 3836 2196 3844
rect 2444 3836 2452 3844
rect 2508 3836 2516 3844
rect 2556 3836 2564 3844
rect 2764 3836 2772 3844
rect 3052 3836 3060 3844
rect 3532 3836 3540 3844
rect 3580 3836 3588 3844
rect 4156 3836 4164 3844
rect 4332 3836 4340 3844
rect 4380 3836 4388 3844
rect 4524 3836 4532 3844
rect 4620 3836 4628 3844
rect 4972 3836 4980 3844
rect 5116 3836 5124 3844
rect 6060 3836 6068 3844
rect 6092 3836 6100 3844
rect 6236 3836 6244 3844
rect 6316 3836 6324 3844
rect 6380 3836 6388 3844
rect 6412 3836 6420 3844
rect 6444 3836 6452 3844
rect 6508 3836 6516 3844
rect 6572 3836 6580 3844
rect 3310 3806 3318 3814
rect 3324 3806 3332 3814
rect 3338 3806 3346 3814
rect 12 3776 20 3784
rect 316 3776 324 3784
rect 764 3776 772 3784
rect 956 3776 964 3784
rect 1660 3776 1668 3784
rect 1676 3776 1684 3784
rect 2204 3776 2212 3784
rect 3260 3776 3268 3784
rect 3372 3776 3380 3784
rect 3420 3776 3428 3784
rect 3484 3776 3492 3784
rect 3644 3776 3652 3784
rect 3916 3776 3924 3784
rect 4108 3776 4116 3784
rect 4748 3776 4756 3784
rect 4780 3776 4788 3784
rect 5004 3776 5012 3784
rect 5068 3776 5076 3784
rect 5212 3776 5220 3784
rect 5996 3776 6004 3784
rect 6540 3776 6548 3784
rect 620 3756 628 3764
rect 892 3756 900 3764
rect 1692 3756 1700 3764
rect 1708 3756 1716 3764
rect 2076 3756 2084 3764
rect 2188 3756 2196 3764
rect 2716 3756 2724 3764
rect 2860 3756 2868 3764
rect 2988 3756 2996 3764
rect 3276 3756 3284 3764
rect 3356 3756 3364 3764
rect 3388 3756 3396 3764
rect 3404 3756 3412 3764
rect 124 3736 132 3744
rect 204 3736 212 3744
rect 268 3736 276 3744
rect 300 3736 308 3744
rect 412 3736 420 3744
rect 508 3736 516 3744
rect 604 3736 612 3744
rect 652 3736 660 3744
rect 748 3736 756 3744
rect 1004 3736 1012 3744
rect 1052 3736 1060 3744
rect 1148 3736 1156 3744
rect 1164 3736 1172 3744
rect 1260 3736 1268 3744
rect 1324 3736 1332 3744
rect 1340 3736 1348 3744
rect 1404 3736 1412 3744
rect 1468 3736 1476 3744
rect 1740 3736 1748 3744
rect 1996 3736 2004 3744
rect 2060 3736 2068 3744
rect 2172 3736 2180 3744
rect 2316 3736 2324 3744
rect 2396 3736 2404 3744
rect 2460 3736 2468 3744
rect 2556 3736 2564 3744
rect 2652 3736 2660 3744
rect 2876 3736 2884 3744
rect 2940 3736 2948 3744
rect 3020 3736 3028 3744
rect 3100 3736 3108 3744
rect 3436 3736 3444 3744
rect 3660 3756 3668 3764
rect 3676 3756 3684 3764
rect 4668 3756 4676 3764
rect 4684 3756 4692 3764
rect 4764 3756 4772 3764
rect 4924 3756 4932 3764
rect 5580 3756 5588 3764
rect 5964 3756 5972 3764
rect 6380 3756 6388 3764
rect 6412 3756 6420 3764
rect 3564 3736 3572 3744
rect 3628 3736 3636 3744
rect 3724 3736 3732 3744
rect 3788 3736 3796 3744
rect 3948 3736 3956 3744
rect 4220 3736 4228 3744
rect 4268 3736 4276 3744
rect 4284 3736 4292 3744
rect 4316 3736 4324 3744
rect 4332 3736 4340 3744
rect 4396 3736 4404 3744
rect 4460 3736 4468 3744
rect 4540 3736 4548 3744
rect 4700 3736 4708 3744
rect 4860 3736 4868 3744
rect 4924 3736 4932 3744
rect 140 3718 148 3726
rect 220 3716 228 3724
rect 428 3716 436 3724
rect 524 3716 532 3724
rect 268 3696 276 3704
rect 572 3696 580 3704
rect 684 3696 692 3704
rect 716 3716 724 3724
rect 732 3716 740 3724
rect 876 3716 884 3724
rect 956 3696 964 3704
rect 1036 3696 1044 3704
rect 1084 3696 1092 3704
rect 1308 3716 1316 3724
rect 1356 3716 1364 3724
rect 1388 3716 1396 3724
rect 1420 3716 1428 3724
rect 1452 3716 1460 3724
rect 1564 3716 1572 3724
rect 1596 3716 1604 3724
rect 1964 3718 1972 3726
rect 2124 3716 2132 3724
rect 2332 3718 2340 3726
rect 2412 3716 2420 3724
rect 2428 3716 2436 3724
rect 2508 3716 2516 3724
rect 1276 3696 1284 3704
rect 1628 3696 1636 3704
rect 1740 3696 1748 3704
rect 1772 3696 1780 3704
rect 2028 3696 2036 3704
rect 2108 3696 2116 3704
rect 2492 3696 2500 3704
rect 2588 3696 2596 3704
rect 2636 3716 2644 3724
rect 2732 3716 2740 3724
rect 2764 3716 2772 3724
rect 2892 3716 2900 3724
rect 2924 3716 2932 3724
rect 2956 3716 2964 3724
rect 3036 3716 3044 3724
rect 3052 3716 3060 3724
rect 3132 3718 3140 3726
rect 3340 3716 3348 3724
rect 3452 3716 3460 3724
rect 3500 3716 3508 3724
rect 3548 3716 3556 3724
rect 3596 3716 3604 3724
rect 3612 3716 3620 3724
rect 3708 3716 3716 3724
rect 3804 3716 3812 3724
rect 3996 3716 4004 3724
rect 4140 3716 4148 3724
rect 4348 3716 4356 3724
rect 4412 3716 4420 3724
rect 4444 3716 4452 3724
rect 4508 3716 4516 3724
rect 4556 3716 4564 3724
rect 4636 3716 4644 3724
rect 4716 3716 4724 3724
rect 4796 3716 4804 3724
rect 4940 3716 4948 3724
rect 4972 3736 4980 3744
rect 5020 3736 5028 3744
rect 5052 3736 5060 3744
rect 5084 3736 5092 3744
rect 5100 3736 5108 3744
rect 5132 3736 5140 3744
rect 5244 3736 5252 3744
rect 5388 3736 5396 3744
rect 5548 3736 5556 3744
rect 4972 3716 4980 3724
rect 5036 3716 5044 3724
rect 5212 3716 5220 3724
rect 5436 3716 5444 3724
rect 5500 3716 5508 3724
rect 5532 3716 5540 3724
rect 5580 3716 5588 3724
rect 5628 3716 5636 3724
rect 5676 3716 5684 3724
rect 5756 3716 5764 3724
rect 5788 3736 5796 3744
rect 5916 3736 5924 3744
rect 6172 3736 6180 3744
rect 6364 3736 6372 3744
rect 5868 3716 5876 3724
rect 5932 3716 5940 3724
rect 6028 3716 6036 3724
rect 6092 3716 6100 3724
rect 6140 3716 6148 3724
rect 6220 3716 6228 3724
rect 6284 3716 6292 3724
rect 6332 3716 6340 3724
rect 6348 3716 6356 3724
rect 6364 3716 6372 3724
rect 6444 3716 6452 3724
rect 6508 3736 6516 3744
rect 6604 3736 6612 3744
rect 2812 3696 2820 3704
rect 2892 3696 2900 3704
rect 3068 3696 3076 3704
rect 3516 3696 3524 3704
rect 3548 3696 3556 3704
rect 3580 3696 3588 3704
rect 3676 3696 3684 3704
rect 4124 3696 4132 3704
rect 4188 3696 4196 3704
rect 4236 3696 4244 3704
rect 4316 3696 4324 3704
rect 4444 3696 4452 3704
rect 4524 3696 4532 3704
rect 4588 3696 4596 3704
rect 4652 3696 4660 3704
rect 4748 3696 4756 3704
rect 4908 3696 4916 3704
rect 5052 3696 5060 3704
rect 5132 3696 5140 3704
rect 5228 3696 5236 3704
rect 5276 3696 5284 3704
rect 5452 3696 5460 3704
rect 5516 3696 5524 3704
rect 5596 3696 5604 3704
rect 5644 3696 5652 3704
rect 5660 3696 5668 3704
rect 5724 3696 5732 3704
rect 5804 3696 5812 3704
rect 5820 3696 5828 3704
rect 5884 3696 5892 3704
rect 6044 3696 6052 3704
rect 6124 3696 6132 3704
rect 6236 3696 6244 3704
rect 6284 3696 6292 3704
rect 6316 3696 6324 3704
rect 652 3676 660 3684
rect 1740 3676 1748 3684
rect 1836 3676 1844 3684
rect 2140 3676 2148 3684
rect 2236 3676 2244 3684
rect 2860 3676 2868 3684
rect 4156 3676 4164 3684
rect 4380 3676 4388 3684
rect 4492 3676 4500 3684
rect 4620 3676 4628 3684
rect 4652 3676 4660 3684
rect 5164 3676 5172 3684
rect 5196 3676 5204 3684
rect 5420 3676 5428 3684
rect 5484 3676 5492 3684
rect 5612 3676 5620 3684
rect 5852 3676 5860 3684
rect 5916 3676 5924 3684
rect 6044 3676 6052 3684
rect 6076 3676 6084 3684
rect 6156 3676 6164 3684
rect 6204 3676 6212 3684
rect 6268 3676 6276 3684
rect 6300 3676 6308 3684
rect 5500 3656 5508 3664
rect 6028 3656 6036 3664
rect 6284 3656 6292 3664
rect 524 3636 532 3644
rect 764 3636 772 3644
rect 1020 3636 1028 3644
rect 1132 3636 1140 3644
rect 1308 3636 1316 3644
rect 1452 3636 1460 3644
rect 1676 3636 1684 3644
rect 2044 3636 2052 3644
rect 2124 3636 2132 3644
rect 2540 3636 2548 3644
rect 2636 3636 2644 3644
rect 4140 3636 4148 3644
rect 4252 3636 4260 3644
rect 4508 3636 4516 3644
rect 4556 3636 4564 3644
rect 4636 3636 4644 3644
rect 5116 3636 5124 3644
rect 5356 3636 5364 3644
rect 5436 3636 5444 3644
rect 5708 3636 5716 3644
rect 5756 3636 5764 3644
rect 5868 3636 5876 3644
rect 5980 3636 5988 3644
rect 6092 3636 6100 3644
rect 6220 3636 6228 3644
rect 6460 3636 6468 3644
rect 1774 3606 1782 3614
rect 1788 3606 1796 3614
rect 1802 3606 1810 3614
rect 4830 3606 4838 3614
rect 4844 3606 4852 3614
rect 4858 3606 4866 3614
rect 204 3576 212 3584
rect 716 3576 724 3584
rect 2588 3576 2596 3584
rect 3244 3576 3252 3584
rect 3452 3576 3460 3584
rect 4188 3576 4196 3584
rect 4348 3576 4356 3584
rect 4476 3576 4484 3584
rect 4796 3576 4804 3584
rect 5404 3576 5412 3584
rect 5516 3576 5524 3584
rect 5644 3576 5652 3584
rect 5852 3576 5860 3584
rect 6092 3576 6100 3584
rect 6188 3576 6196 3584
rect 5580 3556 5588 3564
rect 1612 3536 1620 3544
rect 2204 3536 2212 3544
rect 3020 3536 3028 3544
rect 3660 3536 3668 3544
rect 3948 3536 3956 3544
rect 4012 3536 4020 3544
rect 5500 3536 5508 3544
rect 5596 3536 5604 3544
rect 5660 3536 5668 3544
rect 5836 3536 5844 3544
rect 6028 3536 6036 3544
rect 6108 3536 6116 3544
rect 6172 3536 6180 3544
rect 6332 3536 6340 3544
rect 6588 3536 6596 3544
rect 268 3516 276 3524
rect 76 3496 84 3504
rect 124 3496 132 3504
rect 348 3516 356 3524
rect 428 3516 436 3524
rect 652 3516 660 3524
rect 812 3516 820 3524
rect 844 3516 852 3524
rect 876 3516 884 3524
rect 316 3496 324 3504
rect 428 3496 436 3504
rect 524 3496 532 3504
rect 748 3496 756 3504
rect 940 3496 948 3504
rect 1052 3516 1060 3524
rect 1100 3516 1108 3524
rect 1628 3516 1636 3524
rect 1676 3516 1684 3524
rect 1756 3516 1764 3524
rect 2028 3516 2036 3524
rect 2044 3516 2052 3524
rect 2092 3516 2100 3524
rect 2156 3516 2164 3524
rect 2220 3516 2228 3524
rect 2316 3516 2324 3524
rect 2524 3516 2532 3524
rect 2812 3516 2820 3524
rect 2956 3516 2964 3524
rect 3052 3516 3060 3524
rect 3340 3516 3348 3524
rect 3372 3516 3380 3524
rect 3420 3516 3428 3524
rect 3676 3516 3684 3524
rect 4028 3516 4036 3524
rect 4284 3516 4292 3524
rect 4380 3516 4388 3524
rect 4444 3516 4452 3524
rect 4460 3516 4468 3524
rect 4604 3516 4612 3524
rect 4636 3516 4644 3524
rect 4780 3516 4788 3524
rect 4924 3516 4932 3524
rect 5468 3516 5476 3524
rect 5548 3516 5556 3524
rect 5564 3516 5572 3524
rect 5628 3516 5636 3524
rect 5804 3516 5812 3524
rect 5868 3516 5876 3524
rect 6060 3516 6068 3524
rect 6076 3516 6084 3524
rect 6140 3516 6148 3524
rect 6268 3516 6276 3524
rect 6364 3516 6372 3524
rect 6540 3516 6548 3524
rect 6556 3516 6564 3524
rect 1020 3496 1028 3504
rect 1180 3496 1188 3504
rect 1324 3496 1332 3504
rect 1484 3494 1492 3502
rect 268 3476 276 3484
rect 348 3476 356 3484
rect 380 3476 388 3484
rect 444 3476 452 3484
rect 508 3476 516 3484
rect 684 3476 692 3484
rect 764 3476 772 3484
rect 796 3476 804 3484
rect 844 3476 852 3484
rect 924 3476 932 3484
rect 988 3476 996 3484
rect 1068 3476 1076 3484
rect 1164 3476 1172 3484
rect 1196 3476 1204 3484
rect 1404 3476 1412 3484
rect 1516 3476 1524 3484
rect 1660 3476 1668 3484
rect 1708 3476 1716 3484
rect 1820 3496 1828 3504
rect 2124 3496 2132 3504
rect 2140 3496 2148 3504
rect 2460 3494 2468 3502
rect 2524 3496 2532 3504
rect 2556 3496 2564 3504
rect 2700 3496 2708 3504
rect 2828 3496 2836 3504
rect 2892 3496 2900 3504
rect 3020 3496 3028 3504
rect 3116 3494 3124 3502
rect 3260 3496 3268 3504
rect 3532 3494 3540 3502
rect 3692 3496 3700 3504
rect 3820 3494 3828 3502
rect 4028 3496 4036 3504
rect 4108 3496 4116 3504
rect 4220 3496 4228 3504
rect 4348 3496 4356 3504
rect 4412 3496 4420 3504
rect 4540 3496 4548 3504
rect 4556 3496 4564 3504
rect 4652 3496 4660 3504
rect 4716 3496 4724 3504
rect 4732 3496 4740 3504
rect 4796 3496 4804 3504
rect 5052 3496 5060 3504
rect 5324 3496 5332 3504
rect 5340 3496 5348 3504
rect 5420 3496 5428 3504
rect 5484 3496 5492 3504
rect 5580 3496 5588 3504
rect 5644 3496 5652 3504
rect 5772 3496 5780 3504
rect 5804 3496 5812 3504
rect 5852 3496 5860 3504
rect 5932 3496 5940 3504
rect 5996 3496 6004 3504
rect 6044 3496 6052 3504
rect 6092 3496 6100 3504
rect 6156 3496 6164 3504
rect 6348 3496 6356 3504
rect 6380 3496 6388 3504
rect 6492 3496 6500 3504
rect 6572 3496 6580 3504
rect 1836 3476 1844 3484
rect 1868 3476 1876 3484
rect 1980 3476 1988 3484
rect 1996 3476 2004 3484
rect 2028 3476 2036 3484
rect 2076 3476 2084 3484
rect 2156 3476 2164 3484
rect 2188 3476 2196 3484
rect 2284 3476 2292 3484
rect 2428 3476 2436 3484
rect 2572 3476 2580 3484
rect 2684 3476 2692 3484
rect 2748 3476 2756 3484
rect 2780 3476 2788 3484
rect 2860 3476 2868 3484
rect 2940 3476 2948 3484
rect 2988 3476 2996 3484
rect 3084 3476 3092 3484
rect 3260 3476 3268 3484
rect 3388 3476 3396 3484
rect 3468 3476 3476 3484
rect 3580 3476 3588 3484
rect 3724 3476 3732 3484
rect 3788 3476 3796 3484
rect 4092 3476 4100 3484
rect 4156 3480 4164 3488
rect 4172 3476 4180 3484
rect 4236 3476 4244 3484
rect 4252 3476 4260 3484
rect 4332 3476 4340 3484
rect 4396 3476 4404 3484
rect 4428 3476 4436 3484
rect 4492 3476 4500 3484
rect 4540 3476 4548 3484
rect 4652 3476 4660 3484
rect 4700 3476 4708 3484
rect 4716 3476 4724 3484
rect 4892 3476 4900 3484
rect 4940 3476 4948 3484
rect 5036 3476 5044 3484
rect 5180 3476 5188 3484
rect 5196 3476 5204 3484
rect 5292 3476 5300 3484
rect 220 3456 228 3464
rect 812 3456 820 3464
rect 876 3456 884 3464
rect 892 3456 900 3464
rect 1052 3456 1060 3464
rect 1228 3456 1236 3464
rect 1868 3456 1876 3464
rect 2220 3456 2228 3464
rect 2972 3456 2980 3464
rect 3420 3456 3428 3464
rect 3532 3456 3540 3464
rect 3756 3456 3764 3464
rect 3964 3456 3972 3464
rect 3996 3456 4004 3464
rect 4060 3456 4068 3464
rect 4300 3456 4308 3464
rect 4508 3456 4516 3464
rect 4700 3456 4708 3464
rect 4828 3456 4836 3464
rect 5068 3456 5076 3464
rect 5388 3476 5396 3484
rect 5692 3476 5700 3484
rect 5916 3476 5924 3484
rect 5980 3476 5988 3484
rect 6236 3476 6244 3484
rect 6300 3476 6308 3484
rect 6396 3476 6404 3484
rect 5420 3456 5428 3464
rect 5452 3456 5460 3464
rect 5532 3456 5540 3464
rect 5740 3456 5748 3464
rect 5884 3456 5892 3464
rect 5948 3456 5956 3464
rect 6204 3456 6212 3464
rect 6348 3456 6356 3464
rect 6428 3456 6436 3464
rect 6476 3476 6484 3484
rect 6508 3476 6516 3484
rect 188 3436 196 3444
rect 636 3436 644 3444
rect 668 3436 676 3444
rect 908 3436 916 3444
rect 956 3436 964 3444
rect 1212 3436 1220 3444
rect 1244 3436 1252 3444
rect 1628 3436 1636 3444
rect 1676 3436 1684 3444
rect 1740 3436 1748 3444
rect 1852 3436 1860 3444
rect 1916 3436 1924 3444
rect 2012 3436 2020 3444
rect 2092 3436 2100 3444
rect 2236 3436 2244 3444
rect 2300 3436 2308 3444
rect 2332 3436 2340 3444
rect 2796 3436 2804 3444
rect 3244 3436 3252 3444
rect 3436 3436 3444 3444
rect 3980 3436 3988 3444
rect 4076 3436 4084 3444
rect 4124 3436 4132 3444
rect 4188 3436 4196 3444
rect 4268 3436 4276 3444
rect 4620 3436 4628 3444
rect 4780 3436 4788 3444
rect 4908 3436 4916 3444
rect 5004 3436 5012 3444
rect 5116 3436 5124 3444
rect 5228 3436 5236 3444
rect 5356 3436 5364 3444
rect 5436 3436 5444 3444
rect 5724 3436 5732 3444
rect 5900 3436 5908 3444
rect 5964 3436 5972 3444
rect 6220 3436 6228 3444
rect 6460 3436 6468 3444
rect 6524 3436 6532 3444
rect 6604 3436 6612 3444
rect 3310 3406 3318 3414
rect 3324 3406 3332 3414
rect 3338 3406 3346 3414
rect 124 3376 132 3384
rect 332 3376 340 3384
rect 652 3376 660 3384
rect 940 3376 948 3384
rect 1260 3376 1268 3384
rect 1932 3376 1940 3384
rect 2540 3376 2548 3384
rect 2668 3376 2676 3384
rect 2956 3376 2964 3384
rect 3356 3376 3364 3384
rect 3532 3376 3540 3384
rect 3740 3376 3748 3384
rect 4140 3376 4148 3384
rect 5004 3376 5012 3384
rect 5180 3376 5188 3384
rect 5420 3376 5428 3384
rect 5628 3376 5636 3384
rect 380 3356 388 3364
rect 540 3356 548 3364
rect 556 3356 564 3364
rect 748 3356 756 3364
rect 908 3356 916 3364
rect 1500 3356 1508 3364
rect 1596 3356 1604 3364
rect 1644 3356 1652 3364
rect 2428 3356 2436 3364
rect 2572 3356 2580 3364
rect 2940 3356 2948 3364
rect 3164 3356 3172 3364
rect 3900 3356 3908 3364
rect 4780 3356 4788 3364
rect 5100 3356 5108 3364
rect 5372 3356 5380 3364
rect 5612 3356 5620 3364
rect 5788 3356 5796 3364
rect 5836 3356 5844 3364
rect 12 3336 20 3344
rect 172 3336 180 3344
rect 476 3336 484 3344
rect 524 3336 532 3344
rect 588 3336 596 3344
rect 620 3336 628 3344
rect 636 3336 644 3344
rect 780 3336 788 3344
rect 924 3336 932 3344
rect 956 3336 964 3344
rect 972 3336 980 3344
rect 1036 3336 1044 3344
rect 1068 3336 1076 3344
rect 1100 3336 1108 3344
rect 1372 3336 1380 3344
rect 1388 3336 1396 3344
rect 1468 3336 1476 3344
rect 1644 3336 1652 3344
rect 1708 3336 1716 3344
rect 1724 3332 1732 3340
rect 1772 3336 1780 3344
rect 1868 3336 1876 3344
rect 1916 3336 1924 3344
rect 2060 3336 2068 3344
rect 2124 3336 2132 3344
rect 2156 3336 2164 3344
rect 2220 3336 2228 3344
rect 2252 3336 2260 3344
rect 2348 3336 2356 3344
rect 2460 3336 2468 3344
rect 2524 3336 2532 3344
rect 2604 3336 2612 3344
rect 2908 3336 2916 3344
rect 3116 3336 3124 3344
rect 3164 3336 3172 3344
rect 3404 3336 3412 3344
rect 3580 3336 3588 3344
rect 3980 3336 3988 3344
rect 4092 3336 4100 3344
rect 4188 3336 4196 3344
rect 4204 3336 4212 3344
rect 4364 3336 4372 3344
rect 4524 3336 4532 3344
rect 4572 3336 4580 3344
rect 4748 3336 4756 3344
rect 4940 3336 4948 3344
rect 5340 3336 5348 3344
rect 5372 3336 5380 3344
rect 5452 3336 5460 3344
rect 5548 3336 5556 3344
rect 5596 3336 5604 3344
rect 5644 3336 5652 3344
rect 5676 3336 5684 3344
rect 5772 3336 5780 3344
rect 5900 3336 5908 3344
rect 5932 3336 5940 3344
rect 5980 3336 5988 3344
rect 6028 3356 6036 3364
rect 6092 3356 6100 3364
rect 6108 3356 6116 3364
rect 6428 3356 6436 3364
rect 6044 3336 6052 3344
rect 6172 3336 6180 3344
rect 6460 3336 6468 3344
rect 236 3316 244 3324
rect 380 3316 388 3324
rect 412 3316 420 3324
rect 460 3316 468 3324
rect 460 3296 468 3304
rect 524 3316 532 3324
rect 604 3316 612 3324
rect 732 3316 740 3324
rect 764 3316 772 3324
rect 796 3316 804 3324
rect 844 3316 852 3324
rect 876 3316 884 3324
rect 988 3316 996 3324
rect 1132 3318 1140 3326
rect 572 3296 580 3304
rect 668 3296 676 3304
rect 700 3296 708 3304
rect 860 3296 868 3304
rect 924 3296 932 3304
rect 1196 3316 1204 3324
rect 1036 3296 1044 3304
rect 1308 3296 1316 3304
rect 1372 3316 1380 3324
rect 1404 3316 1412 3324
rect 1452 3316 1460 3324
rect 1484 3316 1492 3324
rect 1548 3316 1556 3324
rect 1612 3316 1620 3324
rect 1804 3316 1812 3324
rect 1852 3316 1860 3324
rect 1356 3296 1364 3304
rect 1436 3296 1444 3304
rect 1564 3296 1572 3304
rect 1660 3296 1668 3304
rect 1820 3296 1828 3304
rect 2044 3316 2052 3324
rect 2156 3296 2164 3304
rect 2204 3316 2212 3324
rect 2300 3316 2308 3324
rect 2492 3316 2500 3324
rect 2652 3316 2660 3324
rect 2732 3316 2740 3324
rect 2764 3316 2772 3324
rect 3068 3316 3076 3324
rect 3228 3318 3236 3326
rect 3292 3316 3300 3324
rect 3612 3318 3620 3326
rect 3788 3316 3796 3324
rect 3852 3316 3860 3324
rect 3900 3316 3908 3324
rect 3996 3316 4004 3324
rect 4076 3316 4084 3324
rect 4108 3316 4116 3324
rect 4236 3316 4244 3324
rect 4284 3316 4292 3324
rect 4332 3316 4340 3324
rect 4348 3316 4356 3324
rect 4412 3316 4420 3324
rect 4460 3316 4468 3324
rect 4540 3316 4548 3324
rect 4636 3316 4644 3324
rect 4684 3316 4692 3324
rect 4732 3316 4740 3324
rect 4828 3316 4836 3324
rect 4940 3316 4948 3324
rect 5004 3316 5012 3324
rect 5068 3316 5076 3324
rect 5148 3316 5156 3324
rect 5228 3316 5236 3324
rect 5292 3316 5300 3324
rect 5324 3316 5332 3324
rect 5420 3316 5428 3324
rect 5468 3316 5476 3324
rect 2508 3296 2516 3304
rect 2556 3296 2564 3304
rect 2652 3296 2660 3304
rect 2860 3296 2868 3304
rect 2892 3296 2900 3304
rect 3804 3296 3812 3304
rect 3868 3296 3876 3304
rect 3916 3296 3924 3304
rect 4028 3296 4036 3304
rect 4044 3296 4052 3304
rect 4156 3296 4164 3304
rect 4236 3296 4244 3304
rect 4284 3296 4292 3304
rect 4316 3296 4324 3304
rect 4444 3296 4452 3304
rect 4556 3296 4564 3304
rect 4588 3296 4596 3304
rect 4652 3296 4660 3304
rect 4668 3296 4676 3304
rect 4844 3296 4852 3304
rect 4956 3296 4964 3304
rect 5020 3296 5028 3304
rect 5244 3296 5252 3304
rect 5308 3296 5316 3304
rect 5436 3296 5444 3304
rect 5500 3296 5508 3304
rect 5660 3316 5668 3324
rect 5900 3316 5908 3324
rect 5980 3316 5988 3324
rect 6156 3316 6164 3324
rect 6220 3316 6228 3324
rect 6348 3316 6356 3324
rect 5788 3296 5796 3304
rect 5932 3296 5940 3304
rect 5964 3296 5972 3304
rect 5996 3296 6004 3304
rect 6124 3296 6132 3304
rect 6156 3296 6164 3304
rect 6252 3296 6260 3304
rect 6524 3300 6532 3308
rect 828 3276 836 3284
rect 1516 3276 1524 3284
rect 1532 3276 1540 3284
rect 1916 3276 1924 3284
rect 2428 3276 2436 3284
rect 3772 3276 3780 3284
rect 3804 3276 3812 3284
rect 3836 3276 3844 3284
rect 3996 3276 4004 3284
rect 4268 3276 4276 3284
rect 4396 3276 4404 3284
rect 4476 3276 4484 3284
rect 4524 3276 4532 3284
rect 4620 3276 4628 3284
rect 4812 3276 4820 3284
rect 4924 3276 4932 3284
rect 5004 3276 5012 3284
rect 5052 3276 5060 3284
rect 5164 3276 5172 3284
rect 5212 3276 5220 3284
rect 5276 3276 5284 3284
rect 5404 3276 5412 3284
rect 5884 3276 5892 3284
rect 6204 3276 6212 3284
rect 4412 3256 4420 3264
rect 4780 3256 4788 3264
rect 4828 3256 4836 3264
rect 5068 3256 5076 3264
rect 5228 3256 5236 3264
rect 5292 3256 5300 3264
rect 6524 3254 6532 3262
rect 124 3236 132 3244
rect 812 3236 820 3244
rect 1260 3236 1268 3244
rect 1404 3236 1412 3244
rect 1580 3236 1588 3244
rect 1628 3236 1636 3244
rect 1900 3236 1908 3244
rect 3148 3236 3156 3244
rect 3756 3236 3764 3244
rect 4076 3236 4084 3244
rect 4172 3236 4180 3244
rect 4284 3236 4292 3244
rect 4460 3236 4468 3244
rect 4636 3236 4644 3244
rect 4716 3236 4724 3244
rect 5580 3236 5588 3244
rect 5740 3236 5748 3244
rect 6076 3236 6084 3244
rect 6220 3236 6228 3244
rect 6268 3236 6276 3244
rect 1774 3206 1782 3214
rect 1788 3206 1796 3214
rect 1802 3206 1810 3214
rect 4830 3206 4838 3214
rect 4844 3206 4852 3214
rect 4858 3206 4866 3214
rect 188 3176 196 3184
rect 572 3176 580 3184
rect 924 3176 932 3184
rect 1212 3176 1220 3184
rect 2012 3176 2020 3184
rect 2444 3176 2452 3184
rect 3100 3176 3108 3184
rect 4060 3176 4068 3184
rect 4700 3176 4708 3184
rect 4892 3176 4900 3184
rect 5052 3176 5060 3184
rect 5132 3176 5140 3184
rect 5900 3176 5908 3184
rect 6028 3176 6036 3184
rect 6268 3176 6276 3184
rect 6508 3176 6516 3184
rect 2492 3156 2500 3164
rect 4380 3156 4388 3164
rect 4572 3156 4580 3164
rect 4636 3156 4644 3164
rect 4764 3156 4772 3164
rect 5564 3156 5572 3164
rect 668 3136 676 3144
rect 1628 3136 1636 3144
rect 2828 3136 2836 3144
rect 3452 3136 3460 3144
rect 4092 3136 4100 3144
rect 4284 3136 4292 3144
rect 4364 3136 4372 3144
rect 4556 3136 4564 3144
rect 4620 3136 4628 3144
rect 4684 3136 4692 3144
rect 4748 3136 4756 3144
rect 4796 3136 4804 3144
rect 4940 3136 4948 3144
rect 5068 3136 5076 3144
rect 5116 3136 5124 3144
rect 5580 3136 5588 3144
rect 5628 3136 5636 3144
rect 5708 3136 5716 3144
rect 5820 3136 5828 3144
rect 5884 3136 5892 3144
rect 5964 3136 5972 3144
rect 6012 3136 6020 3144
rect 6092 3136 6100 3144
rect 6108 3136 6116 3144
rect 6140 3136 6148 3144
rect 636 3116 644 3124
rect 972 3116 980 3124
rect 988 3116 996 3124
rect 1020 3116 1028 3124
rect 1052 3116 1060 3124
rect 1292 3116 1300 3124
rect 1324 3116 1332 3124
rect 1388 3116 1396 3124
rect 1436 3116 1444 3124
rect 1532 3116 1540 3124
rect 1580 3116 1588 3124
rect 1708 3116 1716 3124
rect 2428 3116 2436 3124
rect 2540 3116 2548 3124
rect 76 3096 84 3104
rect 124 3096 132 3104
rect 300 3096 308 3104
rect 364 3094 372 3102
rect 508 3096 516 3104
rect 652 3096 660 3104
rect 700 3096 708 3104
rect 732 3096 740 3104
rect 796 3094 804 3102
rect 860 3096 868 3104
rect 1052 3096 1060 3104
rect 1100 3096 1108 3104
rect 1340 3096 1348 3104
rect 1356 3096 1364 3104
rect 1500 3096 1508 3104
rect 1612 3096 1620 3104
rect 1676 3096 1684 3104
rect 1724 3096 1732 3104
rect 1756 3096 1764 3104
rect 1980 3096 1988 3104
rect 2108 3096 2116 3104
rect 2156 3096 2164 3104
rect 2316 3096 2324 3104
rect 2940 3116 2948 3124
rect 3052 3116 3060 3124
rect 2572 3096 2580 3104
rect 2700 3094 2708 3102
rect 2844 3096 2852 3104
rect 2956 3096 2964 3104
rect 3132 3116 3140 3124
rect 3692 3116 3700 3124
rect 3740 3116 3748 3124
rect 3788 3116 3796 3124
rect 3868 3116 3876 3124
rect 3964 3116 3972 3124
rect 4108 3116 4116 3124
rect 4172 3116 4180 3124
rect 4220 3116 4228 3124
rect 4396 3116 4404 3124
rect 4588 3116 4596 3124
rect 4652 3116 4660 3124
rect 4716 3116 4724 3124
rect 4780 3116 4788 3124
rect 4908 3116 4916 3124
rect 5020 3116 5028 3124
rect 5036 3116 5044 3124
rect 5148 3116 5156 3124
rect 5516 3116 5524 3124
rect 5596 3116 5604 3124
rect 5708 3116 5716 3124
rect 5788 3116 5796 3124
rect 5852 3116 5860 3124
rect 6060 3116 6068 3124
rect 6172 3116 6180 3124
rect 6220 3116 6228 3124
rect 3100 3096 3108 3104
rect 3148 3096 3156 3104
rect 3324 3094 3332 3102
rect 3388 3096 3396 3104
rect 3548 3096 3556 3104
rect 3580 3096 3588 3104
rect 3916 3096 3924 3104
rect 3980 3096 3988 3104
rect 4044 3096 4052 3104
rect 4092 3096 4100 3104
rect 4124 3096 4132 3104
rect 4172 3096 4180 3104
rect 4268 3096 4276 3104
rect 4332 3096 4340 3104
rect 4380 3096 4388 3104
rect 4412 3096 4420 3104
rect 4492 3096 4500 3104
rect 4572 3096 4580 3104
rect 4636 3096 4644 3104
rect 4700 3096 4708 3104
rect 4764 3096 4772 3104
rect 4812 3096 4820 3104
rect 4924 3096 4932 3104
rect 4972 3096 4980 3104
rect 4988 3096 4996 3104
rect 5052 3096 5060 3104
rect 5132 3096 5140 3104
rect 5164 3096 5172 3104
rect 5228 3096 5236 3104
rect 5324 3096 5332 3104
rect 5404 3096 5412 3104
rect 5516 3096 5524 3104
rect 5564 3096 5572 3104
rect 5612 3096 5620 3104
rect 5692 3096 5700 3104
rect 5724 3096 5732 3104
rect 5788 3096 5796 3104
rect 5820 3096 5828 3104
rect 5868 3096 5876 3104
rect 5932 3096 5940 3104
rect 5964 3096 5972 3104
rect 6028 3096 6036 3104
rect 6076 3096 6084 3104
rect 6156 3096 6164 3104
rect 6236 3096 6244 3104
rect 6348 3096 6356 3104
rect 6476 3096 6484 3104
rect 204 3076 212 3084
rect 300 3076 308 3084
rect 332 3076 340 3084
rect 940 3076 948 3084
rect 1036 3076 1044 3084
rect 1084 3076 1092 3084
rect 1148 3076 1156 3084
rect 1244 3076 1252 3084
rect 1292 3076 1300 3084
rect 1324 3076 1332 3084
rect 1468 3076 1476 3084
rect 1484 3076 1492 3084
rect 1532 3076 1540 3084
rect 1548 3076 1556 3084
rect 1740 3076 1748 3084
rect 1836 3076 1844 3084
rect 1964 3076 1972 3084
rect 2060 3076 2068 3084
rect 2252 3076 2260 3084
rect 2460 3076 2468 3084
rect 2508 3076 2516 3084
rect 2604 3076 2612 3084
rect 2732 3076 2740 3084
rect 2860 3076 2868 3084
rect 2908 3076 2916 3084
rect 3020 3076 3028 3084
rect 3116 3076 3124 3084
rect 3180 3076 3188 3084
rect 3292 3076 3300 3084
rect 3484 3076 3492 3084
rect 3660 3076 3668 3084
rect 3708 3076 3716 3084
rect 3756 3076 3764 3084
rect 3836 3076 3844 3084
rect 3932 3076 3940 3084
rect 3996 3076 4004 3084
rect 4028 3076 4036 3084
rect 4124 3076 4132 3084
rect 4316 3076 4324 3084
rect 4428 3076 4436 3084
rect 540 3056 548 3064
rect 588 3056 596 3064
rect 604 3056 612 3064
rect 620 3056 628 3064
rect 732 3056 740 3064
rect 1132 3056 1140 3064
rect 1260 3056 1268 3064
rect 1404 3056 1412 3064
rect 1772 3056 1780 3064
rect 2476 3056 2484 3064
rect 2636 3056 2644 3064
rect 2892 3056 2900 3064
rect 2988 3056 2996 3064
rect 3260 3056 3268 3064
rect 3788 3056 3796 3064
rect 3820 3056 3828 3064
rect 3884 3056 3892 3064
rect 4028 3056 4036 3064
rect 4236 3056 4244 3064
rect 4460 3056 4468 3064
rect 4508 3076 4516 3084
rect 4972 3076 4980 3084
rect 5180 3076 5188 3084
rect 5228 3076 5236 3084
rect 5244 3076 5252 3084
rect 5292 3076 5300 3084
rect 5388 3076 5396 3084
rect 5452 3076 5460 3084
rect 5740 3076 5748 3084
rect 5836 3076 5844 3084
rect 5916 3076 5924 3084
rect 5980 3076 5988 3084
rect 6156 3076 6164 3084
rect 6188 3076 6196 3084
rect 6300 3076 6308 3084
rect 6364 3076 6372 3084
rect 6524 3076 6532 3084
rect 6620 3076 6628 3084
rect 5212 3056 5220 3064
rect 5276 3056 5284 3064
rect 5452 3056 5460 3064
rect 5772 3056 5780 3064
rect 492 3036 500 3044
rect 684 3036 692 3044
rect 972 3036 980 3044
rect 1068 3036 1076 3044
rect 1116 3036 1124 3044
rect 1388 3036 1396 3044
rect 1420 3036 1428 3044
rect 1580 3036 1588 3044
rect 1708 3036 1716 3044
rect 2220 3036 2228 3044
rect 2412 3036 2420 3044
rect 2428 3036 2436 3044
rect 2540 3036 2548 3044
rect 2876 3036 2884 3044
rect 2940 3036 2948 3044
rect 3036 3036 3044 3044
rect 3644 3036 3652 3044
rect 3692 3036 3700 3044
rect 3740 3036 3748 3044
rect 3804 3036 3812 3044
rect 3900 3036 3908 3044
rect 3948 3036 3956 3044
rect 5020 3036 5028 3044
rect 5356 3036 5364 3044
rect 5644 3036 5652 3044
rect 5692 3036 5700 3044
rect 6220 3036 6228 3044
rect 6460 3036 6468 3044
rect 6556 3036 6564 3044
rect 3310 3006 3318 3014
rect 3324 3006 3332 3014
rect 3338 3006 3346 3014
rect 220 2976 228 2984
rect 540 2976 548 2984
rect 620 2976 628 2984
rect 796 2976 804 2984
rect 1164 2976 1172 2984
rect 1228 2976 1236 2984
rect 1516 2976 1524 2984
rect 2332 2976 2340 2984
rect 2524 2976 2532 2984
rect 2908 2976 2916 2984
rect 3372 2976 3380 2984
rect 3756 2976 3764 2984
rect 4012 2976 4020 2984
rect 4220 2976 4228 2984
rect 5500 2976 5508 2984
rect 5836 2976 5844 2984
rect 5900 2976 5908 2984
rect 5948 2976 5956 2984
rect 6044 2976 6052 2984
rect 6156 2976 6164 2984
rect 6380 2976 6388 2984
rect 6476 2976 6484 2984
rect 6572 2976 6580 2984
rect 380 2956 388 2964
rect 524 2956 532 2964
rect 636 2956 644 2964
rect 716 2956 724 2964
rect 780 2956 788 2964
rect 908 2956 916 2964
rect 1004 2956 1012 2964
rect 1084 2956 1092 2964
rect 1612 2956 1620 2964
rect 1900 2956 1908 2964
rect 1964 2956 1972 2964
rect 2060 2956 2068 2964
rect 2412 2956 2420 2964
rect 2780 2956 2788 2964
rect 2828 2956 2836 2964
rect 2860 2956 2868 2964
rect 2892 2956 2900 2964
rect 3100 2956 3108 2964
rect 3564 2956 3572 2964
rect 4076 2956 4084 2964
rect 4140 2956 4148 2964
rect 4492 2956 4500 2964
rect 4652 2956 4660 2964
rect 5244 2956 5252 2964
rect 5388 2956 5396 2964
rect 5404 2956 5412 2964
rect 5516 2956 5524 2964
rect 5660 2956 5668 2964
rect 5756 2956 5764 2964
rect 5852 2956 5860 2964
rect 6028 2956 6036 2964
rect 44 2936 52 2944
rect 172 2936 180 2944
rect 204 2936 212 2944
rect 412 2936 420 2944
rect 428 2936 436 2944
rect 492 2936 500 2944
rect 604 2936 612 2944
rect 812 2936 820 2944
rect 940 2936 948 2944
rect 988 2936 996 2944
rect 1068 2936 1076 2944
rect 1260 2936 1268 2944
rect 1500 2936 1508 2944
rect 1548 2936 1556 2944
rect 1692 2936 1700 2944
rect 1932 2936 1940 2944
rect 1964 2936 1972 2944
rect 2012 2936 2020 2944
rect 2316 2936 2324 2944
rect 2380 2936 2388 2944
rect 2460 2936 2468 2944
rect 2476 2936 2484 2944
rect 2684 2936 2692 2944
rect 2716 2936 2724 2944
rect 2764 2936 2772 2944
rect 2828 2936 2836 2944
rect 3020 2936 3028 2944
rect 3132 2936 3140 2944
rect 3212 2936 3220 2944
rect 3500 2936 3508 2944
rect 3532 2936 3540 2944
rect 3596 2936 3604 2944
rect 3692 2936 3700 2944
rect 3820 2936 3828 2944
rect 3852 2936 3860 2944
rect 4044 2936 4052 2944
rect 4060 2936 4068 2944
rect 4156 2936 4164 2944
rect 4252 2936 4260 2944
rect 4268 2936 4276 2944
rect 4364 2936 4372 2944
rect 4460 2936 4468 2944
rect 4508 2936 4516 2944
rect 4572 2936 4580 2944
rect 4876 2936 4884 2944
rect 4972 2936 4980 2944
rect 5020 2936 5028 2944
rect 5052 2936 5060 2944
rect 5068 2936 5076 2944
rect 5164 2936 5172 2944
rect 5276 2936 5284 2944
rect 5340 2936 5348 2944
rect 5356 2936 5364 2944
rect 5420 2936 5428 2944
rect 5484 2936 5492 2944
rect 5596 2936 5604 2944
rect 5756 2936 5764 2944
rect 5788 2936 5796 2944
rect 5964 2936 5972 2944
rect 6028 2936 6036 2944
rect 6060 2936 6068 2944
rect 6188 2936 6196 2944
rect 6284 2936 6292 2944
rect 6300 2936 6308 2944
rect 44 2916 52 2924
rect 108 2916 116 2924
rect 172 2916 180 2924
rect 268 2916 276 2924
rect 332 2916 340 2924
rect 444 2916 452 2924
rect 476 2916 484 2924
rect 588 2916 596 2924
rect 652 2916 660 2924
rect 684 2916 692 2924
rect 748 2916 756 2924
rect 828 2916 836 2924
rect 908 2916 916 2924
rect 940 2916 948 2924
rect 1100 2916 1108 2924
rect 1196 2916 1204 2924
rect 1340 2916 1348 2924
rect 1580 2916 1588 2924
rect 1676 2918 1684 2926
rect 1868 2916 1876 2924
rect 1996 2916 2004 2924
rect 2140 2916 2148 2924
rect 2204 2918 2212 2926
rect 2268 2916 2276 2924
rect 2300 2916 2308 2924
rect 2508 2916 2516 2924
rect 2652 2918 2660 2926
rect 2748 2916 2756 2924
rect 2812 2916 2820 2924
rect 2860 2916 2868 2924
rect 3004 2916 3012 2924
rect 3180 2916 3188 2924
rect 3244 2918 3252 2926
rect 3388 2916 3396 2924
rect 3628 2918 3636 2926
rect 3804 2916 3812 2924
rect 3884 2918 3892 2926
rect 4060 2916 4068 2924
rect 4412 2916 4420 2924
rect 4444 2916 4452 2924
rect 4524 2916 4532 2924
rect 4588 2916 4596 2924
rect 4620 2916 4628 2924
rect 4652 2916 4660 2924
rect 4684 2916 4692 2924
rect 4748 2916 4756 2924
rect 4812 2916 4820 2924
rect 4924 2916 4932 2924
rect 4972 2916 4980 2924
rect 5020 2916 5028 2924
rect 5212 2916 5220 2924
rect 5260 2916 5268 2924
rect 5292 2916 5300 2924
rect 5356 2916 5364 2924
rect 5468 2916 5476 2924
rect 5548 2916 5556 2924
rect 5612 2916 5620 2924
rect 5644 2916 5652 2924
rect 5708 2916 5716 2924
rect 5804 2916 5812 2924
rect 5884 2916 5892 2924
rect 6076 2916 6084 2924
rect 6108 2916 6116 2924
rect 6252 2918 6260 2926
rect 6396 2916 6404 2924
rect 6444 2916 6452 2924
rect 6492 2916 6500 2924
rect 6540 2916 6548 2924
rect 6588 2916 6596 2924
rect 60 2896 68 2904
rect 124 2896 132 2904
rect 188 2896 196 2904
rect 236 2896 244 2904
rect 252 2896 260 2904
rect 316 2896 324 2904
rect 380 2896 388 2904
rect 444 2896 452 2904
rect 540 2896 548 2904
rect 700 2896 708 2904
rect 764 2896 772 2904
rect 844 2896 852 2904
rect 940 2896 948 2904
rect 1212 2896 1220 2904
rect 1228 2896 1236 2904
rect 1260 2896 1268 2904
rect 1356 2896 1364 2904
rect 1516 2896 1524 2904
rect 1612 2896 1620 2904
rect 2268 2896 2276 2904
rect 2332 2896 2340 2904
rect 2412 2896 2420 2904
rect 2508 2896 2516 2904
rect 2716 2896 2724 2904
rect 3180 2896 3188 2904
rect 3484 2896 3492 2904
rect 3772 2896 3780 2904
rect 4028 2896 4036 2904
rect 4332 2896 4340 2904
rect 4428 2896 4436 2904
rect 4556 2896 4564 2904
rect 4668 2896 4676 2904
rect 4732 2896 4740 2904
rect 4796 2896 4804 2904
rect 4892 2896 4900 2904
rect 5004 2896 5012 2904
rect 5052 2896 5060 2904
rect 5132 2896 5140 2904
rect 5228 2896 5236 2904
rect 5308 2896 5316 2904
rect 5388 2896 5396 2904
rect 5532 2896 5540 2904
rect 5580 2896 5588 2904
rect 5660 2896 5668 2904
rect 5756 2896 5764 2904
rect 5868 2896 5876 2904
rect 6012 2896 6020 2904
rect 6092 2896 6100 2904
rect 28 2876 36 2884
rect 92 2876 100 2884
rect 156 2876 164 2884
rect 252 2876 260 2884
rect 284 2876 292 2884
rect 316 2876 324 2884
rect 524 2876 532 2884
rect 668 2876 676 2884
rect 732 2876 740 2884
rect 956 2876 964 2884
rect 1020 2876 1028 2884
rect 1356 2876 1364 2884
rect 1804 2876 1812 2884
rect 3468 2876 3476 2884
rect 4396 2876 4404 2884
rect 4700 2876 4708 2884
rect 4748 2876 4756 2884
rect 4764 2876 4772 2884
rect 4828 2876 4836 2884
rect 4940 2876 4948 2884
rect 5196 2876 5204 2884
rect 5564 2876 5572 2884
rect 5724 2876 5732 2884
rect 5900 2876 5908 2884
rect 6092 2876 6100 2884
rect 6428 2876 6436 2884
rect 3804 2856 3812 2864
rect 4412 2856 4420 2864
rect 4748 2856 4756 2864
rect 5212 2856 5220 2864
rect 108 2836 116 2844
rect 220 2836 228 2844
rect 332 2836 340 2844
rect 1116 2836 1124 2844
rect 1388 2836 1396 2844
rect 1964 2836 1972 2844
rect 2076 2836 2084 2844
rect 2444 2836 2452 2844
rect 2860 2836 2868 2844
rect 4124 2836 4132 2844
rect 4524 2836 4532 2844
rect 6524 2836 6532 2844
rect 6620 2836 6628 2844
rect 1774 2806 1782 2814
rect 1788 2806 1796 2814
rect 1802 2806 1810 2814
rect 4830 2806 4838 2814
rect 4844 2806 4852 2814
rect 4858 2806 4866 2814
rect 76 2776 84 2784
rect 492 2776 500 2784
rect 636 2776 644 2784
rect 716 2776 724 2784
rect 908 2776 916 2784
rect 940 2776 948 2784
rect 1116 2776 1124 2784
rect 1212 2776 1220 2784
rect 1324 2776 1332 2784
rect 1356 2776 1364 2784
rect 1452 2776 1460 2784
rect 2892 2776 2900 2784
rect 5644 2776 5652 2784
rect 5884 2776 5892 2784
rect 6124 2776 6132 2784
rect 6364 2776 6372 2784
rect 6412 2776 6420 2784
rect 620 2736 628 2744
rect 732 2736 740 2744
rect 844 2736 852 2744
rect 1260 2756 1268 2764
rect 2108 2756 2116 2764
rect 892 2736 900 2744
rect 2620 2736 2628 2744
rect 4092 2736 4100 2744
rect 5452 2736 5460 2744
rect 6076 2736 6084 2744
rect 124 2716 132 2724
rect 252 2716 260 2724
rect 364 2716 372 2724
rect 524 2716 532 2724
rect 700 2716 708 2724
rect 876 2716 884 2724
rect 924 2716 932 2724
rect 1036 2716 1044 2724
rect 1180 2716 1188 2724
rect 1244 2716 1252 2724
rect 1292 2716 1300 2724
rect 1836 2716 1844 2724
rect 1916 2716 1924 2724
rect 2076 2716 2084 2724
rect 2188 2716 2196 2724
rect 2588 2716 2596 2724
rect 3004 2716 3012 2724
rect 3036 2716 3044 2724
rect 3116 2716 3124 2724
rect 172 2696 180 2704
rect 300 2696 308 2704
rect 396 2696 404 2704
rect 476 2696 484 2704
rect 492 2696 500 2704
rect 524 2696 532 2704
rect 588 2696 596 2704
rect 636 2696 644 2704
rect 684 2696 692 2704
rect 716 2696 724 2704
rect 764 2696 772 2704
rect 796 2696 804 2704
rect 860 2696 868 2704
rect 972 2696 980 2704
rect 1068 2696 1076 2704
rect 1116 2696 1124 2704
rect 1212 2696 1220 2704
rect 1324 2696 1332 2704
rect 1564 2696 1572 2704
rect 1628 2694 1636 2702
rect 1756 2696 1764 2704
rect 1980 2696 1988 2704
rect 2092 2696 2100 2704
rect 2156 2696 2164 2704
rect 2300 2696 2308 2704
rect 2460 2696 2468 2704
rect 2524 2694 2532 2702
rect 2636 2696 2644 2704
rect 2764 2696 2772 2704
rect 2796 2696 2804 2704
rect 2828 2696 2836 2704
rect 2924 2696 2932 2704
rect 3036 2696 3044 2704
rect 3052 2696 3060 2704
rect 3100 2696 3108 2704
rect 12 2676 20 2684
rect 172 2676 180 2684
rect 188 2676 196 2684
rect 220 2676 228 2684
rect 284 2676 292 2684
rect 316 2676 324 2684
rect 476 2676 484 2684
rect 572 2676 580 2684
rect 780 2676 788 2684
rect 892 2676 900 2684
rect 988 2676 996 2684
rect 1020 2676 1028 2684
rect 1084 2676 1092 2684
rect 1196 2676 1204 2684
rect 1276 2676 1284 2684
rect 1340 2676 1348 2684
rect 1372 2676 1380 2684
rect 1388 2676 1396 2684
rect 1484 2676 1492 2684
rect 1692 2676 1700 2684
rect 1724 2676 1732 2684
rect 1868 2676 1876 2684
rect 1948 2676 1956 2684
rect 2028 2676 2036 2684
rect 2140 2676 2148 2684
rect 2188 2676 2196 2684
rect 2636 2676 2644 2684
rect 2748 2676 2756 2684
rect 2780 2676 2788 2684
rect 2812 2676 2820 2684
rect 3052 2676 3060 2684
rect 3068 2676 3076 2684
rect 3132 2676 3140 2684
rect 3148 2680 3156 2688
rect 3212 2696 3220 2704
rect 3260 2716 3268 2724
rect 4300 2716 4308 2724
rect 4348 2716 4356 2724
rect 4444 2716 4452 2724
rect 4476 2716 4484 2724
rect 4540 2716 4548 2724
rect 4924 2716 4932 2724
rect 3260 2696 3268 2704
rect 3276 2696 3284 2704
rect 3564 2696 3572 2704
rect 3692 2694 3700 2702
rect 3836 2696 3844 2704
rect 3964 2696 3972 2704
rect 4124 2696 4132 2704
rect 4156 2696 4164 2704
rect 4204 2696 4212 2704
rect 3244 2676 3252 2684
rect 3308 2676 3316 2684
rect 3404 2676 3412 2684
rect 3612 2676 3620 2684
rect 3756 2676 3764 2684
rect 3916 2676 3924 2684
rect 4124 2676 4132 2684
rect 252 2656 260 2664
rect 348 2656 356 2664
rect 428 2656 436 2664
rect 540 2656 548 2664
rect 668 2656 676 2664
rect 684 2656 692 2664
rect 812 2656 820 2664
rect 1004 2656 1012 2664
rect 1036 2656 1044 2664
rect 1164 2656 1172 2664
rect 1692 2656 1700 2664
rect 1788 2656 1796 2664
rect 1996 2656 2004 2664
rect 2124 2656 2132 2664
rect 2332 2656 2340 2664
rect 2828 2656 2836 2664
rect 2860 2656 2868 2664
rect 3388 2656 3396 2664
rect 3692 2656 3700 2664
rect 4092 2656 4100 2664
rect 4156 2656 4164 2664
rect 4172 2656 4180 2664
rect 4236 2656 4244 2664
rect 4268 2676 4276 2684
rect 4316 2676 4324 2684
rect 4364 2680 4372 2688
rect 4476 2696 4484 2704
rect 4588 2696 4596 2704
rect 4620 2696 4628 2704
rect 4716 2694 4724 2702
rect 4780 2696 4788 2704
rect 4940 2696 4948 2704
rect 4956 2696 4964 2704
rect 4988 2696 4996 2704
rect 5068 2696 5076 2704
rect 5132 2694 5140 2702
rect 5196 2696 5204 2704
rect 5324 2694 5332 2702
rect 5388 2696 5396 2704
rect 5516 2694 5524 2702
rect 5708 2694 5716 2702
rect 5852 2696 5860 2704
rect 5948 2694 5956 2702
rect 6092 2696 6100 2704
rect 6140 2696 6148 2704
rect 6236 2694 6244 2702
rect 6380 2696 6388 2704
rect 6492 2696 6500 2704
rect 4428 2676 4436 2684
rect 4492 2676 4500 2684
rect 4508 2676 4516 2684
rect 4572 2676 4580 2684
rect 5100 2676 5108 2684
rect 5292 2676 5300 2684
rect 5484 2676 5492 2684
rect 5740 2676 5748 2684
rect 6012 2676 6020 2684
rect 6172 2676 6180 2684
rect 6204 2676 6212 2684
rect 6284 2676 6292 2684
rect 6444 2676 6452 2684
rect 4316 2656 4324 2664
rect 4652 2656 4660 2664
rect 4908 2656 4916 2664
rect 4988 2656 4996 2664
rect 5036 2656 5044 2664
rect 5068 2656 5076 2664
rect 5948 2656 5956 2664
rect 140 2636 148 2644
rect 204 2636 212 2644
rect 332 2636 340 2644
rect 1500 2636 1508 2644
rect 1916 2636 1924 2644
rect 2076 2636 2084 2644
rect 2204 2636 2212 2644
rect 2396 2636 2404 2644
rect 2700 2636 2708 2644
rect 2972 2636 2980 2644
rect 3436 2636 3444 2644
rect 3452 2636 3460 2644
rect 3820 2636 3828 2644
rect 3868 2636 3876 2644
rect 4140 2636 4148 2644
rect 4396 2636 4404 2644
rect 4844 2636 4852 2644
rect 4972 2636 4980 2644
rect 5260 2636 5268 2644
rect 5836 2636 5844 2644
rect 6620 2636 6628 2644
rect 3310 2606 3318 2614
rect 3324 2606 3332 2614
rect 3338 2606 3346 2614
rect 6060 2596 6068 2604
rect 6172 2596 6180 2604
rect 28 2576 36 2584
rect 588 2576 596 2584
rect 620 2576 628 2584
rect 668 2576 676 2584
rect 716 2576 724 2584
rect 1116 2576 1124 2584
rect 1164 2576 1172 2584
rect 1212 2576 1220 2584
rect 1308 2576 1316 2584
rect 1372 2576 1380 2584
rect 1404 2576 1412 2584
rect 1436 2576 1444 2584
rect 1628 2576 1636 2584
rect 1868 2576 1876 2584
rect 2172 2576 2180 2584
rect 2236 2576 2244 2584
rect 2428 2576 2436 2584
rect 2476 2576 2484 2584
rect 2668 2576 2676 2584
rect 2972 2576 2980 2584
rect 3516 2576 3524 2584
rect 3532 2576 3540 2584
rect 3852 2576 3860 2584
rect 4220 2576 4228 2584
rect 4492 2576 4500 2584
rect 5324 2576 5332 2584
rect 5836 2576 5844 2584
rect 6028 2576 6036 2584
rect 6108 2576 6116 2584
rect 6604 2576 6612 2584
rect 76 2556 84 2564
rect 316 2556 324 2564
rect 364 2556 372 2564
rect 12 2536 20 2544
rect 108 2536 116 2544
rect 204 2536 212 2544
rect 236 2536 244 2544
rect 268 2536 276 2544
rect 300 2536 308 2544
rect 796 2556 804 2564
rect 828 2556 836 2564
rect 1004 2556 1012 2564
rect 1084 2556 1092 2564
rect 1196 2556 1204 2564
rect 1276 2556 1284 2564
rect 1324 2556 1332 2564
rect 444 2536 452 2544
rect 476 2536 484 2544
rect 540 2536 548 2544
rect 108 2516 116 2524
rect 188 2516 196 2524
rect 204 2516 212 2524
rect 284 2516 292 2524
rect 396 2516 404 2524
rect 428 2516 436 2524
rect 524 2516 532 2524
rect 652 2536 660 2544
rect 732 2536 740 2544
rect 812 2536 820 2544
rect 860 2536 868 2544
rect 956 2536 964 2544
rect 988 2536 996 2544
rect 1340 2536 1348 2544
rect 1372 2536 1380 2544
rect 1564 2556 1572 2564
rect 1692 2556 1700 2564
rect 2188 2556 2196 2564
rect 2492 2556 2500 2564
rect 2540 2556 2548 2564
rect 2588 2556 2596 2564
rect 2620 2556 2628 2564
rect 2684 2556 2692 2564
rect 1852 2536 1860 2544
rect 2028 2536 2036 2544
rect 2108 2536 2116 2544
rect 2124 2536 2132 2544
rect 2204 2536 2212 2544
rect 2236 2536 2244 2544
rect 2332 2536 2340 2544
rect 2444 2536 2452 2544
rect 2620 2536 2628 2544
rect 2684 2536 2692 2544
rect 2796 2556 2804 2564
rect 2844 2556 2852 2564
rect 3068 2556 3076 2564
rect 3660 2556 3668 2564
rect 4012 2556 4020 2564
rect 4076 2556 4084 2564
rect 4140 2556 4148 2564
rect 4236 2556 4244 2564
rect 4332 2556 4340 2564
rect 4348 2556 4356 2564
rect 4364 2556 4372 2564
rect 2748 2536 2756 2544
rect 2828 2536 2836 2544
rect 2876 2536 2884 2544
rect 2956 2536 2964 2544
rect 2988 2536 2996 2544
rect 3116 2536 3124 2544
rect 3164 2536 3172 2544
rect 732 2516 740 2524
rect 844 2516 852 2524
rect 972 2516 980 2524
rect 1036 2516 1044 2524
rect 1052 2516 1060 2524
rect 44 2496 52 2504
rect 76 2496 84 2504
rect 236 2496 244 2504
rect 332 2496 340 2504
rect 492 2496 500 2504
rect 588 2496 596 2504
rect 604 2496 612 2504
rect 684 2496 692 2504
rect 700 2496 708 2504
rect 844 2496 852 2504
rect 1132 2516 1140 2524
rect 1228 2516 1236 2524
rect 1292 2516 1300 2524
rect 1420 2516 1428 2524
rect 1564 2518 1572 2526
rect 1708 2516 1716 2524
rect 1756 2518 1764 2526
rect 1996 2518 2004 2526
rect 2060 2516 2068 2524
rect 2316 2516 2324 2524
rect 2524 2516 2532 2524
rect 2636 2516 2644 2524
rect 2652 2516 2660 2524
rect 2732 2516 2740 2524
rect 2796 2516 2804 2524
rect 2828 2516 2836 2524
rect 2860 2516 2868 2524
rect 2892 2516 2900 2524
rect 2940 2516 2948 2524
rect 3052 2516 3060 2524
rect 3084 2516 3092 2524
rect 3100 2516 3108 2524
rect 3132 2516 3140 2524
rect 3164 2516 3172 2524
rect 3244 2536 3252 2544
rect 3324 2536 3332 2544
rect 3564 2536 3572 2544
rect 3628 2536 3636 2544
rect 3692 2536 3700 2544
rect 3884 2536 3892 2544
rect 3916 2536 3924 2544
rect 3996 2536 4004 2544
rect 4076 2536 4084 2544
rect 4108 2536 4116 2544
rect 4172 2536 4180 2544
rect 4300 2536 4308 2544
rect 4348 2536 4356 2544
rect 4396 2536 4404 2544
rect 4444 2556 4452 2564
rect 4508 2556 4516 2564
rect 4748 2556 4756 2564
rect 5132 2556 5140 2564
rect 5196 2556 5204 2564
rect 5276 2556 5284 2564
rect 5308 2556 5316 2564
rect 6172 2556 6180 2564
rect 4444 2536 4452 2544
rect 3196 2516 3204 2524
rect 3388 2518 3396 2526
rect 1372 2496 1380 2504
rect 2156 2496 2164 2504
rect 2236 2496 2244 2504
rect 2476 2496 2484 2504
rect 2556 2496 2564 2504
rect 2780 2496 2788 2504
rect 2908 2496 2916 2504
rect 3020 2496 3028 2504
rect 3164 2496 3172 2504
rect 3452 2516 3460 2524
rect 3596 2516 3604 2524
rect 3724 2518 3732 2526
rect 3868 2516 3876 2524
rect 3932 2516 3940 2524
rect 3980 2516 3988 2524
rect 4044 2516 4052 2524
rect 4060 2516 4068 2524
rect 4204 2516 4212 2524
rect 4236 2516 4244 2524
rect 4284 2516 4292 2524
rect 4396 2516 4404 2524
rect 4444 2516 4452 2524
rect 4476 2536 4484 2544
rect 4524 2536 4532 2544
rect 4588 2536 4596 2544
rect 4652 2536 4660 2544
rect 4700 2536 4708 2544
rect 4764 2536 4772 2544
rect 4924 2536 4932 2544
rect 4956 2536 4964 2544
rect 4524 2516 4532 2524
rect 4604 2516 4612 2524
rect 4716 2516 4724 2524
rect 4780 2516 4788 2524
rect 4796 2516 4804 2524
rect 5116 2536 5124 2544
rect 5164 2536 5172 2544
rect 5180 2536 5188 2544
rect 5388 2536 5396 2544
rect 5484 2536 5492 2544
rect 5516 2536 5524 2544
rect 5644 2536 5652 2544
rect 5676 2536 5684 2544
rect 5868 2536 5876 2544
rect 5948 2536 5956 2544
rect 6108 2536 6116 2544
rect 6284 2556 6292 2564
rect 6444 2536 6452 2544
rect 3244 2496 3252 2504
rect 3532 2496 3540 2504
rect 3580 2496 3588 2504
rect 3948 2496 3956 2504
rect 4012 2496 4020 2504
rect 4572 2496 4580 2504
rect 4604 2496 4612 2504
rect 4636 2496 4644 2504
rect 4652 2496 4660 2504
rect 5196 2516 5204 2524
rect 5292 2516 5300 2524
rect 5420 2516 5428 2524
rect 5708 2518 5716 2526
rect 5900 2518 5908 2526
rect 6140 2516 6148 2524
rect 6204 2516 6212 2524
rect 6220 2516 6228 2524
rect 6284 2518 6292 2526
rect 6476 2518 6484 2526
rect 4876 2496 4884 2504
rect 4908 2496 4916 2504
rect 5084 2496 5092 2504
rect 6060 2496 6068 2504
rect 124 2476 132 2484
rect 2748 2476 2756 2484
rect 4540 2456 4548 2464
rect 5132 2456 5140 2464
rect 60 2436 68 2444
rect 188 2436 196 2444
rect 524 2436 532 2444
rect 1260 2436 1268 2444
rect 2140 2436 2148 2444
rect 2508 2436 2516 2444
rect 2940 2436 2948 2444
rect 3916 2436 3924 2444
rect 3980 2436 3988 2444
rect 4716 2436 4724 2444
rect 5004 2436 5012 2444
rect 6044 2436 6052 2444
rect 6412 2436 6420 2444
rect 1774 2406 1782 2414
rect 1788 2406 1796 2414
rect 1802 2406 1810 2414
rect 4830 2406 4838 2414
rect 4844 2406 4852 2414
rect 4858 2406 4866 2414
rect 252 2376 260 2384
rect 300 2376 308 2384
rect 364 2376 372 2384
rect 684 2376 692 2384
rect 1148 2376 1156 2384
rect 1516 2376 1524 2384
rect 4188 2376 4196 2384
rect 4252 2376 4260 2384
rect 4492 2376 4500 2384
rect 5100 2376 5108 2384
rect 5564 2376 5572 2384
rect 5900 2376 5908 2384
rect 172 2356 180 2364
rect 5452 2356 5460 2364
rect 188 2336 196 2344
rect 236 2336 244 2344
rect 316 2336 324 2344
rect 348 2336 356 2344
rect 380 2336 388 2344
rect 444 2336 452 2344
rect 492 2336 500 2344
rect 1820 2336 1828 2344
rect 2892 2336 2900 2344
rect 3372 2336 3380 2344
rect 5292 2336 5300 2344
rect 5436 2336 5444 2344
rect 5868 2336 5876 2344
rect 12 2316 20 2324
rect 156 2316 164 2324
rect 284 2316 292 2324
rect 348 2316 356 2324
rect 412 2316 420 2324
rect 524 2316 532 2324
rect 604 2316 612 2324
rect 700 2316 708 2324
rect 844 2316 852 2324
rect 924 2316 932 2324
rect 1020 2316 1028 2324
rect 1036 2316 1044 2324
rect 1116 2316 1124 2324
rect 1212 2316 1220 2324
rect 172 2296 180 2304
rect 252 2296 260 2304
rect 300 2296 308 2304
rect 364 2296 372 2304
rect 492 2296 500 2304
rect 524 2296 532 2304
rect 572 2296 580 2304
rect 636 2296 644 2304
rect 972 2296 980 2304
rect 1068 2296 1076 2304
rect 1100 2296 1108 2304
rect 1180 2296 1188 2304
rect 1260 2316 1268 2324
rect 1436 2316 1444 2324
rect 1596 2316 1604 2324
rect 1644 2316 1652 2324
rect 1724 2316 1732 2324
rect 2028 2316 2036 2324
rect 2060 2316 2068 2324
rect 2156 2316 2164 2324
rect 2444 2316 2452 2324
rect 1340 2296 1348 2304
rect 1404 2296 1412 2304
rect 1436 2296 1444 2304
rect 1852 2296 1860 2304
rect 1916 2294 1924 2302
rect 2252 2296 2260 2304
rect 2300 2294 2308 2302
rect 2428 2296 2436 2304
rect 2476 2296 2484 2304
rect 2524 2316 2532 2324
rect 2604 2316 2612 2324
rect 2732 2316 2740 2324
rect 2876 2316 2884 2324
rect 2924 2316 2932 2324
rect 3132 2316 3140 2324
rect 3292 2316 3300 2324
rect 3404 2316 3412 2324
rect 3532 2316 3540 2324
rect 4092 2316 4100 2324
rect 4284 2316 4292 2324
rect 4556 2316 4564 2324
rect 2652 2296 2660 2304
rect 2684 2296 2692 2304
rect 2716 2296 2724 2304
rect 3004 2296 3012 2304
rect 3020 2296 3028 2304
rect 3100 2296 3108 2304
rect 3148 2296 3156 2304
rect 3196 2296 3204 2304
rect 3356 2296 3364 2304
rect 3484 2296 3492 2304
rect 3612 2296 3620 2304
rect 3676 2294 3684 2302
rect 3820 2296 3828 2304
rect 3964 2296 3972 2304
rect 3996 2296 4004 2304
rect 44 2276 52 2284
rect 124 2276 132 2284
rect 460 2276 468 2284
rect 588 2276 596 2284
rect 604 2276 612 2284
rect 652 2276 660 2284
rect 764 2276 772 2284
rect 812 2276 820 2284
rect 876 2276 884 2284
rect 892 2276 900 2284
rect 972 2276 980 2284
rect 1068 2276 1076 2284
rect 1132 2276 1140 2284
rect 1164 2276 1172 2284
rect 1324 2276 1332 2284
rect 1500 2276 1508 2284
rect 1532 2276 1540 2284
rect 1580 2276 1588 2284
rect 1676 2276 1684 2284
rect 2012 2276 2020 2284
rect 2108 2276 2116 2284
rect 2332 2276 2340 2284
rect 2396 2276 2404 2284
rect 2460 2276 2468 2284
rect 2492 2276 2500 2284
rect 2556 2276 2564 2284
rect 2572 2276 2580 2284
rect 2636 2276 2644 2284
rect 2780 2276 2788 2284
rect 2828 2276 2836 2284
rect 2956 2276 2964 2284
rect 3084 2276 3092 2284
rect 3116 2276 3124 2284
rect 3212 2276 3220 2284
rect 3260 2276 3268 2284
rect 3356 2276 3364 2284
rect 3484 2276 3492 2284
rect 3500 2276 3508 2284
rect 3772 2280 3780 2288
rect 3788 2276 3796 2284
rect 4140 2296 4148 2304
rect 4252 2296 4260 2304
rect 4300 2296 4308 2304
rect 4332 2296 4340 2304
rect 4412 2296 4420 2304
rect 4476 2296 4484 2304
rect 4524 2296 4532 2304
rect 4588 2296 4596 2304
rect 4636 2316 4644 2324
rect 5148 2316 5156 2324
rect 4732 2294 4740 2302
rect 4796 2296 4804 2304
rect 4972 2294 4980 2302
rect 5036 2296 5044 2304
rect 5164 2296 5172 2304
rect 5228 2296 5236 2304
rect 5340 2316 5348 2324
rect 5468 2316 5476 2324
rect 5516 2316 5524 2324
rect 5948 2316 5956 2324
rect 6028 2316 6036 2324
rect 6092 2316 6100 2324
rect 6156 2316 6164 2324
rect 5404 2296 5412 2304
rect 5452 2296 5460 2304
rect 5532 2296 5540 2304
rect 5772 2294 5780 2302
rect 6012 2296 6020 2304
rect 6108 2296 6116 2304
rect 6188 2296 6196 2304
rect 6268 2294 6276 2302
rect 6508 2296 6516 2304
rect 4236 2276 4244 2284
rect 4316 2276 4324 2284
rect 4396 2276 4404 2284
rect 4636 2276 4644 2284
rect 4668 2276 4676 2284
rect 4700 2276 4708 2284
rect 4876 2276 4884 2284
rect 5116 2276 5124 2284
rect 5180 2276 5188 2284
rect 5212 2276 5220 2284
rect 668 2256 676 2264
rect 716 2256 724 2264
rect 828 2256 836 2264
rect 940 2256 948 2264
rect 956 2256 964 2264
rect 1052 2256 1060 2264
rect 1228 2256 1236 2264
rect 1340 2256 1348 2264
rect 1372 2256 1380 2264
rect 1468 2256 1476 2264
rect 1484 2256 1492 2264
rect 1548 2256 1556 2264
rect 1644 2256 1652 2264
rect 1980 2256 1988 2264
rect 2076 2256 2084 2264
rect 2364 2256 2372 2264
rect 2716 2256 2724 2264
rect 2812 2256 2820 2264
rect 2892 2256 2900 2264
rect 2972 2256 2980 2264
rect 3068 2256 3076 2264
rect 3180 2256 3188 2264
rect 3244 2256 3252 2264
rect 3420 2256 3428 2264
rect 3436 2256 3444 2264
rect 3452 2256 3460 2264
rect 3532 2256 3540 2264
rect 3804 2256 3812 2264
rect 3836 2256 3844 2264
rect 3916 2256 3924 2264
rect 3948 2256 3956 2264
rect 3964 2256 3972 2264
rect 4044 2256 4052 2264
rect 4108 2256 4116 2264
rect 4220 2256 4228 2264
rect 4348 2256 4356 2264
rect 4364 2256 4372 2264
rect 4460 2256 4468 2264
rect 5276 2276 5284 2284
rect 5372 2276 5380 2284
rect 5484 2276 5492 2284
rect 5580 2276 5588 2284
rect 5708 2276 5716 2284
rect 5740 2276 5748 2284
rect 5916 2276 5924 2284
rect 5948 2276 5956 2284
rect 6092 2276 6100 2284
rect 6172 2276 6180 2284
rect 6204 2276 6212 2284
rect 6236 2276 6244 2284
rect 6428 2276 6436 2284
rect 5388 2256 5396 2264
rect 6140 2256 6148 2264
rect 12 2236 20 2244
rect 108 2236 116 2244
rect 732 2236 740 2244
rect 780 2236 788 2244
rect 844 2236 852 2244
rect 908 2236 916 2244
rect 1004 2236 1012 2244
rect 1148 2236 1156 2244
rect 1436 2236 1444 2244
rect 1516 2236 1524 2244
rect 1772 2236 1780 2244
rect 1788 2236 1796 2244
rect 2156 2236 2164 2244
rect 2172 2236 2180 2244
rect 2876 2236 2884 2244
rect 2940 2236 2948 2244
rect 3052 2236 3060 2244
rect 3228 2236 3236 2244
rect 3548 2236 3556 2244
rect 3740 2236 3748 2244
rect 3852 2236 3860 2244
rect 4028 2236 4036 2244
rect 4380 2236 4388 2244
rect 4860 2236 4868 2244
rect 5148 2236 5156 2244
rect 5180 2236 5188 2244
rect 5516 2236 5524 2244
rect 5948 2236 5956 2244
rect 6076 2236 6084 2244
rect 6396 2236 6404 2244
rect 6588 2236 6596 2244
rect 3310 2206 3318 2214
rect 3324 2206 3332 2214
rect 3338 2206 3346 2214
rect 5964 2196 5972 2204
rect 108 2176 116 2184
rect 364 2176 372 2184
rect 412 2176 420 2184
rect 508 2176 516 2184
rect 860 2176 868 2184
rect 1004 2176 1012 2184
rect 1388 2176 1396 2184
rect 1420 2176 1428 2184
rect 1468 2176 1476 2184
rect 1660 2176 1668 2184
rect 1900 2176 1908 2184
rect 2092 2176 2100 2184
rect 2572 2176 2580 2184
rect 2764 2176 2772 2184
rect 2924 2176 2932 2184
rect 3164 2176 3172 2184
rect 3212 2176 3220 2184
rect 3276 2176 3284 2184
rect 3388 2176 3396 2184
rect 3420 2176 3428 2184
rect 3964 2176 3972 2184
rect 4268 2176 4276 2184
rect 4732 2176 4740 2184
rect 5388 2176 5396 2184
rect 5820 2176 5828 2184
rect 5868 2176 5876 2184
rect 5916 2176 5924 2184
rect 5932 2176 5940 2184
rect 6044 2176 6052 2184
rect 6108 2176 6116 2184
rect 124 2156 132 2164
rect 188 2156 196 2164
rect 588 2156 596 2164
rect 716 2156 724 2164
rect 844 2156 852 2164
rect 956 2156 964 2164
rect 1132 2156 1140 2164
rect 2780 2156 2788 2164
rect 2812 2156 2820 2164
rect 2860 2156 2868 2164
rect 2908 2156 2916 2164
rect 2940 2156 2948 2164
rect 2972 2156 2980 2164
rect 2988 2156 2996 2164
rect 3036 2156 3044 2164
rect 3132 2156 3140 2164
rect 3148 2156 3156 2164
rect 3260 2156 3268 2164
rect 3372 2156 3380 2164
rect 4252 2156 4260 2164
rect 5228 2156 5236 2164
rect 5340 2156 5348 2164
rect 5372 2156 5380 2164
rect 6060 2156 6068 2164
rect 6156 2156 6164 2164
rect 6236 2156 6244 2164
rect 6300 2156 6308 2164
rect 6380 2156 6388 2164
rect 6460 2156 6468 2164
rect 6492 2156 6500 2164
rect 92 2136 100 2144
rect 156 2136 164 2144
rect 252 2136 260 2144
rect 332 2136 340 2144
rect 396 2136 404 2144
rect 428 2136 436 2144
rect 476 2136 484 2144
rect 572 2136 580 2144
rect 636 2136 644 2144
rect 684 2136 692 2144
rect 700 2136 708 2144
rect 828 2136 836 2144
rect 44 2116 52 2124
rect 76 2116 84 2124
rect 140 2116 148 2124
rect 220 2116 228 2124
rect 284 2116 292 2124
rect 380 2116 388 2124
rect 444 2116 452 2124
rect 460 2116 468 2124
rect 524 2116 532 2124
rect 604 2116 612 2124
rect 748 2116 756 2124
rect 988 2136 996 2144
rect 1100 2136 1108 2144
rect 1180 2136 1188 2144
rect 1244 2136 1252 2144
rect 1452 2136 1460 2144
rect 1628 2136 1636 2144
rect 1820 2136 1828 2144
rect 2204 2136 2212 2144
rect 2252 2136 2260 2144
rect 2284 2136 2292 2144
rect 2316 2136 2324 2144
rect 2380 2136 2388 2144
rect 2460 2136 2468 2144
rect 2604 2136 2612 2144
rect 2780 2136 2788 2144
rect 3036 2136 3044 2144
rect 3100 2136 3108 2144
rect 3180 2136 3188 2144
rect 3244 2136 3252 2144
rect 3580 2136 3588 2144
rect 3612 2136 3620 2144
rect 3660 2136 3668 2144
rect 3708 2136 3716 2144
rect 3772 2136 3780 2144
rect 4028 2136 4036 2144
rect 4188 2136 4196 2144
rect 4252 2136 4260 2144
rect 4300 2136 4308 2144
rect 4316 2136 4324 2144
rect 4444 2136 4452 2144
rect 4508 2136 4516 2144
rect 4540 2136 4548 2144
rect 4572 2136 4580 2144
rect 4780 2136 4788 2144
rect 4812 2136 4820 2144
rect 4828 2136 4836 2144
rect 4908 2136 4916 2144
rect 4924 2136 4932 2144
rect 5020 2136 5028 2144
rect 5036 2136 5044 2144
rect 5132 2136 5140 2144
rect 5148 2136 5156 2144
rect 5212 2136 5220 2144
rect 5308 2136 5316 2144
rect 5420 2136 5428 2144
rect 5500 2136 5508 2144
rect 5596 2136 5604 2144
rect 5628 2136 5636 2144
rect 5708 2136 5716 2144
rect 5852 2136 5860 2144
rect 5916 2136 5924 2144
rect 6044 2136 6052 2144
rect 6268 2136 6276 2144
rect 6332 2136 6340 2144
rect 6572 2136 6580 2144
rect 892 2116 900 2124
rect 1068 2116 1076 2124
rect 1084 2116 1092 2124
rect 1164 2116 1172 2124
rect 1196 2116 1204 2124
rect 1260 2116 1268 2124
rect 1292 2116 1300 2124
rect 1324 2116 1332 2124
rect 1596 2118 1604 2126
rect 1772 2116 1780 2124
rect 1964 2116 1972 2124
rect 2028 2118 2036 2126
rect 2220 2118 2228 2126
rect 60 2096 68 2104
rect 268 2096 276 2104
rect 332 2096 340 2104
rect 364 2096 372 2104
rect 604 2096 612 2104
rect 652 2096 660 2104
rect 796 2096 804 2104
rect 812 2096 820 2104
rect 1036 2096 1044 2104
rect 1228 2096 1236 2104
rect 1292 2096 1300 2104
rect 1308 2096 1316 2104
rect 1404 2096 1412 2104
rect 1420 2096 1428 2104
rect 2316 2096 2324 2104
rect 2364 2116 2372 2124
rect 2492 2116 2500 2124
rect 2652 2116 2660 2124
rect 2812 2116 2820 2124
rect 2892 2116 2900 2124
rect 2940 2116 2948 2124
rect 3020 2116 3028 2124
rect 3068 2116 3076 2124
rect 3084 2116 3092 2124
rect 3308 2116 3316 2124
rect 3404 2116 3412 2124
rect 3548 2118 3556 2126
rect 2540 2096 2548 2104
rect 3212 2096 3220 2104
rect 3644 2096 3652 2104
rect 3756 2116 3764 2124
rect 3852 2116 3860 2124
rect 3884 2116 3892 2124
rect 4028 2116 4036 2124
rect 4044 2116 4052 2124
rect 4364 2116 4372 2124
rect 4460 2116 4468 2124
rect 4604 2118 4612 2126
rect 3724 2096 3732 2104
rect 4012 2096 4020 2104
rect 4076 2096 4084 2104
rect 4204 2096 4212 2104
rect 4668 2116 4676 2124
rect 5164 2116 5172 2124
rect 5196 2116 5204 2124
rect 5260 2116 5268 2124
rect 5292 2116 5300 2124
rect 5452 2116 5460 2124
rect 5548 2116 5556 2124
rect 5596 2116 5604 2124
rect 5660 2116 5668 2124
rect 5868 2116 5876 2124
rect 5916 2116 5924 2124
rect 5948 2116 5956 2124
rect 6060 2116 6068 2124
rect 6188 2116 6196 2124
rect 6284 2116 6292 2124
rect 6332 2116 6340 2124
rect 6412 2116 6420 2124
rect 6460 2116 6468 2124
rect 6524 2116 6532 2124
rect 4508 2096 4516 2104
rect 4796 2096 4804 2104
rect 5372 2096 5380 2104
rect 5484 2096 5492 2104
rect 5580 2096 5588 2104
rect 5628 2096 5636 2104
rect 5900 2096 5908 2104
rect 5996 2096 6004 2104
rect 6012 2096 6020 2104
rect 6172 2096 6180 2104
rect 6316 2096 6324 2104
rect 6396 2096 6404 2104
rect 6444 2096 6452 2104
rect 6556 2096 6564 2104
rect 28 2076 36 2084
rect 236 2076 244 2084
rect 300 2076 308 2084
rect 764 2076 772 2084
rect 1196 2076 1204 2084
rect 1340 2076 1348 2084
rect 5372 2076 5380 2084
rect 6204 2076 6212 2084
rect 6412 2076 6420 2084
rect 6428 2076 6436 2084
rect 44 2056 52 2064
rect 540 2036 548 2044
rect 668 2036 676 2044
rect 780 2036 788 2044
rect 1116 2036 1124 2044
rect 1148 2036 1156 2044
rect 1324 2036 1332 2044
rect 1660 2036 1668 2044
rect 1900 2036 1908 2044
rect 2876 2036 2884 2044
rect 3052 2036 3060 2044
rect 3132 2036 3140 2044
rect 4124 2036 4132 2044
rect 4220 2036 4228 2044
rect 4764 2036 4772 2044
rect 4892 2036 4900 2044
rect 4956 2036 4964 2044
rect 5068 2036 5076 2044
rect 5164 2036 5172 2044
rect 5324 2036 5332 2044
rect 5452 2036 5460 2044
rect 5516 2036 5524 2044
rect 5612 2036 5620 2044
rect 5692 2036 5700 2044
rect 5932 2036 5940 2044
rect 5964 2036 5972 2044
rect 6028 2036 6036 2044
rect 6076 2036 6084 2044
rect 6188 2036 6196 2044
rect 6236 2036 6244 2044
rect 6460 2036 6468 2044
rect 6524 2036 6532 2044
rect 6588 2036 6596 2044
rect 1774 2006 1782 2014
rect 1788 2006 1796 2014
rect 1802 2006 1810 2014
rect 4830 2006 4838 2014
rect 4844 2006 4852 2014
rect 4858 2006 4866 2014
rect 28 1976 36 1984
rect 108 1976 116 1984
rect 156 1976 164 1984
rect 268 1976 276 1984
rect 348 1976 356 1984
rect 588 1976 596 1984
rect 668 1976 676 1984
rect 924 1976 932 1984
rect 1260 1976 1268 1984
rect 1276 1976 1284 1984
rect 2364 1976 2372 1984
rect 3068 1976 3076 1984
rect 3196 1976 3204 1984
rect 3948 1976 3956 1984
rect 4396 1976 4404 1984
rect 4588 1976 4596 1984
rect 6572 1976 6580 1984
rect 44 1936 52 1944
rect 92 1936 100 1944
rect 172 1936 180 1944
rect 236 1936 244 1944
rect 284 1936 292 1944
rect 364 1936 372 1944
rect 2556 1936 2564 1944
rect 2572 1936 2580 1944
rect 5020 1936 5028 1944
rect 5708 1936 5716 1944
rect 6476 1936 6484 1944
rect 12 1916 20 1924
rect 124 1916 132 1924
rect 204 1916 212 1924
rect 332 1916 340 1924
rect 460 1916 468 1924
rect 492 1916 500 1924
rect 524 1916 532 1924
rect 796 1916 804 1924
rect 812 1916 820 1924
rect 956 1916 964 1924
rect 1020 1916 1028 1924
rect 1308 1916 1316 1924
rect 1388 1916 1396 1924
rect 1532 1916 1540 1924
rect 1628 1916 1636 1924
rect 1836 1916 1844 1924
rect 1900 1916 1908 1924
rect 2044 1916 2052 1924
rect 3148 1916 3156 1924
rect 28 1896 36 1904
rect 108 1896 116 1904
rect 156 1896 164 1904
rect 220 1896 228 1904
rect 300 1896 308 1904
rect 348 1896 356 1904
rect 396 1896 404 1904
rect 492 1896 500 1904
rect 556 1896 564 1904
rect 636 1896 644 1904
rect 428 1876 436 1884
rect 508 1876 516 1884
rect 556 1876 564 1884
rect 588 1876 596 1884
rect 620 1876 628 1884
rect 716 1896 724 1904
rect 860 1896 868 1904
rect 908 1896 916 1904
rect 988 1896 996 1904
rect 1052 1896 1060 1904
rect 1116 1896 1124 1904
rect 1164 1896 1172 1904
rect 1196 1896 1204 1904
rect 1404 1896 1412 1904
rect 1452 1896 1460 1904
rect 1676 1896 1684 1904
rect 1740 1896 1748 1904
rect 1884 1896 1892 1904
rect 2108 1896 2116 1904
rect 2156 1896 2164 1904
rect 2252 1896 2260 1904
rect 2444 1896 2452 1904
rect 668 1876 676 1884
rect 700 1876 708 1884
rect 764 1876 772 1884
rect 876 1876 884 1884
rect 972 1876 980 1884
rect 1004 1876 1012 1884
rect 444 1856 452 1864
rect 732 1856 740 1864
rect 748 1856 756 1864
rect 1180 1876 1188 1884
rect 1228 1876 1236 1884
rect 1244 1876 1252 1884
rect 1340 1876 1348 1884
rect 1420 1876 1428 1884
rect 1564 1876 1572 1884
rect 1580 1876 1588 1884
rect 2700 1894 2708 1902
rect 2812 1896 2820 1904
rect 2956 1896 2964 1904
rect 3004 1896 3012 1904
rect 3052 1896 3060 1904
rect 3116 1896 3124 1904
rect 3692 1916 3700 1924
rect 4204 1916 4212 1924
rect 4684 1916 4692 1924
rect 4716 1916 4724 1924
rect 4796 1916 4804 1924
rect 4940 1916 4948 1924
rect 5052 1916 5060 1924
rect 5068 1916 5076 1924
rect 5180 1916 5188 1924
rect 3196 1896 3204 1904
rect 3260 1896 3268 1904
rect 3420 1896 3428 1904
rect 3548 1896 3556 1904
rect 3660 1896 3668 1904
rect 3756 1896 3764 1904
rect 3852 1896 3860 1904
rect 3884 1896 3892 1904
rect 3980 1896 3988 1904
rect 3996 1896 4004 1904
rect 4172 1896 4180 1904
rect 4268 1894 4276 1902
rect 4332 1896 4340 1904
rect 4460 1894 4468 1902
rect 4508 1896 4516 1904
rect 4636 1896 4644 1904
rect 4684 1896 4692 1904
rect 4892 1896 4900 1904
rect 4956 1896 4964 1904
rect 4972 1896 4980 1904
rect 4988 1896 4996 1904
rect 5260 1896 5268 1904
rect 5292 1896 5300 1904
rect 5324 1896 5332 1904
rect 5356 1896 5364 1904
rect 5404 1916 5412 1924
rect 5500 1916 5508 1924
rect 5516 1916 5524 1924
rect 5612 1916 5620 1924
rect 5740 1916 5748 1924
rect 5788 1916 5796 1924
rect 5932 1916 5940 1924
rect 6140 1916 6148 1924
rect 6460 1916 6468 1924
rect 6524 1916 6532 1924
rect 6540 1916 6548 1924
rect 6588 1916 6596 1924
rect 5468 1896 5476 1904
rect 5548 1896 5556 1904
rect 5804 1896 5812 1904
rect 5868 1896 5876 1904
rect 6012 1896 6020 1904
rect 6108 1896 6116 1904
rect 6220 1896 6228 1904
rect 6252 1896 6260 1904
rect 6300 1896 6308 1904
rect 6332 1896 6340 1904
rect 6380 1896 6388 1904
rect 6412 1896 6420 1904
rect 6460 1896 6468 1904
rect 1692 1876 1700 1884
rect 1724 1876 1732 1884
rect 1804 1876 1812 1884
rect 1900 1876 1908 1884
rect 1948 1876 1956 1884
rect 1996 1876 2004 1884
rect 2076 1876 2084 1884
rect 2172 1876 2180 1884
rect 2204 1876 2212 1884
rect 2252 1876 2260 1884
rect 2348 1876 2356 1884
rect 2444 1876 2452 1884
rect 2460 1876 2468 1884
rect 2732 1876 2740 1884
rect 2812 1876 2820 1884
rect 2908 1876 2916 1884
rect 892 1856 900 1864
rect 940 1856 948 1864
rect 1084 1856 1092 1864
rect 1292 1856 1300 1864
rect 1356 1856 1364 1864
rect 1452 1856 1460 1864
rect 1516 1856 1524 1864
rect 1964 1856 1972 1864
rect 2060 1856 2068 1864
rect 2764 1856 2772 1864
rect 2924 1856 2932 1864
rect 2956 1856 2964 1864
rect 2988 1856 2996 1864
rect 3036 1856 3044 1864
rect 3100 1876 3108 1884
rect 3212 1876 3220 1884
rect 3260 1876 3268 1884
rect 3324 1876 3332 1884
rect 3644 1876 3652 1884
rect 3708 1876 3716 1884
rect 3724 1880 3732 1888
rect 4028 1876 4036 1884
rect 4140 1876 4148 1884
rect 4156 1876 4164 1884
rect 4204 1876 4212 1884
rect 4652 1876 4660 1884
rect 4668 1876 4676 1884
rect 4764 1876 4772 1884
rect 4876 1876 4884 1884
rect 4988 1876 4996 1884
rect 5004 1876 5012 1884
rect 5100 1876 5108 1884
rect 5116 1876 5124 1884
rect 5340 1876 5348 1884
rect 5404 1876 5412 1884
rect 5436 1876 5444 1884
rect 5452 1876 5460 1884
rect 5532 1876 5540 1884
rect 5564 1876 5572 1884
rect 5644 1876 5652 1884
rect 5708 1876 5716 1884
rect 5740 1876 5748 1884
rect 5756 1876 5764 1884
rect 5820 1876 5828 1884
rect 5884 1876 5892 1884
rect 3228 1856 3236 1864
rect 3276 1856 3284 1864
rect 3340 1856 3348 1864
rect 3404 1856 3412 1864
rect 3436 1856 3444 1864
rect 3580 1856 3588 1864
rect 3692 1856 3700 1864
rect 3964 1856 3972 1864
rect 4028 1856 4036 1864
rect 4732 1856 4740 1864
rect 4892 1856 4900 1864
rect 4924 1856 4932 1864
rect 5084 1856 5092 1864
rect 5228 1856 5236 1864
rect 5260 1856 5268 1864
rect 5292 1856 5300 1864
rect 5676 1856 5684 1864
rect 5852 1856 5860 1864
rect 5996 1876 6004 1884
rect 6092 1876 6100 1884
rect 6156 1876 6164 1884
rect 6236 1876 6244 1884
rect 6268 1876 6276 1884
rect 6316 1876 6324 1884
rect 6348 1876 6356 1884
rect 6364 1876 6372 1884
rect 6396 1876 6404 1884
rect 6428 1876 6436 1884
rect 6508 1876 6516 1884
rect 6556 1876 6564 1884
rect 5932 1856 5940 1864
rect 6076 1856 6084 1864
rect 6188 1856 6196 1864
rect 252 1836 260 1844
rect 524 1836 532 1844
rect 588 1836 596 1844
rect 780 1836 788 1844
rect 812 1836 820 1844
rect 924 1836 932 1844
rect 1020 1836 1028 1844
rect 1132 1836 1140 1844
rect 1212 1836 1220 1844
rect 1260 1836 1268 1844
rect 1308 1836 1316 1844
rect 1532 1836 1540 1844
rect 1596 1836 1604 1844
rect 1628 1836 1636 1844
rect 1692 1836 1700 1844
rect 1820 1836 1828 1844
rect 1852 1836 1860 1844
rect 1916 1836 1924 1844
rect 2044 1836 2052 1844
rect 2124 1836 2132 1844
rect 2780 1836 2788 1844
rect 2876 1836 2884 1844
rect 3068 1836 3076 1844
rect 3452 1836 3460 1844
rect 3948 1836 3956 1844
rect 4076 1836 4084 1844
rect 4604 1836 4612 1844
rect 4748 1836 4756 1844
rect 4812 1836 4820 1844
rect 5276 1836 5284 1844
rect 5308 1836 5316 1844
rect 5404 1836 5412 1844
rect 5500 1836 5508 1844
rect 5612 1836 5620 1844
rect 5836 1836 5844 1844
rect 5980 1836 5988 1844
rect 6060 1836 6068 1844
rect 6460 1836 6468 1844
rect 6588 1836 6596 1844
rect 3310 1806 3318 1814
rect 3324 1806 3332 1814
rect 3338 1806 3346 1814
rect 172 1776 180 1784
rect 252 1776 260 1784
rect 364 1776 372 1784
rect 668 1776 676 1784
rect 1852 1776 1860 1784
rect 2220 1776 2228 1784
rect 2252 1776 2260 1784
rect 2684 1776 2692 1784
rect 3740 1776 3748 1784
rect 4508 1776 4516 1784
rect 5468 1776 5476 1784
rect 5548 1776 5556 1784
rect 5724 1776 5732 1784
rect 108 1756 116 1764
rect 300 1756 308 1764
rect 380 1756 388 1764
rect 428 1756 436 1764
rect 780 1756 788 1764
rect 1004 1756 1012 1764
rect 1212 1756 1220 1764
rect 1468 1756 1476 1764
rect 1516 1756 1524 1764
rect 3116 1756 3124 1764
rect 3164 1756 3172 1764
rect 3180 1756 3188 1764
rect 3196 1756 3204 1764
rect 3356 1756 3364 1764
rect 3436 1756 3444 1764
rect 3548 1756 3556 1764
rect 4220 1756 4228 1764
rect 4684 1756 4692 1764
rect 4892 1756 4900 1764
rect 5020 1756 5028 1764
rect 5116 1756 5124 1764
rect 5676 1756 5684 1764
rect 5772 1756 5780 1764
rect 5788 1756 5796 1764
rect 5900 1756 5908 1764
rect 5916 1756 5924 1764
rect 5932 1756 5940 1764
rect 6012 1756 6020 1764
rect 6300 1756 6308 1764
rect 6348 1756 6356 1764
rect 6364 1756 6372 1764
rect 6588 1756 6596 1764
rect 12 1736 20 1744
rect 44 1736 52 1744
rect 108 1736 116 1744
rect 188 1736 196 1744
rect 348 1736 356 1744
rect 508 1736 516 1744
rect 540 1736 548 1744
rect 556 1736 564 1744
rect 636 1736 644 1744
rect 124 1716 132 1724
rect 140 1716 148 1724
rect 172 1716 180 1724
rect 220 1716 228 1724
rect 268 1716 276 1724
rect 396 1716 404 1724
rect 460 1716 468 1724
rect 764 1736 772 1744
rect 908 1736 916 1744
rect 924 1736 932 1744
rect 956 1736 964 1744
rect 1052 1736 1060 1744
rect 1068 1736 1076 1744
rect 1324 1736 1332 1744
rect 44 1696 52 1704
rect 252 1696 260 1704
rect 316 1696 324 1704
rect 348 1696 356 1704
rect 444 1696 452 1704
rect 508 1696 516 1704
rect 572 1696 580 1704
rect 716 1716 724 1724
rect 828 1716 836 1724
rect 876 1716 884 1724
rect 892 1716 900 1724
rect 972 1716 980 1724
rect 1084 1716 1092 1724
rect 1148 1716 1156 1724
rect 1260 1716 1268 1724
rect 1372 1716 1380 1724
rect 1420 1716 1428 1724
rect 1532 1736 1540 1744
rect 1596 1736 1604 1744
rect 1628 1736 1636 1744
rect 1644 1736 1652 1744
rect 1740 1736 1748 1744
rect 1836 1736 1844 1744
rect 2364 1736 2372 1744
rect 2572 1736 2580 1744
rect 2604 1736 2612 1744
rect 2668 1736 2676 1744
rect 2748 1736 2756 1744
rect 2844 1736 2852 1744
rect 2876 1736 2884 1744
rect 2940 1736 2948 1744
rect 2972 1736 2980 1744
rect 3004 1736 3012 1744
rect 3100 1736 3108 1744
rect 3244 1736 3252 1744
rect 3580 1736 3588 1744
rect 3884 1736 3892 1744
rect 3900 1736 3908 1744
rect 3996 1736 4004 1744
rect 4012 1736 4020 1744
rect 4108 1736 4116 1744
rect 4156 1736 4164 1744
rect 4204 1736 4212 1744
rect 4236 1736 4244 1744
rect 4332 1736 4340 1744
rect 4348 1736 4356 1744
rect 4444 1736 4452 1744
rect 4476 1736 4484 1744
rect 4492 1736 4500 1744
rect 4604 1736 4612 1744
rect 4908 1736 4916 1744
rect 5004 1736 5012 1744
rect 1612 1716 1620 1724
rect 1980 1718 1988 1726
rect 2124 1716 2132 1724
rect 2156 1716 2164 1724
rect 2444 1716 2452 1724
rect 2508 1718 2516 1726
rect 604 1696 612 1704
rect 700 1696 708 1704
rect 844 1696 852 1704
rect 860 1696 868 1704
rect 956 1696 964 1704
rect 1020 1696 1028 1704
rect 1116 1696 1124 1704
rect 1132 1696 1140 1704
rect 1212 1696 1220 1704
rect 1276 1696 1284 1704
rect 1292 1696 1300 1704
rect 1404 1696 1412 1704
rect 1788 1696 1796 1704
rect 2604 1696 2612 1704
rect 2652 1716 2660 1724
rect 2812 1718 2820 1726
rect 2908 1716 2916 1724
rect 2988 1716 2996 1724
rect 3052 1716 3060 1724
rect 3132 1716 3140 1724
rect 3260 1716 3268 1724
rect 3356 1716 3364 1724
rect 3388 1716 3396 1724
rect 3452 1716 3460 1724
rect 3484 1716 3492 1724
rect 3516 1716 3524 1724
rect 3612 1718 3620 1726
rect 3676 1716 3684 1724
rect 3756 1716 3764 1724
rect 4332 1716 4340 1724
rect 4620 1716 4628 1724
rect 4652 1716 4660 1724
rect 4716 1716 4724 1724
rect 4796 1716 4804 1724
rect 4828 1716 4836 1724
rect 5212 1736 5220 1744
rect 5276 1736 5284 1744
rect 5292 1736 5300 1744
rect 5308 1736 5316 1744
rect 5324 1736 5332 1744
rect 5356 1732 5364 1740
rect 5404 1736 5412 1744
rect 5500 1736 5508 1744
rect 5516 1736 5524 1744
rect 5564 1736 5572 1744
rect 5660 1736 5668 1744
rect 5692 1736 5700 1744
rect 5740 1736 5748 1744
rect 5836 1736 5844 1744
rect 5980 1736 5988 1744
rect 6492 1736 6500 1744
rect 5148 1716 5156 1724
rect 5196 1716 5204 1724
rect 5244 1716 5252 1724
rect 5260 1716 5268 1724
rect 5804 1716 5812 1724
rect 5820 1716 5828 1724
rect 5852 1716 5860 1724
rect 5884 1716 5892 1724
rect 6012 1716 6020 1724
rect 6044 1716 6052 1724
rect 6108 1716 6116 1724
rect 6172 1716 6180 1724
rect 6236 1716 6244 1724
rect 6428 1716 6436 1724
rect 6540 1716 6548 1724
rect 2876 1696 2884 1704
rect 2940 1696 2948 1704
rect 2956 1696 2964 1704
rect 3292 1696 3300 1704
rect 4124 1696 4132 1704
rect 4524 1696 4532 1704
rect 4540 1696 4548 1704
rect 4652 1696 4660 1704
rect 4684 1696 4692 1704
rect 4812 1696 4820 1704
rect 5164 1696 5172 1704
rect 5228 1696 5236 1704
rect 5324 1696 5332 1704
rect 5548 1696 5556 1704
rect 5772 1696 5780 1704
rect 5900 1696 5908 1704
rect 6028 1696 6036 1704
rect 6140 1696 6148 1704
rect 6156 1696 6164 1704
rect 6220 1696 6228 1704
rect 6284 1696 6292 1704
rect 6444 1696 6452 1704
rect 6460 1696 6468 1704
rect 6476 1696 6484 1704
rect 268 1676 276 1684
rect 732 1676 740 1684
rect 780 1676 788 1684
rect 812 1676 820 1684
rect 1164 1676 1172 1684
rect 1244 1676 1252 1684
rect 1436 1676 1444 1684
rect 1564 1676 1572 1684
rect 3228 1676 3236 1684
rect 4700 1676 4708 1684
rect 4780 1676 4788 1684
rect 5068 1676 5076 1684
rect 5132 1676 5140 1684
rect 5388 1676 5396 1684
rect 6060 1676 6068 1684
rect 6108 1676 6116 1684
rect 6172 1676 6180 1684
rect 6188 1676 6196 1684
rect 6252 1676 6260 1684
rect 6348 1676 6356 1684
rect 6412 1676 6420 1684
rect 6508 1676 6516 1684
rect 6524 1676 6532 1684
rect 6556 1676 6564 1684
rect 716 1656 724 1664
rect 2380 1656 2388 1664
rect 5084 1656 5092 1664
rect 332 1636 340 1644
rect 940 1636 948 1644
rect 1084 1636 1092 1644
rect 1148 1636 1156 1644
rect 1260 1636 1268 1644
rect 1308 1636 1316 1644
rect 1340 1636 1348 1644
rect 1420 1636 1428 1644
rect 1484 1636 1492 1644
rect 1676 1636 1684 1644
rect 1852 1636 1860 1644
rect 2220 1636 2228 1644
rect 3036 1636 3044 1644
rect 3932 1636 3940 1644
rect 4044 1636 4052 1644
rect 4140 1636 4148 1644
rect 4172 1636 4180 1644
rect 4284 1636 4292 1644
rect 4460 1636 4468 1644
rect 4572 1636 4580 1644
rect 4620 1636 4628 1644
rect 4716 1636 4724 1644
rect 4764 1636 4772 1644
rect 4972 1636 4980 1644
rect 5036 1636 5044 1644
rect 5196 1636 5204 1644
rect 5628 1636 5636 1644
rect 6044 1636 6052 1644
rect 6092 1636 6100 1644
rect 6172 1636 6180 1644
rect 6236 1636 6244 1644
rect 6396 1636 6404 1644
rect 1774 1606 1782 1614
rect 1788 1606 1796 1614
rect 1802 1606 1810 1614
rect 4830 1606 4838 1614
rect 4844 1606 4852 1614
rect 4858 1606 4866 1614
rect 12 1576 20 1584
rect 140 1576 148 1584
rect 188 1576 196 1584
rect 236 1576 244 1584
rect 524 1576 532 1584
rect 636 1576 644 1584
rect 684 1576 692 1584
rect 1404 1576 1412 1584
rect 2988 1576 2996 1584
rect 3292 1576 3300 1584
rect 3548 1576 3556 1584
rect 4508 1576 4516 1584
rect 4540 1576 4548 1584
rect 4924 1576 4932 1584
rect 5084 1576 5092 1584
rect 5276 1576 5284 1584
rect 5324 1576 5332 1584
rect 6268 1576 6276 1584
rect 6412 1576 6420 1584
rect 6476 1576 6484 1584
rect 6508 1576 6516 1584
rect 4396 1556 4404 1564
rect 28 1536 36 1544
rect 92 1536 100 1544
rect 124 1536 132 1544
rect 204 1536 212 1544
rect 252 1536 260 1544
rect 508 1536 516 1544
rect 908 1536 916 1544
rect 972 1536 980 1544
rect 1228 1536 1236 1544
rect 2268 1536 2276 1544
rect 4028 1536 4036 1544
rect 4156 1536 4164 1544
rect 4380 1536 4388 1544
rect 4524 1536 4532 1544
rect 4556 1536 4564 1544
rect 60 1516 68 1524
rect 156 1516 164 1524
rect 284 1516 292 1524
rect 476 1516 484 1524
rect 540 1516 548 1524
rect 716 1516 724 1524
rect 764 1516 772 1524
rect 828 1516 836 1524
rect 940 1516 948 1524
rect 1004 1516 1012 1524
rect 1164 1516 1172 1524
rect 1260 1516 1268 1524
rect 44 1496 52 1504
rect 140 1496 148 1504
rect 188 1496 196 1504
rect 268 1496 276 1504
rect 300 1496 308 1504
rect 428 1496 436 1504
rect 524 1496 532 1504
rect 604 1496 612 1504
rect 620 1496 628 1504
rect 652 1496 660 1504
rect 684 1496 692 1504
rect 716 1496 724 1504
rect 860 1496 868 1504
rect 924 1496 932 1504
rect 972 1496 980 1504
rect 1084 1496 1092 1504
rect 1148 1496 1156 1504
rect 1196 1496 1204 1504
rect 1244 1496 1252 1504
rect 1276 1496 1284 1504
rect 1340 1496 1348 1504
rect 1436 1516 1444 1524
rect 1548 1516 1556 1524
rect 1596 1516 1604 1524
rect 1660 1516 1668 1524
rect 1676 1516 1684 1524
rect 1756 1516 1764 1524
rect 1980 1516 1988 1524
rect 2012 1516 2020 1524
rect 2092 1516 2100 1524
rect 2204 1516 2212 1524
rect 2476 1516 2484 1524
rect 2588 1516 2596 1524
rect 2636 1516 2644 1524
rect 2732 1516 2740 1524
rect 2892 1516 2900 1524
rect 2908 1516 2916 1524
rect 3404 1516 3412 1524
rect 3436 1516 3444 1524
rect 3676 1516 3684 1524
rect 3724 1516 3732 1524
rect 3772 1516 3780 1524
rect 3900 1516 3908 1524
rect 3916 1516 3924 1524
rect 4108 1516 4116 1524
rect 4140 1516 4148 1524
rect 4412 1516 4420 1524
rect 4460 1516 4468 1524
rect 4492 1516 4500 1524
rect 4524 1516 4532 1524
rect 1484 1496 1492 1504
rect 1532 1496 1540 1504
rect 1964 1496 1972 1504
rect 2060 1496 2068 1504
rect 2188 1496 2196 1504
rect 2252 1496 2260 1504
rect 2268 1496 2276 1504
rect 2300 1496 2308 1504
rect 2348 1496 2356 1504
rect 2412 1496 2420 1504
rect 2556 1496 2564 1504
rect 2620 1496 2628 1504
rect 2668 1496 2676 1504
rect 2796 1496 2804 1504
rect 3052 1494 3060 1502
rect 3116 1496 3124 1504
rect 3276 1496 3284 1504
rect 3324 1496 3332 1504
rect 3436 1496 3444 1504
rect 3452 1496 3460 1504
rect 3644 1496 3652 1504
rect 3852 1496 3860 1504
rect 4140 1496 4148 1504
rect 4348 1496 4356 1504
rect 4396 1496 4404 1504
rect 316 1476 324 1484
rect 76 1456 84 1464
rect 348 1456 356 1464
rect 380 1456 388 1464
rect 444 1476 452 1484
rect 588 1476 596 1484
rect 668 1476 676 1484
rect 780 1476 788 1484
rect 812 1476 820 1484
rect 876 1476 884 1484
rect 956 1476 964 1484
rect 1036 1476 1044 1484
rect 1068 1476 1076 1484
rect 1132 1476 1140 1484
rect 1196 1476 1204 1484
rect 1276 1476 1284 1484
rect 1324 1476 1332 1484
rect 1388 1476 1396 1484
rect 1420 1476 1428 1484
rect 1500 1476 1508 1484
rect 1564 1476 1572 1484
rect 1612 1476 1620 1484
rect 1708 1476 1716 1484
rect 1724 1476 1732 1484
rect 1820 1476 1828 1484
rect 1916 1476 1924 1484
rect 1932 1476 1940 1484
rect 2012 1476 2020 1484
rect 2092 1476 2100 1484
rect 2108 1476 2116 1484
rect 2124 1476 2132 1484
rect 2172 1476 2180 1484
rect 2220 1476 2228 1484
rect 2252 1476 2260 1484
rect 2364 1476 2372 1484
rect 2444 1476 2452 1484
rect 2508 1476 2516 1484
rect 2572 1476 2580 1484
rect 2620 1476 2628 1484
rect 2684 1476 2692 1484
rect 2700 1476 2708 1484
rect 2780 1476 2788 1484
rect 2924 1476 2932 1484
rect 3228 1476 3236 1484
rect 3244 1476 3252 1484
rect 3260 1476 3268 1484
rect 3372 1476 3380 1484
rect 3404 1476 3412 1484
rect 3484 1476 3492 1484
rect 3500 1476 3508 1484
rect 3596 1476 3604 1484
rect 556 1456 564 1464
rect 652 1456 660 1464
rect 748 1456 756 1464
rect 892 1456 900 1464
rect 1100 1456 1108 1464
rect 1436 1456 1444 1464
rect 1692 1456 1700 1464
rect 2140 1456 2148 1464
rect 2300 1456 2308 1464
rect 2380 1456 2388 1464
rect 2588 1456 2596 1464
rect 2748 1456 2756 1464
rect 2812 1456 2820 1464
rect 2876 1456 2884 1464
rect 2972 1456 2980 1464
rect 3324 1456 3332 1464
rect 3484 1456 3492 1464
rect 3644 1476 3652 1484
rect 3676 1476 3684 1484
rect 3692 1476 3700 1484
rect 3740 1476 3748 1484
rect 3804 1476 3812 1484
rect 3836 1476 3844 1484
rect 3868 1476 3876 1484
rect 3948 1476 3956 1484
rect 3964 1476 3972 1484
rect 4060 1476 4068 1484
rect 4076 1476 4084 1484
rect 4252 1476 4260 1484
rect 4332 1476 4340 1484
rect 4508 1496 4516 1504
rect 4620 1536 4628 1544
rect 4636 1536 4644 1544
rect 4732 1536 4740 1544
rect 4748 1536 4756 1544
rect 4908 1536 4916 1544
rect 5068 1536 5076 1544
rect 5484 1536 5492 1544
rect 5644 1536 5652 1544
rect 6044 1536 6052 1544
rect 6252 1536 6260 1544
rect 6284 1536 6292 1544
rect 6316 1536 6324 1544
rect 6332 1536 6340 1544
rect 6524 1536 6532 1544
rect 6588 1536 6596 1544
rect 4588 1516 4596 1524
rect 4620 1516 4628 1524
rect 4700 1516 4708 1524
rect 4716 1516 4724 1524
rect 4940 1516 4948 1524
rect 5036 1516 5044 1524
rect 5100 1516 5108 1524
rect 5212 1516 5220 1524
rect 5292 1516 5300 1524
rect 5484 1516 5492 1524
rect 5676 1516 5684 1524
rect 6204 1516 6212 1524
rect 6284 1516 6292 1524
rect 6348 1516 6356 1524
rect 6364 1516 6372 1524
rect 6396 1516 6404 1524
rect 6492 1516 6500 1524
rect 6556 1516 6564 1524
rect 4620 1496 4628 1504
rect 4652 1496 4660 1504
rect 4732 1496 4740 1504
rect 4780 1496 4788 1504
rect 4924 1496 4932 1504
rect 4956 1496 4964 1504
rect 5084 1496 5092 1504
rect 5164 1496 5172 1504
rect 5228 1496 5236 1504
rect 5324 1496 5332 1504
rect 5340 1496 5348 1504
rect 5468 1496 5476 1504
rect 5564 1496 5572 1504
rect 5644 1496 5652 1504
rect 5756 1496 5764 1504
rect 5772 1496 5780 1504
rect 5804 1496 5812 1504
rect 5852 1496 5860 1504
rect 5932 1496 5940 1504
rect 5964 1496 5972 1504
rect 6012 1496 6020 1504
rect 6044 1496 6052 1504
rect 6076 1496 6084 1504
rect 6124 1496 6132 1504
rect 6172 1496 6180 1504
rect 6220 1496 6228 1504
rect 6268 1496 6276 1504
rect 6332 1496 6340 1504
rect 6380 1496 6388 1504
rect 6428 1496 6436 1504
rect 6508 1496 6516 1504
rect 6572 1496 6580 1504
rect 4668 1476 4676 1484
rect 4796 1476 4804 1484
rect 4972 1476 4980 1484
rect 3916 1456 3924 1464
rect 4108 1456 4116 1464
rect 4188 1456 4196 1464
rect 4268 1456 4276 1464
rect 4844 1456 4852 1464
rect 5148 1476 5156 1484
rect 5180 1476 5188 1484
rect 5244 1476 5252 1484
rect 5340 1476 5348 1484
rect 5372 1476 5380 1484
rect 5404 1476 5412 1484
rect 5628 1476 5636 1484
rect 5740 1476 5748 1484
rect 5772 1476 5780 1484
rect 5836 1476 5844 1484
rect 5868 1476 5876 1484
rect 5916 1476 5924 1484
rect 5980 1476 5988 1484
rect 5996 1476 6004 1484
rect 6060 1476 6068 1484
rect 6076 1476 6084 1484
rect 6140 1476 6148 1484
rect 6220 1476 6228 1484
rect 6444 1476 6452 1484
rect 5020 1456 5028 1464
rect 5116 1456 5124 1464
rect 5276 1456 5284 1464
rect 5596 1456 5604 1464
rect 5788 1456 5796 1464
rect 5900 1456 5908 1464
rect 6124 1456 6132 1464
rect 6332 1456 6340 1464
rect 6476 1456 6484 1464
rect 332 1436 340 1444
rect 412 1436 420 1444
rect 460 1436 468 1444
rect 572 1436 580 1444
rect 1036 1436 1044 1444
rect 1116 1436 1124 1444
rect 1212 1436 1220 1444
rect 1292 1436 1300 1444
rect 1356 1436 1364 1444
rect 1580 1436 1588 1444
rect 1660 1436 1668 1444
rect 1676 1436 1684 1444
rect 1740 1436 1748 1444
rect 1852 1436 1860 1444
rect 1948 1436 1956 1444
rect 2156 1436 2164 1444
rect 2396 1436 2404 1444
rect 2524 1436 2532 1444
rect 2716 1436 2724 1444
rect 2764 1436 2772 1444
rect 2828 1436 2836 1444
rect 2956 1436 2964 1444
rect 3180 1436 3188 1444
rect 3196 1436 3204 1444
rect 3372 1436 3380 1444
rect 3388 1436 3396 1444
rect 3404 1436 3412 1444
rect 3724 1436 3732 1444
rect 3836 1436 3844 1444
rect 3900 1436 3908 1444
rect 4172 1436 4180 1444
rect 4236 1436 4244 1444
rect 4316 1436 4324 1444
rect 4460 1436 4468 1444
rect 4684 1436 4692 1444
rect 4764 1436 4772 1444
rect 4812 1436 4820 1444
rect 4988 1436 4996 1444
rect 5132 1436 5140 1444
rect 5212 1436 5220 1444
rect 5404 1436 5412 1444
rect 5580 1436 5588 1444
rect 5820 1436 5828 1444
rect 5884 1436 5892 1444
rect 5932 1436 5940 1444
rect 6380 1436 6388 1444
rect 6572 1436 6580 1444
rect 5228 1416 5236 1424
rect 3310 1406 3318 1414
rect 3324 1406 3332 1414
rect 3338 1406 3346 1414
rect 108 1376 116 1384
rect 156 1376 164 1384
rect 204 1376 212 1384
rect 252 1376 260 1384
rect 316 1376 324 1384
rect 396 1376 404 1384
rect 860 1376 868 1384
rect 1724 1376 1732 1384
rect 2188 1376 2196 1384
rect 2316 1376 2324 1384
rect 3020 1376 3028 1384
rect 4092 1376 4100 1384
rect 4252 1376 4260 1384
rect 4332 1376 4340 1384
rect 4716 1376 4724 1384
rect 4924 1376 4932 1384
rect 4988 1376 4996 1384
rect 5260 1376 5268 1384
rect 5356 1376 5364 1384
rect 5500 1376 5508 1384
rect 5612 1376 5620 1384
rect 5660 1376 5668 1384
rect 5836 1376 5844 1384
rect 5900 1376 5908 1384
rect 6172 1376 6180 1384
rect 6396 1376 6404 1384
rect 124 1356 132 1364
rect 412 1356 420 1364
rect 572 1356 580 1364
rect 780 1356 788 1364
rect 1052 1356 1060 1364
rect 1932 1356 1940 1364
rect 2012 1356 2020 1364
rect 2156 1356 2164 1364
rect 2220 1356 2228 1364
rect 2700 1356 2708 1364
rect 2988 1356 2996 1364
rect 3116 1356 3124 1364
rect 3164 1356 3172 1364
rect 3308 1356 3316 1364
rect 3388 1356 3396 1364
rect 3468 1356 3476 1364
rect 3500 1356 3508 1364
rect 3516 1356 3524 1364
rect 3548 1356 3556 1364
rect 3756 1356 3764 1364
rect 3964 1356 3972 1364
rect 4028 1356 4036 1364
rect 4140 1356 4148 1364
rect 4188 1356 4196 1364
rect 4700 1356 4708 1364
rect 5132 1356 5140 1364
rect 44 1336 52 1344
rect 92 1336 100 1344
rect 172 1336 180 1344
rect 220 1336 228 1344
rect 380 1336 388 1344
rect 668 1336 676 1344
rect 684 1336 692 1344
rect 764 1336 772 1344
rect 812 1336 820 1344
rect 44 1316 52 1324
rect 76 1316 84 1324
rect 252 1316 260 1324
rect 332 1316 340 1324
rect 364 1316 372 1324
rect 460 1316 468 1324
rect 524 1316 532 1324
rect 604 1316 612 1324
rect 60 1296 68 1304
rect 140 1296 148 1304
rect 188 1296 196 1304
rect 236 1296 244 1304
rect 348 1296 356 1304
rect 476 1296 484 1304
rect 540 1296 548 1304
rect 588 1296 596 1304
rect 652 1296 660 1304
rect 796 1316 804 1324
rect 1148 1336 1156 1344
rect 1212 1336 1220 1344
rect 1324 1336 1332 1344
rect 1420 1336 1428 1344
rect 1564 1336 1572 1344
rect 1660 1336 1668 1344
rect 1708 1336 1716 1344
rect 1756 1336 1764 1344
rect 1772 1336 1780 1344
rect 1868 1336 1876 1344
rect 1900 1336 1908 1344
rect 1996 1336 2004 1344
rect 2092 1336 2100 1344
rect 2204 1336 2212 1344
rect 2252 1336 2260 1344
rect 2364 1336 2372 1344
rect 2444 1336 2452 1344
rect 2540 1336 2548 1344
rect 2620 1336 2628 1344
rect 2668 1336 2676 1344
rect 2732 1336 2740 1344
rect 2780 1336 2788 1344
rect 2892 1336 2900 1344
rect 2924 1336 2932 1344
rect 2940 1336 2948 1344
rect 3068 1336 3076 1344
rect 3292 1336 3300 1344
rect 3404 1336 3412 1344
rect 3580 1336 3588 1344
rect 3612 1336 3620 1344
rect 3644 1336 3652 1344
rect 3708 1336 3716 1344
rect 3788 1336 3796 1344
rect 3996 1336 4004 1344
rect 4060 1336 4068 1344
rect 4092 1336 4100 1344
rect 4124 1336 4132 1344
rect 4188 1336 4196 1344
rect 4236 1336 4244 1344
rect 4284 1336 4292 1344
rect 4300 1336 4308 1344
rect 4396 1336 4404 1344
rect 4412 1336 4420 1344
rect 4476 1336 4484 1344
rect 4748 1336 4756 1344
rect 940 1316 948 1324
rect 1004 1316 1012 1324
rect 1084 1316 1092 1324
rect 1116 1316 1124 1324
rect 1292 1316 1300 1324
rect 1340 1316 1348 1324
rect 1468 1316 1476 1324
rect 1532 1316 1540 1324
rect 1660 1316 1668 1324
rect 1932 1316 1940 1324
rect 2060 1316 2068 1324
rect 2108 1316 2116 1324
rect 2348 1316 2356 1324
rect 2364 1316 2372 1324
rect 2412 1316 2420 1324
rect 2492 1316 2500 1324
rect 2540 1316 2548 1324
rect 2588 1316 2596 1324
rect 2620 1316 2628 1324
rect 2652 1316 2660 1324
rect 2684 1316 2692 1324
rect 2796 1316 2804 1324
rect 2812 1316 2820 1324
rect 2940 1316 2948 1324
rect 3052 1316 3060 1324
rect 3132 1316 3140 1324
rect 3212 1316 3220 1324
rect 3276 1316 3284 1324
rect 3404 1316 3412 1324
rect 3420 1316 3428 1324
rect 3468 1316 3476 1324
rect 3548 1316 3556 1324
rect 3564 1316 3572 1324
rect 3596 1316 3604 1324
rect 3628 1316 3636 1324
rect 3660 1316 3668 1324
rect 3756 1316 3764 1324
rect 3852 1316 3860 1324
rect 3932 1316 3940 1324
rect 4012 1316 4020 1324
rect 4044 1316 4052 1324
rect 4108 1316 4116 1324
rect 4428 1316 4436 1324
rect 4492 1316 4500 1324
rect 4524 1316 4532 1324
rect 4556 1316 4564 1324
rect 4620 1316 4628 1324
rect 4668 1316 4676 1324
rect 4860 1336 4868 1344
rect 4956 1332 4964 1340
rect 4988 1336 4996 1344
rect 5020 1336 5028 1344
rect 5068 1336 5076 1344
rect 5116 1336 5124 1344
rect 5196 1356 5204 1364
rect 5276 1356 5284 1364
rect 5308 1356 5316 1364
rect 5420 1356 5428 1364
rect 5436 1356 5444 1364
rect 5212 1336 5220 1344
rect 5260 1336 5268 1344
rect 5340 1336 5348 1344
rect 5372 1336 5380 1344
rect 5644 1356 5652 1364
rect 5804 1356 5812 1364
rect 5820 1356 5828 1364
rect 5948 1356 5956 1364
rect 6044 1356 6052 1364
rect 6060 1356 6068 1364
rect 6076 1356 6084 1364
rect 6156 1356 6164 1364
rect 6524 1356 6532 1364
rect 5564 1336 5572 1344
rect 5660 1336 5668 1344
rect 5756 1336 5764 1344
rect 5852 1336 5860 1344
rect 5884 1336 5892 1344
rect 6108 1336 6116 1344
rect 6172 1336 6180 1344
rect 876 1296 884 1304
rect 924 1296 932 1304
rect 988 1296 996 1304
rect 1084 1296 1092 1304
rect 1196 1296 1204 1304
rect 1244 1296 1252 1304
rect 1308 1296 1316 1304
rect 1484 1296 1492 1304
rect 1548 1296 1556 1304
rect 1676 1296 1684 1304
rect 1724 1296 1732 1304
rect 1756 1296 1764 1304
rect 1820 1296 1828 1304
rect 1868 1296 1876 1304
rect 1948 1296 1956 1304
rect 2124 1296 2132 1304
rect 2172 1296 2180 1304
rect 2300 1296 2308 1304
rect 2316 1296 2324 1304
rect 2380 1296 2388 1304
rect 2508 1296 2516 1304
rect 2604 1296 2612 1304
rect 2828 1296 2836 1304
rect 2844 1296 2852 1304
rect 2956 1296 2964 1304
rect 2972 1296 2980 1304
rect 3020 1296 3028 1304
rect 3228 1296 3236 1304
rect 3244 1296 3252 1304
rect 3452 1296 3460 1304
rect 3692 1296 3700 1304
rect 3708 1296 3716 1304
rect 3820 1296 3828 1304
rect 3836 1296 3844 1304
rect 3900 1296 3908 1304
rect 4236 1296 4244 1304
rect 4460 1296 4468 1304
rect 4540 1296 4548 1304
rect 4604 1296 4612 1304
rect 4860 1316 4868 1324
rect 4876 1316 4884 1324
rect 5180 1316 5188 1324
rect 5308 1316 5316 1324
rect 5324 1316 5332 1324
rect 5436 1316 5444 1324
rect 5484 1316 5492 1324
rect 5580 1316 5588 1324
rect 4876 1296 4884 1304
rect 4908 1296 4916 1304
rect 4988 1296 4996 1304
rect 5036 1296 5044 1304
rect 5228 1296 5236 1304
rect 5644 1316 5652 1324
rect 5676 1316 5684 1324
rect 5772 1316 5780 1324
rect 5868 1316 5876 1324
rect 5884 1316 5892 1324
rect 5932 1316 5940 1324
rect 5964 1316 5972 1324
rect 6012 1316 6020 1324
rect 6124 1316 6132 1324
rect 6188 1316 6196 1324
rect 6284 1316 6292 1324
rect 6348 1316 6356 1324
rect 6428 1316 6436 1324
rect 6492 1316 6500 1324
rect 6556 1316 6564 1324
rect 5804 1296 5812 1304
rect 5948 1296 5956 1304
rect 6268 1296 6276 1304
rect 6332 1296 6340 1304
rect 6444 1296 6452 1304
rect 6508 1296 6516 1304
rect 28 1276 36 1284
rect 268 1276 276 1284
rect 316 1276 324 1284
rect 444 1276 452 1284
rect 508 1276 516 1284
rect 620 1276 628 1284
rect 956 1276 964 1284
rect 1020 1276 1028 1284
rect 1276 1276 1284 1284
rect 1388 1276 1396 1284
rect 1452 1276 1460 1284
rect 1548 1276 1556 1284
rect 1932 1276 1940 1284
rect 2572 1276 2580 1284
rect 2764 1276 2772 1284
rect 3148 1276 3156 1284
rect 3196 1276 3204 1284
rect 3484 1276 3492 1284
rect 3804 1276 3812 1284
rect 4556 1276 4564 1284
rect 4636 1276 4644 1284
rect 4844 1276 4852 1284
rect 5500 1276 5508 1284
rect 5532 1276 5540 1284
rect 5996 1276 6004 1284
rect 6300 1276 6308 1284
rect 6364 1276 6372 1284
rect 6412 1276 6420 1284
rect 6572 1276 6580 1284
rect 604 1256 612 1264
rect 1468 1256 1476 1264
rect 3772 1256 3780 1264
rect 3980 1256 3988 1264
rect 428 1236 436 1244
rect 492 1236 500 1244
rect 556 1236 564 1244
rect 892 1236 900 1244
rect 972 1236 980 1244
rect 1004 1236 1012 1244
rect 1116 1236 1124 1244
rect 1164 1236 1172 1244
rect 1228 1236 1236 1244
rect 1260 1236 1268 1244
rect 1404 1236 1412 1244
rect 1500 1236 1508 1244
rect 1596 1236 1604 1244
rect 1884 1236 1892 1244
rect 2188 1236 2196 1244
rect 2268 1236 2276 1244
rect 2460 1236 2468 1244
rect 2876 1236 2884 1244
rect 3004 1236 3012 1244
rect 3100 1236 3108 1244
rect 3212 1236 3220 1244
rect 3276 1236 3284 1244
rect 3884 1236 3892 1244
rect 3932 1236 3940 1244
rect 4028 1236 4036 1244
rect 4428 1236 4436 1244
rect 4556 1236 4564 1244
rect 4652 1236 4660 1244
rect 5084 1236 5092 1244
rect 5164 1236 5172 1244
rect 5244 1236 5252 1244
rect 5308 1236 5316 1244
rect 6012 1236 6020 1244
rect 6076 1236 6084 1244
rect 6284 1236 6292 1244
rect 6380 1236 6388 1244
rect 6396 1236 6404 1244
rect 6460 1236 6468 1244
rect 6556 1236 6564 1244
rect 1774 1206 1782 1214
rect 1788 1206 1796 1214
rect 1802 1206 1810 1214
rect 4830 1206 4838 1214
rect 4844 1206 4852 1214
rect 4858 1206 4866 1214
rect 44 1176 52 1184
rect 156 1176 164 1184
rect 220 1176 228 1184
rect 284 1176 292 1184
rect 348 1176 356 1184
rect 684 1176 692 1184
rect 1964 1176 1972 1184
rect 2284 1176 2292 1184
rect 4972 1176 4980 1184
rect 6252 1176 6260 1184
rect 6300 1176 6308 1184
rect 2124 1156 2132 1164
rect 2956 1156 2964 1164
rect 4476 1156 4484 1164
rect 4604 1156 4612 1164
rect 5356 1156 5364 1164
rect 28 1136 36 1144
rect 172 1136 180 1144
rect 236 1136 244 1144
rect 300 1136 308 1144
rect 364 1136 372 1144
rect 636 1136 644 1144
rect 1916 1136 1924 1144
rect 2140 1136 2148 1144
rect 2188 1136 2196 1144
rect 2972 1136 2980 1144
rect 3020 1136 3028 1144
rect 3548 1136 3556 1144
rect 4348 1136 4356 1144
rect 4396 1136 4404 1144
rect 4460 1136 4468 1144
rect 4668 1136 4676 1144
rect 5724 1136 5732 1144
rect 5900 1136 5908 1144
rect 5964 1136 5972 1144
rect 6044 1136 6052 1144
rect 6364 1136 6372 1144
rect 60 1116 68 1124
rect 76 1116 84 1124
rect 140 1116 148 1124
rect 204 1116 212 1124
rect 268 1116 276 1124
rect 332 1116 340 1124
rect 428 1116 436 1124
rect 444 1116 452 1124
rect 44 1096 52 1104
rect 76 1096 84 1104
rect 108 1096 116 1104
rect 156 1096 164 1104
rect 220 1096 228 1104
rect 284 1096 292 1104
rect 348 1096 356 1104
rect 476 1096 484 1104
rect 492 1096 500 1104
rect 556 1116 564 1124
rect 668 1116 676 1124
rect 716 1116 724 1124
rect 764 1116 772 1124
rect 812 1116 820 1124
rect 940 1116 948 1124
rect 988 1116 996 1124
rect 1036 1116 1044 1124
rect 1420 1116 1428 1124
rect 1468 1116 1476 1124
rect 1484 1116 1492 1124
rect 1532 1116 1540 1124
rect 1548 1116 1556 1124
rect 1580 1116 1588 1124
rect 1628 1116 1636 1124
rect 1852 1116 1860 1124
rect 1948 1116 1956 1124
rect 2060 1116 2068 1124
rect 2108 1116 2116 1124
rect 2172 1116 2180 1124
rect 2300 1116 2308 1124
rect 2396 1116 2404 1124
rect 2476 1116 2484 1124
rect 2668 1116 2676 1124
rect 2764 1116 2772 1124
rect 2844 1116 2852 1124
rect 2924 1116 2932 1124
rect 2940 1116 2948 1124
rect 3052 1116 3060 1124
rect 3084 1116 3092 1124
rect 3116 1116 3124 1124
rect 3388 1116 3396 1124
rect 3468 1116 3476 1124
rect 3580 1116 3588 1124
rect 3612 1116 3620 1124
rect 3628 1116 3636 1124
rect 124 1076 132 1084
rect 396 1076 404 1084
rect 492 1076 500 1084
rect 588 1096 596 1104
rect 796 1096 804 1104
rect 860 1096 868 1104
rect 924 1096 932 1104
rect 1116 1096 1124 1104
rect 1148 1096 1156 1104
rect 1244 1096 1252 1104
rect 1292 1096 1300 1104
rect 1372 1096 1380 1104
rect 1676 1096 1684 1104
rect 1820 1096 1828 1104
rect 1884 1096 1892 1104
rect 1932 1096 1940 1104
rect 2028 1096 2036 1104
rect 2124 1096 2132 1104
rect 2188 1096 2196 1104
rect 2236 1096 2244 1104
rect 2332 1096 2340 1104
rect 2508 1096 2516 1104
rect 2556 1096 2564 1104
rect 2924 1096 2932 1104
rect 2956 1096 2964 1104
rect 3036 1096 3044 1104
rect 3084 1096 3092 1104
rect 3180 1096 3188 1104
rect 3244 1096 3252 1104
rect 3340 1096 3348 1104
rect 3372 1096 3380 1104
rect 3564 1096 3572 1104
rect 3692 1116 3700 1124
rect 3932 1116 3940 1124
rect 620 1076 628 1084
rect 748 1076 756 1084
rect 796 1076 804 1084
rect 876 1076 884 1084
rect 908 1076 916 1084
rect 972 1076 980 1084
rect 1020 1076 1028 1084
rect 1068 1076 1076 1084
rect 1132 1076 1140 1084
rect 1164 1076 1172 1084
rect 700 1056 708 1064
rect 764 1056 772 1064
rect 1308 1076 1316 1084
rect 1356 1076 1364 1084
rect 1372 1076 1380 1084
rect 1436 1076 1444 1084
rect 1468 1076 1476 1084
rect 1516 1076 1524 1084
rect 1564 1076 1572 1084
rect 1692 1076 1700 1084
rect 1852 1076 1860 1084
rect 2060 1076 2068 1084
rect 2092 1076 2100 1084
rect 2252 1076 2260 1084
rect 2428 1076 2436 1084
rect 2572 1076 2580 1084
rect 2700 1076 2708 1084
rect 2716 1076 2724 1084
rect 2876 1076 2884 1084
rect 3116 1076 3124 1084
rect 3148 1076 3156 1084
rect 3196 1076 3204 1084
rect 3420 1076 3428 1084
rect 3436 1076 3444 1084
rect 3484 1076 3492 1084
rect 3548 1076 3556 1084
rect 3724 1096 3732 1104
rect 3788 1096 3796 1104
rect 3868 1096 3876 1104
rect 3980 1116 3988 1124
rect 4124 1116 4132 1124
rect 4172 1116 4180 1124
rect 4204 1116 4212 1124
rect 4428 1116 4436 1124
rect 4492 1116 4500 1124
rect 4588 1116 4596 1124
rect 4636 1116 4644 1124
rect 5292 1116 5300 1124
rect 5436 1116 5444 1124
rect 5484 1116 5492 1124
rect 5532 1116 5540 1124
rect 5628 1116 5636 1124
rect 5740 1116 5748 1124
rect 6012 1116 6020 1124
rect 6060 1116 6068 1124
rect 6076 1116 6084 1124
rect 6140 1116 6148 1124
rect 6284 1116 6292 1124
rect 6332 1116 6340 1124
rect 6508 1116 6516 1124
rect 6636 1116 6644 1124
rect 4012 1096 4020 1104
rect 4092 1096 4100 1104
rect 4204 1096 4212 1104
rect 4252 1096 4260 1104
rect 3644 1076 3652 1084
rect 3740 1076 3748 1084
rect 1212 1056 1220 1064
rect 1324 1056 1332 1064
rect 1468 1056 1476 1064
rect 1724 1056 1732 1064
rect 1980 1056 1988 1064
rect 2284 1056 2292 1064
rect 2348 1056 2356 1064
rect 2652 1056 2660 1064
rect 2828 1056 2836 1064
rect 3004 1056 3012 1064
rect 3164 1056 3172 1064
rect 3228 1056 3236 1064
rect 3276 1056 3284 1064
rect 3372 1056 3380 1064
rect 3884 1076 3892 1084
rect 3932 1076 3940 1084
rect 4124 1076 4132 1084
rect 4156 1076 4164 1084
rect 4220 1076 4228 1084
rect 4236 1076 4244 1084
rect 4476 1096 4484 1104
rect 4588 1096 4596 1104
rect 4652 1096 4660 1104
rect 4700 1096 4708 1104
rect 5004 1096 5012 1104
rect 5084 1096 5092 1104
rect 5164 1096 5172 1104
rect 5244 1096 5252 1104
rect 5260 1096 5268 1104
rect 5324 1096 5332 1104
rect 5372 1096 5380 1104
rect 5580 1096 5588 1104
rect 5612 1096 5620 1104
rect 5660 1096 5668 1104
rect 5724 1096 5732 1104
rect 5884 1096 5892 1104
rect 5980 1096 5988 1104
rect 6028 1096 6036 1104
rect 6124 1096 6132 1104
rect 6172 1096 6180 1104
rect 6204 1096 6212 1104
rect 6268 1096 6276 1104
rect 6348 1096 6356 1104
rect 6396 1096 6404 1104
rect 6508 1096 6516 1104
rect 6572 1096 6580 1104
rect 6588 1096 6596 1104
rect 4524 1076 4532 1084
rect 4556 1076 4564 1084
rect 4620 1076 4628 1084
rect 4716 1076 4724 1084
rect 4812 1076 4820 1084
rect 4828 1076 4836 1084
rect 4956 1076 4964 1084
rect 5132 1076 5140 1084
rect 5228 1076 5236 1084
rect 5292 1076 5300 1084
rect 5340 1076 5348 1084
rect 3820 1056 3828 1064
rect 3836 1056 3844 1064
rect 3852 1056 3860 1064
rect 4060 1056 4068 1064
rect 4652 1056 4660 1064
rect 4748 1056 4756 1064
rect 4796 1056 4804 1064
rect 4988 1056 4996 1064
rect 5004 1056 5012 1064
rect 5052 1056 5060 1064
rect 5084 1056 5092 1064
rect 5116 1056 5124 1064
rect 5212 1056 5220 1064
rect 5388 1076 5396 1084
rect 5436 1076 5444 1084
rect 5452 1076 5460 1084
rect 5500 1076 5508 1084
rect 5532 1076 5540 1084
rect 5676 1076 5684 1084
rect 5724 1076 5732 1084
rect 5772 1076 5780 1084
rect 5820 1080 5828 1088
rect 5932 1076 5940 1084
rect 5980 1076 5988 1084
rect 6124 1076 6132 1084
rect 6156 1076 6164 1084
rect 6188 1076 6196 1084
rect 6204 1076 6212 1084
rect 6284 1076 6292 1084
rect 6316 1076 6324 1084
rect 6412 1076 6420 1084
rect 6444 1076 6452 1084
rect 6556 1076 6564 1084
rect 5692 1056 5700 1064
rect 5852 1056 5860 1064
rect 5884 1056 5892 1064
rect 6444 1056 6452 1064
rect 6524 1056 6532 1064
rect 412 1036 420 1044
rect 444 1036 452 1044
rect 524 1036 532 1044
rect 684 1036 692 1044
rect 716 1036 724 1044
rect 876 1036 884 1044
rect 956 1036 964 1044
rect 988 1036 996 1044
rect 1036 1036 1044 1044
rect 1084 1036 1092 1044
rect 1180 1036 1188 1044
rect 1260 1036 1268 1044
rect 1340 1036 1348 1044
rect 1404 1036 1412 1044
rect 1596 1036 1604 1044
rect 1628 1036 1636 1044
rect 1708 1036 1716 1044
rect 1740 1036 1748 1044
rect 1852 1036 1860 1044
rect 1996 1036 2004 1044
rect 2060 1036 2068 1044
rect 2204 1036 2212 1044
rect 2300 1036 2308 1044
rect 2396 1036 2404 1044
rect 2460 1036 2468 1044
rect 2508 1036 2516 1044
rect 2620 1036 2628 1044
rect 2684 1036 2692 1044
rect 2700 1036 2708 1044
rect 2716 1036 2724 1044
rect 2732 1036 2740 1044
rect 2764 1036 2772 1044
rect 2780 1036 2788 1044
rect 2860 1036 2868 1044
rect 3132 1036 3140 1044
rect 3260 1036 3268 1044
rect 3420 1036 3428 1044
rect 3452 1036 3460 1044
rect 3500 1036 3508 1044
rect 3676 1036 3684 1044
rect 3772 1036 3780 1044
rect 3916 1036 3924 1044
rect 3948 1036 3956 1044
rect 4204 1036 4212 1044
rect 4284 1036 4292 1044
rect 4300 1036 4308 1044
rect 4540 1036 4548 1044
rect 4892 1036 4900 1044
rect 5100 1036 5108 1044
rect 5196 1036 5204 1044
rect 5468 1036 5476 1044
rect 5596 1036 5604 1044
rect 5788 1036 5796 1044
rect 5868 1036 5876 1044
rect 5932 1036 5940 1044
rect 6076 1036 6084 1044
rect 6348 1036 6356 1044
rect 6428 1036 6436 1044
rect 6540 1036 6548 1044
rect 3036 1016 3044 1024
rect 3820 1016 3828 1024
rect 4060 1016 4068 1024
rect 5164 1016 5172 1024
rect 5692 1016 5700 1024
rect 3310 1006 3318 1014
rect 3324 1006 3332 1014
rect 3338 1006 3346 1014
rect 2668 996 2676 1004
rect 3388 996 3396 1004
rect 3420 996 3428 1004
rect 3516 996 3524 1004
rect 3628 996 3636 1004
rect 4428 996 4436 1004
rect 5420 996 5428 1004
rect 44 976 52 984
rect 92 976 100 984
rect 172 976 180 984
rect 332 976 340 984
rect 412 976 420 984
rect 1020 976 1028 984
rect 2300 976 2308 984
rect 2892 976 2900 984
rect 2924 976 2932 984
rect 2956 976 2964 984
rect 3068 976 3076 984
rect 3116 976 3124 984
rect 3164 976 3172 984
rect 3596 976 3604 984
rect 3708 976 3716 984
rect 4268 976 4276 984
rect 4364 976 4372 984
rect 4476 976 4484 984
rect 4604 976 4612 984
rect 4668 976 4676 984
rect 4716 976 4724 984
rect 5324 976 5332 984
rect 5452 976 5460 984
rect 5580 976 5588 984
rect 5772 976 5780 984
rect 5804 976 5812 984
rect 6188 976 6196 984
rect 60 956 68 964
rect 76 956 84 964
rect 1100 956 1108 964
rect 1132 956 1140 964
rect 1516 956 1524 964
rect 1900 956 1908 964
rect 2188 956 2196 964
rect 2220 956 2228 964
rect 2284 956 2292 964
rect 2348 956 2356 964
rect 2364 956 2372 964
rect 2636 956 2644 964
rect 2684 956 2692 964
rect 3100 956 3108 964
rect 3148 956 3156 964
rect 3212 956 3220 964
rect 3420 956 3428 964
rect 3516 956 3524 964
rect 3628 956 3636 964
rect 3756 956 3764 964
rect 3836 956 3844 964
rect 4012 956 4020 964
rect 4188 956 4196 964
rect 28 936 36 944
rect 108 936 116 944
rect 316 936 324 944
rect 380 936 388 944
rect 460 936 468 944
rect 12 916 20 924
rect 172 916 180 924
rect 236 916 244 924
rect 300 916 308 924
rect 364 916 372 924
rect 412 916 420 924
rect 492 936 500 944
rect 556 936 564 944
rect 620 936 628 944
rect 652 936 660 944
rect 700 936 708 944
rect 972 936 980 944
rect 1180 936 1188 944
rect 1196 936 1204 944
rect 1276 936 1284 944
rect 1404 936 1412 944
rect 1468 936 1476 944
rect 2300 936 2308 944
rect 2364 936 2372 944
rect 2428 936 2436 944
rect 2444 936 2452 944
rect 2540 936 2548 944
rect 2604 936 2612 944
rect 2780 936 2788 944
rect 2812 936 2820 944
rect 2844 932 2852 940
rect 2924 936 2932 944
rect 2956 936 2964 944
rect 3036 936 3044 944
rect 3068 936 3076 944
rect 3132 936 3140 944
rect 508 916 516 924
rect 572 916 580 924
rect 604 916 612 924
rect 636 916 644 924
rect 700 916 708 924
rect 732 916 740 924
rect 812 916 820 924
rect 860 916 868 924
rect 924 916 932 924
rect 988 916 996 924
rect 1052 916 1060 924
rect 1100 916 1108 924
rect 1132 916 1140 924
rect 188 896 196 904
rect 252 896 260 904
rect 268 896 276 904
rect 332 896 340 904
rect 396 896 404 904
rect 540 896 548 904
rect 716 896 724 904
rect 844 896 852 904
rect 908 896 916 904
rect 1020 896 1028 904
rect 1036 896 1044 904
rect 1148 896 1156 904
rect 1324 916 1332 924
rect 1372 916 1380 924
rect 1388 916 1396 924
rect 1436 916 1444 924
rect 1452 916 1460 924
rect 1484 916 1492 924
rect 1500 916 1508 924
rect 1564 916 1572 924
rect 1612 916 1620 924
rect 1692 916 1700 924
rect 1740 916 1748 924
rect 1852 916 1860 924
rect 1932 916 1940 924
rect 1964 916 1972 924
rect 2012 916 2020 924
rect 2092 916 2100 924
rect 2156 916 2164 924
rect 2300 916 2308 924
rect 2364 916 2372 924
rect 2412 916 2420 924
rect 2492 916 2500 924
rect 2556 916 2564 924
rect 2668 916 2676 924
rect 2732 916 2740 924
rect 3052 916 3060 924
rect 3180 916 3188 924
rect 3596 936 3604 944
rect 3756 936 3764 944
rect 3788 936 3796 944
rect 3852 936 3860 944
rect 3948 936 3956 944
rect 4028 936 4036 944
rect 4156 936 4164 944
rect 4332 956 4340 964
rect 4348 956 4356 964
rect 4412 956 4420 964
rect 4300 936 4308 944
rect 4540 956 4548 964
rect 4556 956 4564 964
rect 4684 956 4692 964
rect 4812 956 4820 964
rect 5036 956 5044 964
rect 5132 956 5140 964
rect 5228 956 5236 964
rect 5292 956 5300 964
rect 5420 956 5428 964
rect 5436 956 5444 964
rect 5740 956 5748 964
rect 5884 956 5892 964
rect 6476 956 6484 964
rect 6556 956 6564 964
rect 4524 936 4532 944
rect 4572 936 4580 944
rect 4636 936 4644 944
rect 4732 936 4740 944
rect 4908 936 4916 944
rect 5004 936 5012 944
rect 5020 936 5028 944
rect 5100 936 5108 944
rect 3372 916 3380 924
rect 3420 916 3428 924
rect 3468 916 3476 924
rect 3564 916 3572 924
rect 3596 916 3604 924
rect 3932 916 3940 924
rect 3996 916 4004 924
rect 4108 916 4116 924
rect 4140 916 4148 924
rect 4236 916 4244 924
rect 4252 916 4260 924
rect 4444 916 4452 924
rect 4460 916 4468 924
rect 4508 916 4516 924
rect 4652 916 4660 924
rect 4780 916 4788 924
rect 4908 916 4916 924
rect 4956 916 4964 924
rect 5196 936 5204 944
rect 5212 936 5220 944
rect 5276 936 5284 944
rect 5388 936 5396 944
rect 5404 936 5412 944
rect 5484 936 5492 944
rect 5660 936 5668 944
rect 5676 936 5684 944
rect 5724 936 5732 944
rect 5772 936 5780 944
rect 6156 936 6164 944
rect 6300 936 6308 944
rect 6444 936 6452 944
rect 6588 936 6596 944
rect 5036 916 5044 924
rect 5068 916 5076 924
rect 5100 916 5108 924
rect 5132 916 5140 924
rect 5228 916 5236 924
rect 5260 916 5268 924
rect 5372 916 5380 924
rect 5500 916 5508 924
rect 5548 916 5556 924
rect 5612 916 5620 924
rect 5708 916 5716 924
rect 5820 916 5828 924
rect 5932 916 5940 924
rect 5980 916 5988 924
rect 6044 916 6052 924
rect 6108 916 6116 924
rect 6236 916 6244 924
rect 6300 916 6308 924
rect 6348 916 6356 924
rect 6428 916 6436 924
rect 6524 916 6532 924
rect 6604 916 6612 924
rect 1244 896 1252 904
rect 1340 896 1348 904
rect 1356 896 1364 904
rect 1420 896 1428 904
rect 1580 896 1588 904
rect 1724 896 1732 904
rect 1820 896 1828 904
rect 1980 896 1988 904
rect 156 876 164 884
rect 220 876 228 884
rect 428 876 436 884
rect 748 876 756 884
rect 828 876 836 884
rect 876 876 884 884
rect 940 876 948 884
rect 1068 876 1076 884
rect 1308 876 1316 884
rect 236 856 244 864
rect 1628 876 1636 884
rect 1676 876 1684 884
rect 1756 876 1764 884
rect 1788 876 1796 884
rect 1868 876 1876 884
rect 1948 876 1956 884
rect 1980 876 1988 884
rect 2108 896 2116 904
rect 2172 896 2180 904
rect 2188 896 2196 904
rect 2268 896 2276 904
rect 2380 896 2388 904
rect 2412 896 2420 904
rect 2476 896 2484 904
rect 2780 896 2788 904
rect 2812 896 2820 904
rect 2892 896 2900 904
rect 3388 896 3396 904
rect 3532 896 3540 904
rect 3820 896 3828 904
rect 3900 896 3908 904
rect 3996 896 4004 904
rect 4124 896 4132 904
rect 4332 896 4340 904
rect 4604 896 4612 904
rect 4700 896 4708 904
rect 4732 896 4740 904
rect 4812 896 4820 904
rect 4956 896 4964 904
rect 5116 896 5124 904
rect 5148 896 5156 904
rect 5340 896 5348 904
rect 5532 896 5540 904
rect 5628 896 5636 904
rect 5676 896 5684 904
rect 5740 896 5748 904
rect 5868 896 5876 904
rect 5948 896 5956 904
rect 5964 896 5972 904
rect 6028 896 6036 904
rect 6092 896 6100 904
rect 6156 896 6164 904
rect 6188 896 6196 904
rect 6252 896 6260 904
rect 6316 896 6324 904
rect 6492 896 6500 904
rect 2028 876 2036 884
rect 2060 876 2068 884
rect 2076 876 2084 884
rect 2140 876 2148 884
rect 2748 876 2756 884
rect 2988 876 2996 884
rect 3100 876 3108 884
rect 3196 876 3204 884
rect 3244 876 3252 884
rect 3356 876 3364 884
rect 3452 876 3460 884
rect 3516 876 3524 884
rect 3564 876 3572 884
rect 4060 876 4068 884
rect 4092 876 4100 884
rect 4764 876 4772 884
rect 4924 876 4932 884
rect 5804 876 5812 884
rect 5996 876 6004 884
rect 6060 876 6068 884
rect 6124 876 6132 884
rect 6220 876 6228 884
rect 6284 876 6292 884
rect 6348 876 6356 884
rect 6380 876 6388 884
rect 6524 876 6532 884
rect 6556 876 6564 884
rect 2012 856 2020 864
rect 300 836 308 844
rect 508 836 516 844
rect 588 836 596 844
rect 684 836 692 844
rect 732 836 740 844
rect 812 836 820 844
rect 860 836 868 844
rect 924 836 932 844
rect 1084 836 1092 844
rect 1212 836 1220 844
rect 1292 836 1300 844
rect 1564 836 1572 844
rect 1612 836 1620 844
rect 1692 836 1700 844
rect 1740 836 1748 844
rect 1916 836 1924 844
rect 2124 836 2132 844
rect 2252 836 2260 844
rect 2508 836 2516 844
rect 2572 836 2580 844
rect 2668 836 2676 844
rect 2796 836 2804 844
rect 2876 836 2884 844
rect 3004 836 3012 844
rect 3116 836 3124 844
rect 3260 836 3268 844
rect 3372 836 3380 844
rect 3436 836 3444 844
rect 3772 836 3780 844
rect 3804 836 3812 844
rect 3884 836 3892 844
rect 3932 836 3940 844
rect 4108 836 4116 844
rect 5404 836 5412 844
rect 5852 836 5860 844
rect 5932 836 5940 844
rect 5980 836 5988 844
rect 6044 836 6052 844
rect 6236 836 6244 844
rect 6332 836 6340 844
rect 6460 836 6468 844
rect 6540 836 6548 844
rect 1774 806 1782 814
rect 1788 806 1796 814
rect 1802 806 1810 814
rect 4830 806 4838 814
rect 4844 806 4852 814
rect 4858 806 4866 814
rect 28 776 36 784
rect 76 776 84 784
rect 156 776 164 784
rect 252 776 260 784
rect 412 776 420 784
rect 476 776 484 784
rect 556 776 564 784
rect 1532 776 1540 784
rect 1932 776 1940 784
rect 1996 776 2004 784
rect 2476 776 2484 784
rect 4412 776 4420 784
rect 4604 776 4612 784
rect 5020 776 5028 784
rect 5180 776 5188 784
rect 5292 776 5300 784
rect 5708 776 5716 784
rect 5740 776 5748 784
rect 6108 776 6116 784
rect 6348 776 6356 784
rect 652 756 660 764
rect 1468 756 1476 764
rect 92 736 100 744
rect 236 736 244 744
rect 428 736 436 744
rect 492 736 500 744
rect 572 736 580 744
rect 604 736 612 744
rect 668 736 676 744
rect 700 736 708 744
rect 1228 736 1236 744
rect 1260 736 1268 744
rect 1372 736 1380 744
rect 1420 736 1428 744
rect 1484 736 1492 744
rect 1516 736 1524 744
rect 1612 736 1620 744
rect 1916 736 1924 744
rect 1948 736 1956 744
rect 2012 736 2020 744
rect 3068 736 3076 744
rect 3196 736 3204 744
rect 4044 736 4052 744
rect 4892 736 4900 744
rect 4972 736 4980 744
rect 5036 736 5044 744
rect 5164 736 5172 744
rect 5964 736 5972 744
rect 6092 736 6100 744
rect 6492 736 6500 744
rect 60 716 68 724
rect 124 716 132 724
rect 188 716 196 724
rect 220 716 228 724
rect 300 716 308 724
rect 460 716 468 724
rect 524 716 532 724
rect 540 716 548 724
rect 1068 716 1076 724
rect 1084 716 1092 724
rect 1196 716 1204 724
rect 1340 716 1348 724
rect 1404 716 1412 724
rect 1452 716 1460 724
rect 1516 716 1524 724
rect 1580 716 1588 724
rect 1692 716 1700 724
rect 1788 716 1796 724
rect 1916 716 1924 724
rect 1980 716 1988 724
rect 2044 716 2052 724
rect 2252 716 2260 724
rect 2364 716 2372 724
rect 2460 716 2468 724
rect 2620 716 2628 724
rect 2732 716 2740 724
rect 2876 716 2884 724
rect 3036 716 3044 724
rect 3164 716 3172 724
rect 3228 716 3236 724
rect 3468 716 3476 724
rect 3548 716 3556 724
rect 3612 716 3620 724
rect 3676 716 3684 724
rect 3692 716 3700 724
rect 3772 716 3780 724
rect 3804 716 3812 724
rect 28 696 36 704
rect 108 696 116 704
rect 156 696 164 704
rect 252 696 260 704
rect 348 696 356 704
rect 444 696 452 704
rect 508 696 516 704
rect 556 696 564 704
rect 652 696 660 704
rect 956 696 964 704
rect 1036 696 1044 704
rect 1148 696 1156 704
rect 1212 696 1220 704
rect 1308 696 1316 704
rect 1388 696 1396 704
rect 1468 696 1476 704
rect 1532 696 1540 704
rect 1596 696 1604 704
rect 1756 696 1764 704
rect 1900 696 1908 704
rect 1932 696 1940 704
rect 1996 696 2004 704
rect 2076 696 2084 704
rect 2268 696 2276 704
rect 2348 696 2356 704
rect 2476 696 2484 704
rect 2604 696 2612 704
rect 2652 696 2660 704
rect 12 676 20 684
rect 140 676 148 684
rect 204 676 212 684
rect 332 676 340 684
rect 364 676 372 684
rect 828 676 836 684
rect 940 676 948 684
rect 972 676 980 684
rect 1020 676 1028 684
rect 1084 676 1092 684
rect 1116 676 1124 684
rect 1132 676 1140 684
rect 1292 676 1300 684
rect 1644 676 1652 684
rect 1724 676 1732 684
rect 1836 676 1844 684
rect 1884 676 1892 684
rect 2092 676 2100 684
rect 2108 676 2116 684
rect 2204 676 2212 684
rect 2220 676 2228 684
rect 2252 676 2260 684
rect 2396 676 2404 684
rect 2412 676 2420 684
rect 2444 676 2452 684
rect 220 656 228 664
rect 396 656 404 664
rect 604 656 612 664
rect 700 656 708 664
rect 1004 656 1012 664
rect 1260 656 1268 664
rect 1340 656 1348 664
rect 1420 656 1428 664
rect 1852 656 1860 664
rect 2300 656 2308 664
rect 2316 656 2324 664
rect 2364 656 2372 664
rect 2508 656 2516 664
rect 2556 676 2564 684
rect 2588 676 2596 684
rect 2604 676 2612 684
rect 2668 676 2676 684
rect 2700 696 2708 704
rect 2796 696 2804 704
rect 2892 696 2900 704
rect 2972 696 2980 704
rect 3052 696 3060 704
rect 3148 696 3156 704
rect 3180 696 3188 704
rect 3260 696 3268 704
rect 3580 696 3588 704
rect 3948 716 3956 724
rect 4028 716 4036 724
rect 4156 716 4164 724
rect 4460 716 4468 724
rect 4540 716 4548 724
rect 4636 716 4644 724
rect 4652 716 4660 724
rect 4732 716 4740 724
rect 4780 716 4788 724
rect 4908 716 4916 724
rect 4956 716 4964 724
rect 5004 716 5012 724
rect 5068 716 5076 724
rect 5468 716 5476 724
rect 5548 716 5556 724
rect 5580 716 5588 724
rect 5644 716 5652 724
rect 5772 716 5780 724
rect 5996 716 6004 724
rect 6124 716 6132 724
rect 6380 716 6388 724
rect 6460 716 6468 724
rect 6524 716 6532 724
rect 6556 716 6564 724
rect 6572 716 6580 724
rect 4108 696 4116 704
rect 4220 696 4228 704
rect 4252 696 4260 704
rect 4348 696 4356 704
rect 4380 696 4388 704
rect 4508 696 4516 704
rect 4604 696 4612 704
rect 4844 696 4852 704
rect 4892 696 4900 704
rect 4924 696 4932 704
rect 5020 696 5028 704
rect 5164 696 5172 704
rect 5228 696 5236 704
rect 5372 696 5380 704
rect 5436 696 5444 704
rect 5500 696 5508 704
rect 5612 696 5620 704
rect 5820 696 5828 704
rect 5980 696 5988 704
rect 6028 696 6036 704
rect 6060 696 6068 704
rect 6108 696 6116 704
rect 6188 696 6196 704
rect 6252 696 6260 704
rect 6348 696 6356 704
rect 6380 696 6388 704
rect 6444 696 6452 704
rect 6476 696 6484 704
rect 2780 676 2788 684
rect 2844 676 2852 684
rect 2924 676 2932 684
rect 3084 676 3092 684
rect 3132 676 3140 684
rect 3244 676 3252 684
rect 3276 676 3284 684
rect 3500 676 3508 684
rect 3516 676 3524 684
rect 3564 676 3572 684
rect 3628 676 3636 684
rect 3644 676 3652 684
rect 3660 676 3668 684
rect 3724 676 3732 684
rect 3772 676 3780 684
rect 3980 676 3988 684
rect 4124 676 4132 684
rect 4332 676 4340 684
rect 4364 676 4372 684
rect 4428 676 4436 684
rect 4524 676 4532 684
rect 4572 676 4580 684
rect 4588 676 4596 684
rect 4684 676 4692 684
rect 4700 676 4708 684
rect 4732 676 4740 684
rect 4748 676 4756 684
rect 4828 676 4836 684
rect 5100 676 5108 684
rect 5196 676 5204 684
rect 2556 656 2564 664
rect 2748 656 2756 664
rect 2764 656 2772 664
rect 2956 656 2964 664
rect 3020 656 3028 664
rect 3100 656 3108 664
rect 3356 656 3364 664
rect 3708 656 3716 664
rect 3884 656 3892 664
rect 4060 656 4068 664
rect 4076 656 4084 664
rect 4108 656 4116 664
rect 4172 656 4180 664
rect 4268 656 4276 664
rect 4460 656 4468 664
rect 4796 656 4804 664
rect 4988 656 4996 664
rect 5116 656 5124 664
rect 5212 656 5220 664
rect 5260 676 5268 684
rect 5308 676 5316 684
rect 5372 676 5380 684
rect 5404 676 5412 684
rect 5548 676 5556 684
rect 5644 676 5652 684
rect 5676 676 5684 684
rect 5756 676 5764 684
rect 5788 676 5796 684
rect 5804 676 5812 684
rect 5276 656 5284 664
rect 5404 656 5412 664
rect 5660 656 5668 664
rect 5820 656 5828 664
rect 5852 656 5860 664
rect 5932 676 5940 684
rect 6044 676 6052 684
rect 6172 676 6180 684
rect 6188 676 6196 684
rect 6236 676 6244 684
rect 6332 676 6340 684
rect 6428 676 6436 684
rect 6524 676 6532 684
rect 6604 676 6612 684
rect 6012 656 6020 664
rect 6140 656 6148 664
rect 6220 656 6228 664
rect 6396 656 6404 664
rect 300 636 308 644
rect 380 636 388 644
rect 764 636 772 644
rect 876 636 884 644
rect 988 636 996 644
rect 1084 636 1092 644
rect 1180 636 1188 644
rect 1212 636 1220 644
rect 1276 636 1284 644
rect 1356 636 1364 644
rect 1596 636 1604 644
rect 1660 636 1668 644
rect 1692 636 1700 644
rect 2044 636 2052 644
rect 2140 636 2148 644
rect 2236 636 2244 644
rect 2348 636 2356 644
rect 2396 636 2404 644
rect 2572 636 2580 644
rect 2780 636 2788 644
rect 3004 636 3012 644
rect 3116 636 3124 644
rect 3180 636 3188 644
rect 3372 636 3380 644
rect 3468 636 3476 644
rect 3548 636 3556 644
rect 3612 636 3620 644
rect 3644 636 3652 644
rect 3788 636 3796 644
rect 3820 636 3828 644
rect 3932 636 3940 644
rect 3948 636 3956 644
rect 4012 636 4020 644
rect 4156 636 4164 644
rect 4188 636 4196 644
rect 4316 636 4324 644
rect 4476 636 4484 644
rect 4556 636 4564 644
rect 4652 636 4660 644
rect 4780 636 4788 644
rect 4812 636 4820 644
rect 4940 636 4948 644
rect 5084 636 5092 644
rect 5132 636 5140 644
rect 5164 636 5172 644
rect 5196 636 5204 644
rect 5436 636 5444 644
rect 5548 636 5556 644
rect 5564 636 5572 644
rect 5884 636 5892 644
rect 5916 636 5924 644
rect 5948 636 5956 644
rect 6108 636 6116 644
rect 6156 636 6164 644
rect 6268 636 6276 644
rect 6540 636 6548 644
rect 6572 636 6580 644
rect 2316 616 2324 624
rect 5276 616 5284 624
rect 5324 616 5332 624
rect 5404 616 5412 624
rect 3310 606 3318 614
rect 3324 606 3332 614
rect 3338 606 3346 614
rect 4700 596 4708 604
rect 4972 596 4980 604
rect 5836 596 5844 604
rect 60 576 68 584
rect 236 576 244 584
rect 316 576 324 584
rect 556 576 564 584
rect 2044 576 2052 584
rect 2620 576 2628 584
rect 3532 576 3540 584
rect 3596 576 3604 584
rect 4172 576 4180 584
rect 4620 576 4628 584
rect 5180 576 5188 584
rect 5356 576 5364 584
rect 5452 576 5460 584
rect 5596 576 5604 584
rect 6012 576 6020 584
rect 188 556 196 564
rect 252 556 260 564
rect 332 556 340 564
rect 540 556 548 564
rect 1228 556 1236 564
rect 1484 556 1492 564
rect 1628 556 1636 564
rect 1996 556 2004 564
rect 12 536 20 544
rect 108 536 116 544
rect 140 536 148 544
rect 204 536 212 544
rect 300 536 308 544
rect 364 536 372 544
rect 572 536 580 544
rect 588 536 596 544
rect 700 536 708 544
rect 972 536 980 544
rect 1068 536 1076 544
rect 1132 536 1140 544
rect 1452 536 1460 544
rect 1660 536 1668 544
rect 1868 536 1876 544
rect 2012 536 2020 544
rect 2108 536 2116 544
rect 2124 536 2132 544
rect 2220 536 2228 544
rect 2604 556 2612 564
rect 2812 556 2820 564
rect 2892 556 2900 564
rect 3148 556 3156 564
rect 3164 556 3172 564
rect 3196 556 3204 564
rect 3228 556 3236 564
rect 3260 556 3268 564
rect 4204 556 4212 564
rect 4300 556 4308 564
rect 4316 556 4324 564
rect 4364 556 4372 564
rect 4668 556 4676 564
rect 4684 556 4692 564
rect 4700 556 4708 564
rect 4716 556 4724 564
rect 4764 556 4772 564
rect 4812 556 4820 564
rect 4972 556 4980 564
rect 5036 556 5044 564
rect 5292 556 5300 564
rect 5308 556 5316 564
rect 5340 556 5348 564
rect 5372 556 5380 564
rect 5484 556 5492 564
rect 5500 556 5508 564
rect 5740 556 5748 564
rect 6108 556 6116 564
rect 6236 556 6244 564
rect 6300 556 6308 564
rect 2268 536 2276 544
rect 2300 536 2308 544
rect 2428 536 2436 544
rect 2460 536 2468 544
rect 2524 536 2532 544
rect 2684 536 2692 544
rect 2748 536 2756 544
rect 2812 536 2820 544
rect 2844 536 2852 544
rect 2956 536 2964 544
rect 3340 536 3348 544
rect 3420 536 3428 544
rect 3452 536 3460 544
rect 3468 536 3476 544
rect 3532 536 3540 544
rect 3548 536 3556 544
rect 3628 536 3636 544
rect 3692 536 3700 544
rect 3708 536 3716 544
rect 3772 536 3780 544
rect 3836 536 3844 544
rect 3900 536 3908 544
rect 4156 536 4164 544
rect 4332 536 4340 544
rect 4396 536 4404 544
rect 4540 536 4548 544
rect 4652 536 4660 544
rect 4908 536 4916 544
rect 5004 536 5012 544
rect 284 516 292 524
rect 364 516 372 524
rect 444 516 452 524
rect 508 516 516 524
rect 588 516 596 524
rect 604 516 612 524
rect 748 516 756 524
rect 796 516 804 524
rect 860 516 868 524
rect 940 516 948 524
rect 124 496 132 504
rect 236 496 244 504
rect 348 496 356 504
rect 460 496 468 504
rect 524 496 532 504
rect 764 496 772 504
rect 780 496 788 504
rect 844 496 852 504
rect 956 496 964 504
rect 1052 516 1060 524
rect 1100 516 1108 524
rect 1116 516 1124 524
rect 1180 516 1188 524
rect 1260 516 1268 524
rect 1340 516 1348 524
rect 1388 516 1396 524
rect 1436 516 1444 524
rect 1516 516 1524 524
rect 1596 516 1604 524
rect 1676 516 1684 524
rect 1708 516 1716 524
rect 1836 516 1844 524
rect 2380 516 2388 524
rect 2508 516 2516 524
rect 2556 516 2564 524
rect 2604 516 2612 524
rect 2652 516 2660 524
rect 2668 516 2676 524
rect 2732 516 2740 524
rect 2860 516 2868 524
rect 2940 516 2948 524
rect 2988 516 2996 524
rect 3052 516 3060 524
rect 3196 516 3204 524
rect 3324 516 3332 524
rect 3356 516 3364 524
rect 3404 516 3412 524
rect 3468 516 3476 524
rect 3484 516 3492 524
rect 3548 516 3556 524
rect 3564 516 3572 524
rect 3628 516 3636 524
rect 3676 516 3684 524
rect 3724 516 3732 524
rect 3788 516 3796 524
rect 3836 516 3844 524
rect 3852 516 3860 524
rect 3900 516 3908 524
rect 3996 516 4004 524
rect 4060 516 4068 524
rect 4124 516 4132 524
rect 4220 516 4228 524
rect 4268 516 4276 524
rect 4348 516 4356 524
rect 4380 516 4388 524
rect 4412 516 4420 524
rect 4444 516 4452 524
rect 4524 516 4532 524
rect 4556 516 4564 524
rect 4668 516 4676 524
rect 4748 516 4756 524
rect 4796 516 4804 524
rect 4924 516 4932 524
rect 5068 516 5076 524
rect 5084 516 5092 524
rect 5116 536 5124 544
rect 5356 536 5364 544
rect 5420 536 5428 544
rect 5516 536 5524 544
rect 5596 536 5604 544
rect 5708 536 5716 544
rect 5740 536 5748 544
rect 5820 536 5828 544
rect 5884 536 5892 544
rect 5948 536 5956 544
rect 5964 536 5972 544
rect 6188 536 6196 544
rect 6204 536 6212 544
rect 6236 536 6244 544
rect 6444 536 6452 544
rect 5132 516 5140 524
rect 5212 516 5220 524
rect 5404 516 5412 524
rect 5596 516 5604 524
rect 5660 516 5668 524
rect 5692 516 5700 524
rect 5836 516 5844 524
rect 5884 516 5892 524
rect 5916 516 5924 524
rect 5948 516 5956 524
rect 5980 516 5988 524
rect 6060 516 6068 524
rect 6156 516 6164 524
rect 6188 516 6196 524
rect 6316 516 6324 524
rect 6444 516 6452 524
rect 6556 516 6564 524
rect 1020 496 1028 504
rect 1084 496 1092 504
rect 1196 496 1204 504
rect 1244 496 1252 504
rect 1372 496 1380 504
rect 1500 496 1508 504
rect 1612 496 1620 504
rect 1692 496 1700 504
rect 1852 496 1860 504
rect 2268 496 2276 504
rect 2300 496 2308 504
rect 2316 496 2324 504
rect 2364 496 2372 504
rect 2428 496 2436 504
rect 2476 496 2484 504
rect 2540 496 2548 504
rect 2636 496 2644 504
rect 2700 496 2708 504
rect 2764 496 2772 504
rect 2876 496 2884 504
rect 2892 496 2900 504
rect 2972 496 2980 504
rect 3036 496 3044 504
rect 3644 496 3652 504
rect 3756 496 3764 504
rect 3820 496 3828 504
rect 3884 496 3892 504
rect 3916 496 3924 504
rect 3948 496 3956 504
rect 4012 496 4020 504
rect 4076 496 4084 504
rect 4140 496 4148 504
rect 4188 496 4196 504
rect 4284 496 4292 504
rect 4428 496 4436 504
rect 4492 496 4500 504
rect 4956 496 4964 504
rect 5052 496 5060 504
rect 5132 496 5140 504
rect 5164 496 5172 504
rect 5180 496 5188 504
rect 5244 496 5252 504
rect 5324 496 5332 504
rect 5612 496 5620 504
rect 5676 496 5684 504
rect 5756 496 5764 504
rect 5868 496 5876 504
rect 6076 496 6084 504
rect 6124 496 6132 504
rect 268 476 276 484
rect 380 476 388 484
rect 412 476 420 484
rect 428 476 436 484
rect 492 476 500 484
rect 812 476 820 484
rect 876 476 884 484
rect 924 476 932 484
rect 1164 476 1172 484
rect 1180 476 1188 484
rect 1276 476 1284 484
rect 1324 476 1332 484
rect 1340 476 1348 484
rect 1404 476 1412 484
rect 1532 476 1540 484
rect 1580 476 1588 484
rect 1692 476 1700 484
rect 1820 476 1828 484
rect 1900 476 1908 484
rect 2396 476 2404 484
rect 2572 476 2580 484
rect 2732 476 2740 484
rect 2796 476 2804 484
rect 3004 476 3012 484
rect 3068 476 3076 484
rect 3420 476 3428 484
rect 3980 476 3988 484
rect 4044 476 4052 484
rect 4108 476 4116 484
rect 4252 476 4260 484
rect 4460 476 4468 484
rect 5004 476 5012 484
rect 5276 476 5284 484
rect 5548 476 5556 484
rect 5580 476 5588 484
rect 5644 476 5652 484
rect 508 456 516 464
rect 2556 456 2564 464
rect 3052 456 3060 464
rect 3244 456 3252 464
rect 3724 456 3732 464
rect 4268 456 4276 464
rect 716 436 724 444
rect 796 436 804 444
rect 860 436 868 444
rect 908 436 916 444
rect 988 436 996 444
rect 1148 436 1156 444
rect 1260 436 1268 444
rect 1308 436 1316 444
rect 1388 436 1396 444
rect 1484 436 1492 444
rect 1516 436 1524 444
rect 1596 436 1604 444
rect 1628 436 1636 444
rect 1708 436 1716 444
rect 1836 436 1844 444
rect 2156 436 2164 444
rect 2284 436 2292 444
rect 2380 436 2388 444
rect 2812 436 2820 444
rect 2940 436 2948 444
rect 2988 436 2996 444
rect 3100 436 3108 444
rect 3196 436 3204 444
rect 3676 436 3684 444
rect 3852 436 3860 444
rect 3996 436 4004 444
rect 4028 436 4036 444
rect 4124 436 4132 444
rect 4476 436 4484 444
rect 4524 436 4532 444
rect 4732 436 4740 444
rect 4796 436 4804 444
rect 4828 436 4836 444
rect 4924 436 4932 444
rect 5404 436 5412 444
rect 5660 436 5668 444
rect 5740 436 5748 444
rect 5836 436 5844 444
rect 6060 436 6068 444
rect 6156 436 6164 444
rect 6428 436 6436 444
rect 6620 436 6628 444
rect 1774 406 1782 414
rect 1788 406 1796 414
rect 1802 406 1810 414
rect 4830 406 4838 414
rect 4844 406 4852 414
rect 4858 406 4866 414
rect 12 376 20 384
rect 156 376 164 384
rect 220 376 228 384
rect 284 376 292 384
rect 476 376 484 384
rect 1388 376 1396 384
rect 1628 376 1636 384
rect 2732 376 2740 384
rect 3292 376 3300 384
rect 3420 376 3428 384
rect 4348 376 4356 384
rect 5100 376 5108 384
rect 5628 376 5636 384
rect 5724 376 5732 384
rect 5804 376 5812 384
rect 6012 376 6020 384
rect 6412 376 6420 384
rect 6604 376 6612 384
rect 140 336 148 344
rect 204 336 212 344
rect 380 356 388 364
rect 572 356 580 364
rect 348 336 356 344
rect 396 336 404 344
rect 556 336 564 344
rect 588 336 596 344
rect 652 336 660 344
rect 668 336 676 344
rect 1068 356 1076 364
rect 1692 356 1700 364
rect 1868 356 1876 364
rect 2092 356 2100 364
rect 2476 356 2484 364
rect 2812 356 2820 364
rect 3468 356 3476 364
rect 3596 356 3604 364
rect 3948 356 3956 364
rect 732 336 740 344
rect 796 336 804 344
rect 956 336 964 344
rect 1324 336 1332 344
rect 1340 336 1348 344
rect 1404 336 1412 344
rect 1612 336 1620 344
rect 1708 336 1716 344
rect 1756 336 1764 344
rect 1852 336 1860 344
rect 2076 336 2084 344
rect 2364 336 2372 344
rect 2460 336 2468 344
rect 2716 336 2724 344
rect 2796 336 2804 344
rect 2860 336 2868 344
rect 3100 336 3108 344
rect 3132 336 3140 344
rect 3276 336 3284 344
rect 3404 336 3412 344
rect 3452 336 3460 344
rect 3532 336 3540 344
rect 3580 336 3588 344
rect 3900 336 3908 344
rect 3964 336 3972 344
rect 4172 336 4180 344
rect 4220 336 4228 344
rect 4284 336 4292 344
rect 4300 336 4308 344
rect 4396 336 4404 344
rect 4588 336 4596 344
rect 5820 336 5828 344
rect 6012 336 6020 344
rect 6028 336 6036 344
rect 76 316 84 324
rect 172 316 180 324
rect 236 316 244 324
rect 268 316 276 324
rect 300 316 308 324
rect 316 316 324 324
rect 428 316 436 324
rect 460 316 468 324
rect 492 316 500 324
rect 556 316 564 324
rect 620 316 628 324
rect 684 316 692 324
rect 700 316 708 324
rect 764 316 772 324
rect 828 316 836 324
rect 876 316 884 324
rect 1036 316 1044 324
rect 1100 316 1108 324
rect 1212 316 1220 324
rect 1260 316 1268 324
rect 1372 316 1380 324
rect 1436 316 1444 324
rect 1644 316 1652 324
rect 1708 316 1716 324
rect 1724 316 1732 324
rect 1884 316 1892 324
rect 2012 316 2020 324
rect 2028 316 2036 324
rect 2108 316 2116 324
rect 2188 316 2196 324
rect 2284 316 2292 324
rect 2492 316 2500 324
rect 2572 316 2580 324
rect 2748 316 2756 324
rect 2828 316 2836 324
rect 156 296 164 304
rect 220 296 228 304
rect 284 296 292 304
rect 332 296 340 304
rect 412 296 420 304
rect 476 296 484 304
rect 540 296 548 304
rect 604 296 612 304
rect 668 296 676 304
rect 716 296 724 304
rect 780 296 788 304
rect 908 296 916 304
rect 924 296 932 304
rect 972 296 980 304
rect 1068 296 1076 304
rect 1196 296 1204 304
rect 1340 296 1348 304
rect 1388 296 1396 304
rect 1484 296 1492 304
rect 1580 296 1588 304
rect 1628 296 1636 304
rect 1692 296 1700 304
rect 1740 296 1748 304
rect 1868 296 1876 304
rect 2092 296 2100 304
rect 2124 296 2132 304
rect 2252 296 2260 304
rect 2476 296 2484 304
rect 2508 296 2516 304
rect 2572 296 2580 304
rect 2604 296 2612 304
rect 2684 296 2692 304
rect 2732 296 2740 304
rect 2780 296 2788 304
rect 2860 296 2868 304
rect 2956 316 2964 324
rect 3116 316 3124 324
rect 3308 316 3316 324
rect 3484 316 3492 324
rect 3612 316 3620 324
rect 3628 316 3636 324
rect 3644 316 3652 324
rect 3756 316 3764 324
rect 3804 316 3812 324
rect 3868 316 3876 324
rect 3932 316 3940 324
rect 4028 316 4036 324
rect 4124 316 4132 324
rect 4140 316 4148 324
rect 4252 316 4260 324
rect 4268 316 4276 324
rect 4428 316 4436 324
rect 4540 316 4548 324
rect 4556 316 4564 324
rect 4780 316 4788 324
rect 5036 316 5044 324
rect 5180 316 5188 324
rect 5276 316 5284 324
rect 5292 316 5300 324
rect 3004 296 3012 304
rect 3100 296 3108 304
rect 3148 296 3156 304
rect 3244 296 3252 304
rect 3292 296 3300 304
rect 3388 296 3396 304
rect 3468 296 3476 304
rect 3516 296 3524 304
rect 3596 296 3604 304
rect 3660 296 3668 304
rect 3724 296 3732 304
rect 3852 296 3860 304
rect 3884 296 3892 304
rect 3948 296 3956 304
rect 4076 296 4084 304
rect 4156 296 4164 304
rect 4188 296 4196 304
rect 4236 296 4244 304
rect 4284 296 4292 304
rect 4332 296 4340 304
rect 4412 296 4420 304
rect 4572 296 4580 304
rect 4652 296 4660 304
rect 4732 296 4740 304
rect 4956 296 4964 304
rect 5244 296 5252 304
rect 5388 296 5396 304
rect 44 276 52 284
rect 108 276 116 284
rect 924 276 932 284
rect 1084 276 1092 284
rect 1132 276 1140 284
rect 1148 276 1156 284
rect 1212 276 1220 284
rect 1244 276 1252 284
rect 1292 276 1300 284
rect 1500 276 1508 284
rect 1516 276 1524 284
rect 1564 276 1572 284
rect 1820 276 1828 284
rect 1900 276 1908 284
rect 1996 276 2004 284
rect 2044 276 2052 284
rect 2140 276 2148 284
rect 2172 276 2180 284
rect 2284 276 2292 284
rect 2316 276 2324 284
rect 2332 276 2340 284
rect 2428 276 2436 284
rect 2524 276 2532 284
rect 2620 276 2628 284
rect 2668 276 2676 284
rect 2876 276 2884 284
rect 2940 276 2948 284
rect 2956 276 2964 284
rect 2988 276 2996 284
rect 3020 276 3028 284
rect 3228 276 3236 284
rect 3660 276 3668 284
rect 3708 276 3716 284
rect 3772 276 3780 284
rect 3804 276 3812 284
rect 4060 276 4068 284
rect 4092 276 4100 284
rect 4108 276 4116 284
rect 4236 276 4244 284
rect 4332 276 4340 284
rect 4460 276 4468 284
rect 4508 276 4516 284
rect 4652 276 4660 284
rect 4684 276 4692 284
rect 4716 276 4724 284
rect 5452 294 5460 302
rect 5516 296 5524 304
rect 5724 296 5732 304
rect 5788 316 5796 324
rect 5932 316 5940 324
rect 5996 316 6004 324
rect 6124 316 6132 324
rect 5772 296 5780 304
rect 5804 296 5812 304
rect 5852 296 5860 304
rect 6012 296 6020 304
rect 6108 296 6116 304
rect 6284 296 6292 304
rect 6396 296 6404 304
rect 6476 296 6484 304
rect 6524 296 6532 304
rect 4764 276 4772 284
rect 5068 276 5076 284
rect 5148 276 5156 284
rect 5212 276 5220 284
rect 5228 276 5236 284
rect 5308 276 5316 284
rect 5324 276 5332 284
rect 5372 276 5380 284
rect 5612 276 5620 284
rect 5660 276 5668 284
rect 12 256 20 264
rect 780 256 788 264
rect 1020 256 1028 264
rect 1100 256 1108 264
rect 1148 256 1156 264
rect 1532 256 1540 264
rect 1548 256 1556 264
rect 2204 256 2212 264
rect 2556 256 2564 264
rect 2572 256 2580 264
rect 2636 256 2644 264
rect 3052 256 3060 264
rect 3180 256 3188 264
rect 3196 256 3204 264
rect 3692 256 3700 264
rect 3820 256 3828 264
rect 3996 256 4004 264
rect 4492 256 4500 264
rect 4540 256 4548 264
rect 4972 256 4980 264
rect 5084 256 5092 264
rect 5164 256 5172 264
rect 5276 256 5284 264
rect 5340 256 5348 264
rect 5356 256 5364 264
rect 5596 256 5604 264
rect 5676 256 5684 264
rect 5772 276 5780 284
rect 5868 276 5876 284
rect 5836 256 5844 264
rect 5900 256 5908 264
rect 6092 276 6100 284
rect 6156 276 6164 284
rect 6300 276 6308 284
rect 5964 256 5972 264
rect 6060 256 6068 264
rect 6620 256 6628 264
rect 92 236 100 244
rect 636 236 644 244
rect 828 236 836 244
rect 1212 236 1220 244
rect 1260 236 1268 244
rect 1308 236 1316 244
rect 1436 236 1444 244
rect 1932 236 1940 244
rect 2220 236 2228 244
rect 2284 236 2292 244
rect 2652 236 2660 244
rect 3036 236 3044 244
rect 3084 236 3092 244
rect 3212 236 3220 244
rect 3260 236 3268 244
rect 3548 236 3556 244
rect 3756 236 3764 244
rect 3788 236 3796 244
rect 3884 236 3892 244
rect 4476 236 4484 244
rect 4620 236 4628 244
rect 4684 236 4692 244
rect 4844 236 4852 244
rect 5036 236 5044 244
rect 5068 236 5076 244
rect 5116 236 5124 244
rect 5180 236 5188 244
rect 5324 236 5332 244
rect 5580 236 5588 244
rect 6076 236 6084 244
rect 6124 236 6132 244
rect 6172 236 6180 244
rect 6364 236 6372 244
rect 3310 206 3318 214
rect 3324 206 3332 214
rect 3338 206 3346 214
rect 76 176 84 184
rect 156 176 164 184
rect 364 176 372 184
rect 428 176 436 184
rect 492 176 500 184
rect 1260 176 1268 184
rect 2588 176 2596 184
rect 3116 176 3124 184
rect 3228 176 3236 184
rect 4124 176 4132 184
rect 5004 176 5012 184
rect 6076 176 6084 184
rect 6156 176 6164 184
rect 6332 176 6340 184
rect 6412 176 6420 184
rect 6492 176 6500 184
rect 6556 176 6564 184
rect 12 156 20 164
rect 92 136 100 144
rect 188 136 196 144
rect 220 136 228 144
rect 236 136 244 144
rect 268 156 276 164
rect 444 156 452 164
rect 892 156 900 164
rect 1068 156 1076 164
rect 1164 156 1172 164
rect 1292 156 1300 164
rect 1404 156 1412 164
rect 1612 156 1620 164
rect 2012 156 2020 164
rect 2300 156 2308 164
rect 2524 156 2532 164
rect 2604 156 2612 164
rect 3708 156 3716 164
rect 300 136 308 144
rect 412 136 420 144
rect 460 136 468 144
rect 716 136 724 144
rect 844 136 852 144
rect 1004 136 1012 144
rect 1020 136 1028 144
rect 1036 136 1044 144
rect 1100 136 1108 144
rect 1196 136 1204 144
rect 1260 136 1268 144
rect 1388 136 1396 144
rect 1484 136 1492 144
rect 1564 136 1572 144
rect 1580 136 1588 144
rect 1676 136 1684 144
rect 1948 136 1956 144
rect 2028 136 2036 144
rect 2156 136 2164 144
rect 2252 136 2260 144
rect 2524 136 2532 144
rect 2556 136 2564 144
rect 2764 136 2772 144
rect 2796 136 2804 144
rect 2844 136 2852 144
rect 2876 136 2884 144
rect 2924 136 2932 144
rect 2956 136 2964 144
rect 3004 136 3012 144
rect 3036 136 3044 144
rect 3068 136 3076 144
rect 3132 136 3140 144
rect 3420 136 3428 144
rect 3676 136 3684 144
rect 3804 156 3812 164
rect 3868 156 3876 164
rect 4876 156 4884 164
rect 5660 156 5668 164
rect 6028 156 6036 164
rect 3772 136 3780 144
rect 3788 136 3796 144
rect 3836 136 3844 144
rect 3868 136 3876 144
rect 3996 136 4004 144
rect 4012 136 4020 144
rect 4156 136 4164 144
rect 4428 136 4436 144
rect 4668 136 4676 144
rect 4700 136 4708 144
rect 4796 136 4804 144
rect 4876 136 4884 144
rect 4972 136 4980 144
rect 5020 136 5028 144
rect 5052 136 5060 144
rect 5308 136 5316 144
rect 5420 136 5428 144
rect 5788 136 5796 144
rect 5884 136 5892 144
rect 5916 136 5924 144
rect 6012 136 6020 144
rect 6044 136 6052 144
rect 6124 136 6132 144
rect 6508 136 6516 144
rect 6524 136 6532 144
rect 6620 136 6628 144
rect 204 116 212 124
rect 316 116 324 124
rect 364 116 372 124
rect 396 116 404 124
rect 540 116 548 124
rect 604 116 612 124
rect 668 116 676 124
rect 732 116 740 124
rect 796 116 804 124
rect 828 116 836 124
rect 892 116 900 124
rect 956 116 964 124
rect 988 116 996 124
rect 76 96 84 104
rect 380 96 388 104
rect 492 96 500 104
rect 556 96 564 104
rect 620 96 628 104
rect 684 96 692 104
rect 748 96 756 104
rect 812 96 820 104
rect 348 76 356 84
rect 524 76 532 84
rect 588 76 596 84
rect 652 76 660 84
rect 716 76 724 84
rect 780 76 788 84
rect 812 76 820 84
rect 908 76 916 84
rect 940 76 948 84
rect 1244 116 1252 124
rect 1372 116 1380 124
rect 1404 116 1412 124
rect 972 96 980 104
rect 1068 96 1076 104
rect 1100 96 1108 104
rect 1340 98 1348 106
rect 1468 116 1476 124
rect 1564 116 1572 124
rect 1644 116 1652 124
rect 1708 116 1716 124
rect 1820 116 1828 124
rect 1900 116 1908 124
rect 1932 116 1940 124
rect 1996 116 2004 124
rect 2044 116 2052 124
rect 2076 116 2084 124
rect 2108 116 2116 124
rect 2300 116 2308 124
rect 2364 116 2372 124
rect 2428 116 2436 124
rect 2492 116 2500 124
rect 2636 116 2644 124
rect 2716 116 2724 124
rect 2748 116 2756 124
rect 2812 116 2820 124
rect 2828 116 2836 124
rect 2892 116 2900 124
rect 2908 116 2916 124
rect 2972 116 2980 124
rect 2988 116 2996 124
rect 3052 116 3060 124
rect 3068 116 3076 124
rect 3116 116 3124 124
rect 3276 116 3284 124
rect 3372 116 3380 124
rect 3500 116 3508 124
rect 3564 116 3572 124
rect 3628 116 3636 124
rect 3660 116 3668 124
rect 3772 116 3780 124
rect 3820 116 3828 124
rect 3916 116 3924 124
rect 3980 116 3988 124
rect 4204 116 4212 124
rect 4252 116 4260 124
rect 4396 118 4404 126
rect 4492 116 4500 124
rect 4636 118 4644 126
rect 4764 116 4772 124
rect 4908 116 4916 124
rect 1468 96 1476 104
rect 1548 96 1556 104
rect 1676 96 1684 104
rect 1692 96 1700 104
rect 1804 96 1812 104
rect 1916 96 1924 104
rect 1980 96 1988 104
rect 2076 96 2084 104
rect 2092 96 2100 104
rect 2316 96 2324 104
rect 2380 96 2388 104
rect 2444 96 2452 104
rect 2508 96 2516 104
rect 2636 96 2644 104
rect 2668 96 2676 104
rect 2732 96 2740 104
rect 3116 96 3124 104
rect 3180 96 3188 104
rect 3228 96 3236 104
rect 3356 96 3364 104
rect 3452 96 3460 104
rect 3516 96 3524 104
rect 3580 96 3588 104
rect 3644 96 3652 104
rect 3932 96 3940 104
rect 3948 96 3956 104
rect 4044 96 4052 104
rect 4892 96 4900 104
rect 5052 116 5060 124
rect 5100 116 5108 124
rect 5276 118 5284 126
rect 5404 116 5412 124
rect 5532 116 5540 124
rect 5580 116 5588 124
rect 5628 116 5636 124
rect 5644 116 5652 124
rect 5708 116 5716 124
rect 5852 118 5860 126
rect 5916 116 5924 124
rect 6092 116 6100 124
rect 6172 116 6180 124
rect 6204 116 6212 124
rect 6252 116 6260 124
rect 6316 116 6324 124
rect 6396 116 6404 124
rect 6444 116 6452 124
rect 4940 96 4948 104
rect 4988 96 4996 104
rect 5036 96 5044 104
rect 6188 96 6196 104
rect 6300 96 6308 104
rect 6460 96 6468 104
rect 6476 96 6484 104
rect 972 76 980 84
rect 1724 76 1732 84
rect 1772 76 1780 84
rect 1884 76 1892 84
rect 2124 76 2132 84
rect 2140 76 2148 84
rect 2284 76 2292 84
rect 2348 76 2356 84
rect 540 56 548 64
rect 668 56 676 64
rect 796 56 804 64
rect 956 56 964 64
rect 1788 56 1796 64
rect 1900 56 1908 64
rect 2188 56 2196 64
rect 2380 76 2388 84
rect 2412 76 2420 84
rect 2476 76 2484 84
rect 2700 76 2708 84
rect 3388 76 3396 84
rect 3420 76 3428 84
rect 3484 76 3492 84
rect 3548 76 3556 84
rect 3612 76 3620 84
rect 3900 76 3908 84
rect 4268 76 4276 84
rect 4508 76 4516 84
rect 5068 76 5076 84
rect 5148 76 5156 84
rect 5516 76 5524 84
rect 5724 76 5732 84
rect 6156 76 6164 84
rect 6316 76 6324 84
rect 6332 76 6340 84
rect 6428 76 6436 84
rect 2492 56 2500 64
rect 2716 56 2724 64
rect 3244 56 3252 64
rect 3500 56 3508 64
rect 3564 56 3572 64
rect 3628 56 3636 64
rect 3916 56 3924 64
rect 604 36 612 44
rect 1820 36 1828 44
rect 2428 36 2436 44
rect 2796 36 2804 44
rect 2876 36 2884 44
rect 2956 36 2964 44
rect 3036 36 3044 44
rect 3372 36 3380 44
rect 3724 36 3732 44
rect 3980 36 3988 44
rect 4172 36 4180 44
rect 4220 36 4228 44
rect 4460 36 4468 44
rect 5132 36 5140 44
rect 5564 36 5572 44
rect 5612 36 5620 44
rect 5676 36 5684 44
rect 6236 36 6244 44
rect 6364 36 6372 44
rect 1774 6 1782 14
rect 1788 6 1796 14
rect 1802 6 1810 14
rect 4830 6 4838 14
rect 4844 6 4852 14
rect 4858 6 4866 14
<< metal2 >>
rect 2957 4857 3011 4863
rect 109 4684 115 4736
rect 13 4584 19 4676
rect 205 4664 211 4843
rect 253 4744 259 4843
rect 813 4757 915 4763
rect 381 4684 387 4736
rect 493 4684 499 4716
rect 509 4704 515 4736
rect 557 4684 563 4736
rect 621 4684 627 4756
rect 813 4744 819 4757
rect 909 4744 915 4757
rect 348 4664 356 4670
rect 13 4504 19 4536
rect 45 4524 51 4536
rect 77 4524 83 4636
rect 141 4543 147 4636
rect 173 4624 179 4636
rect 132 4537 147 4543
rect 157 4523 163 4556
rect 148 4517 163 4523
rect 77 4504 83 4516
rect 13 4364 19 4476
rect 45 4324 51 4436
rect 29 4264 35 4296
rect 61 4284 67 4496
rect 141 4304 147 4436
rect 13 4184 19 4256
rect 45 4124 51 4236
rect 13 3904 19 4036
rect 93 3904 99 4276
rect 141 4264 147 4276
rect 189 4224 195 4576
rect 205 4543 211 4656
rect 221 4564 227 4636
rect 253 4544 259 4656
rect 269 4544 275 4636
rect 317 4584 323 4664
rect 205 4537 227 4543
rect 221 4524 227 4537
rect 205 4484 211 4516
rect 253 4503 259 4536
rect 333 4524 339 4616
rect 349 4504 355 4636
rect 381 4564 387 4676
rect 429 4664 435 4676
rect 541 4664 547 4676
rect 621 4664 627 4676
rect 669 4664 675 4676
rect 685 4644 691 4696
rect 701 4644 707 4656
rect 413 4543 419 4636
rect 413 4537 428 4543
rect 445 4524 451 4556
rect 493 4544 499 4636
rect 388 4517 403 4523
rect 244 4497 259 4503
rect 356 4497 364 4503
rect 381 4484 387 4496
rect 397 4484 403 4517
rect 589 4523 595 4636
rect 621 4584 627 4636
rect 781 4584 787 4716
rect 621 4564 627 4576
rect 637 4544 643 4576
rect 813 4544 819 4716
rect 829 4704 835 4736
rect 957 4704 963 4736
rect 957 4684 963 4696
rect 909 4664 915 4676
rect 925 4644 931 4656
rect 941 4564 947 4656
rect 957 4644 963 4656
rect 973 4540 979 4656
rect 765 4524 771 4536
rect 589 4517 611 4523
rect 253 4264 259 4316
rect 301 4284 307 4456
rect 317 4304 323 4316
rect 397 4304 403 4316
rect 301 4264 307 4276
rect 349 4244 355 4276
rect 317 4184 323 4236
rect 301 4177 316 4183
rect 301 4144 307 4177
rect 333 4163 339 4196
rect 397 4164 403 4236
rect 324 4157 339 4163
rect 413 4144 419 4436
rect 429 4304 435 4316
rect 509 4304 515 4516
rect 573 4504 579 4516
rect 605 4504 611 4517
rect 797 4504 803 4536
rect 973 4524 979 4532
rect 573 4424 579 4436
rect 557 4284 563 4296
rect 589 4284 595 4496
rect 653 4304 659 4336
rect 429 4164 435 4216
rect 445 4204 451 4276
rect 461 4224 467 4276
rect 605 4264 611 4276
rect 621 4184 627 4296
rect 653 4224 659 4236
rect 125 3864 131 4136
rect 413 4123 419 4136
rect 605 4124 611 4136
rect 621 4124 627 4176
rect 653 4164 659 4216
rect 669 4184 675 4296
rect 685 4244 691 4316
rect 717 4304 723 4436
rect 717 4244 723 4276
rect 749 4264 755 4316
rect 765 4284 771 4356
rect 781 4304 787 4336
rect 733 4184 739 4236
rect 669 4144 675 4176
rect 765 4144 771 4176
rect 404 4117 419 4123
rect 141 3924 147 4076
rect 237 3963 243 4036
rect 221 3957 243 3963
rect 157 3924 163 3936
rect 189 3863 195 3876
rect 173 3857 195 3863
rect 45 3784 51 3856
rect 125 3744 131 3856
rect 125 3504 131 3736
rect 141 3726 147 3836
rect 173 3704 179 3857
rect 205 3724 211 3736
rect 221 3724 227 3957
rect 237 3904 243 3936
rect 269 3904 275 3916
rect 253 3884 259 3896
rect 365 3884 371 3894
rect 333 3864 339 3876
rect 301 3783 307 3856
rect 413 3844 419 3876
rect 301 3777 316 3783
rect 301 3744 307 3777
rect 205 3584 211 3696
rect 125 3384 131 3496
rect 221 3444 227 3456
rect 125 3344 131 3376
rect 237 3324 243 3536
rect 269 3524 275 3696
rect 333 3523 339 3816
rect 413 3744 419 3836
rect 477 3824 483 4036
rect 509 3924 515 3936
rect 509 3864 515 3916
rect 573 3884 579 3976
rect 589 3904 595 3936
rect 701 3844 707 3896
rect 349 3524 355 3696
rect 413 3564 419 3736
rect 429 3724 435 3736
rect 317 3517 339 3523
rect 317 3504 323 3517
rect 269 3484 275 3496
rect 333 3384 339 3496
rect 349 3484 355 3516
rect 429 3484 435 3496
rect 445 3484 451 3696
rect 381 3444 387 3476
rect 381 3364 387 3436
rect 413 3324 419 3356
rect 477 3344 483 3796
rect 509 3704 515 3736
rect 525 3724 531 3816
rect 557 3784 563 3836
rect 717 3824 723 4036
rect 781 3984 787 4156
rect 813 4144 819 4276
rect 829 4264 835 4276
rect 845 4143 851 4436
rect 861 4304 867 4316
rect 957 4263 963 4316
rect 989 4284 995 4843
rect 1021 4837 1043 4843
rect 1005 4644 1011 4656
rect 1021 4584 1027 4716
rect 1037 4563 1043 4837
rect 2189 4837 2211 4843
rect 1768 4806 1774 4814
rect 1782 4806 1788 4814
rect 1796 4806 1802 4814
rect 1810 4806 1816 4814
rect 1741 4783 1747 4796
rect 1741 4777 1779 4783
rect 1261 4717 1347 4723
rect 1053 4583 1059 4716
rect 1165 4704 1171 4716
rect 1181 4704 1187 4716
rect 1069 4684 1075 4696
rect 1101 4684 1107 4696
rect 1069 4664 1075 4676
rect 1101 4664 1107 4676
rect 1117 4644 1123 4676
rect 1229 4664 1235 4676
rect 1245 4623 1251 4656
rect 1261 4644 1267 4717
rect 1277 4664 1283 4696
rect 1341 4684 1347 4717
rect 1245 4617 1267 4623
rect 1053 4577 1075 4583
rect 1069 4564 1075 4577
rect 1085 4564 1091 4576
rect 1021 4557 1043 4563
rect 1021 4464 1027 4557
rect 1101 4504 1107 4596
rect 1261 4584 1267 4617
rect 1293 4603 1299 4676
rect 1309 4644 1315 4676
rect 1293 4597 1315 4603
rect 1245 4564 1251 4576
rect 1213 4524 1219 4536
rect 989 4264 995 4276
rect 1037 4264 1043 4376
rect 1181 4344 1187 4496
rect 1085 4304 1091 4316
rect 1117 4284 1123 4316
rect 1165 4304 1171 4336
rect 1069 4264 1075 4276
rect 1133 4264 1139 4296
rect 1197 4283 1203 4516
rect 1213 4324 1219 4356
rect 1229 4304 1235 4496
rect 1309 4464 1315 4597
rect 1325 4544 1331 4636
rect 1341 4564 1347 4656
rect 1389 4644 1395 4696
rect 1437 4644 1443 4656
rect 1405 4584 1411 4616
rect 1469 4584 1475 4696
rect 1485 4644 1491 4676
rect 1501 4644 1507 4716
rect 1517 4664 1523 4716
rect 1533 4644 1539 4676
rect 1373 4564 1379 4576
rect 1405 4564 1411 4576
rect 1501 4564 1507 4576
rect 1533 4563 1539 4636
rect 1549 4603 1555 4696
rect 1581 4644 1587 4736
rect 1629 4724 1635 4736
rect 1773 4704 1779 4777
rect 1837 4704 1843 4796
rect 2189 4724 2195 4837
rect 1869 4704 1875 4716
rect 1917 4704 1923 4716
rect 1981 4703 1987 4716
rect 2093 4704 2099 4716
rect 1981 4697 1996 4703
rect 2148 4697 2172 4703
rect 1597 4664 1603 4696
rect 1629 4664 1635 4696
rect 1741 4664 1747 4696
rect 1997 4684 2003 4696
rect 1837 4664 1843 4676
rect 1549 4597 1564 4603
rect 1581 4584 1587 4636
rect 1677 4584 1683 4636
rect 1725 4604 1731 4656
rect 1524 4557 1539 4563
rect 1341 4544 1347 4556
rect 1453 4544 1459 4556
rect 1469 4544 1475 4556
rect 1245 4304 1251 4336
rect 1277 4324 1283 4456
rect 1325 4443 1331 4536
rect 1453 4524 1459 4536
rect 1341 4484 1347 4516
rect 1309 4437 1331 4443
rect 1309 4324 1315 4437
rect 1325 4324 1331 4416
rect 1229 4284 1235 4296
rect 1188 4277 1203 4283
rect 1309 4264 1315 4316
rect 1453 4304 1459 4436
rect 1501 4383 1507 4516
rect 1485 4377 1507 4383
rect 948 4257 963 4263
rect 861 4204 867 4236
rect 957 4204 963 4236
rect 829 4137 851 4143
rect 765 3902 771 3916
rect 829 3904 835 4137
rect 861 4124 867 4196
rect 909 4144 915 4196
rect 1117 4184 1123 4236
rect 1101 4164 1107 4176
rect 845 3924 851 4116
rect 861 3904 867 3936
rect 621 3764 627 3796
rect 765 3764 771 3776
rect 829 3764 835 3876
rect 909 3844 915 3876
rect 893 3764 899 3836
rect 957 3784 963 3916
rect 989 3904 995 4136
rect 1005 4124 1011 4136
rect 1133 4084 1139 4236
rect 1149 4144 1155 4176
rect 1165 4164 1171 4256
rect 1213 4124 1219 4236
rect 1277 4144 1283 4156
rect 1325 4144 1331 4196
rect 1341 4144 1347 4276
rect 1357 4204 1363 4296
rect 1389 4284 1395 4296
rect 1485 4284 1491 4377
rect 1517 4264 1523 4516
rect 1421 4224 1427 4236
rect 1245 4104 1251 4136
rect 1101 3924 1107 4036
rect 1133 3924 1139 3956
rect 1005 3804 1011 3836
rect 653 3744 659 3756
rect 509 3484 515 3556
rect 525 3544 531 3636
rect 525 3504 531 3516
rect 605 3504 611 3736
rect 733 3724 739 3736
rect 653 3524 659 3676
rect 685 3584 691 3696
rect 749 3584 755 3736
rect 957 3724 963 3756
rect 1005 3744 1011 3796
rect 1053 3744 1059 3916
rect 957 3704 963 3716
rect 733 3557 748 3563
rect 541 3364 547 3396
rect 605 3324 611 3496
rect 653 3484 659 3516
rect 685 3484 691 3496
rect 621 3344 627 3476
rect 653 3384 659 3416
rect 637 3324 643 3336
rect 125 3104 131 3236
rect 637 3124 643 3316
rect 669 3304 675 3436
rect 733 3324 739 3557
rect 749 3504 755 3556
rect 765 3484 771 3636
rect 957 3623 963 3696
rect 957 3617 979 3623
rect 765 3364 771 3476
rect 749 3344 755 3356
rect 781 3344 787 3536
rect 813 3464 819 3516
rect 813 3444 819 3456
rect 845 3404 851 3476
rect 941 3464 947 3496
rect 653 3104 659 3296
rect 669 3144 675 3156
rect 765 3144 771 3316
rect 781 3284 787 3336
rect 845 3324 851 3376
rect 877 3324 883 3436
rect 893 3424 899 3456
rect 909 3403 915 3436
rect 893 3397 915 3403
rect 893 3324 899 3397
rect 909 3364 915 3376
rect 925 3344 931 3396
rect 941 3384 947 3416
rect 957 3344 963 3356
rect 973 3344 979 3617
rect 1005 3484 1011 3736
rect 1085 3704 1091 3756
rect 1021 3584 1027 3636
rect 1021 3504 1027 3516
rect 1037 3504 1043 3696
rect 1053 3524 1059 3576
rect 1117 3544 1123 3876
rect 1149 3864 1155 3916
rect 1181 3904 1187 3976
rect 1197 3924 1203 3936
rect 1213 3824 1219 3836
rect 1245 3804 1251 4096
rect 1277 3964 1283 4076
rect 1261 3843 1267 3856
rect 1261 3837 1276 3843
rect 1149 3744 1155 3776
rect 1165 3744 1171 3756
rect 1309 3724 1315 4056
rect 1325 3984 1331 4136
rect 1357 4084 1363 4156
rect 1485 4124 1491 4136
rect 1325 3744 1331 3796
rect 1341 3744 1347 3896
rect 1357 3764 1363 4076
rect 1405 3864 1411 3894
rect 1437 3884 1443 4116
rect 1469 3924 1475 3936
rect 1389 3737 1404 3743
rect 1325 3724 1331 3736
rect 1389 3724 1395 3737
rect 1421 3724 1427 3776
rect 1133 3504 1139 3636
rect 1021 3384 1027 3496
rect 1069 3484 1075 3496
rect 1197 3404 1203 3476
rect 1213 3404 1219 3436
rect 1069 3344 1075 3376
rect 1245 3364 1251 3436
rect 1277 3424 1283 3696
rect 1437 3684 1443 3876
rect 1469 3744 1475 3916
rect 1501 3883 1507 4236
rect 1533 3904 1539 4536
rect 1549 4524 1555 4576
rect 1565 4524 1571 4556
rect 1677 4544 1683 4576
rect 1629 4524 1635 4536
rect 1661 4524 1667 4536
rect 1757 4524 1763 4636
rect 1773 4564 1779 4656
rect 1885 4644 1891 4656
rect 2061 4644 2067 4696
rect 2157 4644 2163 4676
rect 2173 4664 2179 4676
rect 2109 4584 2115 4636
rect 1885 4524 1891 4556
rect 1901 4544 1907 4556
rect 2061 4544 2067 4576
rect 2157 4564 2163 4576
rect 2205 4564 2211 4716
rect 2221 4664 2227 4776
rect 2237 4724 2243 4843
rect 2333 4684 2339 4776
rect 2365 4724 2371 4776
rect 2365 4704 2371 4716
rect 2285 4664 2291 4676
rect 2365 4664 2371 4696
rect 2237 4544 2243 4636
rect 2301 4564 2307 4636
rect 1677 4504 1683 4516
rect 1565 4484 1571 4496
rect 1693 4484 1699 4496
rect 1768 4406 1774 4414
rect 1782 4406 1788 4414
rect 1796 4406 1802 4414
rect 1810 4406 1816 4414
rect 1597 4284 1603 4316
rect 1661 4304 1667 4316
rect 1549 4244 1555 4276
rect 1549 4183 1555 4236
rect 1549 4177 1571 4183
rect 1565 4104 1571 4177
rect 1613 4144 1619 4156
rect 1549 3904 1555 3916
rect 1565 3884 1571 4096
rect 1581 3904 1587 4116
rect 1629 4064 1635 4236
rect 1661 4124 1667 4156
rect 1677 4124 1683 4136
rect 1725 4104 1731 4376
rect 1741 4304 1747 4376
rect 1853 4304 1859 4376
rect 1885 4317 1900 4323
rect 1757 4144 1763 4276
rect 1853 4124 1859 4296
rect 1869 4224 1875 4236
rect 1885 4184 1891 4317
rect 1917 4284 1923 4436
rect 1933 4304 1939 4516
rect 1949 4284 1955 4536
rect 2045 4524 2051 4536
rect 2301 4524 2307 4556
rect 2349 4544 2355 4636
rect 2365 4524 2371 4556
rect 2381 4544 2387 4676
rect 2413 4564 2419 4576
rect 1997 4304 2003 4496
rect 2045 4364 2051 4436
rect 2029 4304 2035 4316
rect 2077 4304 2083 4316
rect 1885 4164 1891 4176
rect 1901 4144 1907 4156
rect 1917 4144 1923 4276
rect 1997 4264 2003 4296
rect 2093 4284 2099 4296
rect 1965 4244 1971 4256
rect 2029 4244 2035 4256
rect 2077 4164 2083 4256
rect 2013 4144 2019 4156
rect 2077 4144 2083 4156
rect 1821 4044 1827 4096
rect 1613 3944 1619 4036
rect 1597 3884 1603 3916
rect 1613 3884 1619 3936
rect 1629 3924 1635 4036
rect 1693 3904 1699 4036
rect 1768 4006 1774 4014
rect 1782 4006 1788 4014
rect 1796 4006 1802 4014
rect 1810 4006 1816 4014
rect 1501 3877 1516 3883
rect 1485 3784 1491 3876
rect 1501 3724 1507 3877
rect 1629 3864 1635 3896
rect 1837 3884 1843 4116
rect 1917 4104 1923 4136
rect 2109 4124 2115 4276
rect 2141 4264 2147 4516
rect 2269 4504 2275 4516
rect 2333 4484 2339 4496
rect 2269 4383 2275 4436
rect 2269 4377 2291 4383
rect 2189 4304 2195 4336
rect 2205 4244 2211 4276
rect 2125 4204 2131 4236
rect 2205 4164 2211 4236
rect 2237 4224 2243 4296
rect 2269 4284 2275 4356
rect 2157 4144 2163 4156
rect 2077 4104 2083 4116
rect 2221 4104 2227 4136
rect 2253 4103 2259 4196
rect 2285 4144 2291 4377
rect 2333 4324 2339 4356
rect 2301 4224 2307 4296
rect 2349 4284 2355 4516
rect 2397 4324 2403 4516
rect 2413 4504 2419 4556
rect 2477 4524 2483 4696
rect 2493 4564 2499 4676
rect 2509 4664 2515 4796
rect 2653 4743 2659 4843
rect 2957 4837 2963 4857
rect 2973 4837 2995 4843
rect 2973 4823 2979 4837
rect 3005 4823 3011 4857
rect 2909 4817 2979 4823
rect 2989 4817 3011 4823
rect 2541 4737 2579 4743
rect 2653 4737 2675 4743
rect 2541 4724 2547 4737
rect 2573 4723 2579 4737
rect 2573 4717 2588 4723
rect 2605 4683 2611 4716
rect 2596 4677 2611 4683
rect 2589 4664 2595 4676
rect 2557 4584 2563 4636
rect 2525 4544 2531 4556
rect 2621 4544 2627 4636
rect 2669 4564 2675 4737
rect 2685 4684 2691 4716
rect 2733 4664 2739 4796
rect 2909 4783 2915 4817
rect 2989 4803 2995 4817
rect 2893 4777 2915 4783
rect 2957 4797 2995 4803
rect 2861 4684 2867 4696
rect 2749 4584 2755 4676
rect 2861 4624 2867 4656
rect 2813 4584 2819 4616
rect 2445 4284 2451 4516
rect 2493 4464 2499 4536
rect 2685 4524 2691 4556
rect 2701 4524 2707 4536
rect 2557 4504 2563 4516
rect 2653 4504 2659 4516
rect 2461 4324 2467 4336
rect 2541 4304 2547 4316
rect 2493 4284 2499 4296
rect 2333 4164 2339 4236
rect 2301 4124 2307 4136
rect 2253 4097 2268 4103
rect 2333 4064 2339 4116
rect 2349 4084 2355 4136
rect 1949 3904 1955 4036
rect 1565 3724 1571 3836
rect 1677 3784 1683 3856
rect 1693 3764 1699 3776
rect 1453 3704 1459 3716
rect 1597 3684 1603 3716
rect 1309 3503 1315 3636
rect 1309 3497 1324 3503
rect 1405 3484 1411 3676
rect 1453 3624 1459 3636
rect 1485 3502 1491 3616
rect 1613 3484 1619 3536
rect 1629 3524 1635 3696
rect 1677 3524 1683 3636
rect 1709 3484 1715 3756
rect 1741 3744 1747 3776
rect 1837 3684 1843 3696
rect 1853 3684 1859 3896
rect 1933 3804 1939 3876
rect 1997 3844 2003 3916
rect 2029 3884 2035 3936
rect 2045 3824 2051 3856
rect 2061 3744 2067 4056
rect 2093 3984 2099 4016
rect 2109 3904 2115 4036
rect 2109 3884 2115 3896
rect 1741 3523 1747 3676
rect 1768 3606 1774 3614
rect 1782 3606 1788 3614
rect 1796 3606 1802 3614
rect 1810 3606 1816 3614
rect 1741 3517 1756 3523
rect 1517 3464 1523 3476
rect 877 3303 883 3316
rect 973 3304 979 3336
rect 868 3297 883 3303
rect 813 3164 819 3236
rect 925 3184 931 3196
rect 1101 3124 1107 3336
rect 1133 3326 1139 3336
rect 1197 3324 1203 3336
rect 1213 3184 1219 3216
rect 1028 3117 1052 3123
rect 861 3104 867 3116
rect 45 2824 51 2916
rect 61 2904 67 2956
rect 77 2784 83 3096
rect 125 3084 131 3096
rect 205 3043 211 3076
rect 205 3037 227 3043
rect 93 2884 99 3016
rect 221 2984 227 3037
rect 301 3024 307 3076
rect 509 3004 515 3096
rect 701 3064 707 3096
rect 628 3057 643 3063
rect 589 3024 595 3056
rect 541 2984 547 2996
rect 621 2984 627 3016
rect 637 2964 643 3057
rect 941 3063 947 3076
rect 973 3064 979 3116
rect 925 3057 947 3063
rect 685 3004 691 3036
rect 797 2984 803 3056
rect 109 2924 115 2936
rect 93 2744 99 2876
rect 125 2844 131 2896
rect 189 2844 195 2876
rect 237 2844 243 2896
rect 109 2723 115 2836
rect 109 2717 124 2723
rect 173 2704 179 2736
rect 221 2704 227 2836
rect 269 2804 275 2916
rect 317 2904 323 2936
rect 381 2924 387 2956
rect 525 2944 531 2956
rect 301 2704 307 2796
rect 189 2684 195 2696
rect 13 2643 19 2676
rect 173 2664 179 2676
rect 13 2637 35 2643
rect 29 2584 35 2637
rect 77 2564 83 2636
rect 77 2504 83 2556
rect 109 2504 115 2516
rect 45 2464 51 2496
rect 125 2484 131 2536
rect 141 2484 147 2636
rect 205 2544 211 2636
rect 221 2564 227 2676
rect 285 2564 291 2676
rect 269 2544 275 2556
rect 301 2544 307 2696
rect 317 2684 323 2876
rect 317 2623 323 2676
rect 349 2664 355 2876
rect 413 2844 419 2936
rect 605 2924 611 2936
rect 397 2704 403 2716
rect 429 2684 435 2916
rect 445 2884 451 2896
rect 477 2704 483 2916
rect 525 2884 531 2916
rect 541 2904 547 2916
rect 493 2784 499 2796
rect 525 2724 531 2876
rect 541 2804 547 2896
rect 685 2884 691 2916
rect 701 2904 707 2936
rect 749 2924 755 2936
rect 781 2904 787 2956
rect 829 2884 835 2916
rect 845 2904 851 2956
rect 909 2924 915 2956
rect 669 2844 675 2876
rect 637 2784 643 2836
rect 589 2704 595 2736
rect 701 2724 707 2816
rect 717 2784 723 2876
rect 925 2844 931 3057
rect 973 2943 979 3036
rect 989 2984 995 3116
rect 973 2937 988 2943
rect 973 2924 979 2937
rect 909 2784 915 2836
rect 525 2684 531 2696
rect 429 2664 435 2676
rect 317 2617 339 2623
rect 285 2524 291 2536
rect 205 2504 211 2516
rect 237 2504 243 2516
rect 45 2284 51 2296
rect 13 1944 19 2236
rect 61 2164 67 2436
rect 125 2284 131 2336
rect 109 2204 115 2236
rect 61 2104 67 2156
rect 93 2124 99 2136
rect 141 2124 147 2456
rect 189 2364 195 2436
rect 173 2324 179 2356
rect 157 2264 163 2316
rect 189 2164 195 2176
rect 77 2104 83 2116
rect 29 2084 35 2096
rect 29 1984 35 2076
rect 45 2064 51 2076
rect 93 2004 99 2116
rect 109 1984 115 2096
rect 141 2084 147 2116
rect 157 1984 163 1996
rect 13 1924 19 1936
rect 45 1924 51 1936
rect 93 1924 99 1936
rect 125 1924 131 1956
rect 173 1924 179 1936
rect 13 1764 19 1916
rect 29 1743 35 1896
rect 45 1744 51 1756
rect 20 1737 35 1743
rect 13 1584 19 1736
rect 45 1684 51 1696
rect 93 1684 99 1916
rect 189 1903 195 2116
rect 205 2104 211 2496
rect 301 2464 307 2536
rect 333 2504 339 2617
rect 365 2524 371 2556
rect 429 2544 435 2656
rect 573 2604 579 2676
rect 589 2584 595 2696
rect 621 2584 627 2676
rect 637 2604 643 2696
rect 685 2664 691 2696
rect 717 2684 723 2696
rect 733 2684 739 2736
rect 765 2684 771 2696
rect 717 2644 723 2676
rect 733 2623 739 2676
rect 781 2644 787 2676
rect 877 2624 883 2716
rect 893 2684 899 2736
rect 925 2724 931 2796
rect 941 2784 947 2896
rect 973 2704 979 2776
rect 1053 2764 1059 3096
rect 1149 3084 1155 3096
rect 1245 3084 1251 3356
rect 1309 3304 1315 3356
rect 1373 3344 1379 3416
rect 1261 3104 1267 3236
rect 1373 3224 1379 3316
rect 1389 3284 1395 3336
rect 1405 3324 1411 3396
rect 1469 3344 1475 3376
rect 1501 3324 1507 3356
rect 1517 3344 1523 3456
rect 1629 3424 1635 3436
rect 1437 3304 1443 3316
rect 1453 3304 1459 3316
rect 1373 3164 1379 3216
rect 1389 3184 1395 3216
rect 1405 3184 1411 3236
rect 1485 3124 1491 3256
rect 1069 3044 1075 3056
rect 1069 2963 1075 3036
rect 1085 3024 1091 3076
rect 1133 3064 1139 3076
rect 1261 3064 1267 3096
rect 1325 3084 1331 3116
rect 1437 3104 1443 3116
rect 1357 3084 1363 3096
rect 1485 3084 1491 3116
rect 1501 3104 1507 3296
rect 1533 3284 1539 3376
rect 1645 3364 1651 3416
rect 1549 3304 1555 3316
rect 1565 3304 1571 3356
rect 1613 3324 1619 3336
rect 1677 3264 1683 3436
rect 1517 3117 1532 3123
rect 1517 3084 1523 3117
rect 1549 3084 1555 3156
rect 1405 3064 1411 3076
rect 1069 2957 1084 2963
rect 1069 2844 1075 2936
rect 1085 2923 1091 2956
rect 1117 2924 1123 3036
rect 1085 2917 1100 2923
rect 1117 2824 1123 2836
rect 1117 2784 1123 2796
rect 1037 2724 1043 2756
rect 1117 2704 1123 2756
rect 1133 2704 1139 3056
rect 1165 2984 1171 3016
rect 1261 2964 1267 3056
rect 1213 2904 1219 2936
rect 1341 2924 1347 2976
rect 1213 2784 1219 2896
rect 717 2617 739 2623
rect 669 2584 675 2596
rect 717 2584 723 2617
rect 893 2584 899 2676
rect 989 2664 995 2676
rect 1005 2624 1011 2656
rect 445 2544 451 2556
rect 525 2524 531 2536
rect 333 2464 339 2496
rect 253 2384 259 2456
rect 301 2384 307 2436
rect 365 2384 371 2456
rect 397 2363 403 2516
rect 429 2484 435 2516
rect 493 2504 499 2516
rect 525 2504 531 2516
rect 653 2503 659 2536
rect 685 2504 691 2536
rect 653 2497 675 2503
rect 589 2484 595 2496
rect 397 2357 412 2363
rect 269 2104 275 2356
rect 324 2337 348 2343
rect 388 2337 403 2343
rect 301 2284 307 2296
rect 349 2264 355 2316
rect 397 2303 403 2337
rect 413 2324 419 2356
rect 461 2303 467 2336
rect 525 2324 531 2436
rect 605 2324 611 2356
rect 397 2297 467 2303
rect 365 2284 371 2296
rect 461 2244 467 2276
rect 413 2184 419 2236
rect 397 2104 403 2136
rect 269 1984 275 2076
rect 349 1984 355 2076
rect 205 1924 211 1936
rect 237 1924 243 1936
rect 173 1897 195 1903
rect 29 1464 35 1536
rect 77 1464 83 1516
rect 109 1384 115 1736
rect 125 1724 131 1736
rect 157 1683 163 1896
rect 173 1784 179 1897
rect 173 1704 179 1716
rect 221 1704 227 1716
rect 141 1677 163 1683
rect 141 1584 147 1677
rect 189 1584 195 1676
rect 205 1544 211 1556
rect 125 1464 131 1536
rect 157 1524 163 1536
rect 221 1523 227 1636
rect 237 1584 243 1916
rect 253 1823 259 1836
rect 269 1823 275 1856
rect 253 1817 275 1823
rect 253 1784 259 1796
rect 269 1724 275 1817
rect 253 1644 259 1696
rect 269 1684 275 1696
rect 285 1644 291 1936
rect 429 1904 435 2136
rect 477 2124 483 2136
rect 445 2004 451 2116
rect 461 2104 467 2116
rect 301 1703 307 1756
rect 349 1744 355 1796
rect 365 1784 371 1876
rect 461 1863 467 1916
rect 452 1857 467 1863
rect 301 1697 316 1703
rect 445 1684 451 1696
rect 253 1544 259 1556
rect 205 1517 227 1523
rect 157 1384 163 1476
rect 205 1384 211 1517
rect 253 1384 259 1536
rect 301 1504 307 1536
rect 333 1524 339 1636
rect 276 1497 291 1503
rect 61 1304 67 1356
rect 157 1337 172 1343
rect 93 1324 99 1336
rect 29 1144 35 1276
rect 45 1184 51 1296
rect 77 1284 83 1316
rect 77 1124 83 1176
rect 29 1063 35 1116
rect 61 1103 67 1116
rect 61 1097 76 1103
rect 45 1084 51 1096
rect 29 1057 51 1063
rect 13 924 19 1036
rect 45 984 51 1057
rect 61 964 67 1097
rect 93 1084 99 1316
rect 141 1304 147 1336
rect 157 1184 163 1337
rect 205 1124 211 1356
rect 221 1184 227 1336
rect 237 1304 243 1336
rect 237 1164 243 1296
rect 141 1104 147 1116
rect 109 1063 115 1096
rect 93 1057 115 1063
rect 93 984 99 1057
rect 77 964 83 976
rect 29 944 35 956
rect 109 944 115 996
rect 173 984 179 1056
rect 221 1023 227 1096
rect 237 1044 243 1136
rect 253 1084 259 1316
rect 285 1264 291 1497
rect 317 1464 323 1476
rect 381 1464 387 1676
rect 445 1484 451 1536
rect 461 1463 467 1716
rect 477 1684 483 2116
rect 493 2084 499 2296
rect 573 2244 579 2296
rect 509 2184 515 2236
rect 589 2204 595 2276
rect 637 2244 643 2296
rect 653 2204 659 2276
rect 669 2264 675 2497
rect 701 2483 707 2496
rect 692 2477 707 2483
rect 685 2384 691 2476
rect 797 2444 803 2556
rect 813 2544 819 2576
rect 861 2544 867 2556
rect 845 2524 851 2536
rect 845 2444 851 2496
rect 957 2444 963 2536
rect 973 2524 979 2536
rect 989 2524 995 2536
rect 1037 2524 1043 2556
rect 1053 2524 1059 2636
rect 1101 2563 1107 2656
rect 1117 2584 1123 2676
rect 1197 2664 1203 2676
rect 1165 2584 1171 2656
rect 1213 2644 1219 2696
rect 1229 2684 1235 2896
rect 1293 2724 1299 2736
rect 1277 2624 1283 2676
rect 1293 2623 1299 2716
rect 1284 2617 1299 2623
rect 1309 2697 1324 2703
rect 1165 2564 1171 2576
rect 1181 2564 1187 2616
rect 1213 2584 1219 2616
rect 1309 2584 1315 2697
rect 1325 2684 1331 2696
rect 1341 2684 1347 2916
rect 1389 2884 1395 3036
rect 1421 2924 1427 3036
rect 1517 2984 1523 3076
rect 1549 2944 1555 2956
rect 1357 2784 1363 2876
rect 1501 2864 1507 2936
rect 1517 2904 1523 2916
rect 1357 2704 1363 2776
rect 1389 2704 1395 2836
rect 1453 2784 1459 2836
rect 1565 2744 1571 3176
rect 1581 3124 1587 3236
rect 1613 3104 1619 3156
rect 1629 3144 1635 3236
rect 1629 3104 1635 3136
rect 1677 3104 1683 3136
rect 1581 2944 1587 3036
rect 1693 2944 1699 3456
rect 1709 3344 1715 3436
rect 1725 3340 1731 3456
rect 1821 3444 1827 3496
rect 1869 3484 1875 3696
rect 1997 3684 2003 3736
rect 2029 3704 2035 3736
rect 2077 3704 2083 3756
rect 2125 3724 2131 3736
rect 1837 3464 1843 3476
rect 1741 3364 1747 3436
rect 1853 3384 1859 3436
rect 1869 3404 1875 3456
rect 1869 3344 1875 3376
rect 1725 3304 1731 3332
rect 1773 3324 1779 3336
rect 1768 3206 1774 3214
rect 1782 3206 1788 3214
rect 1796 3206 1802 3214
rect 1810 3206 1816 3214
rect 1757 3104 1763 3116
rect 1725 3084 1731 3096
rect 1741 3084 1747 3096
rect 1837 3084 1843 3136
rect 1613 2884 1619 2896
rect 1677 2844 1683 2918
rect 1693 2884 1699 2936
rect 1325 2564 1331 2636
rect 1341 2564 1347 2676
rect 1389 2663 1395 2676
rect 1373 2657 1395 2663
rect 1373 2584 1379 2657
rect 1501 2644 1507 2656
rect 1437 2584 1443 2636
rect 1092 2557 1107 2563
rect 829 2317 844 2323
rect 669 2244 675 2256
rect 525 1924 531 1996
rect 541 1904 547 2036
rect 557 1904 563 2116
rect 589 2103 595 2156
rect 589 2097 604 2103
rect 493 1884 499 1896
rect 493 1724 499 1876
rect 509 1864 515 1876
rect 509 1764 515 1856
rect 525 1743 531 1836
rect 516 1737 531 1743
rect 509 1544 515 1656
rect 525 1584 531 1716
rect 541 1684 547 1736
rect 509 1524 515 1536
rect 557 1523 563 1736
rect 573 1704 579 2096
rect 685 2084 691 2136
rect 717 2084 723 2156
rect 781 2103 787 2236
rect 813 2224 819 2276
rect 829 2264 835 2317
rect 973 2304 979 2316
rect 829 2244 835 2256
rect 845 2183 851 2236
rect 861 2184 867 2236
rect 877 2224 883 2276
rect 941 2264 947 2276
rect 829 2177 851 2183
rect 829 2144 835 2177
rect 957 2164 963 2236
rect 829 2124 835 2136
rect 781 2097 796 2103
rect 781 2083 787 2097
rect 772 2077 787 2083
rect 589 1984 595 2076
rect 669 2004 675 2036
rect 589 1884 595 1896
rect 669 1884 675 1896
rect 701 1884 707 1916
rect 717 1904 723 1996
rect 781 1924 787 2036
rect 829 1924 835 2116
rect 548 1517 563 1523
rect 525 1504 531 1516
rect 589 1504 595 1836
rect 621 1724 627 1876
rect 669 1784 675 1876
rect 765 1764 771 1876
rect 797 1844 803 1916
rect 845 1864 851 2156
rect 925 1984 931 2116
rect 957 1964 963 2156
rect 973 2104 979 2276
rect 989 2164 995 2516
rect 1005 2184 1011 2216
rect 1021 2204 1027 2316
rect 1069 2304 1075 2316
rect 1069 2224 1075 2276
rect 1021 2024 1027 2156
rect 1069 2124 1075 2196
rect 1085 2124 1091 2516
rect 1101 2304 1107 2557
rect 1117 2324 1123 2536
rect 1149 2384 1155 2516
rect 1117 2304 1123 2316
rect 1181 2304 1187 2556
rect 1197 2504 1203 2556
rect 1325 2544 1331 2556
rect 1341 2544 1347 2556
rect 1197 2317 1212 2323
rect 1133 2224 1139 2276
rect 1149 2163 1155 2236
rect 1140 2157 1155 2163
rect 877 1904 883 1956
rect 1021 1924 1027 2016
rect 1117 1924 1123 2036
rect 861 1884 867 1896
rect 877 1884 883 1896
rect 909 1884 915 1896
rect 1005 1884 1011 1916
rect 781 1784 787 1836
rect 813 1804 819 1836
rect 637 1704 643 1736
rect 781 1724 787 1756
rect 829 1724 835 1836
rect 701 1704 707 1716
rect 717 1704 723 1716
rect 845 1704 851 1756
rect 861 1704 867 1876
rect 941 1864 947 1876
rect 909 1744 915 1796
rect 925 1744 931 1836
rect 941 1784 947 1856
rect 973 1744 979 1876
rect 1005 1764 1011 1796
rect 1021 1764 1027 1836
rect 1069 1744 1075 1916
rect 1133 1884 1139 2156
rect 1181 2144 1187 2296
rect 1165 2064 1171 2116
rect 1181 2104 1187 2136
rect 1197 2124 1203 2317
rect 1229 2283 1235 2516
rect 1373 2504 1379 2536
rect 1261 2324 1267 2436
rect 1220 2277 1235 2283
rect 1213 2104 1219 2276
rect 1325 2264 1331 2276
rect 1373 2264 1379 2496
rect 1245 2144 1251 2216
rect 1268 2117 1283 2123
rect 1149 2024 1155 2036
rect 1165 1904 1171 2056
rect 1181 1964 1187 2096
rect 1181 1884 1187 1936
rect 1197 1904 1203 1916
rect 1229 1884 1235 2096
rect 1261 1984 1267 2096
rect 1277 2064 1283 2117
rect 1309 2123 1315 2136
rect 1300 2117 1315 2123
rect 1309 2104 1315 2117
rect 1341 2123 1347 2256
rect 1389 2184 1395 2436
rect 1421 2317 1436 2323
rect 1421 2184 1427 2317
rect 1469 2264 1475 2356
rect 1501 2324 1507 2636
rect 1517 2384 1523 2516
rect 1533 2284 1539 2636
rect 1565 2564 1571 2696
rect 1629 2584 1635 2596
rect 1661 2323 1667 2776
rect 1693 2684 1699 2876
rect 1709 2764 1715 3036
rect 1805 2884 1811 2916
rect 1837 2864 1843 3076
rect 1768 2806 1774 2814
rect 1782 2806 1788 2814
rect 1796 2806 1802 2814
rect 1810 2806 1816 2814
rect 1853 2723 1859 3016
rect 1869 2924 1875 2936
rect 1844 2717 1859 2723
rect 1700 2677 1715 2683
rect 1652 2317 1667 2323
rect 1581 2284 1587 2296
rect 1332 2117 1347 2123
rect 1437 2104 1443 2236
rect 1469 2204 1475 2256
rect 1517 2203 1523 2236
rect 1501 2197 1523 2203
rect 1277 1984 1283 2056
rect 1325 1923 1331 2036
rect 1316 1917 1331 1923
rect 1245 1864 1251 1876
rect 1293 1864 1299 1916
rect 1341 1884 1347 2076
rect 1357 1864 1363 2096
rect 1421 2084 1427 2096
rect 1389 1924 1395 1936
rect 1405 1904 1411 1916
rect 1421 1884 1427 2076
rect 1501 1884 1507 2197
rect 1533 1924 1539 2196
rect 1549 2184 1555 2256
rect 1597 2126 1603 2316
rect 1677 2284 1683 2296
rect 1645 2183 1651 2256
rect 1645 2177 1660 2183
rect 1629 2124 1635 2136
rect 1453 1864 1459 1876
rect 1517 1864 1523 1896
rect 1581 1884 1587 1996
rect 1629 1924 1635 1936
rect 1661 1904 1667 2036
rect 1693 1964 1699 2556
rect 1709 2524 1715 2677
rect 1757 2526 1763 2616
rect 1789 2604 1795 2656
rect 1869 2584 1875 2596
rect 1768 2406 1774 2414
rect 1782 2406 1788 2414
rect 1796 2406 1802 2414
rect 1810 2406 1816 2414
rect 1725 2324 1731 2376
rect 1677 1904 1683 1956
rect 1693 1884 1699 1936
rect 1725 1884 1731 1916
rect 1741 1904 1747 2136
rect 1773 2124 1779 2236
rect 1821 2144 1827 2336
rect 1853 2304 1859 2536
rect 1885 2364 1891 3576
rect 2045 3543 2051 3636
rect 2029 3537 2051 3543
rect 2029 3524 2035 3537
rect 1981 3484 1987 3516
rect 2077 3484 2083 3696
rect 2125 3544 2131 3636
rect 2093 3524 2099 3536
rect 2141 3504 2147 3676
rect 2157 3664 2163 3836
rect 2173 3744 2179 3816
rect 2189 3764 2195 3836
rect 2157 3524 2163 3536
rect 2189 3524 2195 3756
rect 2221 3524 2227 3836
rect 1917 3424 1923 3436
rect 1917 3344 1923 3396
rect 1933 3364 1939 3376
rect 1949 3304 1955 3416
rect 1997 3384 2003 3476
rect 2141 3464 2147 3496
rect 2157 3484 2163 3516
rect 2221 3504 2227 3516
rect 2189 3484 2195 3496
rect 2285 3484 2291 3776
rect 2301 3724 2307 4036
rect 2317 3902 2323 3916
rect 2381 3904 2387 4076
rect 2397 3943 2403 4236
rect 2429 4164 2435 4236
rect 2445 4164 2451 4276
rect 2525 4264 2531 4296
rect 2573 4264 2579 4416
rect 2589 4324 2595 4436
rect 2589 4304 2595 4316
rect 2413 4104 2419 4136
rect 2429 4124 2435 4156
rect 2413 4084 2419 4096
rect 2461 4083 2467 4236
rect 2509 4104 2515 4156
rect 2452 4077 2467 4083
rect 2397 3937 2419 3943
rect 2381 3884 2387 3896
rect 2317 3744 2323 3856
rect 2397 3824 2403 3896
rect 2397 3704 2403 3736
rect 2413 3724 2419 3937
rect 2429 3924 2435 4036
rect 2445 3984 2451 4056
rect 2541 3904 2547 4256
rect 2461 3844 2467 3856
rect 2445 3524 2451 3836
rect 2461 3744 2467 3776
rect 2477 3764 2483 3896
rect 2557 3883 2563 4036
rect 2548 3877 2563 3883
rect 2493 3824 2499 3876
rect 2509 3744 2515 3836
rect 2573 3764 2579 4256
rect 2637 4244 2643 4316
rect 2653 4304 2659 4496
rect 2685 4264 2691 4276
rect 2701 4263 2707 4516
rect 2692 4257 2707 4263
rect 2621 4124 2627 4176
rect 2653 4164 2659 4256
rect 2733 4244 2739 4296
rect 2749 4224 2755 4496
rect 2765 4444 2771 4556
rect 2621 3904 2627 4116
rect 2637 4084 2643 4136
rect 2717 4124 2723 4136
rect 2749 4124 2755 4156
rect 2765 4144 2771 4236
rect 2781 4144 2787 4276
rect 2797 4264 2803 4356
rect 2797 4184 2803 4216
rect 2653 4064 2659 4116
rect 2717 4084 2723 4096
rect 2669 3904 2675 4036
rect 2813 3904 2819 4556
rect 2861 4344 2867 4436
rect 2877 4364 2883 4636
rect 2893 4564 2899 4777
rect 2925 4697 2940 4703
rect 2909 4664 2915 4696
rect 2925 4664 2931 4697
rect 2957 4683 2963 4797
rect 3021 4704 3027 4843
rect 3053 4837 3075 4843
rect 2973 4697 3011 4703
rect 2973 4684 2979 4697
rect 2941 4677 2963 4683
rect 2909 4564 2915 4656
rect 2909 4524 2915 4536
rect 2893 4444 2899 4496
rect 2925 4344 2931 4636
rect 2941 4564 2947 4677
rect 3005 4683 3011 4697
rect 3037 4683 3043 4696
rect 3053 4684 3059 4716
rect 3005 4677 3043 4683
rect 2957 4584 2963 4656
rect 2989 4624 2995 4676
rect 2941 4444 2947 4496
rect 2877 4324 2883 4336
rect 2829 4184 2835 4316
rect 2861 4304 2867 4316
rect 2845 4224 2851 4296
rect 2893 4224 2899 4316
rect 2941 4284 2947 4436
rect 2957 4384 2963 4516
rect 3053 4424 3059 4676
rect 3069 4644 3075 4837
rect 3085 4744 3091 4843
rect 3117 4764 3123 4843
rect 3149 4764 3155 4843
rect 3117 4684 3123 4696
rect 3149 4684 3155 4736
rect 3181 4684 3187 4843
rect 3213 4784 3219 4843
rect 3245 4804 3251 4843
rect 4824 4806 4830 4814
rect 4838 4806 4844 4814
rect 4852 4806 4858 4814
rect 4866 4806 4872 4814
rect 4989 4724 4995 4736
rect 4996 4717 5011 4723
rect 3245 4544 3251 4676
rect 3304 4606 3310 4614
rect 3318 4606 3324 4614
rect 3332 4606 3338 4614
rect 3346 4606 3352 4614
rect 3405 4564 3411 4636
rect 3277 4544 3283 4556
rect 3101 4524 3107 4536
rect 3165 4444 3171 4496
rect 2829 4144 2835 4176
rect 2861 4164 2867 4176
rect 2909 4164 2915 4236
rect 2909 4124 2915 4136
rect 2925 4124 2931 4136
rect 2941 4124 2947 4156
rect 2989 4144 2995 4276
rect 2829 4104 2835 4116
rect 2893 3903 2899 4036
rect 2877 3897 2899 3903
rect 2509 3644 2515 3716
rect 2557 3584 2563 3736
rect 2637 3724 2643 3856
rect 2717 3764 2723 3876
rect 2765 3804 2771 3836
rect 2653 3744 2659 3756
rect 2765 3724 2771 3796
rect 2580 3697 2588 3703
rect 2532 3517 2547 3523
rect 2221 3464 2227 3476
rect 2013 3404 2019 3436
rect 1901 2964 1907 3236
rect 1917 2984 1923 3276
rect 2013 3184 2019 3296
rect 2061 3084 2067 3336
rect 2093 3064 2099 3436
rect 2237 3424 2243 3436
rect 2125 3344 2131 3356
rect 2157 3324 2163 3336
rect 2205 3324 2211 3376
rect 2221 3304 2227 3336
rect 2221 3264 2227 3296
rect 2253 3104 2259 3336
rect 2317 3104 2323 3396
rect 2333 3244 2339 3436
rect 2349 3344 2355 3476
rect 2429 3284 2435 3356
rect 2525 3344 2531 3436
rect 2541 3384 2547 3517
rect 2557 3504 2563 3516
rect 2573 3484 2579 3696
rect 2637 3584 2643 3636
rect 2701 3504 2707 3576
rect 2813 3524 2819 3696
rect 2829 3504 2835 3896
rect 2877 3784 2883 3897
rect 2989 3884 2995 4136
rect 3005 4024 3011 4296
rect 3053 4284 3059 4376
rect 3165 4304 3171 4436
rect 3197 4304 3203 4436
rect 3133 4284 3139 4296
rect 3037 4184 3043 4256
rect 3021 4177 3036 4183
rect 3021 4164 3027 4177
rect 3037 3924 3043 3996
rect 2861 3684 2867 3756
rect 2893 3743 2899 3876
rect 3053 3864 3059 4276
rect 3245 4264 3251 4536
rect 3277 4304 3283 4516
rect 3293 4344 3299 4536
rect 3373 4524 3379 4536
rect 3421 4504 3427 4636
rect 3485 4624 3491 4694
rect 3437 4584 3443 4616
rect 3485 4544 3491 4596
rect 3517 4564 3523 4676
rect 3549 4584 3555 4676
rect 3629 4604 3635 4716
rect 3661 4684 3667 4696
rect 3821 4684 3827 4696
rect 3677 4644 3683 4676
rect 3709 4644 3715 4680
rect 3853 4644 3859 4676
rect 3757 4544 3763 4556
rect 3853 4544 3859 4576
rect 3917 4564 3923 4656
rect 4045 4644 4051 4716
rect 4333 4704 4339 4716
rect 3293 4284 3299 4336
rect 3373 4284 3379 4456
rect 3421 4384 3427 4436
rect 3437 4323 3443 4496
rect 3485 4464 3491 4536
rect 3428 4317 3443 4323
rect 3133 4184 3139 4256
rect 3149 4164 3155 4236
rect 3197 4144 3203 4256
rect 3245 4164 3251 4216
rect 3261 4144 3267 4276
rect 3277 4224 3283 4256
rect 3389 4224 3395 4296
rect 3501 4284 3507 4496
rect 3533 4364 3539 4476
rect 3549 4384 3555 4516
rect 3565 4424 3571 4536
rect 3629 4524 3635 4536
rect 3581 4484 3587 4516
rect 3629 4424 3635 4496
rect 3533 4324 3539 4356
rect 3533 4304 3539 4316
rect 3629 4302 3635 4336
rect 3693 4304 3699 4536
rect 3789 4384 3795 4516
rect 3277 4184 3283 4216
rect 3304 4206 3310 4214
rect 3318 4206 3324 4214
rect 3332 4206 3338 4214
rect 3346 4206 3352 4214
rect 2957 3844 2963 3856
rect 2893 3737 2915 3743
rect 2909 3584 2915 3737
rect 2925 3724 2931 3736
rect 2557 3477 2572 3483
rect 2109 3084 2115 3096
rect 2253 3084 2259 3096
rect 1901 2944 1907 2956
rect 1933 2944 1939 2996
rect 1949 2943 1955 2956
rect 1949 2937 1964 2943
rect 1917 2624 1923 2636
rect 1965 2624 1971 2836
rect 1981 2704 1987 2996
rect 2093 2964 2099 3056
rect 2013 2944 2019 2956
rect 1997 2924 2003 2936
rect 1997 2664 2003 2696
rect 1997 2644 2003 2656
rect 2061 2524 2067 2856
rect 2077 2844 2083 2896
rect 2141 2884 2147 2916
rect 2285 2904 2291 2936
rect 2301 2924 2307 3096
rect 2333 2984 2339 3076
rect 2077 2724 2083 2816
rect 2093 2724 2099 2856
rect 2125 2664 2131 2836
rect 2164 2697 2179 2703
rect 2077 2524 2083 2636
rect 2125 2564 2131 2656
rect 2141 2543 2147 2676
rect 2173 2584 2179 2697
rect 2189 2684 2195 2696
rect 2189 2637 2204 2643
rect 2189 2564 2195 2637
rect 2237 2584 2243 2896
rect 2317 2884 2323 2936
rect 2333 2904 2339 2916
rect 2333 2724 2339 2896
rect 2349 2844 2355 3136
rect 2429 3124 2435 3276
rect 2445 3184 2451 3276
rect 2461 3084 2467 3336
rect 2541 3124 2547 3356
rect 2557 3304 2563 3477
rect 2605 3344 2611 3436
rect 2669 3364 2675 3376
rect 2557 3264 2563 3296
rect 2605 3084 2611 3336
rect 2749 3323 2755 3476
rect 2781 3444 2787 3476
rect 2740 3317 2755 3323
rect 2637 3064 2643 3116
rect 2733 3084 2739 3316
rect 2477 3044 2483 3056
rect 2397 3023 2403 3036
rect 2429 3024 2435 3036
rect 2397 3017 2419 3023
rect 2413 2964 2419 3017
rect 2413 2904 2419 2956
rect 2477 2944 2483 2976
rect 2445 2824 2451 2836
rect 2461 2824 2467 2936
rect 2509 2884 2515 2896
rect 2333 2664 2339 2696
rect 2132 2537 2147 2543
rect 2109 2524 2115 2536
rect 1997 2424 2003 2518
rect 1917 2302 1923 2316
rect 2125 2303 2131 2536
rect 2189 2504 2195 2556
rect 2205 2544 2211 2556
rect 2333 2544 2339 2656
rect 2397 2564 2403 2636
rect 2477 2584 2483 2696
rect 2493 2564 2499 2816
rect 2509 2684 2515 2876
rect 2541 2804 2547 3036
rect 2733 2984 2739 3076
rect 2685 2944 2691 2976
rect 2653 2926 2659 2936
rect 2749 2924 2755 3016
rect 2765 2944 2771 3256
rect 2797 3144 2803 3436
rect 2861 3284 2867 3296
rect 2829 3144 2835 3216
rect 2717 2904 2723 2916
rect 2525 2702 2531 2736
rect 2589 2704 2595 2716
rect 2637 2704 2643 2796
rect 2797 2784 2803 3136
rect 2829 3124 2835 3136
rect 2845 3104 2851 3256
rect 2861 3084 2867 3116
rect 2829 2964 2835 3036
rect 2861 2964 2867 3076
rect 2877 3063 2883 3536
rect 2893 3364 2899 3496
rect 2941 3484 2947 3736
rect 2957 3664 2963 3716
rect 2973 3523 2979 3836
rect 3037 3724 3043 3756
rect 3037 3524 3043 3716
rect 3069 3704 3075 4096
rect 3117 3904 3123 4016
rect 3309 3924 3315 4096
rect 3117 3803 3123 3896
rect 3261 3884 3267 3896
rect 3108 3797 3123 3803
rect 3101 3744 3107 3796
rect 3053 3697 3068 3703
rect 3053 3524 3059 3697
rect 2964 3517 2979 3523
rect 3117 3502 3123 3536
rect 2909 3344 2915 3476
rect 2957 3384 2963 3436
rect 2941 3377 2956 3383
rect 2941 3364 2947 3377
rect 2893 3304 2899 3316
rect 2957 3104 2963 3356
rect 2877 3057 2892 3063
rect 2909 3044 2915 3076
rect 2813 2924 2819 2956
rect 2877 2944 2883 3036
rect 2893 2977 2908 2983
rect 2893 2964 2899 2977
rect 2765 2704 2771 2716
rect 2829 2704 2835 2936
rect 2893 2924 2899 2956
rect 2445 2544 2451 2556
rect 2237 2504 2243 2516
rect 2317 2504 2323 2516
rect 2141 2323 2147 2436
rect 2141 2317 2156 2323
rect 2116 2297 2131 2303
rect 1981 2244 1987 2256
rect 1821 2124 1827 2136
rect 1768 2006 1774 2014
rect 1782 2006 1788 2014
rect 1796 2006 1802 2014
rect 1810 2006 1816 2014
rect 1565 1864 1571 1876
rect 1741 1864 1747 1896
rect 1213 1764 1219 1836
rect 1261 1824 1267 1836
rect 605 1664 611 1696
rect 637 1584 643 1636
rect 685 1584 691 1696
rect 717 1664 723 1676
rect 813 1644 819 1676
rect 685 1524 691 1576
rect 621 1484 627 1496
rect 557 1464 563 1476
rect 445 1457 467 1463
rect 317 1384 323 1456
rect 333 1364 339 1436
rect 397 1384 403 1456
rect 413 1364 419 1436
rect 381 1324 387 1336
rect 365 1284 371 1316
rect 413 1304 419 1356
rect 445 1344 451 1457
rect 461 1344 467 1436
rect 269 1124 275 1156
rect 205 1017 227 1023
rect 205 964 211 1017
rect 269 984 275 1116
rect 285 1104 291 1116
rect 317 1103 323 1276
rect 349 1184 355 1256
rect 317 1097 339 1103
rect 285 1064 291 1096
rect 333 984 339 1097
rect 20 917 35 923
rect 29 784 35 917
rect 77 784 83 936
rect 157 784 163 856
rect 205 824 211 956
rect 301 924 307 936
rect 317 924 323 936
rect 237 884 243 916
rect 253 904 259 916
rect 301 903 307 916
rect 301 897 323 903
rect 269 884 275 896
rect 221 764 227 876
rect 253 784 259 816
rect 61 724 67 736
rect 237 724 243 736
rect 301 724 307 836
rect 29 684 35 696
rect 61 584 67 716
rect 125 644 131 716
rect 157 684 163 696
rect 141 664 147 676
rect 221 664 227 716
rect 157 644 163 656
rect 109 544 115 576
rect 13 524 19 536
rect 125 504 131 516
rect 13 384 19 496
rect 157 384 163 636
rect 237 584 243 716
rect 189 564 195 576
rect 221 384 227 536
rect 237 504 243 556
rect 253 404 259 556
rect 285 544 291 696
rect 301 564 307 636
rect 317 584 323 897
rect 349 903 355 1016
rect 365 1004 371 1136
rect 397 1084 403 1156
rect 413 1104 419 1296
rect 429 1164 435 1236
rect 429 1124 435 1136
rect 445 1124 451 1276
rect 461 1084 467 1316
rect 477 1304 483 1316
rect 541 1304 547 1356
rect 557 1304 563 1456
rect 589 1444 595 1476
rect 653 1464 659 1496
rect 669 1464 675 1476
rect 749 1464 755 1596
rect 765 1464 771 1516
rect 573 1384 579 1436
rect 605 1324 611 1436
rect 493 1104 499 1236
rect 541 1124 547 1296
rect 621 1284 627 1416
rect 797 1403 803 1576
rect 845 1544 851 1696
rect 877 1604 883 1716
rect 893 1704 899 1716
rect 957 1704 963 1736
rect 973 1704 979 1716
rect 829 1504 835 1516
rect 861 1504 867 1516
rect 877 1484 883 1556
rect 893 1484 899 1696
rect 941 1584 947 1636
rect 957 1564 963 1656
rect 781 1397 803 1403
rect 765 1344 771 1396
rect 781 1364 787 1397
rect 861 1384 867 1476
rect 909 1444 915 1536
rect 941 1524 947 1536
rect 925 1484 931 1496
rect 957 1484 963 1556
rect 973 1504 979 1516
rect 781 1344 787 1356
rect 685 1324 691 1336
rect 797 1324 803 1376
rect 605 1264 611 1276
rect 557 1124 563 1236
rect 685 1184 691 1296
rect 557 1084 563 1116
rect 621 1084 627 1176
rect 717 1104 723 1116
rect 413 1024 419 1036
rect 365 984 371 996
rect 365 924 371 936
rect 340 897 355 903
rect 333 684 339 716
rect 349 704 355 756
rect 365 684 371 896
rect 381 883 387 936
rect 397 904 403 916
rect 413 904 419 916
rect 381 877 403 883
rect 333 584 339 676
rect 397 664 403 877
rect 413 784 419 876
rect 285 524 291 536
rect 381 524 387 636
rect 397 624 403 656
rect 429 544 435 736
rect 445 724 451 1036
rect 493 944 499 956
rect 525 924 531 1036
rect 509 904 515 916
rect 541 904 547 976
rect 557 964 563 1056
rect 557 944 563 956
rect 605 924 611 996
rect 573 904 579 916
rect 477 784 483 896
rect 509 784 515 836
rect 557 784 563 876
rect 525 724 531 736
rect 573 724 579 736
rect 77 324 83 336
rect 157 264 163 296
rect 173 284 179 316
rect 13 164 19 256
rect 77 184 83 236
rect 93 163 99 236
rect 157 184 163 256
rect 77 157 99 163
rect 77 104 83 157
rect 189 144 195 376
rect 205 324 211 336
rect 205 124 211 316
rect 221 304 227 356
rect 237 324 243 396
rect 285 384 291 496
rect 349 484 355 496
rect 365 484 371 516
rect 413 484 419 516
rect 237 163 243 316
rect 285 304 291 356
rect 301 324 307 476
rect 317 324 323 456
rect 381 444 387 476
rect 397 344 403 356
rect 413 344 419 416
rect 429 364 435 476
rect 445 424 451 516
rect 461 504 467 636
rect 525 563 531 716
rect 541 664 547 716
rect 557 684 563 696
rect 557 584 563 616
rect 525 557 540 563
rect 573 544 579 716
rect 589 544 595 836
rect 621 704 627 936
rect 685 924 691 1036
rect 701 963 707 976
rect 717 963 723 1036
rect 701 957 723 963
rect 701 944 707 957
rect 669 724 675 736
rect 653 684 659 696
rect 685 584 691 836
rect 701 744 707 916
rect 717 904 723 936
rect 733 924 739 1196
rect 813 1184 819 1336
rect 941 1324 947 1336
rect 749 1084 755 1136
rect 813 1104 819 1116
rect 829 884 835 1156
rect 861 1124 867 1256
rect 877 1124 883 1296
rect 893 1144 899 1236
rect 861 1104 867 1116
rect 877 1084 883 1096
rect 909 1084 915 1116
rect 925 1104 931 1296
rect 941 1124 947 1316
rect 989 1304 995 1736
rect 1085 1724 1091 1736
rect 1149 1724 1155 1756
rect 1005 1524 1011 1696
rect 1021 1624 1027 1696
rect 1085 1664 1091 1716
rect 1117 1684 1123 1696
rect 1133 1664 1139 1696
rect 1245 1684 1251 1696
rect 1261 1684 1267 1716
rect 1293 1704 1299 1756
rect 1309 1724 1315 1836
rect 1357 1804 1363 1856
rect 1517 1824 1523 1856
rect 1325 1744 1331 1756
rect 1421 1724 1427 1796
rect 1533 1744 1539 1836
rect 1277 1664 1283 1696
rect 1085 1584 1091 1636
rect 1005 1324 1011 1356
rect 1021 1324 1027 1576
rect 1037 1484 1043 1556
rect 1085 1504 1091 1536
rect 1069 1464 1075 1476
rect 1101 1464 1107 1516
rect 1133 1503 1139 1656
rect 1149 1564 1155 1636
rect 1165 1524 1171 1536
rect 1133 1497 1148 1503
rect 1213 1463 1219 1556
rect 1261 1543 1267 1636
rect 1309 1604 1315 1636
rect 1325 1624 1331 1636
rect 1245 1537 1267 1543
rect 1229 1504 1235 1536
rect 1245 1504 1251 1537
rect 1277 1523 1283 1596
rect 1325 1523 1331 1616
rect 1268 1517 1283 1523
rect 1277 1504 1283 1517
rect 1309 1517 1331 1523
rect 1245 1484 1251 1496
rect 1197 1457 1219 1463
rect 1037 1384 1043 1436
rect 1069 1363 1075 1376
rect 1060 1357 1075 1363
rect 1117 1343 1123 1436
rect 1101 1337 1123 1343
rect 957 1244 963 1276
rect 973 1164 979 1236
rect 989 1143 995 1296
rect 1005 1204 1011 1236
rect 973 1137 995 1143
rect 925 1084 931 1096
rect 973 1084 979 1137
rect 877 1004 883 1036
rect 861 924 867 976
rect 909 904 915 936
rect 925 924 931 976
rect 941 884 947 916
rect 701 664 707 676
rect 701 544 707 616
rect 525 504 531 516
rect 461 464 467 496
rect 477 477 492 483
rect 477 444 483 477
rect 509 464 515 476
rect 477 384 483 436
rect 525 404 531 496
rect 573 484 579 536
rect 733 523 739 836
rect 813 764 819 836
rect 829 684 835 776
rect 765 564 771 636
rect 733 517 748 523
rect 589 504 595 516
rect 765 504 771 536
rect 781 504 787 576
rect 349 324 355 336
rect 317 304 323 316
rect 269 164 275 296
rect 333 264 339 296
rect 317 257 332 263
rect 221 157 243 163
rect 221 144 227 157
rect 317 124 323 257
rect 349 144 355 316
rect 413 304 419 336
rect 445 323 451 376
rect 436 317 451 323
rect 541 304 547 376
rect 557 344 563 396
rect 589 344 595 396
rect 564 317 595 323
rect 477 264 483 296
rect 589 283 595 317
rect 605 304 611 376
rect 621 324 627 356
rect 653 344 659 416
rect 717 384 723 436
rect 797 384 803 436
rect 733 344 739 376
rect 797 344 803 376
rect 669 304 675 336
rect 765 324 771 336
rect 829 324 835 656
rect 845 643 851 756
rect 861 744 867 836
rect 925 744 931 836
rect 957 743 963 1036
rect 989 943 995 1036
rect 1005 984 1011 1156
rect 1021 1084 1027 1096
rect 1037 1064 1043 1116
rect 1037 1004 1043 1036
rect 1053 1024 1059 1316
rect 1085 1284 1091 1296
rect 1085 1184 1091 1276
rect 1069 1084 1075 1136
rect 980 937 995 943
rect 973 904 979 936
rect 1005 923 1011 956
rect 1053 924 1059 996
rect 996 917 1011 923
rect 1021 904 1027 916
rect 1037 864 1043 896
rect 1085 883 1091 1036
rect 1101 1004 1107 1337
rect 1133 1324 1139 1376
rect 1197 1304 1203 1457
rect 1213 1424 1219 1436
rect 1213 1344 1219 1376
rect 1213 1284 1219 1336
rect 1245 1304 1251 1336
rect 1117 1164 1123 1236
rect 1117 1104 1123 1136
rect 1149 1104 1155 1156
rect 1165 1144 1171 1236
rect 1133 1064 1139 1076
rect 1165 944 1171 1076
rect 1213 1064 1219 1216
rect 1229 1184 1235 1236
rect 1229 1103 1235 1176
rect 1245 1144 1251 1296
rect 1277 1284 1283 1416
rect 1293 1404 1299 1436
rect 1293 1324 1299 1356
rect 1309 1304 1315 1517
rect 1341 1504 1347 1636
rect 1373 1624 1379 1716
rect 1405 1664 1411 1696
rect 1373 1564 1379 1616
rect 1405 1584 1411 1656
rect 1421 1544 1427 1636
rect 1437 1544 1443 1616
rect 1437 1524 1443 1536
rect 1485 1524 1491 1636
rect 1501 1604 1507 1736
rect 1485 1504 1491 1516
rect 1325 1484 1331 1496
rect 1389 1484 1395 1496
rect 1501 1484 1507 1596
rect 1325 1344 1331 1416
rect 1325 1304 1331 1336
rect 1261 1164 1267 1236
rect 1277 1124 1283 1276
rect 1309 1264 1315 1296
rect 1293 1104 1299 1136
rect 1229 1097 1244 1103
rect 1197 944 1203 996
rect 1101 904 1107 916
rect 1076 877 1091 883
rect 941 737 963 743
rect 941 684 947 737
rect 957 704 963 716
rect 845 637 867 643
rect 845 504 851 576
rect 861 524 867 637
rect 957 564 963 696
rect 973 684 979 756
rect 1005 664 1011 856
rect 1037 704 1043 796
rect 1085 724 1091 836
rect 1197 724 1203 896
rect 1213 764 1219 836
rect 1229 784 1235 1097
rect 1309 1103 1315 1256
rect 1373 1224 1379 1436
rect 1421 1344 1427 1356
rect 1469 1324 1475 1336
rect 1309 1097 1331 1103
rect 1325 1064 1331 1097
rect 1357 1084 1363 1116
rect 1373 1063 1379 1076
rect 1357 1057 1379 1063
rect 1284 1037 1299 1043
rect 1245 904 1251 976
rect 1261 904 1267 1036
rect 1293 1023 1299 1037
rect 1357 1023 1363 1057
rect 1293 1017 1363 1023
rect 1277 944 1283 1016
rect 1325 924 1331 956
rect 1389 944 1395 1276
rect 1469 1264 1475 1276
rect 1405 1064 1411 1236
rect 1421 1124 1427 1136
rect 1469 1104 1475 1116
rect 1453 1077 1468 1083
rect 1405 1004 1411 1036
rect 1453 964 1459 1077
rect 1485 1024 1491 1096
rect 1485 924 1491 1016
rect 1501 943 1507 1236
rect 1517 1204 1523 1556
rect 1549 1524 1555 1796
rect 1597 1784 1603 1836
rect 1613 1743 1619 1776
rect 1629 1764 1635 1836
rect 1693 1784 1699 1836
rect 1613 1737 1628 1743
rect 1549 1344 1555 1516
rect 1565 1484 1571 1576
rect 1613 1544 1619 1716
rect 1629 1604 1635 1736
rect 1677 1564 1683 1636
rect 1613 1484 1619 1536
rect 1661 1524 1667 1536
rect 1709 1484 1715 1596
rect 1741 1544 1747 1736
rect 1789 1704 1795 1956
rect 1821 1724 1827 1836
rect 1837 1744 1843 1876
rect 1853 1804 1859 1836
rect 1789 1664 1795 1696
rect 1768 1606 1774 1614
rect 1782 1606 1788 1614
rect 1796 1606 1802 1614
rect 1810 1606 1816 1614
rect 1869 1524 1875 2236
rect 1901 1924 1907 2036
rect 1885 1904 1891 1916
rect 1997 1884 2003 2296
rect 2013 2284 2019 2296
rect 2109 2284 2115 2296
rect 2077 2184 2083 2256
rect 2093 2144 2099 2176
rect 2157 2124 2163 2236
rect 2253 2144 2259 2296
rect 2333 2284 2339 2536
rect 2365 2244 2371 2256
rect 2381 2144 2387 2316
rect 2397 2284 2403 2456
rect 2445 2324 2451 2396
rect 2461 2324 2467 2516
rect 2477 2504 2483 2516
rect 2493 2464 2499 2556
rect 2509 2524 2515 2676
rect 2749 2664 2755 2676
rect 2621 2564 2627 2576
rect 2653 2524 2659 2576
rect 2509 2424 2515 2436
rect 2701 2344 2707 2636
rect 2749 2544 2755 2556
rect 2749 2484 2755 2496
rect 2461 2284 2467 2316
rect 2477 2304 2483 2336
rect 2733 2324 2739 2456
rect 2765 2324 2771 2696
rect 2813 2584 2819 2676
rect 2829 2664 2835 2696
rect 2861 2664 2867 2836
rect 2893 2784 2899 2816
rect 2925 2704 2931 2996
rect 2941 2724 2947 3036
rect 2957 3004 2963 3096
rect 3021 3084 3027 3476
rect 3053 3044 3059 3116
rect 3021 2944 3027 2976
rect 3005 2924 3011 2936
rect 3037 2804 3043 3036
rect 3085 2984 3091 3476
rect 3149 3384 3155 3876
rect 3245 3744 3251 3876
rect 3304 3806 3310 3814
rect 3318 3806 3324 3814
rect 3332 3806 3338 3814
rect 3346 3806 3352 3814
rect 3373 3784 3379 4076
rect 3389 4044 3395 4216
rect 3469 4144 3475 4236
rect 3485 4224 3491 4256
rect 3421 3784 3427 4036
rect 3437 4024 3443 4136
rect 3437 3844 3443 3876
rect 3268 3777 3283 3783
rect 3277 3764 3283 3777
rect 3517 3764 3523 4236
rect 3533 4124 3539 4236
rect 3565 4184 3571 4216
rect 3597 4184 3603 4256
rect 3741 4144 3747 4256
rect 3757 4164 3763 4236
rect 3773 4144 3779 4276
rect 3789 4123 3795 4296
rect 3869 4284 3875 4436
rect 3885 4284 3891 4316
rect 3853 4144 3859 4156
rect 3869 4144 3875 4176
rect 3773 4117 3795 4123
rect 3677 4104 3683 4116
rect 3565 3884 3571 4096
rect 3597 4084 3603 4096
rect 3661 3984 3667 4056
rect 3693 3923 3699 4036
rect 3684 3917 3699 3923
rect 3677 3904 3683 3916
rect 3629 3884 3635 3896
rect 3565 3864 3571 3876
rect 3533 3844 3539 3856
rect 3277 3724 3283 3756
rect 3389 3604 3395 3756
rect 3245 3584 3251 3596
rect 3261 3443 3267 3476
rect 3252 3437 3267 3443
rect 3304 3406 3310 3414
rect 3318 3406 3324 3414
rect 3332 3406 3338 3414
rect 3346 3406 3352 3414
rect 3165 3364 3171 3376
rect 3405 3344 3411 3576
rect 3421 3524 3427 3536
rect 3421 3464 3427 3516
rect 3437 3504 3443 3736
rect 3453 3584 3459 3696
rect 3469 3564 3475 3736
rect 3549 3724 3555 3796
rect 3565 3744 3571 3816
rect 3581 3724 3587 3836
rect 3645 3784 3651 3796
rect 3661 3764 3667 3776
rect 3613 3724 3619 3756
rect 3677 3704 3683 3716
rect 3469 3484 3475 3556
rect 3661 3544 3667 3696
rect 3693 3604 3699 3876
rect 3709 3724 3715 3956
rect 3741 3924 3747 4096
rect 3773 4044 3779 4117
rect 3805 4084 3811 4096
rect 3885 4084 3891 4276
rect 3901 4184 3907 4296
rect 3965 4284 3971 4516
rect 4061 4324 4067 4536
rect 4077 4524 4083 4636
rect 4109 4584 4115 4694
rect 4253 4624 4259 4676
rect 4077 4384 4083 4516
rect 4093 4184 4099 4276
rect 3917 4144 3923 4156
rect 4077 4144 4083 4156
rect 3885 3924 3891 4076
rect 3901 4064 3907 4096
rect 4045 4084 4051 4096
rect 3741 3824 3747 3916
rect 3789 3904 3795 3916
rect 3773 3864 3779 3896
rect 3805 3884 3811 3916
rect 3885 3884 3891 3916
rect 3917 3884 3923 3936
rect 3981 3902 3987 3916
rect 3789 3744 3795 3836
rect 3725 3704 3731 3736
rect 3533 3502 3539 3516
rect 3117 3324 3123 3336
rect 3165 3324 3171 3336
rect 3229 3244 3235 3318
rect 3101 3184 3107 3236
rect 3149 3164 3155 3236
rect 3101 3104 3107 3156
rect 3133 3124 3139 3136
rect 3181 3064 3187 3076
rect 3261 3064 3267 3136
rect 3293 3084 3299 3316
rect 3389 3084 3395 3096
rect 3101 2964 3107 3036
rect 3304 3006 3310 3014
rect 3318 3006 3324 3014
rect 3332 3006 3338 3014
rect 3346 3006 3352 3014
rect 3373 2984 3379 3036
rect 3213 2944 3219 2976
rect 3133 2823 3139 2936
rect 3389 2904 3395 2916
rect 3181 2884 3187 2896
rect 3124 2817 3139 2823
rect 3117 2724 3123 2816
rect 3261 2724 3267 2876
rect 3437 2864 3443 3436
rect 3533 3384 3539 3456
rect 3581 3344 3587 3476
rect 3677 3464 3683 3516
rect 3725 3484 3731 3556
rect 3757 3464 3763 3536
rect 3789 3484 3795 3736
rect 3805 3724 3811 3756
rect 3949 3744 3955 3876
rect 3997 3724 4003 4036
rect 4077 3804 4083 4136
rect 4093 4084 4099 4096
rect 4109 3944 4115 4516
rect 4125 4264 4131 4536
rect 4253 4524 4259 4616
rect 4301 4584 4307 4656
rect 4333 4544 4339 4696
rect 4365 4684 4371 4696
rect 4445 4644 4451 4716
rect 4525 4704 4531 4716
rect 4269 4484 4275 4536
rect 4301 4504 4307 4536
rect 4349 4504 4355 4636
rect 4381 4583 4387 4636
rect 4381 4577 4403 4583
rect 4372 4557 4387 4563
rect 4381 4544 4387 4557
rect 4141 4344 4147 4476
rect 4141 4284 4147 4316
rect 4157 4304 4163 4336
rect 4237 4304 4243 4436
rect 4365 4324 4371 4536
rect 4397 4524 4403 4577
rect 4381 4484 4387 4516
rect 4397 4364 4403 4516
rect 4461 4504 4467 4696
rect 4477 4524 4483 4676
rect 4445 4304 4451 4496
rect 4477 4464 4483 4516
rect 4493 4484 4499 4596
rect 4509 4584 4515 4676
rect 4525 4543 4531 4696
rect 4573 4584 4579 4636
rect 4589 4624 4595 4656
rect 4605 4564 4611 4636
rect 4509 4537 4531 4543
rect 4509 4424 4515 4537
rect 4525 4504 4531 4516
rect 4541 4504 4547 4516
rect 4541 4483 4547 4496
rect 4525 4477 4547 4483
rect 4477 4384 4483 4416
rect 4525 4344 4531 4477
rect 4541 4384 4547 4416
rect 4189 4284 4195 4296
rect 4317 4284 4323 4296
rect 4148 4277 4163 4283
rect 4125 4224 4131 4236
rect 4125 4144 4131 4216
rect 4141 4164 4147 4236
rect 4157 4144 4163 4277
rect 4205 4144 4211 4196
rect 4157 4084 4163 4136
rect 4189 3964 4195 4036
rect 4221 3884 4227 4276
rect 4365 4164 4371 4276
rect 4413 4204 4419 4236
rect 4429 4164 4435 4276
rect 4269 4124 4275 4136
rect 4477 4124 4483 4296
rect 4509 4184 4515 4296
rect 4493 4144 4499 4176
rect 4525 4104 4531 4336
rect 4573 4304 4579 4536
rect 4589 4484 4595 4536
rect 4605 4504 4611 4516
rect 4605 4324 4611 4496
rect 4621 4464 4627 4696
rect 4717 4664 4723 4676
rect 4781 4664 4787 4696
rect 4637 4524 4643 4656
rect 4733 4624 4739 4656
rect 4813 4624 4819 4716
rect 4877 4704 4883 4716
rect 4685 4584 4691 4596
rect 4829 4584 4835 4656
rect 4893 4644 4899 4696
rect 4925 4684 4931 4716
rect 4941 4664 4947 4676
rect 4957 4644 4963 4696
rect 5005 4664 5011 4717
rect 5021 4717 5036 4723
rect 5021 4664 5027 4717
rect 5069 4703 5075 4756
rect 5085 4724 5091 4756
rect 5117 4724 5123 4736
rect 5165 4724 5171 4736
rect 5181 4704 5187 4756
rect 5197 4724 5203 4736
rect 5069 4697 5091 4703
rect 5069 4664 5075 4676
rect 5085 4643 5091 4697
rect 5101 4684 5107 4696
rect 5213 4684 5219 4736
rect 5517 4724 5523 4736
rect 5716 4717 5731 4723
rect 5117 4643 5123 4656
rect 5085 4637 5123 4643
rect 4989 4584 4995 4616
rect 5053 4584 5059 4636
rect 5165 4584 5171 4636
rect 4717 4544 4723 4556
rect 4813 4544 4819 4556
rect 4701 4537 4716 4543
rect 4653 4484 4659 4496
rect 4621 4344 4627 4436
rect 4685 4424 4691 4496
rect 4701 4384 4707 4537
rect 4717 4363 4723 4516
rect 4708 4357 4723 4363
rect 4605 4304 4611 4316
rect 4573 4284 4579 4296
rect 4621 4284 4627 4336
rect 4557 4144 4563 4156
rect 4541 4124 4547 4136
rect 4541 4103 4547 4116
rect 4541 4097 4556 4103
rect 4269 4084 4275 4096
rect 4109 3784 4115 3796
rect 4061 3524 4067 3596
rect 3453 3144 3459 3176
rect 3581 3104 3587 3336
rect 3853 3324 3859 3456
rect 4029 3444 4035 3496
rect 4061 3464 4067 3516
rect 4093 3484 4099 3536
rect 4109 3504 4115 3736
rect 4125 3704 4131 3776
rect 4141 3724 4147 3756
rect 4157 3704 4163 3836
rect 3981 3363 3987 3436
rect 3981 3357 4003 3363
rect 3901 3344 3907 3356
rect 3997 3324 4003 3357
rect 3869 3304 3875 3316
rect 3693 3124 3699 3216
rect 3757 3144 3763 3236
rect 3533 2944 3539 3056
rect 3549 2964 3555 3096
rect 3581 2983 3587 3096
rect 3661 3084 3667 3096
rect 3709 3084 3715 3136
rect 3805 3084 3811 3276
rect 3581 2977 3603 2983
rect 3565 2964 3571 2976
rect 3597 2944 3603 2977
rect 3533 2924 3539 2936
rect 3629 2926 3635 2936
rect 3469 2884 3475 2896
rect 3044 2717 3059 2723
rect 2797 2564 2803 2576
rect 2829 2564 2835 2656
rect 2781 2504 2787 2516
rect 2829 2504 2835 2516
rect 2845 2503 2851 2556
rect 2877 2544 2883 2556
rect 2957 2544 2963 2716
rect 3053 2704 3059 2717
rect 3101 2704 3107 2716
rect 3213 2704 3219 2716
rect 2989 2664 2995 2676
rect 2973 2604 2979 2636
rect 2989 2583 2995 2656
rect 3037 2624 3043 2696
rect 3133 2684 3139 2696
rect 3245 2684 3251 2716
rect 3053 2584 3059 2676
rect 2980 2577 2995 2583
rect 2893 2524 2899 2536
rect 2836 2497 2851 2503
rect 2861 2364 2867 2516
rect 2909 2504 2915 2516
rect 2685 2304 2691 2316
rect 2045 1924 2051 1956
rect 2173 1884 2179 1996
rect 2205 1884 2211 2136
rect 2317 2124 2323 2136
rect 2381 2104 2387 2136
rect 1757 1504 1763 1516
rect 1917 1484 1923 1836
rect 1949 1584 1955 1876
rect 1997 1864 2003 1876
rect 1965 1784 1971 1856
rect 2045 1784 2051 1836
rect 2077 1804 2083 1876
rect 1981 1726 1987 1776
rect 2125 1724 2131 1836
rect 2221 1784 2227 1796
rect 2253 1784 2259 1876
rect 2253 1724 2259 1776
rect 2221 1564 2227 1636
rect 1933 1484 1939 1516
rect 1981 1504 1987 1516
rect 2061 1504 2067 1536
rect 2093 1484 2099 1516
rect 2125 1484 2131 1536
rect 2173 1484 2179 1536
rect 2269 1523 2275 1536
rect 2253 1517 2275 1523
rect 2349 1523 2355 1876
rect 2365 1744 2371 1916
rect 2445 1904 2451 1976
rect 2461 1884 2467 2136
rect 2493 2124 2499 2276
rect 2557 2183 2563 2276
rect 2573 2204 2579 2276
rect 2557 2177 2572 2183
rect 2365 1684 2371 1736
rect 2445 1724 2451 1876
rect 2349 1517 2371 1523
rect 2205 1483 2211 1516
rect 2253 1504 2259 1517
rect 2189 1477 2211 1483
rect 1565 1424 1571 1476
rect 1661 1424 1667 1436
rect 1661 1344 1667 1356
rect 1677 1344 1683 1436
rect 1533 1284 1539 1316
rect 1556 1277 1571 1283
rect 1565 1144 1571 1277
rect 1517 1064 1523 1076
rect 1517 964 1523 996
rect 1533 984 1539 1116
rect 1565 1084 1571 1136
rect 1597 1123 1603 1236
rect 1629 1124 1635 1276
rect 1588 1117 1603 1123
rect 1581 1104 1587 1116
rect 1629 1084 1635 1116
rect 1565 1064 1571 1076
rect 1501 937 1523 943
rect 1373 904 1379 916
rect 1309 884 1315 896
rect 1341 884 1347 896
rect 1293 804 1299 836
rect 1085 704 1091 716
rect 877 484 883 556
rect 925 484 931 556
rect 973 544 979 636
rect 957 504 963 536
rect 989 464 995 636
rect 1005 544 1011 656
rect 1021 584 1027 676
rect 1037 624 1043 696
rect 1133 684 1139 696
rect 1149 684 1155 696
rect 1181 644 1187 656
rect 1085 604 1091 636
rect 701 283 707 316
rect 717 304 723 316
rect 781 304 787 316
rect 589 277 803 283
rect 797 264 803 277
rect 365 184 371 196
rect 445 164 451 216
rect 493 184 499 236
rect 365 124 371 156
rect 413 144 419 156
rect 381 137 396 143
rect 381 104 387 137
rect 397 124 403 136
rect 445 84 451 156
rect 493 104 499 156
rect 525 84 531 176
rect 637 144 643 236
rect 813 223 819 276
rect 765 217 819 223
rect 541 84 547 116
rect 653 84 659 176
rect 733 144 739 196
rect 669 84 675 116
rect 749 104 755 196
rect 765 144 771 217
rect 829 164 835 236
rect 845 204 851 416
rect 861 404 867 436
rect 893 303 899 456
rect 909 324 915 436
rect 957 344 963 396
rect 989 344 995 436
rect 973 304 979 316
rect 893 297 908 303
rect 989 284 995 336
rect 1037 324 1043 516
rect 1053 484 1059 516
rect 1085 504 1091 556
rect 1181 524 1187 596
rect 1197 564 1203 716
rect 1101 324 1107 516
rect 1117 484 1123 516
rect 1197 504 1203 516
rect 1021 317 1036 323
rect 1021 264 1027 317
rect 1133 284 1139 336
rect 1149 324 1155 436
rect 1021 217 1091 223
rect 1021 204 1027 217
rect 845 144 851 156
rect 797 124 803 136
rect 813 104 819 136
rect 861 124 867 196
rect 1037 144 1043 196
rect 1085 164 1091 217
rect 1101 144 1107 196
rect 1117 164 1123 256
rect 1149 244 1155 256
rect 1165 243 1171 476
rect 1197 304 1203 496
rect 1213 324 1219 596
rect 1229 564 1235 696
rect 1229 524 1235 556
rect 1245 504 1251 776
rect 1261 664 1267 716
rect 1293 684 1299 776
rect 1309 704 1315 716
rect 1341 704 1347 716
rect 1357 664 1363 896
rect 1389 704 1395 756
rect 1405 724 1411 756
rect 1421 744 1427 896
rect 1437 744 1443 916
rect 1517 744 1523 937
rect 1533 784 1539 876
rect 1421 724 1427 736
rect 1453 664 1459 716
rect 1533 704 1539 716
rect 1261 544 1267 656
rect 1277 484 1283 636
rect 1357 604 1363 636
rect 1325 484 1331 576
rect 1341 484 1347 516
rect 1373 504 1379 596
rect 1389 524 1395 536
rect 1405 484 1411 556
rect 1261 344 1267 436
rect 1197 284 1203 296
rect 1213 284 1219 316
rect 1261 284 1267 316
rect 1293 284 1299 456
rect 1325 344 1331 476
rect 1389 424 1395 436
rect 1421 343 1427 616
rect 1549 584 1555 1016
rect 1565 924 1571 976
rect 1453 524 1459 536
rect 1437 484 1443 516
rect 1485 503 1491 556
rect 1517 524 1523 536
rect 1485 497 1500 503
rect 1412 337 1427 343
rect 1341 304 1347 336
rect 1389 304 1395 336
rect 1437 324 1443 356
rect 1485 304 1491 436
rect 1517 364 1523 436
rect 1501 284 1507 296
rect 1293 264 1299 276
rect 1533 264 1539 416
rect 1565 324 1571 836
rect 1581 784 1587 896
rect 1581 724 1587 776
rect 1597 724 1603 1036
rect 1629 1004 1635 1036
rect 1661 984 1667 1316
rect 1677 1104 1683 1236
rect 1693 1104 1699 1436
rect 1709 1384 1715 1476
rect 1725 1384 1731 1476
rect 1821 1464 1827 1476
rect 1853 1363 1859 1436
rect 1837 1357 1859 1363
rect 1757 1304 1763 1336
rect 1821 1284 1827 1296
rect 1768 1206 1774 1214
rect 1782 1206 1788 1214
rect 1796 1206 1802 1214
rect 1810 1206 1816 1214
rect 1837 1064 1843 1357
rect 1901 1344 1907 1436
rect 1917 1364 1923 1476
rect 1949 1424 1955 1436
rect 1933 1364 1939 1396
rect 1997 1344 2003 1396
rect 2013 1364 2019 1476
rect 2141 1444 2147 1456
rect 2157 1404 2163 1436
rect 2189 1384 2195 1477
rect 2253 1464 2259 1476
rect 2157 1364 2163 1376
rect 2013 1344 2019 1356
rect 2205 1344 2211 1356
rect 1853 1124 1859 1316
rect 1956 1297 1971 1303
rect 1885 1144 1891 1236
rect 1853 1084 1859 1116
rect 1933 1104 1939 1276
rect 1965 1184 1971 1297
rect 2061 1124 2067 1156
rect 1949 1064 1955 1116
rect 2061 1084 2067 1116
rect 2093 1104 2099 1336
rect 2125 1124 2131 1156
rect 2189 1144 2195 1236
rect 2205 1144 2211 1336
rect 2221 1324 2227 1356
rect 2253 1344 2259 1376
rect 2269 1304 2275 1496
rect 2301 1464 2307 1496
rect 2349 1484 2355 1496
rect 2365 1484 2371 1517
rect 2381 1484 2387 1556
rect 2445 1484 2451 1556
rect 2477 1484 2483 1516
rect 2301 1364 2307 1456
rect 2317 1384 2323 1436
rect 2301 1304 2307 1336
rect 2317 1304 2323 1316
rect 2269 1164 2275 1236
rect 2285 1184 2291 1276
rect 2093 1084 2099 1096
rect 1629 884 1635 956
rect 1613 744 1619 836
rect 1613 664 1619 736
rect 1645 684 1651 976
rect 1709 944 1715 1036
rect 1741 1024 1747 1036
rect 1677 884 1683 916
rect 1693 904 1699 916
rect 1741 884 1747 916
rect 1821 884 1827 896
rect 1581 484 1587 656
rect 1597 604 1603 636
rect 1613 577 1628 583
rect 1597 524 1603 536
rect 1613 504 1619 577
rect 1629 564 1635 576
rect 1661 564 1667 636
rect 1661 524 1667 536
rect 1677 524 1683 856
rect 1693 743 1699 836
rect 1693 737 1715 743
rect 1693 624 1699 636
rect 1677 483 1683 516
rect 1693 504 1699 576
rect 1709 524 1715 737
rect 1725 704 1731 876
rect 1757 844 1763 876
rect 1789 864 1795 876
rect 1821 864 1827 876
rect 1725 684 1731 696
rect 1741 544 1747 836
rect 1768 806 1774 814
rect 1782 806 1788 814
rect 1796 806 1802 814
rect 1810 806 1816 814
rect 1789 724 1795 776
rect 1757 704 1763 716
rect 1837 684 1843 896
rect 1853 884 1859 916
rect 1869 884 1875 936
rect 1853 844 1859 876
rect 1901 844 1907 956
rect 1997 944 2003 1036
rect 1965 884 1971 916
rect 1981 904 1987 916
rect 2061 904 2067 1036
rect 2093 924 2099 996
rect 2109 904 2115 1116
rect 2141 884 2147 976
rect 2157 924 2163 996
rect 2173 923 2179 1116
rect 2189 923 2195 956
rect 2205 924 2211 1036
rect 2221 964 2227 1136
rect 2301 1124 2307 1136
rect 2333 1104 2339 1336
rect 2349 1324 2355 1376
rect 2365 1364 2371 1476
rect 2381 1464 2387 1476
rect 2397 1424 2403 1436
rect 2397 1343 2403 1416
rect 2429 1364 2435 1396
rect 2397 1337 2419 1343
rect 2413 1324 2419 1337
rect 2173 917 2195 923
rect 2173 904 2179 917
rect 2253 904 2259 1076
rect 2301 1004 2307 1036
rect 2365 984 2371 1316
rect 2397 1124 2403 1196
rect 2429 1084 2435 1356
rect 2445 1344 2451 1436
rect 2461 1104 2467 1236
rect 2477 1204 2483 1476
rect 2525 1463 2531 1496
rect 2541 1484 2547 2096
rect 2557 1924 2563 1936
rect 2637 1904 2643 2276
rect 2733 2164 2739 2316
rect 2765 2304 2771 2316
rect 2781 2284 2787 2336
rect 2861 2323 2867 2356
rect 2893 2344 2899 2456
rect 2925 2344 2931 2536
rect 2941 2524 2947 2536
rect 3069 2464 3075 2556
rect 3117 2544 3123 2576
rect 3133 2524 3139 2616
rect 3149 2604 3155 2656
rect 3101 2484 3107 2516
rect 2925 2324 2931 2336
rect 2861 2317 2876 2323
rect 2813 2264 2819 2296
rect 2829 2244 2835 2276
rect 2893 2264 2899 2296
rect 2941 2264 2947 2436
rect 3133 2364 3139 2516
rect 3149 2503 3155 2596
rect 3261 2584 3267 2696
rect 3309 2664 3315 2676
rect 3405 2624 3411 2676
rect 3453 2644 3459 2656
rect 3304 2606 3310 2614
rect 3318 2606 3324 2614
rect 3332 2606 3338 2614
rect 3346 2606 3352 2614
rect 3149 2497 3164 2503
rect 3021 2304 3027 2316
rect 3101 2304 3107 2356
rect 3149 2304 3155 2336
rect 2957 2284 2963 2296
rect 2973 2244 2979 2256
rect 2877 2204 2883 2236
rect 3005 2224 3011 2296
rect 3069 2264 3075 2276
rect 3085 2224 3091 2276
rect 2813 2164 2819 2176
rect 2909 2164 2915 2176
rect 3037 2164 3043 2176
rect 2653 2124 2659 2136
rect 2813 2124 2819 2136
rect 2893 2124 2899 2156
rect 2941 2124 2947 2156
rect 2989 2144 2995 2156
rect 3021 2124 3027 2156
rect 3069 2124 3075 2136
rect 3085 2124 3091 2196
rect 3165 2184 3171 2316
rect 3181 2304 3187 2576
rect 3325 2544 3331 2556
rect 3197 2524 3203 2536
rect 3245 2524 3251 2536
rect 3437 2524 3443 2636
rect 3453 2524 3459 2536
rect 3197 2324 3203 2476
rect 3437 2404 3443 2516
rect 3485 2444 3491 2896
rect 3645 2824 3651 3036
rect 3549 2604 3555 2636
rect 3517 2564 3523 2576
rect 3565 2544 3571 2636
rect 3613 2544 3619 2676
rect 3629 2544 3635 2616
rect 3661 2584 3667 3076
rect 3821 3064 3827 3256
rect 3837 3084 3843 3156
rect 3853 3124 3859 3276
rect 3901 3144 3907 3316
rect 3917 3304 3923 3316
rect 4045 3304 4051 3456
rect 4109 3444 4115 3496
rect 4077 3344 4083 3436
rect 4093 3344 4099 3356
rect 4077 3324 4083 3336
rect 4093 3304 4099 3336
rect 4109 3324 4115 3376
rect 4125 3324 4131 3436
rect 4141 3424 4147 3636
rect 4173 3484 4179 3836
rect 4237 3784 4243 3916
rect 4269 3804 4275 3876
rect 4285 3864 4291 3896
rect 4301 3884 4307 3916
rect 4365 3904 4371 3916
rect 4573 3904 4579 4156
rect 4605 3944 4611 4136
rect 4637 4124 4643 4316
rect 4701 4304 4707 4356
rect 4733 4303 4739 4536
rect 4781 4504 4787 4536
rect 4797 4424 4803 4516
rect 4845 4504 4851 4536
rect 4941 4504 4947 4516
rect 4957 4484 4963 4576
rect 4824 4406 4830 4414
rect 4838 4406 4844 4414
rect 4852 4406 4858 4414
rect 4866 4406 4872 4414
rect 4781 4324 4787 4336
rect 4724 4297 4739 4303
rect 4669 4144 4675 4296
rect 4701 4264 4707 4296
rect 4717 4284 4723 4296
rect 4797 4284 4803 4296
rect 4717 4124 4723 4276
rect 4804 4257 4819 4263
rect 4733 4144 4739 4176
rect 4285 3844 4291 3856
rect 4221 3744 4227 3756
rect 4285 3744 4291 3816
rect 4269 3724 4275 3736
rect 4301 3723 4307 3876
rect 4333 3804 4339 3836
rect 4349 3824 4355 3876
rect 4365 3844 4371 3896
rect 4397 3864 4403 3876
rect 4301 3717 4323 3723
rect 4317 3704 4323 3717
rect 4333 3704 4339 3736
rect 4189 3684 4195 3696
rect 4189 3584 4195 3676
rect 4253 3564 4259 3636
rect 4317 3544 4323 3696
rect 4349 3584 4355 3716
rect 4365 3604 4371 3836
rect 4381 3743 4387 3836
rect 4397 3744 4403 3756
rect 4381 3737 4396 3743
rect 4413 3724 4419 3736
rect 4429 3663 4435 3876
rect 4573 3844 4579 3876
rect 4525 3804 4531 3836
rect 4605 3824 4611 3916
rect 4445 3724 4451 3796
rect 4468 3737 4483 3743
rect 4429 3657 4451 3663
rect 4157 3444 4163 3480
rect 4157 3404 4163 3436
rect 4125 3304 4131 3316
rect 3981 3124 3987 3256
rect 3885 3064 3891 3076
rect 3693 3004 3699 3036
rect 3805 2924 3811 3036
rect 3901 2964 3907 3036
rect 3917 3024 3923 3096
rect 3821 2924 3827 2936
rect 3773 2844 3779 2896
rect 3837 2744 3843 2876
rect 3885 2864 3891 2918
rect 3949 2884 3955 3036
rect 3965 3024 3971 3116
rect 3981 3104 3987 3116
rect 3997 3084 4003 3236
rect 4029 3084 4035 3176
rect 4045 3104 4051 3276
rect 4077 3104 4083 3236
rect 4093 3144 4099 3296
rect 4173 3284 4179 3476
rect 4221 3464 4227 3496
rect 4237 3484 4243 3496
rect 4189 3344 4195 3436
rect 4205 3344 4211 3396
rect 4205 3264 4211 3336
rect 4221 3244 4227 3456
rect 4237 3404 4243 3476
rect 4237 3244 4243 3296
rect 4253 3284 4259 3476
rect 4285 3444 4291 3516
rect 4317 3464 4323 3536
rect 4381 3524 4387 3536
rect 4333 3444 4339 3476
rect 4269 3364 4275 3436
rect 4285 3324 4291 3436
rect 4269 3284 4275 3316
rect 4317 3304 4323 3356
rect 4349 3324 4355 3496
rect 4397 3484 4403 3536
rect 4445 3524 4451 3657
rect 4477 3584 4483 3737
rect 4509 3724 4515 3776
rect 4541 3744 4547 3756
rect 4564 3737 4579 3743
rect 4557 3724 4563 3736
rect 4509 3584 4515 3636
rect 4557 3624 4563 3636
rect 4477 3524 4483 3576
rect 4557 3544 4563 3556
rect 4557 3504 4563 3536
rect 4365 3344 4371 3436
rect 4413 3344 4419 3496
rect 4493 3484 4499 3496
rect 4285 3284 4291 3296
rect 4173 3204 4179 3236
rect 4125 3124 4131 3196
rect 4173 3124 4179 3196
rect 4269 3144 4275 3276
rect 4285 3224 4291 3236
rect 4109 3097 4124 3103
rect 4093 3084 4099 3096
rect 4109 3063 4115 3097
rect 4036 3057 4115 3063
rect 4221 3024 4227 3116
rect 4237 3064 4243 3136
rect 4317 3084 4323 3256
rect 4333 3104 4339 3316
rect 4397 3204 4403 3276
rect 4413 3264 4419 3276
rect 4365 3144 4371 3196
rect 4413 3163 4419 3196
rect 4429 3164 4435 3476
rect 4541 3464 4547 3476
rect 4573 3344 4579 3737
rect 4589 3704 4595 3716
rect 4605 3524 4611 3776
rect 4621 3724 4627 3836
rect 4637 3724 4643 3956
rect 4653 3904 4659 4076
rect 4701 3923 4707 4116
rect 4685 3917 4707 3923
rect 4653 3884 4659 3896
rect 4669 3844 4675 3916
rect 4685 3784 4691 3917
rect 4717 3864 4723 4096
rect 4749 3904 4755 4136
rect 4765 4084 4771 4116
rect 4797 4104 4803 4196
rect 4813 4164 4819 4257
rect 4829 4184 4835 4376
rect 4941 4324 4947 4436
rect 4957 4384 4963 4456
rect 4989 4384 4995 4496
rect 4877 4284 4883 4316
rect 5005 4304 5011 4496
rect 5021 4464 5027 4536
rect 5021 4404 5027 4456
rect 5037 4384 5043 4536
rect 5149 4524 5155 4536
rect 5133 4484 5139 4516
rect 5181 4504 5187 4556
rect 5197 4544 5203 4676
rect 5245 4664 5251 4716
rect 5261 4704 5267 4716
rect 5245 4564 5251 4636
rect 5277 4564 5283 4696
rect 5309 4684 5315 4716
rect 5325 4704 5331 4716
rect 5293 4584 5299 4676
rect 5341 4644 5347 4716
rect 5277 4524 5283 4556
rect 5341 4544 5347 4596
rect 5357 4584 5363 4596
rect 5229 4484 5235 4516
rect 5101 4424 5107 4436
rect 5037 4264 5043 4296
rect 4941 4244 4947 4256
rect 4925 4164 4931 4236
rect 4941 4204 4947 4236
rect 4845 4144 4851 4156
rect 4813 4084 4819 4116
rect 4973 4064 4979 4096
rect 4765 3984 4771 4036
rect 4824 4006 4830 4014
rect 4838 4006 4844 4014
rect 4852 4006 4858 4014
rect 4866 4006 4872 4014
rect 4765 3904 4771 3916
rect 4797 3904 4803 3916
rect 4909 3904 4915 3916
rect 4925 3904 4931 4016
rect 4701 3744 4707 3856
rect 4717 3824 4723 3856
rect 4717 3724 4723 3816
rect 4637 3664 4643 3716
rect 4660 3697 4675 3703
rect 4621 3484 4627 3556
rect 4637 3524 4643 3636
rect 4653 3504 4659 3676
rect 4525 3324 4531 3336
rect 4445 3264 4451 3296
rect 4461 3264 4467 3316
rect 4397 3157 4419 3163
rect 4381 3124 4387 3156
rect 4397 3124 4403 3157
rect 4429 3123 4435 3156
rect 4429 3117 4451 3123
rect 4365 3083 4371 3116
rect 4397 3084 4403 3116
rect 4413 3104 4419 3116
rect 4429 3084 4435 3096
rect 4365 3077 4387 3083
rect 3997 3017 4083 3023
rect 3997 3004 4003 3017
rect 4077 3004 4083 3017
rect 4013 2984 4019 2996
rect 4013 2883 4019 2936
rect 4029 2904 4035 2976
rect 4061 2944 4067 2996
rect 4221 2984 4227 3016
rect 4381 3004 4387 3077
rect 4077 2924 4083 2956
rect 4061 2883 4067 2916
rect 4013 2877 4067 2883
rect 3693 2702 3699 2716
rect 3837 2704 3843 2736
rect 4077 2664 4083 2916
rect 4093 2664 4099 2736
rect 3661 2564 3667 2576
rect 3693 2544 3699 2656
rect 3581 2504 3587 2516
rect 3197 2304 3203 2316
rect 3293 2304 3299 2316
rect 3357 2304 3363 2356
rect 3181 2264 3187 2296
rect 3357 2264 3363 2276
rect 3213 2184 3219 2216
rect 3133 2144 3139 2156
rect 3101 2124 3107 2136
rect 2573 1664 2579 1736
rect 2605 1724 2611 1736
rect 2653 1724 2659 2036
rect 2813 1904 2819 2116
rect 2877 1984 2883 2036
rect 2701 1864 2707 1894
rect 2733 1843 2739 1876
rect 2765 1864 2771 1896
rect 2909 1884 2915 1956
rect 2925 1864 2931 1936
rect 2941 1904 2947 2116
rect 3053 1964 3059 2036
rect 3069 1984 3075 2096
rect 2989 1864 2995 1916
rect 3117 1904 3123 1976
rect 3037 1864 3043 1876
rect 3101 1864 3107 1876
rect 2733 1837 2755 1843
rect 2749 1744 2755 1837
rect 2877 1824 2883 1836
rect 2669 1724 2675 1736
rect 2573 1523 2579 1656
rect 2589 1524 2595 1536
rect 2637 1524 2643 1556
rect 2557 1517 2579 1523
rect 2557 1504 2563 1517
rect 2621 1504 2627 1516
rect 2509 1457 2531 1463
rect 2493 1324 2499 1336
rect 2509 1304 2515 1457
rect 2525 1304 2531 1436
rect 2541 1344 2547 1476
rect 2621 1464 2627 1476
rect 2509 1144 2515 1296
rect 2477 1124 2483 1136
rect 2557 1124 2563 1456
rect 2573 1284 2579 1356
rect 2621 1344 2627 1456
rect 2669 1424 2675 1496
rect 2685 1484 2691 1496
rect 2733 1483 2739 1516
rect 2781 1484 2787 1536
rect 2797 1504 2803 1776
rect 2813 1726 2819 1736
rect 2845 1664 2851 1736
rect 2909 1724 2915 1816
rect 2973 1744 2979 1776
rect 2941 1724 2947 1736
rect 2941 1704 2947 1716
rect 3005 1703 3011 1736
rect 3053 1724 3059 1756
rect 3069 1744 3075 1836
rect 3133 1763 3139 2036
rect 3149 1984 3155 2156
rect 3197 1984 3203 2156
rect 3149 1844 3155 1916
rect 3197 1904 3203 1936
rect 3229 1904 3235 2236
rect 3304 2206 3310 2214
rect 3318 2206 3324 2214
rect 3332 2206 3338 2214
rect 3346 2206 3352 2214
rect 3389 2184 3395 2296
rect 3405 2184 3411 2316
rect 3485 2304 3491 2316
rect 3501 2264 3507 2276
rect 3453 2184 3459 2256
rect 3421 2164 3427 2176
rect 3245 2124 3251 2136
rect 3309 2124 3315 2136
rect 3373 2124 3379 2156
rect 3261 1904 3267 1936
rect 3341 1884 3347 2116
rect 3405 2104 3411 2116
rect 3197 1764 3203 1836
rect 3124 1757 3139 1763
rect 3133 1724 3139 1757
rect 3181 1724 3187 1756
rect 3245 1744 3251 1836
rect 3261 1724 3267 1876
rect 3341 1864 3347 1876
rect 3437 1864 3443 1916
rect 3277 1844 3283 1856
rect 3405 1844 3411 1856
rect 3304 1806 3310 1814
rect 3318 1806 3324 1814
rect 3332 1806 3338 1814
rect 3346 1806 3352 1814
rect 3517 1764 3523 2496
rect 3613 2304 3619 2536
rect 3629 2504 3635 2536
rect 3677 2302 3683 2376
rect 3821 2364 3827 2636
rect 3869 2624 3875 2636
rect 3869 2524 3875 2616
rect 3917 2544 3923 2576
rect 3533 2264 3539 2276
rect 3549 2244 3555 2256
rect 3581 2144 3587 2296
rect 3613 2144 3619 2156
rect 3581 1864 3587 2136
rect 3645 2104 3651 2156
rect 3741 2144 3747 2236
rect 3661 2124 3667 2136
rect 3757 2124 3763 2236
rect 3773 2144 3779 2280
rect 3789 2244 3795 2276
rect 3837 2264 3843 2496
rect 3837 2104 3843 2256
rect 3853 2124 3859 2236
rect 3869 2164 3875 2516
rect 3885 2304 3891 2536
rect 3933 2524 3939 2556
rect 3997 2504 4003 2536
rect 4013 2504 4019 2536
rect 4061 2524 4067 2576
rect 4077 2564 4083 2616
rect 4093 2543 4099 2616
rect 4109 2564 4115 2856
rect 4125 2704 4131 2836
rect 4141 2824 4147 2956
rect 4253 2944 4259 2996
rect 4365 2944 4371 2996
rect 4445 2924 4451 3117
rect 4461 3104 4467 3236
rect 4477 3224 4483 3276
rect 4525 3224 4531 3276
rect 4541 3264 4547 3316
rect 4573 3303 4579 3336
rect 4589 3304 4595 3416
rect 4621 3304 4627 3436
rect 4653 3424 4659 3476
rect 4669 3364 4675 3697
rect 4701 3484 4707 3716
rect 4733 3703 4739 3876
rect 4749 3864 4755 3876
rect 4813 3864 4819 3876
rect 4941 3844 4947 3916
rect 4957 3904 4963 3916
rect 4989 3884 4995 4096
rect 5005 4083 5011 4256
rect 5069 4184 5075 4316
rect 5085 4304 5091 4316
rect 5117 4264 5123 4296
rect 5117 4224 5123 4256
rect 5149 4184 5155 4456
rect 5245 4424 5251 4496
rect 5309 4444 5315 4536
rect 5373 4504 5379 4676
rect 5421 4664 5427 4716
rect 5565 4684 5571 4696
rect 5437 4664 5443 4676
rect 5421 4624 5427 4656
rect 5501 4584 5507 4656
rect 5549 4564 5555 4636
rect 5565 4584 5571 4636
rect 5597 4604 5603 4656
rect 5629 4604 5635 4676
rect 5725 4664 5731 4717
rect 5821 4664 5827 4696
rect 5885 4684 5891 4696
rect 5805 4644 5811 4656
rect 5645 4584 5651 4616
rect 5709 4584 5715 4636
rect 5261 4364 5267 4436
rect 5165 4304 5171 4356
rect 5229 4324 5235 4336
rect 5261 4303 5267 4356
rect 5293 4304 5299 4376
rect 5325 4363 5331 4436
rect 5325 4357 5347 4363
rect 5341 4324 5347 4357
rect 5341 4304 5347 4316
rect 5252 4297 5267 4303
rect 5197 4264 5203 4276
rect 5037 4084 5043 4116
rect 5053 4104 5059 4136
rect 5149 4124 5155 4176
rect 5005 4077 5020 4083
rect 5012 3877 5027 3883
rect 4989 3864 4995 3876
rect 4781 3784 4787 3836
rect 4925 3764 4931 3776
rect 4973 3764 4979 3836
rect 5005 3784 5011 3856
rect 5021 3784 5027 3877
rect 5037 3784 5043 4036
rect 5053 4004 5059 4096
rect 5069 4024 5075 4096
rect 5165 4044 5171 4136
rect 5245 4124 5251 4296
rect 5261 4263 5267 4276
rect 5261 4257 5276 4263
rect 5261 4164 5267 4257
rect 5261 4144 5267 4156
rect 5053 3904 5059 3916
rect 5133 3904 5139 4036
rect 5261 4023 5267 4136
rect 5293 4124 5299 4296
rect 5373 4184 5379 4416
rect 5389 4384 5395 4516
rect 5405 4504 5411 4536
rect 5389 4304 5395 4336
rect 5405 4304 5411 4496
rect 5421 4444 5427 4536
rect 5517 4444 5523 4536
rect 5389 4264 5395 4276
rect 5437 4144 5443 4336
rect 5469 4304 5475 4436
rect 5533 4384 5539 4456
rect 5485 4304 5491 4316
rect 5549 4304 5555 4556
rect 5469 4164 5475 4276
rect 5341 4104 5347 4136
rect 5373 4124 5379 4136
rect 5373 4104 5379 4116
rect 5421 4104 5427 4136
rect 5277 4044 5283 4096
rect 5309 4084 5315 4096
rect 5261 4017 5283 4023
rect 5245 3984 5251 3996
rect 5085 3864 5091 3896
rect 5101 3884 5107 3896
rect 5149 3884 5155 3916
rect 5181 3864 5187 3916
rect 5069 3784 5075 3856
rect 4861 3744 4867 3756
rect 4733 3697 4748 3703
rect 4749 3564 4755 3696
rect 4733 3504 4739 3536
rect 4765 3484 4771 3616
rect 4781 3524 4787 3656
rect 4797 3584 4803 3716
rect 4909 3704 4915 3756
rect 4973 3744 4979 3756
rect 5085 3744 5091 3856
rect 5117 3743 5123 3836
rect 5133 3824 5139 3856
rect 5213 3784 5219 3816
rect 5117 3737 5132 3743
rect 5021 3724 5027 3736
rect 4973 3704 4979 3716
rect 5053 3704 5059 3736
rect 5085 3724 5091 3736
rect 5229 3704 5235 3936
rect 5261 3864 5267 3876
rect 5245 3744 5251 3856
rect 5245 3724 5251 3736
rect 4824 3606 4830 3614
rect 4838 3606 4844 3614
rect 4852 3606 4858 3614
rect 4866 3606 4872 3614
rect 4925 3524 4931 3576
rect 4717 3463 4723 3476
rect 4797 3464 4803 3496
rect 5037 3484 5043 3536
rect 4708 3457 4723 3463
rect 4669 3304 4675 3356
rect 4701 3304 4707 3456
rect 4781 3424 4787 3436
rect 4893 3424 4899 3476
rect 4749 3324 4755 3336
rect 4564 3297 4579 3303
rect 4541 3184 4547 3256
rect 4557 3204 4563 3296
rect 4653 3244 4659 3296
rect 4573 3184 4579 3236
rect 4573 3124 4579 3156
rect 4589 3124 4595 3236
rect 4637 3204 4643 3236
rect 4669 3203 4675 3296
rect 4733 3284 4739 3316
rect 4845 3304 4851 3396
rect 4813 3244 4819 3276
rect 4829 3264 4835 3296
rect 4653 3197 4675 3203
rect 4637 3144 4643 3156
rect 4653 3124 4659 3197
rect 4493 3104 4499 3116
rect 4509 3044 4515 3076
rect 4557 3043 4563 3116
rect 4589 3064 4595 3116
rect 4605 3043 4611 3056
rect 4557 3037 4611 3043
rect 4461 2924 4467 2936
rect 4429 2917 4444 2923
rect 4429 2904 4435 2917
rect 4493 2904 4499 2956
rect 4525 2924 4531 2956
rect 4557 2904 4563 2976
rect 4653 2964 4659 2976
rect 4589 2924 4595 2956
rect 4397 2884 4403 2896
rect 4621 2843 4627 2916
rect 4669 2904 4675 3156
rect 4685 3144 4691 3196
rect 4701 3184 4707 3236
rect 4717 3144 4723 3236
rect 4824 3206 4830 3214
rect 4838 3206 4844 3214
rect 4852 3206 4858 3214
rect 4866 3206 4872 3214
rect 4749 3144 4755 3196
rect 4893 3184 4899 3316
rect 4909 3143 4915 3436
rect 4941 3364 4947 3476
rect 5069 3464 5075 3516
rect 5117 3504 5123 3636
rect 5229 3524 5235 3696
rect 5261 3684 5267 3856
rect 5277 3704 5283 4017
rect 5341 3984 5347 4036
rect 5309 3924 5315 3956
rect 5437 3944 5443 4136
rect 5469 4044 5475 4096
rect 5453 3924 5459 4036
rect 5293 3904 5299 3916
rect 5341 3904 5347 3916
rect 5421 3884 5427 3896
rect 5421 3844 5427 3876
rect 5469 3844 5475 3876
rect 5485 3864 5491 4296
rect 5501 4264 5507 4296
rect 5501 4144 5507 4156
rect 5517 4144 5523 4296
rect 5533 4244 5539 4296
rect 5533 4124 5539 4236
rect 5565 4104 5571 4576
rect 5789 4564 5795 4636
rect 5581 4404 5587 4516
rect 5661 4464 5667 4556
rect 5709 4524 5715 4536
rect 5837 4524 5843 4636
rect 5869 4584 5875 4676
rect 5917 4584 5923 4676
rect 5933 4564 5939 4636
rect 5949 4584 5955 4676
rect 5981 4664 5987 4696
rect 5997 4644 6003 4676
rect 6013 4584 6019 4636
rect 6029 4624 6035 4676
rect 6045 4644 6051 4696
rect 6109 4644 6115 4676
rect 6125 4624 6131 4696
rect 6141 4684 6147 4716
rect 6173 4684 6179 4716
rect 6173 4624 6179 4676
rect 6189 4564 6195 4636
rect 6029 4544 6035 4556
rect 6093 4544 6099 4556
rect 5869 4524 5875 4536
rect 5828 4517 5836 4523
rect 5885 4504 5891 4536
rect 5677 4324 5683 4376
rect 5661 4277 5676 4283
rect 5661 4184 5667 4277
rect 5693 4224 5699 4476
rect 5725 4424 5731 4496
rect 5773 4484 5779 4496
rect 5725 4243 5731 4316
rect 5789 4304 5795 4456
rect 5805 4364 5811 4436
rect 5837 4384 5843 4436
rect 5933 4424 5939 4536
rect 6045 4524 6051 4536
rect 6109 4524 6115 4536
rect 6077 4484 6083 4496
rect 6077 4464 6083 4476
rect 5741 4264 5747 4276
rect 5805 4264 5811 4316
rect 6013 4304 6019 4316
rect 6013 4284 6019 4296
rect 5805 4244 5811 4256
rect 5725 4237 5740 4243
rect 5741 4184 5747 4236
rect 5581 4124 5587 4136
rect 5604 4117 5619 4123
rect 5533 4024 5539 4036
rect 5565 3964 5571 4096
rect 5581 3984 5587 4116
rect 5613 3984 5619 4117
rect 5645 4104 5651 4116
rect 5629 4004 5635 4096
rect 5677 4084 5683 4096
rect 5693 4083 5699 4156
rect 5901 4144 5907 4256
rect 5933 4243 5939 4276
rect 5981 4264 5987 4276
rect 6045 4264 6051 4436
rect 6093 4384 6099 4416
rect 6077 4264 6083 4336
rect 5917 4237 5939 4243
rect 5684 4077 5699 4083
rect 5709 4064 5715 4136
rect 5757 4064 5763 4136
rect 5853 4084 5859 4136
rect 5917 4124 5923 4237
rect 5965 4124 5971 4236
rect 6013 4144 6019 4236
rect 6061 4184 6067 4236
rect 5981 4124 5987 4136
rect 5933 4104 5939 4116
rect 5965 4084 5971 4116
rect 6061 4104 6067 4156
rect 5613 3944 5619 3976
rect 5581 3924 5587 3936
rect 5517 3904 5523 3916
rect 5533 3904 5539 3916
rect 5533 3864 5539 3876
rect 5549 3804 5555 3896
rect 5629 3884 5635 3996
rect 5709 3884 5715 3976
rect 5748 3937 5763 3943
rect 5741 3924 5747 3936
rect 5757 3864 5763 3937
rect 5389 3744 5395 3796
rect 5581 3764 5587 3796
rect 5277 3684 5283 3696
rect 5437 3684 5443 3716
rect 5517 3704 5523 3736
rect 5533 3704 5539 3716
rect 5460 3697 5475 3703
rect 5197 3484 5203 3516
rect 5341 3504 5347 3656
rect 4957 3304 4963 3416
rect 5005 3403 5011 3436
rect 5117 3404 5123 3436
rect 5229 3424 5235 3436
rect 5005 3397 5027 3403
rect 5021 3364 5027 3397
rect 5005 3324 5011 3336
rect 5021 3304 5027 3356
rect 5069 3324 5075 3336
rect 4925 3244 4931 3276
rect 4893 3137 4915 3143
rect 4701 3104 4707 3136
rect 4797 3124 4803 3136
rect 4717 3044 4723 3116
rect 4781 3084 4787 3116
rect 4813 3104 4819 3136
rect 4749 2924 4755 2936
rect 4692 2917 4723 2923
rect 4621 2837 4636 2843
rect 4525 2824 4531 2836
rect 4701 2824 4707 2876
rect 4717 2863 4723 2917
rect 4733 2904 4739 2916
rect 4797 2904 4803 2976
rect 4813 2924 4819 2936
rect 4893 2904 4899 3137
rect 4909 3044 4915 3116
rect 4925 3104 4931 3136
rect 4941 3124 4947 3136
rect 4989 3104 4995 3256
rect 5053 3184 5059 3276
rect 5069 3264 5075 3276
rect 5117 3184 5123 3396
rect 5133 3283 5139 3416
rect 5181 3384 5187 3396
rect 5309 3364 5315 3496
rect 5325 3464 5331 3496
rect 5357 3484 5363 3636
rect 5405 3584 5411 3676
rect 5421 3644 5427 3676
rect 5437 3584 5443 3636
rect 5469 3524 5475 3697
rect 5485 3644 5491 3676
rect 5501 3664 5507 3696
rect 5549 3664 5555 3736
rect 5629 3684 5635 3716
rect 5645 3704 5651 3796
rect 5677 3724 5683 3736
rect 5661 3684 5667 3696
rect 5613 3664 5619 3676
rect 5517 3584 5523 3656
rect 5645 3584 5651 3636
rect 5581 3544 5587 3556
rect 5389 3484 5395 3516
rect 5469 3443 5475 3516
rect 5565 3504 5571 3516
rect 5485 3444 5491 3496
rect 5533 3464 5539 3496
rect 5453 3437 5475 3443
rect 5149 3304 5155 3316
rect 5245 3304 5251 3356
rect 5293 3304 5299 3316
rect 5309 3304 5315 3356
rect 5325 3304 5331 3316
rect 5133 3277 5155 3283
rect 5133 3184 5139 3256
rect 5021 3124 5027 3136
rect 5037 3124 5043 3176
rect 5069 3144 5075 3156
rect 5117 3144 5123 3156
rect 5149 3124 5155 3277
rect 5165 3264 5171 3276
rect 5213 3264 5219 3276
rect 5229 3264 5235 3296
rect 4973 3044 4979 3076
rect 5149 3064 5155 3116
rect 5181 3084 5187 3156
rect 5213 3103 5219 3256
rect 5213 3097 5228 3103
rect 5245 3084 5251 3296
rect 5341 3284 5347 3336
rect 5357 3124 5363 3436
rect 5421 3384 5427 3436
rect 5437 3324 5443 3436
rect 5453 3344 5459 3437
rect 5469 3344 5475 3416
rect 5533 3364 5539 3456
rect 5549 3344 5555 3456
rect 5581 3404 5587 3496
rect 5597 3384 5603 3536
rect 5693 3524 5699 3756
rect 5789 3744 5795 4016
rect 5821 3884 5827 3896
rect 5821 3864 5827 3876
rect 5757 3704 5763 3716
rect 5821 3684 5827 3696
rect 5837 3663 5843 4056
rect 5853 3924 5859 3936
rect 5885 3884 5891 4036
rect 5821 3657 5843 3663
rect 5709 3564 5715 3636
rect 5613 3364 5619 3516
rect 5693 3484 5699 3516
rect 5757 3464 5763 3636
rect 5629 3384 5635 3456
rect 5597 3344 5603 3356
rect 5469 3324 5475 3336
rect 5421 3304 5427 3316
rect 5613 3304 5619 3356
rect 5645 3344 5651 3376
rect 5661 3324 5667 3396
rect 5725 3384 5731 3436
rect 5773 3424 5779 3496
rect 5789 3384 5795 3596
rect 5773 3344 5779 3376
rect 5780 3337 5795 3343
rect 5789 3304 5795 3337
rect 5501 3264 5507 3296
rect 5565 3144 5571 3156
rect 5581 3144 5587 3236
rect 5629 3144 5635 3156
rect 5581 3124 5587 3136
rect 5524 3117 5539 3123
rect 5389 3084 5395 3096
rect 5229 3064 5235 3076
rect 4989 3004 4995 3036
rect 5021 3004 5027 3036
rect 5021 2944 5027 2956
rect 5069 2944 5075 3056
rect 5405 3044 5411 3096
rect 5533 3064 5539 3117
rect 5357 2984 5363 3036
rect 5405 2964 5411 2996
rect 5453 2984 5459 3056
rect 5597 3024 5603 3116
rect 5501 2984 5507 2996
rect 5565 2964 5571 2996
rect 4957 2937 4972 2943
rect 4925 2924 4931 2936
rect 4941 2884 4947 2916
rect 4765 2864 4771 2876
rect 4829 2864 4835 2876
rect 4717 2857 4748 2863
rect 4141 2724 4147 2816
rect 4205 2684 4211 2696
rect 4269 2684 4275 2716
rect 4301 2684 4307 2716
rect 4461 2697 4476 2703
rect 4157 2664 4163 2676
rect 4141 2624 4147 2636
rect 4141 2564 4147 2616
rect 4109 2544 4115 2556
rect 4173 2544 4179 2616
rect 4237 2564 4243 2616
rect 4084 2537 4099 2543
rect 4189 2537 4243 2543
rect 4189 2524 4195 2537
rect 4237 2524 4243 2537
rect 4285 2524 4291 2616
rect 4333 2564 4339 2696
rect 4349 2564 4355 2656
rect 4397 2544 4403 2636
rect 4429 2624 4435 2676
rect 4429 2543 4435 2556
rect 4429 2537 4444 2543
rect 4301 2524 4307 2536
rect 4397 2484 4403 2516
rect 4445 2484 4451 2516
rect 3917 2384 3923 2436
rect 3661 1904 3667 1936
rect 3693 1924 3699 2096
rect 3885 1944 3891 2116
rect 3949 2104 3955 2256
rect 3965 2184 3971 2256
rect 3949 1984 3955 2096
rect 3981 2004 3987 2436
rect 4189 2384 4195 2456
rect 4253 2384 4259 2476
rect 4461 2464 4467 2697
rect 4509 2684 4515 2696
rect 4493 2584 4499 2656
rect 4093 2324 4099 2376
rect 4141 2304 4147 2336
rect 4253 2304 4259 2316
rect 3709 1884 3715 1936
rect 3885 1904 3891 1936
rect 3757 1884 3763 1896
rect 3965 1864 3971 1916
rect 3997 1904 4003 2296
rect 4029 2244 4035 2276
rect 4045 2264 4051 2296
rect 4237 2264 4243 2276
rect 4253 2264 4259 2296
rect 4029 2144 4035 2236
rect 4045 2124 4051 2236
rect 4221 2224 4227 2256
rect 4269 2184 4275 2436
rect 4493 2384 4499 2476
rect 4285 2224 4291 2316
rect 4301 2304 4307 2376
rect 4509 2344 4515 2556
rect 4525 2544 4531 2676
rect 4573 2664 4579 2676
rect 4621 2624 4627 2696
rect 4653 2644 4659 2656
rect 4580 2517 4595 2523
rect 4525 2464 4531 2516
rect 4589 2503 4595 2517
rect 4589 2497 4604 2503
rect 4333 2304 4339 2316
rect 4237 2157 4252 2163
rect 4029 2104 4035 2116
rect 4205 2104 4211 2156
rect 4237 2104 4243 2157
rect 4301 2144 4307 2296
rect 4317 2284 4323 2296
rect 4349 2264 4355 2316
rect 4413 2304 4419 2336
rect 4365 2264 4371 2296
rect 4461 2264 4467 2276
rect 4381 2156 4387 2236
rect 4509 2164 4515 2336
rect 4557 2324 4563 2496
rect 4621 2344 4627 2616
rect 4701 2524 4707 2536
rect 4717 2524 4723 2576
rect 4637 2504 4643 2516
rect 4653 2484 4659 2496
rect 4669 2484 4675 2516
rect 4637 2324 4643 2336
rect 4701 2324 4707 2516
rect 4717 2384 4723 2436
rect 4733 2424 4739 2836
rect 4824 2806 4830 2814
rect 4838 2806 4844 2814
rect 4852 2806 4858 2814
rect 4866 2806 4872 2814
rect 4957 2784 4963 2937
rect 5021 2904 5027 2916
rect 5245 2904 5251 2956
rect 5277 2924 5283 2936
rect 5261 2904 5267 2916
rect 5197 2884 5203 2896
rect 5229 2884 5235 2896
rect 5293 2884 5299 2916
rect 5309 2904 5315 2916
rect 5341 2884 5347 2936
rect 5405 2903 5411 2956
rect 5485 2944 5491 2956
rect 5517 2924 5523 2956
rect 5549 2924 5555 2956
rect 5469 2904 5475 2916
rect 5396 2897 5411 2903
rect 5565 2884 5571 2916
rect 5597 2884 5603 2936
rect 5613 2924 5619 2956
rect 4781 2664 4787 2696
rect 4909 2664 4915 2756
rect 5453 2724 5459 2736
rect 5325 2702 5331 2716
rect 4749 2524 4755 2556
rect 4765 2544 4771 2556
rect 4781 2464 4787 2516
rect 4525 2264 4531 2296
rect 4637 2284 4643 2296
rect 4669 2244 4675 2276
rect 4445 2144 4451 2156
rect 4221 1943 4227 2036
rect 4253 1984 4259 2136
rect 4445 2104 4451 2136
rect 4397 1984 4403 2056
rect 4205 1937 4227 1943
rect 4205 1924 4211 1937
rect 4333 1904 4339 1916
rect 4013 1877 4028 1883
rect 3549 1764 3555 1776
rect 3357 1744 3363 1756
rect 3293 1704 3299 1736
rect 3517 1724 3523 1756
rect 3581 1744 3587 1856
rect 4013 1744 4019 1877
rect 4029 1844 4035 1856
rect 4077 1824 4083 1836
rect 3389 1704 3395 1716
rect 2989 1697 3011 1703
rect 2733 1477 2748 1483
rect 2701 1424 2707 1476
rect 2749 1464 2755 1476
rect 2701 1383 2707 1416
rect 2685 1377 2707 1383
rect 2669 1344 2675 1356
rect 2589 1324 2595 1336
rect 2685 1324 2691 1377
rect 2717 1363 2723 1436
rect 2708 1357 2723 1363
rect 2605 1317 2620 1323
rect 2605 1304 2611 1317
rect 2557 1104 2563 1116
rect 2573 1084 2579 1136
rect 2653 1104 2659 1316
rect 2701 1144 2707 1356
rect 2749 1324 2755 1456
rect 2765 1384 2771 1436
rect 2781 1364 2787 1476
rect 2797 1464 2803 1496
rect 2877 1464 2883 1536
rect 2893 1524 2899 1596
rect 2989 1584 2995 1697
rect 3229 1684 3235 1696
rect 3037 1583 3043 1636
rect 3037 1577 3059 1583
rect 3053 1502 3059 1577
rect 3117 1564 3123 1656
rect 3293 1584 3299 1656
rect 3549 1584 3555 1696
rect 3581 1564 3587 1736
rect 3885 1684 3891 1736
rect 3997 1724 4003 1736
rect 4109 1724 4115 1736
rect 4125 1704 4131 1836
rect 4141 1803 4147 1876
rect 4173 1864 4179 1896
rect 4205 1884 4211 1896
rect 4141 1797 4156 1803
rect 4157 1744 4163 1796
rect 4205 1744 4211 1796
rect 4221 1764 4227 1836
rect 3117 1504 3123 1556
rect 3677 1524 3683 1536
rect 3725 1524 3731 1536
rect 3773 1524 3779 1576
rect 3901 1524 3907 1576
rect 3933 1544 3939 1636
rect 4045 1584 4051 1636
rect 2813 1444 2819 1456
rect 2829 1384 2835 1436
rect 2877 1384 2883 1456
rect 2797 1324 2803 1376
rect 2653 1064 2659 1096
rect 1853 664 1859 736
rect 1901 704 1907 756
rect 1917 744 1923 836
rect 1933 784 1939 876
rect 1917 684 1923 716
rect 1933 704 1939 756
rect 1949 744 1955 876
rect 1981 844 1987 876
rect 1981 744 1987 836
rect 2013 744 2019 756
rect 1949 724 1955 736
rect 1981 724 1987 736
rect 1997 684 2003 696
rect 2109 684 2115 836
rect 2125 764 2131 836
rect 2205 684 2211 816
rect 2221 744 2227 856
rect 2253 743 2259 836
rect 2253 737 2275 743
rect 2221 684 2227 736
rect 2253 684 2259 716
rect 2269 704 2275 737
rect 1869 544 1875 656
rect 2093 644 2099 676
rect 2013 544 2019 636
rect 2045 624 2051 636
rect 2045 584 2051 596
rect 2109 564 2115 676
rect 2140 664 2148 670
rect 2285 664 2291 956
rect 2301 944 2307 976
rect 2349 944 2355 956
rect 2365 944 2371 956
rect 2301 924 2307 936
rect 2365 924 2371 936
rect 2365 683 2371 716
rect 2397 704 2403 1036
rect 2445 944 2451 956
rect 2349 677 2371 683
rect 2301 644 2307 656
rect 2349 644 2355 677
rect 2429 683 2435 936
rect 2445 784 2451 936
rect 2461 844 2467 1036
rect 2493 904 2499 916
rect 2477 784 2483 896
rect 2509 864 2515 1036
rect 2509 764 2515 836
rect 2420 677 2435 683
rect 2397 644 2403 676
rect 2429 664 2435 677
rect 2141 584 2147 636
rect 2125 544 2131 556
rect 2109 504 2115 536
rect 1901 484 1907 496
rect 1677 477 1692 483
rect 2237 444 2243 636
rect 2301 504 2307 516
rect 2317 504 2323 616
rect 2445 564 2451 676
rect 2509 664 2515 736
rect 2525 704 2531 916
rect 2541 904 2547 936
rect 2557 924 2563 936
rect 2605 924 2611 936
rect 2573 724 2579 836
rect 2461 524 2467 536
rect 2429 484 2435 496
rect 1597 404 1603 436
rect 1629 424 1635 436
rect 1581 304 1587 336
rect 1629 324 1635 356
rect 1709 344 1715 436
rect 1768 406 1774 414
rect 1782 406 1788 414
rect 1796 406 1802 414
rect 1810 406 1816 414
rect 1741 324 1747 396
rect 1837 344 1843 436
rect 1869 344 1875 356
rect 1844 337 1852 343
rect 1629 304 1635 316
rect 1645 284 1651 316
rect 1693 304 1699 316
rect 1709 304 1715 316
rect 1725 284 1731 316
rect 1741 304 1747 316
rect 1869 304 1875 316
rect 1901 284 1907 296
rect 1997 284 2003 416
rect 2013 324 2019 436
rect 2013 304 2019 316
rect 2045 284 2051 396
rect 2061 304 2067 356
rect 2077 284 2083 336
rect 1156 237 1171 243
rect 1197 144 1203 256
rect 1213 224 1219 236
rect 1261 204 1267 236
rect 1277 183 1283 196
rect 1268 177 1283 183
rect 1293 164 1299 236
rect 964 117 988 123
rect 701 97 739 103
rect 701 64 707 97
rect 733 84 739 97
rect 749 77 780 83
rect 717 64 723 76
rect 749 63 755 77
rect 797 64 803 96
rect 829 83 835 116
rect 1005 103 1011 136
rect 980 97 1011 103
rect 1076 97 1100 103
rect 820 77 835 83
rect 916 77 940 83
rect 957 64 963 76
rect 733 57 755 63
rect 653 43 659 56
rect 733 43 739 57
rect 973 44 979 76
rect 1309 64 1315 236
rect 1325 224 1331 256
rect 1405 164 1411 216
rect 1437 184 1443 236
rect 1405 124 1411 156
rect 1341 64 1347 98
rect 1485 103 1491 116
rect 1549 104 1555 236
rect 1613 164 1619 176
rect 1476 97 1491 103
rect 1565 84 1571 116
rect 1581 104 1587 136
rect 1661 123 1667 136
rect 1709 124 1715 256
rect 2157 244 2163 436
rect 2205 264 2211 396
rect 2285 324 2291 436
rect 2365 324 2371 336
rect 2221 244 2227 256
rect 1661 117 1699 123
rect 1645 64 1651 116
rect 1693 104 1699 117
rect 1805 104 1811 176
rect 1933 164 1939 236
rect 2013 164 2019 236
rect 1821 104 1827 116
rect 1901 104 1907 116
rect 1917 104 1923 116
rect 1677 64 1683 96
rect 1933 84 1939 116
rect 1949 104 1955 136
rect 1965 83 1971 156
rect 2029 144 2035 196
rect 2109 124 2115 156
rect 2157 144 2163 216
rect 2253 144 2259 236
rect 2045 104 2051 116
rect 2269 104 2275 316
rect 2285 284 2291 316
rect 2381 304 2387 436
rect 2317 284 2323 296
rect 2429 284 2435 436
rect 2493 404 2499 636
rect 2509 524 2515 596
rect 2525 544 2531 696
rect 2541 504 2547 716
rect 2605 704 2611 836
rect 2621 824 2627 1036
rect 2669 1004 2675 1116
rect 2701 1044 2707 1076
rect 2717 1044 2723 1076
rect 2765 1044 2771 1116
rect 2813 1084 2819 1316
rect 2829 1304 2835 1356
rect 2893 1344 2899 1496
rect 2909 1343 2915 1456
rect 2925 1404 2931 1476
rect 2941 1424 2947 1496
rect 2973 1464 2979 1476
rect 2973 1424 2979 1456
rect 2941 1344 2947 1416
rect 2909 1337 2924 1343
rect 2973 1304 2979 1376
rect 2989 1364 2995 1376
rect 3069 1344 3075 1376
rect 3117 1364 3123 1376
rect 3165 1364 3171 1496
rect 3261 1484 3267 1496
rect 3181 1424 3187 1436
rect 3197 1384 3203 1436
rect 3213 1324 3219 1416
rect 3229 1404 3235 1476
rect 3053 1304 3059 1316
rect 3229 1304 3235 1396
rect 3261 1384 3267 1476
rect 3277 1444 3283 1496
rect 3325 1464 3331 1496
rect 3453 1484 3459 1496
rect 3501 1484 3507 1496
rect 3693 1484 3699 1496
rect 3741 1484 3747 1496
rect 3853 1484 3859 1496
rect 3949 1484 3955 1556
rect 4061 1484 4067 1576
rect 4141 1524 4147 1636
rect 4077 1484 4083 1516
rect 4109 1504 4115 1516
rect 4173 1504 4179 1636
rect 4221 1564 4227 1756
rect 4237 1744 4243 1816
rect 4333 1744 4339 1796
rect 4349 1683 4355 1736
rect 4461 1704 4467 1894
rect 4477 1744 4483 1976
rect 4493 1764 4499 2076
rect 4509 1904 4515 1916
rect 4509 1784 4515 1856
rect 4525 1784 4531 2196
rect 4541 2144 4547 2176
rect 4701 2144 4707 2276
rect 4781 2144 4787 2356
rect 4797 2344 4803 2516
rect 4877 2504 4883 2616
rect 4909 2504 4915 2636
rect 4941 2604 4947 2696
rect 5197 2684 5203 2696
rect 5101 2664 5107 2676
rect 4989 2644 4995 2656
rect 4925 2484 4931 2536
rect 4973 2524 4979 2636
rect 5037 2584 5043 2656
rect 5069 2504 5075 2656
rect 5085 2484 5091 2496
rect 4909 2477 4924 2483
rect 4824 2406 4830 2414
rect 4838 2406 4844 2414
rect 4852 2406 4858 2414
rect 4866 2406 4872 2414
rect 4877 2284 4883 2296
rect 4573 1924 4579 2136
rect 4605 2126 4611 2136
rect 4669 2124 4675 2136
rect 4797 2104 4803 2176
rect 4909 2144 4915 2477
rect 4973 2302 4979 2336
rect 5005 2284 5011 2436
rect 5037 2304 5043 2416
rect 5085 2383 5091 2476
rect 5101 2424 5107 2656
rect 5165 2564 5171 2636
rect 5261 2584 5267 2636
rect 5197 2564 5203 2576
rect 5277 2564 5283 2576
rect 5165 2544 5171 2556
rect 5085 2377 5100 2383
rect 5117 2364 5123 2536
rect 5197 2524 5203 2556
rect 5309 2504 5315 2556
rect 5389 2544 5395 2696
rect 5485 2544 5491 2676
rect 5517 2524 5523 2536
rect 5565 2384 5571 2856
rect 5629 2704 5635 3036
rect 5661 2964 5667 3196
rect 5661 2904 5667 2956
rect 5645 2784 5651 2876
rect 5677 2864 5683 3296
rect 5741 3164 5747 3236
rect 5716 3137 5724 3143
rect 5693 3104 5699 3136
rect 5693 3084 5699 3096
rect 5709 3064 5715 3116
rect 5725 3104 5731 3136
rect 5789 3124 5795 3156
rect 5789 3084 5795 3096
rect 5693 2824 5699 3036
rect 5805 2964 5811 3416
rect 5821 3304 5827 3657
rect 5853 3604 5859 3676
rect 5869 3664 5875 3716
rect 5853 3584 5859 3596
rect 5876 3537 5891 3543
rect 5837 3524 5843 3536
rect 5869 3524 5875 3536
rect 5837 3504 5843 3516
rect 5885 3464 5891 3537
rect 5901 3463 5907 4076
rect 5933 3864 5939 3916
rect 5917 3724 5923 3736
rect 5917 3604 5923 3676
rect 5933 3664 5939 3716
rect 5965 3704 5971 3756
rect 5917 3544 5923 3576
rect 5917 3504 5923 3536
rect 5933 3504 5939 3516
rect 5917 3484 5923 3496
rect 5949 3484 5955 3676
rect 5965 3664 5971 3696
rect 5981 3684 5987 3896
rect 5997 3784 6003 3916
rect 6029 3904 6035 3956
rect 6045 3744 6051 3976
rect 6077 3904 6083 4156
rect 6093 4123 6099 4176
rect 6125 4164 6131 4556
rect 6205 4544 6211 4716
rect 6221 4704 6227 4736
rect 6253 4704 6259 4716
rect 6285 4664 6291 4676
rect 6349 4623 6355 4694
rect 6477 4624 6483 4636
rect 6333 4617 6355 4623
rect 6301 4524 6307 4536
rect 6141 4444 6147 4496
rect 6173 4464 6179 4516
rect 6173 4284 6179 4456
rect 6189 4304 6195 4336
rect 6205 4284 6211 4516
rect 6253 4504 6259 4516
rect 6269 4484 6275 4496
rect 6285 4384 6291 4496
rect 6317 4484 6323 4496
rect 6237 4324 6243 4356
rect 6285 4344 6291 4376
rect 6301 4323 6307 4436
rect 6317 4324 6323 4336
rect 6301 4317 6316 4323
rect 6301 4284 6307 4296
rect 6317 4284 6323 4316
rect 6205 4264 6211 4276
rect 6333 4263 6339 4617
rect 6381 4524 6387 4536
rect 6365 4484 6371 4496
rect 6381 4344 6387 4436
rect 6397 4424 6403 4496
rect 6445 4464 6451 4476
rect 6429 4424 6435 4436
rect 6397 4384 6403 4396
rect 6429 4383 6435 4416
rect 6429 4377 6451 4383
rect 6381 4324 6387 4336
rect 6397 4304 6403 4356
rect 6349 4284 6355 4296
rect 6333 4257 6355 4263
rect 6157 4183 6163 4236
rect 6141 4177 6163 4183
rect 6093 4117 6108 4123
rect 6125 4104 6131 4136
rect 6141 3963 6147 4177
rect 6157 4144 6163 4156
rect 6164 4137 6179 4143
rect 6173 4104 6179 4137
rect 6189 4104 6195 4116
rect 6205 4084 6211 4176
rect 6221 4144 6227 4236
rect 6253 4224 6259 4256
rect 6237 4104 6243 4136
rect 6157 4024 6163 4036
rect 6125 3957 6147 3963
rect 6109 3904 6115 3956
rect 6077 3864 6083 3876
rect 6061 3744 6067 3836
rect 6093 3744 6099 3836
rect 6013 3677 6028 3683
rect 5965 3483 5971 3596
rect 5981 3503 5987 3636
rect 5997 3504 6003 3516
rect 5981 3497 5996 3503
rect 5965 3477 5980 3483
rect 5901 3457 5923 3463
rect 5837 3344 5843 3356
rect 5821 3144 5827 3216
rect 5853 3124 5859 3456
rect 5917 3324 5923 3457
rect 5949 3444 5955 3456
rect 5965 3323 5971 3436
rect 6013 3363 6019 3677
rect 6061 3677 6076 3683
rect 6029 3664 6035 3676
rect 6045 3604 6051 3676
rect 6061 3604 6067 3677
rect 6029 3504 6035 3536
rect 6045 3504 6051 3536
rect 6061 3524 6067 3556
rect 6077 3524 6083 3656
rect 6093 3624 6099 3636
rect 6109 3604 6115 3836
rect 6125 3704 6131 3957
rect 6141 3864 6147 3936
rect 6157 3924 6163 3956
rect 6237 3944 6243 4096
rect 6269 3944 6275 4236
rect 6285 4184 6291 4256
rect 6317 4124 6323 4216
rect 6333 4184 6339 4236
rect 6285 4064 6291 4096
rect 6317 4084 6323 4116
rect 6349 4083 6355 4257
rect 6365 4104 6371 4156
rect 6349 4077 6371 4083
rect 6253 3904 6259 3936
rect 6317 3904 6323 4036
rect 6333 4004 6339 4056
rect 6253 3884 6259 3896
rect 6269 3864 6275 3896
rect 6189 3824 6195 3856
rect 6141 3644 6147 3716
rect 6189 3677 6204 3683
rect 6157 3664 6163 3676
rect 6189 3664 6195 3677
rect 6221 3664 6227 3716
rect 6269 3703 6275 3796
rect 6285 3744 6291 3896
rect 6333 3884 6339 3996
rect 6349 3904 6355 4016
rect 6365 3883 6371 4077
rect 6381 4064 6387 4176
rect 6397 4164 6403 4296
rect 6413 4264 6419 4316
rect 6429 4184 6435 4316
rect 6445 4304 6451 4377
rect 6461 4363 6467 4396
rect 6477 4384 6483 4496
rect 6493 4464 6499 4476
rect 6509 4444 6515 4636
rect 6557 4544 6563 4696
rect 6525 4497 6540 4503
rect 6493 4364 6499 4436
rect 6461 4357 6483 4363
rect 6477 4323 6483 4357
rect 6509 4323 6515 4336
rect 6525 4324 6531 4497
rect 6541 4344 6547 4476
rect 6557 4424 6563 4516
rect 6461 4317 6483 4323
rect 6493 4317 6515 4323
rect 6461 4284 6467 4317
rect 6445 4184 6451 4276
rect 6445 4144 6451 4156
rect 6397 4104 6403 4116
rect 6413 4084 6419 4136
rect 6349 3877 6371 3883
rect 6285 3724 6291 3736
rect 6269 3697 6284 3703
rect 6093 3584 6099 3596
rect 6109 3544 6115 3556
rect 6093 3504 6099 3536
rect 6125 3504 6131 3616
rect 6189 3584 6195 3656
rect 6157 3544 6163 3576
rect 6173 3544 6179 3556
rect 6189 3544 6195 3576
rect 6221 3564 6227 3636
rect 6157 3504 6163 3536
rect 6045 3364 6051 3476
rect 6109 3364 6115 3456
rect 6013 3357 6028 3363
rect 6013 3324 6019 3357
rect 6045 3344 6051 3356
rect 5949 3317 5971 3323
rect 5949 3303 5955 3317
rect 5940 3297 5955 3303
rect 5885 3224 5891 3276
rect 5901 3184 5907 3296
rect 5821 3004 5827 3096
rect 5837 2984 5843 3076
rect 5853 3064 5859 3116
rect 5837 2964 5843 2976
rect 5853 2964 5859 2976
rect 5709 2924 5715 2936
rect 5757 2904 5763 2916
rect 5725 2884 5731 2896
rect 5149 2264 5155 2316
rect 5229 2304 5235 2356
rect 5165 2284 5171 2296
rect 5181 2263 5187 2276
rect 5213 2264 5219 2276
rect 5165 2257 5187 2263
rect 5149 2164 5155 2236
rect 5165 2204 5171 2257
rect 5181 2184 5187 2236
rect 5341 2204 5347 2316
rect 4829 2084 4835 2136
rect 5021 2104 5027 2136
rect 4589 1984 4595 1996
rect 4637 1904 4643 1936
rect 4653 1884 4659 1916
rect 4685 1864 4691 1896
rect 4605 1804 4611 1836
rect 4493 1744 4499 1756
rect 4349 1677 4371 1683
rect 3373 1444 3379 1476
rect 3405 1444 3411 1476
rect 3304 1406 3310 1414
rect 3318 1406 3324 1414
rect 3332 1406 3338 1414
rect 3346 1406 3352 1414
rect 3389 1404 3395 1436
rect 3245 1304 3251 1376
rect 3293 1344 3299 1376
rect 3405 1344 3411 1376
rect 3421 1324 3427 1456
rect 3453 1364 3459 1476
rect 3485 1304 3491 1456
rect 3645 1424 3651 1476
rect 3837 1464 3843 1476
rect 3517 1364 3523 1396
rect 3725 1384 3731 1436
rect 3613 1324 3619 1336
rect 3629 1324 3635 1356
rect 3645 1344 3651 1376
rect 3661 1324 3667 1336
rect 3565 1304 3571 1316
rect 2845 1284 2851 1296
rect 3021 1264 3027 1296
rect 2845 1124 2851 1156
rect 2877 1124 2883 1236
rect 2941 1084 2947 1116
rect 2957 1104 2963 1116
rect 3005 1084 3011 1236
rect 3101 1123 3107 1236
rect 3213 1184 3219 1236
rect 3101 1117 3116 1123
rect 3085 1084 3091 1096
rect 3117 1084 3123 1096
rect 3229 1084 3235 1256
rect 3277 1144 3283 1236
rect 3469 1124 3475 1156
rect 3005 1064 3011 1076
rect 2685 983 2691 1036
rect 2733 984 2739 1036
rect 2669 977 2691 983
rect 2637 964 2643 976
rect 2669 924 2675 977
rect 2653 704 2659 736
rect 2669 704 2675 836
rect 2685 744 2691 956
rect 2781 944 2787 1036
rect 2813 904 2819 936
rect 2829 924 2835 1056
rect 2733 724 2739 776
rect 2749 724 2755 876
rect 2573 624 2579 636
rect 2605 623 2611 676
rect 2765 664 2771 736
rect 2781 684 2787 776
rect 2797 744 2803 836
rect 2861 644 2867 1036
rect 2893 984 2899 1056
rect 2925 944 2931 976
rect 2957 944 2963 976
rect 3037 944 3043 1016
rect 3117 984 3123 1076
rect 3229 1064 3235 1076
rect 3069 944 3075 976
rect 3133 944 3139 1036
rect 3165 984 3171 1056
rect 3165 944 3171 976
rect 2893 904 2899 916
rect 3037 884 3043 936
rect 3053 924 3059 936
rect 2877 724 2883 836
rect 3005 764 3011 836
rect 2589 617 2611 623
rect 2557 464 2563 476
rect 2573 444 2579 476
rect 2589 424 2595 617
rect 2605 564 2611 596
rect 2621 584 2627 616
rect 2781 604 2787 636
rect 2973 624 2979 696
rect 3021 664 3027 736
rect 3117 724 3123 836
rect 3133 744 3139 936
rect 3213 924 3219 956
rect 3181 824 3187 916
rect 3261 884 3267 1036
rect 3197 844 3203 876
rect 3277 864 3283 1056
rect 3304 1006 3310 1014
rect 3318 1006 3324 1014
rect 3332 1006 3338 1014
rect 3346 1006 3352 1014
rect 3373 984 3379 1056
rect 3389 1004 3395 1116
rect 3437 1084 3443 1116
rect 3421 1044 3427 1076
rect 3421 964 3427 996
rect 3357 884 3363 956
rect 3437 944 3443 1076
rect 3373 924 3379 936
rect 3453 903 3459 1036
rect 3469 964 3475 1116
rect 3485 1084 3491 1176
rect 3549 1144 3555 1176
rect 3581 1124 3587 1136
rect 3501 963 3507 1036
rect 3524 997 3539 1003
rect 3501 957 3516 963
rect 3469 924 3475 936
rect 3501 904 3507 957
rect 3533 904 3539 997
rect 3565 944 3571 1096
rect 3597 1004 3603 1316
rect 3613 1284 3619 1316
rect 3709 1304 3715 1316
rect 3693 1264 3699 1296
rect 3629 1124 3635 1176
rect 3741 1084 3747 1396
rect 3837 1344 3843 1436
rect 3869 1424 3875 1476
rect 3965 1444 3971 1476
rect 3901 1404 3907 1436
rect 4141 1403 4147 1476
rect 4189 1464 4195 1536
rect 4157 1423 4163 1436
rect 4205 1423 4211 1456
rect 4157 1417 4211 1423
rect 4141 1397 4163 1403
rect 4013 1343 4019 1396
rect 4061 1344 4067 1376
rect 4093 1344 4099 1356
rect 4013 1337 4035 1343
rect 3821 1304 3827 1316
rect 3837 1304 3843 1316
rect 3853 1297 3900 1303
rect 3853 1283 3859 1297
rect 3997 1284 4003 1336
rect 4029 1323 4035 1337
rect 4109 1324 4115 1396
rect 4157 1344 4163 1397
rect 4221 1364 4227 1556
rect 4269 1464 4275 1516
rect 4237 1363 4243 1436
rect 4253 1384 4259 1396
rect 4285 1383 4291 1636
rect 4333 1484 4339 1496
rect 4349 1464 4355 1496
rect 4365 1484 4371 1677
rect 4461 1584 4467 1636
rect 4493 1584 4499 1736
rect 4525 1704 4531 1776
rect 4605 1744 4611 1776
rect 4637 1664 4643 1816
rect 4669 1703 4675 1736
rect 4685 1704 4691 1756
rect 4701 1704 4707 2036
rect 4765 1924 4771 2036
rect 4824 2006 4830 2014
rect 4838 2006 4844 2014
rect 4852 2006 4858 2014
rect 4866 2006 4872 2014
rect 4893 1964 4899 2036
rect 4941 1924 4947 1936
rect 4765 1884 4771 1916
rect 4893 1904 4899 1916
rect 4957 1904 4963 1916
rect 4989 1904 4995 1956
rect 4877 1884 4883 1896
rect 4925 1864 4931 1896
rect 4973 1864 4979 1896
rect 4989 1884 4995 1896
rect 4733 1804 4739 1856
rect 4813 1764 4819 1836
rect 4893 1804 4899 1856
rect 4893 1764 4899 1796
rect 4660 1697 4675 1703
rect 4701 1684 4707 1696
rect 4781 1684 4787 1736
rect 4813 1704 4819 1756
rect 4909 1744 4915 1856
rect 5005 1744 5011 1856
rect 5021 1764 5027 1896
rect 5037 1684 5043 2036
rect 5053 1924 5059 2076
rect 5085 2044 5091 2116
rect 5133 2104 5139 2136
rect 5181 2123 5187 2176
rect 5229 2164 5235 2176
rect 5373 2164 5379 2196
rect 5389 2184 5395 2256
rect 5213 2144 5219 2156
rect 5309 2144 5315 2156
rect 5341 2144 5347 2156
rect 5172 2117 5187 2123
rect 5261 2104 5267 2116
rect 5069 1924 5075 2016
rect 5101 1884 5107 2056
rect 5165 1904 5171 2036
rect 5309 1984 5315 2136
rect 5373 2104 5379 2156
rect 5389 2124 5395 2176
rect 5421 2164 5427 2356
rect 5517 2324 5523 2336
rect 5421 2144 5427 2156
rect 5453 2144 5459 2276
rect 5453 2124 5459 2136
rect 5485 2104 5491 2276
rect 5501 2144 5507 2156
rect 5517 2124 5523 2236
rect 5117 1864 5123 1876
rect 5149 1724 5155 1776
rect 5197 1724 5203 1776
rect 5213 1764 5219 1936
rect 5325 1904 5331 2036
rect 5341 1884 5347 1896
rect 5389 1864 5395 2016
rect 5405 1884 5411 1896
rect 5437 1884 5443 2096
rect 5533 2044 5539 2296
rect 5581 2284 5587 2516
rect 5709 2484 5715 2518
rect 5581 2224 5587 2276
rect 5597 2144 5603 2356
rect 5741 2284 5747 2676
rect 5773 2364 5779 2956
rect 5869 2944 5875 3096
rect 5885 3044 5891 3136
rect 5917 3104 5923 3156
rect 5933 3084 5939 3096
rect 5901 2984 5907 3016
rect 5917 2984 5923 3076
rect 5949 3024 5955 3297
rect 5965 3084 5971 3096
rect 5981 3084 5987 3196
rect 6029 3184 6035 3276
rect 5949 2984 5955 2996
rect 5789 2904 5795 2936
rect 5885 2924 5891 2976
rect 5965 2944 5971 2956
rect 5885 2784 5891 2896
rect 5901 2884 5907 2916
rect 5949 2702 5955 2736
rect 5853 2583 5859 2696
rect 5844 2577 5859 2583
rect 5949 2544 5955 2656
rect 5869 2344 5875 2536
rect 5949 2303 5955 2316
rect 5949 2297 5971 2303
rect 5709 2144 5715 2216
rect 5629 2124 5635 2136
rect 5661 2124 5667 2136
rect 5549 2084 5555 2116
rect 5581 2104 5587 2116
rect 5629 2104 5635 2116
rect 5453 1944 5459 2036
rect 5517 2024 5523 2036
rect 5469 1904 5475 1976
rect 5501 1924 5507 1976
rect 5517 1924 5523 1936
rect 5613 1924 5619 2036
rect 5661 1944 5667 2116
rect 5693 1924 5699 2036
rect 5549 1904 5555 1916
rect 5757 1884 5763 1936
rect 5549 1877 5564 1883
rect 5437 1864 5443 1876
rect 5229 1844 5235 1856
rect 5261 1844 5267 1856
rect 5261 1784 5267 1836
rect 5277 1763 5283 1836
rect 5405 1764 5411 1836
rect 5261 1757 5283 1763
rect 5213 1744 5219 1756
rect 5261 1724 5267 1757
rect 5501 1763 5507 1836
rect 5501 1757 5523 1763
rect 5293 1744 5299 1756
rect 5357 1740 5363 1756
rect 5517 1744 5523 1757
rect 5325 1704 5331 1736
rect 5501 1724 5507 1736
rect 5172 1697 5187 1703
rect 5085 1664 5091 1696
rect 4509 1584 4515 1596
rect 4461 1564 4467 1576
rect 4397 1544 4403 1556
rect 4525 1544 4531 1636
rect 4541 1584 4547 1596
rect 4557 1544 4563 1616
rect 4381 1464 4387 1536
rect 4461 1524 4467 1536
rect 4573 1524 4579 1636
rect 4493 1504 4499 1516
rect 4509 1504 4515 1516
rect 4525 1504 4531 1516
rect 4589 1504 4595 1516
rect 4605 1503 4611 1616
rect 4621 1544 4627 1636
rect 4717 1624 4723 1636
rect 4621 1524 4627 1536
rect 4605 1497 4620 1503
rect 4269 1377 4291 1383
rect 4237 1357 4259 1363
rect 4029 1317 4044 1323
rect 3812 1277 3859 1283
rect 3773 1124 3779 1256
rect 3837 1064 3843 1076
rect 3565 924 3571 936
rect 3453 897 3475 903
rect 3101 717 3116 723
rect 3037 664 3043 716
rect 3053 624 3059 696
rect 3101 664 3107 717
rect 3197 704 3203 736
rect 3229 724 3235 736
rect 3181 684 3187 696
rect 2669 524 2675 556
rect 2637 504 2643 516
rect 2653 504 2659 516
rect 2685 503 2691 536
rect 2733 524 2739 576
rect 2813 564 2819 576
rect 2749 544 2755 556
rect 2893 544 2899 556
rect 2685 497 2700 503
rect 2765 484 2771 496
rect 2477 324 2483 356
rect 2493 324 2499 396
rect 2493 304 2499 316
rect 2509 304 2515 376
rect 2525 284 2531 336
rect 2605 304 2611 316
rect 2621 297 2659 303
rect 2333 264 2339 276
rect 2557 264 2563 296
rect 2285 204 2291 236
rect 2333 224 2339 256
rect 2525 164 2531 216
rect 2589 184 2595 296
rect 2621 284 2627 297
rect 2621 264 2627 276
rect 2637 264 2643 276
rect 2653 263 2659 297
rect 2669 284 2675 356
rect 2685 284 2691 296
rect 2717 284 2723 336
rect 2733 304 2739 356
rect 2749 324 2755 336
rect 2781 304 2787 356
rect 2797 344 2803 476
rect 2813 464 2819 536
rect 2861 484 2867 516
rect 2893 504 2899 536
rect 2941 524 2947 576
rect 2957 544 2963 556
rect 2989 524 2995 596
rect 3037 504 3043 536
rect 3053 524 3059 596
rect 3117 564 3123 636
rect 3181 604 3187 636
rect 3229 564 3235 676
rect 3149 524 3155 556
rect 3245 484 3251 676
rect 3261 644 3267 696
rect 3277 684 3283 796
rect 3357 664 3363 736
rect 3373 684 3379 836
rect 3373 664 3379 676
rect 3304 606 3310 614
rect 3318 606 3324 614
rect 3332 606 3338 614
rect 3346 606 3352 614
rect 3373 584 3379 636
rect 3325 484 3331 516
rect 3341 504 3347 536
rect 3357 524 3363 556
rect 3389 484 3395 576
rect 3405 524 3411 636
rect 3421 544 3427 596
rect 3437 544 3443 836
rect 3469 724 3475 897
rect 3501 684 3507 896
rect 3517 684 3523 876
rect 3565 684 3571 816
rect 3581 704 3587 976
rect 3597 944 3603 976
rect 3629 964 3635 996
rect 3677 984 3683 1036
rect 3709 984 3715 1016
rect 3757 964 3763 1016
rect 3773 943 3779 1036
rect 3821 1024 3827 1056
rect 3789 944 3795 996
rect 3764 937 3779 943
rect 3821 904 3827 976
rect 3837 964 3843 976
rect 3853 944 3859 996
rect 3869 924 3875 1096
rect 3885 1084 3891 1236
rect 3933 1124 3939 1236
rect 3997 1104 4003 1276
rect 4013 1124 4019 1316
rect 4237 1304 4243 1336
rect 4253 1284 4259 1357
rect 4269 1344 4275 1377
rect 4285 1344 4291 1356
rect 4301 1344 4307 1416
rect 4317 1404 4323 1436
rect 4333 1384 4339 1456
rect 4397 1344 4403 1476
rect 4413 1344 4419 1376
rect 4461 1344 4467 1436
rect 4477 1344 4483 1376
rect 4029 1144 4035 1236
rect 4013 1104 4019 1116
rect 4093 1104 4099 1136
rect 3885 903 3891 1076
rect 4157 1064 4163 1076
rect 4173 1063 4179 1116
rect 4253 1104 4259 1116
rect 4164 1057 4179 1063
rect 3917 943 3923 1036
rect 3949 944 3955 1036
rect 4061 1024 4067 1056
rect 4221 1043 4227 1076
rect 4212 1037 4227 1043
rect 4285 964 4291 1036
rect 3917 937 3939 943
rect 3933 924 3939 937
rect 3933 904 3939 916
rect 3885 897 3900 903
rect 4013 903 4019 956
rect 4125 904 4131 956
rect 4301 944 4307 1036
rect 4365 984 4371 1236
rect 4397 1144 4403 1336
rect 4461 1304 4467 1336
rect 4429 1144 4435 1236
rect 4397 1084 4403 1136
rect 4429 1004 4435 1116
rect 4461 1083 4467 1136
rect 4477 1124 4483 1156
rect 4525 1144 4531 1316
rect 4541 1304 4547 1396
rect 4557 1324 4563 1436
rect 4589 1404 4595 1496
rect 4637 1464 4643 1536
rect 4669 1484 4675 1576
rect 4701 1524 4707 1556
rect 4717 1524 4723 1576
rect 4749 1544 4755 1656
rect 4824 1606 4830 1614
rect 4838 1606 4844 1614
rect 4852 1606 4858 1614
rect 4866 1606 4872 1614
rect 4925 1584 4931 1596
rect 4973 1584 4979 1636
rect 4733 1504 4739 1536
rect 4797 1484 4803 1516
rect 4669 1384 4675 1476
rect 4845 1464 4851 1556
rect 4861 1504 4867 1576
rect 4685 1364 4691 1436
rect 4717 1384 4723 1416
rect 4813 1384 4819 1436
rect 4701 1344 4707 1356
rect 4621 1324 4627 1336
rect 4605 1304 4611 1316
rect 4749 1264 4755 1336
rect 4877 1324 4883 1576
rect 4909 1484 4915 1536
rect 4941 1524 4947 1556
rect 4925 1504 4931 1516
rect 4957 1484 4963 1496
rect 4973 1484 4979 1516
rect 5021 1464 5027 1556
rect 5037 1543 5043 1636
rect 5085 1584 5091 1616
rect 5037 1537 5059 1543
rect 4925 1384 4931 1456
rect 4989 1424 4995 1436
rect 4989 1384 4995 1396
rect 4957 1340 4963 1356
rect 5021 1344 5027 1356
rect 5053 1343 5059 1537
rect 5108 1517 5123 1523
rect 5117 1464 5123 1517
rect 5133 1483 5139 1496
rect 5149 1484 5155 1516
rect 5165 1504 5171 1536
rect 5181 1504 5187 1697
rect 5133 1477 5148 1483
rect 5197 1483 5203 1636
rect 5213 1524 5219 1696
rect 5229 1504 5235 1536
rect 5261 1524 5267 1576
rect 5245 1484 5251 1516
rect 5188 1477 5203 1483
rect 5133 1404 5139 1436
rect 5053 1337 5068 1343
rect 4861 1303 4867 1316
rect 4989 1304 4995 1336
rect 4861 1297 4876 1303
rect 4493 1124 4499 1136
rect 4557 1104 4563 1236
rect 4637 1124 4643 1136
rect 4653 1104 4659 1236
rect 4824 1206 4830 1214
rect 4838 1206 4844 1214
rect 4852 1206 4858 1214
rect 4866 1206 4872 1214
rect 4525 1084 4531 1096
rect 4461 1077 4483 1083
rect 4477 984 4483 1077
rect 4557 1064 4563 1076
rect 4349 964 4355 976
rect 4157 924 4163 936
rect 4461 924 4467 976
rect 4509 924 4515 1056
rect 4541 1024 4547 1036
rect 4589 944 4595 1096
rect 4621 1064 4627 1076
rect 4669 1044 4675 1136
rect 4717 1084 4723 1136
rect 4909 1104 4915 1296
rect 4973 1184 4979 1256
rect 4957 1084 4963 1176
rect 4973 1144 4979 1176
rect 4989 1123 4995 1296
rect 5037 1284 5043 1296
rect 5133 1284 5139 1356
rect 5085 1124 5091 1236
rect 4989 1117 5004 1123
rect 5005 1104 5011 1116
rect 5085 1104 5091 1116
rect 4749 1044 4755 1056
rect 4669 984 4675 996
rect 4717 984 4723 1036
rect 4797 1024 4803 1056
rect 4813 1024 4819 1076
rect 4989 1064 4995 1096
rect 5053 1064 5059 1076
rect 4893 984 4899 1036
rect 4813 964 4819 976
rect 4004 897 4019 903
rect 4141 884 4147 916
rect 3597 664 3603 876
rect 3661 684 3667 756
rect 3693 724 3699 856
rect 3773 764 3779 836
rect 3805 784 3811 836
rect 3677 684 3683 716
rect 3693 683 3699 716
rect 3725 684 3731 756
rect 3885 744 3891 836
rect 3933 724 3939 836
rect 4013 737 4044 743
rect 4013 723 4019 737
rect 3956 717 4019 723
rect 3693 677 3715 683
rect 3453 624 3459 656
rect 3549 644 3555 656
rect 3645 644 3651 676
rect 3709 664 3715 677
rect 3981 664 3987 676
rect 3453 544 3459 616
rect 3469 584 3475 636
rect 3469 544 3475 576
rect 3549 544 3555 636
rect 3437 504 3443 536
rect 3485 524 3491 536
rect 3469 504 3475 516
rect 2941 343 2947 436
rect 2941 337 2963 343
rect 2797 324 2803 336
rect 2957 324 2963 337
rect 2797 297 2860 303
rect 2797 283 2803 297
rect 2941 284 2947 316
rect 2973 284 2979 316
rect 2989 284 2995 436
rect 3005 304 3011 336
rect 3021 284 3027 376
rect 3101 344 3107 436
rect 2733 277 2803 283
rect 2733 263 2739 277
rect 2877 264 2883 276
rect 3053 264 3059 316
rect 3085 303 3091 336
rect 3117 324 3123 376
rect 3085 297 3100 303
rect 3133 303 3139 336
rect 3108 297 3139 303
rect 3149 284 3155 296
rect 3197 284 3203 436
rect 3533 404 3539 536
rect 3565 524 3571 616
rect 3597 584 3603 616
rect 3613 524 3619 636
rect 3645 544 3651 616
rect 3677 524 3683 616
rect 3693 544 3699 656
rect 3789 624 3795 636
rect 3837 603 3843 636
rect 3821 597 3843 603
rect 3821 564 3827 597
rect 3837 564 3843 576
rect 3709 544 3715 556
rect 3773 544 3779 556
rect 3837 544 3843 556
rect 3885 544 3891 576
rect 3917 564 3923 636
rect 3901 544 3907 556
rect 3725 524 3731 536
rect 3549 504 3555 516
rect 3725 504 3731 516
rect 3757 504 3763 536
rect 3789 504 3795 516
rect 3821 504 3827 536
rect 3837 504 3843 516
rect 3645 464 3651 496
rect 3853 484 3859 516
rect 3885 504 3891 536
rect 3901 484 3907 516
rect 3229 284 3235 356
rect 3277 324 3283 336
rect 3309 324 3315 356
rect 3533 344 3539 376
rect 3581 344 3587 376
rect 3597 344 3603 356
rect 3245 304 3251 316
rect 3389 304 3395 316
rect 3293 284 3299 296
rect 3405 284 3411 316
rect 3485 304 3491 316
rect 3517 304 3523 316
rect 3597 304 3603 316
rect 3197 264 3203 276
rect 2653 257 2739 263
rect 2605 164 2611 236
rect 2093 84 2099 96
rect 1949 77 1971 83
rect 1725 44 1731 76
rect 1949 63 1955 77
rect 1908 57 1955 63
rect 2109 63 2115 96
rect 2125 84 2131 96
rect 2285 84 2291 136
rect 2301 64 2307 116
rect 2349 84 2355 136
rect 2365 64 2371 116
rect 2381 104 2387 136
rect 2445 104 2451 136
rect 2557 124 2563 136
rect 2637 124 2643 196
rect 2653 184 2659 236
rect 2669 184 2675 216
rect 2669 104 2675 136
rect 2701 84 2707 136
rect 2733 104 2739 236
rect 2797 144 2803 196
rect 2893 184 2899 256
rect 3037 224 3043 236
rect 2381 64 2387 76
rect 2717 64 2723 96
rect 2749 64 2755 116
rect 2765 84 2771 136
rect 2109 57 2188 63
rect 2813 44 2819 116
rect 2829 64 2835 116
rect 2845 84 2851 136
rect 2877 84 2883 136
rect 2893 124 2899 156
rect 2925 144 2931 176
rect 2909 64 2915 116
rect 653 37 739 43
rect 2941 43 2947 176
rect 3037 164 3043 196
rect 2957 84 2963 136
rect 2973 124 2979 156
rect 3005 144 3011 156
rect 3021 123 3027 156
rect 3037 144 3043 156
rect 3069 144 3075 196
rect 3085 144 3091 236
rect 3213 224 3219 236
rect 3117 184 3123 196
rect 3133 144 3139 176
rect 2996 117 3027 123
rect 3101 117 3116 123
rect 2973 84 2979 116
rect 2957 64 2963 76
rect 3053 44 3059 116
rect 2884 37 2947 43
rect 2797 24 2803 36
rect 2957 24 2963 36
rect 3037 24 3043 36
rect 3069 23 3075 116
rect 3101 24 3107 117
rect 3149 103 3155 176
rect 3124 97 3155 103
rect 3213 103 3219 196
rect 3229 184 3235 216
rect 3261 124 3267 236
rect 3304 206 3310 214
rect 3318 206 3324 214
rect 3332 206 3338 214
rect 3346 206 3352 214
rect 3357 104 3363 176
rect 3373 124 3379 256
rect 3421 163 3427 276
rect 3469 204 3475 296
rect 3613 244 3619 316
rect 3629 304 3635 316
rect 3677 283 3683 436
rect 3709 304 3715 456
rect 3933 404 3939 636
rect 3949 604 3955 636
rect 3949 504 3955 556
rect 3997 524 4003 536
rect 4013 524 4019 636
rect 4029 624 4035 716
rect 4077 684 4083 836
rect 4109 783 4115 836
rect 4109 777 4131 783
rect 4109 704 4115 756
rect 4125 704 4131 777
rect 4237 764 4243 916
rect 4253 904 4259 916
rect 4509 904 4515 916
rect 4573 884 4579 936
rect 4413 784 4419 796
rect 4605 784 4611 896
rect 4637 884 4643 936
rect 4157 724 4163 756
rect 4077 664 4083 676
rect 4061 624 4067 656
rect 4061 524 4067 536
rect 3997 504 4003 516
rect 4077 504 4083 516
rect 4109 504 4115 656
rect 4157 644 4163 676
rect 4157 544 4163 636
rect 4173 584 4179 636
rect 3997 424 4003 436
rect 3725 304 3731 396
rect 3709 284 3715 296
rect 3668 277 3683 283
rect 3693 264 3699 276
rect 3757 264 3763 316
rect 3853 304 3859 396
rect 3885 304 3891 356
rect 3821 264 3827 296
rect 3917 264 3923 356
rect 3933 284 3939 316
rect 4013 304 4019 496
rect 4029 364 4035 436
rect 4061 284 4067 456
rect 4109 444 4115 476
rect 4125 464 4131 516
rect 4189 504 4195 636
rect 4205 564 4211 716
rect 4221 684 4227 696
rect 4253 684 4259 696
rect 4269 664 4275 736
rect 4333 684 4339 776
rect 4349 684 4355 696
rect 4365 684 4371 736
rect 4381 704 4387 776
rect 4317 584 4323 636
rect 4365 564 4371 616
rect 4269 524 4275 536
rect 4301 523 4307 556
rect 4397 544 4403 756
rect 4429 684 4435 776
rect 4461 724 4467 736
rect 4548 717 4563 723
rect 4509 664 4515 696
rect 4525 644 4531 676
rect 4477 604 4483 636
rect 4413 524 4419 576
rect 4525 524 4531 556
rect 4541 544 4547 696
rect 4557 684 4563 717
rect 4589 684 4595 736
rect 4573 664 4579 676
rect 4557 544 4563 636
rect 4605 624 4611 696
rect 4621 584 4627 836
rect 4637 724 4643 736
rect 4653 724 4659 796
rect 4653 564 4659 636
rect 4669 564 4675 956
rect 4781 924 4787 956
rect 4765 884 4771 916
rect 4813 904 4819 956
rect 5005 944 5011 1056
rect 5021 944 5027 976
rect 5037 944 5043 956
rect 5101 944 5107 996
rect 5133 984 5139 1076
rect 5133 944 5139 956
rect 4925 923 4931 936
rect 5005 924 5011 936
rect 5069 924 5075 936
rect 5101 924 5107 936
rect 5149 924 5155 1456
rect 5213 1364 5219 1436
rect 5197 1324 5203 1356
rect 5181 1284 5187 1316
rect 5229 1304 5235 1416
rect 5261 1404 5267 1476
rect 5277 1464 5283 1556
rect 5261 1344 5267 1376
rect 5277 1364 5283 1396
rect 5309 1364 5315 1696
rect 5325 1584 5331 1696
rect 5341 1504 5347 1616
rect 5373 1484 5379 1596
rect 5533 1564 5539 1876
rect 5549 1784 5555 1877
rect 5565 1864 5571 1876
rect 5709 1864 5715 1876
rect 5773 1863 5779 2294
rect 5933 2277 5948 2283
rect 5821 2184 5827 2236
rect 5917 2184 5923 2276
rect 5933 2184 5939 2277
rect 5853 2177 5868 2183
rect 5853 2144 5859 2177
rect 5901 2177 5916 2183
rect 5869 2104 5875 2116
rect 5901 2104 5907 2177
rect 5917 2144 5923 2176
rect 5949 2164 5955 2236
rect 5965 2204 5971 2297
rect 5949 2124 5955 2156
rect 5997 2143 6003 3176
rect 6013 3004 6019 3136
rect 6045 3084 6051 3296
rect 6077 3104 6083 3236
rect 6093 3144 6099 3336
rect 6125 3304 6131 3336
rect 6141 3317 6156 3323
rect 6141 3304 6147 3317
rect 6029 2964 6035 3016
rect 6077 2924 6083 3036
rect 6013 2904 6019 2916
rect 6077 2883 6083 2916
rect 6093 2904 6099 3016
rect 6109 2924 6115 2936
rect 6077 2877 6092 2883
rect 6125 2784 6131 3256
rect 6173 3204 6179 3336
rect 6189 3264 6195 3516
rect 6237 3484 6243 3696
rect 6301 3684 6307 3876
rect 6317 3724 6323 3836
rect 6333 3744 6339 3856
rect 6349 3824 6355 3877
rect 6365 3844 6371 3856
rect 6381 3804 6387 3836
rect 6381 3744 6387 3756
rect 6317 3684 6323 3696
rect 6285 3664 6291 3676
rect 6221 3344 6227 3436
rect 6221 3304 6227 3316
rect 6253 3304 6259 3576
rect 6269 3524 6275 3536
rect 6285 3404 6291 3636
rect 6301 3484 6307 3656
rect 6317 3604 6323 3676
rect 6333 3584 6339 3716
rect 6333 3544 6339 3556
rect 6349 3523 6355 3536
rect 6365 3524 6371 3716
rect 6397 3624 6403 4056
rect 6413 3864 6419 4016
rect 6445 3984 6451 4036
rect 6445 3924 6451 3936
rect 6429 3864 6435 3916
rect 6413 3764 6419 3836
rect 6429 3744 6435 3796
rect 6445 3724 6451 3836
rect 6333 3517 6355 3523
rect 6221 3124 6227 3236
rect 6157 3104 6163 3116
rect 6237 3104 6243 3236
rect 6269 3224 6275 3236
rect 6285 3203 6291 3276
rect 6269 3197 6291 3203
rect 6269 3184 6275 3197
rect 6301 3184 6307 3436
rect 6317 3224 6323 3356
rect 6157 2984 6163 2996
rect 6189 2824 6195 2936
rect 6221 2784 6227 3036
rect 6253 2844 6259 2918
rect 6077 2724 6083 2736
rect 6061 2504 6067 2596
rect 6093 2584 6099 2696
rect 6109 2544 6115 2576
rect 6045 2323 6051 2436
rect 6036 2317 6051 2323
rect 6013 2304 6019 2316
rect 6093 2284 6099 2316
rect 5981 2137 6003 2143
rect 5917 2104 5923 2116
rect 5933 1964 5939 2036
rect 5805 1904 5811 1916
rect 5869 1904 5875 1916
rect 5757 1857 5779 1863
rect 5565 1744 5571 1776
rect 5492 1537 5507 1543
rect 5405 1484 5411 1536
rect 5341 1404 5347 1476
rect 5357 1384 5363 1476
rect 5165 1104 5171 1236
rect 5245 1124 5251 1236
rect 5229 1117 5244 1123
rect 5229 1104 5235 1117
rect 5261 1104 5267 1176
rect 5229 1084 5235 1096
rect 5213 1064 5219 1076
rect 5277 1064 5283 1356
rect 5341 1344 5347 1356
rect 5405 1344 5411 1436
rect 5437 1364 5443 1436
rect 5469 1404 5475 1496
rect 5485 1464 5491 1516
rect 5501 1384 5507 1537
rect 5549 1444 5555 1696
rect 5677 1684 5683 1756
rect 5693 1724 5699 1736
rect 5629 1604 5635 1636
rect 5629 1504 5635 1556
rect 5565 1484 5571 1496
rect 5677 1484 5683 1516
rect 5661 1444 5667 1476
rect 5581 1364 5587 1436
rect 5613 1384 5619 1396
rect 5645 1364 5651 1436
rect 5661 1384 5667 1436
rect 5325 1324 5331 1336
rect 5373 1284 5379 1336
rect 5421 1264 5427 1356
rect 5549 1284 5555 1336
rect 5309 1184 5315 1236
rect 5293 1124 5299 1156
rect 5325 1084 5331 1096
rect 5341 1084 5347 1096
rect 5373 1084 5379 1096
rect 4916 917 4931 923
rect 4925 864 4931 876
rect 4824 806 4830 814
rect 4838 806 4844 814
rect 4852 806 4858 814
rect 4866 806 4872 814
rect 4733 724 4739 796
rect 5021 784 5027 876
rect 5133 864 5139 916
rect 5165 744 5171 1016
rect 5181 943 5187 1036
rect 5197 963 5203 1036
rect 5277 964 5283 996
rect 5197 957 5219 963
rect 5213 944 5219 957
rect 5277 944 5283 956
rect 5293 944 5299 956
rect 5181 937 5196 943
rect 5197 924 5203 936
rect 5261 924 5267 936
rect 5181 784 5187 916
rect 5293 784 5299 856
rect 4685 644 4691 676
rect 4701 564 4707 596
rect 4717 564 4723 696
rect 4749 644 4755 676
rect 4781 664 4787 716
rect 4797 664 4803 716
rect 4893 704 4899 736
rect 5069 724 5075 736
rect 5005 704 5011 716
rect 5021 704 5027 716
rect 4845 684 4851 696
rect 4829 644 4835 676
rect 4813 624 4819 636
rect 4292 517 4307 523
rect 4285 504 4291 516
rect 4381 504 4387 516
rect 4253 484 4259 496
rect 4269 464 4275 476
rect 4093 284 4099 436
rect 4125 344 4131 436
rect 4141 304 4147 316
rect 4157 304 4163 456
rect 4173 344 4179 436
rect 4221 344 4227 356
rect 4301 344 4307 356
rect 4269 304 4275 316
rect 4285 304 4291 336
rect 4381 324 4387 496
rect 4413 484 4419 516
rect 4397 344 4403 356
rect 4413 304 4419 416
rect 4445 344 4451 516
rect 4461 424 4467 476
rect 4429 324 4435 336
rect 4461 284 4467 416
rect 4477 324 4483 436
rect 3405 157 3427 163
rect 3405 124 3411 157
rect 3421 104 3427 136
rect 3437 124 3443 156
rect 3501 104 3507 116
rect 3517 104 3523 176
rect 3213 97 3228 103
rect 3181 24 3187 96
rect 3453 84 3459 96
rect 3549 84 3555 236
rect 3565 104 3571 116
rect 3581 104 3587 196
rect 3629 124 3635 156
rect 3645 104 3651 136
rect 3661 124 3667 156
rect 3709 144 3715 156
rect 3565 64 3571 76
rect 3613 64 3619 76
rect 3629 64 3635 96
rect 3677 64 3683 136
rect 3757 124 3763 236
rect 3773 144 3779 236
rect 3789 224 3795 236
rect 3805 164 3811 216
rect 3869 164 3875 216
rect 3885 164 3891 236
rect 3773 104 3779 116
rect 3773 64 3779 96
rect 3837 84 3843 136
rect 3917 124 3923 256
rect 3933 184 3939 276
rect 4093 264 4099 276
rect 4493 264 4499 496
rect 4525 364 4531 436
rect 4509 284 4515 336
rect 4541 324 4547 416
rect 4557 384 4563 516
rect 4653 344 4659 536
rect 4669 524 4675 536
rect 4797 524 4803 596
rect 4829 524 4835 616
rect 4909 564 4915 676
rect 4925 644 4931 696
rect 4989 664 4995 696
rect 4909 544 4915 556
rect 4941 504 4947 636
rect 4973 564 4979 596
rect 5037 564 5043 656
rect 5069 584 5075 716
rect 5101 684 5107 716
rect 5309 684 5315 1056
rect 5373 984 5379 1076
rect 5389 1004 5395 1076
rect 5421 1024 5427 1156
rect 5437 1124 5443 1136
rect 5485 1124 5491 1136
rect 5444 1117 5459 1123
rect 5453 1084 5459 1117
rect 5332 977 5347 983
rect 5341 904 5347 977
rect 5373 924 5379 976
rect 5389 944 5395 996
rect 5421 964 5427 996
rect 5437 964 5443 996
rect 5453 984 5459 1016
rect 5469 924 5475 1036
rect 5485 1024 5491 1116
rect 5501 1084 5507 1116
rect 5501 1024 5507 1076
rect 5485 944 5491 996
rect 5501 924 5507 976
rect 5405 704 5411 836
rect 5469 724 5475 756
rect 5517 704 5523 1196
rect 5533 1124 5539 1136
rect 5565 1083 5571 1336
rect 5645 1324 5651 1356
rect 5581 1264 5587 1316
rect 5581 1104 5587 1256
rect 5629 1124 5635 1136
rect 5613 1084 5619 1096
rect 5565 1077 5587 1083
rect 5533 904 5539 1016
rect 5581 984 5587 1077
rect 5597 964 5603 1036
rect 5629 904 5635 1116
rect 5645 824 5651 1256
rect 5677 1063 5683 1076
rect 5677 1057 5692 1063
rect 5693 1024 5699 1056
rect 5709 1024 5715 1816
rect 5757 1764 5763 1857
rect 5821 1844 5827 1876
rect 5853 1864 5859 1896
rect 5885 1844 5891 1876
rect 5933 1864 5939 1896
rect 5837 1804 5843 1836
rect 5725 1224 5731 1756
rect 5741 1724 5747 1736
rect 5789 1724 5795 1756
rect 5773 1684 5779 1696
rect 5821 1684 5827 1716
rect 5885 1704 5891 1716
rect 5901 1704 5907 1756
rect 5933 1744 5939 1756
rect 5741 1484 5747 1516
rect 5805 1504 5811 1516
rect 5757 1363 5763 1496
rect 5773 1444 5779 1476
rect 5789 1464 5795 1476
rect 5821 1444 5827 1456
rect 5757 1357 5779 1363
rect 5773 1324 5779 1357
rect 5725 1123 5731 1136
rect 5725 1117 5740 1123
rect 5661 944 5667 956
rect 5677 924 5683 936
rect 5709 924 5715 976
rect 5725 944 5731 996
rect 5741 964 5747 1116
rect 5789 1064 5795 1436
rect 5821 1364 5827 1436
rect 5837 1384 5843 1456
rect 5853 1384 5859 1496
rect 5901 1484 5907 1636
rect 5869 1404 5875 1476
rect 5901 1464 5907 1476
rect 5917 1464 5923 1476
rect 5821 1344 5827 1356
rect 5869 1324 5875 1376
rect 5885 1344 5891 1416
rect 5933 1404 5939 1436
rect 5949 1384 5955 1936
rect 5965 1644 5971 2036
rect 5981 1944 5987 2137
rect 5997 2104 6003 2116
rect 6013 2104 6019 2196
rect 6045 2144 6051 2176
rect 6061 2144 6067 2156
rect 6061 2124 6067 2136
rect 6077 2124 6083 2236
rect 6109 2184 6115 2296
rect 6029 1984 6035 2036
rect 6077 2004 6083 2036
rect 5997 1884 6003 1896
rect 6013 1884 6019 1896
rect 5981 1824 5987 1836
rect 6093 1804 6099 1876
rect 6109 1824 6115 1896
rect 5981 1744 5987 1776
rect 6045 1724 6051 1756
rect 6109 1724 6115 1756
rect 6125 1684 6131 2756
rect 6173 2684 6179 2696
rect 6237 2604 6243 2694
rect 6173 2564 6179 2596
rect 6141 2344 6147 2516
rect 6221 2504 6227 2516
rect 6253 2383 6259 2776
rect 6269 2644 6275 3116
rect 6301 2944 6307 3076
rect 6333 3024 6339 3517
rect 6365 3504 6371 3516
rect 6381 3504 6387 3556
rect 6413 3444 6419 3676
rect 6461 3664 6467 4176
rect 6477 4124 6483 4156
rect 6477 3944 6483 4036
rect 6493 3984 6499 4317
rect 6525 4284 6531 4296
rect 6525 4124 6531 4156
rect 6541 4044 6547 4276
rect 6557 4264 6563 4316
rect 6557 4184 6563 4236
rect 6557 4144 6563 4156
rect 6573 4064 6579 4776
rect 6717 4764 6723 4816
rect 6589 4324 6595 4436
rect 6605 4304 6611 4316
rect 6589 4204 6595 4276
rect 6621 4244 6627 4736
rect 6637 4544 6643 4636
rect 6589 4104 6595 4116
rect 6477 3884 6483 3896
rect 6493 3864 6499 3916
rect 6541 3904 6547 3936
rect 6525 3884 6531 3896
rect 6557 3884 6563 3996
rect 6573 3884 6579 3896
rect 6477 3644 6483 3856
rect 6509 3844 6515 3876
rect 6509 3744 6515 3836
rect 6541 3784 6547 3816
rect 6589 3783 6595 3936
rect 6605 3904 6611 4236
rect 6621 3904 6627 4036
rect 6621 3804 6627 3896
rect 6589 3777 6611 3783
rect 6605 3764 6611 3777
rect 6461 3544 6467 3636
rect 6493 3523 6499 3656
rect 6477 3517 6499 3523
rect 6429 3464 6435 3496
rect 6477 3484 6483 3517
rect 6461 3424 6467 3436
rect 6477 3424 6483 3476
rect 6493 3464 6499 3496
rect 6509 3484 6515 3596
rect 6525 3504 6531 3636
rect 6573 3523 6579 3576
rect 6573 3517 6595 3523
rect 6541 3464 6547 3516
rect 6525 3344 6531 3436
rect 6365 3084 6371 3216
rect 6381 3044 6387 3176
rect 6429 3023 6435 3296
rect 6445 3144 6451 3216
rect 6461 3124 6467 3336
rect 6525 3262 6531 3300
rect 6509 3184 6515 3216
rect 6477 3064 6483 3096
rect 6413 3017 6435 3023
rect 6381 2944 6387 2976
rect 6285 2684 6291 2936
rect 6397 2784 6403 2916
rect 6413 2784 6419 3017
rect 6461 2984 6467 3036
rect 6477 2984 6483 3036
rect 6493 3004 6499 3176
rect 6541 3143 6547 3416
rect 6557 3144 6563 3496
rect 6525 3137 6547 3143
rect 6509 3044 6515 3136
rect 6525 3084 6531 3137
rect 6573 3104 6579 3456
rect 6589 3104 6595 3517
rect 6605 3464 6611 3716
rect 6621 3704 6627 3776
rect 6605 3144 6611 3436
rect 6621 3304 6627 3616
rect 6621 3104 6627 3156
rect 6445 2924 6451 2936
rect 6493 2924 6499 2976
rect 6429 2884 6435 2896
rect 6381 2704 6387 2716
rect 6493 2704 6499 2776
rect 6285 2564 6291 2676
rect 6445 2544 6451 2676
rect 6285 2504 6291 2518
rect 6253 2377 6275 2383
rect 6269 2302 6275 2377
rect 6413 2364 6419 2436
rect 6173 2184 6179 2276
rect 6205 2264 6211 2276
rect 6237 2244 6243 2276
rect 6173 2123 6179 2176
rect 6173 2117 6188 2123
rect 6205 2084 6211 2116
rect 6141 1764 6147 1916
rect 6189 1864 6195 2036
rect 6141 1704 6147 1716
rect 6173 1704 6179 1716
rect 6189 1684 6195 1716
rect 6045 1624 6051 1636
rect 5965 1504 5971 1556
rect 5981 1484 5987 1536
rect 6029 1503 6035 1576
rect 6061 1504 6067 1636
rect 6077 1504 6083 1556
rect 6029 1497 6044 1503
rect 5997 1464 6003 1476
rect 6061 1424 6067 1476
rect 5805 1304 5811 1316
rect 5885 1284 5891 1316
rect 5901 1144 5907 1376
rect 5949 1344 5955 1356
rect 5821 1088 5827 1096
rect 5805 1080 5820 1083
rect 5805 1077 5827 1080
rect 5789 984 5795 1036
rect 5805 984 5811 1077
rect 5773 944 5779 976
rect 5821 924 5827 1056
rect 5869 944 5875 1036
rect 5709 784 5715 856
rect 5741 784 5747 836
rect 5652 717 5667 723
rect 5405 684 5411 696
rect 5197 644 5203 676
rect 5309 664 5315 676
rect 5085 624 5091 636
rect 5133 604 5139 636
rect 5005 484 5011 496
rect 4653 304 4659 336
rect 4685 284 4691 376
rect 3949 123 3955 216
rect 4125 184 4131 256
rect 3997 144 4003 176
rect 4157 144 4163 236
rect 3981 124 3987 136
rect 3933 117 3955 123
rect 3933 104 3939 117
rect 4013 104 4019 136
rect 4205 124 4211 236
rect 4477 224 4483 236
rect 4429 144 4435 156
rect 4621 144 4627 236
rect 4685 184 4691 236
rect 4669 144 4675 156
rect 4701 144 4707 436
rect 4733 304 4739 436
rect 4717 264 4723 276
rect 4781 264 4787 316
rect 4797 304 4803 436
rect 4824 406 4830 414
rect 4838 406 4844 414
rect 4852 406 4858 414
rect 4866 406 4872 414
rect 4797 144 4803 176
rect 4877 164 4883 316
rect 4925 264 4931 436
rect 5037 324 5043 556
rect 5085 524 5091 576
rect 4973 164 4979 256
rect 5005 184 5011 236
rect 5037 184 5043 236
rect 4877 144 4883 156
rect 5053 144 5059 456
rect 5069 324 5075 516
rect 5117 304 5123 536
rect 5133 524 5139 536
rect 5165 504 5171 636
rect 5277 624 5283 656
rect 5405 624 5411 656
rect 5181 584 5187 616
rect 5213 524 5219 556
rect 5293 544 5299 556
rect 5181 464 5187 496
rect 5213 324 5219 516
rect 5325 504 5331 616
rect 5421 603 5427 696
rect 5437 644 5443 696
rect 5501 684 5507 696
rect 5405 597 5427 603
rect 5357 544 5363 576
rect 5373 564 5379 596
rect 5245 444 5251 496
rect 5277 324 5283 476
rect 5293 324 5299 436
rect 5165 317 5180 323
rect 5069 244 5075 276
rect 5165 264 5171 317
rect 5229 284 5235 296
rect 5277 284 5283 316
rect 5389 304 5395 536
rect 5405 524 5411 597
rect 5453 584 5459 656
rect 5549 644 5555 676
rect 5421 544 5427 576
rect 5501 564 5507 576
rect 5517 544 5523 616
rect 5565 544 5571 636
rect 5581 583 5587 716
rect 5581 577 5596 583
rect 5613 564 5619 696
rect 5661 664 5667 717
rect 5805 704 5811 876
rect 5885 864 5891 956
rect 5821 704 5827 716
rect 5677 664 5683 676
rect 5789 624 5795 676
rect 5805 644 5811 676
rect 5661 524 5667 616
rect 5741 524 5747 536
rect 5405 464 5411 516
rect 5620 497 5635 503
rect 5405 344 5411 436
rect 5629 384 5635 497
rect 5661 424 5667 436
rect 5725 384 5731 496
rect 5629 344 5635 376
rect 5741 364 5747 436
rect 5805 384 5811 556
rect 5821 544 5827 656
rect 5837 604 5843 696
rect 5853 683 5859 836
rect 5853 677 5875 683
rect 5853 644 5859 656
rect 5869 584 5875 677
rect 5885 544 5891 636
rect 5901 564 5907 1116
rect 5917 663 5923 1176
rect 5933 1104 5939 1316
rect 5949 1304 5955 1336
rect 5933 1044 5939 1076
rect 5965 1044 5971 1136
rect 5981 1124 5987 1376
rect 5997 1284 6003 1396
rect 5965 904 5971 936
rect 5997 903 6003 1196
rect 6013 1124 6019 1236
rect 6029 1123 6035 1376
rect 6061 1364 6067 1416
rect 6077 1324 6083 1356
rect 6077 1224 6083 1236
rect 6045 1144 6051 1156
rect 6077 1124 6083 1156
rect 6029 1117 6051 1123
rect 6045 984 6051 1117
rect 6061 1044 6067 1096
rect 6093 984 6099 1636
rect 6109 1444 6115 1516
rect 6141 1484 6147 1516
rect 6125 1464 6131 1476
rect 6157 1463 6163 1676
rect 6205 1663 6211 2056
rect 6221 2024 6227 2216
rect 6237 2104 6243 2156
rect 6269 2144 6275 2176
rect 6301 2104 6307 2156
rect 6333 2144 6339 2176
rect 6365 2064 6371 2356
rect 6429 2244 6435 2276
rect 6397 2224 6403 2236
rect 6381 2104 6387 2156
rect 6413 2124 6419 2176
rect 6461 2164 6467 2256
rect 6461 2124 6467 2136
rect 6429 2084 6435 2116
rect 6237 1903 6243 2036
rect 6413 1924 6419 2076
rect 6253 1904 6259 1916
rect 6301 1904 6307 1916
rect 6333 1904 6339 1916
rect 6413 1904 6419 1916
rect 6429 1904 6435 1936
rect 6228 1897 6243 1903
rect 6221 1884 6227 1896
rect 6349 1884 6355 1896
rect 6221 1704 6227 1736
rect 6237 1724 6243 1876
rect 6269 1844 6275 1876
rect 6237 1704 6243 1716
rect 6253 1684 6259 1716
rect 6189 1657 6211 1663
rect 6173 1564 6179 1636
rect 6141 1457 6163 1463
rect 6109 1344 6115 1356
rect 6125 1324 6131 1396
rect 6141 1264 6147 1457
rect 6157 1364 6163 1416
rect 6189 1384 6195 1657
rect 6269 1624 6275 1736
rect 6317 1684 6323 1876
rect 6349 1764 6355 1816
rect 6365 1804 6371 1876
rect 6381 1824 6387 1896
rect 6429 1884 6435 1896
rect 6221 1504 6227 1576
rect 6173 1364 6179 1376
rect 6109 1084 6115 1136
rect 6125 1104 6131 1216
rect 6157 1184 6163 1296
rect 6189 1284 6195 1316
rect 6205 1244 6211 1456
rect 6221 1424 6227 1476
rect 6237 1243 6243 1616
rect 6269 1584 6275 1596
rect 6349 1544 6355 1676
rect 6292 1537 6316 1543
rect 6253 1524 6259 1536
rect 6349 1524 6355 1536
rect 6365 1524 6371 1756
rect 6381 1543 6387 1776
rect 6397 1724 6403 1876
rect 6429 1724 6435 1736
rect 6445 1724 6451 2076
rect 6461 1924 6467 2036
rect 6477 1944 6483 2436
rect 6509 2304 6515 3016
rect 6525 2863 6531 3056
rect 6541 2884 6547 2916
rect 6525 2857 6547 2863
rect 6509 2004 6515 2236
rect 6525 2144 6531 2836
rect 6541 2584 6547 2857
rect 6557 2784 6563 3036
rect 6573 2984 6579 3016
rect 6589 2924 6595 3036
rect 6605 2603 6611 3036
rect 6621 3004 6627 3076
rect 6637 3024 6643 4256
rect 6717 3224 6723 4696
rect 6637 2864 6643 2936
rect 6621 2664 6627 2836
rect 6589 2597 6611 2603
rect 6589 2263 6595 2597
rect 6589 2257 6611 2263
rect 6525 1984 6531 2036
rect 6541 1964 6547 2216
rect 6573 2103 6579 2136
rect 6564 2097 6579 2103
rect 6573 1984 6579 2076
rect 6477 1904 6483 1936
rect 6541 1924 6547 1936
rect 6509 1884 6515 1916
rect 6461 1744 6467 1836
rect 6525 1744 6531 1916
rect 6541 1724 6547 1896
rect 6557 1884 6563 1976
rect 6461 1683 6467 1696
rect 6525 1684 6531 1716
rect 6461 1677 6483 1683
rect 6397 1564 6403 1636
rect 6381 1537 6419 1543
rect 6269 1404 6275 1496
rect 6381 1484 6387 1496
rect 6269 1304 6275 1316
rect 6221 1237 6243 1243
rect 6141 1104 6147 1116
rect 6173 1104 6179 1216
rect 6205 1104 6211 1136
rect 6189 1084 6195 1096
rect 6125 1064 6131 1076
rect 6205 1044 6211 1076
rect 6029 904 6035 936
rect 5997 897 6019 903
rect 5965 864 5971 896
rect 5933 744 5939 836
rect 5981 764 5987 836
rect 6013 744 6019 897
rect 6061 884 6067 976
rect 6125 884 6131 976
rect 6157 924 6163 936
rect 5965 684 5971 736
rect 6045 724 6051 836
rect 5981 704 5987 716
rect 5997 704 6003 716
rect 6004 697 6019 703
rect 6013 664 6019 697
rect 6045 703 6051 716
rect 6045 697 6060 703
rect 5917 657 5939 663
rect 5917 624 5923 636
rect 5917 544 5923 616
rect 5837 524 5843 536
rect 5885 504 5891 516
rect 5837 384 5843 436
rect 5453 302 5459 336
rect 5325 244 5331 276
rect 3917 64 3923 96
rect 4045 64 4051 96
rect 4253 83 4259 116
rect 4253 77 4268 83
rect 4493 83 4499 116
rect 4989 104 4995 116
rect 5101 104 5107 116
rect 4941 84 4947 96
rect 5117 84 5123 236
rect 5181 124 5187 236
rect 5517 164 5523 296
rect 5677 244 5683 256
rect 5725 244 5731 296
rect 5309 144 5315 156
rect 5421 144 5427 156
rect 5581 124 5587 236
rect 5629 124 5635 216
rect 5741 184 5747 356
rect 5789 324 5795 376
rect 5869 343 5875 496
rect 5933 464 5939 657
rect 5949 544 5955 636
rect 6013 584 6019 636
rect 5949 504 5955 516
rect 5965 484 5971 536
rect 6061 524 6067 536
rect 6077 524 6083 816
rect 6109 784 6115 796
rect 6173 784 6179 936
rect 6093 624 6099 736
rect 6109 704 6115 756
rect 6173 684 6179 756
rect 6189 724 6195 896
rect 6189 704 6195 716
rect 6109 583 6115 636
rect 6093 577 6115 583
rect 6093 503 6099 577
rect 6084 497 6099 503
rect 6109 503 6115 556
rect 6125 504 6131 656
rect 6141 624 6147 656
rect 6157 644 6163 676
rect 6109 497 6124 503
rect 5860 337 5875 343
rect 5789 284 5795 316
rect 5853 304 5859 336
rect 5869 284 5875 296
rect 5661 164 5667 176
rect 5741 144 5747 176
rect 5789 144 5795 156
rect 5885 144 5891 336
rect 5917 284 5923 456
rect 5997 324 6003 416
rect 6013 384 6019 476
rect 6029 344 6035 376
rect 6013 304 6019 336
rect 6061 324 6067 436
rect 6077 304 6083 336
rect 5901 264 5907 276
rect 6013 264 6019 296
rect 6093 284 6099 376
rect 6109 304 6115 497
rect 6125 424 6131 496
rect 6013 144 6019 236
rect 6077 224 6083 236
rect 6077 184 6083 196
rect 6141 164 6147 556
rect 6157 524 6163 636
rect 6157 444 6163 496
rect 6157 284 6163 436
rect 6173 324 6179 576
rect 6189 544 6195 676
rect 6205 643 6211 1016
rect 6221 964 6227 1237
rect 6237 943 6243 1216
rect 6253 944 6259 1156
rect 6269 1104 6275 1296
rect 6285 1284 6291 1316
rect 6333 1304 6339 1356
rect 6365 1303 6371 1456
rect 6381 1304 6387 1436
rect 6397 1384 6403 1496
rect 6413 1344 6419 1537
rect 6429 1484 6435 1496
rect 6445 1484 6451 1516
rect 6397 1337 6412 1343
rect 6349 1297 6371 1303
rect 6285 1224 6291 1236
rect 6301 1184 6307 1276
rect 6333 1244 6339 1296
rect 6317 1103 6323 1216
rect 6349 1164 6355 1297
rect 6397 1263 6403 1337
rect 6461 1263 6467 1636
rect 6477 1584 6483 1677
rect 6525 1663 6531 1676
rect 6509 1657 6531 1663
rect 6509 1584 6515 1657
rect 6541 1604 6547 1716
rect 6477 1464 6483 1536
rect 6493 1524 6499 1536
rect 6525 1524 6531 1536
rect 6557 1524 6563 1676
rect 6573 1523 6579 1956
rect 6589 1944 6595 2036
rect 6589 1764 6595 1836
rect 6589 1644 6595 1756
rect 6589 1544 6595 1576
rect 6573 1517 6595 1523
rect 6509 1484 6515 1496
rect 6573 1464 6579 1496
rect 6557 1324 6563 1336
rect 6397 1257 6419 1263
rect 6381 1144 6387 1236
rect 6397 1164 6403 1236
rect 6317 1097 6339 1103
rect 6285 1084 6291 1096
rect 6221 937 6243 943
rect 6221 884 6227 937
rect 6253 844 6259 896
rect 6237 824 6243 836
rect 6269 804 6275 1056
rect 6285 1044 6291 1076
rect 6317 923 6323 956
rect 6308 917 6323 923
rect 6333 863 6339 1097
rect 6349 1084 6355 1096
rect 6365 1044 6371 1136
rect 6397 1104 6403 1116
rect 6413 1104 6419 1257
rect 6445 1257 6467 1263
rect 6349 964 6355 1036
rect 6349 924 6355 936
rect 6317 857 6339 863
rect 6237 684 6243 696
rect 6253 684 6259 696
rect 6269 684 6275 776
rect 6237 644 6243 676
rect 6205 637 6227 643
rect 6189 364 6195 516
rect 6205 504 6211 536
rect 6221 484 6227 637
rect 6269 564 6275 636
rect 6301 564 6307 696
rect 6157 184 6163 256
rect 6093 124 6099 136
rect 6125 124 6131 136
rect 6173 124 6179 136
rect 6205 124 6211 236
rect 6237 144 6243 396
rect 6253 124 6259 476
rect 5149 84 5155 96
rect 4493 77 4508 83
rect 5533 83 5539 116
rect 5524 77 5539 83
rect 5709 83 5715 116
rect 5709 77 5724 83
rect 3261 24 3267 56
rect 3981 24 3987 36
rect 3053 17 3075 23
rect 1768 6 1774 14
rect 1782 6 1788 14
rect 1796 6 1802 14
rect 1810 6 1816 14
rect 2941 3 2947 16
rect 3053 3 3059 17
rect 2941 -3 3059 3
rect 4173 -17 4179 36
rect 4221 -17 4227 36
rect 4461 -17 4467 36
rect 4824 6 4830 14
rect 4838 6 4844 14
rect 4852 6 4858 14
rect 4866 6 4872 14
rect 5133 -17 5139 36
rect 5565 -17 5571 36
rect 5613 24 5619 36
rect 4173 -23 4195 -17
rect 4221 -23 4243 -17
rect 4461 -23 4483 -17
rect 5117 -23 5139 -17
rect 5549 -23 5571 -17
rect 5677 -17 5683 36
rect 6269 24 6275 536
rect 6301 304 6307 556
rect 6317 544 6323 857
rect 6333 744 6339 836
rect 6349 784 6355 876
rect 6333 664 6339 676
rect 6285 284 6291 296
rect 6301 284 6307 296
rect 6333 184 6339 536
rect 6349 344 6355 676
rect 6365 664 6371 1016
rect 6381 924 6387 1096
rect 6429 1083 6435 1176
rect 6445 1104 6451 1257
rect 6461 1224 6467 1236
rect 6429 1077 6444 1083
rect 6429 1063 6435 1077
rect 6413 1057 6435 1063
rect 6381 844 6387 876
rect 6397 764 6403 976
rect 6413 944 6419 1057
rect 6445 1044 6451 1056
rect 6429 924 6435 1036
rect 6445 963 6451 996
rect 6461 984 6467 1176
rect 6493 1123 6499 1316
rect 6573 1284 6579 1436
rect 6557 1184 6563 1236
rect 6573 1204 6579 1276
rect 6509 1124 6515 1136
rect 6477 1117 6499 1123
rect 6477 1004 6483 1117
rect 6445 957 6467 963
rect 6397 684 6403 756
rect 6397 644 6403 656
rect 6365 324 6371 596
rect 6285 103 6291 156
rect 6301 124 6307 156
rect 6285 97 6300 103
rect 6333 84 6339 136
rect 6349 104 6355 236
rect 5677 -23 5699 -17
rect 6253 -37 6259 16
rect 6285 -17 6291 56
rect 6317 24 6323 76
rect 6365 64 6371 236
rect 6381 43 6387 416
rect 6413 404 6419 916
rect 6445 704 6451 896
rect 6461 864 6467 957
rect 6493 923 6499 1096
rect 6525 1083 6531 1116
rect 6477 917 6499 923
rect 6509 1077 6531 1083
rect 6477 723 6483 917
rect 6493 824 6499 896
rect 6493 744 6499 756
rect 6477 717 6499 723
rect 6445 624 6451 676
rect 6461 644 6467 716
rect 6429 463 6435 576
rect 6445 544 6451 616
rect 6493 584 6499 717
rect 6509 584 6515 1077
rect 6541 1064 6547 1096
rect 6557 1084 6563 1136
rect 6573 1104 6579 1156
rect 6589 1104 6595 1517
rect 6525 924 6531 1036
rect 6541 963 6547 1036
rect 6541 957 6556 963
rect 6605 944 6611 2257
rect 6541 683 6547 836
rect 6557 724 6563 736
rect 6573 724 6579 916
rect 6532 677 6547 683
rect 6541 604 6547 636
rect 6429 457 6451 463
rect 6429 364 6435 436
rect 6397 304 6403 356
rect 6413 184 6419 276
rect 6397 124 6403 176
rect 6429 123 6435 336
rect 6445 144 6451 457
rect 6429 117 6444 123
rect 6477 104 6483 276
rect 6493 184 6499 496
rect 6372 37 6387 43
rect 6269 -23 6291 -17
rect 6301 -23 6307 16
rect 6317 -23 6339 -17
rect 6317 -37 6323 -23
rect 6253 -43 6323 -37
rect 6349 -37 6355 16
rect 6365 -23 6371 16
rect 6381 -37 6387 16
rect 6397 -23 6403 96
rect 6493 44 6499 156
rect 6509 144 6515 316
rect 6525 304 6531 476
rect 6541 364 6547 576
rect 6557 524 6563 696
rect 6589 684 6595 936
rect 6605 684 6611 716
rect 6621 704 6627 2636
rect 6637 1144 6643 2716
rect 6573 564 6579 636
rect 6605 384 6611 656
rect 6557 184 6563 216
rect 6605 184 6611 356
rect 6621 284 6627 436
rect 6637 264 6643 1076
rect 6717 544 6723 3196
rect 6621 204 6627 256
rect 6525 144 6531 156
rect 6461 -23 6467 36
rect 6493 -23 6499 16
rect 6541 -23 6547 16
rect 6573 -23 6579 76
rect 6605 -23 6611 56
rect 6637 -23 6643 36
rect 6349 -43 6387 -37
<< m3contact >>
rect 108 4736 116 4744
rect 620 4756 628 4764
rect 252 4736 260 4744
rect 380 4736 388 4744
rect 460 4736 468 4744
rect 508 4736 516 4744
rect 556 4736 564 4744
rect 636 4736 644 4744
rect 812 4736 820 4744
rect 828 4736 836 4744
rect 892 4736 900 4744
rect 908 4736 916 4744
rect 956 4736 964 4744
rect 428 4676 436 4684
rect 460 4676 468 4684
rect 492 4676 500 4684
rect 540 4676 548 4684
rect 620 4676 628 4684
rect 124 4656 132 4664
rect 252 4656 260 4664
rect 12 4576 20 4584
rect 12 4536 20 4544
rect 44 4536 52 4544
rect 92 4536 100 4544
rect 172 4616 180 4624
rect 188 4576 196 4584
rect 156 4556 164 4564
rect 76 4516 84 4524
rect 12 4496 20 4504
rect 60 4496 68 4504
rect 172 4496 180 4504
rect 12 4476 20 4484
rect 28 4476 36 4484
rect 12 4356 20 4364
rect 28 4296 36 4304
rect 44 4296 52 4304
rect 124 4316 132 4324
rect 76 4296 84 4304
rect 140 4296 148 4304
rect 172 4296 180 4304
rect 60 4276 68 4284
rect 92 4276 100 4284
rect 28 4256 36 4264
rect 44 4116 52 4124
rect 28 3936 36 3944
rect 108 4256 116 4264
rect 140 4256 148 4264
rect 220 4556 228 4564
rect 348 4656 356 4664
rect 332 4616 340 4624
rect 316 4576 324 4584
rect 268 4536 276 4544
rect 316 4536 324 4544
rect 204 4516 212 4524
rect 268 4516 276 4524
rect 332 4516 340 4524
rect 396 4656 404 4664
rect 524 4656 532 4664
rect 636 4656 644 4664
rect 668 4656 676 4664
rect 732 4676 740 4684
rect 732 4656 740 4664
rect 764 4656 772 4664
rect 620 4636 628 4644
rect 684 4636 692 4644
rect 700 4636 708 4644
rect 380 4556 388 4564
rect 444 4556 452 4564
rect 428 4536 436 4544
rect 476 4536 484 4544
rect 492 4536 500 4544
rect 300 4496 308 4504
rect 348 4496 356 4504
rect 636 4576 644 4584
rect 620 4556 628 4564
rect 860 4696 868 4704
rect 972 4696 980 4704
rect 828 4676 836 4684
rect 908 4676 916 4684
rect 956 4676 964 4684
rect 908 4656 916 4664
rect 940 4656 948 4664
rect 924 4636 932 4644
rect 956 4636 964 4644
rect 940 4556 948 4564
rect 636 4536 644 4544
rect 652 4536 660 4544
rect 796 4536 804 4544
rect 268 4476 276 4484
rect 380 4476 388 4484
rect 396 4476 404 4484
rect 220 4456 228 4464
rect 300 4456 308 4464
rect 252 4316 260 4324
rect 268 4316 276 4324
rect 380 4316 388 4324
rect 316 4296 324 4304
rect 396 4296 404 4304
rect 204 4256 212 4264
rect 300 4256 308 4264
rect 236 4236 244 4244
rect 284 4236 292 4244
rect 348 4236 356 4244
rect 188 4216 196 4224
rect 332 4196 340 4204
rect 316 4176 324 4184
rect 396 4156 404 4164
rect 428 4316 436 4324
rect 764 4516 772 4524
rect 972 4516 980 4524
rect 524 4496 532 4504
rect 572 4496 580 4504
rect 556 4476 564 4484
rect 572 4416 580 4424
rect 572 4336 580 4344
rect 508 4296 516 4304
rect 556 4296 564 4304
rect 668 4356 676 4364
rect 652 4296 660 4304
rect 588 4276 596 4284
rect 428 4216 436 4224
rect 572 4256 580 4264
rect 604 4256 612 4264
rect 492 4236 500 4244
rect 460 4216 468 4224
rect 444 4196 452 4204
rect 652 4236 660 4244
rect 652 4216 660 4224
rect 620 4176 628 4184
rect 556 4156 564 4164
rect 204 4136 212 4144
rect 348 4136 356 4144
rect 412 4136 420 4144
rect 540 4136 548 4144
rect 604 4136 612 4144
rect 108 4116 116 4124
rect 92 3896 100 3904
rect 764 4356 772 4364
rect 812 4356 820 4364
rect 748 4316 756 4324
rect 700 4296 708 4304
rect 716 4296 724 4304
rect 780 4336 788 4344
rect 812 4276 820 4284
rect 748 4256 756 4264
rect 684 4236 692 4244
rect 716 4236 724 4244
rect 668 4176 676 4184
rect 732 4176 740 4184
rect 764 4176 772 4184
rect 652 4156 660 4164
rect 572 4116 580 4124
rect 140 4076 148 4084
rect 156 3936 164 3944
rect 140 3916 148 3924
rect 204 3916 212 3924
rect 172 3876 180 3884
rect 204 3876 212 3884
rect 124 3856 132 3864
rect 12 3776 20 3784
rect 44 3776 52 3784
rect 236 3936 244 3944
rect 268 3916 276 3924
rect 252 3896 260 3904
rect 300 3896 308 3904
rect 364 3876 372 3884
rect 332 3856 340 3864
rect 412 3836 420 3844
rect 332 3816 340 3824
rect 268 3736 276 3744
rect 204 3716 212 3724
rect 172 3696 180 3704
rect 204 3696 212 3704
rect 268 3696 276 3704
rect 236 3536 244 3544
rect 76 3496 84 3504
rect 188 3436 196 3444
rect 220 3436 228 3444
rect 12 3336 20 3344
rect 124 3336 132 3344
rect 172 3336 180 3344
rect 572 3976 580 3984
rect 636 3976 644 3984
rect 524 3936 532 3944
rect 508 3916 516 3924
rect 540 3916 548 3924
rect 588 3936 596 3944
rect 620 3876 628 3884
rect 700 3836 708 3844
rect 476 3816 484 3824
rect 524 3816 532 3824
rect 476 3796 484 3804
rect 428 3736 436 3744
rect 348 3696 356 3704
rect 444 3696 452 3704
rect 412 3556 420 3564
rect 428 3516 436 3524
rect 268 3496 276 3504
rect 332 3496 340 3504
rect 428 3476 436 3484
rect 380 3436 388 3444
rect 412 3356 420 3364
rect 828 4256 836 4264
rect 924 4316 932 4324
rect 860 4296 868 4304
rect 908 4296 916 4304
rect 876 4256 884 4264
rect 908 4256 916 4264
rect 940 4256 948 4264
rect 1004 4636 1012 4644
rect 1020 4576 1028 4584
rect 1774 4806 1782 4814
rect 1788 4806 1796 4814
rect 1802 4806 1810 4814
rect 1740 4796 1748 4804
rect 1836 4796 1844 4804
rect 1068 4696 1076 4704
rect 1164 4696 1172 4704
rect 1180 4696 1188 4704
rect 1212 4696 1220 4704
rect 1100 4676 1108 4684
rect 1068 4656 1076 4664
rect 1164 4656 1172 4664
rect 1228 4656 1236 4664
rect 1116 4636 1124 4644
rect 1180 4636 1188 4644
rect 1324 4696 1332 4704
rect 1516 4716 1524 4724
rect 1388 4696 1396 4704
rect 1372 4680 1380 4684
rect 1372 4676 1380 4680
rect 1276 4656 1284 4664
rect 1260 4636 1268 4644
rect 1100 4596 1108 4604
rect 1084 4576 1092 4584
rect 1052 4556 1060 4564
rect 1036 4536 1044 4544
rect 1340 4656 1348 4664
rect 1308 4636 1316 4644
rect 1324 4636 1332 4644
rect 1244 4576 1252 4584
rect 1292 4576 1300 4584
rect 1148 4536 1156 4544
rect 1212 4536 1220 4544
rect 1132 4516 1140 4524
rect 1276 4516 1284 4524
rect 1100 4496 1108 4504
rect 1100 4476 1108 4484
rect 1020 4456 1028 4464
rect 1036 4376 1044 4384
rect 1004 4296 1012 4304
rect 1164 4336 1172 4344
rect 1084 4316 1092 4324
rect 1068 4296 1076 4304
rect 1132 4296 1140 4304
rect 1116 4276 1124 4284
rect 1228 4496 1236 4504
rect 1292 4496 1300 4504
rect 1212 4356 1220 4364
rect 1420 4676 1428 4684
rect 1452 4676 1460 4684
rect 1388 4636 1396 4644
rect 1404 4636 1412 4644
rect 1436 4636 1444 4644
rect 1404 4616 1412 4624
rect 1532 4676 1540 4684
rect 1484 4636 1492 4644
rect 1500 4636 1508 4644
rect 1372 4576 1380 4584
rect 1404 4576 1412 4584
rect 1468 4576 1476 4584
rect 1500 4576 1508 4584
rect 1452 4556 1460 4564
rect 1468 4556 1476 4564
rect 1516 4556 1524 4564
rect 1612 4716 1620 4724
rect 1628 4716 1636 4724
rect 2220 4776 2228 4784
rect 1868 4716 1876 4724
rect 1916 4716 1924 4724
rect 1980 4716 1988 4724
rect 2028 4716 2036 4724
rect 2092 4716 2100 4724
rect 2188 4716 2196 4724
rect 1836 4676 1844 4684
rect 1932 4676 1940 4684
rect 1996 4676 2004 4684
rect 1596 4656 1604 4664
rect 1692 4656 1700 4664
rect 1740 4656 1748 4664
rect 1772 4656 1780 4664
rect 1884 4656 1892 4664
rect 1580 4636 1588 4644
rect 1564 4596 1572 4604
rect 1724 4596 1732 4604
rect 1548 4576 1556 4584
rect 1676 4576 1684 4584
rect 1340 4536 1348 4544
rect 1452 4536 1460 4544
rect 1532 4536 1540 4544
rect 1276 4456 1284 4464
rect 1308 4456 1316 4464
rect 1244 4356 1252 4364
rect 1244 4336 1252 4344
rect 1372 4516 1380 4524
rect 1500 4516 1508 4524
rect 1420 4496 1428 4504
rect 1484 4496 1492 4504
rect 1340 4476 1348 4484
rect 1324 4416 1332 4424
rect 1308 4316 1316 4324
rect 1228 4296 1236 4304
rect 1244 4296 1252 4304
rect 1276 4296 1284 4304
rect 1388 4296 1396 4304
rect 1452 4296 1460 4304
rect 988 4256 996 4264
rect 1020 4256 1028 4264
rect 1036 4256 1044 4264
rect 1068 4256 1076 4264
rect 1132 4236 1140 4244
rect 860 4196 868 4204
rect 908 4196 916 4204
rect 956 4196 964 4204
rect 780 3976 788 3984
rect 764 3916 772 3924
rect 876 4156 884 4164
rect 1116 4176 1124 4184
rect 1100 4156 1108 4164
rect 1004 4136 1012 4144
rect 860 4096 868 4104
rect 860 3936 868 3944
rect 844 3916 852 3924
rect 876 3916 884 3924
rect 956 3916 964 3924
rect 860 3896 868 3904
rect 876 3896 884 3904
rect 940 3902 948 3904
rect 940 3896 948 3902
rect 716 3816 724 3824
rect 620 3796 628 3804
rect 556 3776 564 3784
rect 892 3836 900 3844
rect 908 3836 916 3844
rect 1116 4096 1124 4104
rect 1148 4176 1156 4184
rect 1164 4136 1172 4144
rect 1324 4196 1332 4204
rect 1276 4156 1284 4164
rect 1372 4276 1380 4284
rect 1420 4216 1428 4224
rect 1356 4196 1364 4204
rect 1340 4136 1348 4144
rect 1180 4096 1188 4104
rect 1260 4096 1268 4104
rect 1132 4076 1140 4084
rect 1180 3976 1188 3984
rect 1132 3956 1140 3964
rect 1052 3916 1060 3924
rect 1100 3916 1108 3924
rect 1148 3916 1156 3924
rect 1004 3836 1012 3844
rect 1004 3796 1012 3804
rect 652 3756 660 3764
rect 764 3756 772 3764
rect 828 3756 836 3764
rect 956 3756 964 3764
rect 732 3736 740 3744
rect 508 3696 516 3704
rect 572 3696 580 3704
rect 508 3556 516 3564
rect 524 3536 532 3544
rect 524 3516 532 3524
rect 716 3716 724 3724
rect 684 3696 692 3704
rect 1100 3896 1108 3904
rect 1132 3896 1140 3904
rect 1084 3876 1092 3884
rect 1068 3836 1076 3844
rect 1084 3756 1092 3764
rect 1052 3736 1060 3744
rect 876 3716 884 3724
rect 956 3716 964 3724
rect 684 3576 692 3584
rect 716 3576 724 3584
rect 748 3576 756 3584
rect 604 3496 612 3504
rect 540 3396 548 3404
rect 540 3356 548 3364
rect 556 3356 564 3364
rect 476 3336 484 3344
rect 524 3336 532 3344
rect 588 3336 596 3344
rect 684 3496 692 3504
rect 620 3476 628 3484
rect 652 3476 660 3484
rect 636 3436 644 3444
rect 652 3416 660 3424
rect 380 3316 388 3324
rect 460 3316 468 3324
rect 524 3316 532 3324
rect 636 3316 644 3324
rect 460 3296 468 3304
rect 572 3296 580 3304
rect 188 3176 196 3184
rect 572 3176 580 3184
rect 748 3556 756 3564
rect 780 3536 788 3544
rect 764 3356 772 3364
rect 844 3516 852 3524
rect 876 3516 884 3524
rect 796 3476 804 3484
rect 924 3476 932 3484
rect 812 3436 820 3444
rect 876 3456 884 3464
rect 940 3456 948 3464
rect 876 3436 884 3444
rect 844 3396 852 3404
rect 844 3376 852 3384
rect 748 3336 756 3344
rect 652 3296 660 3304
rect 700 3296 708 3304
rect 668 3156 676 3164
rect 956 3436 964 3444
rect 892 3416 900 3424
rect 940 3416 948 3424
rect 924 3396 932 3404
rect 908 3376 916 3384
rect 956 3356 964 3364
rect 1020 3576 1028 3584
rect 1020 3516 1028 3524
rect 1052 3576 1060 3584
rect 1196 3936 1204 3944
rect 1212 3816 1220 3824
rect 1308 4056 1316 4064
rect 1276 3956 1284 3964
rect 1260 3916 1268 3924
rect 1244 3796 1252 3804
rect 1148 3776 1156 3784
rect 1164 3756 1172 3764
rect 1260 3736 1268 3744
rect 1484 4136 1492 4144
rect 1324 3976 1332 3984
rect 1340 3896 1348 3904
rect 1324 3796 1332 3804
rect 1468 3936 1476 3944
rect 1404 3856 1412 3864
rect 1420 3776 1428 3784
rect 1356 3756 1364 3764
rect 1324 3716 1332 3724
rect 1356 3716 1364 3724
rect 1116 3536 1124 3544
rect 1100 3516 1108 3524
rect 1036 3496 1044 3504
rect 1068 3496 1076 3504
rect 1132 3496 1140 3504
rect 1180 3496 1188 3504
rect 988 3476 996 3484
rect 1004 3476 1012 3484
rect 1164 3476 1172 3484
rect 1052 3456 1060 3464
rect 1228 3456 1236 3464
rect 1196 3396 1204 3404
rect 1212 3396 1220 3404
rect 1020 3376 1028 3384
rect 1068 3376 1076 3384
rect 1660 4536 1668 4544
rect 1676 4536 1684 4544
rect 1724 4536 1732 4544
rect 2172 4656 2180 4664
rect 2060 4636 2068 4644
rect 2156 4636 2164 4644
rect 1836 4576 1844 4584
rect 2060 4576 2068 4584
rect 2108 4576 2116 4584
rect 2156 4576 2164 4584
rect 1820 4556 1828 4564
rect 1852 4556 1860 4564
rect 1884 4556 1892 4564
rect 2508 4796 2516 4804
rect 2332 4776 2340 4784
rect 2364 4776 2372 4784
rect 2236 4716 2244 4724
rect 2428 4716 2436 4724
rect 2476 4716 2484 4724
rect 2220 4656 2228 4664
rect 2284 4656 2292 4664
rect 2316 4656 2324 4664
rect 2364 4656 2372 4664
rect 2252 4636 2260 4644
rect 2108 4556 2116 4564
rect 2140 4556 2148 4564
rect 2204 4556 2212 4564
rect 2300 4556 2308 4564
rect 1900 4536 1908 4544
rect 1948 4536 1956 4544
rect 2044 4536 2052 4544
rect 2108 4536 2116 4544
rect 2188 4536 2196 4544
rect 2220 4536 2228 4544
rect 2236 4536 2244 4544
rect 2284 4536 2292 4544
rect 1564 4516 1572 4524
rect 1628 4516 1636 4524
rect 1708 4516 1716 4524
rect 1756 4516 1764 4524
rect 1564 4496 1572 4504
rect 1596 4496 1604 4504
rect 1676 4496 1684 4504
rect 1692 4476 1700 4484
rect 1756 4476 1764 4484
rect 1774 4406 1782 4414
rect 1788 4406 1796 4414
rect 1802 4406 1810 4414
rect 1724 4376 1732 4384
rect 1740 4376 1748 4384
rect 1852 4376 1860 4384
rect 1596 4316 1604 4324
rect 1660 4316 1668 4324
rect 1708 4316 1716 4324
rect 1580 4296 1588 4304
rect 1548 4276 1556 4284
rect 1692 4276 1700 4284
rect 1612 4156 1620 4164
rect 1596 4116 1604 4124
rect 1548 3916 1556 3924
rect 1532 3896 1540 3904
rect 1660 4156 1668 4164
rect 1676 4116 1684 4124
rect 1772 4316 1780 4324
rect 1836 4256 1844 4264
rect 1756 4136 1764 4144
rect 1868 4216 1876 4224
rect 2364 4556 2372 4564
rect 2412 4576 2420 4584
rect 2444 4556 2452 4564
rect 2380 4536 2388 4544
rect 1964 4516 1972 4524
rect 2092 4516 2100 4524
rect 2140 4516 2148 4524
rect 1980 4336 1988 4344
rect 2044 4356 2052 4364
rect 2028 4316 2036 4324
rect 2076 4316 2084 4324
rect 1916 4276 1924 4284
rect 1884 4156 1892 4164
rect 2092 4276 2100 4284
rect 2108 4276 2116 4284
rect 1996 4256 2004 4264
rect 1964 4236 1972 4244
rect 2028 4236 2036 4244
rect 2012 4156 2020 4164
rect 1868 4136 1876 4144
rect 1900 4136 1908 4144
rect 2028 4136 2036 4144
rect 2060 4136 2068 4144
rect 2076 4136 2084 4144
rect 1628 4056 1636 4064
rect 1612 4036 1620 4044
rect 1820 4036 1828 4044
rect 1612 3936 1620 3944
rect 1596 3916 1604 3924
rect 1628 3916 1636 3924
rect 1774 4006 1782 4014
rect 1788 4006 1796 4014
rect 1802 4006 1810 4014
rect 1660 3896 1668 3904
rect 1692 3896 1700 3904
rect 1804 3896 1812 3904
rect 1484 3776 1492 3784
rect 1532 3876 1540 3884
rect 1564 3876 1572 3884
rect 2188 4496 2196 4504
rect 2268 4496 2276 4504
rect 2220 4476 2228 4484
rect 2332 4476 2340 4484
rect 2268 4356 2276 4364
rect 2188 4336 2196 4344
rect 2252 4336 2260 4344
rect 2156 4316 2164 4324
rect 2204 4276 2212 4284
rect 2188 4256 2196 4264
rect 2220 4256 2228 4264
rect 2124 4196 2132 4204
rect 2236 4216 2244 4224
rect 2252 4196 2260 4204
rect 2156 4156 2164 4164
rect 2124 4136 2132 4144
rect 2140 4116 2148 4124
rect 2236 4116 2244 4124
rect 1916 4096 1924 4104
rect 2060 4096 2068 4104
rect 2076 4096 2084 4104
rect 2220 4096 2228 4104
rect 2332 4356 2340 4364
rect 2732 4796 2740 4804
rect 2540 4716 2548 4724
rect 2556 4716 2564 4724
rect 2604 4716 2612 4724
rect 2508 4656 2516 4664
rect 2588 4656 2596 4664
rect 2652 4656 2660 4664
rect 2556 4576 2564 4584
rect 2492 4556 2500 4564
rect 2636 4576 2644 4584
rect 2684 4716 2692 4724
rect 2860 4676 2868 4684
rect 2812 4616 2820 4624
rect 2860 4616 2868 4624
rect 2652 4556 2660 4564
rect 2668 4556 2676 4564
rect 2684 4556 2692 4564
rect 2764 4556 2772 4564
rect 2796 4556 2804 4564
rect 2812 4556 2820 4564
rect 2492 4536 2500 4544
rect 2524 4536 2532 4544
rect 2620 4536 2628 4544
rect 2428 4516 2436 4524
rect 2476 4516 2484 4524
rect 2396 4316 2404 4324
rect 2524 4516 2532 4524
rect 2620 4516 2628 4524
rect 2700 4516 2708 4524
rect 2556 4496 2564 4504
rect 2652 4496 2660 4504
rect 2492 4456 2500 4464
rect 2572 4416 2580 4424
rect 2508 4356 2516 4364
rect 2460 4336 2468 4344
rect 2540 4316 2548 4324
rect 2492 4296 2500 4304
rect 2524 4296 2532 4304
rect 2428 4236 2436 4244
rect 2300 4216 2308 4224
rect 2332 4156 2340 4164
rect 2300 4136 2308 4144
rect 2364 4136 2372 4144
rect 2268 4116 2276 4124
rect 2364 4096 2372 4104
rect 2348 4076 2356 4084
rect 2380 4076 2388 4084
rect 2060 4056 2068 4064
rect 2332 4056 2340 4064
rect 1916 3936 1924 3944
rect 2028 3936 2036 3944
rect 1964 3896 1972 3904
rect 1676 3876 1684 3884
rect 1836 3876 1844 3884
rect 1580 3856 1588 3864
rect 1628 3856 1636 3864
rect 1676 3856 1684 3864
rect 1564 3836 1572 3844
rect 1660 3836 1668 3844
rect 1660 3776 1668 3784
rect 1692 3776 1700 3784
rect 1740 3776 1748 3784
rect 1500 3716 1508 3724
rect 1452 3696 1460 3704
rect 1404 3676 1412 3684
rect 1436 3676 1444 3684
rect 1596 3676 1604 3684
rect 1452 3616 1460 3624
rect 1484 3616 1492 3624
rect 1740 3696 1748 3704
rect 1772 3696 1780 3704
rect 1836 3696 1844 3704
rect 1996 3836 2004 3844
rect 2044 3816 2052 3824
rect 1932 3796 1940 3804
rect 2108 4036 2116 4044
rect 2092 4016 2100 4024
rect 2108 3896 2116 3904
rect 2220 3836 2228 3844
rect 2028 3736 2036 3744
rect 1964 3718 1972 3724
rect 1964 3716 1972 3718
rect 1868 3696 1876 3704
rect 1852 3676 1860 3684
rect 1774 3606 1782 3614
rect 1788 3606 1796 3614
rect 1802 3606 1810 3614
rect 1612 3476 1620 3484
rect 1660 3476 1668 3484
rect 1708 3476 1716 3484
rect 1516 3456 1524 3464
rect 1692 3456 1700 3464
rect 1724 3456 1732 3464
rect 1276 3416 1284 3424
rect 1372 3416 1380 3424
rect 1260 3376 1268 3384
rect 1244 3356 1252 3364
rect 1308 3356 1316 3364
rect 1036 3336 1044 3344
rect 1132 3336 1140 3344
rect 1196 3336 1204 3344
rect 796 3316 804 3324
rect 892 3316 900 3324
rect 988 3316 996 3324
rect 924 3296 932 3304
rect 972 3296 980 3304
rect 1036 3296 1044 3304
rect 780 3276 788 3284
rect 828 3276 836 3284
rect 924 3196 932 3204
rect 812 3156 820 3164
rect 764 3136 772 3144
rect 1212 3216 1220 3224
rect 860 3116 868 3124
rect 1100 3116 1108 3124
rect 300 3096 308 3104
rect 364 3102 372 3104
rect 364 3096 372 3102
rect 732 3096 740 3104
rect 796 3102 804 3104
rect 796 3096 804 3102
rect 60 2956 68 2964
rect 44 2936 52 2944
rect 44 2916 52 2924
rect 28 2876 36 2884
rect 44 2816 52 2824
rect 124 3076 132 3084
rect 332 3076 340 3084
rect 92 3016 100 3024
rect 492 3036 500 3044
rect 300 3016 308 3024
rect 540 3056 548 3064
rect 604 3056 612 3064
rect 588 3016 596 3024
rect 620 3016 628 3024
rect 508 2996 516 3004
rect 540 2996 548 3004
rect 700 3056 708 3064
rect 732 3056 740 3064
rect 796 3056 804 3064
rect 684 2996 692 3004
rect 636 2956 644 2964
rect 716 2956 724 2964
rect 844 2956 852 2964
rect 108 2936 116 2944
rect 172 2936 180 2944
rect 204 2936 212 2944
rect 316 2936 324 2944
rect 172 2916 180 2924
rect 268 2916 276 2924
rect 188 2896 196 2904
rect 252 2896 260 2904
rect 156 2876 164 2884
rect 188 2876 196 2884
rect 252 2876 260 2884
rect 124 2836 132 2844
rect 188 2836 196 2844
rect 236 2836 244 2844
rect 92 2736 100 2744
rect 172 2736 180 2744
rect 428 2936 436 2944
rect 492 2936 500 2944
rect 524 2936 532 2944
rect 700 2936 708 2944
rect 748 2936 756 2944
rect 332 2916 340 2924
rect 380 2916 388 2924
rect 380 2896 388 2904
rect 284 2876 292 2884
rect 316 2876 324 2884
rect 348 2876 356 2884
rect 268 2796 276 2804
rect 300 2796 308 2804
rect 252 2716 260 2724
rect 188 2696 196 2704
rect 220 2696 228 2704
rect 172 2656 180 2664
rect 76 2636 84 2644
rect 12 2536 20 2544
rect 108 2536 116 2544
rect 124 2536 132 2544
rect 108 2496 116 2504
rect 252 2656 260 2664
rect 220 2556 228 2564
rect 268 2556 276 2564
rect 284 2556 292 2564
rect 332 2836 340 2844
rect 428 2916 436 2924
rect 444 2916 452 2924
rect 524 2916 532 2924
rect 540 2916 548 2924
rect 588 2916 596 2924
rect 604 2916 612 2924
rect 652 2916 660 2924
rect 412 2836 420 2844
rect 364 2716 372 2724
rect 396 2716 404 2724
rect 444 2876 452 2884
rect 492 2796 500 2804
rect 812 2936 820 2944
rect 764 2896 772 2904
rect 780 2896 788 2904
rect 684 2876 692 2884
rect 716 2876 724 2884
rect 732 2876 740 2884
rect 828 2876 836 2884
rect 636 2836 644 2844
rect 668 2836 676 2844
rect 540 2796 548 2804
rect 700 2816 708 2824
rect 588 2736 596 2744
rect 620 2736 628 2744
rect 524 2716 532 2724
rect 972 3056 980 3064
rect 940 2936 948 2944
rect 1052 3096 1060 3104
rect 1100 3096 1108 3104
rect 1148 3096 1156 3104
rect 1036 3076 1044 3084
rect 988 2976 996 2984
rect 1004 2956 1012 2964
rect 940 2916 948 2924
rect 972 2916 980 2924
rect 908 2836 916 2844
rect 924 2836 932 2844
rect 924 2796 932 2804
rect 844 2736 852 2744
rect 492 2696 500 2704
rect 428 2676 436 2684
rect 476 2676 484 2684
rect 524 2676 532 2684
rect 540 2656 548 2664
rect 332 2636 340 2644
rect 316 2556 324 2564
rect 236 2536 244 2544
rect 284 2536 292 2544
rect 188 2516 196 2524
rect 236 2516 244 2524
rect 204 2496 212 2504
rect 140 2476 148 2484
rect 44 2456 52 2464
rect 140 2456 148 2464
rect 12 2316 20 2324
rect 44 2296 52 2304
rect 124 2336 132 2344
rect 108 2196 116 2204
rect 108 2176 116 2184
rect 60 2156 68 2164
rect 124 2156 132 2164
rect 44 2116 52 2124
rect 188 2356 196 2364
rect 188 2336 196 2344
rect 172 2316 180 2324
rect 172 2296 180 2304
rect 156 2256 164 2264
rect 188 2176 196 2184
rect 156 2136 164 2144
rect 92 2116 100 2124
rect 188 2116 196 2124
rect 28 2096 36 2104
rect 76 2096 84 2104
rect 44 2076 52 2084
rect 108 2096 116 2104
rect 92 1996 100 2004
rect 140 2076 148 2084
rect 156 1996 164 2004
rect 124 1956 132 1964
rect 12 1936 20 1944
rect 44 1916 52 1924
rect 92 1916 100 1924
rect 172 1916 180 1924
rect 28 1896 36 1904
rect 12 1756 20 1764
rect 44 1756 52 1764
rect 108 1896 116 1904
rect 156 1896 164 1904
rect 572 2596 580 2604
rect 620 2676 628 2684
rect 796 2696 804 2704
rect 860 2696 868 2704
rect 716 2676 724 2684
rect 732 2676 740 2684
rect 764 2676 772 2684
rect 668 2656 676 2664
rect 684 2656 692 2664
rect 716 2636 724 2644
rect 812 2656 820 2664
rect 780 2636 788 2644
rect 956 2876 964 2884
rect 1020 2876 1028 2884
rect 972 2776 980 2784
rect 1404 3396 1412 3404
rect 1356 3296 1364 3304
rect 1468 3376 1476 3384
rect 1628 3416 1636 3424
rect 1644 3416 1652 3424
rect 1532 3376 1540 3384
rect 1516 3336 1524 3344
rect 1436 3316 1444 3324
rect 1484 3316 1492 3324
rect 1500 3316 1508 3324
rect 1452 3296 1460 3304
rect 1500 3296 1508 3304
rect 1388 3276 1396 3284
rect 1484 3256 1492 3264
rect 1372 3216 1380 3224
rect 1388 3216 1396 3224
rect 1388 3176 1396 3184
rect 1404 3176 1412 3184
rect 1372 3156 1380 3164
rect 1292 3116 1300 3124
rect 1324 3116 1332 3124
rect 1388 3116 1396 3124
rect 1484 3116 1492 3124
rect 1260 3096 1268 3104
rect 1132 3076 1140 3084
rect 1244 3076 1252 3084
rect 1068 3056 1076 3064
rect 1340 3096 1348 3104
rect 1436 3096 1444 3104
rect 1564 3356 1572 3364
rect 1596 3356 1604 3364
rect 1612 3336 1620 3344
rect 1644 3336 1652 3344
rect 1548 3296 1556 3304
rect 1660 3296 1668 3304
rect 1516 3276 1524 3284
rect 1676 3256 1684 3264
rect 1564 3176 1572 3184
rect 1548 3156 1556 3164
rect 1292 3076 1300 3084
rect 1356 3076 1364 3084
rect 1404 3076 1412 3084
rect 1468 3076 1476 3084
rect 1516 3076 1524 3084
rect 1532 3076 1540 3084
rect 1084 3016 1092 3024
rect 1116 2916 1124 2924
rect 1068 2836 1076 2844
rect 1116 2816 1124 2824
rect 1116 2796 1124 2804
rect 1036 2756 1044 2764
rect 1052 2756 1060 2764
rect 1116 2756 1124 2764
rect 1164 3016 1172 3024
rect 1228 2976 1236 2984
rect 1340 2976 1348 2984
rect 1260 2956 1268 2964
rect 1212 2936 1220 2944
rect 1260 2936 1268 2944
rect 1196 2916 1204 2924
rect 1260 2896 1268 2904
rect 1180 2716 1188 2724
rect 1068 2696 1076 2704
rect 1132 2696 1140 2704
rect 1020 2676 1028 2684
rect 1084 2676 1092 2684
rect 1116 2676 1124 2684
rect 636 2596 644 2604
rect 668 2596 676 2604
rect 876 2616 884 2624
rect 988 2656 996 2664
rect 1036 2656 1044 2664
rect 1100 2656 1108 2664
rect 1052 2636 1060 2644
rect 1004 2616 1012 2624
rect 812 2576 820 2584
rect 892 2576 900 2584
rect 444 2556 452 2564
rect 428 2536 436 2544
rect 476 2536 484 2544
rect 524 2536 532 2544
rect 540 2536 548 2544
rect 652 2536 660 2544
rect 684 2536 692 2544
rect 732 2536 740 2544
rect 364 2516 372 2524
rect 492 2516 500 2524
rect 252 2456 260 2464
rect 300 2456 308 2464
rect 332 2456 340 2464
rect 364 2456 372 2464
rect 300 2436 308 2444
rect 268 2356 276 2364
rect 524 2496 532 2504
rect 604 2496 612 2504
rect 732 2516 740 2524
rect 428 2476 436 2484
rect 588 2476 596 2484
rect 412 2356 420 2364
rect 236 2336 244 2344
rect 252 2296 260 2304
rect 252 2136 260 2144
rect 220 2116 228 2124
rect 284 2316 292 2324
rect 300 2276 308 2284
rect 444 2336 452 2344
rect 460 2336 468 2344
rect 492 2336 500 2344
rect 604 2356 612 2364
rect 524 2296 532 2304
rect 364 2276 372 2284
rect 348 2256 356 2264
rect 412 2236 420 2244
rect 460 2236 468 2244
rect 364 2176 372 2184
rect 332 2136 340 2144
rect 284 2116 292 2124
rect 380 2116 388 2124
rect 204 2096 212 2104
rect 332 2096 340 2104
rect 364 2096 372 2104
rect 396 2096 404 2104
rect 236 2076 244 2084
rect 268 2076 276 2084
rect 300 2076 308 2084
rect 348 2076 356 2084
rect 204 1936 212 1944
rect 364 1936 372 1944
rect 236 1916 244 1924
rect 108 1756 116 1764
rect 124 1736 132 1744
rect 44 1676 52 1684
rect 92 1676 100 1684
rect 92 1536 100 1544
rect 60 1516 68 1524
rect 76 1516 84 1524
rect 44 1496 52 1504
rect 28 1456 36 1464
rect 140 1716 148 1724
rect 220 1896 228 1904
rect 188 1736 196 1744
rect 172 1696 180 1704
rect 220 1696 228 1704
rect 188 1676 196 1684
rect 220 1636 228 1644
rect 204 1556 212 1564
rect 156 1536 164 1544
rect 268 1856 276 1864
rect 252 1796 260 1804
rect 268 1696 276 1704
rect 332 1916 340 1924
rect 476 2116 484 2124
rect 460 2096 468 2104
rect 444 1996 452 2004
rect 300 1896 308 1904
rect 348 1896 356 1904
rect 396 1896 404 1904
rect 428 1896 436 1904
rect 364 1876 372 1884
rect 428 1876 436 1884
rect 348 1796 356 1804
rect 444 1856 452 1864
rect 380 1756 388 1764
rect 428 1756 436 1764
rect 396 1716 404 1724
rect 316 1696 324 1704
rect 348 1696 356 1704
rect 380 1676 388 1684
rect 444 1676 452 1684
rect 252 1636 260 1644
rect 284 1636 292 1644
rect 252 1556 260 1564
rect 300 1536 308 1544
rect 140 1496 148 1504
rect 188 1496 196 1504
rect 156 1476 164 1484
rect 124 1456 132 1464
rect 284 1516 292 1524
rect 332 1516 340 1524
rect 268 1496 276 1504
rect 60 1356 68 1364
rect 124 1356 132 1364
rect 204 1356 212 1364
rect 44 1336 52 1344
rect 44 1316 52 1324
rect 140 1336 148 1344
rect 92 1316 100 1324
rect 44 1296 52 1304
rect 28 1276 36 1284
rect 76 1276 84 1284
rect 76 1176 84 1184
rect 28 1136 36 1144
rect 28 1116 36 1124
rect 44 1076 52 1084
rect 12 1036 20 1044
rect 76 1096 84 1104
rect 188 1296 196 1304
rect 172 1136 180 1144
rect 236 1336 244 1344
rect 252 1316 260 1324
rect 236 1156 244 1164
rect 236 1136 244 1144
rect 140 1096 148 1104
rect 156 1096 164 1104
rect 220 1096 228 1104
rect 92 1076 100 1084
rect 124 1076 132 1084
rect 172 1056 180 1064
rect 108 996 116 1004
rect 76 976 84 984
rect 28 956 36 964
rect 268 1276 276 1284
rect 444 1536 452 1544
rect 428 1496 436 1504
rect 316 1456 324 1464
rect 348 1456 356 1464
rect 396 1456 404 1464
rect 604 2276 612 2284
rect 508 2236 516 2244
rect 572 2236 580 2244
rect 636 2236 644 2244
rect 684 2476 692 2484
rect 828 2556 836 2564
rect 860 2556 868 2564
rect 1004 2556 1012 2564
rect 1036 2556 1044 2564
rect 844 2536 852 2544
rect 972 2536 980 2544
rect 1196 2656 1204 2664
rect 1324 2776 1332 2784
rect 1260 2756 1268 2764
rect 1292 2736 1300 2744
rect 1244 2716 1252 2724
rect 1228 2676 1236 2684
rect 1212 2636 1220 2644
rect 1180 2616 1188 2624
rect 1212 2616 1220 2624
rect 1276 2616 1284 2624
rect 1356 2896 1364 2904
rect 1548 2956 1556 2964
rect 1420 2916 1428 2924
rect 1388 2876 1396 2884
rect 1516 2916 1524 2924
rect 1500 2856 1508 2864
rect 1452 2836 1460 2844
rect 1612 3156 1620 3164
rect 1676 3136 1684 3144
rect 1628 3096 1636 3104
rect 1612 2956 1620 2964
rect 1708 3436 1716 3444
rect 2124 3736 2132 3744
rect 2076 3696 2084 3704
rect 2108 3696 2116 3704
rect 1996 3676 2004 3684
rect 1884 3576 1892 3584
rect 1836 3456 1844 3464
rect 1820 3436 1828 3444
rect 1868 3396 1876 3404
rect 1852 3376 1860 3384
rect 1868 3376 1876 3384
rect 1740 3356 1748 3364
rect 1772 3316 1780 3324
rect 1804 3316 1812 3324
rect 1852 3316 1860 3324
rect 1724 3296 1732 3304
rect 1820 3296 1828 3304
rect 1774 3206 1782 3214
rect 1788 3206 1796 3214
rect 1802 3206 1810 3214
rect 1836 3136 1844 3144
rect 1708 3116 1716 3124
rect 1756 3116 1764 3124
rect 1740 3096 1748 3104
rect 1724 3076 1732 3084
rect 1772 3056 1780 3064
rect 1580 2936 1588 2944
rect 1580 2916 1588 2924
rect 1612 2876 1620 2884
rect 1692 2876 1700 2884
rect 1676 2836 1684 2844
rect 1660 2776 1668 2784
rect 1564 2736 1572 2744
rect 1356 2696 1364 2704
rect 1388 2696 1396 2704
rect 1564 2696 1572 2704
rect 1628 2702 1636 2704
rect 1628 2696 1636 2702
rect 1324 2676 1332 2684
rect 1372 2676 1380 2684
rect 1484 2676 1492 2684
rect 1324 2636 1332 2644
rect 1500 2656 1508 2664
rect 1436 2636 1444 2644
rect 1532 2636 1540 2644
rect 1404 2576 1412 2584
rect 988 2516 996 2524
rect 1052 2516 1060 2524
rect 1084 2516 1092 2524
rect 796 2436 804 2444
rect 844 2436 852 2444
rect 956 2436 964 2444
rect 700 2316 708 2324
rect 764 2276 772 2284
rect 716 2256 724 2264
rect 668 2236 676 2244
rect 732 2236 740 2244
rect 588 2196 596 2204
rect 652 2196 660 2204
rect 572 2136 580 2144
rect 524 2116 532 2124
rect 556 2116 564 2124
rect 492 2076 500 2084
rect 524 1996 532 2004
rect 492 1916 500 1924
rect 572 2096 580 2104
rect 636 2136 644 2144
rect 700 2136 708 2144
rect 604 2116 612 2124
rect 604 2096 612 2104
rect 652 2096 660 2104
rect 492 1896 500 1904
rect 540 1896 548 1904
rect 492 1876 500 1884
rect 556 1876 564 1884
rect 508 1856 516 1864
rect 508 1756 516 1764
rect 556 1736 564 1744
rect 492 1716 500 1724
rect 524 1716 532 1724
rect 508 1696 516 1704
rect 476 1676 484 1684
rect 508 1656 516 1664
rect 540 1676 548 1684
rect 476 1516 484 1524
rect 508 1516 516 1524
rect 524 1516 532 1524
rect 748 2116 756 2124
rect 924 2316 932 2324
rect 972 2316 980 2324
rect 892 2276 900 2284
rect 940 2276 948 2284
rect 828 2236 836 2244
rect 860 2236 868 2244
rect 812 2216 820 2224
rect 956 2256 964 2264
rect 908 2236 916 2244
rect 956 2236 964 2244
rect 876 2216 884 2224
rect 828 2116 836 2124
rect 588 2076 596 2084
rect 684 2076 692 2084
rect 716 2076 724 2084
rect 812 2096 820 2104
rect 668 1996 676 2004
rect 716 1996 724 2004
rect 668 1976 676 1984
rect 700 1916 708 1924
rect 588 1896 596 1904
rect 636 1896 644 1904
rect 668 1896 676 1904
rect 780 1916 788 1924
rect 812 1916 820 1924
rect 828 1916 836 1924
rect 700 1876 708 1884
rect 572 1696 580 1704
rect 732 1856 740 1864
rect 748 1856 756 1864
rect 892 2116 900 2124
rect 924 2116 932 2124
rect 1036 2316 1044 2324
rect 1068 2316 1076 2324
rect 1004 2236 1012 2244
rect 1004 2216 1012 2224
rect 1052 2256 1060 2264
rect 1068 2216 1076 2224
rect 1020 2196 1028 2204
rect 1068 2196 1076 2204
rect 988 2156 996 2164
rect 1020 2156 1028 2164
rect 988 2136 996 2144
rect 972 2096 980 2104
rect 1164 2556 1172 2564
rect 1180 2556 1188 2564
rect 1276 2556 1284 2564
rect 1340 2556 1348 2564
rect 1116 2536 1124 2544
rect 1132 2516 1140 2524
rect 1148 2516 1156 2524
rect 1324 2536 1332 2544
rect 1292 2516 1300 2524
rect 1196 2496 1204 2504
rect 1116 2296 1124 2304
rect 1164 2276 1172 2284
rect 1132 2216 1140 2224
rect 1100 2136 1108 2144
rect 1036 2096 1044 2104
rect 1020 2016 1028 2024
rect 876 1956 884 1964
rect 956 1956 964 1964
rect 956 1916 964 1924
rect 1004 1916 1012 1924
rect 1068 1916 1076 1924
rect 1116 1916 1124 1924
rect 876 1896 884 1904
rect 988 1896 996 1904
rect 1052 1896 1060 1904
rect 860 1876 868 1884
rect 908 1876 916 1884
rect 940 1876 948 1884
rect 844 1856 852 1864
rect 796 1836 804 1844
rect 828 1836 836 1844
rect 812 1796 820 1804
rect 780 1776 788 1784
rect 764 1756 772 1764
rect 764 1736 772 1744
rect 620 1716 628 1724
rect 844 1756 852 1764
rect 700 1716 708 1724
rect 780 1716 788 1724
rect 892 1856 900 1864
rect 908 1796 916 1804
rect 940 1776 948 1784
rect 1004 1796 1012 1804
rect 1020 1756 1028 1764
rect 1116 1896 1124 1904
rect 1212 2276 1220 2284
rect 1420 2516 1428 2524
rect 1372 2496 1380 2504
rect 1340 2296 1348 2304
rect 1196 2116 1204 2124
rect 1388 2436 1396 2444
rect 1228 2256 1236 2264
rect 1324 2256 1332 2264
rect 1372 2256 1380 2264
rect 1244 2216 1252 2224
rect 1308 2136 1316 2144
rect 1180 2096 1188 2104
rect 1212 2096 1220 2104
rect 1260 2096 1268 2104
rect 1164 2056 1172 2064
rect 1148 2016 1156 2024
rect 1196 2076 1204 2084
rect 1180 1956 1188 1964
rect 1180 1936 1188 1944
rect 1196 1916 1204 1924
rect 1324 2116 1332 2124
rect 1468 2356 1476 2364
rect 1404 2296 1412 2304
rect 1436 2296 1444 2304
rect 1516 2516 1524 2524
rect 1500 2316 1508 2324
rect 1628 2596 1636 2604
rect 1564 2518 1572 2524
rect 1564 2516 1572 2518
rect 1804 2916 1812 2924
rect 1852 3016 1860 3024
rect 1836 2856 1844 2864
rect 1774 2806 1782 2814
rect 1788 2806 1796 2814
rect 1802 2806 1810 2814
rect 1708 2756 1716 2764
rect 1868 2936 1876 2944
rect 1756 2696 1764 2704
rect 1692 2656 1700 2664
rect 1580 2296 1588 2304
rect 1500 2276 1508 2284
rect 1484 2256 1492 2264
rect 1468 2196 1476 2204
rect 1468 2176 1476 2184
rect 1452 2136 1460 2144
rect 1292 2096 1300 2104
rect 1356 2096 1364 2104
rect 1404 2096 1412 2104
rect 1436 2096 1444 2104
rect 1340 2076 1348 2084
rect 1276 2056 1284 2064
rect 1292 1916 1300 1924
rect 1132 1876 1140 1884
rect 1180 1876 1188 1884
rect 1420 2076 1428 2084
rect 1388 1936 1396 1944
rect 1404 1916 1412 1924
rect 1452 1896 1460 1904
rect 1532 2196 1540 2204
rect 1548 2176 1556 2184
rect 1676 2296 1684 2304
rect 1628 2116 1636 2124
rect 1580 1996 1588 2004
rect 1532 1916 1540 1924
rect 1516 1896 1524 1904
rect 1452 1876 1460 1884
rect 1500 1876 1508 1884
rect 1628 1936 1636 1944
rect 1724 2676 1732 2684
rect 1868 2676 1876 2684
rect 1756 2616 1764 2624
rect 1788 2596 1796 2604
rect 1868 2596 1876 2604
rect 1774 2406 1782 2414
rect 1788 2406 1796 2414
rect 1802 2406 1810 2414
rect 1724 2376 1732 2384
rect 1788 2236 1796 2244
rect 1740 2136 1748 2144
rect 1676 1956 1684 1964
rect 1692 1956 1700 1964
rect 1692 1936 1700 1944
rect 1660 1896 1668 1904
rect 1724 1916 1732 1924
rect 1980 3516 1988 3524
rect 2044 3516 2052 3524
rect 2092 3536 2100 3544
rect 2124 3536 2132 3544
rect 2172 3816 2180 3824
rect 2204 3776 2212 3784
rect 2172 3736 2180 3744
rect 2156 3656 2164 3664
rect 2156 3536 2164 3544
rect 2204 3536 2212 3544
rect 2284 3776 2292 3784
rect 2236 3676 2244 3684
rect 2188 3516 2196 3524
rect 2124 3496 2132 3504
rect 1996 3476 2004 3484
rect 2028 3476 2036 3484
rect 1916 3416 1924 3424
rect 1948 3416 1956 3424
rect 1916 3396 1924 3404
rect 1932 3356 1940 3364
rect 2188 3496 2196 3504
rect 2220 3496 2228 3504
rect 2316 3916 2324 3924
rect 2588 4316 2596 4324
rect 2588 4296 2596 4304
rect 2604 4296 2612 4304
rect 2588 4276 2596 4284
rect 2428 4156 2436 4164
rect 2444 4156 2452 4164
rect 2412 4136 2420 4144
rect 2412 4076 2420 4084
rect 2476 4156 2484 4164
rect 2508 4096 2516 4104
rect 2444 4056 2452 4064
rect 2396 3916 2404 3924
rect 2380 3896 2388 3904
rect 2348 3876 2356 3884
rect 2396 3816 2404 3824
rect 2300 3716 2308 3724
rect 2332 3718 2340 3724
rect 2332 3716 2340 3718
rect 2460 3836 2468 3844
rect 2428 3716 2436 3724
rect 2396 3696 2404 3704
rect 2460 3776 2468 3784
rect 2556 3836 2564 3844
rect 2492 3816 2500 3824
rect 2476 3756 2484 3764
rect 2652 4296 2660 4304
rect 2684 4276 2692 4284
rect 2636 4236 2644 4244
rect 2620 4176 2628 4184
rect 2588 4136 2596 4144
rect 2732 4236 2740 4244
rect 2796 4536 2804 4544
rect 2764 4436 2772 4444
rect 2796 4356 2804 4364
rect 2748 4216 2756 4224
rect 2652 4156 2660 4164
rect 2748 4156 2756 4164
rect 2636 4136 2644 4144
rect 2700 4136 2708 4144
rect 2796 4216 2804 4224
rect 2764 4136 2772 4144
rect 2684 4116 2692 4124
rect 2716 4116 2724 4124
rect 2636 4076 2644 4084
rect 2780 4096 2788 4104
rect 2716 4076 2724 4084
rect 2652 4056 2660 4064
rect 2844 4536 2852 4544
rect 2860 4516 2868 4524
rect 3036 4716 3044 4724
rect 3052 4716 3060 4724
rect 2924 4656 2932 4664
rect 2892 4556 2900 4564
rect 2908 4536 2916 4544
rect 2892 4436 2900 4444
rect 2876 4356 2884 4364
rect 2972 4676 2980 4684
rect 3020 4696 3028 4704
rect 3036 4656 3044 4664
rect 2988 4616 2996 4624
rect 2956 4576 2964 4584
rect 2940 4516 2948 4524
rect 2956 4516 2964 4524
rect 3036 4518 3044 4524
rect 3036 4516 3044 4518
rect 2940 4496 2948 4504
rect 2940 4436 2948 4444
rect 2860 4336 2868 4344
rect 2876 4336 2884 4344
rect 2924 4336 2932 4344
rect 2828 4316 2836 4324
rect 2860 4316 2868 4324
rect 3116 4756 3124 4764
rect 3148 4756 3156 4764
rect 3084 4736 3092 4744
rect 3148 4736 3156 4744
rect 3116 4716 3124 4724
rect 3116 4696 3124 4704
rect 6716 4816 6724 4824
rect 4830 4806 4838 4814
rect 4844 4806 4852 4814
rect 4858 4806 4866 4814
rect 3244 4796 3252 4804
rect 3212 4776 3220 4784
rect 6572 4776 6580 4784
rect 4892 4756 4900 4764
rect 5068 4756 5076 4764
rect 5084 4756 5092 4764
rect 5180 4756 5188 4764
rect 3340 4736 3348 4744
rect 4988 4736 4996 4744
rect 3820 4716 3828 4724
rect 4044 4716 4052 4724
rect 4284 4716 4292 4724
rect 4332 4716 4340 4724
rect 4524 4716 4532 4724
rect 4572 4716 4580 4724
rect 4876 4716 4884 4724
rect 3212 4702 3220 4704
rect 3212 4696 3220 4702
rect 3180 4676 3188 4684
rect 3244 4676 3252 4684
rect 3068 4636 3076 4644
rect 3180 4556 3188 4564
rect 3404 4636 3412 4644
rect 3310 4606 3318 4614
rect 3324 4606 3332 4614
rect 3338 4606 3346 4614
rect 3276 4556 3284 4564
rect 3404 4556 3412 4564
rect 3100 4536 3108 4544
rect 3244 4536 3252 4544
rect 3292 4536 3300 4544
rect 3372 4536 3380 4544
rect 3388 4536 3396 4544
rect 3212 4516 3220 4524
rect 3164 4496 3172 4504
rect 3228 4496 3236 4504
rect 3052 4416 3060 4424
rect 3052 4376 3060 4384
rect 3020 4356 3028 4364
rect 2988 4316 2996 4324
rect 2956 4296 2964 4304
rect 2940 4276 2948 4284
rect 2988 4276 2996 4284
rect 2844 4216 2852 4224
rect 2892 4216 2900 4224
rect 2828 4176 2836 4184
rect 2860 4176 2868 4184
rect 2876 4156 2884 4164
rect 2908 4156 2916 4164
rect 2940 4156 2948 4164
rect 2908 4136 2916 4144
rect 2988 4136 2996 4144
rect 2876 4116 2884 4124
rect 2924 4116 2932 4124
rect 2956 4116 2964 4124
rect 2828 4096 2836 4104
rect 2620 3896 2628 3904
rect 2812 3896 2820 3904
rect 2828 3896 2836 3904
rect 2620 3876 2628 3884
rect 2636 3856 2644 3864
rect 2572 3756 2580 3764
rect 2508 3736 2516 3744
rect 2492 3696 2500 3704
rect 2508 3636 2516 3644
rect 2540 3636 2548 3644
rect 2764 3796 2772 3804
rect 2652 3756 2660 3764
rect 2732 3716 2740 3724
rect 2572 3696 2580 3704
rect 2556 3576 2564 3584
rect 2316 3516 2324 3524
rect 2444 3516 2452 3524
rect 2460 3502 2468 3504
rect 2460 3496 2468 3502
rect 2524 3496 2532 3504
rect 2220 3476 2228 3484
rect 2284 3476 2292 3484
rect 2348 3476 2356 3484
rect 2428 3476 2436 3484
rect 2140 3456 2148 3464
rect 2300 3436 2308 3444
rect 2332 3436 2340 3444
rect 2012 3396 2020 3404
rect 1996 3376 2004 3384
rect 2044 3316 2052 3324
rect 1948 3296 1956 3304
rect 2012 3296 2020 3304
rect 1980 3096 1988 3104
rect 1964 3076 1972 3084
rect 2060 3076 2068 3084
rect 2236 3416 2244 3424
rect 2316 3396 2324 3404
rect 2204 3376 2212 3384
rect 2124 3356 2132 3364
rect 2156 3316 2164 3324
rect 2156 3296 2164 3304
rect 2220 3296 2228 3304
rect 2220 3256 2228 3264
rect 2300 3316 2308 3324
rect 2524 3436 2532 3444
rect 2556 3516 2564 3524
rect 2588 3576 2596 3584
rect 2636 3576 2644 3584
rect 2700 3576 2708 3584
rect 2940 3896 2948 3904
rect 3068 4336 3076 4344
rect 3132 4296 3140 4304
rect 3164 4296 3172 4304
rect 3100 4276 3108 4284
rect 3164 4276 3172 4284
rect 3004 4016 3012 4024
rect 3036 3996 3044 4004
rect 3036 3896 3044 3904
rect 2908 3876 2916 3884
rect 2988 3876 2996 3884
rect 2876 3776 2884 3784
rect 2876 3736 2884 3744
rect 3260 4516 3268 4524
rect 3276 4516 3284 4524
rect 3260 4496 3268 4504
rect 3516 4676 3524 4684
rect 3548 4676 3556 4684
rect 3436 4616 3444 4624
rect 3484 4616 3492 4624
rect 3484 4596 3492 4604
rect 3612 4636 3620 4644
rect 3644 4696 3652 4704
rect 3772 4696 3780 4704
rect 3820 4696 3828 4704
rect 3916 4702 3924 4704
rect 3916 4696 3924 4702
rect 3660 4676 3668 4684
rect 3692 4676 3700 4684
rect 3980 4676 3988 4684
rect 3676 4636 3684 4644
rect 3708 4636 3716 4644
rect 3852 4636 3860 4644
rect 3628 4596 3636 4604
rect 3516 4556 3524 4564
rect 3756 4556 3764 4564
rect 4332 4696 4340 4704
rect 4076 4676 4084 4684
rect 4044 4636 4052 4644
rect 4076 4636 4084 4644
rect 3916 4556 3924 4564
rect 3516 4536 3524 4544
rect 3660 4536 3668 4544
rect 3852 4536 3860 4544
rect 3436 4516 3444 4524
rect 3468 4516 3476 4524
rect 3340 4496 3348 4504
rect 3420 4496 3428 4504
rect 3372 4476 3380 4484
rect 3372 4456 3380 4464
rect 3292 4336 3300 4344
rect 3420 4376 3428 4384
rect 3388 4336 3396 4344
rect 3420 4316 3428 4324
rect 3516 4516 3524 4524
rect 3548 4516 3556 4524
rect 3500 4496 3508 4504
rect 3484 4456 3492 4464
rect 3436 4296 3444 4304
rect 3260 4276 3268 4284
rect 3372 4276 3380 4284
rect 3196 4256 3204 4264
rect 3244 4256 3252 4264
rect 3132 4176 3140 4184
rect 3148 4156 3156 4164
rect 3244 4236 3252 4244
rect 3244 4216 3252 4224
rect 3228 4176 3236 4184
rect 3628 4516 3636 4524
rect 3580 4476 3588 4484
rect 3564 4416 3572 4424
rect 3628 4416 3636 4424
rect 3532 4356 3540 4364
rect 3628 4336 3636 4344
rect 3532 4296 3540 4304
rect 3724 4518 3732 4524
rect 3724 4516 3732 4518
rect 3788 4516 3796 4524
rect 3916 4518 3924 4524
rect 3916 4516 3924 4518
rect 3868 4436 3876 4444
rect 3836 4316 3844 4324
rect 3452 4276 3460 4284
rect 3500 4276 3508 4284
rect 3564 4256 3572 4264
rect 3596 4256 3604 4264
rect 3740 4256 3748 4264
rect 3276 4216 3284 4224
rect 3388 4216 3396 4224
rect 3310 4206 3318 4214
rect 3324 4206 3332 4214
rect 3338 4206 3346 4214
rect 3276 4176 3284 4184
rect 3260 4136 3268 4144
rect 3148 4116 3156 4124
rect 3356 4116 3364 4124
rect 3068 4096 3076 4104
rect 3308 4096 3316 4104
rect 3052 3856 3060 3864
rect 2956 3836 2964 3844
rect 2972 3836 2980 3844
rect 3052 3836 3060 3844
rect 2892 3716 2900 3724
rect 2892 3696 2900 3704
rect 2924 3736 2932 3744
rect 2940 3736 2948 3744
rect 2908 3576 2916 3584
rect 2876 3536 2884 3544
rect 2828 3496 2836 3504
rect 2540 3356 2548 3364
rect 2444 3276 2452 3284
rect 2332 3236 2340 3244
rect 2348 3136 2356 3144
rect 2156 3096 2164 3104
rect 2252 3096 2260 3104
rect 2300 3096 2308 3104
rect 2108 3076 2116 3084
rect 2092 3056 2100 3064
rect 1932 2996 1940 3004
rect 1980 2996 1988 3004
rect 1916 2976 1924 2984
rect 1948 2956 1956 2964
rect 1964 2956 1972 2964
rect 1900 2936 1908 2944
rect 1916 2716 1924 2724
rect 1948 2676 1956 2684
rect 2220 3036 2228 3044
rect 2012 2956 2020 2964
rect 2060 2956 2068 2964
rect 2092 2956 2100 2964
rect 1996 2936 2004 2944
rect 2284 2936 2292 2944
rect 2204 2918 2212 2924
rect 2204 2916 2212 2918
rect 2268 2916 2276 2924
rect 2076 2896 2084 2904
rect 2060 2856 2068 2864
rect 1996 2696 2004 2704
rect 2028 2676 2036 2684
rect 1996 2636 2004 2644
rect 1916 2616 1924 2624
rect 1964 2616 1972 2624
rect 2028 2536 2036 2544
rect 2332 3076 2340 3084
rect 2236 2896 2244 2904
rect 2268 2896 2276 2904
rect 2284 2896 2292 2904
rect 2140 2876 2148 2884
rect 2092 2856 2100 2864
rect 2076 2836 2084 2844
rect 2076 2816 2084 2824
rect 2124 2836 2132 2844
rect 2108 2756 2116 2764
rect 2092 2716 2100 2724
rect 2092 2696 2100 2704
rect 2188 2716 2196 2724
rect 2140 2676 2148 2684
rect 2124 2556 2132 2564
rect 2188 2696 2196 2704
rect 2332 2916 2340 2924
rect 2316 2876 2324 2884
rect 2492 3316 2500 3324
rect 2508 3296 2516 3304
rect 2492 3156 2500 3164
rect 2684 3476 2692 3484
rect 2780 3476 2788 3484
rect 2860 3476 2868 3484
rect 2604 3436 2612 3444
rect 2572 3356 2580 3364
rect 2668 3356 2676 3364
rect 2556 3256 2564 3264
rect 2572 3096 2580 3104
rect 2652 3316 2660 3324
rect 2780 3436 2788 3444
rect 2764 3316 2772 3324
rect 2652 3296 2660 3304
rect 2636 3116 2644 3124
rect 2460 3076 2468 3084
rect 2508 3076 2516 3084
rect 2604 3076 2612 3084
rect 2700 3102 2708 3104
rect 2700 3096 2708 3102
rect 2764 3256 2772 3264
rect 2396 3036 2404 3044
rect 2412 3036 2420 3044
rect 2476 3036 2484 3044
rect 2428 3016 2436 3024
rect 2476 2976 2484 2984
rect 2524 2976 2532 2984
rect 2380 2936 2388 2944
rect 2460 2936 2468 2944
rect 2348 2836 2356 2844
rect 2444 2836 2452 2844
rect 2508 2916 2516 2924
rect 2508 2876 2516 2884
rect 2444 2816 2452 2824
rect 2460 2816 2468 2824
rect 2492 2816 2500 2824
rect 2332 2716 2340 2724
rect 2300 2696 2308 2704
rect 2332 2696 2340 2704
rect 2460 2696 2468 2704
rect 2476 2696 2484 2704
rect 2204 2556 2212 2564
rect 2076 2516 2084 2524
rect 2108 2516 2116 2524
rect 1996 2416 2004 2424
rect 1884 2356 1892 2364
rect 1916 2316 1924 2324
rect 2028 2316 2036 2324
rect 2060 2316 2068 2324
rect 1996 2296 2004 2304
rect 2012 2296 2020 2304
rect 2108 2296 2116 2304
rect 2428 2576 2436 2584
rect 2748 3016 2756 3024
rect 2684 2976 2692 2984
rect 2732 2976 2740 2984
rect 2652 2936 2660 2944
rect 2716 2936 2724 2944
rect 2860 3276 2868 3284
rect 2844 3256 2852 3264
rect 2828 3216 2836 3224
rect 2796 3136 2804 3144
rect 2780 2956 2788 2964
rect 2716 2916 2724 2924
rect 2540 2796 2548 2804
rect 2636 2796 2644 2804
rect 2524 2736 2532 2744
rect 2620 2736 2628 2744
rect 2828 3116 2836 3124
rect 2860 3116 2868 3124
rect 2828 3036 2836 3044
rect 2892 3496 2900 3504
rect 2956 3656 2964 3664
rect 2988 3756 2996 3764
rect 3036 3756 3044 3764
rect 3020 3736 3028 3744
rect 3052 3716 3060 3724
rect 3020 3536 3028 3544
rect 3116 4016 3124 4024
rect 3372 4076 3380 4084
rect 3148 3896 3156 3904
rect 3340 3896 3348 3904
rect 3100 3796 3108 3804
rect 3148 3876 3156 3884
rect 3260 3876 3268 3884
rect 3132 3718 3140 3724
rect 3132 3716 3140 3718
rect 3116 3536 3124 3544
rect 3036 3516 3044 3524
rect 3052 3516 3060 3524
rect 3020 3496 3028 3504
rect 2908 3476 2916 3484
rect 2988 3476 2996 3484
rect 3020 3476 3028 3484
rect 2892 3356 2900 3364
rect 2972 3456 2980 3464
rect 2956 3436 2964 3444
rect 2956 3356 2964 3364
rect 2892 3316 2900 3324
rect 2940 3116 2948 3124
rect 2908 3036 2916 3044
rect 2812 2956 2820 2964
rect 2860 2956 2868 2964
rect 2924 2996 2932 3004
rect 2876 2936 2884 2944
rect 2796 2776 2804 2784
rect 2764 2716 2772 2724
rect 2860 2916 2868 2924
rect 2892 2916 2900 2924
rect 2588 2696 2596 2704
rect 2796 2696 2804 2704
rect 2508 2676 2516 2684
rect 2636 2676 2644 2684
rect 2396 2556 2404 2564
rect 2444 2556 2452 2564
rect 2492 2556 2500 2564
rect 2236 2536 2244 2544
rect 2236 2516 2244 2524
rect 2156 2496 2164 2504
rect 2188 2496 2196 2504
rect 2316 2496 2324 2504
rect 2140 2436 2148 2444
rect 2300 2302 2308 2304
rect 2300 2296 2308 2302
rect 1868 2236 1876 2244
rect 1980 2236 1988 2244
rect 1820 2116 1828 2124
rect 1774 2006 1782 2014
rect 1788 2006 1796 2014
rect 1802 2006 1810 2014
rect 1788 1956 1796 1964
rect 1580 1876 1588 1884
rect 1084 1856 1092 1864
rect 1244 1856 1252 1864
rect 1564 1856 1572 1864
rect 1740 1856 1748 1864
rect 1132 1836 1140 1844
rect 1260 1816 1268 1824
rect 1148 1756 1156 1764
rect 1212 1756 1220 1764
rect 1292 1756 1300 1764
rect 972 1736 980 1744
rect 988 1736 996 1744
rect 1052 1736 1060 1744
rect 1084 1736 1092 1744
rect 636 1696 644 1704
rect 684 1696 692 1704
rect 716 1696 724 1704
rect 604 1656 612 1664
rect 636 1636 644 1644
rect 716 1676 724 1684
rect 732 1676 740 1684
rect 780 1676 788 1684
rect 812 1636 820 1644
rect 748 1596 756 1604
rect 684 1516 692 1524
rect 716 1516 724 1524
rect 588 1496 596 1504
rect 604 1496 612 1504
rect 684 1496 692 1504
rect 716 1496 724 1504
rect 556 1476 564 1484
rect 620 1476 628 1484
rect 332 1356 340 1364
rect 332 1316 340 1324
rect 380 1316 388 1324
rect 348 1296 356 1304
rect 540 1356 548 1364
rect 444 1336 452 1344
rect 460 1336 468 1344
rect 476 1316 484 1324
rect 524 1316 532 1324
rect 412 1296 420 1304
rect 316 1276 324 1284
rect 364 1276 372 1284
rect 284 1256 292 1264
rect 284 1176 292 1184
rect 268 1156 276 1164
rect 300 1136 308 1144
rect 284 1116 292 1124
rect 252 1076 260 1084
rect 236 1036 244 1044
rect 348 1256 356 1264
rect 396 1156 404 1164
rect 364 1136 372 1144
rect 332 1116 340 1124
rect 284 1056 292 1064
rect 348 1096 356 1104
rect 348 1016 356 1024
rect 268 976 276 984
rect 204 956 212 964
rect 76 936 84 944
rect 172 916 180 924
rect 188 896 196 904
rect 156 876 164 884
rect 156 856 164 864
rect 300 936 308 944
rect 236 916 244 924
rect 252 916 260 924
rect 316 916 324 924
rect 220 876 228 884
rect 236 876 244 884
rect 268 876 276 884
rect 204 816 212 824
rect 236 856 244 864
rect 252 816 260 824
rect 220 756 228 764
rect 60 736 68 744
rect 92 736 100 744
rect 188 716 196 724
rect 236 716 244 724
rect 12 676 20 684
rect 28 676 36 684
rect 108 696 116 704
rect 156 676 164 684
rect 204 676 212 684
rect 140 656 148 664
rect 156 656 164 664
rect 220 656 228 664
rect 124 636 132 644
rect 156 636 164 644
rect 108 576 116 584
rect 140 536 148 544
rect 12 516 20 524
rect 124 516 132 524
rect 12 496 20 504
rect 252 696 260 704
rect 284 696 292 704
rect 188 576 196 584
rect 236 556 244 564
rect 204 536 212 544
rect 220 536 228 544
rect 332 896 340 904
rect 444 1276 452 1284
rect 428 1156 436 1164
rect 428 1136 436 1144
rect 412 1096 420 1104
rect 796 1576 804 1584
rect 780 1476 788 1484
rect 668 1456 676 1464
rect 764 1456 772 1464
rect 588 1436 596 1444
rect 604 1436 612 1444
rect 572 1376 580 1384
rect 572 1356 580 1364
rect 620 1416 628 1424
rect 556 1296 564 1304
rect 588 1296 596 1304
rect 508 1276 516 1284
rect 764 1396 772 1404
rect 892 1696 900 1704
rect 972 1696 980 1704
rect 876 1596 884 1604
rect 876 1556 884 1564
rect 844 1536 852 1544
rect 860 1516 868 1524
rect 828 1496 836 1504
rect 956 1656 964 1664
rect 940 1576 948 1584
rect 956 1556 964 1564
rect 940 1536 948 1544
rect 812 1476 820 1484
rect 860 1476 868 1484
rect 892 1476 900 1484
rect 892 1456 900 1464
rect 972 1536 980 1544
rect 972 1516 980 1524
rect 924 1476 932 1484
rect 908 1436 916 1444
rect 796 1376 804 1384
rect 668 1336 676 1344
rect 780 1336 788 1344
rect 940 1336 948 1344
rect 684 1316 692 1324
rect 652 1296 660 1304
rect 684 1296 692 1304
rect 604 1276 612 1284
rect 732 1196 740 1204
rect 620 1176 628 1184
rect 540 1116 548 1124
rect 476 1096 484 1104
rect 588 1096 596 1104
rect 636 1136 644 1144
rect 668 1116 676 1124
rect 716 1096 724 1104
rect 460 1076 468 1084
rect 492 1076 500 1084
rect 556 1076 564 1084
rect 556 1056 564 1064
rect 700 1056 708 1064
rect 412 1016 420 1024
rect 364 996 372 1004
rect 364 976 372 984
rect 412 976 420 984
rect 364 936 372 944
rect 364 896 372 904
rect 348 756 356 764
rect 332 716 340 724
rect 396 916 404 924
rect 412 896 420 904
rect 412 876 420 884
rect 428 876 436 884
rect 428 736 436 744
rect 332 576 340 584
rect 300 556 308 564
rect 332 556 340 564
rect 284 536 292 544
rect 300 536 308 544
rect 364 536 372 544
rect 396 616 404 624
rect 492 956 500 964
rect 460 936 468 944
rect 540 976 548 984
rect 524 916 532 924
rect 604 996 612 1004
rect 556 956 564 964
rect 652 936 660 944
rect 476 896 484 904
rect 508 896 516 904
rect 572 896 580 904
rect 556 876 564 884
rect 508 776 516 784
rect 492 736 500 744
rect 524 736 532 744
rect 444 716 452 724
rect 460 716 468 724
rect 540 716 548 724
rect 572 716 580 724
rect 444 696 452 704
rect 508 696 516 704
rect 460 636 468 644
rect 428 536 436 544
rect 380 516 388 524
rect 412 516 420 524
rect 284 496 292 504
rect 268 476 276 484
rect 236 396 244 404
rect 252 396 260 404
rect 188 376 196 384
rect 76 336 84 344
rect 140 336 148 344
rect 44 276 52 284
rect 108 276 116 284
rect 172 276 180 284
rect 12 256 20 264
rect 156 256 164 264
rect 76 236 84 244
rect 220 356 228 364
rect 204 316 212 324
rect 92 136 100 144
rect 300 476 308 484
rect 348 476 356 484
rect 364 476 372 484
rect 412 476 420 484
rect 284 356 292 364
rect 268 316 276 324
rect 316 456 324 464
rect 380 436 388 444
rect 412 416 420 424
rect 380 356 388 364
rect 396 356 404 364
rect 556 676 564 684
rect 540 656 548 664
rect 556 616 564 624
rect 604 736 612 744
rect 700 976 708 984
rect 716 936 724 944
rect 636 916 644 924
rect 684 916 692 924
rect 652 756 660 764
rect 668 716 676 724
rect 620 696 628 704
rect 652 676 660 684
rect 604 656 612 664
rect 860 1256 868 1264
rect 812 1176 820 1184
rect 828 1156 836 1164
rect 748 1136 756 1144
rect 764 1116 772 1124
rect 796 1096 804 1104
rect 812 1096 820 1104
rect 796 1076 804 1084
rect 764 1056 772 1064
rect 732 916 740 924
rect 812 916 820 924
rect 892 1136 900 1144
rect 860 1116 868 1124
rect 876 1116 884 1124
rect 908 1116 916 1124
rect 876 1096 884 1104
rect 1004 1696 1012 1704
rect 1212 1696 1220 1704
rect 1244 1696 1252 1704
rect 1116 1676 1124 1684
rect 1516 1816 1524 1824
rect 1356 1796 1364 1804
rect 1420 1796 1428 1804
rect 1324 1756 1332 1764
rect 1468 1756 1476 1764
rect 1516 1756 1524 1764
rect 1548 1796 1556 1804
rect 1500 1736 1508 1744
rect 1308 1716 1316 1724
rect 1164 1676 1172 1684
rect 1260 1676 1268 1684
rect 1084 1656 1092 1664
rect 1132 1656 1140 1664
rect 1276 1656 1284 1664
rect 1020 1616 1028 1624
rect 1020 1576 1028 1584
rect 1084 1576 1092 1584
rect 1004 1356 1012 1364
rect 1036 1556 1044 1564
rect 1084 1536 1092 1544
rect 1100 1516 1108 1524
rect 1036 1476 1044 1484
rect 1324 1636 1332 1644
rect 1148 1556 1156 1564
rect 1212 1556 1220 1564
rect 1164 1536 1172 1544
rect 1196 1496 1204 1504
rect 1132 1476 1140 1484
rect 1196 1476 1204 1484
rect 1068 1456 1076 1464
rect 1324 1616 1332 1624
rect 1276 1596 1284 1604
rect 1308 1596 1316 1604
rect 1228 1496 1236 1504
rect 1244 1476 1252 1484
rect 1276 1476 1284 1484
rect 1036 1376 1044 1384
rect 1068 1376 1076 1384
rect 1052 1356 1060 1364
rect 1132 1376 1140 1384
rect 1020 1316 1028 1324
rect 1052 1316 1060 1324
rect 1084 1316 1092 1324
rect 988 1296 996 1304
rect 956 1236 964 1244
rect 972 1156 980 1164
rect 1020 1276 1028 1284
rect 1004 1196 1012 1204
rect 1004 1156 1012 1164
rect 988 1116 996 1124
rect 924 1076 932 1084
rect 876 996 884 1004
rect 860 976 868 984
rect 924 976 932 984
rect 908 936 916 944
rect 940 916 948 924
rect 844 896 852 904
rect 748 876 756 884
rect 828 876 836 884
rect 876 876 884 884
rect 940 876 948 884
rect 700 676 708 684
rect 700 616 708 624
rect 684 576 692 584
rect 588 536 596 544
rect 508 516 516 524
rect 524 516 532 524
rect 460 456 468 464
rect 508 476 516 484
rect 476 436 484 444
rect 444 416 452 424
rect 604 516 612 524
rect 828 776 836 784
rect 812 756 820 764
rect 844 756 852 764
rect 828 656 836 664
rect 780 576 788 584
rect 764 556 772 564
rect 764 536 772 544
rect 748 516 756 524
rect 796 516 804 524
rect 588 496 596 504
rect 572 476 580 484
rect 812 476 820 484
rect 652 416 660 424
rect 524 396 532 404
rect 556 396 564 404
rect 588 396 596 404
rect 444 376 452 384
rect 540 376 548 384
rect 428 356 436 364
rect 412 336 420 344
rect 348 316 356 324
rect 268 296 276 304
rect 316 296 324 304
rect 236 136 244 144
rect 300 136 308 144
rect 332 256 340 264
rect 460 316 468 324
rect 492 316 500 324
rect 572 356 580 364
rect 604 376 612 384
rect 620 356 628 364
rect 716 376 724 384
rect 732 376 740 384
rect 796 376 804 384
rect 668 336 676 344
rect 764 336 772 344
rect 860 736 868 744
rect 924 736 932 744
rect 1020 1096 1028 1104
rect 1036 1056 1044 1064
rect 1084 1276 1092 1284
rect 1084 1176 1092 1184
rect 1068 1136 1076 1144
rect 1052 1016 1060 1024
rect 1036 996 1044 1004
rect 1052 996 1060 1004
rect 1004 976 1012 984
rect 1020 976 1028 984
rect 1004 956 1012 964
rect 1020 916 1028 924
rect 972 896 980 904
rect 1148 1336 1156 1344
rect 1116 1316 1124 1324
rect 1132 1316 1140 1324
rect 1212 1416 1220 1424
rect 1276 1416 1284 1424
rect 1212 1376 1220 1384
rect 1244 1336 1252 1344
rect 1212 1276 1220 1284
rect 1116 1156 1124 1164
rect 1148 1156 1156 1164
rect 1116 1136 1124 1144
rect 1212 1216 1220 1224
rect 1164 1136 1172 1144
rect 1132 1056 1140 1064
rect 1100 996 1108 1004
rect 1100 956 1108 964
rect 1132 956 1140 964
rect 1228 1176 1236 1184
rect 1292 1396 1300 1404
rect 1292 1356 1300 1364
rect 1436 1676 1444 1684
rect 1404 1656 1412 1664
rect 1372 1616 1380 1624
rect 1372 1556 1380 1564
rect 1436 1616 1444 1624
rect 1420 1536 1428 1544
rect 1436 1536 1444 1544
rect 1500 1596 1508 1604
rect 1484 1516 1492 1524
rect 1324 1496 1332 1504
rect 1388 1496 1396 1504
rect 1516 1556 1524 1564
rect 1420 1476 1428 1484
rect 1500 1476 1508 1484
rect 1436 1456 1444 1464
rect 1356 1436 1364 1444
rect 1372 1436 1380 1444
rect 1324 1416 1332 1424
rect 1340 1316 1348 1324
rect 1324 1296 1332 1304
rect 1260 1156 1268 1164
rect 1244 1136 1252 1144
rect 1308 1256 1316 1264
rect 1292 1136 1300 1144
rect 1276 1116 1284 1124
rect 1180 1036 1188 1044
rect 1196 996 1204 1004
rect 1164 936 1172 944
rect 1180 936 1188 944
rect 1132 916 1140 924
rect 1100 896 1108 904
rect 1148 896 1156 904
rect 1196 896 1204 904
rect 1004 856 1012 864
rect 1036 856 1044 864
rect 972 756 980 764
rect 956 716 964 724
rect 940 676 948 684
rect 844 576 852 584
rect 876 636 884 644
rect 1036 796 1044 804
rect 1420 1356 1428 1364
rect 1468 1336 1476 1344
rect 1484 1296 1492 1304
rect 1388 1276 1396 1284
rect 1452 1276 1460 1284
rect 1468 1276 1476 1284
rect 1372 1216 1380 1224
rect 1356 1116 1364 1124
rect 1308 1076 1316 1084
rect 1372 1096 1380 1104
rect 1372 1076 1380 1084
rect 1276 1036 1284 1044
rect 1244 976 1252 984
rect 1276 1016 1284 1024
rect 1340 1036 1348 1044
rect 1324 956 1332 964
rect 1420 1136 1428 1144
rect 1484 1116 1492 1124
rect 1468 1096 1476 1104
rect 1484 1096 1492 1104
rect 1436 1076 1444 1084
rect 1404 1056 1412 1064
rect 1404 996 1412 1004
rect 1468 1056 1476 1064
rect 1484 1016 1492 1024
rect 1452 956 1460 964
rect 1388 936 1396 944
rect 1404 936 1412 944
rect 1468 936 1476 944
rect 1596 1776 1604 1784
rect 1612 1776 1620 1784
rect 1596 1736 1604 1744
rect 1692 1776 1700 1784
rect 1628 1756 1636 1764
rect 1644 1736 1652 1744
rect 1612 1716 1620 1724
rect 1564 1676 1572 1684
rect 1564 1576 1572 1584
rect 1532 1496 1540 1504
rect 1628 1596 1636 1604
rect 1708 1596 1716 1604
rect 1676 1556 1684 1564
rect 1612 1536 1620 1544
rect 1660 1536 1668 1544
rect 1596 1516 1604 1524
rect 1676 1516 1684 1524
rect 1836 1916 1844 1924
rect 1804 1876 1812 1884
rect 1836 1876 1844 1884
rect 1852 1796 1860 1804
rect 1852 1776 1860 1784
rect 1820 1716 1828 1724
rect 1788 1656 1796 1664
rect 1852 1636 1860 1644
rect 1774 1606 1782 1614
rect 1788 1606 1796 1614
rect 1802 1606 1810 1614
rect 1740 1536 1748 1544
rect 1900 2176 1908 2184
rect 1964 2116 1972 2124
rect 1884 1916 1892 1924
rect 2172 2236 2180 2244
rect 2076 2176 2084 2184
rect 2092 2136 2100 2144
rect 2460 2516 2468 2524
rect 2476 2516 2484 2524
rect 2396 2456 2404 2464
rect 2380 2316 2388 2324
rect 2364 2236 2372 2244
rect 2444 2396 2452 2404
rect 2700 2656 2708 2664
rect 2748 2656 2756 2664
rect 2620 2576 2628 2584
rect 2652 2576 2660 2584
rect 2668 2576 2676 2584
rect 2540 2556 2548 2564
rect 2588 2556 2596 2564
rect 2620 2536 2628 2544
rect 2684 2556 2692 2564
rect 2684 2536 2692 2544
rect 2508 2516 2516 2524
rect 2524 2516 2532 2524
rect 2636 2516 2644 2524
rect 2556 2496 2564 2504
rect 2492 2456 2500 2464
rect 2508 2416 2516 2424
rect 2748 2556 2756 2564
rect 2732 2516 2740 2524
rect 2748 2496 2756 2504
rect 2732 2456 2740 2464
rect 2476 2336 2484 2344
rect 2700 2336 2708 2344
rect 2460 2316 2468 2324
rect 2428 2296 2436 2304
rect 2780 2676 2788 2684
rect 2812 2676 2820 2684
rect 2892 2816 2900 2824
rect 3068 3316 3076 3324
rect 3020 3076 3028 3084
rect 2988 3056 2996 3064
rect 3052 3036 3060 3044
rect 2956 2996 2964 3004
rect 3020 2976 3028 2984
rect 3004 2936 3012 2944
rect 3310 3806 3318 3814
rect 3324 3806 3332 3814
rect 3338 3806 3346 3814
rect 3516 4236 3524 4244
rect 3484 4216 3492 4224
rect 3468 4136 3476 4144
rect 3420 4118 3428 4124
rect 3420 4116 3428 4118
rect 3388 4036 3396 4044
rect 3420 4036 3428 4044
rect 3404 3902 3412 3904
rect 3404 3896 3412 3902
rect 3436 4016 3444 4024
rect 3436 3836 3444 3844
rect 3484 3776 3492 3784
rect 3564 4216 3572 4224
rect 3548 4176 3556 4184
rect 3580 4156 3588 4164
rect 3644 4156 3652 4164
rect 3724 4156 3732 4164
rect 3756 4156 3764 4164
rect 3532 4116 3540 4124
rect 3692 4116 3700 4124
rect 3756 4116 3764 4124
rect 3884 4316 3892 4324
rect 3932 4316 3940 4324
rect 3932 4296 3940 4304
rect 3804 4176 3812 4184
rect 3868 4176 3876 4184
rect 3852 4156 3860 4164
rect 3564 4096 3572 4104
rect 3676 4096 3684 4104
rect 3740 4096 3748 4104
rect 3596 4076 3604 4084
rect 3660 4056 3668 4064
rect 3708 3956 3716 3964
rect 3628 3896 3636 3904
rect 3676 3896 3684 3904
rect 3548 3876 3556 3884
rect 3612 3880 3620 3884
rect 3612 3876 3620 3880
rect 3644 3876 3652 3884
rect 3532 3856 3540 3864
rect 3564 3856 3572 3864
rect 3564 3816 3572 3824
rect 3548 3796 3556 3804
rect 3356 3756 3364 3764
rect 3404 3756 3412 3764
rect 3516 3756 3524 3764
rect 3244 3736 3252 3744
rect 3276 3716 3284 3724
rect 3340 3716 3348 3724
rect 3468 3736 3476 3744
rect 3244 3596 3252 3604
rect 3388 3596 3396 3604
rect 3404 3576 3412 3584
rect 3340 3516 3348 3524
rect 3372 3516 3380 3524
rect 3260 3496 3268 3504
rect 3388 3476 3396 3484
rect 3310 3406 3318 3414
rect 3324 3406 3332 3414
rect 3338 3406 3346 3414
rect 3148 3376 3156 3384
rect 3164 3376 3172 3384
rect 3356 3376 3364 3384
rect 3420 3536 3428 3544
rect 3452 3716 3460 3724
rect 3452 3696 3460 3704
rect 3564 3736 3572 3744
rect 3644 3796 3652 3804
rect 3660 3776 3668 3784
rect 3612 3756 3620 3764
rect 3676 3756 3684 3764
rect 3628 3736 3636 3744
rect 3500 3716 3508 3724
rect 3580 3716 3588 3724
rect 3596 3716 3604 3724
rect 3676 3716 3684 3724
rect 3516 3696 3524 3704
rect 3548 3696 3556 3704
rect 3580 3696 3588 3704
rect 3660 3696 3668 3704
rect 3468 3556 3476 3564
rect 3436 3496 3444 3504
rect 3836 4116 3844 4124
rect 3788 4096 3796 4104
rect 4044 4436 4052 4444
rect 4316 4676 4324 4684
rect 4236 4636 4244 4644
rect 4300 4656 4308 4664
rect 4252 4616 4260 4624
rect 4108 4516 4116 4524
rect 4076 4376 4084 4384
rect 4060 4316 4068 4324
rect 3996 4302 4004 4304
rect 3996 4296 4004 4302
rect 4060 4296 4068 4304
rect 4092 4276 4100 4284
rect 3916 4156 3924 4164
rect 4076 4156 4084 4164
rect 3980 4136 3988 4144
rect 3932 4116 3940 4124
rect 3964 4096 3972 4104
rect 3804 4076 3812 4084
rect 3884 4076 3892 4084
rect 3772 4036 3780 4044
rect 4044 4076 4052 4084
rect 3900 4056 3908 4064
rect 3916 3936 3924 3944
rect 3788 3916 3796 3924
rect 3820 3896 3828 3904
rect 3980 3916 3988 3924
rect 3804 3876 3812 3884
rect 3900 3876 3908 3884
rect 3772 3856 3780 3864
rect 3788 3836 3796 3844
rect 3740 3816 3748 3824
rect 3916 3776 3924 3784
rect 3804 3756 3812 3764
rect 3788 3736 3796 3744
rect 3724 3696 3732 3704
rect 3692 3596 3700 3604
rect 3724 3556 3732 3564
rect 3660 3536 3668 3544
rect 3532 3516 3540 3524
rect 3468 3476 3476 3484
rect 3580 3476 3588 3484
rect 3116 3316 3124 3324
rect 3164 3316 3172 3324
rect 3100 3236 3108 3244
rect 3228 3236 3236 3244
rect 3100 3156 3108 3164
rect 3148 3156 3156 3164
rect 3132 3136 3140 3144
rect 3260 3136 3268 3144
rect 3148 3096 3156 3104
rect 3116 3076 3124 3084
rect 3324 3102 3332 3104
rect 3324 3096 3332 3102
rect 3388 3076 3396 3084
rect 3180 3056 3188 3064
rect 3100 3036 3108 3044
rect 3372 3036 3380 3044
rect 3084 2976 3092 2984
rect 3310 3006 3318 3014
rect 3324 3006 3332 3014
rect 3338 3006 3346 3014
rect 3212 2976 3220 2984
rect 3116 2816 3124 2824
rect 3180 2916 3188 2924
rect 3244 2918 3252 2924
rect 3244 2916 3252 2918
rect 3388 2896 3396 2904
rect 3180 2876 3188 2884
rect 3260 2876 3268 2884
rect 3036 2796 3044 2804
rect 3692 3496 3700 3504
rect 3756 3536 3764 3544
rect 3948 3736 3956 3744
rect 4092 4076 4100 4084
rect 4364 4676 4372 4684
rect 4396 4656 4404 4664
rect 4444 4636 4452 4644
rect 4300 4536 4308 4544
rect 4252 4516 4260 4524
rect 4316 4516 4324 4524
rect 4364 4536 4372 4544
rect 4380 4536 4388 4544
rect 4348 4496 4356 4504
rect 4140 4476 4148 4484
rect 4268 4476 4276 4484
rect 4156 4336 4164 4344
rect 4204 4336 4212 4344
rect 4140 4316 4148 4324
rect 4444 4576 4452 4584
rect 4380 4476 4388 4484
rect 4492 4656 4500 4664
rect 4492 4596 4500 4604
rect 4396 4356 4404 4364
rect 4364 4316 4372 4324
rect 4396 4316 4404 4324
rect 4508 4576 4516 4584
rect 4508 4556 4516 4564
rect 4604 4636 4612 4644
rect 4588 4616 4596 4624
rect 4572 4576 4580 4584
rect 4476 4456 4484 4464
rect 4572 4536 4580 4544
rect 4588 4536 4596 4544
rect 4524 4516 4532 4524
rect 4540 4496 4548 4504
rect 4476 4416 4484 4424
rect 4508 4416 4516 4424
rect 4556 4476 4564 4484
rect 4540 4456 4548 4464
rect 4540 4416 4548 4424
rect 4460 4336 4468 4344
rect 4524 4336 4532 4344
rect 4492 4316 4500 4324
rect 4236 4296 4244 4304
rect 4268 4296 4276 4304
rect 4444 4296 4452 4304
rect 4508 4296 4516 4304
rect 4124 4256 4132 4264
rect 4140 4236 4148 4244
rect 4124 4216 4132 4224
rect 4188 4276 4196 4284
rect 4316 4276 4324 4284
rect 4204 4196 4212 4204
rect 4156 4076 4164 4084
rect 4188 3956 4196 3964
rect 4108 3936 4116 3944
rect 4412 4196 4420 4204
rect 4428 4156 4436 4164
rect 4300 4136 4308 4144
rect 4492 4136 4500 4144
rect 4268 4116 4276 4124
rect 4364 4118 4372 4124
rect 4364 4116 4372 4118
rect 4476 4116 4484 4124
rect 4556 4316 4564 4324
rect 4604 4516 4612 4524
rect 4588 4476 4596 4484
rect 4684 4676 4692 4684
rect 4716 4656 4724 4664
rect 4780 4656 4788 4664
rect 4876 4676 4884 4684
rect 4828 4656 4836 4664
rect 4732 4616 4740 4624
rect 4812 4616 4820 4624
rect 4684 4596 4692 4604
rect 4924 4676 4932 4684
rect 4940 4656 4948 4664
rect 5084 4716 5092 4724
rect 5116 4716 5124 4724
rect 5164 4716 5172 4724
rect 5196 4736 5204 4744
rect 5276 4736 5284 4744
rect 5484 4736 5492 4744
rect 5516 4736 5524 4744
rect 5548 4736 5556 4744
rect 6172 4736 6180 4744
rect 6220 4736 6228 4744
rect 6524 4736 6532 4744
rect 5036 4676 5044 4684
rect 4988 4656 4996 4664
rect 5020 4656 5028 4664
rect 5068 4656 5076 4664
rect 4892 4636 4900 4644
rect 4956 4636 4964 4644
rect 5260 4716 5268 4724
rect 5340 4716 5348 4724
rect 5372 4716 5380 4724
rect 5420 4716 5428 4724
rect 5500 4716 5508 4724
rect 5660 4716 5668 4724
rect 5708 4716 5716 4724
rect 5100 4676 5108 4684
rect 5196 4676 5204 4684
rect 5100 4656 5108 4664
rect 5116 4656 5124 4664
rect 5164 4636 5172 4644
rect 4988 4616 4996 4624
rect 4956 4576 4964 4584
rect 5052 4576 5060 4584
rect 4716 4556 4724 4564
rect 4812 4556 4820 4564
rect 4652 4496 4660 4504
rect 4668 4496 4676 4504
rect 4620 4456 4628 4464
rect 4620 4436 4628 4444
rect 4684 4416 4692 4424
rect 4780 4536 4788 4544
rect 4700 4356 4708 4364
rect 4620 4336 4628 4344
rect 4604 4316 4612 4324
rect 4540 4296 4548 4304
rect 4572 4296 4580 4304
rect 4636 4316 4644 4324
rect 4668 4316 4676 4324
rect 4556 4156 4564 4164
rect 4572 4156 4580 4164
rect 4620 4156 4628 4164
rect 4540 4136 4548 4144
rect 4556 4136 4564 4144
rect 4524 4096 4532 4104
rect 4268 4076 4276 4084
rect 4300 3916 4308 3924
rect 4444 3916 4452 3924
rect 4124 3876 4132 3884
rect 4172 3836 4180 3844
rect 4076 3796 4084 3804
rect 4108 3796 4116 3804
rect 4124 3776 4132 3784
rect 4108 3736 4116 3744
rect 4060 3596 4068 3604
rect 3948 3536 3956 3544
rect 4012 3536 4020 3544
rect 4092 3536 4100 3544
rect 4028 3516 4036 3524
rect 4060 3516 4068 3524
rect 3820 3502 3828 3504
rect 3820 3496 3828 3502
rect 3788 3476 3796 3484
rect 3676 3456 3684 3464
rect 3852 3456 3860 3464
rect 3964 3456 3972 3464
rect 3996 3456 4004 3464
rect 3740 3376 3748 3384
rect 3452 3176 3460 3184
rect 3452 3136 3460 3144
rect 4140 3756 4148 3764
rect 4156 3696 4164 3704
rect 4156 3676 4164 3684
rect 4044 3456 4052 3464
rect 4028 3436 4036 3444
rect 3900 3336 3908 3344
rect 3980 3336 3988 3344
rect 3612 3318 3620 3324
rect 3612 3316 3620 3318
rect 3788 3316 3796 3324
rect 3852 3316 3860 3324
rect 3868 3316 3876 3324
rect 3916 3316 3924 3324
rect 3804 3296 3812 3304
rect 3772 3276 3780 3284
rect 3836 3276 3844 3284
rect 3852 3276 3860 3284
rect 3692 3216 3700 3224
rect 3708 3136 3716 3144
rect 3756 3136 3764 3144
rect 3660 3096 3668 3104
rect 3484 3076 3492 3084
rect 3532 3056 3540 3064
rect 3564 2976 3572 2984
rect 3740 3116 3748 3124
rect 3788 3116 3796 3124
rect 3820 3256 3828 3264
rect 3756 3076 3764 3084
rect 3804 3076 3812 3084
rect 3548 2956 3556 2964
rect 3500 2936 3508 2944
rect 3628 2936 3636 2944
rect 3532 2916 3540 2924
rect 3468 2896 3476 2904
rect 3436 2856 3444 2864
rect 2940 2716 2948 2724
rect 2956 2716 2964 2724
rect 3004 2716 3012 2724
rect 2796 2576 2804 2584
rect 2812 2576 2820 2584
rect 2828 2556 2836 2564
rect 2876 2556 2884 2564
rect 2828 2536 2836 2544
rect 2780 2516 2788 2524
rect 2796 2516 2804 2524
rect 2828 2496 2836 2504
rect 3100 2716 3108 2724
rect 3212 2716 3220 2724
rect 3244 2716 3252 2724
rect 3052 2696 3060 2704
rect 3132 2696 3140 2704
rect 2988 2676 2996 2684
rect 2988 2656 2996 2664
rect 2972 2596 2980 2604
rect 3276 2696 3284 2704
rect 3068 2676 3076 2684
rect 3148 2680 3156 2684
rect 3148 2676 3156 2680
rect 3036 2616 3044 2624
rect 3148 2656 3156 2664
rect 3132 2616 3140 2624
rect 3052 2576 3060 2584
rect 3116 2576 3124 2584
rect 2892 2536 2900 2544
rect 2924 2536 2932 2544
rect 2940 2536 2948 2544
rect 2988 2536 2996 2544
rect 2908 2516 2916 2524
rect 2892 2456 2900 2464
rect 2860 2356 2868 2364
rect 2780 2336 2788 2344
rect 2524 2316 2532 2324
rect 2604 2316 2612 2324
rect 2684 2316 2692 2324
rect 2764 2316 2772 2324
rect 2652 2296 2660 2304
rect 2716 2296 2724 2304
rect 2284 2136 2292 2144
rect 2460 2136 2468 2144
rect 2028 2118 2036 2124
rect 2028 2116 2036 2118
rect 2156 2116 2164 2124
rect 2172 1996 2180 2004
rect 2044 1956 2052 1964
rect 2108 1896 2116 1904
rect 2156 1896 2164 1904
rect 2220 2118 2228 2124
rect 2220 2116 2228 2118
rect 2316 2116 2324 2124
rect 2364 2116 2372 2124
rect 2316 2096 2324 2104
rect 2380 2096 2388 2104
rect 2364 1976 2372 1984
rect 2444 1976 2452 1984
rect 2364 1916 2372 1924
rect 2252 1896 2260 1904
rect 1900 1876 1908 1884
rect 1868 1516 1876 1524
rect 1756 1496 1764 1504
rect 1996 1856 2004 1864
rect 2060 1856 2068 1864
rect 2076 1796 2084 1804
rect 1964 1776 1972 1784
rect 1980 1776 1988 1784
rect 2044 1776 2052 1784
rect 2220 1796 2228 1804
rect 2156 1716 2164 1724
rect 2252 1716 2260 1724
rect 1948 1576 1956 1584
rect 2220 1556 2228 1564
rect 2060 1536 2068 1544
rect 2124 1536 2132 1544
rect 2172 1536 2180 1544
rect 1932 1516 1940 1524
rect 2012 1516 2020 1524
rect 2092 1516 2100 1524
rect 1964 1496 1972 1504
rect 1980 1496 1988 1504
rect 2572 2196 2580 2204
rect 2604 2136 2612 2144
rect 2444 1716 2452 1724
rect 2508 1718 2516 1724
rect 2508 1716 2516 1718
rect 2364 1676 2372 1684
rect 2380 1656 2388 1664
rect 2380 1556 2388 1564
rect 2444 1556 2452 1564
rect 2188 1496 2196 1504
rect 2012 1476 2020 1484
rect 2108 1476 2116 1484
rect 1692 1456 1700 1464
rect 1580 1436 1588 1444
rect 1692 1436 1700 1444
rect 1564 1416 1572 1424
rect 1660 1416 1668 1424
rect 1660 1356 1668 1364
rect 1548 1336 1556 1344
rect 1564 1336 1572 1344
rect 1676 1336 1684 1344
rect 1548 1296 1556 1304
rect 1532 1276 1540 1284
rect 1516 1196 1524 1204
rect 1628 1276 1636 1284
rect 1564 1136 1572 1144
rect 1548 1116 1556 1124
rect 1516 1056 1524 1064
rect 1516 996 1524 1004
rect 1580 1096 1588 1104
rect 1628 1076 1636 1084
rect 1564 1056 1572 1064
rect 1548 1016 1556 1024
rect 1532 976 1540 984
rect 1388 916 1396 924
rect 1452 916 1460 924
rect 1500 916 1508 924
rect 1260 896 1268 904
rect 1308 896 1316 904
rect 1372 896 1380 904
rect 1340 876 1348 884
rect 1292 796 1300 804
rect 1228 776 1236 784
rect 1244 776 1252 784
rect 1292 776 1300 784
rect 1212 756 1220 764
rect 1228 736 1236 744
rect 1068 716 1076 724
rect 1084 696 1092 704
rect 1132 696 1140 704
rect 972 636 980 644
rect 876 556 884 564
rect 924 556 932 564
rect 956 556 964 564
rect 860 516 868 524
rect 956 536 964 544
rect 940 516 948 524
rect 1084 676 1092 684
rect 1116 676 1124 684
rect 1148 676 1156 684
rect 1180 656 1188 664
rect 1036 616 1044 624
rect 1084 596 1092 604
rect 1180 596 1188 604
rect 1020 576 1028 584
rect 1084 556 1092 564
rect 1004 536 1012 544
rect 1068 536 1076 544
rect 1036 516 1044 524
rect 1020 496 1028 504
rect 892 456 900 464
rect 988 456 996 464
rect 844 416 852 424
rect 684 316 692 324
rect 716 316 724 324
rect 780 316 788 324
rect 812 276 820 284
rect 476 256 484 264
rect 780 256 788 264
rect 796 256 804 264
rect 492 236 500 244
rect 444 216 452 224
rect 364 196 372 204
rect 428 176 436 184
rect 524 176 532 184
rect 364 156 372 164
rect 412 156 420 164
rect 492 156 500 164
rect 348 136 356 144
rect 396 136 404 144
rect 460 136 468 144
rect 732 196 740 204
rect 748 196 756 204
rect 652 176 660 184
rect 636 136 644 144
rect 604 116 612 124
rect 556 96 564 104
rect 620 96 628 104
rect 716 136 724 144
rect 732 136 740 144
rect 732 116 740 124
rect 860 396 868 404
rect 876 316 884 324
rect 956 396 964 404
rect 988 336 996 344
rect 908 316 916 324
rect 972 316 980 324
rect 924 296 932 304
rect 1132 536 1140 544
rect 1212 696 1220 704
rect 1228 696 1236 704
rect 1212 636 1220 644
rect 1212 596 1220 604
rect 1196 556 1204 564
rect 1196 516 1204 524
rect 1052 476 1060 484
rect 1068 356 1076 364
rect 1116 476 1124 484
rect 1180 476 1188 484
rect 1132 336 1140 344
rect 924 276 932 284
rect 988 276 996 284
rect 1068 296 1076 304
rect 1148 316 1156 324
rect 1084 276 1092 284
rect 1148 276 1156 284
rect 1100 256 1108 264
rect 1116 256 1124 264
rect 844 196 852 204
rect 860 196 868 204
rect 1020 196 1028 204
rect 1036 196 1044 204
rect 828 156 836 164
rect 844 156 852 164
rect 764 136 772 144
rect 796 136 804 144
rect 812 136 820 144
rect 892 156 900 164
rect 1100 196 1108 204
rect 1068 156 1076 164
rect 1084 156 1092 164
rect 1148 236 1156 244
rect 1228 516 1236 524
rect 1260 736 1268 744
rect 1260 716 1268 724
rect 1308 716 1316 724
rect 1340 696 1348 704
rect 1388 756 1396 764
rect 1404 756 1412 764
rect 1372 736 1380 744
rect 1468 756 1476 764
rect 1532 876 1540 884
rect 1436 736 1444 744
rect 1484 736 1492 744
rect 1516 736 1524 744
rect 1420 716 1428 724
rect 1516 716 1524 724
rect 1532 716 1540 724
rect 1468 696 1476 704
rect 1532 696 1540 704
rect 1340 656 1348 664
rect 1356 656 1364 664
rect 1420 656 1428 664
rect 1452 656 1460 664
rect 1260 536 1268 544
rect 1260 516 1268 524
rect 1244 496 1252 504
rect 1420 616 1428 624
rect 1356 596 1364 604
rect 1372 596 1380 604
rect 1324 576 1332 584
rect 1404 556 1412 564
rect 1388 536 1396 544
rect 1292 456 1300 464
rect 1260 336 1268 344
rect 1308 436 1316 444
rect 1388 416 1396 424
rect 1388 376 1396 384
rect 1388 336 1396 344
rect 1564 976 1572 984
rect 1580 896 1588 904
rect 1548 576 1556 584
rect 1452 516 1460 524
rect 1516 536 1524 544
rect 1516 516 1524 524
rect 1500 496 1508 504
rect 1436 476 1444 484
rect 1532 476 1540 484
rect 1436 356 1444 364
rect 1372 316 1380 324
rect 1532 416 1540 424
rect 1516 356 1524 364
rect 1500 296 1508 304
rect 1196 276 1204 284
rect 1244 276 1252 284
rect 1260 276 1268 284
rect 1516 276 1524 284
rect 1580 776 1588 784
rect 1628 996 1636 1004
rect 1676 1296 1684 1304
rect 1676 1236 1684 1244
rect 1820 1456 1828 1464
rect 1740 1436 1748 1444
rect 1900 1436 1908 1444
rect 1708 1376 1716 1384
rect 1708 1336 1716 1344
rect 1772 1336 1780 1344
rect 1724 1296 1732 1304
rect 1820 1276 1828 1284
rect 1774 1206 1782 1214
rect 1788 1206 1796 1214
rect 1802 1206 1810 1214
rect 1692 1096 1700 1104
rect 1820 1096 1828 1104
rect 1692 1076 1700 1084
rect 1948 1416 1956 1424
rect 1932 1396 1940 1404
rect 1996 1396 2004 1404
rect 1916 1356 1924 1364
rect 2140 1436 2148 1444
rect 2156 1396 2164 1404
rect 2220 1476 2228 1484
rect 2252 1456 2260 1464
rect 2156 1376 2164 1384
rect 2252 1376 2260 1384
rect 2204 1356 2212 1364
rect 1868 1336 1876 1344
rect 2012 1336 2020 1344
rect 1852 1316 1860 1324
rect 1932 1316 1940 1324
rect 2060 1316 2068 1324
rect 1868 1296 1876 1304
rect 1884 1136 1892 1144
rect 1916 1136 1924 1144
rect 2060 1156 2068 1164
rect 1884 1096 1892 1104
rect 2028 1096 2036 1104
rect 2108 1316 2116 1324
rect 2124 1296 2132 1304
rect 2172 1296 2180 1304
rect 2220 1316 2228 1324
rect 2412 1496 2420 1504
rect 2524 1496 2532 1504
rect 2348 1476 2356 1484
rect 2380 1476 2388 1484
rect 2476 1476 2484 1484
rect 2508 1476 2516 1484
rect 2316 1436 2324 1444
rect 2348 1376 2356 1384
rect 2300 1356 2308 1364
rect 2300 1336 2308 1344
rect 2332 1336 2340 1344
rect 2316 1316 2324 1324
rect 2268 1296 2276 1304
rect 2284 1276 2292 1284
rect 2268 1156 2276 1164
rect 2140 1136 2148 1144
rect 2188 1136 2196 1144
rect 2204 1136 2212 1144
rect 2220 1136 2228 1144
rect 2300 1136 2308 1144
rect 2124 1116 2132 1124
rect 2172 1116 2180 1124
rect 2092 1096 2100 1104
rect 1724 1056 1732 1064
rect 1836 1056 1844 1064
rect 1948 1056 1956 1064
rect 1980 1056 1988 1064
rect 1852 1036 1860 1044
rect 1644 976 1652 984
rect 1660 976 1668 984
rect 1628 956 1636 964
rect 1612 916 1620 924
rect 1596 716 1604 724
rect 1596 696 1604 704
rect 1740 1016 1748 1024
rect 1708 936 1716 944
rect 1868 936 1876 944
rect 1676 916 1684 924
rect 1692 896 1700 904
rect 1724 896 1732 904
rect 1836 896 1844 904
rect 1724 876 1732 884
rect 1740 876 1748 884
rect 1820 876 1828 884
rect 1676 856 1684 864
rect 1580 656 1588 664
rect 1612 656 1620 664
rect 1596 596 1604 604
rect 1596 536 1604 544
rect 1628 576 1636 584
rect 1660 556 1668 564
rect 1692 716 1700 724
rect 1692 616 1700 624
rect 1692 576 1700 584
rect 1660 516 1668 524
rect 1580 476 1588 484
rect 1788 856 1796 864
rect 1820 856 1828 864
rect 1756 836 1764 844
rect 1724 696 1732 704
rect 1774 806 1782 814
rect 1788 806 1796 814
rect 1802 806 1810 814
rect 1788 776 1796 784
rect 1756 716 1764 724
rect 1852 876 1860 884
rect 1996 936 2004 944
rect 1932 916 1940 924
rect 1980 916 1988 924
rect 2012 916 2020 924
rect 2092 996 2100 1004
rect 2124 1096 2132 1104
rect 2156 996 2164 1004
rect 2140 976 2148 984
rect 2060 896 2068 904
rect 2108 896 2116 904
rect 2188 1096 2196 1104
rect 2444 1436 2452 1444
rect 2396 1416 2404 1424
rect 2364 1356 2372 1364
rect 2364 1336 2372 1344
rect 2428 1396 2436 1404
rect 2428 1356 2436 1364
rect 2236 1096 2244 1104
rect 2204 916 2212 924
rect 2284 1056 2292 1064
rect 2348 1056 2356 1064
rect 2300 996 2308 1004
rect 2380 1296 2388 1304
rect 2396 1196 2404 1204
rect 2572 1936 2580 1944
rect 2556 1916 2564 1924
rect 2716 2256 2724 2264
rect 2764 2296 2772 2304
rect 3052 2516 3060 2524
rect 3020 2496 3028 2504
rect 3148 2596 3156 2604
rect 3084 2516 3092 2524
rect 3100 2476 3108 2484
rect 3068 2456 3076 2464
rect 2892 2336 2900 2344
rect 2924 2336 2932 2344
rect 2812 2296 2820 2304
rect 2892 2296 2900 2304
rect 3308 2676 3316 2684
rect 3404 2676 3412 2684
rect 3308 2656 3316 2664
rect 3388 2656 3396 2664
rect 3452 2656 3460 2664
rect 3404 2616 3412 2624
rect 3310 2606 3318 2614
rect 3324 2606 3332 2614
rect 3338 2606 3346 2614
rect 3180 2576 3188 2584
rect 3260 2576 3268 2584
rect 3164 2536 3172 2544
rect 3164 2516 3172 2524
rect 3100 2356 3108 2364
rect 3132 2356 3140 2364
rect 3020 2316 3028 2324
rect 3148 2336 3156 2344
rect 3132 2316 3140 2324
rect 3164 2316 3172 2324
rect 2956 2296 2964 2304
rect 2892 2256 2900 2264
rect 2940 2256 2948 2264
rect 2828 2236 2836 2244
rect 2940 2236 2948 2244
rect 2972 2236 2980 2244
rect 3068 2276 3076 2284
rect 3116 2276 3124 2284
rect 3052 2236 3060 2244
rect 3004 2216 3012 2224
rect 3084 2216 3092 2224
rect 2876 2196 2884 2204
rect 3084 2196 3092 2204
rect 2764 2176 2772 2184
rect 2812 2176 2820 2184
rect 2908 2176 2916 2184
rect 2924 2176 2932 2184
rect 3036 2176 3044 2184
rect 2732 2156 2740 2164
rect 2780 2156 2788 2164
rect 2860 2156 2868 2164
rect 2892 2156 2900 2164
rect 2972 2156 2980 2164
rect 3020 2156 3028 2164
rect 2652 2136 2660 2144
rect 2780 2136 2788 2144
rect 2812 2136 2820 2144
rect 2988 2136 2996 2144
rect 3036 2136 3044 2144
rect 3068 2136 3076 2144
rect 3324 2556 3332 2564
rect 3196 2536 3204 2544
rect 3452 2536 3460 2544
rect 3244 2516 3252 2524
rect 3388 2518 3396 2524
rect 3388 2516 3396 2518
rect 3436 2516 3444 2524
rect 3244 2496 3252 2504
rect 3196 2476 3204 2484
rect 3644 2816 3652 2824
rect 3564 2696 3572 2704
rect 3548 2636 3556 2644
rect 3564 2636 3572 2644
rect 3548 2596 3556 2604
rect 3532 2576 3540 2584
rect 3516 2556 3524 2564
rect 3628 2616 3636 2624
rect 3836 3156 3844 3164
rect 4108 3436 4116 3444
rect 4108 3376 4116 3384
rect 4092 3356 4100 3364
rect 4076 3336 4084 3344
rect 4252 3876 4260 3884
rect 4604 4136 4612 4144
rect 4668 4296 4676 4304
rect 4716 4296 4724 4304
rect 4764 4516 4772 4524
rect 4860 4516 4868 4524
rect 4844 4496 4852 4504
rect 4940 4496 4948 4504
rect 5036 4536 5044 4544
rect 4988 4516 4996 4524
rect 5004 4496 5012 4504
rect 4956 4456 4964 4464
rect 4796 4416 4804 4424
rect 4830 4406 4838 4414
rect 4844 4406 4852 4414
rect 4858 4406 4866 4414
rect 4828 4376 4836 4384
rect 4780 4336 4788 4344
rect 4796 4296 4804 4304
rect 4652 4276 4660 4284
rect 4652 4256 4660 4264
rect 4700 4256 4708 4264
rect 4796 4196 4804 4204
rect 4732 4176 4740 4184
rect 4748 4136 4756 4144
rect 4620 4116 4628 4124
rect 4636 4116 4644 4124
rect 4652 4116 4660 4124
rect 4620 4096 4628 4104
rect 4684 4096 4692 4104
rect 4652 4076 4660 4084
rect 4636 3956 4644 3964
rect 4604 3936 4612 3944
rect 4492 3896 4500 3904
rect 4284 3856 4292 3864
rect 4284 3836 4292 3844
rect 4284 3816 4292 3824
rect 4268 3796 4276 3804
rect 4236 3776 4244 3784
rect 4220 3756 4228 3764
rect 4284 3736 4292 3744
rect 4268 3716 4276 3724
rect 4428 3876 4436 3884
rect 4460 3876 4468 3884
rect 4396 3856 4404 3864
rect 4364 3836 4372 3844
rect 4348 3816 4356 3824
rect 4332 3796 4340 3804
rect 4316 3736 4324 3744
rect 4348 3716 4356 3724
rect 4236 3696 4244 3704
rect 4332 3696 4340 3704
rect 4188 3676 4196 3684
rect 4252 3556 4260 3564
rect 4396 3756 4404 3764
rect 4412 3736 4420 3744
rect 4380 3676 4388 3684
rect 4572 3836 4580 3844
rect 4604 3816 4612 3824
rect 4444 3796 4452 3804
rect 4524 3796 4532 3804
rect 4508 3776 4516 3784
rect 4604 3776 4612 3784
rect 4444 3696 4452 3704
rect 4364 3596 4372 3604
rect 4316 3536 4324 3544
rect 4380 3536 4388 3544
rect 4396 3536 4404 3544
rect 4284 3516 4292 3524
rect 4236 3496 4244 3504
rect 4156 3436 4164 3444
rect 4140 3416 4148 3424
rect 4156 3396 4164 3404
rect 4140 3376 4148 3384
rect 4124 3316 4132 3324
rect 4028 3296 4036 3304
rect 4092 3296 4100 3304
rect 4124 3296 4132 3304
rect 4156 3296 4164 3304
rect 3996 3276 4004 3284
rect 4044 3276 4052 3284
rect 3980 3256 3988 3264
rect 3900 3136 3908 3144
rect 3996 3236 4004 3244
rect 3852 3116 3860 3124
rect 3868 3116 3876 3124
rect 3980 3116 3988 3124
rect 3884 3076 3892 3084
rect 3788 3056 3796 3064
rect 3740 3036 3748 3044
rect 3692 2996 3700 3004
rect 3756 2976 3764 2984
rect 3692 2936 3700 2944
rect 3932 3076 3940 3084
rect 3916 3016 3924 3024
rect 3900 2956 3908 2964
rect 3852 2936 3860 2944
rect 3820 2916 3828 2924
rect 3836 2876 3844 2884
rect 3804 2856 3812 2864
rect 3772 2836 3780 2844
rect 4028 3176 4036 3184
rect 4060 3176 4068 3184
rect 4220 3456 4228 3464
rect 4204 3396 4212 3404
rect 4172 3276 4180 3284
rect 4204 3256 4212 3264
rect 4236 3396 4244 3404
rect 4236 3316 4244 3324
rect 4300 3456 4308 3464
rect 4316 3456 4324 3464
rect 4284 3436 4292 3444
rect 4332 3436 4340 3444
rect 4268 3356 4276 3364
rect 4316 3356 4324 3364
rect 4268 3316 4276 3324
rect 4540 3756 4548 3764
rect 4556 3736 4564 3744
rect 4524 3696 4532 3704
rect 4492 3676 4500 3684
rect 4556 3616 4564 3624
rect 4508 3576 4516 3584
rect 4556 3556 4564 3564
rect 4556 3536 4564 3544
rect 4460 3516 4468 3524
rect 4476 3516 4484 3524
rect 4492 3496 4500 3504
rect 4540 3496 4548 3504
rect 4364 3436 4372 3444
rect 4492 3476 4500 3484
rect 4412 3336 4420 3344
rect 4332 3316 4340 3324
rect 4412 3316 4420 3324
rect 4252 3276 4260 3284
rect 4284 3276 4292 3284
rect 4220 3236 4228 3244
rect 4236 3236 4244 3244
rect 4124 3196 4132 3204
rect 4172 3196 4180 3204
rect 4316 3256 4324 3264
rect 4284 3216 4292 3224
rect 4236 3136 4244 3144
rect 4268 3136 4276 3144
rect 4284 3136 4292 3144
rect 4108 3116 4116 3124
rect 4124 3116 4132 3124
rect 4044 3096 4052 3104
rect 4076 3096 4084 3104
rect 3996 3076 4004 3084
rect 4092 3076 4100 3084
rect 4172 3096 4180 3104
rect 4124 3076 4132 3084
rect 4268 3096 4276 3104
rect 4412 3276 4420 3284
rect 4364 3196 4372 3204
rect 4396 3196 4404 3204
rect 4412 3196 4420 3204
rect 4508 3456 4516 3464
rect 4540 3456 4548 3464
rect 4588 3716 4596 3724
rect 4716 4096 4724 4104
rect 4652 3896 4660 3904
rect 4668 3836 4676 3844
rect 4700 3896 4708 3904
rect 4700 3876 4708 3884
rect 4988 4376 4996 4384
rect 4876 4316 4884 4324
rect 5020 4456 5028 4464
rect 5020 4396 5028 4404
rect 5100 4516 5108 4524
rect 5148 4516 5156 4524
rect 5052 4496 5060 4504
rect 5116 4496 5124 4504
rect 5276 4696 5284 4704
rect 5260 4676 5268 4684
rect 5244 4656 5252 4664
rect 5324 4696 5332 4704
rect 5292 4676 5300 4684
rect 5308 4676 5316 4684
rect 5388 4676 5396 4684
rect 5340 4636 5348 4644
rect 5340 4596 5348 4604
rect 5356 4596 5364 4604
rect 5244 4556 5252 4564
rect 5276 4516 5284 4524
rect 5180 4496 5188 4504
rect 5084 4476 5092 4484
rect 5132 4476 5140 4484
rect 5228 4476 5236 4484
rect 5148 4456 5156 4464
rect 5100 4416 5108 4424
rect 5084 4316 5092 4324
rect 4892 4296 4900 4304
rect 4860 4256 4868 4264
rect 4972 4256 4980 4264
rect 5036 4256 5044 4264
rect 4940 4236 4948 4244
rect 4940 4196 4948 4204
rect 4924 4156 4932 4164
rect 4844 4136 4852 4144
rect 4972 4116 4980 4124
rect 4972 4096 4980 4104
rect 4764 4076 4772 4084
rect 4812 4076 4820 4084
rect 4924 4076 4932 4084
rect 4956 4076 4964 4084
rect 4764 4036 4772 4044
rect 4924 4016 4932 4024
rect 4830 4006 4838 4014
rect 4844 4006 4852 4014
rect 4858 4006 4866 4014
rect 4764 3916 4772 3924
rect 4908 3916 4916 3924
rect 4956 3916 4964 3924
rect 4748 3896 4756 3904
rect 4796 3896 4804 3904
rect 4732 3876 4740 3884
rect 4892 3876 4900 3884
rect 4700 3856 4708 3864
rect 4684 3776 4692 3784
rect 4668 3756 4676 3764
rect 4684 3756 4692 3764
rect 4716 3816 4724 3824
rect 4620 3716 4628 3724
rect 4700 3716 4708 3724
rect 4620 3676 4628 3684
rect 4652 3696 4660 3704
rect 4636 3656 4644 3664
rect 4620 3556 4628 3564
rect 4620 3476 4628 3484
rect 4588 3416 4596 3424
rect 4524 3316 4532 3324
rect 4444 3296 4452 3304
rect 4444 3256 4452 3264
rect 4460 3256 4468 3264
rect 4428 3156 4436 3164
rect 4364 3116 4372 3124
rect 4380 3116 4388 3124
rect 4412 3116 4420 3124
rect 4332 3096 4340 3104
rect 4380 3096 4388 3104
rect 4428 3096 4436 3104
rect 3964 3016 3972 3024
rect 4220 3016 4228 3024
rect 3996 2996 4004 3004
rect 4012 2996 4020 3004
rect 4060 2996 4068 3004
rect 4076 2996 4084 3004
rect 4028 2976 4036 2984
rect 4012 2936 4020 2944
rect 3948 2876 3956 2884
rect 4396 3076 4404 3084
rect 4252 2996 4260 3004
rect 4364 2996 4372 3004
rect 4380 2996 4388 3004
rect 4044 2936 4052 2944
rect 4076 2916 4084 2924
rect 3884 2856 3892 2864
rect 3836 2736 3844 2744
rect 3692 2716 3700 2724
rect 3964 2696 3972 2704
rect 3756 2676 3764 2684
rect 3916 2676 3924 2684
rect 4108 2856 4116 2864
rect 4076 2656 4084 2664
rect 3660 2576 3668 2584
rect 3820 2636 3828 2644
rect 3612 2536 3620 2544
rect 3692 2536 3700 2544
rect 3580 2516 3588 2524
rect 3596 2516 3604 2524
rect 3516 2496 3524 2504
rect 3532 2496 3540 2504
rect 3484 2436 3492 2444
rect 3436 2396 3444 2404
rect 3356 2356 3364 2364
rect 3196 2316 3204 2324
rect 3372 2336 3380 2344
rect 3484 2316 3492 2324
rect 3180 2296 3188 2304
rect 3292 2296 3300 2304
rect 3388 2296 3396 2304
rect 3212 2276 3220 2284
rect 3260 2276 3268 2284
rect 3244 2256 3252 2264
rect 3356 2256 3364 2264
rect 3212 2216 3220 2224
rect 3196 2156 3204 2164
rect 3132 2136 3140 2144
rect 3100 2116 3108 2124
rect 2652 2036 2660 2044
rect 2636 1896 2644 1904
rect 2876 1976 2884 1984
rect 2908 1956 2916 1964
rect 2764 1896 2772 1904
rect 2700 1856 2708 1864
rect 2924 1936 2932 1944
rect 2812 1876 2820 1884
rect 3068 2096 3076 2104
rect 3116 1976 3124 1984
rect 3052 1956 3060 1964
rect 2988 1916 2996 1924
rect 2940 1896 2948 1904
rect 2956 1896 2964 1904
rect 3004 1896 3012 1904
rect 3052 1896 3060 1904
rect 3116 1896 3124 1904
rect 3036 1876 3044 1884
rect 2956 1856 2964 1864
rect 3100 1856 3108 1864
rect 2684 1776 2692 1784
rect 2780 1836 2788 1844
rect 2876 1816 2884 1824
rect 2908 1816 2916 1824
rect 2796 1776 2804 1784
rect 2604 1716 2612 1724
rect 2668 1716 2676 1724
rect 2604 1696 2612 1704
rect 2572 1656 2580 1664
rect 2636 1556 2644 1564
rect 2588 1536 2596 1544
rect 2780 1536 2788 1544
rect 2620 1516 2628 1524
rect 2636 1516 2644 1524
rect 2556 1496 2564 1504
rect 2684 1496 2692 1504
rect 2540 1476 2548 1484
rect 2572 1476 2580 1484
rect 2492 1336 2500 1344
rect 2556 1456 2564 1464
rect 2588 1456 2596 1464
rect 2620 1456 2628 1464
rect 2540 1316 2548 1324
rect 2524 1296 2532 1304
rect 2476 1196 2484 1204
rect 2476 1136 2484 1144
rect 2508 1136 2516 1144
rect 2572 1356 2580 1364
rect 2700 1476 2708 1484
rect 2812 1736 2820 1744
rect 2876 1736 2884 1744
rect 2972 1776 2980 1784
rect 3052 1756 3060 1764
rect 2940 1716 2948 1724
rect 2988 1716 2996 1724
rect 2876 1696 2884 1704
rect 2956 1696 2964 1704
rect 3180 2136 3188 2144
rect 3212 2096 3220 2104
rect 3148 1976 3156 1984
rect 3196 1936 3204 1944
rect 3310 2206 3318 2214
rect 3324 2206 3332 2214
rect 3338 2206 3346 2214
rect 3484 2276 3492 2284
rect 3420 2256 3428 2264
rect 3436 2256 3444 2264
rect 3500 2256 3508 2264
rect 3276 2176 3284 2184
rect 3404 2176 3412 2184
rect 3452 2176 3460 2184
rect 3260 2156 3268 2164
rect 3420 2156 3428 2164
rect 3308 2136 3316 2144
rect 3244 2116 3252 2124
rect 3340 2116 3348 2124
rect 3372 2116 3380 2124
rect 3260 1936 3268 1944
rect 3228 1896 3236 1904
rect 3260 1896 3268 1904
rect 3404 2096 3412 2104
rect 3436 1916 3444 1924
rect 3420 1896 3428 1904
rect 3212 1876 3220 1884
rect 3324 1876 3332 1884
rect 3340 1876 3348 1884
rect 3228 1856 3236 1864
rect 3148 1836 3156 1844
rect 3196 1836 3204 1844
rect 3244 1836 3252 1844
rect 3068 1736 3076 1744
rect 3100 1736 3108 1744
rect 3164 1756 3172 1764
rect 3180 1756 3188 1764
rect 3276 1836 3284 1844
rect 3404 1836 3412 1844
rect 3452 1836 3460 1844
rect 3310 1806 3318 1814
rect 3324 1806 3332 1814
rect 3338 1806 3346 1814
rect 3532 2316 3540 2324
rect 3724 2518 3732 2524
rect 3724 2516 3732 2518
rect 3628 2496 3636 2504
rect 3676 2376 3684 2384
rect 3580 2296 3588 2304
rect 3612 2296 3620 2304
rect 3868 2616 3876 2624
rect 4076 2616 4084 2624
rect 4092 2616 4100 2624
rect 3852 2576 3860 2584
rect 3916 2576 3924 2584
rect 4060 2576 4068 2584
rect 3932 2556 3940 2564
rect 4012 2556 4020 2564
rect 3836 2496 3844 2504
rect 3820 2356 3828 2364
rect 3532 2276 3540 2284
rect 3548 2256 3556 2264
rect 3820 2296 3828 2304
rect 3756 2236 3764 2244
rect 3612 2156 3620 2164
rect 3644 2156 3652 2164
rect 3548 2118 3556 2124
rect 3548 2116 3556 2118
rect 3548 1896 3556 1904
rect 3708 2136 3716 2144
rect 3740 2136 3748 2144
rect 3804 2256 3812 2264
rect 3788 2236 3796 2244
rect 3772 2136 3780 2144
rect 3660 2116 3668 2124
rect 4012 2536 4020 2544
rect 3980 2516 3988 2524
rect 4156 2936 4164 2944
rect 4268 2936 4276 2944
rect 4652 3416 4660 3424
rect 4748 3856 4756 3864
rect 4812 3856 4820 3864
rect 5116 4296 5124 4304
rect 5132 4256 5140 4264
rect 5116 4216 5124 4224
rect 5292 4456 5300 4464
rect 5676 4696 5684 4704
rect 5484 4676 5492 4684
rect 5564 4676 5572 4684
rect 5612 4676 5620 4684
rect 5676 4676 5684 4684
rect 5436 4656 5444 4664
rect 5500 4656 5508 4664
rect 5420 4616 5428 4624
rect 5548 4636 5556 4644
rect 6108 4716 6116 4724
rect 6204 4716 6212 4724
rect 5964 4696 5972 4704
rect 6060 4696 6068 4704
rect 5740 4676 5748 4684
rect 5772 4676 5780 4684
rect 5836 4676 5844 4684
rect 5884 4676 5892 4684
rect 5916 4676 5924 4684
rect 5948 4676 5956 4684
rect 5708 4656 5716 4664
rect 5820 4656 5828 4664
rect 5708 4636 5716 4644
rect 5804 4636 5812 4644
rect 5644 4616 5652 4624
rect 5596 4596 5604 4604
rect 5628 4596 5636 4604
rect 5564 4576 5572 4584
rect 5372 4496 5380 4504
rect 5308 4436 5316 4444
rect 5244 4416 5252 4424
rect 5292 4376 5300 4384
rect 5164 4356 5172 4364
rect 5260 4356 5268 4364
rect 5228 4336 5236 4344
rect 5372 4416 5380 4424
rect 5324 4336 5332 4344
rect 5340 4316 5348 4324
rect 5324 4296 5332 4304
rect 5180 4276 5188 4284
rect 5196 4256 5204 4264
rect 5228 4256 5236 4264
rect 5148 4176 5156 4184
rect 5116 4156 5124 4164
rect 5052 4136 5060 4144
rect 5100 4136 5108 4144
rect 5228 4136 5236 4144
rect 4988 3876 4996 3884
rect 5004 3856 5012 3864
rect 4780 3836 4788 3844
rect 4940 3836 4948 3844
rect 4748 3776 4756 3784
rect 4924 3776 4932 3784
rect 5260 4276 5268 4284
rect 5260 4156 5268 4164
rect 5196 4096 5204 4104
rect 5164 4036 5172 4044
rect 5068 4016 5076 4024
rect 5052 3996 5060 4004
rect 5068 3956 5076 3964
rect 5052 3916 5060 3924
rect 5404 4496 5412 4504
rect 5388 4376 5396 4384
rect 5388 4336 5396 4344
rect 5436 4516 5444 4524
rect 5468 4496 5476 4504
rect 5532 4456 5540 4464
rect 5420 4436 5428 4444
rect 5468 4436 5476 4444
rect 5516 4436 5524 4444
rect 5436 4336 5444 4344
rect 5452 4336 5460 4344
rect 5420 4316 5428 4324
rect 5404 4296 5412 4304
rect 5388 4276 5396 4284
rect 5404 4256 5412 4264
rect 5484 4296 5492 4304
rect 5500 4296 5508 4304
rect 5516 4296 5524 4304
rect 5548 4296 5556 4304
rect 5468 4276 5476 4284
rect 5468 4156 5476 4164
rect 5420 4136 5428 4144
rect 5324 4116 5332 4124
rect 5372 4116 5380 4124
rect 5308 4096 5316 4104
rect 5340 4096 5348 4104
rect 5404 4076 5412 4084
rect 5276 4036 5284 4044
rect 5340 4036 5348 4044
rect 5244 3996 5252 4004
rect 5228 3936 5236 3944
rect 5148 3916 5156 3924
rect 5196 3916 5204 3924
rect 5084 3896 5092 3904
rect 5132 3896 5140 3904
rect 5164 3896 5172 3904
rect 5100 3876 5108 3884
rect 5212 3896 5220 3904
rect 5068 3856 5076 3864
rect 5180 3856 5188 3864
rect 5020 3776 5028 3784
rect 5036 3776 5044 3784
rect 4764 3756 4772 3764
rect 4860 3756 4868 3764
rect 4908 3756 4916 3764
rect 4972 3756 4980 3764
rect 4748 3696 4756 3704
rect 4780 3656 4788 3664
rect 4764 3616 4772 3624
rect 4748 3556 4756 3564
rect 4732 3536 4740 3544
rect 4716 3496 4724 3504
rect 4924 3736 4932 3744
rect 5100 3736 5108 3744
rect 5132 3816 5140 3824
rect 5212 3816 5220 3824
rect 5132 3736 5140 3744
rect 4940 3716 4948 3724
rect 5020 3716 5028 3724
rect 5036 3716 5044 3724
rect 5084 3716 5092 3724
rect 5212 3716 5220 3724
rect 5260 3896 5268 3904
rect 5260 3876 5268 3884
rect 5244 3856 5252 3864
rect 5244 3716 5252 3724
rect 4972 3696 4980 3704
rect 5132 3696 5140 3704
rect 5164 3676 5172 3684
rect 5196 3676 5204 3684
rect 4830 3606 4838 3614
rect 4844 3606 4852 3614
rect 4858 3606 4866 3614
rect 4924 3576 4932 3584
rect 5036 3536 5044 3544
rect 4764 3476 4772 3484
rect 4700 3456 4708 3464
rect 5068 3516 5076 3524
rect 5052 3496 5060 3504
rect 4796 3456 4804 3464
rect 4828 3456 4836 3464
rect 4668 3356 4676 3364
rect 4636 3316 4644 3324
rect 4684 3316 4692 3324
rect 4780 3416 4788 3424
rect 4892 3416 4900 3424
rect 4844 3396 4852 3404
rect 4780 3356 4788 3364
rect 4748 3316 4756 3324
rect 4828 3316 4836 3324
rect 4588 3296 4596 3304
rect 4620 3296 4628 3304
rect 4652 3296 4660 3304
rect 4700 3296 4708 3304
rect 4540 3256 4548 3264
rect 4476 3216 4484 3224
rect 4524 3216 4532 3224
rect 4620 3276 4628 3284
rect 4572 3236 4580 3244
rect 4588 3236 4596 3244
rect 4652 3236 4660 3244
rect 4556 3196 4564 3204
rect 4540 3176 4548 3184
rect 4572 3176 4580 3184
rect 4556 3136 4564 3144
rect 4636 3196 4644 3204
rect 4892 3316 4900 3324
rect 4828 3296 4836 3304
rect 4732 3276 4740 3284
rect 4780 3256 4788 3264
rect 4700 3236 4708 3244
rect 4812 3236 4820 3244
rect 4620 3136 4628 3144
rect 4636 3136 4644 3144
rect 4684 3196 4692 3204
rect 4668 3156 4676 3164
rect 4492 3116 4500 3124
rect 4556 3116 4564 3124
rect 4572 3116 4580 3124
rect 4460 3096 4468 3104
rect 4508 3076 4516 3084
rect 4460 3056 4468 3064
rect 4508 3036 4516 3044
rect 4572 3096 4580 3104
rect 4636 3096 4644 3104
rect 4588 3056 4596 3064
rect 4604 3056 4612 3064
rect 4556 2976 4564 2984
rect 4652 2976 4660 2984
rect 4524 2956 4532 2964
rect 4412 2916 4420 2924
rect 4460 2916 4468 2924
rect 4508 2936 4516 2944
rect 4588 2956 4596 2964
rect 4572 2936 4580 2944
rect 4652 2916 4660 2924
rect 4332 2896 4340 2904
rect 4396 2896 4404 2904
rect 4492 2896 4500 2904
rect 4412 2856 4420 2864
rect 4830 3206 4838 3214
rect 4844 3206 4852 3214
rect 4858 3206 4866 3214
rect 4748 3196 4756 3204
rect 4764 3156 4772 3164
rect 4700 3136 4708 3144
rect 4716 3136 4724 3144
rect 4812 3136 4820 3144
rect 5308 3956 5316 3964
rect 5468 4036 5476 4044
rect 5436 3936 5444 3944
rect 5292 3916 5300 3924
rect 5340 3916 5348 3924
rect 5452 3916 5460 3924
rect 5420 3876 5428 3884
rect 5452 3876 5460 3884
rect 5372 3856 5380 3864
rect 5500 4156 5508 4164
rect 5548 4276 5556 4284
rect 5532 4236 5540 4244
rect 5516 4116 5524 4124
rect 5580 4556 5588 4564
rect 5612 4556 5620 4564
rect 5708 4536 5716 4544
rect 5740 4536 5748 4544
rect 5980 4656 5988 4664
rect 6012 4656 6020 4664
rect 5996 4636 6004 4644
rect 6012 4636 6020 4644
rect 6076 4676 6084 4684
rect 6044 4636 6052 4644
rect 6108 4636 6116 4644
rect 6028 4616 6036 4624
rect 6124 4616 6132 4624
rect 6172 4616 6180 4624
rect 5948 4576 5956 4584
rect 5932 4556 5940 4564
rect 6028 4556 6036 4564
rect 6092 4556 6100 4564
rect 6124 4556 6132 4564
rect 6188 4556 6196 4564
rect 5868 4536 5876 4544
rect 5884 4536 5892 4544
rect 5964 4536 5972 4544
rect 6044 4536 6052 4544
rect 6108 4536 6116 4544
rect 5836 4516 5844 4524
rect 5756 4496 5764 4504
rect 5900 4496 5908 4504
rect 5692 4476 5700 4484
rect 5660 4456 5668 4464
rect 5580 4396 5588 4404
rect 5676 4376 5684 4384
rect 5612 4336 5620 4344
rect 5580 4316 5588 4324
rect 5596 4276 5604 4284
rect 5644 4276 5652 4284
rect 5628 4256 5636 4264
rect 5676 4276 5684 4284
rect 5676 4256 5684 4264
rect 5772 4476 5780 4484
rect 5852 4476 5860 4484
rect 5788 4456 5796 4464
rect 5724 4416 5732 4424
rect 5836 4436 5844 4444
rect 6012 4496 6020 4504
rect 6076 4476 6084 4484
rect 6076 4456 6084 4464
rect 5932 4416 5940 4424
rect 5804 4356 5812 4364
rect 5932 4316 5940 4324
rect 5964 4316 5972 4324
rect 5756 4296 5764 4304
rect 6012 4296 6020 4304
rect 5868 4276 5876 4284
rect 5740 4256 5748 4264
rect 5900 4256 5908 4264
rect 5916 4256 5924 4264
rect 5740 4236 5748 4244
rect 5804 4236 5812 4244
rect 5692 4216 5700 4224
rect 5868 4156 5876 4164
rect 5644 4136 5652 4144
rect 5580 4116 5588 4124
rect 5532 4016 5540 4024
rect 5644 4096 5652 4104
rect 5676 4076 5684 4084
rect 6092 4416 6100 4424
rect 6092 4376 6100 4384
rect 6076 4336 6084 4344
rect 6060 4316 6068 4324
rect 5980 4256 5988 4264
rect 6044 4256 6052 4264
rect 6108 4256 6116 4264
rect 5708 4136 5716 4144
rect 5804 4116 5812 4124
rect 5932 4156 5940 4164
rect 6060 4176 6068 4184
rect 6092 4176 6100 4184
rect 6076 4156 6084 4164
rect 5980 4136 5988 4144
rect 6012 4136 6020 4144
rect 5916 4116 5924 4124
rect 5932 4116 5940 4124
rect 5964 4116 5972 4124
rect 6012 4116 6020 4124
rect 6044 4116 6052 4124
rect 5996 4096 6004 4104
rect 6060 4096 6068 4104
rect 5852 4076 5860 4084
rect 5900 4076 5908 4084
rect 5708 4056 5716 4064
rect 5756 4056 5764 4064
rect 5836 4056 5844 4064
rect 5788 4016 5796 4024
rect 5628 3996 5636 4004
rect 5580 3976 5588 3984
rect 5564 3956 5572 3964
rect 5580 3936 5588 3944
rect 5612 3936 5620 3944
rect 5532 3916 5540 3924
rect 5596 3916 5604 3924
rect 5516 3896 5524 3904
rect 5596 3896 5604 3904
rect 5484 3856 5492 3864
rect 5532 3856 5540 3864
rect 5420 3836 5428 3844
rect 5468 3836 5476 3844
rect 5708 3976 5716 3984
rect 5692 3916 5700 3924
rect 5660 3896 5668 3904
rect 5740 3936 5748 3944
rect 5644 3876 5652 3884
rect 5708 3876 5716 3884
rect 5772 3876 5780 3884
rect 5740 3856 5748 3864
rect 5388 3796 5396 3804
rect 5548 3796 5556 3804
rect 5580 3796 5588 3804
rect 5644 3796 5652 3804
rect 5388 3736 5396 3744
rect 5516 3736 5524 3744
rect 5436 3716 5444 3724
rect 5500 3716 5508 3724
rect 5452 3696 5460 3704
rect 5260 3676 5268 3684
rect 5276 3676 5284 3684
rect 5404 3676 5412 3684
rect 5436 3676 5444 3684
rect 5340 3656 5348 3664
rect 5196 3516 5204 3524
rect 5228 3516 5236 3524
rect 5116 3496 5124 3504
rect 5308 3496 5316 3504
rect 5324 3496 5332 3504
rect 5180 3476 5188 3484
rect 5292 3476 5300 3484
rect 4956 3416 4964 3424
rect 4940 3356 4948 3364
rect 4940 3336 4948 3344
rect 4940 3316 4948 3324
rect 5132 3416 5140 3424
rect 5228 3416 5236 3424
rect 5004 3376 5012 3384
rect 5116 3396 5124 3404
rect 5020 3356 5028 3364
rect 5100 3356 5108 3364
rect 5004 3336 5012 3344
rect 5068 3336 5076 3344
rect 5004 3276 5012 3284
rect 5052 3276 5060 3284
rect 5068 3276 5076 3284
rect 4988 3256 4996 3264
rect 4924 3236 4932 3244
rect 4796 3116 4804 3124
rect 4700 3096 4708 3104
rect 4764 3096 4772 3104
rect 4780 3076 4788 3084
rect 4716 3036 4724 3044
rect 4796 2976 4804 2984
rect 4748 2936 4756 2944
rect 4636 2836 4644 2844
rect 4732 2916 4740 2924
rect 4812 2936 4820 2944
rect 4876 2936 4884 2944
rect 4924 3136 4932 3144
rect 4940 3116 4948 3124
rect 5180 3396 5188 3404
rect 5420 3636 5428 3644
rect 5436 3576 5444 3584
rect 5500 3696 5508 3704
rect 5532 3696 5540 3704
rect 5580 3716 5588 3724
rect 5596 3696 5604 3704
rect 5692 3756 5700 3764
rect 5676 3736 5684 3744
rect 5628 3676 5636 3684
rect 5660 3676 5668 3684
rect 5516 3656 5524 3664
rect 5548 3656 5556 3664
rect 5612 3656 5620 3664
rect 5484 3636 5492 3644
rect 5644 3636 5652 3644
rect 5500 3536 5508 3544
rect 5580 3536 5588 3544
rect 5596 3536 5604 3544
rect 5660 3536 5668 3544
rect 5388 3516 5396 3524
rect 5548 3516 5556 3524
rect 5420 3496 5428 3504
rect 5356 3476 5364 3484
rect 5324 3456 5332 3464
rect 5420 3456 5428 3464
rect 5452 3456 5460 3464
rect 5420 3436 5428 3444
rect 5532 3496 5540 3504
rect 5564 3496 5572 3504
rect 5580 3496 5588 3504
rect 5548 3456 5556 3464
rect 5244 3356 5252 3364
rect 5308 3356 5316 3364
rect 5148 3316 5156 3324
rect 5228 3316 5236 3324
rect 5148 3296 5156 3304
rect 5228 3296 5236 3304
rect 5292 3296 5300 3304
rect 5324 3296 5332 3304
rect 5132 3256 5140 3264
rect 5036 3176 5044 3184
rect 5116 3176 5124 3184
rect 5020 3136 5028 3144
rect 5068 3156 5076 3164
rect 5116 3156 5124 3164
rect 5164 3256 5172 3264
rect 5212 3256 5220 3264
rect 5180 3156 5188 3164
rect 4972 3096 4980 3104
rect 5052 3096 5060 3104
rect 5132 3096 5140 3104
rect 5164 3096 5172 3104
rect 5276 3276 5284 3284
rect 5340 3276 5348 3284
rect 5292 3256 5300 3264
rect 5372 3356 5380 3364
rect 5372 3336 5380 3344
rect 5484 3436 5492 3444
rect 5468 3416 5476 3424
rect 5532 3356 5540 3364
rect 5580 3396 5588 3404
rect 5820 3936 5828 3944
rect 5820 3896 5828 3904
rect 5820 3856 5828 3864
rect 5724 3696 5732 3704
rect 5756 3696 5764 3704
rect 5804 3696 5812 3704
rect 5820 3676 5828 3684
rect 5852 3936 5860 3944
rect 5884 3876 5892 3884
rect 5884 3856 5892 3864
rect 5868 3716 5876 3724
rect 5708 3556 5716 3564
rect 5612 3516 5620 3524
rect 5628 3516 5636 3524
rect 5692 3516 5700 3524
rect 5596 3376 5604 3384
rect 5644 3496 5652 3504
rect 5788 3596 5796 3604
rect 5628 3456 5636 3464
rect 5740 3456 5748 3464
rect 5756 3456 5764 3464
rect 5660 3396 5668 3404
rect 5644 3376 5652 3384
rect 5596 3356 5604 3364
rect 5468 3336 5476 3344
rect 5548 3336 5556 3344
rect 5436 3316 5444 3324
rect 5772 3416 5780 3424
rect 5804 3516 5812 3524
rect 5804 3496 5812 3504
rect 5804 3416 5812 3424
rect 5724 3376 5732 3384
rect 5772 3376 5780 3384
rect 5788 3376 5796 3384
rect 5788 3356 5796 3364
rect 5676 3336 5684 3344
rect 5420 3296 5428 3304
rect 5436 3296 5444 3304
rect 5612 3296 5620 3304
rect 5676 3296 5684 3304
rect 5404 3276 5412 3284
rect 5500 3256 5508 3264
rect 5660 3196 5668 3204
rect 5628 3156 5636 3164
rect 5564 3136 5572 3144
rect 5356 3116 5364 3124
rect 5324 3096 5332 3104
rect 5388 3096 5396 3104
rect 5516 3096 5524 3104
rect 5292 3076 5300 3084
rect 5068 3056 5076 3064
rect 5148 3056 5156 3064
rect 5212 3056 5220 3064
rect 5228 3056 5236 3064
rect 5276 3056 5284 3064
rect 4908 3036 4916 3044
rect 4972 3036 4980 3044
rect 4988 3036 4996 3044
rect 4988 2996 4996 3004
rect 5020 2996 5028 3004
rect 5020 2956 5028 2964
rect 5452 3076 5460 3084
rect 5580 3116 5588 3124
rect 5564 3096 5572 3104
rect 5532 3056 5540 3064
rect 5404 3036 5412 3044
rect 5404 2996 5412 3004
rect 5356 2976 5364 2984
rect 5612 3096 5620 3104
rect 5628 3036 5636 3044
rect 5644 3036 5652 3044
rect 5596 3016 5604 3024
rect 5500 2996 5508 3004
rect 5564 2996 5572 3004
rect 5452 2976 5460 2984
rect 5388 2956 5396 2964
rect 5484 2956 5492 2964
rect 5548 2956 5556 2964
rect 5564 2956 5572 2964
rect 5612 2956 5620 2964
rect 4924 2936 4932 2944
rect 4940 2916 4948 2924
rect 4748 2876 4756 2884
rect 4764 2856 4772 2864
rect 4828 2856 4836 2864
rect 4732 2836 4740 2844
rect 4140 2816 4148 2824
rect 4524 2816 4532 2824
rect 4700 2816 4708 2824
rect 4140 2716 4148 2724
rect 4268 2716 4276 2724
rect 4348 2716 4356 2724
rect 4444 2716 4452 2724
rect 4476 2716 4484 2724
rect 4540 2716 4548 2724
rect 4156 2696 4164 2704
rect 4332 2696 4340 2704
rect 4124 2676 4132 2684
rect 4156 2676 4164 2684
rect 4204 2676 4212 2684
rect 4300 2676 4308 2684
rect 4316 2676 4324 2684
rect 4172 2656 4180 2664
rect 4236 2656 4244 2664
rect 4316 2656 4324 2664
rect 4140 2616 4148 2624
rect 4172 2616 4180 2624
rect 4236 2616 4244 2624
rect 4284 2616 4292 2624
rect 4108 2556 4116 2564
rect 4220 2576 4228 2584
rect 4364 2680 4372 2684
rect 4364 2676 4372 2680
rect 4428 2676 4436 2684
rect 4348 2656 4356 2664
rect 4332 2556 4340 2564
rect 4364 2556 4372 2564
rect 4428 2616 4436 2624
rect 4428 2556 4436 2564
rect 4444 2556 4452 2564
rect 4348 2536 4356 2544
rect 4044 2516 4052 2524
rect 4188 2516 4196 2524
rect 4204 2516 4212 2524
rect 4300 2516 4308 2524
rect 3948 2496 3956 2504
rect 3996 2496 4004 2504
rect 4252 2476 4260 2484
rect 4396 2476 4404 2484
rect 4444 2476 4452 2484
rect 4188 2456 4196 2464
rect 3916 2376 3924 2384
rect 3884 2296 3892 2304
rect 3964 2296 3972 2304
rect 3916 2256 3924 2264
rect 3964 2256 3972 2264
rect 3868 2156 3876 2164
rect 3692 2096 3700 2104
rect 3724 2096 3732 2104
rect 3836 2096 3844 2104
rect 3660 1936 3668 1944
rect 3948 2096 3956 2104
rect 4508 2696 4516 2704
rect 4588 2696 4596 2704
rect 4716 2702 4724 2704
rect 4716 2696 4724 2702
rect 4492 2676 4500 2684
rect 4524 2676 4532 2684
rect 4492 2656 4500 2664
rect 4476 2536 4484 2544
rect 4492 2476 4500 2484
rect 4460 2456 4468 2464
rect 4268 2436 4276 2444
rect 4092 2376 4100 2384
rect 4140 2336 4148 2344
rect 4252 2316 4260 2324
rect 4044 2296 4052 2304
rect 3980 1996 3988 2004
rect 3708 1936 3716 1944
rect 3884 1936 3892 1944
rect 3692 1916 3700 1924
rect 3964 1916 3972 1924
rect 3852 1896 3860 1904
rect 3644 1876 3652 1884
rect 3724 1880 3732 1884
rect 3724 1876 3732 1880
rect 3756 1876 3764 1884
rect 4028 2276 4036 2284
rect 4108 2256 4116 2264
rect 4236 2256 4244 2264
rect 4252 2256 4260 2264
rect 4044 2236 4052 2244
rect 4028 2136 4036 2144
rect 4220 2216 4228 2224
rect 4300 2376 4308 2384
rect 4284 2316 4292 2324
rect 4572 2656 4580 2664
rect 4652 2636 4660 2644
rect 4620 2616 4628 2624
rect 4588 2536 4596 2544
rect 4572 2516 4580 2524
rect 4556 2496 4564 2504
rect 4572 2496 4580 2504
rect 4604 2516 4612 2524
rect 4524 2456 4532 2464
rect 4540 2456 4548 2464
rect 4412 2336 4420 2344
rect 4508 2336 4516 2344
rect 4332 2316 4340 2324
rect 4348 2316 4356 2324
rect 4316 2296 4324 2304
rect 4284 2216 4292 2224
rect 4204 2156 4212 2164
rect 4188 2136 4196 2144
rect 4364 2296 4372 2304
rect 4476 2296 4484 2304
rect 4396 2276 4404 2284
rect 4460 2276 4468 2284
rect 4716 2576 4724 2584
rect 4652 2536 4660 2544
rect 4636 2516 4644 2524
rect 4668 2516 4676 2524
rect 4700 2516 4708 2524
rect 4652 2476 4660 2484
rect 4668 2476 4676 2484
rect 4620 2336 4628 2344
rect 4636 2336 4644 2344
rect 4830 2806 4838 2814
rect 4844 2806 4852 2814
rect 4858 2806 4866 2814
rect 5052 2936 5060 2944
rect 5164 2936 5172 2944
rect 4972 2916 4980 2924
rect 5212 2916 5220 2924
rect 5356 2936 5364 2944
rect 5276 2916 5284 2924
rect 5308 2916 5316 2924
rect 5004 2896 5012 2904
rect 5020 2896 5028 2904
rect 5052 2896 5060 2904
rect 5132 2896 5140 2904
rect 5196 2896 5204 2904
rect 5244 2896 5252 2904
rect 5260 2896 5268 2904
rect 5356 2916 5364 2924
rect 5420 2936 5428 2944
rect 5516 2916 5524 2924
rect 5564 2916 5572 2924
rect 5468 2896 5476 2904
rect 5532 2896 5540 2904
rect 5580 2896 5588 2904
rect 5228 2876 5236 2884
rect 5292 2876 5300 2884
rect 5340 2876 5348 2884
rect 5596 2876 5604 2884
rect 5212 2856 5220 2864
rect 5564 2856 5572 2864
rect 4956 2776 4964 2784
rect 4908 2756 4916 2764
rect 4924 2716 4932 2724
rect 5324 2716 5332 2724
rect 5452 2716 5460 2724
rect 4956 2696 4964 2704
rect 4988 2696 4996 2704
rect 5068 2696 5076 2704
rect 5132 2702 5140 2704
rect 5132 2696 5140 2702
rect 4780 2656 4788 2664
rect 4844 2636 4852 2644
rect 4908 2636 4916 2644
rect 4876 2616 4884 2624
rect 4764 2556 4772 2564
rect 4748 2516 4756 2524
rect 4780 2456 4788 2464
rect 4732 2416 4740 2424
rect 4716 2376 4724 2384
rect 4780 2356 4788 2364
rect 4700 2316 4708 2324
rect 4588 2296 4596 2304
rect 4636 2296 4644 2304
rect 4732 2302 4740 2304
rect 4732 2296 4740 2302
rect 4524 2256 4532 2264
rect 4668 2236 4676 2244
rect 4524 2196 4532 2204
rect 4444 2156 4452 2164
rect 4508 2156 4516 2164
rect 4316 2136 4324 2144
rect 4508 2136 4516 2144
rect 4012 2096 4020 2104
rect 4028 2096 4036 2104
rect 4076 2096 4084 2104
rect 4236 2096 4244 2104
rect 4124 2036 4132 2044
rect 4364 2116 4372 2124
rect 4460 2116 4468 2124
rect 4444 2096 4452 2104
rect 4508 2096 4516 2104
rect 4492 2076 4500 2084
rect 4396 2056 4404 2064
rect 4252 1976 4260 1984
rect 4396 1976 4404 1984
rect 4476 1976 4484 1984
rect 4332 1916 4340 1924
rect 3980 1896 3988 1904
rect 4204 1896 4212 1904
rect 4268 1902 4276 1904
rect 4268 1896 4276 1902
rect 3692 1856 3700 1864
rect 3548 1776 3556 1784
rect 3436 1756 3444 1764
rect 3516 1756 3524 1764
rect 3292 1736 3300 1744
rect 3356 1736 3364 1744
rect 3180 1716 3188 1724
rect 3948 1836 3956 1844
rect 3740 1776 3748 1784
rect 4156 1876 4164 1884
rect 4028 1836 4036 1844
rect 4124 1836 4132 1844
rect 4076 1816 4084 1824
rect 3900 1736 3908 1744
rect 4012 1736 4020 1744
rect 3356 1716 3364 1724
rect 3452 1716 3460 1724
rect 3484 1716 3492 1724
rect 2844 1656 2852 1664
rect 2892 1596 2900 1604
rect 2876 1536 2884 1544
rect 2748 1476 2756 1484
rect 2668 1416 2676 1424
rect 2700 1416 2708 1424
rect 2668 1356 2676 1364
rect 2588 1336 2596 1344
rect 2620 1336 2628 1344
rect 2620 1316 2628 1324
rect 2572 1136 2580 1144
rect 2556 1116 2564 1124
rect 2460 1096 2468 1104
rect 2508 1096 2516 1104
rect 2732 1336 2740 1344
rect 2764 1376 2772 1384
rect 3228 1696 3236 1704
rect 3388 1696 3396 1704
rect 3548 1696 3556 1704
rect 3116 1656 3124 1664
rect 3292 1656 3300 1664
rect 2908 1516 2916 1524
rect 2892 1496 2900 1504
rect 2940 1496 2948 1504
rect 3612 1718 3620 1724
rect 3612 1716 3620 1718
rect 3676 1716 3684 1724
rect 3756 1716 3764 1724
rect 3996 1716 4004 1724
rect 4108 1716 4116 1724
rect 4172 1856 4180 1864
rect 4220 1836 4228 1844
rect 4156 1796 4164 1804
rect 4204 1796 4212 1804
rect 4236 1816 4244 1824
rect 3884 1676 3892 1684
rect 3772 1576 3780 1584
rect 3900 1576 3908 1584
rect 3116 1556 3124 1564
rect 3580 1556 3588 1564
rect 3676 1536 3684 1544
rect 3724 1536 3732 1544
rect 4044 1576 4052 1584
rect 4060 1576 4068 1584
rect 3948 1556 3956 1564
rect 3932 1536 3940 1544
rect 3404 1516 3412 1524
rect 3436 1516 3444 1524
rect 3916 1516 3924 1524
rect 2796 1456 2804 1464
rect 2812 1436 2820 1444
rect 2796 1376 2804 1384
rect 2828 1376 2836 1384
rect 2876 1376 2884 1384
rect 2780 1356 2788 1364
rect 2780 1336 2788 1344
rect 2828 1356 2836 1364
rect 2748 1316 2756 1324
rect 2764 1276 2772 1284
rect 2700 1136 2708 1144
rect 2652 1096 2660 1104
rect 2364 976 2372 984
rect 2284 956 2292 964
rect 2188 896 2196 904
rect 2252 896 2260 904
rect 2268 896 2276 904
rect 1932 876 1940 884
rect 1964 876 1972 884
rect 2028 876 2036 884
rect 2060 876 2068 884
rect 2076 876 2084 884
rect 2140 876 2148 884
rect 1852 836 1860 844
rect 1900 836 1908 844
rect 1900 756 1908 764
rect 1852 736 1860 744
rect 1932 756 1940 764
rect 2012 856 2020 864
rect 2220 856 2228 864
rect 1980 836 1988 844
rect 2108 836 2116 844
rect 1996 776 2004 784
rect 2012 756 2020 764
rect 1980 736 1988 744
rect 1948 716 1956 724
rect 2044 716 2052 724
rect 2076 696 2084 704
rect 2204 816 2212 824
rect 2124 756 2132 764
rect 2220 736 2228 744
rect 2268 696 2276 704
rect 1884 676 1892 684
rect 1916 676 1924 684
rect 1996 676 2004 684
rect 1868 656 1876 664
rect 2012 636 2020 644
rect 2092 636 2100 644
rect 1996 556 2004 564
rect 2044 616 2052 624
rect 2044 596 2052 604
rect 2348 936 2356 944
rect 2380 896 2388 904
rect 2348 696 2356 704
rect 2444 956 2452 964
rect 2428 936 2436 944
rect 2412 916 2420 924
rect 2412 896 2420 904
rect 2396 696 2404 704
rect 2140 656 2148 664
rect 2284 656 2292 664
rect 2316 656 2324 664
rect 2492 896 2500 904
rect 2460 836 2468 844
rect 2556 936 2564 944
rect 2524 916 2532 924
rect 2508 856 2516 864
rect 2444 776 2452 784
rect 2508 756 2516 764
rect 2508 736 2516 744
rect 2460 716 2468 724
rect 2476 696 2484 704
rect 2364 656 2372 664
rect 2428 656 2436 664
rect 2300 636 2308 644
rect 2140 576 2148 584
rect 2108 556 2116 564
rect 2124 556 2132 564
rect 1740 536 1748 544
rect 2220 536 2228 544
rect 1708 516 1716 524
rect 1836 516 1844 524
rect 1852 496 1860 504
rect 1900 496 1908 504
rect 2108 496 2116 504
rect 1692 476 1700 484
rect 1820 476 1828 484
rect 2268 536 2276 544
rect 2300 536 2308 544
rect 2300 516 2308 524
rect 2604 916 2612 924
rect 2540 896 2548 904
rect 2604 836 2612 844
rect 2540 716 2548 724
rect 2572 716 2580 724
rect 2524 696 2532 704
rect 2508 656 2516 664
rect 2492 636 2500 644
rect 2444 556 2452 564
rect 2428 536 2436 544
rect 2380 516 2388 524
rect 2460 516 2468 524
rect 2268 496 2276 504
rect 2364 496 2372 504
rect 2476 496 2484 504
rect 2396 476 2404 484
rect 2428 476 2436 484
rect 2012 436 2020 444
rect 2236 436 2244 444
rect 2428 436 2436 444
rect 1628 416 1636 424
rect 1596 396 1604 404
rect 1628 376 1636 384
rect 1628 356 1636 364
rect 1692 356 1700 364
rect 1580 336 1588 344
rect 1612 336 1620 344
rect 1564 316 1572 324
rect 1774 406 1782 414
rect 1788 406 1796 414
rect 1802 406 1810 414
rect 1740 396 1748 404
rect 1708 336 1716 344
rect 1996 416 2004 424
rect 1756 336 1764 344
rect 1836 336 1844 344
rect 1868 336 1876 344
rect 1628 316 1636 324
rect 1692 316 1700 324
rect 1740 316 1748 324
rect 1868 316 1876 324
rect 1884 316 1892 324
rect 1708 296 1716 304
rect 1900 296 1908 304
rect 2044 396 2052 404
rect 2028 316 2036 324
rect 2012 296 2020 304
rect 2060 356 2068 364
rect 2092 356 2100 364
rect 2060 296 2068 304
rect 2108 316 2116 324
rect 2092 296 2100 304
rect 2124 296 2132 304
rect 1564 276 1572 284
rect 1644 276 1652 284
rect 1724 276 1732 284
rect 1820 276 1828 284
rect 2076 276 2084 284
rect 2140 276 2148 284
rect 1196 256 1204 264
rect 1292 256 1300 264
rect 1324 256 1332 264
rect 1548 256 1556 264
rect 1708 256 1716 264
rect 1116 156 1124 164
rect 1164 156 1172 164
rect 1292 236 1300 244
rect 1212 216 1220 224
rect 1260 196 1268 204
rect 1276 196 1284 204
rect 1004 136 1012 144
rect 1020 136 1028 144
rect 1260 136 1268 144
rect 860 116 868 124
rect 892 116 900 124
rect 684 96 692 104
rect 348 76 356 84
rect 444 76 452 84
rect 540 76 548 84
rect 588 76 596 84
rect 668 76 676 84
rect 748 96 756 104
rect 796 96 804 104
rect 716 76 724 84
rect 732 76 740 84
rect 540 56 548 64
rect 652 56 660 64
rect 668 56 676 64
rect 700 56 708 64
rect 716 56 724 64
rect 1244 116 1252 124
rect 956 76 964 84
rect 604 36 612 44
rect 1548 236 1556 244
rect 1324 216 1332 224
rect 1404 216 1412 224
rect 1436 176 1444 184
rect 1388 136 1396 144
rect 1484 136 1492 144
rect 1372 116 1380 124
rect 1468 116 1476 124
rect 1484 116 1492 124
rect 1612 176 1620 184
rect 1564 136 1572 144
rect 1660 136 1668 144
rect 1676 136 1684 144
rect 2204 396 2212 404
rect 2188 316 2196 324
rect 2172 276 2180 284
rect 2268 316 2276 324
rect 2364 316 2372 324
rect 2252 296 2260 304
rect 2220 256 2228 264
rect 2012 236 2020 244
rect 2156 236 2164 244
rect 2252 236 2260 244
rect 1804 176 1812 184
rect 1580 96 1588 104
rect 1564 76 1572 84
rect 2156 216 2164 224
rect 2028 196 2036 204
rect 1932 156 1940 164
rect 1964 156 1972 164
rect 1916 116 1924 124
rect 1820 96 1828 104
rect 1900 96 1908 104
rect 1948 96 1956 104
rect 1772 76 1780 84
rect 1884 76 1892 84
rect 1932 76 1940 84
rect 2108 156 2116 164
rect 1996 116 2004 124
rect 2076 116 2084 124
rect 2316 296 2324 304
rect 2380 296 2388 304
rect 2508 596 2516 604
rect 2908 1456 2916 1464
rect 2892 1336 2900 1344
rect 3164 1496 3172 1504
rect 3260 1496 3268 1504
rect 3436 1496 3444 1504
rect 3500 1496 3508 1504
rect 3644 1496 3652 1504
rect 3692 1496 3700 1504
rect 3740 1496 3748 1504
rect 2972 1476 2980 1484
rect 2956 1436 2964 1444
rect 2940 1416 2948 1424
rect 2972 1416 2980 1424
rect 2924 1396 2932 1404
rect 2972 1376 2980 1384
rect 2988 1376 2996 1384
rect 3020 1376 3028 1384
rect 3068 1376 3076 1384
rect 3116 1376 3124 1384
rect 2940 1316 2948 1324
rect 3244 1476 3252 1484
rect 3180 1416 3188 1424
rect 3212 1416 3220 1424
rect 3196 1376 3204 1384
rect 3228 1396 3236 1404
rect 3132 1316 3140 1324
rect 4028 1536 4036 1544
rect 4156 1536 4164 1544
rect 4076 1516 4084 1524
rect 4140 1516 4148 1524
rect 4332 1796 4340 1804
rect 4236 1736 4244 1744
rect 4444 1736 4452 1744
rect 4332 1716 4340 1724
rect 4508 1916 4516 1924
rect 4508 1856 4516 1864
rect 4540 2176 4548 2184
rect 4732 2176 4740 2184
rect 5516 2702 5524 2704
rect 5516 2696 5524 2702
rect 5196 2676 5204 2684
rect 5292 2676 5300 2684
rect 5100 2656 5108 2664
rect 4988 2636 4996 2644
rect 4940 2596 4948 2604
rect 4956 2536 4964 2544
rect 5036 2576 5044 2584
rect 4972 2516 4980 2524
rect 5068 2496 5076 2504
rect 4830 2406 4838 2414
rect 4844 2406 4852 2414
rect 4858 2406 4866 2414
rect 4796 2336 4804 2344
rect 4796 2296 4804 2304
rect 4876 2296 4884 2304
rect 4860 2236 4868 2244
rect 4796 2176 4804 2184
rect 4604 2136 4612 2144
rect 4668 2136 4676 2144
rect 4700 2136 4708 2144
rect 4924 2476 4932 2484
rect 5084 2476 5092 2484
rect 4972 2336 4980 2344
rect 5036 2416 5044 2424
rect 5164 2636 5172 2644
rect 5196 2576 5204 2584
rect 5260 2576 5268 2584
rect 5276 2576 5284 2584
rect 5324 2576 5332 2584
rect 5132 2556 5140 2564
rect 5164 2556 5172 2564
rect 5276 2556 5284 2564
rect 5180 2536 5188 2544
rect 5100 2416 5108 2424
rect 5292 2516 5300 2524
rect 5484 2536 5492 2544
rect 5420 2516 5428 2524
rect 5516 2516 5524 2524
rect 5308 2496 5316 2504
rect 5132 2456 5140 2464
rect 5644 2916 5652 2924
rect 5644 2876 5652 2884
rect 5740 3156 5748 3164
rect 5788 3156 5796 3164
rect 5692 3136 5700 3144
rect 5724 3136 5732 3144
rect 5692 3076 5700 3084
rect 5740 3076 5748 3084
rect 5788 3076 5796 3084
rect 5708 3056 5716 3064
rect 5772 3056 5780 3064
rect 5676 2856 5684 2864
rect 5884 3696 5892 3704
rect 5868 3656 5876 3664
rect 5868 3636 5876 3644
rect 5852 3596 5860 3604
rect 5868 3536 5876 3544
rect 5836 3516 5844 3524
rect 5836 3496 5844 3504
rect 5852 3496 5860 3504
rect 5852 3456 5860 3464
rect 5980 4056 5988 4064
rect 6044 3976 6052 3984
rect 6028 3956 6036 3964
rect 5980 3936 5988 3944
rect 5996 3936 6004 3944
rect 5932 3916 5940 3924
rect 5948 3916 5956 3924
rect 5996 3916 6004 3924
rect 5964 3896 5972 3904
rect 5980 3896 5988 3904
rect 5916 3716 5924 3724
rect 5964 3696 5972 3704
rect 5948 3676 5956 3684
rect 5932 3656 5940 3664
rect 5916 3596 5924 3604
rect 5916 3576 5924 3584
rect 5916 3536 5924 3544
rect 5932 3516 5940 3524
rect 5916 3496 5924 3504
rect 5932 3496 5940 3504
rect 6012 3876 6020 3884
rect 6060 3916 6068 3924
rect 6492 4716 6500 4724
rect 6252 4696 6260 4704
rect 6508 4696 6516 4704
rect 6316 4676 6324 4684
rect 6284 4656 6292 4664
rect 6140 4536 6148 4544
rect 6300 4536 6308 4544
rect 6188 4516 6196 4524
rect 6204 4516 6212 4524
rect 6172 4456 6180 4464
rect 6140 4436 6148 4444
rect 6188 4336 6196 4344
rect 6252 4496 6260 4504
rect 6316 4496 6324 4504
rect 6268 4476 6276 4484
rect 6284 4376 6292 4384
rect 6236 4356 6244 4364
rect 6284 4336 6292 4344
rect 6316 4336 6324 4344
rect 6300 4276 6308 4284
rect 6204 4256 6212 4264
rect 6284 4256 6292 4264
rect 6476 4616 6484 4624
rect 6380 4536 6388 4544
rect 6428 4516 6436 4524
rect 6492 4516 6500 4524
rect 6364 4496 6372 4504
rect 6444 4456 6452 4464
rect 6396 4416 6404 4424
rect 6428 4416 6436 4424
rect 6396 4396 6404 4404
rect 6460 4396 6468 4404
rect 6396 4356 6404 4364
rect 6380 4316 6388 4324
rect 6428 4316 6436 4324
rect 6348 4296 6356 4304
rect 6348 4276 6356 4284
rect 6124 4156 6132 4164
rect 6108 4136 6116 4144
rect 6124 4096 6132 4104
rect 6108 3956 6116 3964
rect 6204 4176 6212 4184
rect 6156 4136 6164 4144
rect 6188 4096 6196 4104
rect 6252 4216 6260 4224
rect 6220 4136 6228 4144
rect 6252 4116 6260 4124
rect 6236 4096 6244 4104
rect 6220 4076 6228 4084
rect 6156 4016 6164 4024
rect 6076 3896 6084 3904
rect 6076 3876 6084 3884
rect 6108 3836 6116 3844
rect 6044 3736 6052 3744
rect 6060 3736 6068 3744
rect 6092 3736 6100 3744
rect 6028 3716 6036 3724
rect 6092 3716 6100 3724
rect 6044 3696 6052 3704
rect 5980 3676 5988 3684
rect 5964 3656 5972 3664
rect 5964 3596 5972 3604
rect 5948 3476 5956 3484
rect 5996 3516 6004 3524
rect 5836 3336 5844 3344
rect 5820 3296 5828 3304
rect 5820 3216 5828 3224
rect 5820 3136 5828 3144
rect 5900 3436 5908 3444
rect 5900 3336 5908 3344
rect 5948 3436 5956 3444
rect 5932 3336 5940 3344
rect 5900 3316 5908 3324
rect 5916 3316 5924 3324
rect 6028 3676 6036 3684
rect 6076 3656 6084 3664
rect 6044 3596 6052 3604
rect 6060 3596 6068 3604
rect 6060 3556 6068 3564
rect 6044 3536 6052 3544
rect 6092 3616 6100 3624
rect 6316 4216 6324 4224
rect 6332 4176 6340 4184
rect 6300 4096 6308 4104
rect 6332 4076 6340 4084
rect 6380 4176 6388 4184
rect 6364 4096 6372 4104
rect 6284 4056 6292 4064
rect 6332 4056 6340 4064
rect 6236 3936 6244 3944
rect 6252 3936 6260 3944
rect 6268 3936 6276 3944
rect 6156 3916 6164 3924
rect 6348 4016 6356 4024
rect 6332 3996 6340 4004
rect 6156 3896 6164 3904
rect 6252 3896 6260 3904
rect 6316 3896 6324 3904
rect 6140 3856 6148 3864
rect 6268 3856 6276 3864
rect 6236 3836 6244 3844
rect 6188 3816 6196 3824
rect 6268 3796 6276 3804
rect 6172 3736 6180 3744
rect 6140 3716 6148 3724
rect 6220 3716 6228 3724
rect 6236 3696 6244 3704
rect 6412 4256 6420 4264
rect 6492 4456 6500 4464
rect 6556 4536 6564 4544
rect 6508 4436 6516 4444
rect 6476 4376 6484 4384
rect 6460 4336 6468 4344
rect 6492 4356 6500 4364
rect 6556 4416 6564 4424
rect 6540 4336 6548 4344
rect 6444 4296 6452 4304
rect 6476 4296 6484 4304
rect 6444 4276 6452 4284
rect 6460 4276 6468 4284
rect 6444 4176 6452 4184
rect 6460 4176 6468 4184
rect 6396 4156 6404 4164
rect 6444 4136 6452 4144
rect 6396 4096 6404 4104
rect 6412 4076 6420 4084
rect 6380 4056 6388 4064
rect 6396 4056 6404 4064
rect 6284 3736 6292 3744
rect 6156 3656 6164 3664
rect 6188 3656 6196 3664
rect 6220 3656 6228 3664
rect 6140 3636 6148 3644
rect 6124 3616 6132 3624
rect 6092 3596 6100 3604
rect 6108 3596 6116 3604
rect 6108 3556 6116 3564
rect 6092 3536 6100 3544
rect 6156 3576 6164 3584
rect 6172 3556 6180 3564
rect 6220 3556 6228 3564
rect 6156 3536 6164 3544
rect 6188 3536 6196 3544
rect 6140 3516 6148 3524
rect 6188 3516 6196 3524
rect 6028 3496 6036 3504
rect 6124 3496 6132 3504
rect 6044 3476 6052 3484
rect 6108 3456 6116 3464
rect 5980 3336 5988 3344
rect 6044 3356 6052 3364
rect 6092 3356 6100 3364
rect 6092 3336 6100 3344
rect 6124 3336 6132 3344
rect 6172 3336 6180 3344
rect 5900 3296 5908 3304
rect 5980 3316 5988 3324
rect 6012 3316 6020 3324
rect 5884 3216 5892 3224
rect 5916 3156 5924 3164
rect 5820 2996 5828 3004
rect 5852 3056 5860 3064
rect 5852 2976 5860 2984
rect 5756 2956 5764 2964
rect 5772 2956 5780 2964
rect 5804 2956 5812 2964
rect 5836 2956 5844 2964
rect 5708 2936 5716 2944
rect 5756 2936 5764 2944
rect 5756 2916 5764 2924
rect 5724 2896 5732 2904
rect 5692 2816 5700 2824
rect 5628 2696 5636 2704
rect 5708 2702 5716 2704
rect 5708 2696 5716 2702
rect 5644 2536 5652 2544
rect 5676 2536 5684 2544
rect 5580 2516 5588 2524
rect 5116 2356 5124 2364
rect 5228 2356 5236 2364
rect 5420 2356 5428 2364
rect 5452 2356 5460 2364
rect 5004 2276 5012 2284
rect 5116 2276 5124 2284
rect 5292 2336 5300 2344
rect 5164 2276 5172 2284
rect 5276 2276 5284 2284
rect 5148 2256 5156 2264
rect 5212 2256 5220 2264
rect 5164 2196 5172 2204
rect 5404 2296 5412 2304
rect 5372 2276 5380 2284
rect 5340 2196 5348 2204
rect 5372 2196 5380 2204
rect 5180 2176 5188 2184
rect 5228 2176 5236 2184
rect 5148 2156 5156 2164
rect 4812 2136 4820 2144
rect 4924 2136 4932 2144
rect 5036 2136 5044 2144
rect 5148 2136 5156 2144
rect 5084 2116 5092 2124
rect 5020 2096 5028 2104
rect 4828 2076 4836 2084
rect 5052 2076 5060 2084
rect 4700 2036 4708 2044
rect 4956 2036 4964 2044
rect 5036 2036 5044 2044
rect 4588 1996 4596 2004
rect 4636 1936 4644 1944
rect 4572 1916 4580 1924
rect 4652 1916 4660 1924
rect 4684 1916 4692 1924
rect 4668 1876 4676 1884
rect 4684 1856 4692 1864
rect 4636 1816 4644 1824
rect 4604 1796 4612 1804
rect 4524 1776 4532 1784
rect 4604 1776 4612 1784
rect 4492 1756 4500 1764
rect 4476 1736 4484 1744
rect 4460 1696 4468 1704
rect 4220 1556 4228 1564
rect 4188 1536 4196 1544
rect 4108 1496 4116 1504
rect 4140 1496 4148 1504
rect 4172 1496 4180 1504
rect 3452 1476 3460 1484
rect 3484 1476 3492 1484
rect 3596 1476 3604 1484
rect 3676 1476 3684 1484
rect 3804 1476 3812 1484
rect 3852 1476 3860 1484
rect 4140 1476 4148 1484
rect 3420 1456 3428 1464
rect 3276 1436 3284 1444
rect 3310 1406 3318 1414
rect 3324 1406 3332 1414
rect 3338 1406 3346 1414
rect 3388 1396 3396 1404
rect 3244 1376 3252 1384
rect 3260 1376 3268 1384
rect 3292 1376 3300 1384
rect 3404 1376 3412 1384
rect 3308 1356 3316 1364
rect 3388 1356 3396 1364
rect 3452 1356 3460 1364
rect 3468 1356 3476 1364
rect 3276 1316 3284 1324
rect 3404 1316 3412 1324
rect 3468 1316 3476 1324
rect 3836 1456 3844 1464
rect 3644 1416 3652 1424
rect 3516 1396 3524 1404
rect 3740 1396 3748 1404
rect 3644 1376 3652 1384
rect 3724 1376 3732 1384
rect 3500 1356 3508 1364
rect 3548 1356 3556 1364
rect 3628 1356 3636 1364
rect 3580 1336 3588 1344
rect 3660 1336 3668 1344
rect 3708 1336 3716 1344
rect 3548 1316 3556 1324
rect 3612 1316 3620 1324
rect 3708 1316 3716 1324
rect 2956 1296 2964 1304
rect 3052 1296 3060 1304
rect 3228 1296 3236 1304
rect 3452 1296 3460 1304
rect 3484 1296 3492 1304
rect 3564 1296 3572 1304
rect 2844 1276 2852 1284
rect 3148 1276 3156 1284
rect 3196 1276 3204 1284
rect 3484 1276 3492 1284
rect 3020 1256 3028 1264
rect 3228 1256 3236 1264
rect 2844 1156 2852 1164
rect 2956 1156 2964 1164
rect 2972 1136 2980 1144
rect 2876 1116 2884 1124
rect 2924 1116 2932 1124
rect 2956 1116 2964 1124
rect 2924 1096 2932 1104
rect 3020 1136 3028 1144
rect 3052 1116 3060 1124
rect 3084 1116 3092 1124
rect 3212 1176 3220 1184
rect 3036 1096 3044 1104
rect 3116 1096 3124 1104
rect 3180 1096 3188 1104
rect 3484 1176 3492 1184
rect 3548 1176 3556 1184
rect 3468 1156 3476 1164
rect 3276 1136 3284 1144
rect 3436 1116 3444 1124
rect 3244 1096 3252 1104
rect 3340 1096 3348 1104
rect 3372 1096 3380 1104
rect 2812 1076 2820 1084
rect 2876 1076 2884 1084
rect 2940 1076 2948 1084
rect 3004 1076 3012 1084
rect 3084 1076 3092 1084
rect 3148 1076 3156 1084
rect 3196 1076 3204 1084
rect 3228 1076 3236 1084
rect 2828 1056 2836 1064
rect 2892 1056 2900 1064
rect 2636 976 2644 984
rect 2732 976 2740 984
rect 2668 916 2676 924
rect 2620 816 2628 824
rect 2652 736 2660 744
rect 2620 716 2628 724
rect 2780 936 2788 944
rect 2732 916 2740 924
rect 2844 940 2852 944
rect 2844 936 2852 940
rect 2828 916 2836 924
rect 2780 896 2788 904
rect 2812 896 2820 904
rect 2732 776 2740 784
rect 2684 736 2692 744
rect 2780 776 2788 784
rect 2764 736 2772 744
rect 2748 716 2756 724
rect 2668 696 2676 704
rect 2700 696 2708 704
rect 2556 676 2564 684
rect 2588 676 2596 684
rect 2668 676 2676 684
rect 2556 656 2564 664
rect 2572 616 2580 624
rect 2796 736 2804 744
rect 2796 696 2804 704
rect 2844 676 2852 684
rect 2748 656 2756 664
rect 3100 956 3108 964
rect 3148 956 3156 964
rect 3052 936 3060 944
rect 3164 936 3172 944
rect 2892 916 2900 924
rect 2988 876 2996 884
rect 3036 876 3044 884
rect 3100 876 3108 884
rect 3004 756 3012 764
rect 3020 736 3028 744
rect 3068 736 3076 744
rect 2892 696 2900 704
rect 2924 676 2932 684
rect 2956 656 2964 664
rect 2860 636 2868 644
rect 2556 516 2564 524
rect 2556 476 2564 484
rect 2572 436 2580 444
rect 2620 616 2628 624
rect 2604 596 2612 604
rect 3212 916 3220 924
rect 3196 876 3204 884
rect 3244 876 3252 884
rect 3260 876 3268 884
rect 3310 1006 3318 1014
rect 3324 1006 3332 1014
rect 3338 1006 3346 1014
rect 3372 976 3380 984
rect 3356 956 3364 964
rect 3372 936 3380 944
rect 3436 936 3444 944
rect 3420 916 3428 924
rect 3388 896 3396 904
rect 3580 1136 3588 1144
rect 3548 1076 3556 1084
rect 3468 956 3476 964
rect 3468 936 3476 944
rect 3612 1276 3620 1284
rect 3692 1256 3700 1264
rect 3628 1176 3636 1184
rect 3612 1116 3620 1124
rect 3692 1116 3700 1124
rect 3724 1096 3732 1104
rect 3756 1356 3764 1364
rect 3916 1456 3924 1464
rect 4108 1456 4116 1464
rect 3964 1436 3972 1444
rect 3868 1416 3876 1424
rect 3900 1396 3908 1404
rect 4012 1396 4020 1404
rect 4108 1396 4116 1404
rect 4204 1456 4212 1464
rect 4156 1436 4164 1444
rect 4172 1436 4180 1444
rect 3964 1356 3972 1364
rect 3788 1336 3796 1344
rect 3836 1336 3844 1344
rect 4060 1376 4068 1384
rect 4092 1376 4100 1384
rect 4028 1356 4036 1364
rect 4092 1356 4100 1364
rect 3756 1316 3764 1324
rect 3820 1316 3828 1324
rect 3836 1316 3844 1324
rect 3852 1316 3860 1324
rect 3932 1316 3940 1324
rect 4012 1316 4020 1324
rect 4140 1356 4148 1364
rect 4268 1516 4276 1524
rect 4252 1476 4260 1484
rect 4188 1356 4196 1364
rect 4220 1356 4228 1364
rect 4252 1396 4260 1404
rect 4332 1496 4340 1504
rect 4620 1716 4628 1724
rect 4540 1696 4548 1704
rect 4684 1756 4692 1764
rect 4668 1736 4676 1744
rect 4652 1716 4660 1724
rect 4830 2006 4838 2014
rect 4844 2006 4852 2014
rect 4858 2006 4866 2014
rect 4892 1956 4900 1964
rect 4988 1956 4996 1964
rect 4940 1936 4948 1944
rect 4716 1916 4724 1924
rect 4764 1916 4772 1924
rect 4796 1916 4804 1924
rect 4892 1916 4900 1924
rect 4956 1916 4964 1924
rect 5020 1936 5028 1944
rect 4876 1896 4884 1904
rect 4924 1896 4932 1904
rect 5020 1896 5028 1904
rect 4988 1876 4996 1884
rect 5004 1876 5012 1884
rect 4908 1856 4916 1864
rect 4972 1856 4980 1864
rect 5004 1856 5012 1864
rect 4748 1836 4756 1844
rect 4732 1796 4740 1804
rect 4892 1796 4900 1804
rect 4812 1756 4820 1764
rect 4780 1736 4788 1744
rect 4716 1716 4724 1724
rect 4700 1696 4708 1704
rect 4796 1716 4804 1724
rect 4828 1716 4836 1724
rect 5212 2156 5220 2164
rect 5308 2156 5316 2164
rect 5340 2136 5348 2144
rect 5196 2116 5204 2124
rect 5292 2116 5300 2124
rect 5132 2096 5140 2104
rect 5260 2096 5268 2104
rect 5100 2056 5108 2064
rect 5068 2036 5076 2044
rect 5084 2036 5092 2044
rect 5068 2016 5076 2024
rect 5436 2336 5444 2344
rect 5516 2336 5524 2344
rect 5468 2316 5476 2324
rect 5452 2296 5460 2304
rect 5452 2276 5460 2284
rect 5420 2156 5428 2164
rect 5452 2136 5460 2144
rect 5388 2116 5396 2124
rect 5500 2156 5508 2164
rect 5516 2116 5524 2124
rect 5436 2096 5444 2104
rect 5372 2076 5380 2084
rect 5308 1976 5316 1984
rect 5212 1936 5220 1944
rect 5180 1916 5188 1924
rect 5164 1896 5172 1904
rect 5084 1856 5092 1864
rect 5116 1856 5124 1864
rect 5148 1776 5156 1784
rect 5196 1776 5204 1784
rect 5116 1756 5124 1764
rect 5388 2016 5396 2024
rect 5260 1896 5268 1904
rect 5292 1896 5300 1904
rect 5340 1896 5348 1904
rect 5356 1896 5364 1904
rect 5404 1916 5412 1924
rect 5404 1896 5412 1904
rect 5708 2476 5716 2484
rect 5596 2356 5604 2364
rect 5580 2216 5588 2224
rect 5916 3096 5924 3104
rect 5932 3076 5940 3084
rect 5884 3036 5892 3044
rect 5900 3016 5908 3024
rect 5964 3296 5972 3304
rect 5996 3296 6004 3304
rect 6044 3296 6052 3304
rect 6028 3276 6036 3284
rect 5980 3196 5988 3204
rect 5964 3136 5972 3144
rect 5996 3176 6004 3184
rect 5964 3076 5972 3084
rect 5948 3016 5956 3024
rect 5948 2996 5956 3004
rect 5884 2976 5892 2984
rect 5916 2976 5924 2984
rect 5788 2936 5796 2944
rect 5868 2936 5876 2944
rect 5964 2956 5972 2964
rect 5804 2916 5812 2924
rect 5900 2916 5908 2924
rect 5788 2896 5796 2904
rect 5868 2896 5876 2904
rect 5884 2896 5892 2904
rect 5948 2736 5956 2744
rect 5836 2636 5844 2644
rect 5772 2356 5780 2364
rect 5900 2518 5908 2524
rect 5900 2516 5908 2518
rect 5900 2376 5908 2384
rect 5708 2276 5716 2284
rect 5740 2276 5748 2284
rect 5708 2216 5716 2224
rect 5596 2136 5604 2144
rect 5660 2136 5668 2144
rect 5580 2116 5588 2124
rect 5596 2116 5604 2124
rect 5628 2116 5636 2124
rect 5548 2076 5556 2084
rect 5532 2036 5540 2044
rect 5516 2016 5524 2024
rect 5468 1976 5476 1984
rect 5500 1976 5508 1984
rect 5452 1936 5460 1944
rect 5516 1936 5524 1944
rect 5660 1936 5668 1944
rect 5708 1936 5716 1944
rect 5756 1936 5764 1944
rect 5548 1916 5556 1924
rect 5612 1916 5620 1924
rect 5692 1916 5700 1924
rect 5740 1916 5748 1924
rect 5452 1876 5460 1884
rect 5292 1856 5300 1864
rect 5388 1856 5396 1864
rect 5436 1856 5444 1864
rect 5228 1836 5236 1844
rect 5260 1836 5268 1844
rect 5308 1836 5316 1844
rect 5260 1776 5268 1784
rect 5212 1756 5220 1764
rect 5468 1776 5476 1784
rect 5292 1756 5300 1764
rect 5356 1756 5364 1764
rect 5404 1756 5412 1764
rect 5276 1736 5284 1744
rect 5308 1736 5316 1744
rect 5244 1716 5252 1724
rect 5404 1736 5412 1744
rect 5500 1716 5508 1724
rect 5084 1696 5092 1704
rect 4780 1676 4788 1684
rect 5036 1676 5044 1684
rect 5068 1676 5076 1684
rect 5132 1676 5140 1684
rect 4636 1656 4644 1664
rect 4748 1656 4756 1664
rect 4524 1636 4532 1644
rect 4508 1596 4516 1604
rect 4460 1576 4468 1584
rect 4492 1576 4500 1584
rect 4460 1556 4468 1564
rect 4556 1616 4564 1624
rect 4540 1596 4548 1604
rect 4396 1536 4404 1544
rect 4460 1536 4468 1544
rect 4364 1476 4372 1484
rect 4604 1616 4612 1624
rect 4412 1516 4420 1524
rect 4508 1516 4516 1524
rect 4572 1516 4580 1524
rect 4396 1496 4404 1504
rect 4492 1496 4500 1504
rect 4524 1496 4532 1504
rect 4588 1496 4596 1504
rect 4716 1616 4724 1624
rect 4668 1576 4676 1584
rect 4716 1576 4724 1584
rect 4396 1476 4404 1484
rect 4332 1456 4340 1464
rect 4348 1456 4356 1464
rect 4380 1456 4388 1464
rect 4300 1416 4308 1424
rect 4124 1336 4132 1344
rect 4156 1336 4164 1344
rect 4188 1336 4196 1344
rect 4236 1336 4244 1344
rect 3996 1276 4004 1284
rect 3772 1256 3780 1264
rect 3980 1256 3988 1264
rect 3772 1116 3780 1124
rect 3788 1096 3796 1104
rect 3644 1076 3652 1084
rect 3740 1076 3748 1084
rect 3836 1076 3844 1084
rect 3852 1056 3860 1064
rect 3596 996 3604 1004
rect 3580 976 3588 984
rect 3564 936 3572 944
rect 3356 876 3364 884
rect 3452 876 3460 884
rect 3276 856 3284 864
rect 3196 836 3204 844
rect 3260 836 3268 844
rect 3180 816 3188 824
rect 3276 796 3284 804
rect 3132 736 3140 744
rect 3228 736 3236 744
rect 3036 656 3044 664
rect 3004 636 3012 644
rect 3084 676 3092 684
rect 3116 716 3124 724
rect 3164 716 3172 724
rect 3148 696 3156 704
rect 3196 696 3204 704
rect 3132 676 3140 684
rect 3180 676 3188 684
rect 3228 676 3236 684
rect 2972 616 2980 624
rect 3052 616 3060 624
rect 2780 596 2788 604
rect 2988 596 2996 604
rect 3052 596 3060 604
rect 2732 576 2740 584
rect 2812 576 2820 584
rect 2940 576 2948 584
rect 2668 556 2676 564
rect 2604 516 2612 524
rect 2636 516 2644 524
rect 2652 496 2660 504
rect 2748 556 2756 564
rect 2844 536 2852 544
rect 2892 536 2900 544
rect 2700 496 2708 504
rect 2732 476 2740 484
rect 2764 476 2772 484
rect 2588 416 2596 424
rect 2492 396 2500 404
rect 2460 336 2468 344
rect 2508 376 2516 384
rect 2732 376 2740 384
rect 2476 316 2484 324
rect 2668 356 2676 364
rect 2732 356 2740 364
rect 2780 356 2788 364
rect 2524 336 2532 344
rect 2476 296 2484 304
rect 2492 296 2500 304
rect 2572 316 2580 324
rect 2604 316 2612 324
rect 2556 296 2564 304
rect 2572 296 2580 304
rect 2588 296 2596 304
rect 2332 256 2340 264
rect 2572 256 2580 264
rect 2332 216 2340 224
rect 2524 216 2532 224
rect 2284 196 2292 204
rect 2636 276 2644 284
rect 2620 256 2628 264
rect 2636 256 2644 264
rect 2748 336 2756 344
rect 2956 556 2964 564
rect 3036 536 3044 544
rect 2988 516 2996 524
rect 3180 596 3188 604
rect 3116 556 3124 564
rect 3164 556 3172 564
rect 3196 556 3204 564
rect 3148 516 3156 524
rect 3196 516 3204 524
rect 2876 496 2884 504
rect 2972 496 2980 504
rect 3356 736 3364 744
rect 3372 676 3380 684
rect 3372 656 3380 664
rect 3260 636 3268 644
rect 3404 636 3412 644
rect 3310 606 3318 614
rect 3324 606 3332 614
rect 3338 606 3346 614
rect 3372 576 3380 584
rect 3388 576 3396 584
rect 3260 556 3268 564
rect 3356 556 3364 564
rect 3356 516 3364 524
rect 3340 496 3348 504
rect 3420 596 3428 604
rect 3500 896 3508 904
rect 3468 716 3476 724
rect 3564 876 3572 884
rect 3564 816 3572 824
rect 3548 716 3556 724
rect 3708 1016 3716 1024
rect 3756 1016 3764 1024
rect 3676 976 3684 984
rect 3756 936 3764 944
rect 3788 996 3796 1004
rect 3852 996 3860 1004
rect 3820 976 3828 984
rect 3836 976 3844 984
rect 3596 916 3604 924
rect 3980 1116 3988 1124
rect 4284 1356 4292 1364
rect 4316 1396 4324 1404
rect 4556 1436 4564 1444
rect 4412 1376 4420 1384
rect 4540 1396 4548 1404
rect 4476 1376 4484 1384
rect 4268 1336 4276 1344
rect 4460 1336 4468 1344
rect 4252 1276 4260 1284
rect 4364 1236 4372 1244
rect 4028 1136 4036 1144
rect 4092 1136 4100 1144
rect 4348 1136 4356 1144
rect 4012 1116 4020 1124
rect 4124 1116 4132 1124
rect 4204 1116 4212 1124
rect 4252 1116 4260 1124
rect 3996 1096 4004 1104
rect 3932 1076 3940 1084
rect 4124 1076 4132 1084
rect 3868 916 3876 924
rect 4156 1056 4164 1064
rect 4204 1096 4212 1104
rect 4236 1076 4244 1084
rect 4268 976 4276 984
rect 4124 956 4132 964
rect 4188 956 4196 964
rect 4284 956 4292 964
rect 3948 936 3956 944
rect 3996 916 4004 924
rect 3932 896 3940 904
rect 3996 896 4004 904
rect 4028 936 4036 944
rect 4108 916 4116 924
rect 4428 1316 4436 1324
rect 4492 1316 4500 1324
rect 4428 1136 4436 1144
rect 4396 1076 4404 1084
rect 4652 1496 4660 1504
rect 4700 1556 4708 1564
rect 4764 1636 4772 1644
rect 4830 1606 4838 1614
rect 4844 1606 4852 1614
rect 4858 1606 4866 1614
rect 4924 1596 4932 1604
rect 4860 1576 4868 1584
rect 4876 1576 4884 1584
rect 4972 1576 4980 1584
rect 4844 1556 4852 1564
rect 4796 1516 4804 1524
rect 4780 1496 4788 1504
rect 4796 1476 4804 1484
rect 4636 1456 4644 1464
rect 4588 1396 4596 1404
rect 4860 1496 4868 1504
rect 4764 1436 4772 1444
rect 4668 1376 4676 1384
rect 4716 1416 4724 1424
rect 4812 1376 4820 1384
rect 4684 1356 4692 1364
rect 4620 1336 4628 1344
rect 4700 1336 4708 1344
rect 4860 1336 4868 1344
rect 4556 1316 4564 1324
rect 4604 1316 4612 1324
rect 4668 1316 4676 1324
rect 4556 1276 4564 1284
rect 4636 1276 4644 1284
rect 4940 1556 4948 1564
rect 5020 1556 5028 1564
rect 4924 1516 4932 1524
rect 4972 1516 4980 1524
rect 4908 1476 4916 1484
rect 4956 1476 4964 1484
rect 5084 1616 5092 1624
rect 5036 1516 5044 1524
rect 4924 1456 4932 1464
rect 4988 1416 4996 1424
rect 4988 1396 4996 1404
rect 4956 1356 4964 1364
rect 5020 1356 5028 1364
rect 5068 1536 5076 1544
rect 5164 1536 5172 1544
rect 5100 1516 5108 1524
rect 5084 1496 5092 1504
rect 5148 1516 5156 1524
rect 5132 1496 5140 1504
rect 5212 1696 5220 1704
rect 5228 1696 5236 1704
rect 5308 1696 5316 1704
rect 5180 1496 5188 1504
rect 5260 1576 5268 1584
rect 5276 1576 5284 1584
rect 5228 1536 5236 1544
rect 5276 1556 5284 1564
rect 5244 1516 5252 1524
rect 5260 1516 5268 1524
rect 5260 1476 5268 1484
rect 5148 1456 5156 1464
rect 5132 1396 5140 1404
rect 5068 1336 5076 1344
rect 5116 1336 5124 1344
rect 4876 1316 4884 1324
rect 4844 1276 4852 1284
rect 4748 1256 4756 1264
rect 4492 1136 4500 1144
rect 4524 1136 4532 1144
rect 4476 1116 4484 1124
rect 4604 1156 4612 1164
rect 4636 1136 4644 1144
rect 4588 1116 4596 1124
rect 4830 1206 4838 1214
rect 4844 1206 4852 1214
rect 4858 1206 4866 1214
rect 4716 1136 4724 1144
rect 4476 1096 4484 1104
rect 4524 1096 4532 1104
rect 4556 1096 4564 1104
rect 4652 1096 4660 1104
rect 4508 1056 4516 1064
rect 4556 1056 4564 1064
rect 4348 976 4356 984
rect 4460 976 4468 984
rect 4332 956 4340 964
rect 4412 956 4420 964
rect 4540 1016 4548 1024
rect 4540 956 4548 964
rect 4556 956 4564 964
rect 4620 1056 4628 1064
rect 4652 1056 4660 1064
rect 4700 1096 4708 1104
rect 4972 1256 4980 1264
rect 4956 1176 4964 1184
rect 4908 1096 4916 1104
rect 4972 1136 4980 1144
rect 5036 1276 5044 1284
rect 5132 1276 5140 1284
rect 5004 1116 5012 1124
rect 5084 1116 5092 1124
rect 4988 1096 4996 1104
rect 4828 1076 4836 1084
rect 4668 1036 4676 1044
rect 4716 1036 4724 1044
rect 4748 1036 4756 1044
rect 4668 996 4676 1004
rect 5052 1076 5060 1084
rect 5084 1056 5092 1064
rect 5116 1056 5124 1064
rect 4796 1016 4804 1024
rect 4812 1016 4820 1024
rect 4604 976 4612 984
rect 4812 976 4820 984
rect 4892 976 4900 984
rect 4668 956 4676 964
rect 4684 956 4692 964
rect 4780 956 4788 964
rect 4524 936 4532 944
rect 4588 936 4596 944
rect 4156 916 4164 924
rect 4444 916 4452 924
rect 3596 876 3604 884
rect 4060 876 4068 884
rect 4092 876 4100 884
rect 4140 876 4148 884
rect 3564 676 3572 684
rect 3692 856 3700 864
rect 3660 756 3668 764
rect 3612 716 3620 724
rect 4076 836 4084 844
rect 3804 776 3812 784
rect 3724 756 3732 764
rect 3772 756 3780 764
rect 3676 716 3684 724
rect 3628 676 3636 684
rect 3676 676 3684 684
rect 3884 736 3892 744
rect 3772 716 3780 724
rect 3804 716 3812 724
rect 3932 716 3940 724
rect 3452 656 3460 664
rect 3548 656 3556 664
rect 3596 656 3604 664
rect 3772 676 3780 684
rect 3692 656 3700 664
rect 3884 656 3892 664
rect 3980 656 3988 664
rect 3452 616 3460 624
rect 3468 576 3476 584
rect 3532 576 3540 584
rect 3564 616 3572 624
rect 3596 616 3604 624
rect 3436 536 3444 544
rect 3484 536 3492 544
rect 3532 536 3540 544
rect 3436 496 3444 504
rect 3468 496 3476 504
rect 2860 476 2868 484
rect 3004 476 3012 484
rect 3068 476 3076 484
rect 3244 476 3252 484
rect 3324 476 3332 484
rect 3388 476 3396 484
rect 3420 476 3428 484
rect 2812 456 2820 464
rect 3052 456 3060 464
rect 3244 456 3252 464
rect 2812 436 2820 444
rect 2812 356 2820 364
rect 2860 336 2868 344
rect 2796 316 2804 324
rect 2828 316 2836 324
rect 2940 316 2948 324
rect 2972 316 2980 324
rect 2684 276 2692 284
rect 2716 276 2724 284
rect 3020 376 3028 384
rect 3004 336 3012 344
rect 3116 376 3124 384
rect 3084 336 3092 344
rect 3100 336 3108 344
rect 3052 316 3060 324
rect 2956 276 2964 284
rect 2972 276 2980 284
rect 3644 616 3652 624
rect 3676 616 3684 624
rect 3628 536 3636 544
rect 3644 536 3652 544
rect 3820 636 3828 644
rect 3836 636 3844 644
rect 3916 636 3924 644
rect 3788 616 3796 624
rect 3836 576 3844 584
rect 3884 576 3892 584
rect 3708 556 3716 564
rect 3772 556 3780 564
rect 3820 556 3828 564
rect 3836 556 3844 564
rect 3900 556 3908 564
rect 3916 556 3924 564
rect 3724 536 3732 544
rect 3756 536 3764 544
rect 3820 536 3828 544
rect 3884 536 3892 544
rect 3612 516 3620 524
rect 3628 516 3636 524
rect 3548 496 3556 504
rect 3724 496 3732 504
rect 3788 496 3796 504
rect 3836 496 3844 504
rect 3916 496 3924 504
rect 3852 476 3860 484
rect 3900 476 3908 484
rect 3644 456 3652 464
rect 3708 456 3716 464
rect 3724 456 3732 464
rect 3532 396 3540 404
rect 3292 376 3300 384
rect 3420 376 3428 384
rect 3532 376 3540 384
rect 3580 376 3588 384
rect 3228 356 3236 364
rect 3308 356 3316 364
rect 3468 356 3476 364
rect 3404 336 3412 344
rect 3452 336 3460 344
rect 3596 336 3604 344
rect 3244 316 3252 324
rect 3276 316 3284 324
rect 3388 316 3396 324
rect 3404 316 3412 324
rect 3516 316 3524 324
rect 3596 316 3604 324
rect 3612 316 3620 324
rect 3644 316 3652 324
rect 3484 296 3492 304
rect 3148 276 3156 284
rect 3196 276 3204 284
rect 3292 276 3300 284
rect 3404 276 3412 284
rect 3420 276 3428 284
rect 2876 256 2884 264
rect 2892 256 2900 264
rect 3180 256 3188 264
rect 3372 256 3380 264
rect 2604 236 2612 244
rect 2732 236 2740 244
rect 2636 196 2644 204
rect 2300 156 2308 164
rect 2284 136 2292 144
rect 2348 136 2356 144
rect 2380 136 2388 144
rect 2444 136 2452 144
rect 2524 136 2532 144
rect 1980 96 1988 104
rect 2044 96 2052 104
rect 2076 96 2084 104
rect 2108 96 2116 104
rect 2124 96 2132 104
rect 2268 96 2276 104
rect 1308 56 1316 64
rect 1340 56 1348 64
rect 1644 56 1652 64
rect 1676 56 1684 64
rect 1788 56 1796 64
rect 2092 76 2100 84
rect 2140 76 2148 84
rect 2316 96 2324 104
rect 2428 116 2436 124
rect 2668 216 2676 224
rect 2652 176 2660 184
rect 2668 176 2676 184
rect 2668 136 2676 144
rect 2700 136 2708 144
rect 2492 116 2500 124
rect 2556 116 2564 124
rect 2508 96 2516 104
rect 2636 96 2644 104
rect 2716 116 2724 124
rect 2796 196 2804 204
rect 3036 216 3044 224
rect 3036 196 3044 204
rect 3068 196 3076 204
rect 2892 176 2900 184
rect 2924 176 2932 184
rect 2940 176 2948 184
rect 2892 156 2900 164
rect 2716 96 2724 104
rect 2412 76 2420 84
rect 2476 76 2484 84
rect 2764 76 2772 84
rect 2300 56 2308 64
rect 2364 56 2372 64
rect 2380 56 2388 64
rect 2492 56 2500 64
rect 2748 56 2756 64
rect 2844 76 2852 84
rect 2876 76 2884 84
rect 2828 56 2836 64
rect 2908 56 2916 64
rect 972 36 980 44
rect 1724 36 1732 44
rect 1820 36 1828 44
rect 2428 36 2436 44
rect 2812 36 2820 44
rect 2972 156 2980 164
rect 3004 156 3012 164
rect 3020 156 3028 164
rect 3036 156 3044 164
rect 3212 216 3220 224
rect 3228 216 3236 224
rect 3116 196 3124 204
rect 3212 196 3220 204
rect 3132 176 3140 184
rect 3148 176 3156 184
rect 3084 136 3092 144
rect 2956 76 2964 84
rect 2972 76 2980 84
rect 2956 56 2964 64
rect 3052 36 3060 44
rect 2796 16 2804 24
rect 2940 16 2948 24
rect 2956 16 2964 24
rect 3036 16 3044 24
rect 3310 206 3318 214
rect 3324 206 3332 214
rect 3338 206 3346 214
rect 3356 176 3364 184
rect 3260 116 3268 124
rect 3276 116 3284 124
rect 3628 296 3636 304
rect 3660 296 3668 304
rect 3852 436 3860 444
rect 3948 596 3956 604
rect 3948 556 3956 564
rect 3996 536 4004 544
rect 4108 756 4116 764
rect 4252 896 4260 904
rect 4332 896 4340 904
rect 4508 896 4516 904
rect 4572 876 4580 884
rect 4412 796 4420 804
rect 4652 916 4660 924
rect 4636 876 4644 884
rect 4620 836 4628 844
rect 4332 776 4340 784
rect 4380 776 4388 784
rect 4428 776 4436 784
rect 4156 756 4164 764
rect 4236 756 4244 764
rect 4268 736 4276 744
rect 4204 716 4212 724
rect 4124 696 4132 704
rect 4076 676 4084 684
rect 4124 676 4132 684
rect 4156 676 4164 684
rect 4108 656 4116 664
rect 4028 616 4036 624
rect 4060 616 4068 624
rect 4060 536 4068 544
rect 4012 516 4020 524
rect 4076 516 4084 524
rect 4172 656 4180 664
rect 4172 636 4180 644
rect 3996 496 4004 504
rect 4012 496 4020 504
rect 4108 496 4116 504
rect 3980 476 3988 484
rect 3996 416 4004 424
rect 3724 396 3732 404
rect 3852 396 3860 404
rect 3932 396 3940 404
rect 3756 316 3764 324
rect 3804 316 3812 324
rect 3708 296 3716 304
rect 3692 276 3700 284
rect 3884 356 3892 364
rect 3916 356 3924 364
rect 3948 356 3956 364
rect 3868 316 3876 324
rect 3900 336 3908 344
rect 3820 296 3828 304
rect 3884 296 3892 304
rect 3772 276 3780 284
rect 3804 276 3812 284
rect 3964 336 3972 344
rect 4044 476 4052 484
rect 4060 456 4068 464
rect 4028 356 4036 364
rect 4028 316 4036 324
rect 3948 296 3956 304
rect 4012 296 4020 304
rect 4220 676 4228 684
rect 4252 676 4260 684
rect 4364 736 4372 744
rect 4396 756 4404 764
rect 4348 676 4356 684
rect 4364 616 4372 624
rect 4316 576 4324 584
rect 4316 556 4324 564
rect 4364 556 4372 564
rect 4268 536 4276 544
rect 4220 516 4228 524
rect 4284 516 4292 524
rect 4460 736 4468 744
rect 4588 736 4596 744
rect 4540 696 4548 704
rect 4460 656 4468 664
rect 4508 656 4516 664
rect 4524 636 4532 644
rect 4476 596 4484 604
rect 4412 576 4420 584
rect 4332 536 4340 544
rect 4524 556 4532 564
rect 4556 676 4564 684
rect 4572 656 4580 664
rect 4604 616 4612 624
rect 4652 796 4660 804
rect 4636 736 4644 744
rect 4732 936 4740 944
rect 4764 916 4772 924
rect 4700 896 4708 904
rect 4732 896 4740 904
rect 5100 1036 5108 1044
rect 5100 996 5108 1004
rect 5020 976 5028 984
rect 5132 976 5140 984
rect 4908 936 4916 944
rect 4924 936 4932 944
rect 5036 936 5044 944
rect 5068 936 5076 944
rect 5132 936 5140 944
rect 5212 1356 5220 1364
rect 5212 1336 5220 1344
rect 5196 1316 5204 1324
rect 5292 1516 5300 1524
rect 5260 1396 5268 1404
rect 5276 1396 5284 1404
rect 5388 1676 5396 1684
rect 5340 1616 5348 1624
rect 5372 1596 5380 1604
rect 5324 1496 5332 1504
rect 5644 1876 5652 1884
rect 5740 1876 5748 1884
rect 5564 1856 5572 1864
rect 5676 1856 5684 1864
rect 5708 1856 5716 1864
rect 5820 2236 5828 2244
rect 5964 2196 5972 2204
rect 5948 2156 5956 2164
rect 6028 3096 6036 3104
rect 6060 3116 6068 3124
rect 6140 3296 6148 3304
rect 6156 3296 6164 3304
rect 6124 3256 6132 3264
rect 6108 3136 6116 3144
rect 6076 3096 6084 3104
rect 6044 3076 6052 3084
rect 6076 3036 6084 3044
rect 6028 3016 6036 3024
rect 6012 2996 6020 3004
rect 6044 2976 6052 2984
rect 6028 2936 6036 2944
rect 6060 2936 6068 2944
rect 6092 3016 6100 3024
rect 6012 2916 6020 2924
rect 6108 2936 6116 2944
rect 6332 3856 6340 3864
rect 6364 3836 6372 3844
rect 6348 3816 6356 3824
rect 6380 3796 6388 3804
rect 6332 3736 6340 3744
rect 6364 3736 6372 3744
rect 6380 3736 6388 3744
rect 6316 3716 6324 3724
rect 6348 3716 6356 3724
rect 6268 3676 6276 3684
rect 6284 3676 6292 3684
rect 6316 3676 6324 3684
rect 6300 3656 6308 3664
rect 6284 3636 6292 3644
rect 6252 3576 6260 3584
rect 6204 3456 6212 3464
rect 6220 3336 6228 3344
rect 6268 3536 6276 3544
rect 6316 3596 6324 3604
rect 6332 3576 6340 3584
rect 6332 3556 6340 3564
rect 6348 3536 6356 3544
rect 6412 4016 6420 4024
rect 6444 3976 6452 3984
rect 6444 3936 6452 3944
rect 6428 3916 6436 3924
rect 6412 3856 6420 3864
rect 6428 3796 6436 3804
rect 6428 3736 6436 3744
rect 6412 3676 6420 3684
rect 6396 3616 6404 3624
rect 6380 3556 6388 3564
rect 6300 3436 6308 3444
rect 6284 3396 6292 3404
rect 6220 3296 6228 3304
rect 6204 3276 6212 3284
rect 6284 3276 6292 3284
rect 6188 3256 6196 3264
rect 6236 3236 6244 3244
rect 6172 3196 6180 3204
rect 6140 3136 6148 3144
rect 6156 3116 6164 3124
rect 6172 3116 6180 3124
rect 6268 3216 6276 3224
rect 6316 3356 6324 3364
rect 6316 3216 6324 3224
rect 6300 3176 6308 3184
rect 6268 3116 6276 3124
rect 6156 3076 6164 3084
rect 6188 3076 6196 3084
rect 6156 2996 6164 3004
rect 6188 2816 6196 2824
rect 6252 2836 6260 2844
rect 6220 2776 6228 2784
rect 6252 2776 6260 2784
rect 6124 2756 6132 2764
rect 6076 2716 6084 2724
rect 6012 2676 6020 2684
rect 6028 2576 6036 2584
rect 6092 2576 6100 2584
rect 6012 2316 6020 2324
rect 6108 2296 6116 2304
rect 6012 2196 6020 2204
rect 5868 2096 5876 2104
rect 5916 2096 5924 2104
rect 5932 1956 5940 1964
rect 5948 1936 5956 1944
rect 5788 1916 5796 1924
rect 5804 1916 5812 1924
rect 5868 1916 5876 1924
rect 5932 1916 5940 1924
rect 5852 1896 5860 1904
rect 5932 1896 5940 1904
rect 5612 1836 5620 1844
rect 5708 1816 5716 1824
rect 5564 1776 5572 1784
rect 5660 1736 5668 1744
rect 5532 1556 5540 1564
rect 5404 1536 5412 1544
rect 5356 1476 5364 1484
rect 5340 1396 5348 1404
rect 5436 1436 5444 1444
rect 5340 1356 5348 1364
rect 5180 1276 5188 1284
rect 5260 1176 5268 1184
rect 5244 1116 5252 1124
rect 5228 1096 5236 1104
rect 5244 1096 5252 1104
rect 5212 1076 5220 1084
rect 5484 1456 5492 1464
rect 5468 1396 5476 1404
rect 5692 1716 5700 1724
rect 5676 1676 5684 1684
rect 5628 1596 5636 1604
rect 5628 1556 5636 1564
rect 5644 1536 5652 1544
rect 5628 1496 5636 1504
rect 5644 1496 5652 1504
rect 5564 1476 5572 1484
rect 5628 1476 5636 1484
rect 5660 1476 5668 1484
rect 5676 1476 5684 1484
rect 5596 1456 5604 1464
rect 5548 1436 5556 1444
rect 5644 1436 5652 1444
rect 5660 1436 5668 1444
rect 5500 1376 5508 1384
rect 5612 1396 5620 1404
rect 5580 1356 5588 1364
rect 5324 1336 5332 1344
rect 5404 1336 5412 1344
rect 5308 1316 5316 1324
rect 5372 1276 5380 1284
rect 5548 1336 5556 1344
rect 5564 1336 5572 1344
rect 5436 1316 5444 1324
rect 5484 1316 5492 1324
rect 5500 1276 5508 1284
rect 5532 1276 5540 1284
rect 5548 1276 5556 1284
rect 5420 1256 5428 1264
rect 5516 1196 5524 1204
rect 5308 1176 5316 1184
rect 5292 1156 5300 1164
rect 5356 1156 5364 1164
rect 5420 1156 5428 1164
rect 5324 1096 5332 1104
rect 5340 1096 5348 1104
rect 5292 1076 5300 1084
rect 5324 1076 5332 1084
rect 5372 1076 5380 1084
rect 5276 1056 5284 1064
rect 5308 1056 5316 1064
rect 5180 1036 5188 1044
rect 4956 916 4964 924
rect 5004 916 5012 924
rect 5036 916 5044 924
rect 5148 916 5156 924
rect 4956 896 4964 904
rect 5116 896 5124 904
rect 5020 876 5028 884
rect 4924 856 4932 864
rect 4830 806 4838 814
rect 4844 806 4852 814
rect 4858 806 4866 814
rect 4732 796 4740 804
rect 5148 896 5156 904
rect 5132 856 5140 864
rect 5276 996 5284 1004
rect 5228 956 5236 964
rect 5276 956 5284 964
rect 5260 936 5268 944
rect 5292 936 5300 944
rect 5180 916 5188 924
rect 5196 916 5204 924
rect 5228 916 5236 924
rect 5292 856 5300 864
rect 4972 736 4980 744
rect 5036 736 5044 744
rect 5068 736 5076 744
rect 4796 716 4804 724
rect 4716 696 4724 704
rect 4700 676 4708 684
rect 4684 636 4692 644
rect 4732 676 4740 684
rect 4908 716 4916 724
rect 4956 716 4964 724
rect 5020 716 5028 724
rect 5100 716 5108 724
rect 4988 696 4996 704
rect 5004 696 5012 704
rect 4844 676 4852 684
rect 4908 676 4916 684
rect 4780 656 4788 664
rect 4748 636 4756 644
rect 4780 636 4788 644
rect 4828 636 4836 644
rect 4812 616 4820 624
rect 4828 616 4836 624
rect 4796 596 4804 604
rect 4652 556 4660 564
rect 4684 556 4692 564
rect 4764 556 4772 564
rect 4556 536 4564 544
rect 4668 536 4676 544
rect 4348 516 4356 524
rect 4140 496 4148 504
rect 4188 496 4196 504
rect 4252 496 4260 504
rect 4380 496 4388 504
rect 4268 476 4276 484
rect 4124 456 4132 464
rect 4156 456 4164 464
rect 4092 436 4100 444
rect 4108 436 4116 444
rect 4076 296 4084 304
rect 4124 336 4132 344
rect 4124 316 4132 324
rect 4172 436 4180 444
rect 4348 376 4356 384
rect 4220 356 4228 364
rect 4300 356 4308 364
rect 4252 316 4260 324
rect 4428 496 4436 504
rect 4412 476 4420 484
rect 4412 416 4420 424
rect 4396 356 4404 364
rect 4380 316 4388 324
rect 4492 496 4500 504
rect 4460 416 4468 424
rect 4428 336 4436 344
rect 4444 336 4452 344
rect 4140 296 4148 304
rect 4188 296 4196 304
rect 4236 296 4244 304
rect 4268 296 4276 304
rect 4332 296 4340 304
rect 4476 316 4484 324
rect 3932 276 3940 284
rect 4108 276 4116 284
rect 4236 276 4244 284
rect 4332 276 4340 284
rect 3692 256 3700 264
rect 3756 256 3764 264
rect 3916 256 3924 264
rect 3612 236 3620 244
rect 3772 236 3780 244
rect 3468 196 3476 204
rect 3516 176 3524 184
rect 3436 156 3444 164
rect 3404 116 3412 124
rect 3436 116 3444 124
rect 3420 96 3428 104
rect 3500 96 3508 104
rect 3580 196 3588 204
rect 3628 156 3636 164
rect 3660 156 3668 164
rect 3644 136 3652 144
rect 3708 136 3716 144
rect 3564 96 3572 104
rect 3628 96 3636 104
rect 3388 76 3396 84
rect 3420 76 3428 84
rect 3452 76 3460 84
rect 3484 76 3492 84
rect 3548 76 3556 84
rect 3564 76 3572 84
rect 3788 216 3796 224
rect 3804 216 3812 224
rect 3868 216 3876 224
rect 3884 156 3892 164
rect 3788 136 3796 144
rect 3868 136 3876 144
rect 3756 116 3764 124
rect 3820 116 3828 124
rect 3772 96 3780 104
rect 4540 416 4548 424
rect 4524 356 4532 364
rect 4508 336 4516 344
rect 4556 376 4564 384
rect 4812 556 4820 564
rect 5036 656 5044 664
rect 4924 636 4932 644
rect 4908 556 4916 564
rect 4748 516 4756 524
rect 4828 516 4836 524
rect 4924 516 4932 524
rect 5164 696 5172 704
rect 5228 696 5236 704
rect 5436 1136 5444 1144
rect 5484 1136 5492 1144
rect 5500 1116 5508 1124
rect 5436 1076 5444 1084
rect 5420 1016 5428 1024
rect 5452 1016 5460 1024
rect 5388 996 5396 1004
rect 5436 996 5444 1004
rect 5372 976 5380 984
rect 5404 936 5412 944
rect 5484 1016 5492 1024
rect 5500 1016 5508 1024
rect 5484 996 5492 1004
rect 5500 976 5508 984
rect 5468 916 5476 924
rect 5468 756 5476 764
rect 5532 1136 5540 1144
rect 5532 1076 5540 1084
rect 5660 1336 5668 1344
rect 5580 1316 5588 1324
rect 5676 1316 5684 1324
rect 5580 1256 5588 1264
rect 5644 1256 5652 1264
rect 5628 1136 5636 1144
rect 5532 1016 5540 1024
rect 5612 1076 5620 1084
rect 5596 956 5604 964
rect 5548 916 5556 924
rect 5612 916 5620 924
rect 5660 1096 5668 1104
rect 5724 1776 5732 1784
rect 5932 1856 5940 1864
rect 5820 1836 5828 1844
rect 5884 1836 5892 1844
rect 5836 1796 5844 1804
rect 5724 1756 5732 1764
rect 5756 1756 5764 1764
rect 5772 1756 5780 1764
rect 5900 1756 5908 1764
rect 5916 1756 5924 1764
rect 5836 1736 5844 1744
rect 5740 1716 5748 1724
rect 5788 1716 5796 1724
rect 5804 1716 5812 1724
rect 5852 1716 5860 1724
rect 5932 1736 5940 1744
rect 5884 1696 5892 1704
rect 5772 1676 5780 1684
rect 5820 1676 5828 1684
rect 5900 1636 5908 1644
rect 5740 1516 5748 1524
rect 5804 1516 5812 1524
rect 5756 1496 5764 1504
rect 5772 1496 5780 1504
rect 5788 1476 5796 1484
rect 5836 1476 5844 1484
rect 5820 1456 5828 1464
rect 5836 1456 5844 1464
rect 5772 1436 5780 1444
rect 5788 1436 5796 1444
rect 5756 1336 5764 1344
rect 5724 1216 5732 1224
rect 5724 1096 5732 1104
rect 5724 1076 5732 1084
rect 5708 1016 5716 1024
rect 5724 996 5732 1004
rect 5708 976 5716 984
rect 5660 956 5668 964
rect 5772 1076 5780 1084
rect 5932 1496 5940 1504
rect 5900 1476 5908 1484
rect 5916 1456 5924 1464
rect 5884 1436 5892 1444
rect 5884 1416 5892 1424
rect 5868 1396 5876 1404
rect 5852 1376 5860 1384
rect 5868 1376 5876 1384
rect 5804 1356 5812 1364
rect 5820 1336 5828 1344
rect 5852 1336 5860 1344
rect 5932 1396 5940 1404
rect 5996 2116 6004 2124
rect 6060 2136 6068 2144
rect 6076 2116 6084 2124
rect 6076 1996 6084 2004
rect 6028 1976 6036 1984
rect 5980 1936 5988 1944
rect 5996 1896 6004 1904
rect 6012 1876 6020 1884
rect 6076 1856 6084 1864
rect 6060 1836 6068 1844
rect 5980 1816 5988 1824
rect 6108 1816 6116 1824
rect 6092 1796 6100 1804
rect 5980 1776 5988 1784
rect 6012 1756 6020 1764
rect 6044 1756 6052 1764
rect 6108 1756 6116 1764
rect 6012 1716 6020 1724
rect 6028 1696 6036 1704
rect 6140 2696 6148 2704
rect 6172 2696 6180 2704
rect 6204 2676 6212 2684
rect 6236 2596 6244 2604
rect 6204 2516 6212 2524
rect 6220 2496 6228 2504
rect 6348 3496 6356 3504
rect 6364 3496 6372 3504
rect 6396 3476 6404 3484
rect 6348 3456 6356 3464
rect 6476 4156 6484 4164
rect 6476 4116 6484 4124
rect 6524 4316 6532 4324
rect 6540 4316 6548 4324
rect 6524 4276 6532 4284
rect 6540 4276 6548 4284
rect 6524 4256 6532 4264
rect 6524 4156 6532 4164
rect 6508 4096 6516 4104
rect 6556 4256 6564 4264
rect 6556 4176 6564 4184
rect 6556 4136 6564 4144
rect 6716 4756 6724 4764
rect 6620 4736 6628 4744
rect 6588 4316 6596 4324
rect 6604 4296 6612 4304
rect 6716 4696 6724 4704
rect 6636 4536 6644 4544
rect 6636 4276 6644 4284
rect 6636 4256 6644 4264
rect 6620 4236 6628 4244
rect 6588 4196 6596 4204
rect 6588 4096 6596 4104
rect 6572 4056 6580 4064
rect 6540 4036 6548 4044
rect 6556 3996 6564 4004
rect 6476 3936 6484 3944
rect 6540 3936 6548 3944
rect 6492 3916 6500 3924
rect 6476 3896 6484 3904
rect 6524 3896 6532 3904
rect 6588 3936 6596 3944
rect 6572 3896 6580 3904
rect 6508 3876 6516 3884
rect 6540 3876 6548 3884
rect 6556 3876 6564 3884
rect 6476 3856 6484 3864
rect 6460 3656 6468 3664
rect 6572 3836 6580 3844
rect 6540 3816 6548 3824
rect 6604 3896 6612 3904
rect 6604 3876 6612 3884
rect 6620 3796 6628 3804
rect 6620 3776 6628 3784
rect 6604 3756 6612 3764
rect 6604 3736 6612 3744
rect 6604 3716 6612 3724
rect 6492 3656 6500 3664
rect 6476 3636 6484 3644
rect 6460 3536 6468 3544
rect 6524 3636 6532 3644
rect 6508 3596 6516 3604
rect 6428 3496 6436 3504
rect 6412 3436 6420 3444
rect 6572 3576 6580 3584
rect 6556 3516 6564 3524
rect 6588 3536 6596 3544
rect 6524 3496 6532 3504
rect 6556 3496 6564 3504
rect 6572 3496 6580 3504
rect 6492 3456 6500 3464
rect 6540 3456 6548 3464
rect 6460 3416 6468 3424
rect 6476 3416 6484 3424
rect 6428 3356 6436 3364
rect 6540 3416 6548 3424
rect 6524 3336 6532 3344
rect 6348 3316 6356 3324
rect 6428 3296 6436 3304
rect 6364 3216 6372 3224
rect 6348 3096 6356 3104
rect 6380 3176 6388 3184
rect 6380 3036 6388 3044
rect 6332 3016 6340 3024
rect 6444 3216 6452 3224
rect 6444 3136 6452 3144
rect 6508 3216 6516 3224
rect 6492 3176 6500 3184
rect 6460 3116 6468 3124
rect 6476 3056 6484 3064
rect 6476 3036 6484 3044
rect 6380 2936 6388 2944
rect 6508 3136 6516 3144
rect 6572 3456 6580 3464
rect 6556 3136 6564 3144
rect 6620 3696 6628 3704
rect 6620 3616 6628 3624
rect 6604 3456 6612 3464
rect 6620 3296 6628 3304
rect 6620 3156 6628 3164
rect 6604 3136 6612 3144
rect 6572 3096 6580 3104
rect 6588 3096 6596 3104
rect 6620 3096 6628 3104
rect 6524 3056 6532 3064
rect 6508 3036 6516 3044
rect 6508 3016 6516 3024
rect 6492 2996 6500 3004
rect 6460 2976 6468 2984
rect 6492 2976 6500 2984
rect 6444 2936 6452 2944
rect 6428 2896 6436 2904
rect 6364 2776 6372 2784
rect 6396 2776 6404 2784
rect 6492 2776 6500 2784
rect 6380 2716 6388 2724
rect 6444 2676 6452 2684
rect 6268 2636 6276 2644
rect 6476 2518 6484 2524
rect 6476 2516 6484 2518
rect 6284 2496 6292 2504
rect 6476 2436 6484 2444
rect 6140 2336 6148 2344
rect 6156 2316 6164 2324
rect 6188 2296 6196 2304
rect 6364 2356 6372 2364
rect 6412 2356 6420 2364
rect 6140 2256 6148 2264
rect 6204 2256 6212 2264
rect 6236 2236 6244 2244
rect 6220 2216 6228 2224
rect 6172 2176 6180 2184
rect 6156 2156 6164 2164
rect 6204 2116 6212 2124
rect 6172 2096 6180 2104
rect 6204 2056 6212 2064
rect 6156 1876 6164 1884
rect 6140 1756 6148 1764
rect 6140 1716 6148 1724
rect 6188 1716 6196 1724
rect 6156 1696 6164 1704
rect 6172 1696 6180 1704
rect 6060 1676 6068 1684
rect 6108 1676 6116 1684
rect 6124 1676 6132 1684
rect 6156 1676 6164 1684
rect 6172 1676 6180 1684
rect 5964 1636 5972 1644
rect 6060 1636 6068 1644
rect 6044 1616 6052 1624
rect 6028 1576 6036 1584
rect 5964 1556 5972 1564
rect 5980 1536 5988 1544
rect 6012 1496 6020 1504
rect 6044 1536 6052 1544
rect 6076 1556 6084 1564
rect 6060 1496 6068 1504
rect 5980 1476 5988 1484
rect 6076 1476 6084 1484
rect 5996 1456 6004 1464
rect 6060 1416 6068 1424
rect 5996 1396 6004 1404
rect 5948 1376 5956 1384
rect 5980 1376 5988 1384
rect 5804 1316 5812 1324
rect 5868 1316 5876 1324
rect 5884 1276 5892 1284
rect 5948 1356 5956 1364
rect 5948 1336 5956 1344
rect 5916 1176 5924 1184
rect 5900 1116 5908 1124
rect 5820 1096 5828 1104
rect 5884 1096 5892 1104
rect 5788 1056 5796 1064
rect 5820 1056 5828 1064
rect 5852 1056 5860 1064
rect 5884 1056 5892 1064
rect 5788 976 5796 984
rect 5740 956 5748 964
rect 5724 936 5732 944
rect 5868 936 5876 944
rect 5676 916 5684 924
rect 5676 896 5684 904
rect 5740 896 5748 904
rect 5868 896 5876 904
rect 5708 856 5716 864
rect 5644 816 5652 824
rect 5740 836 5748 844
rect 5548 716 5556 724
rect 5644 716 5652 724
rect 5372 696 5380 704
rect 5404 696 5412 704
rect 5420 696 5428 704
rect 5516 696 5524 704
rect 5260 676 5268 684
rect 5372 676 5380 684
rect 5116 656 5124 664
rect 5212 656 5220 664
rect 5308 656 5316 664
rect 5084 616 5092 624
rect 5132 596 5140 604
rect 5068 576 5076 584
rect 5084 576 5092 584
rect 5004 536 5012 544
rect 4940 496 4948 504
rect 4956 496 4964 504
rect 5004 496 5012 504
rect 4700 436 4708 444
rect 4828 436 4836 444
rect 4684 376 4692 384
rect 4588 336 4596 344
rect 4652 336 4660 344
rect 4556 316 4564 324
rect 4572 296 4580 304
rect 4652 276 4660 284
rect 3996 256 4004 264
rect 4092 256 4100 264
rect 4124 256 4132 264
rect 4540 256 4548 264
rect 3948 216 3956 224
rect 3932 176 3940 184
rect 3916 116 3924 124
rect 4156 236 4164 244
rect 4204 236 4212 244
rect 3996 176 4004 184
rect 3980 136 3988 144
rect 4156 136 4164 144
rect 4476 216 4484 224
rect 4428 156 4436 164
rect 4684 176 4692 184
rect 4668 156 4676 164
rect 4764 276 4772 284
rect 4830 406 4838 414
rect 4844 406 4852 414
rect 4858 406 4866 414
rect 4876 316 4884 324
rect 4796 296 4804 304
rect 4716 256 4724 264
rect 4780 256 4788 264
rect 4844 236 4852 244
rect 4796 176 4804 184
rect 5116 536 5124 544
rect 5132 536 5140 544
rect 5052 496 5060 504
rect 5052 456 5060 464
rect 4956 296 4964 304
rect 4924 256 4932 264
rect 5004 236 5012 244
rect 5036 176 5044 184
rect 4972 156 4980 164
rect 5100 376 5108 384
rect 5068 316 5076 324
rect 5180 616 5188 624
rect 5212 556 5220 564
rect 5308 556 5316 564
rect 5292 536 5300 544
rect 5132 496 5140 504
rect 5180 456 5188 464
rect 5372 596 5380 604
rect 5500 676 5508 684
rect 5452 656 5460 664
rect 5340 556 5348 564
rect 5388 536 5396 544
rect 5244 436 5252 444
rect 5292 436 5300 444
rect 5116 296 5124 304
rect 5148 276 5156 284
rect 5180 316 5188 324
rect 5212 316 5220 324
rect 5228 296 5236 304
rect 5244 296 5252 304
rect 5516 616 5524 624
rect 5420 576 5428 584
rect 5500 576 5508 584
rect 5484 556 5492 564
rect 5644 676 5652 684
rect 5772 716 5780 724
rect 5884 856 5892 864
rect 5820 716 5828 724
rect 5804 696 5812 704
rect 5836 696 5844 704
rect 5756 676 5764 684
rect 5788 676 5796 684
rect 5676 656 5684 664
rect 5804 636 5812 644
rect 5660 616 5668 624
rect 5788 616 5796 624
rect 5612 556 5620 564
rect 5564 536 5572 544
rect 5596 536 5604 544
rect 5740 556 5748 564
rect 5804 556 5812 564
rect 5708 536 5716 544
rect 5596 516 5604 524
rect 5660 516 5668 524
rect 5692 516 5700 524
rect 5740 516 5748 524
rect 5548 476 5556 484
rect 5580 476 5588 484
rect 5404 456 5412 464
rect 5676 496 5684 504
rect 5724 496 5732 504
rect 5756 496 5764 504
rect 5644 476 5652 484
rect 5660 416 5668 424
rect 5852 636 5860 644
rect 5868 576 5876 584
rect 5964 1316 5972 1324
rect 5932 1096 5940 1104
rect 6028 1376 6036 1384
rect 6012 1316 6020 1324
rect 5996 1196 6004 1204
rect 5980 1116 5988 1124
rect 5980 1096 5988 1104
rect 5980 1076 5988 1084
rect 5964 1036 5972 1044
rect 5964 936 5972 944
rect 5932 916 5940 924
rect 5980 916 5988 924
rect 5948 896 5956 904
rect 6044 1356 6052 1364
rect 6076 1316 6084 1324
rect 6076 1216 6084 1224
rect 6044 1156 6052 1164
rect 6076 1156 6084 1164
rect 6028 1096 6036 1104
rect 6060 1116 6068 1124
rect 6060 1096 6068 1104
rect 6060 1036 6068 1044
rect 6076 1036 6084 1044
rect 6108 1516 6116 1524
rect 6140 1516 6148 1524
rect 6124 1496 6132 1504
rect 6124 1476 6132 1484
rect 6268 2176 6276 2184
rect 6332 2176 6340 2184
rect 6284 2116 6292 2124
rect 6332 2116 6340 2124
rect 6236 2096 6244 2104
rect 6300 2096 6308 2104
rect 6316 2096 6324 2104
rect 6460 2256 6468 2264
rect 6428 2236 6436 2244
rect 6396 2216 6404 2224
rect 6412 2176 6420 2184
rect 6460 2136 6468 2144
rect 6428 2116 6436 2124
rect 6460 2116 6468 2124
rect 6380 2096 6388 2104
rect 6396 2096 6404 2104
rect 6444 2096 6452 2104
rect 6444 2076 6452 2084
rect 6364 2056 6372 2064
rect 6220 2016 6228 2024
rect 6428 1936 6436 1944
rect 6252 1916 6260 1924
rect 6300 1916 6308 1924
rect 6332 1916 6340 1924
rect 6412 1916 6420 1924
rect 6348 1896 6356 1904
rect 6428 1896 6436 1904
rect 6220 1876 6228 1884
rect 6220 1736 6228 1744
rect 6268 1836 6276 1844
rect 6300 1756 6308 1764
rect 6268 1736 6276 1744
rect 6252 1716 6260 1724
rect 6236 1696 6244 1704
rect 6172 1556 6180 1564
rect 6172 1496 6180 1504
rect 6108 1436 6116 1444
rect 6124 1396 6132 1404
rect 6108 1356 6116 1364
rect 6156 1416 6164 1424
rect 6236 1636 6244 1644
rect 6284 1696 6292 1704
rect 6348 1816 6356 1824
rect 6380 1816 6388 1824
rect 6364 1796 6372 1804
rect 6380 1776 6388 1784
rect 6364 1756 6372 1764
rect 6316 1676 6324 1684
rect 6236 1616 6244 1624
rect 6268 1616 6276 1624
rect 6220 1576 6228 1584
rect 6204 1516 6212 1524
rect 6204 1456 6212 1464
rect 6188 1376 6196 1384
rect 6172 1356 6180 1364
rect 6172 1336 6180 1344
rect 6156 1296 6164 1304
rect 6140 1256 6148 1264
rect 6124 1216 6132 1224
rect 6108 1136 6116 1144
rect 6188 1276 6196 1284
rect 6220 1416 6228 1424
rect 6204 1236 6212 1244
rect 6268 1596 6276 1604
rect 6332 1536 6340 1544
rect 6348 1536 6356 1544
rect 6428 1736 6436 1744
rect 6588 3036 6596 3044
rect 6604 3036 6612 3044
rect 6540 2876 6548 2884
rect 6508 2236 6516 2244
rect 6492 2156 6500 2164
rect 6572 3016 6580 3024
rect 6556 2776 6564 2784
rect 6716 3216 6724 3224
rect 6716 3196 6724 3204
rect 6636 3016 6644 3024
rect 6620 2996 6628 3004
rect 6636 2936 6644 2944
rect 6636 2856 6644 2864
rect 6636 2716 6644 2724
rect 6620 2656 6628 2664
rect 6540 2576 6548 2584
rect 6604 2576 6612 2584
rect 6588 2236 6596 2244
rect 6540 2216 6548 2224
rect 6524 2136 6532 2144
rect 6524 2116 6532 2124
rect 6508 1996 6516 2004
rect 6524 1976 6532 1984
rect 6556 2096 6564 2104
rect 6572 2076 6580 2084
rect 6556 1976 6564 1984
rect 6540 1956 6548 1964
rect 6540 1936 6548 1944
rect 6460 1916 6468 1924
rect 6508 1916 6516 1924
rect 6524 1916 6532 1924
rect 6460 1896 6468 1904
rect 6476 1896 6484 1904
rect 6540 1896 6548 1904
rect 6460 1736 6468 1744
rect 6492 1736 6500 1744
rect 6524 1736 6532 1744
rect 6572 1956 6580 1964
rect 6396 1716 6404 1724
rect 6444 1716 6452 1724
rect 6524 1716 6532 1724
rect 6444 1696 6452 1704
rect 6476 1696 6484 1704
rect 6412 1676 6420 1684
rect 6460 1636 6468 1644
rect 6412 1576 6420 1584
rect 6396 1556 6404 1564
rect 6252 1516 6260 1524
rect 6284 1516 6292 1524
rect 6364 1516 6372 1524
rect 6396 1516 6404 1524
rect 6268 1496 6276 1504
rect 6332 1496 6340 1504
rect 6396 1496 6404 1504
rect 6380 1476 6388 1484
rect 6332 1456 6340 1464
rect 6364 1456 6372 1464
rect 6268 1396 6276 1404
rect 6332 1356 6340 1364
rect 6268 1316 6276 1324
rect 6172 1216 6180 1224
rect 6156 1176 6164 1184
rect 6204 1136 6212 1144
rect 6140 1096 6148 1104
rect 6188 1096 6196 1104
rect 6108 1076 6116 1084
rect 6156 1076 6164 1084
rect 6124 1056 6132 1064
rect 6204 1036 6212 1044
rect 6204 1016 6212 1024
rect 6044 976 6052 984
rect 6060 976 6068 984
rect 6092 976 6100 984
rect 6124 976 6132 984
rect 6188 976 6196 984
rect 6028 936 6036 944
rect 6044 916 6052 924
rect 5996 876 6004 884
rect 5964 856 5972 864
rect 5980 756 5988 764
rect 6108 916 6116 924
rect 6092 896 6100 904
rect 6172 936 6180 944
rect 6156 916 6164 924
rect 6156 896 6164 904
rect 5932 736 5940 744
rect 5964 736 5972 744
rect 6012 736 6020 744
rect 6076 816 6084 824
rect 5980 716 5988 724
rect 6044 716 6052 724
rect 5996 696 6004 704
rect 5932 676 5940 684
rect 5964 676 5972 684
rect 6028 696 6036 704
rect 6044 676 6052 684
rect 5916 616 5924 624
rect 5900 556 5908 564
rect 5836 536 5844 544
rect 5916 536 5924 544
rect 5916 516 5924 524
rect 5884 496 5892 504
rect 5788 376 5796 384
rect 5836 376 5844 384
rect 5740 356 5748 364
rect 5404 336 5412 344
rect 5452 336 5460 344
rect 5628 336 5636 344
rect 5388 296 5396 304
rect 5212 276 5220 284
rect 5276 276 5284 284
rect 5308 276 5316 284
rect 5372 276 5380 284
rect 5084 256 5092 264
rect 5276 256 5284 264
rect 5340 256 5348 264
rect 5356 256 5364 264
rect 4620 136 4628 144
rect 4972 136 4980 144
rect 5020 136 5028 144
rect 5052 136 5060 144
rect 4396 118 4404 124
rect 4396 116 4404 118
rect 4636 118 4644 124
rect 4636 116 4644 118
rect 4764 116 4772 124
rect 4908 116 4916 124
rect 4988 116 4996 124
rect 5052 116 5060 124
rect 3916 96 3924 104
rect 3948 96 3956 104
rect 4012 96 4020 104
rect 3836 76 3844 84
rect 3900 76 3908 84
rect 4892 96 4900 104
rect 5036 96 5044 104
rect 5100 96 5108 104
rect 5612 276 5620 284
rect 5660 276 5668 284
rect 5596 256 5604 264
rect 5676 236 5684 244
rect 5724 236 5732 244
rect 5308 156 5316 164
rect 5420 156 5428 164
rect 5516 156 5524 164
rect 5628 216 5636 224
rect 5820 336 5828 344
rect 5852 336 5860 344
rect 6012 636 6020 644
rect 5948 536 5956 544
rect 6060 536 6068 544
rect 5948 496 5956 504
rect 6108 796 6116 804
rect 6188 896 6196 904
rect 6172 776 6180 784
rect 6108 756 6116 764
rect 6172 756 6180 764
rect 6124 716 6132 724
rect 6188 716 6196 724
rect 6156 676 6164 684
rect 6124 656 6132 664
rect 6092 616 6100 624
rect 5980 516 5988 524
rect 6076 516 6084 524
rect 6076 496 6084 504
rect 6140 616 6148 624
rect 6140 556 6148 564
rect 5964 476 5972 484
rect 6012 476 6020 484
rect 5916 456 5924 464
rect 5932 456 5940 464
rect 5884 336 5892 344
rect 5772 296 5780 304
rect 5804 296 5812 304
rect 5868 296 5876 304
rect 5772 276 5780 284
rect 5788 276 5796 284
rect 5836 256 5844 264
rect 5660 176 5668 184
rect 5740 176 5748 184
rect 5788 156 5796 164
rect 5996 416 6004 424
rect 6028 376 6036 384
rect 5932 316 5940 324
rect 6092 376 6100 384
rect 6076 336 6084 344
rect 6060 316 6068 324
rect 6076 296 6084 304
rect 5900 276 5908 284
rect 5916 276 5924 284
rect 6124 416 6132 424
rect 6124 316 6132 324
rect 5964 256 5972 264
rect 6012 256 6020 264
rect 6060 256 6068 264
rect 6012 236 6020 244
rect 6124 236 6132 244
rect 6076 216 6084 224
rect 6076 196 6084 204
rect 6172 576 6180 584
rect 6156 496 6164 504
rect 6236 1216 6244 1224
rect 6220 956 6228 964
rect 6252 1176 6260 1184
rect 6252 1156 6260 1164
rect 6348 1316 6356 1324
rect 6444 1516 6452 1524
rect 6428 1476 6436 1484
rect 6284 1276 6292 1284
rect 6284 1216 6292 1224
rect 6332 1236 6340 1244
rect 6316 1216 6324 1224
rect 6284 1116 6292 1124
rect 6284 1096 6292 1104
rect 6380 1296 6388 1304
rect 6364 1276 6372 1284
rect 6412 1336 6420 1344
rect 6428 1316 6436 1324
rect 6444 1296 6452 1304
rect 6412 1276 6420 1284
rect 6508 1676 6516 1684
rect 6540 1596 6548 1604
rect 6476 1536 6484 1544
rect 6492 1536 6500 1544
rect 6524 1516 6532 1524
rect 6588 1936 6596 1944
rect 6588 1916 6596 1924
rect 6588 1636 6596 1644
rect 6588 1576 6596 1584
rect 6508 1476 6516 1484
rect 6572 1456 6580 1464
rect 6524 1356 6532 1364
rect 6556 1336 6564 1344
rect 6348 1156 6356 1164
rect 6396 1156 6404 1164
rect 6364 1136 6372 1144
rect 6380 1136 6388 1144
rect 6332 1116 6340 1124
rect 6316 1076 6324 1084
rect 6268 1056 6276 1064
rect 6252 936 6260 944
rect 6236 916 6244 924
rect 6220 876 6228 884
rect 6252 836 6260 844
rect 6236 816 6244 824
rect 6284 1036 6292 1044
rect 6316 956 6324 964
rect 6300 936 6308 944
rect 6300 916 6308 924
rect 6316 896 6324 904
rect 6284 876 6292 884
rect 6348 1076 6356 1084
rect 6396 1116 6404 1124
rect 6428 1176 6436 1184
rect 6380 1096 6388 1104
rect 6412 1096 6420 1104
rect 6364 1036 6372 1044
rect 6364 1016 6372 1024
rect 6348 956 6356 964
rect 6348 936 6356 944
rect 6268 796 6276 804
rect 6268 776 6276 784
rect 6236 696 6244 704
rect 6300 696 6308 704
rect 6252 676 6260 684
rect 6268 676 6276 684
rect 6220 656 6228 664
rect 6204 496 6212 504
rect 6236 636 6244 644
rect 6236 556 6244 564
rect 6268 556 6276 564
rect 6236 536 6244 544
rect 6268 536 6276 544
rect 6220 476 6228 484
rect 6252 476 6260 484
rect 6236 396 6244 404
rect 6188 356 6196 364
rect 6172 316 6180 324
rect 6156 256 6164 264
rect 6172 236 6180 244
rect 6204 236 6212 244
rect 6028 156 6036 164
rect 6140 156 6148 164
rect 5740 136 5748 144
rect 5916 136 5924 144
rect 6044 136 6052 144
rect 6092 136 6100 144
rect 6172 136 6180 144
rect 6236 136 6244 144
rect 5180 116 5188 124
rect 5276 118 5284 124
rect 5276 116 5284 118
rect 5404 116 5412 124
rect 5644 116 5652 124
rect 5852 118 5860 124
rect 5852 116 5860 118
rect 5916 116 5924 124
rect 6124 116 6132 124
rect 5148 96 5156 104
rect 4940 76 4948 84
rect 5068 76 5076 84
rect 5116 76 5124 84
rect 6188 96 6196 104
rect 6156 76 6164 84
rect 3244 56 3252 64
rect 3260 56 3268 64
rect 3500 56 3508 64
rect 3612 56 3620 64
rect 3676 56 3684 64
rect 3772 56 3780 64
rect 4044 56 4052 64
rect 3372 36 3380 44
rect 3724 36 3732 44
rect 6236 36 6244 44
rect 1774 6 1782 14
rect 1788 6 1796 14
rect 1802 6 1810 14
rect 3100 16 3108 24
rect 3180 16 3188 24
rect 3260 16 3268 24
rect 3980 16 3988 24
rect 4830 6 4838 14
rect 4844 6 4852 14
rect 4858 6 4866 14
rect 5612 16 5620 24
rect 6332 736 6340 744
rect 6348 696 6356 704
rect 6348 676 6356 684
rect 6332 656 6340 664
rect 6316 536 6324 544
rect 6332 536 6340 544
rect 6316 516 6324 524
rect 6300 296 6308 304
rect 6284 276 6292 284
rect 6412 1076 6420 1084
rect 6460 1216 6468 1224
rect 6460 1176 6468 1184
rect 6444 1096 6452 1104
rect 6396 976 6404 984
rect 6380 916 6388 924
rect 6380 836 6388 844
rect 6444 1036 6452 1044
rect 6412 936 6420 944
rect 6444 996 6452 1004
rect 6508 1296 6516 1304
rect 6572 1196 6580 1204
rect 6556 1176 6564 1184
rect 6572 1156 6580 1164
rect 6508 1136 6516 1144
rect 6556 1136 6564 1144
rect 6524 1116 6532 1124
rect 6492 1096 6500 1104
rect 6508 1096 6516 1104
rect 6476 996 6484 1004
rect 6460 976 6468 984
rect 6444 936 6452 944
rect 6412 916 6420 924
rect 6396 756 6404 764
rect 6380 716 6388 724
rect 6380 696 6388 704
rect 6396 676 6404 684
rect 6364 656 6372 664
rect 6396 636 6404 644
rect 6364 596 6372 604
rect 6348 336 6356 344
rect 6380 416 6388 424
rect 6364 316 6372 324
rect 6348 236 6356 244
rect 6284 156 6292 164
rect 6300 156 6308 164
rect 6332 136 6340 144
rect 6300 116 6308 124
rect 6316 116 6324 124
rect 6348 96 6356 104
rect 6284 56 6292 64
rect 6252 16 6260 24
rect 6268 16 6276 24
rect 6364 56 6372 64
rect 6444 896 6452 904
rect 6476 956 6484 964
rect 6540 1096 6548 1104
rect 6460 856 6468 864
rect 6460 836 6468 844
rect 6492 816 6500 824
rect 6492 756 6500 764
rect 6444 696 6452 704
rect 6428 676 6436 684
rect 6444 676 6452 684
rect 6476 696 6484 704
rect 6460 636 6468 644
rect 6444 616 6452 624
rect 6428 576 6436 584
rect 6556 1076 6564 1084
rect 6524 1056 6532 1064
rect 6540 1056 6548 1064
rect 6524 1036 6532 1044
rect 6604 936 6612 944
rect 6572 916 6580 924
rect 6524 876 6532 884
rect 6556 876 6564 884
rect 6524 716 6532 724
rect 6556 736 6564 744
rect 6556 696 6564 704
rect 6540 596 6548 604
rect 6492 576 6500 584
rect 6508 576 6516 584
rect 6540 576 6548 584
rect 6508 556 6516 564
rect 6444 516 6452 524
rect 6492 496 6500 504
rect 6412 396 6420 404
rect 6412 376 6420 384
rect 6396 356 6404 364
rect 6428 356 6436 364
rect 6428 336 6436 344
rect 6412 276 6420 284
rect 6396 176 6404 184
rect 6476 296 6484 304
rect 6476 276 6484 284
rect 6444 136 6452 144
rect 6524 476 6532 484
rect 6508 316 6516 324
rect 6492 156 6500 164
rect 6396 96 6404 104
rect 6460 96 6468 104
rect 6300 16 6308 24
rect 6316 16 6324 24
rect 6348 16 6356 24
rect 6364 16 6372 24
rect 6380 16 6388 24
rect 6428 76 6436 84
rect 6604 916 6612 924
rect 6604 716 6612 724
rect 6636 1136 6644 1144
rect 6636 1116 6644 1124
rect 6636 1076 6644 1084
rect 6620 696 6628 704
rect 6588 676 6596 684
rect 6604 656 6612 664
rect 6572 556 6580 564
rect 6540 356 6548 364
rect 6604 356 6612 364
rect 6556 216 6564 224
rect 6620 276 6628 284
rect 6716 536 6724 544
rect 6636 256 6644 264
rect 6620 196 6628 204
rect 6604 176 6612 184
rect 6524 156 6532 164
rect 6620 136 6628 144
rect 6572 76 6580 84
rect 6460 36 6468 44
rect 6492 36 6500 44
rect 6492 16 6500 24
rect 6540 16 6548 24
rect 6604 56 6612 64
rect 6636 36 6644 44
<< metal3 >>
rect -19 4803 -13 4823
rect 6669 4817 6716 4823
rect 1768 4814 1816 4816
rect 1768 4806 1772 4814
rect 1782 4806 1788 4814
rect 1796 4806 1802 4814
rect 1812 4806 1816 4814
rect 1768 4804 1816 4806
rect 4824 4814 4872 4816
rect 4824 4806 4828 4814
rect 4838 4806 4844 4814
rect 4852 4806 4858 4814
rect 4868 4806 4872 4814
rect 4824 4804 4872 4806
rect -19 4797 1740 4803
rect 1844 4797 2508 4803
rect 2580 4797 2732 4803
rect 2740 4797 3244 4803
rect -19 4777 2220 4783
rect 2228 4777 2332 4783
rect 2372 4777 3212 4783
rect 6580 4777 6675 4783
rect 628 4757 3116 4763
rect 4900 4757 5068 4763
rect 5092 4757 5180 4763
rect 6580 4757 6716 4763
rect -19 4737 12 4743
rect 116 4737 252 4743
rect 260 4737 380 4743
rect 468 4737 508 4743
rect 516 4737 556 4743
rect 644 4737 812 4743
rect 836 4737 892 4743
rect 916 4737 940 4743
rect 964 4737 3084 4743
rect 3156 4737 3340 4743
rect 4996 4737 5196 4743
rect 5204 4737 5276 4743
rect 5492 4737 5516 4743
rect 5524 4737 5548 4743
rect 6180 4737 6220 4743
rect 6324 4737 6524 4743
rect 6628 4737 6675 4743
rect -19 4717 1516 4723
rect -19 4697 -13 4717
rect 1524 4717 1612 4723
rect 1636 4717 1852 4723
rect 1876 4717 1916 4723
rect 1924 4717 1980 4723
rect 2004 4717 2028 4723
rect 2100 4717 2156 4723
rect 2244 4717 2252 4723
rect 2324 4717 2428 4723
rect 2484 4717 2540 4723
rect 2564 4717 2572 4723
rect 2612 4717 2684 4723
rect 2740 4717 2988 4723
rect 3028 4717 3036 4723
rect 3060 4717 3116 4723
rect 3796 4717 3820 4723
rect 4052 4717 4284 4723
rect 4292 4717 4332 4723
rect 4532 4717 4572 4723
rect 4884 4717 5084 4723
rect 5124 4717 5164 4723
rect 5268 4717 5340 4723
rect 5380 4717 5420 4723
rect 5508 4717 5660 4723
rect 5668 4717 5708 4723
rect 6116 4717 6204 4723
rect 6500 4717 6540 4723
rect 20 4697 851 4703
rect -19 4677 428 4683
rect -19 4657 -13 4677
rect 436 4677 460 4683
rect 500 4677 540 4683
rect 548 4677 620 4683
rect 740 4677 828 4683
rect 845 4683 851 4697
rect 868 4697 972 4703
rect 1012 4697 1036 4703
rect 1076 4697 1164 4703
rect 1188 4697 1196 4703
rect 1220 4697 1324 4703
rect 1396 4697 3020 4703
rect 3124 4697 3212 4703
rect 3652 4697 3772 4703
rect 3828 4697 3916 4703
rect 4340 4697 5276 4703
rect 5284 4697 5324 4703
rect 5684 4697 5964 4703
rect 5972 4697 6060 4703
rect 6068 4697 6252 4703
rect 6484 4697 6508 4703
rect 6669 4697 6716 4703
rect 845 4677 892 4683
rect 916 4677 956 4683
rect 973 4683 979 4696
rect 973 4677 1100 4683
rect 1124 4677 1363 4683
rect 84 4657 124 4663
rect 132 4657 252 4663
rect 356 4657 396 4663
rect 532 4657 636 4663
rect 676 4657 732 4663
rect 772 4657 908 4663
rect 948 4657 1068 4663
rect 1172 4657 1228 4663
rect 1284 4657 1340 4663
rect 1357 4663 1363 4677
rect 1380 4677 1420 4683
rect 1460 4677 1532 4683
rect 1549 4677 1836 4683
rect 1549 4663 1555 4677
rect 1844 4677 1932 4683
rect 1956 4677 1980 4683
rect 2004 4677 2732 4683
rect 2868 4677 2972 4683
rect 2996 4677 3180 4683
rect 3252 4677 3516 4683
rect 3556 4677 3660 4683
rect 3668 4677 3692 4683
rect 3988 4677 4076 4683
rect 4324 4677 4364 4683
rect 4692 4677 4876 4683
rect 4932 4677 5036 4683
rect 5044 4677 5100 4683
rect 5108 4677 5196 4683
rect 5268 4677 5292 4683
rect 5316 4677 5388 4683
rect 5396 4677 5484 4683
rect 5492 4677 5564 4683
rect 5620 4677 5676 4683
rect 5684 4677 5740 4683
rect 5780 4677 5836 4683
rect 5844 4677 5868 4683
rect 5892 4677 5916 4683
rect 5956 4677 6076 4683
rect 6164 4677 6316 4683
rect 1357 4657 1555 4663
rect 1604 4657 1692 4663
rect 1748 4657 1772 4663
rect 1780 4657 1884 4663
rect 2180 4657 2220 4663
rect 2292 4657 2316 4663
rect 2324 4657 2364 4663
rect 2516 4657 2588 4663
rect 2644 4657 2652 4663
rect 2932 4657 3036 4663
rect 4308 4657 4396 4663
rect 4500 4657 4716 4663
rect 4788 4657 4828 4663
rect 4877 4663 4883 4676
rect 4877 4657 4940 4663
rect 4996 4657 5020 4663
rect 5076 4657 5100 4663
rect 5124 4657 5244 4663
rect 5444 4657 5500 4663
rect 5716 4657 5820 4663
rect 5828 4657 5980 4663
rect 6020 4657 6028 4663
rect 6077 4663 6083 4676
rect 6077 4657 6284 4663
rect 6612 4657 6675 4663
rect -19 4637 355 4643
rect -19 4617 -13 4637
rect 180 4617 332 4623
rect 349 4623 355 4637
rect 628 4637 684 4643
rect 708 4637 924 4643
rect 964 4637 1004 4643
rect 1012 4637 1116 4643
rect 1188 4637 1260 4643
rect 1300 4637 1308 4643
rect 1332 4637 1388 4643
rect 1412 4637 1420 4643
rect 1444 4637 1484 4643
rect 1508 4637 1580 4643
rect 1604 4637 2060 4643
rect 2164 4637 2252 4643
rect 2797 4637 3068 4643
rect 701 4623 707 4636
rect 349 4617 707 4623
rect 2797 4623 2803 4637
rect 3412 4637 3612 4643
rect 3620 4637 3676 4643
rect 3684 4637 3708 4643
rect 3860 4637 4044 4643
rect 4084 4637 4236 4643
rect 4452 4637 4604 4643
rect 4900 4637 4956 4643
rect 4964 4637 5164 4643
rect 5348 4637 5548 4643
rect 5716 4637 5804 4643
rect 5876 4637 5996 4643
rect 6020 4637 6044 4643
rect 6052 4637 6108 4643
rect 1412 4617 2803 4623
rect 2820 4617 2860 4623
rect 2868 4617 2988 4623
rect 3444 4617 3484 4623
rect 4260 4617 4588 4623
rect 4596 4617 4723 4623
rect 3304 4614 3352 4616
rect 3304 4606 3308 4614
rect 3318 4606 3324 4614
rect 3332 4606 3338 4614
rect 3348 4606 3352 4614
rect 3304 4604 3352 4606
rect -19 4597 1091 4603
rect -19 4577 -13 4597
rect 1085 4584 1091 4597
rect 1108 4597 1548 4603
rect 1572 4597 1724 4603
rect 1732 4597 3148 4603
rect 3492 4597 3628 4603
rect 4500 4597 4684 4603
rect 4717 4603 4723 4617
rect 4740 4617 4812 4623
rect 4820 4617 4988 4623
rect 5428 4617 5644 4623
rect 5805 4623 5811 4636
rect 5805 4617 6028 4623
rect 6036 4617 6124 4623
rect 6132 4617 6172 4623
rect 6452 4617 6476 4623
rect 4717 4597 5340 4603
rect 5364 4597 5596 4603
rect 5604 4597 5628 4603
rect 6669 4603 6675 4623
rect 5876 4597 6675 4603
rect 20 4577 188 4583
rect 196 4577 316 4583
rect 644 4577 1020 4583
rect 1092 4577 1244 4583
rect 1380 4577 1404 4583
rect 1476 4577 1500 4583
rect 1508 4577 1548 4583
rect 1556 4577 1676 4583
rect 1844 4577 2060 4583
rect 2116 4577 2156 4583
rect 2189 4577 2252 4583
rect 164 4557 220 4563
rect 388 4557 444 4563
rect 628 4557 940 4563
rect 1060 4557 1452 4563
rect 1476 4557 1516 4563
rect 1556 4557 1820 4563
rect 1828 4557 1852 4563
rect 1892 4557 2051 4563
rect 2045 4544 2051 4557
rect 2116 4557 2140 4563
rect 2189 4563 2195 4577
rect 2420 4577 2556 4583
rect 2644 4577 2956 4583
rect 4452 4577 4508 4583
rect 4580 4577 4956 4583
rect 5060 4577 5516 4583
rect 5572 4577 5948 4583
rect 6068 4577 6604 4583
rect 6644 4577 6675 4583
rect 2148 4557 2195 4563
rect 2212 4557 2300 4563
rect 2372 4557 2444 4563
rect 2452 4557 2492 4563
rect 2660 4557 2668 4563
rect 2676 4557 2684 4563
rect 2772 4557 2796 4563
rect 2820 4557 2892 4563
rect 3188 4557 3276 4563
rect 3284 4557 3404 4563
rect 3524 4557 3756 4563
rect 3764 4557 3916 4563
rect 4516 4557 4652 4563
rect 4724 4557 4812 4563
rect 5252 4557 5388 4563
rect 5588 4557 5612 4563
rect 5940 4557 6028 4563
rect 6036 4557 6092 4563
rect 6132 4557 6188 4563
rect -19 4537 12 4543
rect 52 4537 92 4543
rect 276 4537 316 4543
rect 436 4537 476 4543
rect 500 4537 636 4543
rect 660 4537 796 4543
rect 804 4537 1036 4543
rect 1044 4537 1148 4543
rect 1220 4537 1340 4543
rect 1460 4537 1532 4543
rect 1540 4537 1660 4543
rect 1684 4537 1724 4543
rect 1908 4537 1948 4543
rect 2052 4537 2108 4543
rect 2196 4537 2220 4543
rect 2244 4537 2284 4543
rect 2292 4537 2380 4543
rect 2500 4537 2524 4543
rect 2628 4537 2668 4543
rect 2804 4537 2844 4543
rect 2852 4537 2908 4543
rect 3108 4537 3244 4543
rect 3300 4537 3372 4543
rect 3396 4537 3516 4543
rect 3668 4537 3852 4543
rect 3860 4537 4300 4543
rect 4308 4537 4364 4543
rect 4388 4537 4572 4543
rect 4596 4537 4780 4543
rect 5044 4537 5708 4543
rect 5716 4537 5740 4543
rect 5748 4537 5868 4543
rect 5892 4537 5964 4543
rect 6036 4537 6044 4543
rect 6052 4537 6108 4543
rect 6148 4537 6300 4543
rect 6308 4537 6380 4543
rect 6564 4537 6604 4543
rect 6644 4537 6675 4543
rect 84 4517 204 4523
rect 276 4517 332 4523
rect 404 4517 595 4523
rect -19 4483 -13 4503
rect 68 4497 172 4503
rect 308 4497 348 4503
rect 372 4497 524 4503
rect 532 4497 572 4503
rect 589 4503 595 4517
rect 772 4517 972 4523
rect 1140 4517 1276 4523
rect 1284 4517 1372 4523
rect 1508 4517 1564 4523
rect 1572 4517 1628 4523
rect 1636 4517 1708 4523
rect 1716 4517 1756 4523
rect 1972 4517 2092 4523
rect 2100 4517 2140 4523
rect 2436 4517 2476 4523
rect 2532 4517 2620 4523
rect 2628 4517 2700 4523
rect 2868 4517 2940 4523
rect 2964 4517 3036 4523
rect 3220 4517 3260 4523
rect 3268 4517 3276 4523
rect 3389 4523 3395 4536
rect 3284 4517 3395 4523
rect 3444 4517 3468 4523
rect 3524 4517 3548 4523
rect 3636 4517 3724 4523
rect 3796 4517 3916 4523
rect 4116 4517 4252 4523
rect 4260 4517 4316 4523
rect 4532 4517 4604 4523
rect 4772 4517 4860 4523
rect 4996 4517 5100 4523
rect 5108 4517 5148 4523
rect 5284 4517 5436 4523
rect 5844 4517 6188 4523
rect 6212 4517 6428 4523
rect 6436 4517 6492 4523
rect 589 4497 1100 4503
rect 1236 4497 1292 4503
rect 1428 4497 1484 4503
rect 1572 4497 1596 4503
rect 1684 4497 2188 4503
rect 2196 4497 2268 4503
rect 2564 4497 2652 4503
rect 2948 4497 3020 4503
rect 3172 4497 3228 4503
rect 3268 4497 3340 4503
rect 3428 4497 3500 4503
rect 4356 4497 4540 4503
rect 4548 4497 4652 4503
rect 4676 4497 4844 4503
rect 4852 4497 4940 4503
rect 5012 4497 5052 4503
rect 5060 4497 5116 4503
rect 5124 4497 5180 4503
rect 5380 4497 5404 4503
rect 5412 4497 5468 4503
rect 5764 4497 5900 4503
rect 5908 4497 6012 4503
rect 6260 4497 6316 4503
rect 6324 4497 6364 4503
rect -19 4477 12 4483
rect 36 4477 268 4483
rect 276 4477 380 4483
rect 404 4477 556 4483
rect 1108 4477 1340 4483
rect 1700 4477 1756 4483
rect 2228 4477 2332 4483
rect 2340 4477 2348 4483
rect 3380 4477 3580 4483
rect 4148 4477 4268 4483
rect 4276 4477 4380 4483
rect 4564 4477 4588 4483
rect 4660 4477 5084 4483
rect 5092 4477 5132 4483
rect 5236 4477 5580 4483
rect 5700 4477 5772 4483
rect 5780 4477 5852 4483
rect 6084 4477 6268 4483
rect -19 4443 -13 4463
rect 228 4457 268 4463
rect 308 4457 1020 4463
rect 1284 4457 1308 4463
rect 1332 4457 2492 4463
rect 3380 4457 3484 4463
rect 4484 4457 4540 4463
rect 4628 4457 4748 4463
rect 4964 4457 5020 4463
rect 5156 4457 5292 4463
rect 5540 4457 5660 4463
rect 5668 4457 5772 4463
rect 5796 4457 6076 4463
rect 6180 4457 6444 4463
rect 6452 4457 6492 4463
rect -19 4437 2764 4443
rect 2900 4437 2940 4443
rect 3876 4437 4044 4443
rect 4052 4437 4620 4443
rect 4628 4437 5308 4443
rect 5316 4437 5420 4443
rect 5428 4437 5468 4443
rect 5476 4437 5516 4443
rect 5844 4437 6140 4443
rect 6420 4437 6508 4443
rect -19 4417 419 4423
rect -19 4397 396 4403
rect -19 4377 -13 4397
rect 413 4403 419 4417
rect 580 4417 1324 4423
rect 2580 4417 2636 4423
rect 2644 4417 3052 4423
rect 3060 4417 3564 4423
rect 3572 4417 3628 4423
rect 3636 4417 3660 4423
rect 3668 4417 3788 4423
rect 4484 4417 4508 4423
rect 4548 4417 4684 4423
rect 4692 4417 4796 4423
rect 5108 4417 5164 4423
rect 5172 4417 5244 4423
rect 5380 4417 5724 4423
rect 5732 4417 5932 4423
rect 6100 4417 6396 4423
rect 6436 4417 6556 4423
rect 1768 4414 1816 4416
rect 1768 4406 1772 4414
rect 1782 4406 1788 4414
rect 1796 4406 1802 4414
rect 1812 4406 1816 4414
rect 1768 4404 1816 4406
rect 4824 4414 4872 4416
rect 4824 4406 4828 4414
rect 4838 4406 4844 4414
rect 4852 4406 4858 4414
rect 4868 4406 4872 4414
rect 4824 4404 4872 4406
rect 413 4397 1324 4403
rect 5028 4397 5580 4403
rect 6404 4397 6460 4403
rect 20 4377 1036 4383
rect 1165 4377 1724 4383
rect 20 4357 44 4363
rect 676 4357 764 4363
rect 1165 4363 1171 4377
rect 1732 4377 1740 4383
rect 1748 4377 1852 4383
rect 3060 4377 3420 4383
rect 4084 4377 4108 4383
rect 4836 4377 4988 4383
rect 5300 4377 5388 4383
rect 5684 4377 6092 4383
rect 6292 4377 6476 4383
rect 820 4357 1171 4363
rect 1220 4357 1244 4363
rect 2052 4357 2268 4363
rect 2340 4357 2508 4363
rect 2804 4357 2876 4363
rect 3028 4357 3532 4363
rect 4404 4357 4700 4363
rect 5172 4357 5260 4363
rect 6244 4357 6396 4363
rect 6404 4357 6492 4363
rect -19 4337 236 4343
rect 580 4337 780 4343
rect 1172 4337 1244 4343
rect 1988 4337 2188 4343
rect 2260 4337 2460 4343
rect 2884 4337 2924 4343
rect 3076 4337 3292 4343
rect 3396 4337 3628 4343
rect 4164 4337 4204 4343
rect 4468 4337 4524 4343
rect 4628 4337 4780 4343
rect 5236 4337 5324 4343
rect 5396 4337 5436 4343
rect 5444 4337 5452 4343
rect 5620 4337 6076 4343
rect 6084 4337 6188 4343
rect 6196 4337 6284 4343
rect 6324 4337 6460 4343
rect 6468 4337 6540 4343
rect 132 4317 252 4323
rect 260 4317 268 4323
rect 388 4317 428 4323
rect 756 4317 924 4323
rect 1092 4317 1308 4323
rect 1604 4317 1660 4323
rect 1716 4317 1772 4323
rect 2036 4317 2076 4323
rect 2084 4317 2156 4323
rect 2404 4317 2540 4323
rect 2596 4317 2828 4323
rect 2868 4317 2988 4323
rect 2996 4317 3212 4323
rect 3220 4317 3420 4323
rect 3844 4317 3884 4323
rect 3940 4317 3948 4323
rect 4068 4317 4140 4323
rect 4372 4317 4396 4323
rect 4500 4317 4556 4323
rect 4564 4317 4604 4323
rect 4644 4317 4668 4323
rect 4884 4317 5084 4323
rect 5092 4317 5340 4323
rect 5428 4317 5580 4323
rect 5940 4317 5964 4323
rect 5972 4317 6060 4323
rect 6292 4317 6380 4323
rect 6436 4317 6524 4323
rect 6548 4317 6588 4323
rect -19 4297 28 4303
rect 52 4297 76 4303
rect 180 4297 316 4303
rect 324 4297 396 4303
rect 516 4297 556 4303
rect 564 4297 652 4303
rect 660 4297 700 4303
rect 868 4297 908 4303
rect 916 4297 1004 4303
rect 1076 4297 1132 4303
rect 1140 4297 1228 4303
rect 1252 4297 1276 4303
rect 1396 4297 1452 4303
rect 1588 4297 2220 4303
rect 2500 4297 2524 4303
rect 2532 4297 2588 4303
rect 2612 4297 2652 4303
rect 2708 4297 2956 4303
rect 2964 4297 3107 4303
rect 3101 4284 3107 4297
rect 3140 4297 3164 4303
rect 3444 4297 3532 4303
rect 3940 4297 3996 4303
rect 4068 4297 4236 4303
rect 4244 4297 4268 4303
rect 4372 4297 4444 4303
rect 4452 4297 4508 4303
rect 4516 4297 4540 4303
rect 4580 4297 4668 4303
rect 4676 4297 4716 4303
rect 4804 4297 4892 4303
rect 5124 4297 5324 4303
rect 5332 4297 5404 4303
rect 5412 4297 5484 4303
rect 5508 4297 5516 4303
rect 5524 4297 5548 4303
rect 5764 4297 6012 4303
rect 6036 4297 6316 4303
rect 6356 4297 6444 4303
rect 6484 4297 6604 4303
rect 68 4277 92 4283
rect 100 4277 588 4283
rect 596 4277 812 4283
rect 820 4277 1116 4283
rect 1124 4277 1372 4283
rect 1380 4277 1548 4283
rect 1700 4277 1916 4283
rect 1924 4277 2092 4283
rect 2116 4277 2204 4283
rect 2596 4277 2684 4283
rect 2948 4277 2988 4283
rect 3108 4277 3164 4283
rect 3268 4277 3372 4283
rect 3460 4277 3500 4283
rect 3956 4277 4092 4283
rect 4196 4277 4316 4283
rect 4660 4277 4716 4283
rect 5188 4277 5260 4283
rect 5268 4277 5388 4283
rect 5476 4277 5548 4283
rect 5604 4277 5644 4283
rect 5684 4277 5868 4283
rect 6308 4277 6348 4283
rect 6468 4277 6524 4283
rect 6548 4277 6636 4283
rect -19 4257 12 4263
rect 36 4257 108 4263
rect 116 4257 140 4263
rect 212 4257 300 4263
rect 340 4257 572 4263
rect 612 4257 748 4263
rect 788 4257 828 4263
rect 836 4257 876 4263
rect 916 4257 940 4263
rect 996 4257 1020 4263
rect 1044 4257 1068 4263
rect 1844 4257 1996 4263
rect 2196 4257 2220 4263
rect 3204 4257 3244 4263
rect 3572 4257 3596 4263
rect 3604 4257 3740 4263
rect 4084 4257 4124 4263
rect 4660 4257 4700 4263
rect 4868 4257 4972 4263
rect 4980 4257 5036 4263
rect 5140 4257 5196 4263
rect 5236 4257 5404 4263
rect 5549 4263 5555 4276
rect 5549 4257 5628 4263
rect 5684 4257 5740 4263
rect 5748 4257 5900 4263
rect 5908 4257 5916 4263
rect 5924 4257 5980 4263
rect 6052 4257 6108 4263
rect 6116 4257 6204 4263
rect 6292 4257 6412 4263
rect 6532 4257 6556 4263
rect 6580 4257 6636 4263
rect 244 4237 268 4243
rect 292 4237 348 4243
rect 436 4237 492 4243
rect 660 4237 684 4243
rect 692 4237 716 4243
rect 1140 4237 1964 4243
rect 1972 4237 2028 4243
rect 2436 4237 2636 4243
rect 2644 4237 2732 4243
rect 3252 4237 3516 4243
rect 3524 4237 4140 4243
rect 4948 4237 5532 4243
rect 5748 4237 5804 4243
rect 5940 4237 6620 4243
rect -19 4217 188 4223
rect 436 4217 460 4223
rect 468 4217 652 4223
rect 1076 4217 1420 4223
rect 1876 4217 2236 4223
rect 2244 4217 2300 4223
rect 2756 4217 2796 4223
rect 2804 4217 2844 4223
rect 2852 4217 2892 4223
rect 3252 4217 3276 4223
rect 3396 4217 3484 4223
rect 3492 4217 3564 4223
rect 4132 4217 5116 4223
rect 5140 4217 5692 4223
rect 6260 4217 6316 4223
rect 3304 4214 3352 4216
rect 3304 4206 3308 4214
rect 3318 4206 3324 4214
rect 3332 4206 3338 4214
rect 3348 4206 3352 4214
rect 3304 4204 3352 4206
rect 340 4197 444 4203
rect 452 4197 860 4203
rect 916 4197 956 4203
rect 1332 4197 1356 4203
rect 2132 4197 2252 4203
rect 3572 4197 4204 4203
rect 4420 4197 4796 4203
rect 4804 4197 4940 4203
rect 6004 4197 6588 4203
rect -19 4177 76 4183
rect 324 4177 620 4183
rect 628 4177 668 4183
rect 740 4177 764 4183
rect 1124 4177 1148 4183
rect 2228 4177 2620 4183
rect 2836 4177 2860 4183
rect 2996 4177 3132 4183
rect 3140 4177 3228 4183
rect 3284 4177 3548 4183
rect 3812 4177 3868 4183
rect 4740 4177 4748 4183
rect 4756 4177 5148 4183
rect 6068 4177 6092 4183
rect 6100 4177 6204 4183
rect 6340 4177 6380 4183
rect 6468 4177 6556 4183
rect 404 4157 556 4163
rect 660 4157 876 4163
rect 1108 4157 1276 4163
rect 1620 4157 1660 4163
rect 1668 4157 1884 4163
rect 2020 4157 2156 4163
rect 2340 4157 2428 4163
rect 2452 4157 2476 4163
rect 2660 4157 2748 4163
rect 2868 4157 2876 4163
rect 2916 4157 2940 4163
rect 3156 4157 3564 4163
rect 3588 4157 3644 4163
rect 3652 4157 3724 4163
rect 3732 4157 3756 4163
rect 3764 4157 3852 4163
rect 3860 4157 3916 4163
rect 4084 4157 4428 4163
rect 4436 4157 4556 4163
rect 4580 4157 4620 4163
rect 4932 4157 5068 4163
rect 5124 4157 5260 4163
rect 5476 4157 5500 4163
rect 5780 4157 5868 4163
rect 5940 4157 6067 4163
rect 212 4137 348 4143
rect 420 4137 540 4143
rect 548 4137 604 4143
rect 1012 4137 1164 4143
rect 1348 4137 1484 4143
rect 1764 4137 1868 4143
rect 1876 4137 1900 4143
rect 1908 4137 2028 4143
rect 2036 4137 2060 4143
rect 2084 4137 2124 4143
rect 2308 4137 2364 4143
rect 2420 4137 2588 4143
rect 2596 4137 2636 4143
rect 2708 4137 2764 4143
rect 2772 4137 2908 4143
rect 2996 4137 3260 4143
rect 3476 4137 3980 4143
rect 4308 4137 4492 4143
rect 4500 4137 4540 4143
rect 4564 4137 4604 4143
rect 4756 4137 4844 4143
rect 5060 4137 5100 4143
rect 5236 4137 5420 4143
rect 5652 4137 5708 4143
rect 5988 4137 6012 4143
rect 6061 4143 6067 4157
rect 6084 4157 6124 4163
rect 6388 4157 6396 4163
rect 6484 4157 6524 4163
rect 6061 4137 6092 4143
rect 6116 4137 6156 4143
rect 6196 4137 6220 4143
rect 6356 4137 6444 4143
rect 6452 4137 6556 4143
rect 52 4117 108 4123
rect 580 4117 1596 4123
rect 1604 4117 1676 4123
rect 1684 4117 2140 4123
rect 2148 4117 2236 4123
rect 2276 4117 2675 4123
rect 20 4097 780 4103
rect 868 4097 1116 4103
rect 1188 4097 1260 4103
rect 1924 4097 2060 4103
rect 2084 4097 2220 4103
rect 2356 4097 2364 4103
rect 2372 4097 2508 4103
rect 2669 4103 2675 4117
rect 2692 4117 2716 4123
rect 2884 4117 2924 4123
rect 2964 4117 3148 4123
rect 3364 4117 3420 4123
rect 3540 4117 3692 4123
rect 3700 4117 3756 4123
rect 3764 4117 3836 4123
rect 3844 4117 3932 4123
rect 4276 4117 4364 4123
rect 4468 4117 4476 4123
rect 4484 4117 4620 4123
rect 4628 4117 4636 4123
rect 4644 4117 4652 4123
rect 4957 4117 4972 4123
rect 2669 4097 2780 4103
rect 2788 4097 2828 4103
rect 3076 4097 3212 4103
rect 3220 4097 3308 4103
rect 3572 4097 3676 4103
rect 3748 4097 3788 4103
rect 3796 4097 3964 4103
rect 4532 4097 4620 4103
rect 4628 4097 4684 4103
rect 4957 4103 4963 4117
rect 5332 4117 5372 4123
rect 5524 4117 5580 4123
rect 5812 4117 5916 4123
rect 5924 4117 5932 4123
rect 5972 4117 6012 4123
rect 6052 4117 6252 4123
rect 6260 4117 6476 4123
rect 4724 4097 4963 4103
rect 4980 4097 5196 4103
rect 5204 4097 5308 4103
rect 5316 4097 5340 4103
rect 5652 4097 5996 4103
rect 6004 4097 6060 4103
rect 6100 4097 6124 4103
rect 6132 4097 6188 4103
rect 6244 4097 6300 4103
rect 6308 4097 6364 4103
rect 6404 4097 6508 4103
rect 6516 4097 6588 4103
rect 244 4077 1132 4083
rect 2356 4077 2380 4083
rect 2388 4077 2412 4083
rect 2644 4077 2716 4083
rect 3380 4077 3596 4083
rect 3677 4083 3683 4096
rect 3677 4077 3804 4083
rect 3892 4077 4044 4083
rect 4052 4077 4092 4083
rect 4100 4077 4156 4083
rect 4164 4077 4268 4083
rect 4660 4077 4764 4083
rect 4772 4077 4812 4083
rect 4932 4077 4956 4083
rect 5412 4077 5676 4083
rect 5684 4077 5852 4083
rect 5908 4077 6028 4083
rect 6228 4077 6332 4083
rect 6340 4077 6412 4083
rect 1316 4057 1628 4063
rect 2068 4057 2332 4063
rect 2452 4057 2652 4063
rect 3668 4057 3900 4063
rect 5012 4057 5708 4063
rect 5716 4057 5756 4063
rect 5844 4057 5868 4063
rect 5988 4057 6284 4063
rect 6340 4057 6380 4063
rect 6404 4057 6572 4063
rect 1620 4037 1820 4043
rect 1828 4037 2108 4043
rect 2516 4037 3388 4043
rect 3428 4037 3772 4043
rect 4772 4037 5164 4043
rect 5172 4037 5276 4043
rect 5348 4037 5468 4043
rect 6228 4037 6540 4043
rect 2100 4017 3004 4023
rect 3124 4017 3436 4023
rect 4932 4017 5068 4023
rect 5540 4017 5788 4023
rect 6164 4017 6348 4023
rect 6420 4017 6444 4023
rect 1768 4014 1816 4016
rect 1768 4006 1772 4014
rect 1782 4006 1788 4014
rect 1796 4006 1802 4014
rect 1812 4006 1816 4014
rect 1768 4004 1816 4006
rect 4824 4014 4872 4016
rect 4824 4006 4828 4014
rect 4838 4006 4844 4014
rect 4852 4006 4858 4014
rect 4868 4006 4872 4014
rect 4824 4004 4872 4006
rect 2676 3997 2860 4003
rect 2868 3997 3036 4003
rect 5044 3997 5052 4003
rect 5252 3997 5628 4003
rect 5780 3997 6332 4003
rect 6340 3997 6556 4003
rect 580 3977 636 3983
rect 644 3977 780 3983
rect 1188 3977 1324 3983
rect 5588 3977 5708 3983
rect 6052 3977 6444 3983
rect 1140 3957 1276 3963
rect 3716 3957 4188 3963
rect 4644 3957 4716 3963
rect 5076 3957 5308 3963
rect 5572 3957 6028 3963
rect 6036 3957 6108 3963
rect 36 3937 156 3943
rect 244 3937 524 3943
rect 532 3937 588 3943
rect 868 3937 1196 3943
rect 1476 3937 1612 3943
rect 1924 3937 2028 3943
rect 3924 3937 4108 3943
rect 4612 3937 5228 3943
rect 5444 3937 5580 3943
rect 5620 3937 5740 3943
rect 5828 3937 5852 3943
rect 5860 3937 5980 3943
rect 6004 3937 6236 3943
rect 6244 3937 6252 3943
rect 6276 3937 6316 3943
rect 6452 3937 6476 3943
rect 6484 3937 6540 3943
rect 6596 3937 6604 3943
rect 148 3917 204 3923
rect 228 3917 268 3923
rect 516 3917 540 3923
rect 772 3917 844 3923
rect 884 3917 956 3923
rect 1060 3917 1100 3923
rect 1108 3917 1148 3923
rect 1268 3917 1548 3923
rect 1604 3917 1628 3923
rect 2324 3917 2396 3923
rect 3796 3917 3980 3923
rect 4308 3917 4444 3923
rect 4772 3917 4908 3923
rect 4916 3917 4956 3923
rect 5060 3917 5148 3923
rect 5156 3917 5196 3923
rect 5220 3917 5283 3923
rect 100 3897 252 3903
rect 308 3897 860 3903
rect 884 3897 940 3903
rect 1108 3897 1132 3903
rect 1348 3897 1532 3903
rect 1668 3897 1692 3903
rect 1812 3897 1964 3903
rect 2116 3897 2380 3903
rect 2628 3897 2812 3903
rect 2820 3897 2828 3903
rect 2836 3897 2940 3903
rect 3044 3897 3148 3903
rect 3348 3897 3404 3903
rect 3636 3897 3676 3903
rect 4500 3897 4652 3903
rect 4708 3897 4748 3903
rect 4756 3897 4796 3903
rect 5092 3897 5132 3903
rect 5172 3897 5196 3903
rect 5220 3897 5260 3903
rect 5277 3903 5283 3917
rect 5300 3917 5340 3923
rect 5348 3917 5452 3923
rect 5540 3917 5596 3923
rect 5700 3917 5932 3923
rect 5940 3917 5948 3923
rect 6004 3917 6060 3923
rect 6164 3917 6428 3923
rect 6436 3917 6492 3923
rect 5277 3897 5516 3903
rect 5604 3897 5660 3903
rect 5828 3897 5964 3903
rect 5988 3897 5996 3903
rect 6084 3897 6092 3903
rect 6164 3897 6252 3903
rect 6324 3897 6476 3903
rect 6484 3897 6524 3903
rect 6580 3897 6604 3903
rect 180 3877 188 3883
rect 212 3877 364 3883
rect 628 3877 1084 3883
rect 1540 3877 1564 3883
rect 1684 3877 1836 3883
rect 2356 3877 2620 3883
rect 2916 3877 2988 3883
rect 3156 3877 3260 3883
rect 3268 3877 3548 3883
rect 3556 3877 3612 3883
rect 3620 3877 3644 3883
rect 3812 3877 3900 3883
rect 4116 3877 4124 3883
rect 4260 3877 4428 3883
rect 4436 3877 4460 3883
rect 4708 3877 4732 3883
rect 4900 3877 4988 3883
rect 4996 3877 5100 3883
rect 5268 3877 5420 3883
rect 5460 3877 5644 3883
rect 5716 3877 5772 3883
rect 5892 3877 6012 3883
rect 6020 3877 6076 3883
rect 6324 3877 6444 3883
rect 6516 3877 6540 3883
rect 6564 3877 6604 3883
rect 132 3857 332 3863
rect 1412 3857 1580 3863
rect 1636 3857 1676 3863
rect 2644 3857 3052 3863
rect 3540 3857 3564 3863
rect 3636 3857 3772 3863
rect 4292 3857 4396 3863
rect 4404 3857 4700 3863
rect 4708 3857 4748 3863
rect 4756 3857 4812 3863
rect 5076 3857 5180 3863
rect 5252 3857 5372 3863
rect 5380 3857 5484 3863
rect 5492 3857 5532 3863
rect 5748 3857 5820 3863
rect 5892 3857 6140 3863
rect 6148 3857 6268 3863
rect 6340 3857 6387 3863
rect 420 3837 700 3843
rect 708 3837 892 3843
rect 900 3837 908 3843
rect 1012 3837 1068 3843
rect 1572 3837 1660 3843
rect 2004 3837 2060 3843
rect 2228 3837 2460 3843
rect 2468 3837 2556 3843
rect 2964 3837 2972 3843
rect 2980 3837 3052 3843
rect 3444 3837 3788 3843
rect 4180 3837 4284 3843
rect 4372 3837 4572 3843
rect 4580 3837 4668 3843
rect 4788 3837 4940 3843
rect 5428 3837 5468 3843
rect 6068 3837 6108 3843
rect 6244 3837 6364 3843
rect 6381 3843 6387 3857
rect 6420 3857 6476 3863
rect 6381 3837 6572 3843
rect 340 3817 476 3823
rect 532 3817 716 3823
rect 1220 3817 2044 3823
rect 2180 3817 2396 3823
rect 2500 3817 2604 3823
rect 3572 3817 3740 3823
rect 4292 3817 4348 3823
rect 4356 3817 4604 3823
rect 4612 3817 4716 3823
rect 5108 3817 5132 3823
rect 5220 3817 6188 3823
rect 6356 3817 6540 3823
rect 6557 3817 6675 3823
rect 3304 3814 3352 3816
rect 3304 3806 3308 3814
rect 3318 3806 3324 3814
rect 3332 3806 3338 3814
rect 3348 3806 3352 3814
rect 3304 3804 3352 3806
rect 484 3797 620 3803
rect 628 3797 1004 3803
rect 1252 3797 1324 3803
rect 1332 3797 1932 3803
rect 2772 3797 3100 3803
rect 3556 3797 3644 3803
rect 4084 3797 4108 3803
rect 4116 3797 4268 3803
rect 4340 3797 4444 3803
rect 4532 3797 4908 3803
rect 5396 3797 5548 3803
rect 5588 3797 5644 3803
rect 5652 3797 6092 3803
rect 6276 3797 6316 3803
rect 6356 3797 6380 3803
rect 6436 3797 6444 3803
rect 6557 3803 6563 3817
rect 6516 3797 6563 3803
rect 6580 3797 6620 3803
rect 20 3777 44 3783
rect 564 3777 1148 3783
rect 1428 3777 1484 3783
rect 1668 3777 1692 3783
rect 1700 3777 1740 3783
rect 2212 3777 2284 3783
rect 2292 3777 2460 3783
rect 2884 3777 2892 3783
rect 3492 3777 3628 3783
rect 3668 3777 3916 3783
rect 3924 3777 4124 3783
rect 4132 3777 4236 3783
rect 4516 3777 4604 3783
rect 4612 3777 4684 3783
rect 4756 3777 4924 3783
rect 4932 3777 5020 3783
rect 5044 3777 5132 3783
rect 5364 3777 6620 3783
rect 6669 3777 6675 3817
rect 660 3757 764 3763
rect 836 3757 956 3763
rect 1092 3757 1164 3763
rect 1172 3757 1356 3763
rect 2484 3757 2572 3763
rect 2580 3757 2652 3763
rect 2660 3757 2988 3763
rect 3044 3757 3356 3763
rect 3364 3757 3404 3763
rect 3524 3757 3612 3763
rect 3684 3757 3804 3763
rect 4148 3757 4220 3763
rect 4228 3757 4364 3763
rect 4404 3757 4540 3763
rect 4548 3757 4668 3763
rect 4692 3757 4764 3763
rect 4772 3757 4860 3763
rect 4916 3757 4972 3763
rect 5517 3757 5692 3763
rect 5517 3744 5523 3757
rect 6452 3757 6508 3763
rect 6589 3757 6604 3763
rect 276 3737 428 3743
rect 724 3737 732 3743
rect 1060 3737 1260 3743
rect 2036 3737 2124 3743
rect 2132 3737 2172 3743
rect 2324 3737 2508 3743
rect 2884 3737 2924 3743
rect 2948 3737 3020 3743
rect 3028 3737 3244 3743
rect 3252 3737 3468 3743
rect 3476 3737 3564 3743
rect 3636 3737 3660 3743
rect 3796 3737 3948 3743
rect 4116 3737 4284 3743
rect 4324 3737 4412 3743
rect 4420 3737 4556 3743
rect 4932 3737 5036 3743
rect 5044 3737 5100 3743
rect 5140 3737 5388 3743
rect 5684 3737 5804 3743
rect 6004 3737 6044 3743
rect 6100 3737 6124 3743
rect 6180 3737 6284 3743
rect 6340 3737 6364 3743
rect 6388 3737 6428 3743
rect 212 3717 275 3723
rect 269 3704 275 3717
rect 724 3717 876 3723
rect 964 3717 1324 3723
rect 1364 3717 1500 3723
rect 1972 3717 2300 3723
rect 2340 3717 2428 3723
rect 2740 3717 2892 3723
rect 3060 3717 3132 3723
rect 3284 3717 3340 3723
rect 3460 3717 3500 3723
rect 3508 3717 3580 3723
rect 3604 3717 3676 3723
rect 4276 3717 4348 3723
rect 4596 3717 4620 3723
rect 4628 3717 4700 3723
rect 4948 3717 5020 3723
rect 5044 3717 5084 3723
rect 5220 3717 5244 3723
rect 5444 3717 5500 3723
rect 5588 3717 5708 3723
rect 5725 3717 5868 3723
rect 5725 3704 5731 3717
rect 5924 3717 6028 3723
rect 6036 3717 6092 3723
rect 6148 3717 6220 3723
rect 6324 3717 6348 3723
rect 6589 3723 6595 3757
rect 6589 3717 6604 3723
rect 6669 3723 6675 3743
rect 6669 3717 6691 3723
rect 180 3697 204 3703
rect 276 3697 348 3703
rect 356 3697 444 3703
rect 452 3697 508 3703
rect 516 3697 572 3703
rect 580 3697 684 3703
rect 1460 3697 1740 3703
rect 1748 3697 1772 3703
rect 1844 3697 1868 3703
rect 1876 3697 2076 3703
rect 2084 3697 2108 3703
rect 2404 3697 2492 3703
rect 2500 3697 2572 3703
rect 2868 3697 2892 3703
rect 3460 3697 3516 3703
rect 3556 3697 3580 3703
rect 3668 3697 3724 3703
rect 4116 3697 4156 3703
rect 4244 3697 4332 3703
rect 4452 3697 4524 3703
rect 4532 3697 4652 3703
rect 4756 3697 4972 3703
rect 4980 3697 5100 3703
rect 5396 3697 5452 3703
rect 5508 3697 5532 3703
rect 5604 3697 5724 3703
rect 5748 3697 5756 3703
rect 5812 3697 5884 3703
rect 5892 3697 5964 3703
rect 6052 3697 6188 3703
rect 6196 3697 6236 3703
rect 6628 3697 6675 3703
rect 1412 3677 1436 3683
rect 1444 3677 1596 3683
rect 1604 3677 1852 3683
rect 1860 3677 1996 3683
rect 2004 3677 2236 3683
rect 4164 3677 4188 3683
rect 4388 3677 4492 3683
rect 4500 3677 4620 3683
rect 5172 3677 5196 3683
rect 5204 3677 5260 3683
rect 5284 3677 5404 3683
rect 5428 3677 5436 3683
rect 5533 3683 5539 3696
rect 5533 3677 5628 3683
rect 5636 3677 5660 3683
rect 5828 3677 5948 3683
rect 5972 3677 5980 3683
rect 6036 3677 6268 3683
rect 6292 3677 6316 3683
rect 6685 3683 6691 3717
rect 6420 3677 6691 3683
rect 2036 3657 2156 3663
rect 2164 3657 2956 3663
rect 2964 3657 3820 3663
rect 4644 3657 4780 3663
rect 5108 3657 5340 3663
rect 5524 3657 5548 3663
rect 5556 3657 5612 3663
rect 5876 3657 5932 3663
rect 5972 3657 6076 3663
rect 6164 3657 6188 3663
rect 6228 3657 6300 3663
rect 6468 3657 6492 3663
rect 212 3637 2508 3643
rect 2548 3637 5356 3643
rect 5428 3637 5484 3643
rect 5492 3637 5644 3643
rect 5876 3637 6140 3643
rect 6292 3637 6444 3643
rect 6484 3637 6524 3643
rect 1460 3617 1484 3623
rect 4564 3617 4764 3623
rect 6100 3617 6124 3623
rect 6228 3617 6316 3623
rect 6404 3617 6620 3623
rect 1768 3614 1816 3616
rect 1768 3606 1772 3614
rect 1782 3606 1788 3614
rect 1796 3606 1802 3614
rect 1812 3606 1816 3614
rect 1768 3604 1816 3606
rect 4824 3614 4872 3616
rect 4824 3606 4828 3614
rect 4838 3606 4844 3614
rect 4852 3606 4858 3614
rect 4868 3606 4872 3614
rect 4824 3604 4872 3606
rect 3252 3597 3388 3603
rect 3396 3597 3692 3603
rect 4068 3597 4364 3603
rect 4980 3597 5788 3603
rect 5860 3597 5916 3603
rect 5924 3597 5964 3603
rect 6052 3597 6060 3603
rect 6068 3597 6092 3603
rect 6116 3597 6188 3603
rect 6324 3597 6508 3603
rect 692 3577 716 3583
rect 724 3577 748 3583
rect 1028 3577 1052 3583
rect 1892 3577 2556 3583
rect 2564 3577 2588 3583
rect 2644 3577 2700 3583
rect 2740 3577 2908 3583
rect 2916 3577 3404 3583
rect 3412 3577 4076 3583
rect 4516 3577 4924 3583
rect 5444 3577 5916 3583
rect 5981 3577 6156 3583
rect 420 3557 508 3563
rect 756 3557 2028 3563
rect 3476 3557 3724 3563
rect 4260 3557 4556 3563
rect 4628 3557 4748 3563
rect 5981 3563 5987 3577
rect 6260 3577 6332 3583
rect 5716 3557 5987 3563
rect 6068 3557 6092 3563
rect 6116 3557 6172 3563
rect 6228 3557 6332 3563
rect 6340 3557 6380 3563
rect 244 3537 524 3543
rect 788 3537 1116 3543
rect 2100 3537 2124 3543
rect 2164 3537 2204 3543
rect 2884 3537 2892 3543
rect 3028 3537 3116 3543
rect 3428 3537 3660 3543
rect 3764 3537 3948 3543
rect 3956 3537 4012 3543
rect 4020 3537 4092 3543
rect 4100 3537 4316 3543
rect 4388 3537 4396 3543
rect 4404 3537 4460 3543
rect 4564 3537 4732 3543
rect 4740 3537 5036 3543
rect 5508 3537 5580 3543
rect 5604 3537 5660 3543
rect 5812 3537 5868 3543
rect 5924 3537 6044 3543
rect 6100 3537 6156 3543
rect 6196 3537 6268 3543
rect 6356 3537 6460 3543
rect 6516 3537 6588 3543
rect 436 3517 524 3523
rect 852 3517 876 3523
rect 1028 3517 1100 3523
rect 1988 3517 2044 3523
rect 2052 3517 2188 3523
rect 2324 3517 2444 3523
rect 2564 3517 3036 3523
rect 3060 3517 3340 3523
rect 3380 3517 3532 3523
rect 3668 3517 4028 3523
rect 4036 3517 4060 3523
rect 4292 3517 4460 3523
rect 4484 3517 5068 3523
rect 5076 3517 5196 3523
rect 5236 3517 5388 3523
rect 5556 3517 5612 3523
rect 5620 3517 5628 3523
rect 5700 3517 5804 3523
rect 5844 3517 5932 3523
rect 6004 3517 6140 3523
rect 6228 3517 6556 3523
rect 84 3497 268 3503
rect 340 3497 604 3503
rect 612 3497 684 3503
rect 692 3497 1036 3503
rect 1044 3497 1068 3503
rect 1140 3497 1180 3503
rect 2132 3497 2188 3503
rect 2196 3497 2220 3503
rect 2468 3497 2524 3503
rect 2836 3497 2892 3503
rect 3028 3497 3084 3503
rect 3092 3497 3260 3503
rect 3268 3497 3436 3503
rect 3700 3497 3820 3503
rect 4244 3497 4492 3503
rect 4548 3497 4707 3503
rect 628 3477 652 3483
rect 804 3477 924 3483
rect 932 3477 988 3483
rect 1012 3477 1164 3483
rect 1620 3477 1660 3483
rect 1668 3477 1708 3483
rect 2004 3477 2028 3483
rect 2228 3477 2284 3483
rect 2356 3477 2428 3483
rect 2436 3477 2684 3483
rect 2788 3477 2860 3483
rect 2868 3477 2908 3483
rect 2916 3477 2988 3483
rect 2996 3477 3020 3483
rect 3396 3477 3468 3483
rect 3588 3477 3788 3483
rect 4500 3477 4620 3483
rect 4701 3483 4707 3497
rect 4724 3497 5052 3503
rect 5124 3497 5308 3503
rect 5332 3497 5420 3503
rect 5540 3497 5564 3503
rect 5588 3497 5644 3503
rect 5812 3497 5836 3503
rect 5860 3497 5916 3503
rect 5940 3497 6028 3503
rect 6132 3497 6348 3503
rect 6372 3497 6428 3503
rect 6532 3497 6556 3503
rect 4701 3477 4755 3483
rect 884 3457 940 3463
rect 1060 3457 1228 3463
rect 1524 3457 1692 3463
rect 1732 3457 1836 3463
rect 1844 3457 2140 3463
rect 2836 3457 2972 3463
rect 2980 3457 3676 3463
rect 3860 3457 3964 3463
rect 3972 3457 3996 3463
rect 4004 3457 4044 3463
rect 4228 3457 4300 3463
rect 4324 3457 4508 3463
rect 4548 3457 4700 3463
rect 4749 3463 4755 3477
rect 4772 3477 5180 3483
rect 5188 3477 5292 3483
rect 5364 3477 5612 3483
rect 5956 3477 6044 3483
rect 6349 3483 6355 3496
rect 6349 3477 6396 3483
rect 4749 3457 4796 3463
rect 4836 3457 5324 3463
rect 5428 3457 5452 3463
rect 5556 3457 5580 3463
rect 5636 3457 5740 3463
rect 5764 3457 5852 3463
rect 6004 3457 6028 3463
rect 6116 3457 6124 3463
rect 6132 3457 6204 3463
rect 6356 3457 6492 3463
rect 6500 3457 6540 3463
rect 6580 3457 6604 3463
rect 196 3437 220 3443
rect 388 3437 636 3443
rect 644 3437 812 3443
rect 884 3437 956 3443
rect 1716 3437 1820 3443
rect 1828 3437 2300 3443
rect 2340 3437 2524 3443
rect 2612 3437 2780 3443
rect 2964 3437 4028 3443
rect 4036 3437 4108 3443
rect 4164 3437 4284 3443
rect 4340 3437 4364 3443
rect 4829 3443 4835 3456
rect 4372 3437 4835 3443
rect 5428 3437 5484 3443
rect 5780 3437 5836 3443
rect 5908 3437 5948 3443
rect 6308 3437 6412 3443
rect 660 3417 892 3423
rect 948 3417 1276 3423
rect 1380 3417 1628 3423
rect 1652 3417 1916 3423
rect 1956 3417 2236 3423
rect 3892 3417 4140 3423
rect 4148 3417 4236 3423
rect 4596 3417 4652 3423
rect 4788 3417 4892 3423
rect 4964 3417 5132 3423
rect 5140 3417 5228 3423
rect 5476 3417 5772 3423
rect 5812 3417 5964 3423
rect 6196 3417 6460 3423
rect 6484 3417 6540 3423
rect 3304 3414 3352 3416
rect 3304 3406 3308 3414
rect 3318 3406 3324 3414
rect 3332 3406 3338 3414
rect 3348 3406 3352 3414
rect 3304 3404 3352 3406
rect 548 3397 844 3403
rect 932 3397 1196 3403
rect 1220 3397 1404 3403
rect 1876 3397 1916 3403
rect 1924 3397 2012 3403
rect 4052 3397 4156 3403
rect 4212 3397 4236 3403
rect 4852 3397 5116 3403
rect 5188 3397 5580 3403
rect 5588 3397 5660 3403
rect 5780 3397 6284 3403
rect 6452 3397 6572 3403
rect 852 3377 908 3383
rect 916 3377 1020 3383
rect 1076 3377 1260 3383
rect 1476 3377 1532 3383
rect 1540 3377 1852 3383
rect 1876 3377 1996 3383
rect 2212 3377 3148 3383
rect 3172 3377 3356 3383
rect 3364 3377 3660 3383
rect 3748 3377 4108 3383
rect 4148 3377 4972 3383
rect 5012 3377 5596 3383
rect 5604 3377 5644 3383
rect 5732 3377 5772 3383
rect 5796 3377 6659 3383
rect 420 3357 540 3363
rect 564 3357 764 3363
rect 964 3357 1244 3363
rect 1252 3357 1308 3363
rect 1572 3357 1596 3363
rect 1604 3357 1740 3363
rect 1940 3357 2124 3363
rect 2548 3357 2572 3363
rect 2580 3357 2668 3363
rect 2900 3357 2956 3363
rect 4100 3357 4268 3363
rect 4276 3357 4316 3363
rect 4676 3357 4780 3363
rect 4788 3357 4940 3363
rect 5028 3357 5100 3363
rect 5108 3357 5244 3363
rect 5316 3357 5372 3363
rect 5380 3357 5532 3363
rect 5604 3357 5788 3363
rect 6052 3357 6092 3363
rect 6164 3357 6316 3363
rect 6324 3357 6428 3363
rect 20 3337 44 3343
rect 132 3337 172 3343
rect 484 3337 524 3343
rect 596 3337 748 3343
rect 1044 3337 1132 3343
rect 1204 3337 1516 3343
rect 1620 3337 1644 3343
rect 1748 3337 3619 3343
rect 3613 3324 3619 3337
rect 3908 3337 3980 3343
rect 3988 3337 4076 3343
rect 4269 3337 4412 3343
rect 4269 3324 4275 3337
rect 4948 3337 5004 3343
rect 5012 3337 5068 3343
rect 5380 3337 5468 3343
rect 5556 3337 5676 3343
rect 5684 3337 5836 3343
rect 5908 3337 5932 3343
rect 5988 3337 6092 3343
rect 6100 3337 6124 3343
rect 6180 3337 6220 3343
rect 6532 3337 6604 3343
rect 388 3317 460 3323
rect 532 3317 636 3323
rect 804 3317 892 3323
rect 996 3317 1068 3323
rect 1444 3317 1484 3323
rect 1508 3317 1772 3323
rect 1812 3317 1852 3323
rect 2052 3317 2156 3323
rect 2308 3317 2492 3323
rect 2660 3317 2764 3323
rect 2900 3317 3068 3323
rect 3124 3317 3164 3323
rect 3796 3317 3852 3323
rect 3876 3317 3916 3323
rect 3924 3317 4124 3323
rect 4244 3317 4268 3323
rect 4340 3317 4412 3323
rect 4532 3317 4636 3323
rect 4644 3317 4684 3323
rect 4692 3317 4748 3323
rect 4836 3317 4892 3323
rect 4900 3317 4940 3323
rect 5156 3317 5228 3323
rect 5444 3317 5708 3323
rect 5748 3317 5900 3323
rect 5924 3317 5964 3323
rect 5988 3317 6012 3323
rect 6356 3317 6572 3323
rect 6653 3323 6659 3377
rect 6669 3337 6691 3343
rect 6653 3317 6675 3323
rect 468 3297 572 3303
rect 580 3297 652 3303
rect 708 3297 924 3303
rect 932 3297 972 3303
rect 980 3297 1036 3303
rect 1364 3297 1452 3303
rect 1508 3297 1548 3303
rect 1668 3297 1724 3303
rect 1828 3297 1948 3303
rect 2020 3297 2060 3303
rect 2068 3297 2156 3303
rect 2164 3297 2220 3303
rect 2484 3297 2508 3303
rect 2516 3297 2652 3303
rect 2660 3297 2668 3303
rect 3812 3297 4028 3303
rect 4036 3297 4092 3303
rect 4132 3297 4156 3303
rect 4452 3297 4588 3303
rect 4660 3297 4700 3303
rect 4836 3297 5148 3303
rect 5236 3297 5292 3303
rect 5300 3297 5324 3303
rect 5332 3297 5420 3303
rect 5444 3297 5612 3303
rect 5684 3297 5820 3303
rect 5908 3297 5964 3303
rect 6004 3297 6044 3303
rect 6052 3297 6140 3303
rect 6164 3297 6220 3303
rect 6436 3297 6620 3303
rect 6669 3297 6675 3317
rect 788 3277 828 3283
rect 1396 3277 1516 3283
rect 2452 3277 2860 3283
rect 3780 3277 3836 3283
rect 3860 3277 3996 3283
rect 4052 3277 4172 3283
rect 4180 3277 4252 3283
rect 4260 3277 4284 3283
rect 4420 3277 4620 3283
rect 4628 3277 4732 3283
rect 5012 3277 5052 3283
rect 5076 3277 5276 3283
rect 5284 3277 5340 3283
rect 5348 3277 5404 3283
rect 6036 3277 6204 3283
rect 6685 3283 6691 3337
rect 6292 3277 6691 3283
rect 1492 3257 1676 3263
rect 2228 3257 2556 3263
rect 2564 3257 2764 3263
rect 2772 3257 2844 3263
rect 3828 3257 3980 3263
rect 3988 3257 4204 3263
rect 4324 3257 4444 3263
rect 4468 3257 4540 3263
rect 4788 3257 4988 3263
rect 5140 3257 5164 3263
rect 5172 3257 5212 3263
rect 5300 3257 5420 3263
rect 5428 3257 5500 3263
rect 6132 3257 6188 3263
rect 884 3237 2332 3243
rect 3108 3237 3228 3243
rect 3693 3237 3996 3243
rect 3693 3224 3699 3237
rect 4004 3237 4220 3243
rect 4228 3237 4236 3243
rect 4253 3237 4572 3243
rect 1220 3217 1372 3223
rect 1396 3217 1740 3223
rect 2836 3217 3692 3223
rect 4253 3223 4259 3237
rect 4596 3237 4652 3243
rect 4708 3237 4812 3243
rect 4820 3237 4924 3243
rect 4948 3237 6236 3243
rect 3732 3217 4259 3223
rect 4292 3217 4476 3223
rect 4484 3217 4524 3223
rect 5828 3217 5884 3223
rect 6132 3217 6268 3223
rect 6324 3217 6364 3223
rect 6516 3217 6716 3223
rect 1768 3214 1816 3216
rect 1768 3206 1772 3214
rect 1782 3206 1788 3214
rect 1796 3206 1802 3214
rect 1812 3206 1816 3214
rect 1768 3204 1816 3206
rect 4824 3214 4872 3216
rect 4824 3206 4828 3214
rect 4838 3206 4844 3214
rect 4852 3206 4858 3214
rect 4868 3206 4872 3214
rect 4824 3204 4872 3206
rect 932 3197 1587 3203
rect 196 3177 204 3183
rect 580 3177 1388 3183
rect 1412 3177 1564 3183
rect 1581 3183 1587 3197
rect 1837 3197 4124 3203
rect 1837 3183 1843 3197
rect 4180 3197 4364 3203
rect 4372 3197 4396 3203
rect 4420 3197 4556 3203
rect 4644 3197 4684 3203
rect 4692 3197 4748 3203
rect 4916 3197 5660 3203
rect 5988 3197 6172 3203
rect 6324 3197 6716 3203
rect 1581 3177 1843 3183
rect 3460 3177 4028 3183
rect 4036 3177 4044 3183
rect 4068 3177 4540 3183
rect 4580 3177 4940 3183
rect 5044 3177 5116 3183
rect 6004 3177 6028 3183
rect 6308 3177 6380 3183
rect 6500 3177 6604 3183
rect 676 3157 812 3163
rect 1380 3157 1548 3163
rect 1556 3157 1612 3163
rect 2500 3157 2604 3163
rect 2612 3157 2764 3163
rect 3108 3157 3148 3163
rect 3844 3157 4428 3163
rect 4628 3157 4668 3163
rect 4772 3157 5068 3163
rect 5076 3157 5116 3163
rect 5124 3157 5180 3163
rect 5636 3157 5740 3163
rect 5748 3157 5788 3163
rect 5924 3157 6620 3163
rect 772 3137 1676 3143
rect 1844 3137 2348 3143
rect 2356 3137 2732 3143
rect 2804 3137 3132 3143
rect 3268 3137 3452 3143
rect 3716 3137 3756 3143
rect 3773 3137 3900 3143
rect 868 3117 1100 3123
rect 1300 3117 1324 3123
rect 1396 3117 1484 3123
rect 1716 3117 1756 3123
rect 2644 3117 2828 3123
rect 2868 3117 2940 3123
rect 2964 3117 3724 3123
rect 3773 3123 3779 3137
rect 4244 3137 4268 3143
rect 4292 3137 4332 3143
rect 4413 3137 4556 3143
rect 4413 3124 4419 3137
rect 4564 3137 4620 3143
rect 4644 3137 4700 3143
rect 4724 3137 4812 3143
rect 4820 3137 4924 3143
rect 4932 3137 5020 3143
rect 5572 3137 5692 3143
rect 5732 3137 5820 3143
rect 5972 3137 6099 3143
rect 3748 3117 3779 3123
rect 3796 3117 3852 3123
rect 3876 3117 3884 3123
rect 3988 3117 4012 3123
rect 4020 3117 4108 3123
rect 4132 3117 4364 3123
rect 4388 3117 4412 3123
rect 4500 3117 4556 3123
rect 4580 3117 4796 3123
rect 4804 3117 4940 3123
rect 5588 3117 5996 3123
rect 6093 3123 6099 3137
rect 6116 3137 6140 3143
rect 6516 3137 6556 3143
rect 6093 3117 6156 3123
rect 6180 3117 6188 3123
rect 6276 3117 6460 3123
rect 308 3097 364 3103
rect 740 3097 796 3103
rect 1060 3097 1100 3103
rect 1156 3097 1260 3103
rect 1348 3097 1436 3103
rect 1636 3097 1740 3103
rect 1988 3097 2028 3103
rect 2164 3097 2252 3103
rect 2308 3097 2508 3103
rect 2580 3097 2700 3103
rect 3156 3097 3324 3103
rect 3668 3097 4044 3103
rect 4340 3097 4380 3103
rect 4436 3097 4460 3103
rect 4468 3097 4572 3103
rect 4580 3097 4636 3103
rect 4708 3097 4764 3103
rect 4980 3097 5052 3103
rect 5060 3097 5132 3103
rect 5140 3097 5164 3103
rect 5332 3097 5388 3103
rect 5524 3097 5564 3103
rect 5572 3097 5612 3103
rect 5677 3097 5916 3103
rect 132 3077 332 3083
rect 1044 3077 1132 3083
rect 1252 3077 1292 3083
rect 1300 3077 1356 3083
rect 1364 3077 1404 3083
rect 1476 3077 1516 3083
rect 1540 3077 1724 3083
rect 1972 3077 2060 3083
rect 2116 3077 2332 3083
rect 2468 3077 2508 3083
rect 2516 3077 2604 3083
rect 3028 3077 3116 3083
rect 3396 3077 3484 3083
rect 3764 3077 3804 3083
rect 3892 3077 3932 3083
rect 4004 3077 4092 3083
rect 4132 3077 4396 3083
rect 4429 3077 4492 3083
rect 548 3057 604 3063
rect 612 3057 700 3063
rect 740 3057 796 3063
rect 980 3057 1068 3063
rect 1780 3057 2092 3063
rect 2109 3057 2956 3063
rect 2109 3043 2115 3057
rect 2996 3057 3180 3063
rect 3188 3057 3532 3063
rect 4429 3063 4435 3077
rect 4516 3077 4780 3083
rect 5076 3077 5292 3083
rect 5677 3083 5683 3097
rect 6036 3097 6076 3103
rect 6525 3097 6572 3103
rect 5460 3077 5683 3083
rect 5700 3077 5740 3083
rect 5796 3077 5932 3083
rect 5972 3077 6044 3083
rect 6164 3077 6188 3083
rect 6525 3064 6531 3097
rect 6596 3097 6611 3103
rect 3796 3057 4435 3063
rect 4468 3057 4588 3063
rect 4612 3057 5068 3063
rect 5156 3057 5212 3063
rect 5236 3057 5276 3063
rect 5540 3057 5644 3063
rect 5716 3057 5772 3063
rect 5780 3057 5852 3063
rect 5908 3057 6476 3063
rect 6605 3044 6611 3097
rect 6628 3097 6675 3103
rect 500 3037 2115 3043
rect 2228 3037 2396 3043
rect 2420 3037 2476 3043
rect 2484 3037 2828 3043
rect 2836 3037 2908 3043
rect 3060 3037 3100 3043
rect 3108 3037 3372 3043
rect 3748 3037 4508 3043
rect 4532 3037 4716 3043
rect 4724 3037 4908 3043
rect 4916 3037 4972 3043
rect 4996 3037 5404 3043
rect 5620 3037 5628 3043
rect 5652 3037 5884 3043
rect 5892 3037 6076 3043
rect 6388 3037 6476 3043
rect 6516 3037 6588 3043
rect 100 3017 300 3023
rect 308 3017 588 3023
rect 596 3017 620 3023
rect 1092 3017 1164 3023
rect 1860 3017 2428 3023
rect 2756 3017 2988 3023
rect 3924 3017 3964 3023
rect 3972 3017 4220 3023
rect 4308 3017 5587 3023
rect 3304 3014 3352 3016
rect 3304 3006 3308 3014
rect 3318 3006 3324 3014
rect 3332 3006 3338 3014
rect 3348 3006 3352 3014
rect 3304 3004 3352 3006
rect 516 2997 540 3003
rect 692 2997 1932 3003
rect 1988 2997 2924 3003
rect 2932 2997 2956 3003
rect 3700 2997 3996 3003
rect 4020 2997 4060 3003
rect 4084 2997 4252 3003
rect 4260 2997 4364 3003
rect 4388 2997 4988 3003
rect 5028 2997 5404 3003
rect 5508 2997 5564 3003
rect 5581 3003 5587 3017
rect 5604 3017 5900 3023
rect 5956 3017 6028 3023
rect 6036 3017 6092 3023
rect 6340 3017 6508 3023
rect 6580 3017 6636 3023
rect 5581 2997 5804 3003
rect 5828 2997 5948 3003
rect 6020 2997 6156 3003
rect 6500 2997 6620 3003
rect 996 2977 1228 2983
rect 1348 2977 1916 2983
rect 2004 2977 2476 2983
rect 2484 2977 2524 2983
rect 2692 2977 2732 2983
rect 2740 2977 3020 2983
rect 3028 2977 3084 2983
rect 3092 2977 3212 2983
rect 3572 2977 3756 2983
rect 3764 2977 4028 2983
rect 4084 2977 4556 2983
rect 4564 2977 4652 2983
rect 4660 2977 4796 2983
rect 5364 2977 5452 2983
rect 5460 2977 5852 2983
rect 5860 2977 5884 2983
rect 5924 2977 6044 2983
rect 6468 2977 6492 2983
rect 68 2957 323 2963
rect 317 2944 323 2957
rect 644 2957 716 2963
rect 852 2957 1004 2963
rect 1268 2957 1548 2963
rect 1620 2957 1948 2963
rect 1972 2957 2012 2963
rect 2068 2957 2092 2963
rect 2772 2957 2780 2963
rect 2820 2957 2860 2963
rect 3556 2957 3875 2963
rect 52 2937 108 2943
rect 180 2937 204 2943
rect 324 2937 428 2943
rect 500 2937 524 2943
rect 532 2937 700 2943
rect 708 2937 748 2943
rect 756 2937 812 2943
rect 820 2937 940 2943
rect 1220 2937 1260 2943
rect 1588 2937 1868 2943
rect 1908 2937 1996 2943
rect 2013 2937 2284 2943
rect 52 2917 172 2923
rect 276 2917 332 2923
rect 388 2917 428 2923
rect 452 2917 524 2923
rect 548 2917 588 2923
rect 612 2917 652 2923
rect 948 2917 972 2923
rect 1124 2917 1196 2923
rect 1428 2917 1516 2923
rect 1524 2917 1580 2923
rect 2013 2923 2019 2937
rect 2388 2937 2460 2943
rect 2660 2937 2716 2943
rect 2884 2937 3004 2943
rect 3508 2937 3628 2943
rect 3700 2937 3852 2943
rect 3869 2943 3875 2957
rect 3908 2957 4524 2963
rect 4532 2957 4588 2963
rect 4628 2957 5020 2963
rect 5396 2957 5484 2963
rect 5492 2957 5548 2963
rect 5572 2957 5612 2963
rect 5652 2957 5756 2963
rect 5780 2957 5804 2963
rect 5844 2957 5964 2963
rect 3869 2937 4012 2943
rect 4052 2937 4156 2943
rect 4164 2937 4268 2943
rect 4340 2937 4492 2943
rect 4516 2937 4572 2943
rect 4724 2937 4748 2943
rect 4756 2937 4812 2943
rect 4884 2937 4924 2943
rect 5060 2937 5164 2943
rect 5172 2937 5356 2943
rect 5364 2937 5420 2943
rect 5556 2937 5708 2943
rect 5764 2937 5788 2943
rect 5876 2937 6028 2943
rect 6036 2937 6060 2943
rect 6068 2937 6108 2943
rect 6388 2937 6444 2943
rect 6644 2937 6675 2943
rect 1812 2917 2019 2923
rect 2212 2917 2268 2923
rect 2340 2917 2476 2923
rect 2516 2917 2716 2923
rect 2868 2917 2892 2923
rect 3188 2917 3244 2923
rect 3540 2917 3820 2923
rect 3828 2917 4076 2923
rect 4244 2917 4412 2923
rect 4420 2917 4460 2923
rect 4660 2917 4732 2923
rect 4756 2917 4940 2923
rect 4980 2917 5212 2923
rect 5220 2917 5276 2923
rect 5284 2917 5308 2923
rect 5364 2917 5516 2923
rect 5524 2917 5564 2923
rect 5652 2917 5756 2923
rect 5764 2917 5804 2923
rect 5812 2917 5900 2923
rect 6004 2917 6012 2923
rect 196 2897 252 2903
rect 260 2897 380 2903
rect 772 2897 780 2903
rect 788 2897 1260 2903
rect 1364 2897 1516 2903
rect 1524 2897 2076 2903
rect 2244 2897 2268 2903
rect 2292 2897 3388 2903
rect 3476 2897 4300 2903
rect 4340 2897 4396 2903
rect 4404 2897 4492 2903
rect 4500 2897 5004 2903
rect 5028 2897 5052 2903
rect 5140 2897 5196 2903
rect 5204 2897 5244 2903
rect 5268 2897 5459 2903
rect 36 2877 156 2883
rect 164 2877 172 2883
rect 196 2877 252 2883
rect 292 2877 316 2883
rect 356 2877 444 2883
rect 452 2877 684 2883
rect 692 2877 716 2883
rect 740 2877 828 2883
rect 964 2877 1020 2883
rect 1396 2877 1612 2883
rect 1700 2877 2140 2883
rect 2324 2877 2508 2883
rect 2676 2877 3180 2883
rect 3188 2877 3260 2883
rect 3828 2877 3836 2883
rect 3956 2877 4716 2883
rect 4756 2877 5228 2883
rect 5236 2877 5292 2883
rect 5300 2877 5340 2883
rect 5453 2883 5459 2897
rect 5476 2897 5532 2903
rect 5588 2897 5724 2903
rect 5796 2897 5868 2903
rect 5892 2897 5932 2903
rect 6436 2897 6675 2903
rect 5453 2877 5596 2883
rect 5652 2877 6540 2883
rect 20 2857 1500 2863
rect 1508 2857 1836 2863
rect 2036 2857 2060 2863
rect 2100 2857 3436 2863
rect 3812 2857 3884 2863
rect 4180 2857 4403 2863
rect 132 2837 188 2843
rect 244 2837 332 2843
rect 420 2837 636 2843
rect 644 2837 668 2843
rect 916 2837 924 2843
rect 932 2837 1068 2843
rect 1460 2837 1676 2843
rect 2084 2837 2124 2843
rect 2452 2837 3772 2843
rect 4397 2843 4403 2857
rect 4420 2857 4764 2863
rect 4772 2857 4828 2863
rect 5220 2857 5548 2863
rect 5572 2857 5676 2863
rect 5812 2857 6636 2863
rect 4397 2837 4620 2843
rect 4644 2837 4716 2843
rect 4740 2837 6252 2843
rect 20 2817 44 2823
rect 708 2817 1116 2823
rect 2084 2817 2444 2823
rect 2468 2817 2492 2823
rect 2500 2817 2892 2823
rect 2900 2817 3116 2823
rect 3652 2817 4140 2823
rect 4532 2817 4700 2823
rect 5700 2817 6188 2823
rect 1768 2814 1816 2816
rect 1768 2806 1772 2814
rect 1782 2806 1788 2814
rect 1796 2806 1802 2814
rect 1812 2806 1816 2814
rect 1768 2804 1816 2806
rect 4824 2814 4872 2816
rect 4824 2806 4828 2814
rect 4838 2806 4844 2814
rect 4852 2806 4858 2814
rect 4868 2806 4872 2814
rect 4824 2804 4872 2806
rect 276 2797 300 2803
rect 500 2797 540 2803
rect 932 2797 1116 2803
rect 2164 2797 2540 2803
rect 2644 2797 2700 2803
rect 2804 2797 3036 2803
rect 980 2777 1324 2783
rect 1668 2777 2796 2783
rect 4500 2777 4956 2783
rect 6228 2777 6252 2783
rect 6372 2777 6396 2783
rect 6500 2777 6556 2783
rect 1044 2757 1052 2763
rect 1060 2757 1116 2763
rect 1124 2757 1260 2763
rect 1716 2757 2092 2763
rect 2116 2757 4908 2763
rect 100 2737 172 2743
rect 596 2737 620 2743
rect 852 2737 1292 2743
rect 1572 2737 2515 2743
rect 260 2717 364 2723
rect 404 2717 524 2723
rect 1188 2717 1244 2723
rect 1924 2717 2092 2723
rect 2196 2717 2332 2723
rect 2509 2723 2515 2737
rect 2532 2737 2620 2743
rect 3060 2737 3836 2743
rect 4276 2737 5948 2743
rect 2509 2717 2764 2723
rect 2948 2717 2956 2723
rect 2964 2717 3004 2723
rect 3108 2717 3212 2723
rect 3252 2717 3692 2723
rect 4148 2717 4268 2723
rect 4356 2717 4444 2723
rect 4484 2717 4540 2723
rect 4932 2717 5324 2723
rect 5460 2717 5731 2723
rect 196 2697 220 2703
rect 500 2697 796 2703
rect 868 2697 876 2703
rect 884 2697 972 2703
rect 1076 2697 1132 2703
rect 1140 2697 1356 2703
rect 1396 2697 1564 2703
rect 1636 2697 1756 2703
rect 2004 2697 2092 2703
rect 2196 2697 2300 2703
rect 2340 2697 2460 2703
rect 2484 2697 2588 2703
rect 2740 2697 2796 2703
rect 3060 2697 3132 2703
rect 3284 2697 3564 2703
rect 3972 2697 4156 2703
rect 4340 2697 4508 2703
rect 4596 2697 4716 2703
rect 4964 2697 4988 2703
rect 5076 2697 5132 2703
rect 5181 2697 5516 2703
rect 436 2677 476 2683
rect 484 2677 524 2683
rect 628 2677 716 2683
rect 740 2677 764 2683
rect 1028 2677 1084 2683
rect 1124 2677 1228 2683
rect 1332 2677 1372 2683
rect 1380 2677 1484 2683
rect 1732 2677 1868 2683
rect 1876 2677 1948 2683
rect 1956 2677 2028 2683
rect 2036 2677 2140 2683
rect 2516 2677 2636 2683
rect 2788 2677 2812 2683
rect 2996 2677 3068 2683
rect 3076 2677 3148 2683
rect 3316 2677 3404 2683
rect 3764 2677 3916 2683
rect 4132 2677 4156 2683
rect 4164 2677 4204 2683
rect 4212 2677 4300 2683
rect 4324 2677 4364 2683
rect 4436 2677 4492 2683
rect 4500 2677 4524 2683
rect 5181 2683 5187 2697
rect 5636 2697 5708 2703
rect 5725 2703 5731 2717
rect 6084 2717 6380 2723
rect 6516 2717 6636 2723
rect 5725 2697 6140 2703
rect 6180 2697 6675 2703
rect 4756 2677 5187 2683
rect 5204 2677 5292 2683
rect 6020 2677 6204 2683
rect 6212 2677 6444 2683
rect 180 2657 252 2663
rect 548 2657 668 2663
rect 692 2657 812 2663
rect 996 2657 1036 2663
rect 1108 2657 1196 2663
rect 1508 2657 1692 2663
rect 2708 2657 2732 2663
rect 2756 2657 2988 2663
rect 3156 2657 3308 2663
rect 3396 2657 3452 2663
rect 4084 2657 4172 2663
rect 4180 2657 4204 2663
rect 4244 2657 4316 2663
rect 4324 2657 4348 2663
rect 4500 2657 4572 2663
rect 4788 2657 5100 2663
rect 6004 2657 6620 2663
rect 84 2637 332 2643
rect 724 2637 780 2643
rect 1060 2637 1212 2643
rect 1332 2637 1436 2643
rect 1444 2637 1532 2643
rect 1540 2637 1996 2643
rect 2420 2637 3548 2643
rect 3572 2637 3820 2643
rect 4660 2637 4844 2643
rect 4852 2637 4908 2643
rect 4996 2637 5164 2643
rect 5844 2637 5868 2643
rect 6164 2637 6268 2643
rect 884 2617 1004 2623
rect 1012 2617 1180 2623
rect 1220 2617 1276 2623
rect 1764 2617 1916 2623
rect 1972 2617 3036 2623
rect 3044 2617 3132 2623
rect 3412 2617 3628 2623
rect 3876 2617 4076 2623
rect 4100 2617 4140 2623
rect 4180 2617 4236 2623
rect 4244 2617 4284 2623
rect 4292 2617 4428 2623
rect 4628 2617 4876 2623
rect 3304 2614 3352 2616
rect 3304 2606 3308 2614
rect 3318 2606 3324 2614
rect 3332 2606 3338 2614
rect 3348 2606 3352 2614
rect 3304 2604 3352 2606
rect 580 2597 636 2603
rect 644 2597 668 2603
rect 1636 2597 1788 2603
rect 1876 2597 2627 2603
rect 2621 2584 2627 2597
rect 2980 2597 3148 2603
rect 3556 2597 4940 2603
rect 4948 2597 6236 2603
rect 820 2577 867 2583
rect 861 2564 867 2577
rect 900 2577 908 2583
rect 1412 2577 2412 2583
rect 2436 2577 2595 2583
rect 2589 2564 2595 2577
rect 2628 2577 2652 2583
rect 2676 2577 2796 2583
rect 2820 2577 3052 2583
rect 3060 2577 3116 2583
rect 3124 2577 3180 2583
rect 3268 2577 3532 2583
rect 3668 2577 3852 2583
rect 3924 2577 4060 2583
rect 4116 2577 4220 2583
rect 4724 2577 5004 2583
rect 5044 2577 5196 2583
rect 5204 2577 5260 2583
rect 5284 2577 5324 2583
rect 6036 2577 6092 2583
rect 6548 2577 6604 2583
rect 228 2557 268 2563
rect 276 2557 284 2563
rect 292 2557 316 2563
rect 452 2557 828 2563
rect 868 2557 1004 2563
rect 1044 2557 1164 2563
rect 1188 2557 1276 2563
rect 1284 2557 1340 2563
rect 2132 2557 2204 2563
rect 2228 2557 2396 2563
rect 2404 2557 2444 2563
rect 2500 2557 2540 2563
rect 2596 2557 2684 2563
rect 2692 2557 2748 2563
rect 2836 2557 2876 2563
rect 3332 2557 3516 2563
rect 3524 2557 3916 2563
rect 3940 2557 4012 2563
rect 4116 2557 4332 2563
rect 4372 2557 4428 2563
rect 4452 2557 4764 2563
rect 5172 2557 5276 2563
rect 20 2537 108 2543
rect 132 2537 236 2543
rect 244 2537 268 2543
rect 292 2537 428 2543
rect 484 2537 524 2543
rect 548 2537 652 2543
rect 692 2537 732 2543
rect 740 2537 844 2543
rect 980 2537 1116 2543
rect 1124 2537 1324 2543
rect 2036 2537 2236 2543
rect 2628 2537 2684 2543
rect 2836 2537 2892 2543
rect 2900 2537 2924 2543
rect 2932 2537 2940 2543
rect 2948 2537 2988 2543
rect 3172 2537 3196 2543
rect 3460 2537 3612 2543
rect 3620 2537 3692 2543
rect 4020 2537 4348 2543
rect 4356 2537 4476 2543
rect 4596 2537 4652 2543
rect 4948 2537 4956 2543
rect 5012 2537 5180 2543
rect 5492 2537 5644 2543
rect 5652 2537 5676 2543
rect 196 2517 236 2523
rect 372 2517 492 2523
rect 500 2517 732 2523
rect 996 2517 1052 2523
rect 1092 2517 1132 2523
rect 1156 2517 1292 2523
rect 1428 2517 1516 2523
rect 1572 2517 2076 2523
rect 2116 2517 2236 2523
rect 2244 2517 2460 2523
rect 2468 2517 2476 2523
rect 2484 2517 2508 2523
rect 2532 2517 2636 2523
rect 2644 2517 2732 2523
rect 2740 2517 2780 2523
rect 2804 2517 2908 2523
rect 3092 2517 3164 2523
rect 3252 2517 3388 2523
rect 3444 2517 3580 2523
rect 3604 2517 3724 2523
rect 3988 2517 4044 2523
rect 4052 2517 4188 2523
rect 4212 2517 4300 2523
rect 4308 2517 4572 2523
rect 4596 2517 4604 2523
rect 4644 2517 4668 2523
rect 4708 2517 4748 2523
rect 4756 2517 4972 2523
rect 5300 2517 5420 2523
rect 5524 2517 5580 2523
rect 5812 2517 5900 2523
rect 6212 2517 6476 2523
rect 116 2497 204 2503
rect 532 2497 604 2503
rect 1204 2497 1372 2503
rect 2164 2497 2188 2503
rect 2324 2497 2556 2503
rect 2756 2497 2828 2503
rect 3028 2497 3244 2503
rect 3252 2497 3516 2503
rect 3524 2497 3532 2503
rect 3636 2497 3836 2503
rect 3844 2497 3948 2503
rect 4004 2497 4108 2503
rect 4212 2497 4556 2503
rect 4564 2497 4572 2503
rect 4580 2497 5068 2503
rect 5076 2497 5308 2503
rect 5316 2497 5580 2503
rect 5684 2497 6220 2503
rect 6228 2497 6284 2503
rect 436 2477 588 2483
rect 596 2477 684 2483
rect 2100 2477 3100 2483
rect 3108 2477 3196 2483
rect 4260 2477 4396 2483
rect 4404 2477 4444 2483
rect 4500 2477 4652 2483
rect 4676 2477 4803 2483
rect 52 2457 140 2463
rect 260 2457 300 2463
rect 340 2457 364 2463
rect 2404 2457 2492 2463
rect 2500 2457 2732 2463
rect 2900 2457 3068 2463
rect 4196 2457 4460 2463
rect 4468 2457 4524 2463
rect 4548 2457 4780 2463
rect 4797 2463 4803 2477
rect 4932 2477 5084 2483
rect 5492 2477 5708 2483
rect 4797 2457 5132 2463
rect 180 2437 300 2443
rect 804 2437 844 2443
rect 852 2437 956 2443
rect 964 2437 1388 2443
rect 2148 2437 3484 2443
rect 4276 2437 5132 2443
rect 2004 2417 2508 2423
rect 2708 2417 4732 2423
rect 5044 2417 5100 2423
rect 1768 2414 1816 2416
rect 1768 2406 1772 2414
rect 1782 2406 1788 2414
rect 1796 2406 1802 2414
rect 1812 2406 1816 2414
rect 1768 2404 1816 2406
rect 4824 2414 4872 2416
rect 4824 2406 4828 2414
rect 4838 2406 4844 2414
rect 4852 2406 4858 2414
rect 4868 2406 4872 2414
rect 4824 2404 4872 2406
rect 2452 2397 3436 2403
rect 4372 2397 4748 2403
rect 1732 2377 2828 2383
rect 3684 2377 3916 2383
rect 4100 2377 4300 2383
rect 4308 2377 4716 2383
rect 196 2357 268 2363
rect 420 2357 604 2363
rect 1476 2357 1884 2363
rect 2868 2357 3100 2363
rect 3140 2357 3356 2363
rect 3828 2357 4780 2363
rect 4788 2357 5116 2363
rect 5124 2357 5228 2363
rect 5236 2357 5420 2363
rect 5460 2357 5596 2363
rect 5652 2357 5772 2363
rect 6372 2357 6412 2363
rect 132 2337 188 2343
rect 196 2337 236 2343
rect 244 2337 444 2343
rect 468 2337 492 2343
rect 2484 2337 2700 2343
rect 2788 2337 2892 2343
rect 2932 2337 3148 2343
rect 3380 2337 4140 2343
rect 4148 2337 4412 2343
rect 4516 2337 4620 2343
rect 4628 2337 4636 2343
rect 4804 2337 4972 2343
rect 5300 2337 5436 2343
rect 5444 2337 5516 2343
rect 6132 2337 6140 2343
rect 20 2317 172 2323
rect 292 2317 700 2323
rect 932 2317 972 2323
rect 980 2317 1036 2323
rect 1076 2317 1420 2323
rect 1428 2317 1500 2323
rect 1924 2317 2028 2323
rect 2068 2317 2156 2323
rect 2388 2317 2460 2323
rect 2468 2317 2524 2323
rect 2532 2317 2604 2323
rect 2692 2317 2764 2323
rect 2772 2317 3020 2323
rect 3140 2317 3164 2323
rect 3204 2317 3484 2323
rect 3540 2317 4252 2323
rect 4292 2317 4332 2323
rect 4356 2317 4700 2323
rect 4948 2317 5468 2323
rect 6020 2317 6156 2323
rect 52 2297 172 2303
rect 180 2297 252 2303
rect 260 2297 524 2303
rect 1044 2297 1116 2303
rect 1348 2297 1404 2303
rect 1412 2297 1436 2303
rect 1588 2297 1676 2303
rect 1684 2297 1996 2303
rect 2004 2297 2012 2303
rect 2020 2297 2108 2303
rect 2308 2297 2428 2303
rect 2660 2297 2716 2303
rect 2772 2297 2812 2303
rect 2900 2297 2956 2303
rect 2964 2297 3180 2303
rect 3300 2297 3388 2303
rect 3588 2297 3612 2303
rect 3828 2297 3884 2303
rect 3972 2297 4044 2303
rect 4052 2297 4316 2303
rect 4324 2297 4364 2303
rect 4484 2297 4588 2303
rect 4644 2297 4732 2303
rect 4804 2297 4876 2303
rect 5412 2297 5452 2303
rect 6116 2297 6188 2303
rect 308 2277 364 2283
rect 372 2277 604 2283
rect 772 2277 876 2283
rect 900 2277 908 2283
rect 916 2277 940 2283
rect 1172 2277 1212 2283
rect 1508 2277 1516 2283
rect 3076 2277 3116 2283
rect 3220 2277 3260 2283
rect 3492 2277 3532 2283
rect 4036 2277 4396 2283
rect 4404 2277 4460 2283
rect 4532 2277 5004 2283
rect 5076 2277 5116 2283
rect 5124 2277 5164 2283
rect 5172 2277 5276 2283
rect 5284 2277 5372 2283
rect 5380 2277 5452 2283
rect 5716 2277 5740 2283
rect 164 2257 348 2263
rect 356 2257 716 2263
rect 724 2257 956 2263
rect 1060 2257 1228 2263
rect 1332 2257 1372 2263
rect 1380 2257 1484 2263
rect 2724 2257 2892 2263
rect 2948 2257 3244 2263
rect 3252 2257 3276 2263
rect 3364 2257 3420 2263
rect 3444 2257 3500 2263
rect 3540 2257 3548 2263
rect 3556 2257 3804 2263
rect 3924 2257 3964 2263
rect 4116 2257 4236 2263
rect 4260 2257 4524 2263
rect 4861 2257 5148 2263
rect 4861 2244 4867 2257
rect 5156 2257 5212 2263
rect 6148 2257 6204 2263
rect 6212 2257 6460 2263
rect 420 2237 460 2243
rect 516 2237 572 2243
rect 580 2237 636 2243
rect 676 2237 732 2243
rect 836 2237 860 2243
rect 884 2237 908 2243
rect 964 2237 1004 2243
rect 1796 2237 1868 2243
rect 1876 2237 1980 2243
rect 2180 2237 2364 2243
rect 2836 2237 2940 2243
rect 2948 2237 2972 2243
rect 3060 2237 3756 2243
rect 3764 2237 3788 2243
rect 3796 2237 4044 2243
rect 4052 2237 4588 2243
rect 4676 2237 4860 2243
rect 5828 2237 6236 2243
rect 6244 2237 6252 2243
rect 6260 2237 6428 2243
rect 6516 2237 6588 2243
rect 820 2217 876 2223
rect 884 2217 1004 2223
rect 1076 2217 1132 2223
rect 1140 2217 1244 2223
rect 1252 2217 1740 2223
rect 2173 2223 2179 2236
rect 1748 2217 2179 2223
rect 3012 2217 3084 2223
rect 3092 2217 3212 2223
rect 4228 2217 4284 2223
rect 4692 2217 5580 2223
rect 5588 2217 5708 2223
rect 6404 2217 6540 2223
rect 3304 2214 3352 2216
rect 3304 2206 3308 2214
rect 3318 2206 3324 2214
rect 3332 2206 3338 2214
rect 3348 2206 3352 2214
rect 3304 2204 3352 2206
rect 596 2197 652 2203
rect 1028 2197 1068 2203
rect 1076 2197 1468 2203
rect 1476 2197 1532 2203
rect 2388 2197 2572 2203
rect 2884 2197 2924 2203
rect 2932 2197 3084 2203
rect 4532 2197 5164 2203
rect 5172 2197 5340 2203
rect 5348 2197 5372 2203
rect 5972 2197 6012 2203
rect 6356 2197 6412 2203
rect 116 2177 188 2183
rect 372 2177 1443 2183
rect 68 2157 124 2163
rect 996 2157 1020 2163
rect 1437 2163 1443 2177
rect 1460 2177 1468 2183
rect 1476 2177 1548 2183
rect 1908 2177 2076 2183
rect 2772 2177 2812 2183
rect 2820 2177 2908 2183
rect 2932 2177 3036 2183
rect 3284 2177 3404 2183
rect 3412 2177 3452 2183
rect 4548 2177 4732 2183
rect 4740 2177 4796 2183
rect 5188 2177 5228 2183
rect 5620 2177 5836 2183
rect 6180 2177 6268 2183
rect 6276 2177 6332 2183
rect 6340 2177 6412 2183
rect 1437 2157 2700 2163
rect 2740 2157 2780 2163
rect 2788 2157 2860 2163
rect 2900 2157 2972 2163
rect 2980 2157 3020 2163
rect 3204 2157 3260 2163
rect 3412 2157 3420 2163
rect 3428 2157 3612 2163
rect 3652 2157 3868 2163
rect 3876 2157 4204 2163
rect 4212 2157 4444 2163
rect 4452 2157 4508 2163
rect 5156 2157 5212 2163
rect 5220 2157 5308 2163
rect 5428 2157 5500 2163
rect 5956 2157 6156 2163
rect 6164 2157 6492 2163
rect 148 2137 156 2143
rect 260 2137 332 2143
rect 580 2137 636 2143
rect 644 2137 700 2143
rect 980 2137 988 2143
rect 996 2137 1100 2143
rect 1108 2137 1132 2143
rect 1316 2137 1452 2143
rect 1748 2137 2092 2143
rect 2100 2137 2284 2143
rect 2468 2137 2604 2143
rect 2660 2137 2780 2143
rect 2820 2137 2988 2143
rect 3044 2137 3068 2143
rect 3076 2137 3132 2143
rect 3140 2137 3180 2143
rect 3284 2137 3308 2143
rect 3716 2137 3740 2143
rect 3780 2137 4028 2143
rect 4196 2137 4316 2143
rect 4516 2137 4604 2143
rect 4676 2137 4700 2143
rect 4820 2137 4924 2143
rect 4932 2137 5036 2143
rect 5044 2137 5148 2143
rect 5348 2137 5452 2143
rect 5604 2137 5660 2143
rect 6068 2137 6460 2143
rect 6516 2137 6524 2143
rect 52 2117 92 2123
rect 196 2117 220 2123
rect 292 2117 300 2123
rect 388 2117 476 2123
rect 532 2117 556 2123
rect 564 2117 604 2123
rect 756 2117 828 2123
rect 900 2117 924 2123
rect 1204 2117 1324 2123
rect 1636 2117 1820 2123
rect 1828 2117 1964 2123
rect 2036 2117 2156 2123
rect 2228 2117 2316 2123
rect 2372 2117 3084 2123
rect 3108 2117 3244 2123
rect 3252 2117 3340 2123
rect 3348 2117 3372 2123
rect 3556 2117 3660 2123
rect 4372 2117 4460 2123
rect 4596 2117 5084 2123
rect 5204 2117 5292 2123
rect 5300 2117 5388 2123
rect 5524 2117 5580 2123
rect 5604 2117 5628 2123
rect 6004 2117 6076 2123
rect 6084 2117 6204 2123
rect 6212 2117 6284 2123
rect 6292 2117 6332 2123
rect 6340 2117 6428 2123
rect 6468 2117 6524 2123
rect 36 2097 76 2103
rect 116 2097 204 2103
rect 340 2097 364 2103
rect 404 2097 460 2103
rect 468 2097 572 2103
rect 612 2097 652 2103
rect 660 2097 812 2103
rect 980 2097 1036 2103
rect 1044 2097 1180 2103
rect 1220 2097 1260 2103
rect 1300 2097 1356 2103
rect 1412 2097 1436 2103
rect 2324 2097 2380 2103
rect 3076 2097 3212 2103
rect 3220 2097 3404 2103
rect 3700 2097 3724 2103
rect 3732 2097 3836 2103
rect 3956 2097 4012 2103
rect 4036 2097 4076 2103
rect 4084 2097 4236 2103
rect 4452 2097 4508 2103
rect 5028 2097 5132 2103
rect 5140 2097 5260 2103
rect 5444 2097 5868 2103
rect 5924 2097 6172 2103
rect 6180 2097 6236 2103
rect 6244 2097 6300 2103
rect 6324 2097 6380 2103
rect 6388 2097 6396 2103
rect 6452 2097 6556 2103
rect 52 2077 140 2083
rect 244 2077 268 2083
rect 308 2077 348 2083
rect 500 2077 588 2083
rect 692 2077 716 2083
rect 724 2077 1196 2083
rect 1348 2077 1420 2083
rect 4500 2077 4828 2083
rect 4836 2077 4940 2083
rect 5060 2077 5372 2083
rect 5380 2077 5548 2083
rect 5972 2077 6444 2083
rect 6548 2077 6572 2083
rect 1172 2057 1276 2063
rect 4404 2057 5068 2063
rect 5076 2057 5100 2063
rect 6212 2057 6364 2063
rect 2660 2037 4124 2043
rect 4708 2037 4956 2043
rect 5044 2037 5068 2043
rect 5092 2037 5532 2043
rect 1028 2017 1148 2023
rect 5076 2017 5388 2023
rect 5396 2017 5516 2023
rect 1768 2014 1816 2016
rect 1768 2006 1772 2014
rect 1782 2006 1788 2014
rect 1796 2006 1802 2014
rect 1812 2006 1816 2014
rect 1768 2004 1816 2006
rect 4824 2014 4872 2016
rect 4824 2006 4828 2014
rect 4838 2006 4844 2014
rect 4852 2006 4858 2014
rect 4868 2006 4872 2014
rect 4824 2004 4872 2006
rect 100 1997 156 2003
rect 452 1997 524 2003
rect 532 1997 668 2003
rect 676 1997 716 2003
rect 1524 1997 1580 2003
rect 2180 1997 3980 2003
rect 5524 1997 6076 2003
rect 6196 1997 6508 2003
rect 660 1977 668 1983
rect 2372 1977 2380 1983
rect 2452 1977 2876 1983
rect 3124 1977 3148 1983
rect 4260 1977 4396 1983
rect 4484 1977 5308 1983
rect 5316 1977 5468 1983
rect 5508 1977 6028 1983
rect 6532 1977 6556 1983
rect 116 1957 124 1963
rect 884 1957 956 1963
rect 1188 1957 1676 1963
rect 1700 1957 1788 1963
rect 2052 1957 2796 1963
rect 2916 1957 3052 1963
rect 4900 1957 4988 1963
rect 5364 1957 5388 1963
rect 5748 1957 5932 1963
rect 6548 1957 6572 1963
rect 20 1937 204 1943
rect 340 1937 364 1943
rect 1188 1937 1388 1943
rect 1636 1937 1692 1943
rect 1700 1937 2220 1943
rect 2580 1937 2924 1943
rect 2932 1937 3196 1943
rect 3268 1937 3660 1943
rect 3668 1937 3708 1943
rect 3892 1937 4339 1943
rect 4333 1924 4339 1937
rect 4644 1937 4940 1943
rect 4948 1937 5020 1943
rect 5220 1937 5452 1943
rect 5524 1937 5660 1943
rect 5716 1937 5756 1943
rect 5956 1937 5980 1943
rect 6436 1937 6540 1943
rect 6548 1937 6588 1943
rect 52 1917 92 1923
rect 180 1917 236 1923
rect 340 1917 492 1923
rect 708 1917 780 1923
rect 788 1917 812 1923
rect 836 1917 956 1923
rect 1012 1917 1068 1923
rect 1076 1917 1116 1923
rect 1124 1917 1196 1923
rect 1300 1917 1388 1923
rect 1396 1917 1404 1923
rect 1412 1917 1420 1923
rect 1540 1917 1724 1923
rect 1844 1917 1884 1923
rect 1892 1917 1996 1923
rect 2356 1917 2364 1923
rect 2564 1917 2771 1923
rect 2765 1904 2771 1917
rect 2996 1917 3436 1923
rect 3444 1917 3692 1923
rect 3700 1917 3964 1923
rect 4340 1917 4508 1923
rect 4516 1917 4572 1923
rect 4660 1917 4684 1923
rect 4724 1917 4764 1923
rect 4804 1917 4892 1923
rect 4900 1917 4956 1923
rect 5188 1917 5404 1923
rect 5556 1917 5612 1923
rect 5700 1917 5740 1923
rect 5748 1917 5788 1923
rect 5812 1917 5868 1923
rect 5940 1917 6252 1923
rect 6260 1917 6300 1923
rect 6340 1917 6412 1923
rect 6468 1917 6508 1923
rect 6532 1917 6588 1923
rect 36 1897 108 1903
rect 164 1897 220 1903
rect 308 1897 348 1903
rect 356 1897 396 1903
rect 436 1897 492 1903
rect 548 1897 588 1903
rect 644 1897 668 1903
rect 884 1897 988 1903
rect 1060 1897 1116 1903
rect 1124 1897 1452 1903
rect 1524 1897 1660 1903
rect 2116 1897 2156 1903
rect 2260 1897 2636 1903
rect 2772 1897 2940 1903
rect 2964 1897 3004 1903
rect 3060 1897 3116 1903
rect 3236 1897 3260 1903
rect 3428 1897 3548 1903
rect 3860 1897 3980 1903
rect 4212 1897 4268 1903
rect 4884 1897 4924 1903
rect 4932 1897 5020 1903
rect 5028 1897 5164 1903
rect 5300 1897 5340 1903
rect 5412 1897 5852 1903
rect 5860 1897 5932 1903
rect 5972 1897 5996 1903
rect 6356 1897 6428 1903
rect 6436 1897 6460 1903
rect 6484 1897 6540 1903
rect 372 1877 428 1883
rect 500 1877 556 1883
rect 564 1877 700 1883
rect 868 1877 908 1883
rect 916 1877 940 1883
rect 1140 1877 1180 1883
rect 1204 1877 1452 1883
rect 1460 1877 1500 1883
rect 1588 1877 1804 1883
rect 1812 1877 1836 1883
rect 1844 1877 1900 1883
rect 2820 1877 2924 1883
rect 3044 1877 3212 1883
rect 3220 1877 3324 1883
rect 3348 1877 3644 1883
rect 3652 1877 3724 1883
rect 3764 1877 4156 1883
rect 4676 1877 4940 1883
rect 4948 1877 4988 1883
rect 5012 1877 5036 1883
rect 5044 1877 5452 1883
rect 5652 1877 5731 1883
rect 276 1857 444 1863
rect 516 1857 732 1863
rect 756 1857 844 1863
rect 852 1857 892 1863
rect 916 1857 1084 1863
rect 1252 1857 1564 1863
rect 1572 1857 1740 1863
rect 2004 1857 2060 1863
rect 2708 1857 2956 1863
rect 3108 1857 3228 1863
rect 3700 1857 4172 1863
rect 4516 1857 4684 1863
rect 4692 1857 4908 1863
rect 4916 1857 4972 1863
rect 5012 1857 5084 1863
rect 5092 1857 5116 1863
rect 5204 1857 5292 1863
rect 5300 1857 5388 1863
rect 5428 1857 5436 1863
rect 5572 1857 5676 1863
rect 5684 1857 5708 1863
rect 5725 1863 5731 1877
rect 5748 1877 6012 1883
rect 6164 1877 6220 1883
rect 5725 1857 5900 1863
rect 5940 1857 6076 1863
rect 804 1837 828 1843
rect 836 1837 1132 1843
rect 2788 1837 3148 1843
rect 3156 1837 3196 1843
rect 3204 1837 3244 1843
rect 3284 1837 3404 1843
rect 3412 1837 3452 1843
rect 3956 1837 4028 1843
rect 4132 1837 4220 1843
rect 4228 1837 4748 1843
rect 4973 1843 4979 1856
rect 4973 1837 5228 1843
rect 5268 1837 5308 1843
rect 5620 1837 5820 1843
rect 5828 1837 5884 1843
rect 6068 1837 6268 1843
rect 852 1817 1260 1823
rect 1300 1817 1516 1823
rect 2884 1817 2908 1823
rect 3956 1817 4076 1823
rect 4244 1817 4524 1823
rect 4644 1817 5676 1823
rect 5716 1817 5772 1823
rect 5988 1817 6108 1823
rect 6116 1817 6348 1823
rect 6356 1817 6380 1823
rect 6484 1817 6508 1823
rect 3304 1814 3352 1816
rect 3304 1806 3308 1814
rect 3318 1806 3324 1814
rect 3332 1806 3338 1814
rect 3348 1806 3352 1814
rect 3304 1804 3352 1806
rect 260 1797 300 1803
rect 356 1797 812 1803
rect 916 1797 1004 1803
rect 1012 1797 1356 1803
rect 1428 1797 1548 1803
rect 1556 1797 1852 1803
rect 2084 1797 2220 1803
rect 4164 1797 4204 1803
rect 4212 1797 4332 1803
rect 4340 1797 4604 1803
rect 4740 1797 4892 1803
rect 5140 1797 5804 1803
rect 5844 1797 6092 1803
rect 6100 1797 6364 1803
rect 724 1777 780 1783
rect 948 1777 1596 1783
rect 1620 1777 1692 1783
rect 1860 1777 1964 1783
rect 1988 1777 2044 1783
rect 2692 1777 2796 1783
rect 2804 1777 2972 1783
rect 3556 1777 3740 1783
rect 3748 1777 4524 1783
rect 4733 1783 4739 1796
rect 4612 1777 4739 1783
rect 5156 1777 5196 1783
rect 5204 1777 5260 1783
rect 5476 1777 5564 1783
rect 5732 1777 5980 1783
rect 6356 1777 6380 1783
rect 20 1757 44 1763
rect 116 1757 380 1763
rect 436 1757 508 1763
rect 772 1757 844 1763
rect 852 1757 1020 1763
rect 1156 1757 1212 1763
rect 1220 1757 1292 1763
rect 1332 1757 1468 1763
rect 1476 1757 1516 1763
rect 1524 1757 1628 1763
rect 3060 1757 3164 1763
rect 3188 1757 3436 1763
rect 3444 1757 3516 1763
rect 3924 1757 4492 1763
rect 4692 1757 4812 1763
rect 5124 1757 5212 1763
rect 5300 1757 5356 1763
rect 5364 1757 5404 1763
rect 5732 1757 5756 1763
rect 5780 1757 5900 1763
rect 5924 1757 6012 1763
rect 6052 1757 6108 1763
rect 6116 1757 6140 1763
rect 6308 1757 6364 1763
rect 132 1737 188 1743
rect 564 1737 764 1743
rect 788 1737 972 1743
rect 996 1737 1036 1743
rect 1044 1737 1052 1743
rect 1092 1737 1500 1743
rect 1604 1737 1644 1743
rect 2820 1737 2876 1743
rect 3076 1737 3100 1743
rect 3108 1737 3292 1743
rect 3300 1737 3356 1743
rect 3908 1737 4012 1743
rect 4020 1737 4236 1743
rect 4452 1737 4476 1743
rect 4676 1737 4780 1743
rect 5044 1737 5276 1743
rect 5316 1737 5404 1743
rect 5668 1737 5804 1743
rect 5812 1737 5836 1743
rect 5844 1737 5932 1743
rect 6141 1737 6220 1743
rect 6141 1724 6147 1737
rect 6276 1737 6284 1743
rect 6436 1737 6460 1743
rect 6500 1737 6508 1743
rect 6516 1737 6524 1743
rect 404 1717 492 1723
rect 532 1717 620 1723
rect 708 1717 780 1723
rect 788 1717 1308 1723
rect 1620 1717 1820 1723
rect 2164 1717 2252 1723
rect 2260 1717 2444 1723
rect 2516 1717 2604 1723
rect 2676 1717 2940 1723
rect 2948 1717 2988 1723
rect 2996 1717 3180 1723
rect 3364 1717 3452 1723
rect 3492 1717 3612 1723
rect 3684 1717 3756 1723
rect 4004 1717 4108 1723
rect 4116 1717 4332 1723
rect 4628 1717 4652 1723
rect 4724 1717 4796 1723
rect 4804 1717 4828 1723
rect 5252 1717 5500 1723
rect 5508 1717 5692 1723
rect 5700 1717 5740 1723
rect 5748 1717 5788 1723
rect 5812 1717 5852 1723
rect 6020 1717 6140 1723
rect 6196 1717 6252 1723
rect 6260 1717 6396 1723
rect 6452 1717 6524 1723
rect 180 1697 220 1703
rect 228 1697 268 1703
rect 324 1697 348 1703
rect 516 1697 572 1703
rect 644 1697 684 1703
rect 692 1697 716 1703
rect 900 1697 972 1703
rect 1012 1697 1212 1703
rect 1220 1697 1244 1703
rect 2669 1703 2675 1716
rect 2612 1697 2675 1703
rect 2884 1697 2956 1703
rect 3236 1697 3388 1703
rect 3556 1697 4460 1703
rect 4548 1697 4700 1703
rect 5092 1697 5212 1703
rect 5220 1697 5228 1703
rect 5316 1697 5420 1703
rect 5892 1697 6028 1703
rect 6036 1697 6156 1703
rect 6180 1697 6236 1703
rect 6244 1697 6284 1703
rect 6452 1697 6476 1703
rect 52 1677 92 1683
rect 100 1677 188 1683
rect 388 1677 444 1683
rect 452 1677 476 1683
rect 484 1677 540 1683
rect 548 1677 716 1683
rect 740 1677 780 1683
rect 1124 1677 1164 1683
rect 1172 1677 1260 1683
rect 1268 1677 1436 1683
rect 1444 1677 1564 1683
rect 2372 1677 3884 1683
rect 3892 1677 4684 1683
rect 4788 1677 5036 1683
rect 5076 1677 5132 1683
rect 5396 1677 5676 1683
rect 5684 1677 5772 1683
rect 5780 1677 5820 1683
rect 6068 1677 6108 1683
rect 6132 1677 6156 1683
rect 6180 1677 6316 1683
rect 6356 1677 6412 1683
rect 6420 1677 6508 1683
rect 516 1657 604 1663
rect 733 1663 739 1676
rect 612 1657 739 1663
rect 964 1657 1084 1663
rect 1140 1657 1276 1663
rect 1284 1657 1404 1663
rect 1492 1657 1788 1663
rect 2388 1657 2572 1663
rect 2852 1657 3116 1663
rect 3300 1657 4636 1663
rect 4756 1657 5516 1663
rect 5588 1657 6028 1663
rect 228 1637 252 1643
rect 260 1637 284 1643
rect 644 1637 812 1643
rect 1332 1637 1852 1643
rect 4532 1637 4764 1643
rect 5108 1637 5484 1643
rect 5908 1637 5964 1643
rect 6068 1637 6236 1643
rect 6468 1637 6476 1643
rect 6548 1637 6588 1643
rect 1028 1617 1324 1623
rect 1380 1617 1436 1623
rect 4564 1617 4604 1623
rect 4612 1617 4716 1623
rect 5092 1617 5340 1623
rect 5972 1617 6044 1623
rect 6244 1617 6268 1623
rect 1768 1614 1816 1616
rect 1768 1606 1772 1614
rect 1782 1606 1788 1614
rect 1796 1606 1802 1614
rect 1812 1606 1816 1614
rect 1768 1604 1816 1606
rect 4824 1614 4872 1616
rect 4824 1606 4828 1614
rect 4838 1606 4844 1614
rect 4852 1606 4858 1614
rect 4868 1606 4872 1614
rect 4824 1604 4872 1606
rect 756 1597 876 1603
rect 1284 1597 1308 1603
rect 1508 1597 1628 1603
rect 1716 1597 1740 1603
rect 2900 1597 3532 1603
rect 4516 1597 4524 1603
rect 4548 1597 4803 1603
rect 804 1577 940 1583
rect 1028 1577 1084 1583
rect 1572 1577 1948 1583
rect 3780 1577 3900 1583
rect 3908 1577 4044 1583
rect 4068 1577 4460 1583
rect 4500 1577 4668 1583
rect 4676 1577 4716 1583
rect 4797 1583 4803 1597
rect 4932 1597 5372 1603
rect 5636 1597 5676 1603
rect 5908 1597 5996 1603
rect 6276 1597 6476 1603
rect 6484 1597 6540 1603
rect 4797 1577 4860 1583
rect 4884 1577 4940 1583
rect 4980 1577 5260 1583
rect 5284 1577 6028 1583
rect 6036 1577 6220 1583
rect 6420 1577 6588 1583
rect 212 1557 252 1563
rect 884 1557 956 1563
rect 1044 1557 1148 1563
rect 1220 1557 1372 1563
rect 1524 1557 1676 1563
rect 2228 1557 2380 1563
rect 2452 1557 2636 1563
rect 3124 1557 3580 1563
rect 3956 1557 4220 1563
rect 4468 1557 4700 1563
rect 4852 1557 4940 1563
rect 4948 1557 5020 1563
rect 5028 1557 5276 1563
rect 5284 1557 5532 1563
rect 5636 1557 5964 1563
rect 5972 1557 6076 1563
rect 6100 1557 6172 1563
rect 6292 1557 6396 1563
rect 100 1537 156 1543
rect 164 1537 300 1543
rect 452 1537 844 1543
rect 948 1537 972 1543
rect 1092 1537 1164 1543
rect 1172 1537 1420 1543
rect 1444 1537 1612 1543
rect 1668 1537 1740 1543
rect 2068 1537 2124 1543
rect 2132 1537 2172 1543
rect 2180 1537 2211 1543
rect 68 1517 76 1523
rect 84 1517 172 1523
rect 180 1517 284 1523
rect 292 1517 332 1523
rect 484 1517 508 1523
rect 532 1517 684 1523
rect 868 1517 972 1523
rect 980 1517 1100 1523
rect 1108 1517 1484 1523
rect 1524 1517 1596 1523
rect 1604 1517 1676 1523
rect 1684 1517 1868 1523
rect 1940 1517 2012 1523
rect 2205 1523 2211 1537
rect 2596 1537 2780 1543
rect 2788 1537 2876 1543
rect 2884 1537 3404 1543
rect 3684 1537 3724 1543
rect 3732 1537 3932 1543
rect 4036 1537 4156 1543
rect 4164 1537 4188 1543
rect 4404 1537 4460 1543
rect 4468 1537 5068 1543
rect 5076 1537 5164 1543
rect 5172 1537 5228 1543
rect 5412 1537 5644 1543
rect 5725 1537 5980 1543
rect 2100 1517 2195 1523
rect 2205 1517 2620 1523
rect 2189 1504 2195 1517
rect 2644 1517 2908 1523
rect 3412 1517 3436 1523
rect 3924 1517 3948 1523
rect 3956 1517 4044 1523
rect 4084 1517 4140 1523
rect 4276 1517 4412 1523
rect 4420 1517 4508 1523
rect 4516 1517 4572 1523
rect 4804 1517 4924 1523
rect 4932 1517 4972 1523
rect 5044 1517 5100 1523
rect 5156 1517 5244 1523
rect 5268 1517 5292 1523
rect 5725 1523 5731 1537
rect 6052 1537 6332 1543
rect 6356 1537 6476 1543
rect 6484 1537 6492 1543
rect 5460 1517 5731 1523
rect 5748 1517 5795 1523
rect 52 1497 140 1503
rect 196 1497 268 1503
rect 436 1497 588 1503
rect 612 1497 620 1503
rect 692 1497 716 1503
rect 836 1497 1139 1503
rect 1133 1484 1139 1497
rect 1204 1497 1228 1503
rect 1332 1497 1388 1503
rect 1396 1497 1532 1503
rect 1764 1497 1964 1503
rect 1988 1497 2131 1503
rect 116 1477 140 1483
rect 164 1477 332 1483
rect 564 1477 620 1483
rect 724 1477 780 1483
rect 820 1477 844 1483
rect 868 1477 892 1483
rect 932 1477 1036 1483
rect 1252 1477 1276 1483
rect 1428 1477 1500 1483
rect 2020 1477 2108 1483
rect 2125 1483 2131 1497
rect 2196 1497 2412 1503
rect 2532 1497 2556 1503
rect 2692 1497 2892 1503
rect 2948 1497 3164 1503
rect 3172 1497 3260 1503
rect 3444 1497 3500 1503
rect 3652 1497 3692 1503
rect 3700 1497 3740 1503
rect 4116 1497 4140 1503
rect 4148 1497 4172 1503
rect 4340 1497 4396 1503
rect 4404 1497 4492 1503
rect 4532 1497 4588 1503
rect 4660 1497 4780 1503
rect 4788 1497 4851 1503
rect 2125 1477 2220 1483
rect 2356 1477 2380 1483
rect 2388 1477 2476 1483
rect 2516 1477 2540 1483
rect 2548 1477 2572 1483
rect 2580 1477 2700 1483
rect 2756 1477 2972 1483
rect 2996 1477 3244 1483
rect 3252 1477 3452 1483
rect 3492 1477 3596 1483
rect 3604 1477 3660 1483
rect 3684 1477 3804 1483
rect 3860 1477 4140 1483
rect 4189 1477 4252 1483
rect 36 1457 124 1463
rect 132 1457 316 1463
rect 356 1457 396 1463
rect 621 1463 627 1476
rect 621 1457 668 1463
rect 772 1457 892 1463
rect 1197 1463 1203 1476
rect 1076 1457 1436 1463
rect 1700 1457 1820 1463
rect 2260 1457 2556 1463
rect 2564 1457 2588 1463
rect 2628 1457 2796 1463
rect 2804 1457 2908 1463
rect 2916 1457 3420 1463
rect 3844 1457 3916 1463
rect 4189 1463 4195 1477
rect 4372 1477 4396 1483
rect 4564 1477 4796 1483
rect 4845 1483 4851 1497
rect 4868 1497 5084 1503
rect 5092 1497 5132 1503
rect 5341 1497 5628 1503
rect 4845 1477 4908 1483
rect 4916 1477 4956 1483
rect 4116 1457 4195 1463
rect 4212 1457 4332 1463
rect 4356 1457 4380 1463
rect 4388 1457 4636 1463
rect 4644 1457 4924 1463
rect 5181 1463 5187 1496
rect 5341 1483 5347 1497
rect 5652 1497 5756 1503
rect 5789 1503 5795 1517
rect 5812 1517 6099 1523
rect 5789 1497 5932 1503
rect 5940 1497 6012 1503
rect 6093 1503 6099 1517
rect 6116 1517 6140 1523
rect 6212 1517 6252 1523
rect 6292 1517 6364 1523
rect 6404 1517 6444 1523
rect 6452 1517 6524 1523
rect 6093 1497 6124 1503
rect 6132 1497 6172 1503
rect 6276 1497 6332 1503
rect 6404 1497 6444 1503
rect 5268 1477 5347 1483
rect 5364 1477 5564 1483
rect 5636 1477 5660 1483
rect 5684 1477 5788 1483
rect 5796 1477 5836 1483
rect 5844 1477 5900 1483
rect 5988 1477 6076 1483
rect 6132 1477 6380 1483
rect 6388 1477 6428 1483
rect 6436 1477 6508 1483
rect 5156 1457 5187 1463
rect 5492 1457 5596 1463
rect 5604 1457 5820 1463
rect 5844 1457 5916 1463
rect 5924 1457 5996 1463
rect 6164 1457 6204 1463
rect 6340 1457 6364 1463
rect 6372 1457 6572 1463
rect 596 1437 604 1443
rect 765 1443 771 1456
rect 612 1437 771 1443
rect 916 1437 1356 1443
rect 1380 1437 1580 1443
rect 1700 1437 1740 1443
rect 1908 1437 2140 1443
rect 2148 1437 2316 1443
rect 2452 1437 2812 1443
rect 2820 1437 2956 1443
rect 2964 1437 3276 1443
rect 3972 1437 4156 1443
rect 4180 1437 4556 1443
rect 4772 1437 5436 1443
rect 5444 1437 5548 1443
rect 5556 1437 5644 1443
rect 5668 1437 5772 1443
rect 5796 1437 5804 1443
rect 5844 1437 5868 1443
rect 5892 1437 6108 1443
rect 628 1417 1212 1423
rect 1284 1417 1292 1423
rect 1332 1417 1564 1423
rect 1588 1417 1660 1423
rect 1684 1417 1948 1423
rect 2404 1417 2668 1423
rect 2708 1417 2940 1423
rect 2980 1417 3180 1423
rect 3188 1417 3212 1423
rect 3652 1417 3868 1423
rect 3876 1417 4300 1423
rect 4308 1417 4716 1423
rect 4996 1417 5884 1423
rect 5892 1417 6060 1423
rect 6068 1417 6156 1423
rect 6164 1417 6220 1423
rect 3304 1414 3352 1416
rect 3304 1406 3308 1414
rect 3318 1406 3324 1414
rect 3332 1406 3338 1414
rect 3348 1406 3352 1414
rect 3304 1404 3352 1406
rect 772 1397 1292 1403
rect 1940 1397 1996 1403
rect 2004 1397 2156 1403
rect 2436 1397 2924 1403
rect 2932 1397 3228 1403
rect 3396 1397 3516 1403
rect 3524 1397 3740 1403
rect 3908 1397 4012 1403
rect 4116 1397 4252 1403
rect 4324 1397 4540 1403
rect 4596 1397 4988 1403
rect 5140 1397 5260 1403
rect 5284 1397 5340 1403
rect 5476 1397 5612 1403
rect 5620 1397 5868 1403
rect 5940 1397 5996 1403
rect 6004 1397 6124 1403
rect 6132 1397 6268 1403
rect 580 1377 588 1383
rect 804 1377 1036 1383
rect 1076 1377 1132 1383
rect 1220 1377 1708 1383
rect 2164 1377 2252 1383
rect 2260 1377 2348 1383
rect 2356 1377 2764 1383
rect 2804 1377 2828 1383
rect 2884 1377 2972 1383
rect 2996 1377 3020 1383
rect 3076 1377 3116 1383
rect 3124 1377 3196 1383
rect 3204 1377 3244 1383
rect 3268 1377 3292 1383
rect 3300 1377 3404 1383
rect 3501 1377 3644 1383
rect 3501 1364 3507 1377
rect 3732 1377 4060 1383
rect 4100 1377 4412 1383
rect 4420 1377 4476 1383
rect 4676 1377 4780 1383
rect 4820 1377 5452 1383
rect 5508 1377 5852 1383
rect 5860 1377 5868 1383
rect 5956 1377 5980 1383
rect 6036 1377 6188 1383
rect 68 1357 124 1363
rect 132 1357 204 1363
rect 212 1357 332 1363
rect 548 1357 572 1363
rect 580 1357 780 1363
rect 1012 1357 1052 1363
rect 1069 1357 1251 1363
rect 52 1337 140 1343
rect 244 1337 444 1343
rect 676 1337 780 1343
rect 1069 1343 1075 1357
rect 1245 1344 1251 1357
rect 1300 1357 1388 1363
rect 1428 1357 1475 1363
rect 1469 1344 1475 1357
rect 1668 1357 1916 1363
rect 2212 1357 2300 1363
rect 2372 1357 2428 1363
rect 2580 1357 2668 1363
rect 2676 1357 2780 1363
rect 2836 1357 3308 1363
rect 3396 1357 3452 1363
rect 3476 1357 3500 1363
rect 3556 1357 3628 1363
rect 3636 1357 3756 1363
rect 3972 1357 4028 1363
rect 4100 1357 4140 1363
rect 4196 1357 4220 1363
rect 4228 1357 4284 1363
rect 4692 1357 4940 1363
rect 4964 1357 5020 1363
rect 5172 1357 5212 1363
rect 5348 1357 5516 1363
rect 5588 1357 5772 1363
rect 5812 1357 5948 1363
rect 6052 1357 6108 1363
rect 6164 1357 6172 1363
rect 6340 1357 6524 1363
rect 948 1337 1075 1343
rect 1156 1337 1196 1343
rect 1252 1337 1452 1343
rect 1476 1337 1548 1343
rect 1572 1337 1676 1343
rect 1716 1337 1772 1343
rect 1876 1337 2012 1343
rect 2308 1337 2332 1343
rect 2340 1337 2364 1343
rect 2372 1337 2492 1343
rect 2596 1337 2620 1343
rect 2740 1337 2780 1343
rect 2900 1337 2988 1343
rect 3469 1337 3580 1343
rect 3469 1324 3475 1337
rect 3588 1337 3660 1343
rect 3716 1337 3788 1343
rect 3796 1337 3820 1343
rect 3844 1337 4035 1343
rect 52 1317 92 1323
rect 260 1317 332 1323
rect 340 1317 380 1323
rect 484 1317 524 1323
rect 532 1317 684 1323
rect 1028 1317 1052 1323
rect 1092 1317 1116 1323
rect 1140 1317 1340 1323
rect 1348 1317 1516 1323
rect 1860 1317 1932 1323
rect 2068 1317 2108 1323
rect 2116 1317 2220 1323
rect 2228 1317 2316 1323
rect 2324 1317 2540 1323
rect 2628 1317 2748 1323
rect 2948 1317 3132 1323
rect 3140 1317 3276 1323
rect 3412 1317 3468 1323
rect 3556 1317 3564 1323
rect 3620 1317 3708 1323
rect 3764 1317 3820 1323
rect 3860 1317 3884 1323
rect 3940 1317 4012 1323
rect 4029 1323 4035 1337
rect 4052 1337 4124 1343
rect 4164 1337 4188 1343
rect 4244 1337 4268 1343
rect 4468 1337 4620 1343
rect 4708 1337 4860 1343
rect 4868 1337 5036 1343
rect 5076 1337 5116 1343
rect 5220 1337 5324 1343
rect 5412 1337 5548 1343
rect 5572 1337 5660 1343
rect 5764 1337 5820 1343
rect 5860 1337 5868 1343
rect 5956 1337 6172 1343
rect 6420 1337 6556 1343
rect 4029 1317 4428 1323
rect 4436 1317 4492 1323
rect 4564 1317 4604 1323
rect 4676 1317 4876 1323
rect 4948 1317 5196 1323
rect 5316 1317 5324 1323
rect 5444 1317 5484 1323
rect 5588 1317 5676 1323
rect 5812 1317 5868 1323
rect 5972 1317 6012 1323
rect 6020 1317 6076 1323
rect 6276 1317 6348 1323
rect 6356 1317 6428 1323
rect 52 1297 188 1303
rect 356 1297 412 1303
rect 564 1297 588 1303
rect 596 1297 652 1303
rect 692 1297 908 1303
rect 996 1297 1324 1303
rect 1556 1297 1580 1303
rect 1732 1297 1868 1303
rect 1876 1297 1932 1303
rect 2132 1297 2172 1303
rect 2180 1297 2268 1303
rect 2276 1297 2380 1303
rect 2388 1297 2524 1303
rect 2964 1297 3052 1303
rect 3236 1297 3452 1303
rect 3460 1297 3484 1303
rect 3492 1297 3564 1303
rect 3572 1297 6124 1303
rect 6164 1297 6380 1303
rect 6452 1297 6508 1303
rect 36 1277 76 1283
rect 276 1277 316 1283
rect 324 1277 364 1283
rect 452 1277 508 1283
rect 516 1277 604 1283
rect 1028 1277 1084 1283
rect 1220 1277 1292 1283
rect 1396 1277 1452 1283
rect 1476 1277 1532 1283
rect 1540 1277 1628 1283
rect 1828 1277 2284 1283
rect 2772 1277 2844 1283
rect 3156 1277 3196 1283
rect 3492 1277 3612 1283
rect 3668 1277 3996 1283
rect 4260 1277 4556 1283
rect 4564 1277 4636 1283
rect 4852 1277 5036 1283
rect 5044 1277 5132 1283
rect 5140 1277 5180 1283
rect 5380 1277 5500 1283
rect 5508 1277 5532 1283
rect 5556 1277 5884 1283
rect 5892 1277 6188 1283
rect 6292 1277 6348 1283
rect 6372 1277 6412 1283
rect 292 1257 348 1263
rect 868 1257 1308 1263
rect 3028 1257 3228 1263
rect 3700 1257 3772 1263
rect 3892 1257 3980 1263
rect 4756 1257 4972 1263
rect 5428 1257 5580 1263
rect 6132 1257 6140 1263
rect 964 1237 1219 1243
rect 1213 1224 1219 1237
rect 1588 1237 1676 1243
rect 4372 1237 5132 1243
rect 5940 1237 6204 1243
rect 6324 1237 6332 1243
rect 1220 1217 1372 1223
rect 5076 1217 5724 1223
rect 6084 1217 6124 1223
rect 6132 1217 6172 1223
rect 6244 1217 6284 1223
rect 6324 1217 6460 1223
rect 1768 1214 1816 1216
rect 1768 1206 1772 1214
rect 1782 1206 1788 1214
rect 1796 1206 1802 1214
rect 1812 1206 1816 1214
rect 1768 1204 1816 1206
rect 4824 1214 4872 1216
rect 4824 1206 4828 1214
rect 4838 1206 4844 1214
rect 4852 1206 4858 1214
rect 4868 1206 4872 1214
rect 4824 1204 4872 1206
rect 740 1197 1004 1203
rect 1140 1197 1516 1203
rect 2404 1197 2476 1203
rect 3252 1197 4364 1203
rect 5524 1197 5708 1203
rect 6004 1197 6572 1203
rect 52 1177 76 1183
rect 84 1177 284 1183
rect 628 1177 812 1183
rect 1092 1177 1228 1183
rect 3220 1177 3484 1183
rect 3492 1177 3548 1183
rect 3556 1177 3628 1183
rect 4964 1177 5260 1183
rect 5316 1177 5420 1183
rect 5924 1177 6156 1183
rect 6260 1177 6428 1183
rect 6468 1177 6556 1183
rect 244 1157 268 1163
rect 404 1157 428 1163
rect 836 1157 972 1163
rect 1012 1157 1116 1163
rect 1124 1157 1148 1163
rect 2068 1157 2268 1163
rect 2852 1157 2956 1163
rect 2964 1157 3468 1163
rect 4612 1157 5260 1163
rect 5300 1157 5356 1163
rect 5428 1157 6044 1163
rect 6052 1157 6076 1163
rect 6260 1157 6348 1163
rect 6404 1157 6572 1163
rect 36 1137 44 1143
rect 180 1137 236 1143
rect 308 1137 364 1143
rect 436 1137 636 1143
rect 756 1137 892 1143
rect 1076 1137 1116 1143
rect 1124 1137 1164 1143
rect 1252 1137 1292 1143
rect 1428 1137 1564 1143
rect 1892 1137 1916 1143
rect 2148 1137 2188 1143
rect 2212 1137 2220 1143
rect 2228 1137 2300 1143
rect 2484 1137 2508 1143
rect 2580 1137 2700 1143
rect 2980 1137 3020 1143
rect 3284 1137 3580 1143
rect 4036 1137 4092 1143
rect 4100 1137 4348 1143
rect 4436 1137 4492 1143
rect 4532 1137 4636 1143
rect 4644 1137 4716 1143
rect 4980 1137 5436 1143
rect 5492 1137 5532 1143
rect 5540 1137 5628 1143
rect 6116 1137 6204 1143
rect 6292 1137 6364 1143
rect 6388 1137 6444 1143
rect 6452 1137 6508 1143
rect 6564 1137 6636 1143
rect 36 1117 108 1123
rect 292 1117 332 1123
rect 548 1117 668 1123
rect 772 1117 860 1123
rect 884 1117 908 1123
rect 916 1117 988 1123
rect 996 1117 1276 1123
rect 1284 1117 1356 1123
rect 1492 1117 1548 1123
rect 2100 1117 2124 1123
rect 2180 1117 2556 1123
rect 2884 1117 2924 1123
rect 2932 1117 2956 1123
rect 3021 1117 3052 1123
rect 84 1097 140 1103
rect 164 1097 220 1103
rect 356 1097 412 1103
rect 484 1097 588 1103
rect 724 1097 796 1103
rect 820 1097 876 1103
rect 884 1097 1020 1103
rect 1028 1097 1372 1103
rect 1380 1097 1388 1103
rect 1476 1097 1484 1103
rect 1492 1097 1580 1103
rect 1700 1097 1708 1103
rect 1828 1097 1884 1103
rect 2036 1097 2092 1103
rect 2132 1097 2188 1103
rect 2196 1097 2236 1103
rect 2244 1097 2460 1103
rect 2516 1097 2652 1103
rect 3021 1103 3027 1117
rect 3092 1117 3436 1123
rect 3620 1117 3692 1123
rect 3780 1117 3980 1123
rect 4020 1117 4124 1123
rect 4212 1117 4252 1123
rect 4484 1117 4588 1123
rect 5012 1117 5084 1123
rect 5252 1117 5500 1123
rect 5908 1117 5980 1123
rect 6068 1117 6284 1123
rect 6292 1117 6332 1123
rect 6340 1117 6396 1123
rect 6532 1117 6636 1123
rect 2932 1097 3027 1103
rect 3044 1097 3116 1103
rect 3188 1097 3244 1103
rect 3348 1097 3372 1103
rect 3732 1097 3788 1103
rect 4004 1097 4204 1103
rect 4484 1097 4524 1103
rect 4532 1097 4556 1103
rect 4660 1097 4700 1103
rect 4916 1097 4988 1103
rect 4996 1097 5228 1103
rect 5252 1097 5324 1103
rect 5348 1097 5660 1103
rect 5668 1097 5724 1103
rect 5732 1097 5740 1103
rect 5828 1097 5884 1103
rect 5940 1097 5980 1103
rect 5988 1097 6028 1103
rect 6068 1097 6140 1103
rect 6164 1097 6188 1103
rect 6292 1097 6348 1103
rect 6388 1097 6412 1103
rect 6452 1097 6492 1103
rect 6516 1097 6540 1103
rect 52 1077 76 1083
rect 84 1077 92 1083
rect 132 1077 172 1083
rect 260 1077 268 1083
rect 468 1077 492 1083
rect 500 1077 556 1083
rect 804 1077 924 1083
rect 932 1077 1292 1083
rect 1300 1077 1308 1083
rect 1380 1077 1436 1083
rect 1636 1077 1692 1083
rect 2820 1077 2876 1083
rect 2884 1077 2940 1083
rect 3012 1077 3084 1083
rect 3156 1077 3196 1083
rect 3341 1083 3347 1096
rect 3236 1077 3347 1083
rect 3556 1077 3644 1083
rect 3748 1077 3836 1083
rect 3924 1077 3932 1083
rect 4132 1077 4236 1083
rect 4404 1077 4828 1083
rect 5060 1077 5212 1083
rect 5220 1077 5292 1083
rect 5332 1077 5372 1083
rect 5444 1077 5532 1083
rect 5620 1077 5724 1083
rect 5780 1077 5859 1083
rect 5853 1064 5859 1077
rect 5988 1077 6108 1083
rect 6164 1077 6316 1083
rect 6324 1077 6348 1083
rect 6356 1077 6412 1083
rect 6564 1077 6636 1083
rect 180 1057 284 1063
rect 564 1057 700 1063
rect 708 1057 764 1063
rect 1044 1057 1132 1063
rect 1140 1057 1404 1063
rect 1476 1057 1516 1063
rect 1572 1057 1724 1063
rect 1732 1057 1836 1063
rect 1956 1057 1980 1063
rect 1988 1057 2028 1063
rect 2292 1057 2348 1063
rect 2836 1057 2892 1063
rect 3860 1057 4156 1063
rect 4516 1057 4556 1063
rect 4628 1057 4652 1063
rect 5092 1057 5116 1063
rect 5284 1057 5308 1063
rect 5780 1057 5788 1063
rect 5828 1057 5836 1063
rect 5860 1057 5884 1063
rect 6132 1057 6156 1063
rect 6228 1057 6268 1063
rect 6276 1057 6524 1063
rect 20 1037 236 1043
rect 1188 1037 1276 1043
rect 1300 1037 1340 1043
rect 1492 1037 1852 1043
rect 4676 1037 4716 1043
rect 4724 1037 4748 1043
rect 5108 1037 5180 1043
rect 5268 1037 5964 1043
rect 5972 1037 6060 1043
rect 6084 1037 6204 1043
rect 6292 1037 6348 1043
rect 6372 1037 6444 1043
rect 6541 1043 6547 1056
rect 6532 1037 6547 1043
rect 356 1017 412 1023
rect 1060 1017 1068 1023
rect 1284 1017 1484 1023
rect 1556 1017 1740 1023
rect 3716 1017 3756 1023
rect 4548 1017 4796 1023
rect 4820 1017 5420 1023
rect 5460 1017 5484 1023
rect 5508 1017 5532 1023
rect 5716 1017 5747 1023
rect 3304 1014 3352 1016
rect 3304 1006 3308 1014
rect 3318 1006 3324 1014
rect 3332 1006 3338 1014
rect 3348 1006 3352 1014
rect 3304 1004 3352 1006
rect 116 997 364 1003
rect 612 997 876 1003
rect 980 997 1036 1003
rect 1060 997 1100 1003
rect 1204 997 1404 1003
rect 1524 997 1628 1003
rect 2100 997 2156 1003
rect 2164 997 2300 1003
rect 3604 997 3788 1003
rect 3796 997 3852 1003
rect 4676 997 5068 1003
rect 5108 997 5276 1003
rect 5396 997 5436 1003
rect 5444 997 5484 1003
rect 5492 997 5724 1003
rect 5741 1003 5747 1017
rect 6196 1017 6204 1023
rect 6372 1017 6572 1023
rect 5741 997 6156 1003
rect 6452 997 6476 1003
rect 84 977 268 983
rect 372 977 412 983
rect 548 977 700 983
rect 868 977 924 983
rect 932 977 1004 983
rect 1028 977 1244 983
rect 1252 977 1532 983
rect 1572 977 1644 983
rect 1652 977 1660 983
rect 2148 977 2364 983
rect 2644 977 2732 983
rect 3149 977 3372 983
rect 3149 964 3155 977
rect 3380 977 3580 983
rect 3684 977 3820 983
rect 3828 977 3836 983
rect 4276 977 4348 983
rect 4468 977 4604 983
rect 4820 977 4892 983
rect 5028 977 5132 983
rect 5380 977 5500 983
rect 5508 977 5708 983
rect 5716 977 5788 983
rect 6004 977 6044 983
rect 6068 977 6092 983
rect 6100 977 6124 983
rect 6196 977 6316 983
rect 6404 977 6460 983
rect 36 957 204 963
rect 500 957 556 963
rect 1012 957 1100 963
rect 1140 957 1187 963
rect 1181 944 1187 957
rect 1332 957 1452 963
rect 1636 957 1875 963
rect 1869 944 1875 957
rect 2292 957 2444 963
rect 3108 957 3148 963
rect 3364 957 3468 963
rect 4132 957 4188 963
rect 4196 957 4284 963
rect 4340 957 4412 963
rect 4420 957 4540 963
rect 4564 957 4668 963
rect 4676 957 4684 963
rect 4788 957 5228 963
rect 5284 957 5596 963
rect 5668 957 5740 963
rect 6228 957 6284 963
rect 6324 957 6348 963
rect 6452 957 6476 963
rect 52 937 76 943
rect 308 937 364 943
rect 468 937 652 943
rect 660 937 716 943
rect 724 937 908 943
rect 916 937 1164 943
rect 1188 937 1388 943
rect 1412 937 1468 943
rect 1476 937 1708 943
rect 1876 937 1996 943
rect 2356 937 2428 943
rect 2564 937 2780 943
rect 2788 937 2844 943
rect 3060 937 3164 943
rect 3380 937 3436 943
rect 3444 937 3468 943
rect 3572 937 3756 943
rect 3956 937 4028 943
rect 4532 937 4588 943
rect 4596 937 4732 943
rect 4740 937 4908 943
rect 4932 937 5036 943
rect 5076 937 5132 943
rect 5140 937 5260 943
rect 5300 937 5404 943
rect 5732 937 5868 943
rect 5972 937 6028 943
rect 6180 937 6252 943
rect 6308 937 6348 943
rect 6420 937 6444 943
rect 6580 937 6604 943
rect 180 917 236 923
rect 260 917 316 923
rect 324 917 396 923
rect 404 917 524 923
rect 644 917 684 923
rect 740 917 812 923
rect 948 917 1020 923
rect 1028 917 1132 923
rect 1396 917 1452 923
rect 1460 917 1500 923
rect 1620 917 1676 923
rect 1684 917 1932 923
rect 1988 917 2012 923
rect 2020 917 2204 923
rect 2420 917 2524 923
rect 2612 917 2668 923
rect 2740 917 2828 923
rect 2900 917 3212 923
rect 3220 917 3420 923
rect 3428 917 3596 923
rect 3604 917 3868 923
rect 4004 917 4108 923
rect 4116 917 4156 923
rect 4452 917 4652 923
rect 4772 917 4956 923
rect 5012 917 5036 923
rect 5156 917 5180 923
rect 5204 917 5228 923
rect 5476 917 5548 923
rect 5620 917 5676 923
rect 5940 917 5964 923
rect 5972 917 5980 923
rect 6052 917 6092 923
rect 6100 917 6108 923
rect 6116 917 6156 923
rect 6244 917 6300 923
rect 6388 917 6412 923
rect 6580 917 6604 923
rect 196 897 332 903
rect 340 897 364 903
rect 420 897 476 903
rect 516 897 572 903
rect 580 897 844 903
rect 852 897 972 903
rect 1108 897 1148 903
rect 1156 897 1196 903
rect 1204 897 1260 903
rect 1316 897 1372 903
rect 1588 897 1692 903
rect 1732 897 1836 903
rect 1844 897 2060 903
rect 2116 897 2188 903
rect 2196 897 2252 903
rect 2276 897 2380 903
rect 2420 897 2492 903
rect 2548 897 2780 903
rect 2788 897 2812 903
rect 3396 897 3500 903
rect 3940 897 3996 903
rect 4260 897 4332 903
rect 4516 897 4700 903
rect 4708 897 4732 903
rect 4964 897 5116 903
rect 5124 897 5148 903
rect 5684 897 5740 903
rect 5876 897 5948 903
rect 5956 897 6092 903
rect 6164 897 6188 903
rect 6324 897 6444 903
rect 164 877 220 883
rect 244 877 268 883
rect 276 877 412 883
rect 436 877 556 883
rect 756 877 828 883
rect 884 877 940 883
rect 1348 877 1532 883
rect 1716 877 1724 883
rect 1748 877 1820 883
rect 1860 877 1932 883
rect 1972 877 2028 883
rect 2036 877 2060 883
rect 2084 877 2140 883
rect 2996 877 3036 883
rect 3044 877 3100 883
rect 3204 877 3244 883
rect 3268 877 3347 883
rect 84 857 156 863
rect 244 857 268 863
rect 1012 857 1036 863
rect 1684 857 1788 863
rect 1828 857 2012 863
rect 2228 857 2508 863
rect 3341 863 3347 877
rect 3364 877 3452 883
rect 3572 877 3596 883
rect 4068 877 4092 883
rect 4100 877 4140 883
rect 4580 877 4636 883
rect 4644 877 5020 883
rect 6004 877 6060 883
rect 6228 877 6284 883
rect 6532 877 6556 883
rect 3341 857 3692 863
rect 4932 857 5132 863
rect 5300 857 5324 863
rect 5716 857 5884 863
rect 5892 857 5964 863
rect 6452 857 6460 863
rect 1764 837 1852 843
rect 1908 837 1980 843
rect 2116 837 2460 843
rect 2612 837 3196 843
rect 3268 837 3916 843
rect 3924 837 4076 843
rect 4628 837 5100 843
rect 5748 837 5772 843
rect 5972 837 5996 843
rect 6260 837 6380 843
rect 6388 837 6460 843
rect 6580 837 6604 843
rect 212 817 252 823
rect 2212 817 2620 823
rect 2708 817 3180 823
rect 3188 817 3564 823
rect 5652 817 6076 823
rect 6244 817 6492 823
rect 1768 814 1816 816
rect 1768 806 1772 814
rect 1782 806 1788 814
rect 1796 806 1802 814
rect 1812 806 1816 814
rect 1768 804 1816 806
rect 4824 814 4872 816
rect 4824 806 4828 814
rect 4838 806 4844 814
rect 4852 806 4858 814
rect 4868 806 4872 814
rect 4824 804 4872 806
rect 372 797 716 803
rect 980 797 1036 803
rect 1204 797 1292 803
rect 2548 797 3276 803
rect 4420 797 4652 803
rect 4660 797 4732 803
rect 6116 797 6268 803
rect 516 777 828 783
rect 1236 777 1244 783
rect 1252 777 1292 783
rect 1588 777 1788 783
rect 1796 777 1996 783
rect 2452 777 2732 783
rect 2740 777 2780 783
rect 3812 777 4332 783
rect 4340 777 4380 783
rect 4388 777 4428 783
rect 6180 777 6268 783
rect 228 757 348 763
rect 356 757 652 763
rect 820 757 844 763
rect 852 757 972 763
rect 1220 757 1388 763
rect 1412 757 1468 763
rect 1908 757 1932 763
rect 1940 757 2012 763
rect 2020 757 2124 763
rect 2516 757 2540 763
rect 3012 757 3660 763
rect 3668 757 3724 763
rect 3780 757 4108 763
rect 4116 757 4156 763
rect 4244 757 4396 763
rect 4404 757 4643 763
rect 4637 744 4643 757
rect 5428 757 5468 763
rect 5988 757 6108 763
rect 6116 757 6172 763
rect 6404 757 6492 763
rect 68 737 92 743
rect 436 737 492 743
rect 532 737 604 743
rect 820 737 860 743
rect 932 737 963 743
rect 957 724 963 737
rect 1236 737 1260 743
rect 1380 737 1436 743
rect 1492 737 1516 743
rect 1860 737 1980 743
rect 1988 737 2220 743
rect 2516 737 2652 743
rect 2660 737 2684 743
rect 2692 737 2764 743
rect 2804 737 3020 743
rect 3028 737 3068 743
rect 3140 737 3228 743
rect 3236 737 3356 743
rect 3892 737 4268 743
rect 4276 737 4364 743
rect 4372 737 4460 743
rect 4564 737 4588 743
rect 4596 737 4620 743
rect 4644 737 4972 743
rect 5044 737 5068 743
rect 5940 737 5964 743
rect 6020 737 6060 743
rect 6340 737 6556 743
rect 196 717 236 723
rect 340 717 444 723
rect 468 717 540 723
rect 580 717 668 723
rect 1268 717 1292 723
rect 1300 717 1308 723
rect 1428 717 1516 723
rect 1540 717 1596 723
rect 1700 717 1756 723
rect 1956 717 2044 723
rect 2468 717 2540 723
rect 2548 717 2572 723
rect 2580 717 2620 723
rect 2628 717 2748 723
rect 3124 717 3164 723
rect 3476 717 3548 723
rect 3620 717 3676 723
rect 3780 717 3804 723
rect 3940 717 4204 723
rect 4212 717 4796 723
rect 4804 717 4908 723
rect 4964 717 5020 723
rect 5028 717 5100 723
rect 5556 717 5644 723
rect 5684 717 5772 723
rect 5780 717 5820 723
rect 5988 717 6044 723
rect 6132 717 6188 723
rect 6388 717 6524 723
rect 6532 717 6604 723
rect 116 697 252 703
rect 292 697 444 703
rect 452 697 508 703
rect 628 697 707 703
rect 701 684 707 697
rect 1092 697 1132 703
rect 1220 697 1228 703
rect 1236 697 1260 703
rect 1268 697 1340 703
rect 1476 697 1532 703
rect 1604 697 1724 703
rect 2084 697 2268 703
rect 2356 697 2396 703
rect 2484 697 2524 703
rect 2532 697 2668 703
rect 2676 697 2700 703
rect 2708 697 2796 703
rect 2900 697 3148 703
rect 3156 697 3196 703
rect 4132 697 4540 703
rect 4548 697 4716 703
rect 4724 697 4988 703
rect 4996 697 5004 703
rect 5044 697 5164 703
rect 5172 697 5228 703
rect 5380 697 5404 703
rect 5428 697 5516 703
rect 5812 697 5836 703
rect 5933 697 5996 703
rect 5933 684 5939 697
rect 6036 697 6236 703
rect 6260 697 6300 703
rect 6356 697 6380 703
rect 6452 697 6476 703
rect 6564 697 6620 703
rect 36 677 156 683
rect 164 677 204 683
rect 564 677 652 683
rect 708 677 940 683
rect 1092 677 1116 683
rect 1124 677 1148 683
rect 1892 677 1916 683
rect 1924 677 1996 683
rect 2004 677 2092 683
rect 2564 677 2588 683
rect 2676 677 2700 683
rect 2852 677 2924 683
rect 3092 677 3132 683
rect 3140 677 3180 683
rect 3236 677 3372 683
rect 3572 677 3628 683
rect 3684 677 3772 683
rect 4084 677 4124 683
rect 4164 677 4220 683
rect 4260 677 4348 683
rect 4356 677 4556 683
rect 4564 677 4700 683
rect 4740 677 4844 683
rect 4916 677 5260 683
rect 5380 677 5500 683
rect 5652 677 5756 683
rect 5796 677 5932 683
rect 5972 677 6044 683
rect 6164 677 6252 683
rect 6276 677 6348 683
rect 6404 677 6428 683
rect 6452 677 6588 683
rect 13 663 19 676
rect 13 657 140 663
rect 164 657 220 663
rect 548 657 604 663
rect 836 657 1180 663
rect 1348 657 1356 663
rect 1364 657 1420 663
rect 1428 657 1452 663
rect 1588 657 1612 663
rect 1876 657 2140 663
rect 2292 657 2316 663
rect 2324 657 2364 663
rect 2436 657 2508 663
rect 2548 657 2556 663
rect 2756 657 2956 663
rect 2964 657 3036 663
rect 3380 657 3452 663
rect 3508 657 3548 663
rect 3604 657 3692 663
rect 3700 657 3884 663
rect 3892 657 3980 663
rect 4116 657 4172 663
rect 4468 657 4508 663
rect 4516 657 4572 663
rect 4580 657 4780 663
rect 5044 657 5116 663
rect 5124 657 5212 663
rect 5220 657 5308 663
rect 5460 657 5676 663
rect 6132 657 6220 663
rect 6260 657 6332 663
rect 6372 657 6604 663
rect 132 637 156 643
rect 468 637 876 643
rect 980 637 1212 643
rect 2020 637 2092 643
rect 2100 637 2300 643
rect 2500 637 2860 643
rect 3012 637 3260 643
rect 3412 637 3820 643
rect 3844 637 3916 643
rect 4180 637 4524 643
rect 4532 637 4684 643
rect 4692 637 4748 643
rect 4788 637 4828 643
rect 4836 637 4924 643
rect 5517 637 5804 643
rect 5517 624 5523 637
rect 5812 637 5852 643
rect 6020 637 6227 643
rect 404 617 556 623
rect 708 617 1036 623
rect 1428 617 1692 623
rect 2052 617 2060 623
rect 2100 617 2572 623
rect 2628 617 2972 623
rect 2980 617 3052 623
rect 3460 617 3564 623
rect 3604 617 3644 623
rect 3684 617 3788 623
rect 3796 617 4028 623
rect 4036 617 4060 623
rect 4372 617 4604 623
rect 4628 617 4812 623
rect 4836 617 5084 623
rect 5188 617 5516 623
rect 5668 617 5788 623
rect 5924 617 6092 623
rect 6100 617 6140 623
rect 6221 623 6227 637
rect 6244 637 6396 643
rect 6404 637 6460 643
rect 6221 617 6444 623
rect 3304 614 3352 616
rect 3304 606 3308 614
rect 3318 606 3324 614
rect 3332 606 3338 614
rect 3348 606 3352 614
rect 3304 604 3352 606
rect 692 597 1084 603
rect 1188 597 1212 603
rect 1220 597 1356 603
rect 1380 597 1596 603
rect 2036 597 2044 603
rect 2516 597 2604 603
rect 2612 597 2780 603
rect 2996 597 3052 603
rect 3060 597 3180 603
rect 3428 597 3948 603
rect 3981 597 4476 603
rect 116 577 188 583
rect 196 577 332 583
rect 692 577 780 583
rect 788 577 844 583
rect 852 577 1020 583
rect 1332 577 1548 583
rect 1636 577 1692 583
rect 1700 577 2140 583
rect 2740 577 2812 583
rect 2820 577 2940 583
rect 2948 577 3372 583
rect 3396 577 3468 583
rect 3540 577 3836 583
rect 3981 583 3987 597
rect 4532 597 4796 603
rect 4804 597 5132 603
rect 5380 597 5388 603
rect 5620 597 6364 603
rect 6548 597 6572 603
rect 3892 577 3987 583
rect 3997 577 4316 583
rect 244 557 300 563
rect 340 557 460 563
rect 532 557 764 563
rect 884 557 924 563
rect 932 557 956 563
rect 1092 557 1196 563
rect 1412 557 1660 563
rect 2004 557 2108 563
rect 2132 557 2444 563
rect 2676 557 2748 563
rect 2756 557 2956 563
rect 2964 557 3116 563
rect 3172 557 3196 563
rect 3268 557 3276 563
rect 3364 557 3708 563
rect 3716 557 3772 563
rect 3789 557 3820 563
rect 148 537 204 543
rect 228 537 284 543
rect 308 537 364 543
rect 372 537 428 543
rect 596 537 764 543
rect 772 537 956 543
rect 964 537 1004 543
rect 1076 537 1132 543
rect 1140 537 1260 543
rect 1396 537 1484 543
rect 1524 537 1596 543
rect 1604 537 1740 543
rect 2228 537 2268 543
rect 2276 537 2300 543
rect 2317 537 2428 543
rect 20 517 124 523
rect 132 517 380 523
rect 420 517 508 523
rect 532 517 604 523
rect 756 517 796 523
rect 868 517 940 523
rect 1044 517 1132 523
rect 1236 517 1260 523
rect 1460 517 1516 523
rect 1668 517 1708 523
rect 1716 517 1836 523
rect 2317 523 2323 537
rect 2852 537 2892 543
rect 2900 537 3036 543
rect 3044 537 3379 543
rect 2308 517 2323 523
rect 2388 517 2460 523
rect 2564 517 2604 523
rect 2644 517 2988 523
rect 3156 517 3196 523
rect 3204 517 3356 523
rect 3373 523 3379 537
rect 3444 537 3484 543
rect 3540 537 3628 543
rect 3652 537 3724 543
rect 3789 543 3795 557
rect 3844 557 3900 563
rect 3924 557 3948 563
rect 3997 563 4003 577
rect 4420 577 5068 583
rect 5092 577 5347 583
rect 5341 564 5347 577
rect 5364 577 5420 583
rect 5508 577 5676 583
rect 5876 577 6172 583
rect 6436 577 6492 583
rect 6516 577 6540 583
rect 3956 557 4003 563
rect 4324 557 4364 563
rect 4532 557 4556 563
rect 4596 557 4652 563
rect 4692 557 4764 563
rect 4788 557 4812 563
rect 4820 557 4908 563
rect 5172 557 5212 563
rect 5316 557 5324 563
rect 5348 557 5484 563
rect 5492 557 5612 563
rect 5748 557 5804 563
rect 5908 557 6140 563
rect 6244 557 6268 563
rect 6516 557 6572 563
rect 3764 537 3795 543
rect 3828 537 3884 543
rect 4004 537 4060 543
rect 4276 537 4332 543
rect 4340 537 4556 543
rect 4781 543 4787 556
rect 4676 537 4787 543
rect 5012 537 5116 543
rect 5140 537 5292 543
rect 5300 537 5388 543
rect 5396 537 5564 543
rect 5604 537 5708 543
rect 5844 537 5916 543
rect 5956 537 6060 543
rect 6244 537 6252 543
rect 6276 537 6316 543
rect 6340 537 6716 543
rect 3373 517 3612 523
rect 3636 517 4012 523
rect 4084 517 4147 523
rect 292 497 588 503
rect 596 497 652 503
rect 1028 497 1244 503
rect 1508 497 1852 503
rect 1860 497 1900 503
rect 2116 497 2268 503
rect 2276 497 2364 503
rect 2388 497 2476 503
rect 2484 497 2652 503
rect 2708 497 2876 503
rect 2884 497 2972 503
rect 3348 497 3436 503
rect 3476 497 3500 503
rect 3629 503 3635 516
rect 4141 504 4147 517
rect 4228 517 4284 523
rect 4356 517 4588 523
rect 4756 517 4828 523
rect 4932 517 5196 523
rect 5604 517 5660 523
rect 5700 517 5740 523
rect 5924 517 5980 523
rect 6084 517 6227 523
rect 3556 497 3635 503
rect 3732 497 3788 503
rect 3844 497 3884 503
rect 3924 497 3996 503
rect 4020 497 4108 503
rect 4148 497 4188 503
rect 4349 503 4355 516
rect 4260 497 4355 503
rect 4388 497 4428 503
rect 4500 497 4940 503
rect 4964 497 5004 503
rect 5060 497 5132 503
rect 5684 497 5724 503
rect 5732 497 5756 503
rect 5764 497 5884 503
rect 5956 497 6076 503
rect 6164 497 6204 503
rect 6221 503 6227 517
rect 6324 517 6444 523
rect 6221 497 6492 503
rect 276 477 300 483
rect 308 477 348 483
rect 372 477 412 483
rect 516 477 572 483
rect 1060 477 1116 483
rect 1124 477 1180 483
rect 1444 477 1532 483
rect 1540 477 1580 483
rect 1700 477 1820 483
rect 2404 477 2428 483
rect 2436 477 2556 483
rect 2740 477 2764 483
rect 2868 477 3004 483
rect 3012 477 3068 483
rect 3076 477 3244 483
rect 3332 477 3388 483
rect 3428 477 3852 483
rect 3860 477 3900 483
rect 3924 477 3980 483
rect 3988 477 4044 483
rect 4276 477 4412 483
rect 5556 477 5580 483
rect 5588 477 5644 483
rect 5972 477 6012 483
rect 6228 477 6252 483
rect 6532 477 6572 483
rect 324 457 460 463
rect 900 457 988 463
rect 1300 457 2092 463
rect 2820 457 3052 463
rect 3252 457 3644 463
rect 3652 457 3708 463
rect 3732 457 4060 463
rect 4068 457 4124 463
rect 4132 457 4156 463
rect 5060 457 5180 463
rect 5412 457 5916 463
rect 5940 457 6188 463
rect 388 437 476 443
rect 596 437 1308 443
rect 1684 437 1868 443
rect 2020 437 2236 443
rect 2436 437 2572 443
rect 2580 437 2812 443
rect 3860 437 4092 443
rect 4100 437 4108 443
rect 4116 437 4172 443
rect 4708 437 4828 443
rect 4836 437 5244 443
rect 5252 437 5292 443
rect 5908 437 6572 443
rect 420 417 444 423
rect 660 417 684 423
rect 852 417 1388 423
rect 1540 417 1628 423
rect 2004 417 2588 423
rect 4004 417 4412 423
rect 4420 417 4460 423
rect 4468 417 4540 423
rect 5668 417 5996 423
rect 6004 417 6124 423
rect 6388 417 6636 423
rect 1768 414 1816 416
rect 1768 406 1772 414
rect 1782 406 1788 414
rect 1796 406 1802 414
rect 1812 406 1816 414
rect 1768 404 1816 406
rect 4824 414 4872 416
rect 4824 406 4828 414
rect 4838 406 4844 414
rect 4852 406 4858 414
rect 4868 406 4872 414
rect 4824 404 4872 406
rect 244 397 252 403
rect 260 397 524 403
rect 564 397 588 403
rect 596 397 860 403
rect 884 397 956 403
rect 1604 397 1740 403
rect 1844 397 2028 403
rect 2052 397 2060 403
rect 2212 397 2492 403
rect 3540 397 3724 403
rect 3732 397 3852 403
rect 3860 397 3932 403
rect 6244 397 6412 403
rect 196 377 364 383
rect 452 377 524 383
rect 548 377 604 383
rect 612 377 716 383
rect 740 377 796 383
rect 820 377 1388 383
rect 1636 377 2476 383
rect 2484 377 2508 383
rect 2740 377 3020 383
rect 3028 377 3116 383
rect 3300 377 3404 383
rect 3428 377 3532 383
rect 3540 377 3580 383
rect 4356 377 4556 383
rect 4564 377 4684 383
rect 5108 377 5788 383
rect 5844 377 6028 383
rect 6036 377 6092 383
rect 6420 377 6444 383
rect 228 357 284 363
rect 292 357 380 363
rect 404 357 428 363
rect 436 357 572 363
rect 628 357 771 363
rect 765 344 771 357
rect 788 357 1068 363
rect 1444 357 1516 363
rect 1524 357 1628 363
rect 1700 357 2060 363
rect 2100 357 2668 363
rect 2676 357 2732 363
rect 2740 357 2780 363
rect 2820 357 3228 363
rect 3236 357 3308 363
rect 3476 357 3884 363
rect 3924 357 3948 363
rect 4036 357 4220 363
rect 4308 357 4396 363
rect 4404 357 4524 363
rect 5748 357 6188 363
rect 6404 357 6428 363
rect 6548 357 6604 363
rect 84 337 140 343
rect 148 337 364 343
rect 420 337 668 343
rect 772 337 988 343
rect 1140 337 1260 343
rect 1396 337 1484 343
rect 1588 337 1612 343
rect 1620 337 1708 343
rect 1764 337 1836 343
rect 1876 337 2460 343
rect 2468 337 2524 343
rect 2573 337 2748 343
rect 2573 324 2579 337
rect 2868 337 3004 343
rect 3012 337 3084 343
rect 3108 337 3404 343
rect 3444 337 3452 343
rect 3604 337 3900 343
rect 3908 337 3964 343
rect 4132 337 4428 343
rect 4436 337 4444 343
rect 4452 337 4508 343
rect 4596 337 4652 343
rect 5412 337 5452 343
rect 5636 337 5820 343
rect 5828 337 5852 343
rect 5892 337 6076 343
rect 6356 337 6428 343
rect 212 317 268 323
rect 356 317 460 323
rect 500 317 524 323
rect 564 317 668 323
rect 692 317 716 323
rect 724 317 780 323
rect 788 317 876 323
rect 884 317 908 323
rect 980 317 1148 323
rect 1380 317 1564 323
rect 1636 317 1692 323
rect 1748 317 1868 323
rect 1892 317 2028 323
rect 2116 317 2188 323
rect 2276 317 2364 323
rect 2484 317 2572 323
rect 2612 317 2796 323
rect 2804 317 2828 323
rect 2948 317 2972 323
rect 3101 323 3107 336
rect 3060 317 3107 323
rect 3156 317 3244 323
rect 3252 317 3276 323
rect 3284 317 3388 323
rect 3412 317 3516 323
rect 3524 317 3596 323
rect 3620 317 3644 323
rect 3764 317 3804 323
rect 3828 317 3868 323
rect 3876 317 4028 323
rect 4132 317 4195 323
rect 276 297 316 303
rect 333 297 924 303
rect 52 277 108 283
rect 116 277 172 283
rect 333 283 339 297
rect 948 297 1068 303
rect 1508 297 1708 303
rect 1885 303 1891 316
rect 4189 304 4195 317
rect 4260 317 4380 323
rect 4484 317 4556 323
rect 4884 317 5068 323
rect 5188 317 5212 323
rect 5332 317 5932 323
rect 6068 317 6124 323
rect 6180 317 6252 323
rect 6372 317 6508 323
rect 1716 297 1891 303
rect 1908 297 2012 303
rect 2068 297 2092 303
rect 2100 297 2124 303
rect 2260 297 2316 303
rect 2324 297 2380 303
rect 2500 297 2556 303
rect 2596 297 3484 303
rect 3636 297 3660 303
rect 3716 297 3820 303
rect 3892 297 3948 303
rect 4020 297 4076 303
rect 4084 297 4140 303
rect 4196 297 4236 303
rect 4244 297 4268 303
rect 4340 297 4572 303
rect 4804 297 4956 303
rect 5124 297 5228 303
rect 5252 297 5388 303
rect 5780 297 5804 303
rect 5812 297 5868 303
rect 6084 297 6300 303
rect 6308 297 6476 303
rect 180 277 339 283
rect 372 277 780 283
rect 820 277 876 283
rect 932 277 988 283
rect 1092 277 1148 283
rect 1204 277 1244 283
rect 1524 277 1564 283
rect 1572 277 1644 283
rect 1652 277 1724 283
rect 1828 277 2076 283
rect 2084 277 2140 283
rect 2180 277 2636 283
rect 2692 277 2716 283
rect 2724 277 2956 283
rect 2980 277 3132 283
rect 3156 277 3196 283
rect 3204 277 3292 283
rect 3357 277 3404 283
rect 20 257 156 263
rect 340 257 476 263
rect 484 257 780 263
rect 804 257 1100 263
rect 1124 257 1187 263
rect 84 237 108 243
rect 500 237 1148 243
rect 1181 243 1187 257
rect 1204 257 1292 263
rect 1332 257 1548 263
rect 1716 257 1836 263
rect 1876 257 2220 263
rect 2340 257 2572 263
rect 2612 257 2620 263
rect 2644 257 2876 263
rect 2900 257 3052 263
rect 3357 263 3363 277
rect 3629 283 3635 296
rect 3428 277 3635 283
rect 3700 277 3772 283
rect 3780 277 3804 283
rect 3940 277 4108 283
rect 4244 277 4332 283
rect 4660 277 4764 283
rect 5156 277 5212 283
rect 5220 277 5276 283
rect 5316 277 5372 283
rect 5620 277 5660 283
rect 5668 277 5772 283
rect 5796 277 5900 283
rect 5924 277 6284 283
rect 6484 277 6604 283
rect 6628 277 6636 283
rect 3188 257 3363 263
rect 3380 257 3692 263
rect 3764 257 3916 263
rect 4004 257 4092 263
rect 4132 257 4268 263
rect 4548 257 4716 263
rect 4724 257 4780 263
rect 4932 257 5084 263
rect 5284 257 5340 263
rect 5364 257 5596 263
rect 5844 257 5964 263
rect 6020 257 6060 263
rect 6164 257 6636 263
rect 1181 237 1235 243
rect 452 217 1212 223
rect 1229 223 1235 237
rect 1300 237 1548 243
rect 1556 237 2012 243
rect 2020 237 2156 243
rect 2260 237 2380 243
rect 2612 237 2732 243
rect 2740 237 3612 243
rect 3780 237 4156 243
rect 4212 237 4844 243
rect 5012 237 5676 243
rect 5684 237 5724 243
rect 6020 237 6124 243
rect 6180 237 6204 243
rect 6260 237 6348 243
rect 1229 217 1324 223
rect 1412 217 2156 223
rect 2164 217 2332 223
rect 2532 217 2668 223
rect 2685 217 3036 223
rect 372 197 732 203
rect 756 197 844 203
rect 868 197 1020 203
rect 1044 197 1100 203
rect 1108 197 1260 203
rect 1284 197 2028 203
rect 2052 197 2284 203
rect 2685 203 2691 217
rect 3060 217 3212 223
rect 3236 217 3244 223
rect 3380 217 3788 223
rect 3812 217 3868 223
rect 3876 217 3948 223
rect 3956 217 4476 223
rect 5636 217 6076 223
rect 6356 217 6556 223
rect 3304 214 3352 216
rect 3304 206 3308 214
rect 3318 206 3324 214
rect 3332 206 3338 214
rect 3348 206 3352 214
rect 3304 204 3352 206
rect 2644 197 2691 203
rect 2804 197 3036 203
rect 3076 197 3084 203
rect 3124 197 3212 203
rect 3412 197 3468 203
rect 3588 197 3820 203
rect 5940 197 6076 203
rect 6164 197 6620 203
rect 436 177 492 183
rect 532 177 652 183
rect 660 177 1436 183
rect 1620 177 1804 183
rect 1812 177 2652 183
rect 2676 177 2892 183
rect 2948 177 3132 183
rect 3156 177 3276 183
rect 3364 177 3516 183
rect 3524 177 3932 183
rect 4004 177 4684 183
rect 4804 177 5036 183
rect 5668 177 5740 183
rect 5972 177 6396 183
rect 372 157 412 163
rect 420 157 492 163
rect 500 157 828 163
rect 900 157 1068 163
rect 1092 157 1116 163
rect 1172 157 1260 163
rect 1268 157 1932 163
rect 1972 157 2108 163
rect 2308 157 2876 163
rect 2900 157 2972 163
rect 2996 157 3004 163
rect 3044 157 3436 163
rect 3636 157 3660 163
rect 3668 157 3884 163
rect 4436 157 4668 163
rect 4676 157 4972 163
rect 4980 157 5308 163
rect 5316 157 5420 163
rect 5428 157 5516 163
rect 5524 157 5788 163
rect 6148 157 6284 163
rect 6308 157 6492 163
rect 6516 157 6524 163
rect 100 137 236 143
rect 308 137 348 143
rect 404 137 460 143
rect 468 137 636 143
rect 740 137 764 143
rect 788 137 796 143
rect 893 143 899 156
rect 820 137 899 143
rect 948 137 1004 143
rect 1028 137 1260 143
rect 1268 137 1388 143
rect 1396 137 1484 143
rect 1588 137 1660 143
rect 1684 137 2284 143
rect 2292 137 2348 143
rect 2388 137 2444 143
rect 2452 137 2524 143
rect 2676 137 2700 143
rect 2708 137 3084 143
rect 3092 137 3436 143
rect 3652 137 3708 143
rect 3716 137 3788 143
rect 3876 137 3980 143
rect 4164 137 4620 143
rect 4980 137 5011 143
rect 612 117 732 123
rect 740 117 860 123
rect 900 117 1244 123
rect 1252 117 1372 123
rect 1380 117 1468 123
rect 1492 117 1516 123
rect 1565 123 1571 136
rect 1565 117 1900 123
rect 1924 117 1996 123
rect 2084 117 2428 123
rect 2436 117 2492 123
rect 2564 117 2716 123
rect 2724 117 3260 123
rect 3284 117 3404 123
rect 3444 117 3756 123
rect 3828 117 3916 123
rect 4404 117 4524 123
rect 4644 117 4764 123
rect 4916 117 4988 123
rect 5005 123 5011 137
rect 5028 137 5052 143
rect 5748 137 5916 143
rect 6052 137 6092 143
rect 6100 137 6124 143
rect 6180 137 6236 143
rect 6292 137 6332 143
rect 6420 137 6444 143
rect 6484 137 6620 143
rect 5005 117 5052 123
rect 5060 117 5180 123
rect 5284 117 5324 123
rect 5412 117 5644 123
rect 5860 117 5916 123
rect 6132 117 6300 123
rect 6324 117 6380 123
rect 564 97 620 103
rect 692 97 748 103
rect 804 97 1580 103
rect 1588 97 1820 103
rect 1828 97 1900 103
rect 1908 97 1948 103
rect 1988 97 2044 103
rect 2084 97 2108 103
rect 2132 97 2268 103
rect 2324 97 2508 103
rect 2516 97 2636 103
rect 2724 97 3420 103
rect 3428 97 3500 103
rect 3508 97 3564 103
rect 3636 97 3772 103
rect 3924 97 3948 103
rect 3956 97 4012 103
rect 4900 97 5036 103
rect 5108 97 5148 103
rect 6196 97 6316 103
rect 6356 97 6396 103
rect 6468 97 6540 103
rect 356 77 444 83
rect 548 77 588 83
rect 676 77 716 83
rect 740 77 940 83
rect 964 77 1564 83
rect 1572 77 1772 83
rect 1780 77 1884 83
rect 1892 77 1932 83
rect 1956 77 2092 83
rect 2148 77 2412 83
rect 2420 77 2476 83
rect 2500 77 2764 83
rect 2772 77 2844 83
rect 2884 77 2956 83
rect 2980 77 3372 83
rect 3396 77 3420 83
rect 3460 77 3484 83
rect 3492 77 3548 83
rect 3572 77 3836 83
rect 3844 77 3900 83
rect 4948 77 5068 83
rect 5076 77 5116 83
rect 6068 77 6156 83
rect 6196 77 6428 83
rect 6580 77 6636 83
rect 548 57 652 63
rect 676 57 700 63
rect 724 57 1308 63
rect 1348 57 1644 63
rect 1796 57 2300 63
rect 2308 57 2364 63
rect 2388 57 2476 63
rect 2500 57 2748 63
rect 2756 57 2828 63
rect 2868 57 2908 63
rect 2916 57 2924 63
rect 2964 57 3244 63
rect 3268 57 3395 63
rect 612 37 972 43
rect 1732 37 1820 43
rect 2436 37 2796 43
rect 2820 37 3052 43
rect 3060 37 3372 43
rect 3389 43 3395 57
rect 3508 57 3612 63
rect 3620 57 3676 63
rect 3780 57 4044 63
rect 6292 57 6364 63
rect 3389 37 3724 43
rect 6244 37 6371 43
rect 6365 24 6371 37
rect 6420 37 6460 43
rect 6500 37 6636 43
rect 2804 17 2940 23
rect 2964 17 3020 23
rect 3044 17 3100 23
rect 3188 17 3260 23
rect 3284 17 3980 23
rect 5620 17 6252 23
rect 6276 17 6300 23
rect 6324 17 6348 23
rect 6388 17 6492 23
rect 6548 17 6572 23
rect 1768 14 1816 16
rect 1768 6 1772 14
rect 1782 6 1788 14
rect 1796 6 1802 14
rect 1812 6 1816 14
rect 1768 4 1816 6
rect 4824 14 4872 16
rect 4824 6 4828 14
rect 4838 6 4844 14
rect 4852 6 4858 14
rect 4868 6 4872 14
rect 4824 4 4872 6
<< m4contact >>
rect 1772 4806 1774 4814
rect 1774 4806 1780 4814
rect 1788 4806 1796 4814
rect 1804 4806 1810 4814
rect 1810 4806 1812 4814
rect 4828 4806 4830 4814
rect 4830 4806 4836 4814
rect 4844 4806 4852 4814
rect 4860 4806 4866 4814
rect 4866 4806 4868 4814
rect 2572 4796 2580 4804
rect 3148 4756 3156 4764
rect 6572 4756 6580 4764
rect 12 4736 20 4744
rect 940 4736 948 4744
rect 6316 4736 6324 4744
rect 1852 4716 1860 4724
rect 1996 4716 2004 4724
rect 2156 4716 2164 4724
rect 2188 4716 2196 4724
rect 2252 4716 2260 4724
rect 2316 4716 2324 4724
rect 2572 4716 2580 4724
rect 2732 4716 2740 4724
rect 2988 4716 2996 4724
rect 3020 4716 3028 4724
rect 3788 4716 3796 4724
rect 5164 4716 5172 4724
rect 6540 4716 6548 4724
rect 12 4696 20 4704
rect 1004 4696 1012 4704
rect 1036 4696 1044 4704
rect 1196 4696 1204 4704
rect 6476 4696 6484 4704
rect 892 4676 900 4684
rect 1116 4676 1124 4684
rect 76 4656 84 4664
rect 1948 4676 1956 4684
rect 1980 4676 1988 4684
rect 2732 4676 2740 4684
rect 2988 4676 2996 4684
rect 5868 4676 5876 4684
rect 6156 4676 6164 4684
rect 2636 4656 2644 4664
rect 6028 4656 6036 4664
rect 6604 4656 6612 4664
rect 1292 4636 1300 4644
rect 1420 4636 1428 4644
rect 1596 4636 1604 4644
rect 5868 4636 5876 4644
rect 3308 4606 3310 4614
rect 3310 4606 3316 4614
rect 3324 4606 3332 4614
rect 3340 4606 3346 4614
rect 3346 4606 3348 4614
rect 1548 4596 1556 4604
rect 3148 4596 3156 4604
rect 6444 4616 6452 4624
rect 5868 4596 5876 4604
rect 1292 4576 1300 4584
rect 1548 4556 1556 4564
rect 2252 4576 2260 4584
rect 5516 4576 5524 4584
rect 6060 4576 6068 4584
rect 6604 4576 6612 4584
rect 6636 4576 6644 4584
rect 4652 4556 4660 4564
rect 5388 4556 5396 4564
rect 2668 4536 2676 4544
rect 6028 4536 6036 4544
rect 6604 4536 6612 4544
rect 396 4516 404 4524
rect 12 4496 20 4504
rect 364 4496 372 4504
rect 3020 4496 3028 4504
rect 2348 4476 2356 4484
rect 4652 4476 4660 4484
rect 5580 4476 5588 4484
rect 268 4456 276 4464
rect 1324 4456 1332 4464
rect 4748 4456 4756 4464
rect 5772 4456 5780 4464
rect 6412 4436 6420 4444
rect 396 4396 404 4404
rect 2636 4416 2644 4424
rect 3660 4416 3668 4424
rect 3788 4416 3796 4424
rect 5164 4416 5172 4424
rect 1772 4406 1774 4414
rect 1774 4406 1780 4414
rect 1788 4406 1796 4414
rect 1804 4406 1810 4414
rect 1810 4406 1812 4414
rect 4828 4406 4830 4414
rect 4830 4406 4836 4414
rect 4844 4406 4852 4414
rect 4860 4406 4866 4414
rect 4866 4406 4868 4414
rect 1324 4396 1332 4404
rect 12 4376 20 4384
rect 44 4356 52 4364
rect 4108 4376 4116 4384
rect 5804 4356 5812 4364
rect 236 4336 244 4344
rect 2860 4336 2868 4344
rect 3212 4316 3220 4324
rect 3948 4316 3956 4324
rect 6284 4316 6292 4324
rect 140 4296 148 4304
rect 716 4296 724 4304
rect 2220 4296 2228 4304
rect 2700 4296 2708 4304
rect 4364 4296 4372 4304
rect 6028 4296 6036 4304
rect 6316 4296 6324 4304
rect 3948 4276 3956 4284
rect 4716 4276 4724 4284
rect 6444 4276 6452 4284
rect 12 4256 20 4264
rect 332 4256 340 4264
rect 780 4256 788 4264
rect 2188 4256 2196 4264
rect 4076 4256 4084 4264
rect 6572 4256 6580 4264
rect 268 4236 276 4244
rect 428 4236 436 4244
rect 5932 4236 5940 4244
rect 1068 4216 1076 4224
rect 5132 4216 5140 4224
rect 3308 4206 3310 4214
rect 3310 4206 3316 4214
rect 3324 4206 3332 4214
rect 3340 4206 3346 4214
rect 3346 4206 3348 4214
rect 3564 4196 3572 4204
rect 5996 4196 6004 4204
rect 76 4176 84 4184
rect 2220 4176 2228 4184
rect 2988 4176 2996 4184
rect 4748 4176 4756 4184
rect 6444 4176 6452 4184
rect 2860 4156 2868 4164
rect 3564 4156 3572 4164
rect 5068 4156 5076 4164
rect 5772 4156 5780 4164
rect 6380 4156 6388 4164
rect 6092 4136 6100 4144
rect 6188 4136 6196 4144
rect 6348 4136 6356 4144
rect 12 4096 20 4104
rect 780 4096 788 4104
rect 2348 4096 2356 4104
rect 4460 4116 4468 4124
rect 3212 4096 3220 4104
rect 6092 4096 6100 4104
rect 140 4076 148 4084
rect 236 4076 244 4084
rect 6028 4076 6036 4084
rect 5004 4056 5012 4064
rect 5868 4056 5876 4064
rect 2508 4036 2516 4044
rect 6220 4036 6228 4044
rect 6348 4016 6356 4024
rect 6444 4016 6452 4024
rect 1772 4006 1774 4014
rect 1774 4006 1780 4014
rect 1788 4006 1796 4014
rect 1804 4006 1810 4014
rect 1810 4006 1812 4014
rect 4828 4006 4830 4014
rect 4830 4006 4836 4014
rect 4844 4006 4852 4014
rect 4860 4006 4866 4014
rect 4866 4006 4868 4014
rect 2668 3996 2676 4004
rect 2860 3996 2868 4004
rect 5036 3996 5044 4004
rect 5772 3996 5780 4004
rect 4716 3956 4724 3964
rect 6316 3936 6324 3944
rect 6604 3936 6612 3944
rect 220 3916 228 3924
rect 5212 3916 5220 3924
rect 3820 3896 3828 3904
rect 5196 3896 5204 3904
rect 5996 3896 6004 3904
rect 6092 3896 6100 3904
rect 6604 3896 6612 3904
rect 188 3876 196 3884
rect 4108 3876 4116 3884
rect 6316 3876 6324 3884
rect 6444 3876 6452 3884
rect 3628 3856 3636 3864
rect 5004 3856 5012 3864
rect 2060 3836 2068 3844
rect 6060 3836 6068 3844
rect 2604 3816 2612 3824
rect 5100 3816 5108 3824
rect 3308 3806 3310 3814
rect 3310 3806 3316 3814
rect 3324 3806 3332 3814
rect 3340 3806 3346 3814
rect 3346 3806 3348 3814
rect 4908 3796 4916 3804
rect 6092 3796 6100 3804
rect 6316 3796 6324 3804
rect 6348 3796 6356 3804
rect 6444 3796 6452 3804
rect 6508 3796 6516 3804
rect 6572 3796 6580 3804
rect 2892 3776 2900 3784
rect 3628 3776 3636 3784
rect 5132 3776 5140 3784
rect 5356 3776 5364 3784
rect 4364 3756 4372 3764
rect 6444 3756 6452 3764
rect 6508 3756 6516 3764
rect 716 3736 724 3744
rect 2316 3736 2324 3744
rect 3660 3736 3668 3744
rect 5036 3736 5044 3744
rect 5516 3736 5524 3744
rect 5804 3736 5812 3744
rect 5996 3736 6004 3744
rect 6060 3736 6068 3744
rect 6124 3736 6132 3744
rect 5708 3716 5716 3724
rect 6604 3736 6612 3744
rect 2860 3696 2868 3704
rect 4108 3696 4116 3704
rect 5100 3696 5108 3704
rect 5132 3696 5140 3704
rect 5388 3696 5396 3704
rect 5740 3696 5748 3704
rect 6188 3696 6196 3704
rect 5420 3676 5428 3684
rect 5964 3676 5972 3684
rect 2028 3656 2036 3664
rect 3820 3656 3828 3664
rect 5100 3656 5108 3664
rect 204 3636 212 3644
rect 5356 3636 5364 3644
rect 6444 3636 6452 3644
rect 6220 3616 6228 3624
rect 6316 3616 6324 3624
rect 1772 3606 1774 3614
rect 1774 3606 1780 3614
rect 1788 3606 1796 3614
rect 1804 3606 1810 3614
rect 1810 3606 1812 3614
rect 4828 3606 4830 3614
rect 4830 3606 4836 3614
rect 4844 3606 4852 3614
rect 4860 3606 4866 3614
rect 4866 3606 4868 3614
rect 4972 3596 4980 3604
rect 6188 3596 6196 3604
rect 2732 3576 2740 3584
rect 4076 3576 4084 3584
rect 2028 3556 2036 3564
rect 6572 3576 6580 3584
rect 6092 3556 6100 3564
rect 2892 3536 2900 3544
rect 4460 3536 4468 3544
rect 5804 3536 5812 3544
rect 6508 3536 6516 3544
rect 3660 3516 3668 3524
rect 6188 3516 6196 3524
rect 6220 3516 6228 3524
rect 3084 3496 3092 3504
rect 428 3476 436 3484
rect 6572 3496 6580 3504
rect 2828 3456 2836 3464
rect 5612 3476 5620 3484
rect 5580 3456 5588 3464
rect 5996 3456 6004 3464
rect 6028 3456 6036 3464
rect 6124 3456 6132 3464
rect 5772 3436 5780 3444
rect 5836 3436 5844 3444
rect 3884 3416 3892 3424
rect 4236 3416 4244 3424
rect 5964 3416 5972 3424
rect 6188 3416 6196 3424
rect 3308 3406 3310 3414
rect 3310 3406 3316 3414
rect 3324 3406 3332 3414
rect 3340 3406 3346 3414
rect 3346 3406 3348 3414
rect 2316 3396 2324 3404
rect 4044 3396 4052 3404
rect 5772 3396 5780 3404
rect 6444 3396 6452 3404
rect 6572 3396 6580 3404
rect 3660 3376 3668 3384
rect 4972 3376 4980 3384
rect 4268 3356 4276 3364
rect 6156 3356 6164 3364
rect 12 3336 20 3344
rect 44 3336 52 3344
rect 1740 3336 1748 3344
rect 6604 3336 6612 3344
rect 1068 3316 1076 3324
rect 5708 3316 5716 3324
rect 5740 3316 5748 3324
rect 5964 3316 5972 3324
rect 6572 3316 6580 3324
rect 2060 3296 2068 3304
rect 2476 3296 2484 3304
rect 2668 3296 2676 3304
rect 4620 3296 4628 3304
rect 5420 3256 5428 3264
rect 876 3236 884 3244
rect 1740 3216 1748 3224
rect 3724 3216 3732 3224
rect 4940 3236 4948 3244
rect 6124 3216 6132 3224
rect 6444 3216 6452 3224
rect 1772 3206 1774 3214
rect 1774 3206 1780 3214
rect 1788 3206 1796 3214
rect 1804 3206 1810 3214
rect 1810 3206 1812 3214
rect 4828 3206 4830 3214
rect 4830 3206 4836 3214
rect 4844 3206 4852 3214
rect 4860 3206 4866 3214
rect 4866 3206 4868 3214
rect 204 3176 212 3184
rect 4908 3196 4916 3204
rect 6316 3196 6324 3204
rect 4044 3176 4052 3184
rect 4940 3176 4948 3184
rect 6028 3176 6036 3184
rect 6604 3176 6612 3184
rect 2604 3156 2612 3164
rect 2764 3156 2772 3164
rect 4620 3156 4628 3164
rect 2732 3136 2740 3144
rect 2956 3116 2964 3124
rect 3724 3116 3732 3124
rect 4332 3136 4340 3144
rect 3884 3116 3892 3124
rect 4012 3116 4020 3124
rect 5356 3116 5364 3124
rect 5996 3116 6004 3124
rect 6060 3116 6068 3124
rect 6444 3136 6452 3144
rect 6604 3136 6612 3144
rect 6188 3116 6196 3124
rect 2028 3096 2036 3104
rect 2508 3096 2516 3104
rect 4076 3096 4084 3104
rect 4172 3096 4180 3104
rect 4268 3096 4276 3104
rect 2956 3056 2964 3064
rect 4492 3076 4500 3084
rect 5068 3076 5076 3084
rect 6348 3096 6356 3104
rect 5740 3076 5748 3084
rect 5644 3056 5652 3064
rect 5900 3056 5908 3064
rect 4524 3036 4532 3044
rect 5612 3036 5620 3044
rect 2988 3016 2996 3024
rect 4300 3016 4308 3024
rect 3308 3006 3310 3014
rect 3310 3006 3316 3014
rect 3324 3006 3332 3014
rect 3340 3006 3346 3014
rect 3346 3006 3348 3014
rect 4012 2996 4020 3004
rect 5804 2996 5812 3004
rect 1996 2976 2004 2984
rect 4076 2976 4084 2984
rect 2764 2956 2772 2964
rect 4620 2956 4628 2964
rect 5644 2956 5652 2964
rect 4332 2936 4340 2944
rect 4492 2936 4500 2944
rect 4716 2936 4724 2944
rect 5548 2936 5556 2944
rect 2476 2916 2484 2924
rect 4236 2916 4244 2924
rect 4748 2916 4756 2924
rect 5996 2916 6004 2924
rect 1516 2896 1524 2904
rect 4300 2896 4308 2904
rect 172 2876 180 2884
rect 2668 2876 2676 2884
rect 3820 2876 3828 2884
rect 4716 2876 4724 2884
rect 5932 2896 5940 2904
rect 12 2856 20 2864
rect 2028 2856 2036 2864
rect 4108 2856 4116 2864
rect 4172 2856 4180 2864
rect 2348 2836 2356 2844
rect 5548 2856 5556 2864
rect 5804 2856 5812 2864
rect 4620 2836 4628 2844
rect 4716 2836 4724 2844
rect 12 2816 20 2824
rect 1772 2806 1774 2814
rect 1774 2806 1780 2814
rect 1788 2806 1796 2814
rect 1804 2806 1810 2814
rect 1810 2806 1812 2814
rect 4828 2806 4830 2814
rect 4830 2806 4836 2814
rect 4844 2806 4852 2814
rect 4860 2806 4866 2814
rect 4866 2806 4868 2814
rect 2156 2796 2164 2804
rect 2700 2796 2708 2804
rect 2796 2796 2804 2804
rect 4492 2776 4500 2784
rect 2092 2756 2100 2764
rect 6124 2756 6132 2764
rect 3052 2736 3060 2744
rect 4268 2736 4276 2744
rect 876 2696 884 2704
rect 972 2696 980 2704
rect 2732 2696 2740 2704
rect 4748 2676 4756 2684
rect 6508 2716 6516 2724
rect 2732 2656 2740 2664
rect 4204 2656 4212 2664
rect 5996 2656 6004 2664
rect 2412 2636 2420 2644
rect 5868 2636 5876 2644
rect 6156 2636 6164 2644
rect 3308 2606 3310 2614
rect 3310 2606 3316 2614
rect 3324 2606 3332 2614
rect 3340 2606 3346 2614
rect 3346 2606 3348 2614
rect 908 2576 916 2584
rect 2412 2576 2420 2584
rect 4108 2576 4116 2584
rect 5004 2576 5012 2584
rect 2220 2556 2228 2564
rect 3916 2556 3924 2564
rect 5132 2556 5140 2564
rect 268 2536 276 2544
rect 4940 2536 4948 2544
rect 5004 2536 5012 2544
rect 3052 2516 3060 2524
rect 4588 2516 4596 2524
rect 5804 2516 5812 2524
rect 4108 2496 4116 2504
rect 4204 2496 4212 2504
rect 5580 2496 5588 2504
rect 5676 2496 5684 2504
rect 140 2476 148 2484
rect 2092 2476 2100 2484
rect 5484 2476 5492 2484
rect 172 2436 180 2444
rect 5132 2436 5140 2444
rect 6476 2436 6484 2444
rect 2700 2416 2708 2424
rect 1772 2406 1774 2414
rect 1774 2406 1780 2414
rect 1788 2406 1796 2414
rect 1804 2406 1810 2414
rect 1810 2406 1812 2414
rect 4828 2406 4830 2414
rect 4830 2406 4836 2414
rect 4844 2406 4852 2414
rect 4860 2406 4866 2414
rect 4866 2406 4868 2414
rect 4364 2396 4372 2404
rect 4748 2396 4756 2404
rect 2828 2376 2836 2384
rect 5900 2376 5908 2384
rect 5644 2356 5652 2364
rect 6124 2336 6132 2344
rect 12 2316 20 2324
rect 1420 2316 1428 2324
rect 2156 2316 2164 2324
rect 4940 2316 4948 2324
rect 1036 2296 1044 2304
rect 876 2276 884 2284
rect 908 2276 916 2284
rect 1516 2276 1524 2284
rect 4524 2276 4532 2284
rect 5068 2276 5076 2284
rect 3276 2256 3284 2264
rect 3532 2256 3540 2264
rect 876 2236 884 2244
rect 4588 2236 4596 2244
rect 6252 2236 6260 2244
rect 1740 2216 1748 2224
rect 4684 2216 4692 2224
rect 6220 2216 6228 2224
rect 3308 2206 3310 2214
rect 3310 2206 3316 2214
rect 3324 2206 3332 2214
rect 3340 2206 3346 2214
rect 3346 2206 3348 2214
rect 108 2196 116 2204
rect 652 2196 660 2204
rect 2380 2196 2388 2204
rect 2924 2196 2932 2204
rect 6348 2196 6356 2204
rect 6412 2196 6420 2204
rect 1452 2176 1460 2184
rect 5612 2176 5620 2184
rect 5836 2176 5844 2184
rect 2700 2156 2708 2164
rect 3404 2156 3412 2164
rect 140 2136 148 2144
rect 972 2136 980 2144
rect 1132 2136 1140 2144
rect 3276 2136 3284 2144
rect 6508 2136 6516 2144
rect 300 2116 308 2124
rect 3084 2116 3092 2124
rect 4588 2116 4596 2124
rect 4940 2076 4948 2084
rect 5964 2076 5972 2084
rect 6540 2076 6548 2084
rect 5068 2056 5076 2064
rect 6220 2016 6228 2024
rect 1772 2006 1774 2014
rect 1774 2006 1780 2014
rect 1788 2006 1796 2014
rect 1804 2006 1810 2014
rect 1810 2006 1812 2014
rect 4828 2006 4830 2014
rect 4830 2006 4836 2014
rect 4844 2006 4852 2014
rect 4860 2006 4866 2014
rect 4866 2006 4868 2014
rect 1516 1996 1524 2004
rect 4588 1996 4596 2004
rect 5516 1996 5524 2004
rect 6188 1996 6196 2004
rect 652 1976 660 1984
rect 2380 1976 2388 1984
rect 108 1956 116 1964
rect 2796 1956 2804 1964
rect 5356 1956 5364 1964
rect 5388 1956 5396 1964
rect 5740 1956 5748 1964
rect 332 1936 340 1944
rect 2220 1936 2228 1944
rect 1388 1916 1396 1924
rect 1420 1916 1428 1924
rect 1996 1916 2004 1924
rect 2348 1916 2356 1924
rect 5260 1896 5268 1904
rect 5356 1896 5364 1904
rect 5964 1896 5972 1904
rect 1196 1876 1204 1884
rect 2924 1876 2932 1884
rect 4940 1876 4948 1884
rect 5036 1876 5044 1884
rect 268 1856 276 1864
rect 908 1856 916 1864
rect 5196 1856 5204 1864
rect 5420 1856 5428 1864
rect 5900 1856 5908 1864
rect 844 1816 852 1824
rect 1292 1816 1300 1824
rect 3948 1816 3956 1824
rect 4524 1816 4532 1824
rect 5676 1816 5684 1824
rect 5772 1816 5780 1824
rect 6476 1816 6484 1824
rect 6508 1816 6516 1824
rect 3308 1806 3310 1814
rect 3310 1806 3316 1814
rect 3324 1806 3332 1814
rect 3340 1806 3346 1814
rect 3346 1806 3348 1814
rect 300 1796 308 1804
rect 5132 1796 5140 1804
rect 5804 1796 5812 1804
rect 716 1776 724 1784
rect 6348 1776 6356 1784
rect 3916 1756 3924 1764
rect 780 1736 788 1744
rect 1036 1736 1044 1744
rect 5036 1736 5044 1744
rect 5804 1736 5812 1744
rect 6284 1736 6292 1744
rect 6508 1736 6516 1744
rect 140 1716 148 1724
rect 5420 1696 5428 1704
rect 4684 1676 4692 1684
rect 6348 1676 6356 1684
rect 1484 1656 1492 1664
rect 5516 1656 5524 1664
rect 5580 1656 5588 1664
rect 6028 1656 6036 1664
rect 5100 1636 5108 1644
rect 5484 1636 5492 1644
rect 6476 1636 6484 1644
rect 6540 1636 6548 1644
rect 5964 1616 5972 1624
rect 1772 1606 1774 1614
rect 1774 1606 1780 1614
rect 1788 1606 1796 1614
rect 1804 1606 1810 1614
rect 1810 1606 1812 1614
rect 4828 1606 4830 1614
rect 4830 1606 4836 1614
rect 4844 1606 4852 1614
rect 4860 1606 4866 1614
rect 4866 1606 4868 1614
rect 1740 1596 1748 1604
rect 3532 1596 3540 1604
rect 4524 1596 4532 1604
rect 5676 1596 5684 1604
rect 5900 1596 5908 1604
rect 5996 1596 6004 1604
rect 6476 1596 6484 1604
rect 4940 1576 4948 1584
rect 6092 1556 6100 1564
rect 6284 1556 6292 1564
rect 172 1516 180 1524
rect 716 1516 724 1524
rect 1516 1516 1524 1524
rect 1932 1516 1940 1524
rect 3404 1536 3412 1544
rect 3948 1516 3956 1524
rect 4044 1516 4052 1524
rect 5452 1516 5460 1524
rect 44 1496 52 1504
rect 620 1496 628 1504
rect 108 1476 116 1484
rect 140 1476 148 1484
rect 332 1476 340 1484
rect 716 1476 724 1484
rect 844 1476 852 1484
rect 1132 1476 1140 1484
rect 2988 1476 2996 1484
rect 3660 1476 3668 1484
rect 4556 1476 4564 1484
rect 5324 1496 5332 1504
rect 5772 1496 5780 1504
rect 6060 1496 6068 1504
rect 6444 1496 6452 1504
rect 6156 1456 6164 1464
rect 5804 1436 5812 1444
rect 5836 1436 5844 1444
rect 5868 1436 5876 1444
rect 620 1416 628 1424
rect 1292 1416 1300 1424
rect 1580 1416 1588 1424
rect 1676 1416 1684 1424
rect 3308 1406 3310 1414
rect 3310 1406 3316 1414
rect 3324 1406 3332 1414
rect 3340 1406 3346 1414
rect 3346 1406 3348 1414
rect 5868 1396 5876 1404
rect 588 1376 596 1384
rect 4780 1376 4788 1384
rect 5452 1376 5460 1384
rect 780 1356 788 1364
rect 460 1336 468 1344
rect 1388 1356 1396 1364
rect 4940 1356 4948 1364
rect 5164 1356 5172 1364
rect 5516 1356 5524 1364
rect 5772 1356 5780 1364
rect 6156 1356 6164 1364
rect 1196 1336 1204 1344
rect 1452 1336 1460 1344
rect 2988 1336 2996 1344
rect 3820 1336 3828 1344
rect 1516 1316 1524 1324
rect 3564 1316 3572 1324
rect 3836 1316 3844 1324
rect 3884 1316 3892 1324
rect 4044 1336 4052 1344
rect 5036 1336 5044 1344
rect 5868 1336 5876 1344
rect 4940 1316 4948 1324
rect 5324 1316 5332 1324
rect 6348 1316 6356 1324
rect 908 1296 916 1304
rect 1484 1296 1492 1304
rect 1580 1296 1588 1304
rect 1676 1296 1684 1304
rect 1932 1296 1940 1304
rect 6124 1296 6132 1304
rect 1292 1276 1300 1284
rect 3660 1276 3668 1284
rect 6348 1276 6356 1284
rect 6412 1276 6420 1284
rect 3884 1256 3892 1264
rect 5644 1256 5652 1264
rect 6124 1256 6132 1264
rect 1580 1236 1588 1244
rect 5132 1236 5140 1244
rect 5932 1236 5940 1244
rect 6316 1236 6324 1244
rect 5068 1216 5076 1224
rect 1772 1206 1774 1214
rect 1774 1206 1780 1214
rect 1788 1206 1796 1214
rect 1804 1206 1810 1214
rect 1810 1206 1812 1214
rect 4828 1206 4830 1214
rect 4830 1206 4836 1214
rect 4844 1206 4852 1214
rect 4860 1206 4866 1214
rect 4866 1206 4868 1214
rect 1132 1196 1140 1204
rect 3244 1196 3252 1204
rect 4364 1196 4372 1204
rect 5708 1196 5716 1204
rect 44 1176 52 1184
rect 5420 1176 5428 1184
rect 1260 1156 1268 1164
rect 5260 1156 5268 1164
rect 44 1136 52 1144
rect 6284 1136 6292 1144
rect 6444 1136 6452 1144
rect 108 1116 116 1124
rect 2092 1116 2100 1124
rect 588 1096 596 1104
rect 1388 1096 1396 1104
rect 1708 1096 1716 1104
rect 5740 1096 5748 1104
rect 6156 1096 6164 1104
rect 6348 1096 6356 1104
rect 76 1076 84 1084
rect 172 1076 180 1084
rect 268 1076 276 1084
rect 1292 1076 1300 1084
rect 3916 1076 3924 1084
rect 2028 1056 2036 1064
rect 5772 1056 5780 1064
rect 5836 1056 5844 1064
rect 6156 1056 6164 1064
rect 6220 1056 6228 1064
rect 1292 1036 1300 1044
rect 1484 1036 1492 1044
rect 5260 1036 5268 1044
rect 6348 1036 6356 1044
rect 1068 1016 1076 1024
rect 3308 1006 3310 1014
rect 3310 1006 3316 1014
rect 3324 1006 3332 1014
rect 3340 1006 3346 1014
rect 3346 1006 3348 1014
rect 972 996 980 1004
rect 5068 996 5076 1004
rect 6188 1016 6196 1024
rect 6572 1016 6580 1024
rect 6156 996 6164 1004
rect 5996 976 6004 984
rect 6316 976 6324 984
rect 6284 956 6292 964
rect 6444 956 6452 964
rect 44 936 52 944
rect 6572 936 6580 944
rect 5964 916 5972 924
rect 6092 916 6100 924
rect 6604 916 6612 924
rect 6444 896 6452 904
rect 1708 876 1716 884
rect 76 856 84 864
rect 268 856 276 864
rect 3276 856 3284 864
rect 6060 876 6068 884
rect 5324 856 5332 864
rect 6444 856 6452 864
rect 3916 836 3924 844
rect 5100 836 5108 844
rect 5772 836 5780 844
rect 5964 836 5972 844
rect 5996 836 6004 844
rect 6572 836 6580 844
rect 6604 836 6612 844
rect 2700 816 2708 824
rect 3564 816 3572 824
rect 1772 806 1774 814
rect 1774 806 1780 814
rect 1788 806 1796 814
rect 1804 806 1810 814
rect 1810 806 1812 814
rect 4828 806 4830 814
rect 4830 806 4836 814
rect 4844 806 4852 814
rect 4860 806 4866 814
rect 4866 806 4868 814
rect 364 796 372 804
rect 716 796 724 804
rect 972 796 980 804
rect 1196 796 1204 804
rect 2540 796 2548 804
rect 2540 756 2548 764
rect 5420 756 5428 764
rect 812 736 820 744
rect 4556 736 4564 744
rect 4620 736 4628 744
rect 6060 736 6068 744
rect 460 716 468 724
rect 1068 716 1076 724
rect 1292 716 1300 724
rect 5676 716 5684 724
rect 108 696 116 704
rect 1260 696 1268 704
rect 5036 696 5044 704
rect 6252 696 6260 704
rect 12 676 20 684
rect 652 676 660 684
rect 2092 676 2100 684
rect 2700 676 2708 684
rect 2540 656 2548 664
rect 3500 656 3508 664
rect 6252 656 6260 664
rect 2060 616 2068 624
rect 2092 616 2100 624
rect 4620 616 4628 624
rect 3308 606 3310 614
rect 3310 606 3316 614
rect 3324 606 3332 614
rect 3340 606 3346 614
rect 3346 606 3348 614
rect 684 596 692 604
rect 2028 596 2036 604
rect 4524 596 4532 604
rect 5388 596 5396 604
rect 5612 596 5620 604
rect 6572 596 6580 604
rect 460 556 468 564
rect 524 556 532 564
rect 3276 556 3284 564
rect 1484 536 1492 544
rect 1132 516 1140 524
rect 1196 516 1204 524
rect 5356 576 5364 584
rect 5676 576 5684 584
rect 4556 556 4564 564
rect 4588 556 4596 564
rect 4780 556 4788 564
rect 5164 556 5172 564
rect 5324 556 5332 564
rect 6252 536 6260 544
rect 12 496 20 504
rect 652 496 660 504
rect 2380 496 2388 504
rect 3500 496 3508 504
rect 4588 516 4596 524
rect 5196 516 5204 524
rect 3884 496 3892 504
rect 812 476 820 484
rect 3916 476 3924 484
rect 6572 476 6580 484
rect 2092 456 2100 464
rect 6188 456 6196 464
rect 588 436 596 444
rect 1676 436 1684 444
rect 1868 436 1876 444
rect 5900 436 5908 444
rect 6572 436 6580 444
rect 684 416 692 424
rect 6636 416 6644 424
rect 1772 406 1774 414
rect 1774 406 1780 414
rect 1788 406 1796 414
rect 1804 406 1810 414
rect 1810 406 1812 414
rect 4828 406 4830 414
rect 4830 406 4836 414
rect 4844 406 4852 414
rect 4860 406 4866 414
rect 4866 406 4868 414
rect 876 396 884 404
rect 1836 396 1844 404
rect 2028 396 2036 404
rect 2060 396 2068 404
rect 364 376 372 384
rect 524 376 532 384
rect 812 376 820 384
rect 2476 376 2484 384
rect 3404 376 3412 384
rect 6444 376 6452 384
rect 780 356 788 364
rect 364 336 372 344
rect 1484 336 1492 344
rect 3436 336 3444 344
rect 524 316 532 324
rect 556 316 564 324
rect 668 316 676 324
rect 3148 316 3156 324
rect 3820 316 3828 324
rect 940 296 948 304
rect 5324 316 5332 324
rect 6252 316 6260 324
rect 2476 296 2484 304
rect 2572 296 2580 304
rect 364 276 372 284
rect 780 276 788 284
rect 876 276 884 284
rect 1260 276 1268 284
rect 3132 276 3140 284
rect 108 236 116 244
rect 1836 256 1844 264
rect 1868 256 1876 264
rect 2604 256 2612 264
rect 3052 256 3060 264
rect 6412 276 6420 284
rect 6604 276 6612 284
rect 6636 276 6644 284
rect 4268 256 4276 264
rect 2380 236 2388 244
rect 6252 236 6260 244
rect 2044 196 2052 204
rect 3052 216 3060 224
rect 3244 216 3252 224
rect 3372 216 3380 224
rect 6348 216 6356 224
rect 3308 206 3310 214
rect 3310 206 3316 214
rect 3324 206 3332 214
rect 3340 206 3346 214
rect 3346 206 3348 214
rect 3084 196 3092 204
rect 3404 196 3412 204
rect 3820 196 3828 204
rect 5932 196 5940 204
rect 6156 196 6164 204
rect 492 176 500 184
rect 2924 176 2932 184
rect 3276 176 3284 184
rect 5964 176 5972 184
rect 6604 176 6612 184
rect 844 156 852 164
rect 1260 156 1268 164
rect 2876 156 2884 164
rect 2988 156 2996 164
rect 3020 156 3028 164
rect 6028 156 6036 164
rect 6508 156 6516 164
rect 716 136 724 144
rect 780 136 788 144
rect 940 136 948 144
rect 1580 136 1588 144
rect 3436 136 3444 144
rect 1516 116 1524 124
rect 1900 116 1908 124
rect 4524 116 4532 124
rect 6124 136 6132 144
rect 6284 136 6292 144
rect 6412 136 6420 144
rect 6476 136 6484 144
rect 5324 116 5332 124
rect 6380 116 6388 124
rect 620 96 628 104
rect 6316 96 6324 104
rect 6540 96 6548 104
rect 588 76 596 84
rect 940 76 948 84
rect 1948 76 1956 84
rect 2492 76 2500 84
rect 3372 76 3380 84
rect 6060 76 6068 84
rect 6188 76 6196 84
rect 6636 76 6644 84
rect 1676 56 1684 64
rect 2476 56 2484 64
rect 2860 56 2868 64
rect 2924 56 2932 64
rect 2796 36 2804 44
rect 6604 56 6612 64
rect 6412 36 6420 44
rect 3020 16 3028 24
rect 3276 16 3284 24
rect 6572 16 6580 24
rect 1772 6 1774 14
rect 1774 6 1780 14
rect 1788 6 1796 14
rect 1804 6 1810 14
rect 1810 6 1812 14
rect 4828 6 4830 14
rect 4830 6 4836 14
rect 4844 6 4852 14
rect 4860 6 4866 14
rect 4866 6 4868 14
<< metal4 >>
rect 1768 4814 1816 4840
rect 1768 4806 1772 4814
rect 1780 4806 1788 4814
rect 1796 4806 1804 4814
rect 1812 4806 1816 4814
rect 938 4754 1078 4766
rect 10 4744 22 4746
rect 10 4736 12 4744
rect 20 4736 22 4744
rect 10 4704 22 4736
rect 938 4744 950 4754
rect 938 4736 940 4744
rect 948 4736 950 4744
rect 938 4734 950 4736
rect 1066 4726 1078 4754
rect 1066 4714 1206 4726
rect 10 4696 12 4704
rect 20 4696 22 4704
rect 10 4694 22 4696
rect 1002 4704 1014 4706
rect 1002 4696 1004 4704
rect 1012 4696 1014 4704
rect 1002 4686 1014 4696
rect 890 4684 1014 4686
rect 890 4676 892 4684
rect 900 4676 1014 4684
rect 890 4674 1014 4676
rect 1034 4704 1046 4706
rect 1034 4696 1036 4704
rect 1044 4696 1046 4704
rect 1034 4686 1046 4696
rect 1194 4704 1206 4714
rect 1194 4696 1196 4704
rect 1204 4696 1206 4704
rect 1194 4694 1206 4696
rect 1418 4714 1526 4726
rect 1034 4684 1126 4686
rect 1034 4676 1116 4684
rect 1124 4676 1126 4684
rect 1034 4674 1126 4676
rect 74 4664 86 4666
rect 74 4656 76 4664
rect 84 4656 86 4664
rect 10 4504 22 4506
rect 10 4496 12 4504
rect 20 4496 22 4504
rect 10 4384 22 4496
rect 10 4376 12 4384
rect 20 4376 22 4384
rect 10 4374 22 4376
rect 42 4364 54 4366
rect 42 4356 44 4364
rect 52 4356 54 4364
rect 10 4264 22 4266
rect 10 4256 12 4264
rect 20 4256 22 4264
rect 10 4104 22 4256
rect 10 4096 12 4104
rect 20 4096 22 4104
rect 10 4094 22 4096
rect 10 3344 22 3346
rect 10 3336 12 3344
rect 20 3336 22 3344
rect 10 2864 22 3336
rect 42 3344 54 4356
rect 74 4184 86 4656
rect 1290 4644 1302 4646
rect 1290 4636 1292 4644
rect 1300 4636 1302 4644
rect 1290 4584 1302 4636
rect 1418 4644 1430 4714
rect 1418 4636 1420 4644
rect 1428 4636 1430 4644
rect 1418 4634 1430 4636
rect 1514 4646 1526 4714
rect 1514 4644 1606 4646
rect 1514 4636 1596 4644
rect 1604 4636 1606 4644
rect 1514 4634 1606 4636
rect 1290 4576 1292 4584
rect 1300 4576 1302 4584
rect 1290 4574 1302 4576
rect 1546 4604 1558 4606
rect 1546 4596 1548 4604
rect 1556 4596 1558 4604
rect 1546 4564 1558 4596
rect 1546 4556 1548 4564
rect 1556 4556 1558 4564
rect 1546 4554 1558 4556
rect 394 4524 406 4526
rect 394 4516 396 4524
rect 404 4516 406 4524
rect 362 4504 374 4506
rect 362 4496 364 4504
rect 372 4496 374 4504
rect 362 4486 374 4496
rect 266 4474 374 4486
rect 266 4464 278 4474
rect 266 4456 268 4464
rect 276 4456 278 4464
rect 266 4454 278 4456
rect 394 4404 406 4516
rect 394 4396 396 4404
rect 404 4396 406 4404
rect 394 4394 406 4396
rect 1322 4464 1334 4466
rect 1322 4456 1324 4464
rect 1332 4456 1334 4464
rect 1322 4404 1334 4456
rect 1322 4396 1324 4404
rect 1332 4396 1334 4404
rect 1322 4394 1334 4396
rect 1768 4414 1816 4806
rect 2570 4804 2582 4806
rect 2570 4796 2572 4804
rect 2580 4796 2582 4804
rect 2154 4754 2326 4766
rect 1850 4724 1878 4726
rect 1850 4716 1852 4724
rect 1860 4716 1878 4724
rect 1850 4714 1878 4716
rect 1866 4686 1878 4714
rect 1994 4724 2006 4726
rect 1994 4716 1996 4724
rect 2004 4716 2006 4724
rect 1994 4686 2006 4716
rect 2154 4724 2166 4754
rect 2154 4716 2156 4724
rect 2164 4716 2166 4724
rect 2154 4714 2166 4716
rect 2186 4724 2198 4726
rect 2186 4716 2188 4724
rect 2196 4716 2198 4724
rect 1866 4684 1958 4686
rect 1866 4676 1948 4684
rect 1956 4676 1958 4684
rect 1866 4674 1958 4676
rect 1978 4684 2006 4686
rect 1978 4676 1980 4684
rect 1988 4676 2006 4684
rect 1978 4674 2006 4676
rect 1768 4406 1772 4414
rect 1780 4406 1788 4414
rect 1796 4406 1804 4414
rect 1812 4406 1816 4414
rect 234 4344 246 4346
rect 234 4336 236 4344
rect 244 4336 246 4344
rect 74 4176 76 4184
rect 84 4176 86 4184
rect 74 4174 86 4176
rect 138 4304 150 4306
rect 138 4296 140 4304
rect 148 4296 150 4304
rect 138 4084 150 4296
rect 138 4076 140 4084
rect 148 4076 150 4084
rect 138 4074 150 4076
rect 234 4084 246 4336
rect 714 4304 726 4306
rect 714 4296 716 4304
rect 724 4296 726 4304
rect 330 4264 342 4266
rect 330 4256 332 4264
rect 340 4256 342 4264
rect 330 4246 342 4256
rect 266 4244 342 4246
rect 266 4236 268 4244
rect 276 4236 342 4244
rect 266 4234 342 4236
rect 426 4244 438 4246
rect 426 4236 428 4244
rect 436 4236 438 4244
rect 234 4076 236 4084
rect 244 4076 246 4084
rect 234 4074 246 4076
rect 202 3924 230 3926
rect 202 3916 220 3924
rect 228 3916 230 3924
rect 202 3914 230 3916
rect 202 3886 214 3914
rect 186 3884 214 3886
rect 186 3876 188 3884
rect 196 3876 214 3884
rect 186 3874 214 3876
rect 42 3336 44 3344
rect 52 3336 54 3344
rect 42 3334 54 3336
rect 202 3644 214 3646
rect 202 3636 204 3644
rect 212 3636 214 3644
rect 202 3184 214 3636
rect 426 3484 438 4236
rect 714 3744 726 4296
rect 778 4264 790 4266
rect 778 4256 780 4264
rect 788 4256 790 4264
rect 778 4104 790 4256
rect 778 4096 780 4104
rect 788 4096 790 4104
rect 778 4094 790 4096
rect 1066 4224 1078 4226
rect 1066 4216 1068 4224
rect 1076 4216 1078 4224
rect 714 3736 716 3744
rect 724 3736 726 3744
rect 714 3734 726 3736
rect 426 3476 428 3484
rect 436 3476 438 3484
rect 426 3474 438 3476
rect 1066 3324 1078 4216
rect 1768 4014 1816 4406
rect 2186 4264 2198 4716
rect 2250 4724 2262 4726
rect 2250 4716 2252 4724
rect 2260 4716 2262 4724
rect 2250 4584 2262 4716
rect 2314 4724 2326 4754
rect 2314 4716 2316 4724
rect 2324 4716 2326 4724
rect 2314 4714 2326 4716
rect 2570 4724 2582 4796
rect 3146 4764 3158 4766
rect 3146 4756 3148 4764
rect 3156 4756 3158 4764
rect 2570 4716 2572 4724
rect 2580 4716 2582 4724
rect 2570 4714 2582 4716
rect 2730 4724 2742 4726
rect 2730 4716 2732 4724
rect 2740 4716 2742 4724
rect 2730 4684 2742 4716
rect 2730 4676 2732 4684
rect 2740 4676 2742 4684
rect 2730 4674 2742 4676
rect 2986 4724 2998 4726
rect 2986 4716 2988 4724
rect 2996 4716 2998 4724
rect 2986 4684 2998 4716
rect 2986 4676 2988 4684
rect 2996 4676 2998 4684
rect 2986 4674 2998 4676
rect 3018 4724 3030 4726
rect 3018 4716 3020 4724
rect 3028 4716 3030 4724
rect 2250 4576 2252 4584
rect 2260 4576 2262 4584
rect 2250 4574 2262 4576
rect 2634 4664 2646 4666
rect 2634 4656 2636 4664
rect 2644 4656 2646 4664
rect 2346 4484 2358 4486
rect 2346 4476 2348 4484
rect 2356 4476 2358 4484
rect 2186 4256 2188 4264
rect 2196 4256 2198 4264
rect 2186 4254 2198 4256
rect 2218 4304 2230 4306
rect 2218 4296 2220 4304
rect 2228 4296 2230 4304
rect 2218 4184 2230 4296
rect 2218 4176 2220 4184
rect 2228 4176 2230 4184
rect 2218 4174 2230 4176
rect 2346 4104 2358 4476
rect 2634 4424 2646 4656
rect 2634 4416 2636 4424
rect 2644 4416 2646 4424
rect 2634 4414 2646 4416
rect 2666 4544 2678 4546
rect 2666 4536 2668 4544
rect 2676 4536 2678 4544
rect 2346 4096 2348 4104
rect 2356 4096 2358 4104
rect 2346 4094 2358 4096
rect 1768 4006 1772 4014
rect 1780 4006 1788 4014
rect 1796 4006 1804 4014
rect 1812 4006 1816 4014
rect 1768 3614 1816 4006
rect 2506 4044 2518 4046
rect 2506 4036 2508 4044
rect 2516 4036 2518 4044
rect 2058 3844 2070 3846
rect 2058 3836 2060 3844
rect 2068 3836 2070 3844
rect 1768 3606 1772 3614
rect 1780 3606 1788 3614
rect 1796 3606 1804 3614
rect 1812 3606 1816 3614
rect 1066 3316 1068 3324
rect 1076 3316 1078 3324
rect 1066 3314 1078 3316
rect 1738 3344 1750 3346
rect 1738 3336 1740 3344
rect 1748 3336 1750 3344
rect 202 3176 204 3184
rect 212 3176 214 3184
rect 202 3174 214 3176
rect 874 3244 886 3246
rect 874 3236 876 3244
rect 884 3236 886 3244
rect 10 2856 12 2864
rect 20 2856 22 2864
rect 10 2854 22 2856
rect 170 2884 182 2886
rect 170 2876 172 2884
rect 180 2876 182 2884
rect 10 2824 22 2826
rect 10 2816 12 2824
rect 20 2816 22 2824
rect 10 2324 22 2816
rect 10 2316 12 2324
rect 20 2316 22 2324
rect 10 2314 22 2316
rect 138 2484 150 2486
rect 138 2476 140 2484
rect 148 2476 150 2484
rect 106 2204 118 2206
rect 106 2196 108 2204
rect 116 2196 118 2204
rect 106 1964 118 2196
rect 138 2144 150 2476
rect 170 2444 182 2876
rect 874 2704 886 3236
rect 1738 3224 1750 3336
rect 1738 3216 1740 3224
rect 1748 3216 1750 3224
rect 1738 3214 1750 3216
rect 1768 3214 1816 3606
rect 1768 3206 1772 3214
rect 1780 3206 1788 3214
rect 1796 3206 1804 3214
rect 1812 3206 1816 3214
rect 1514 2904 1526 2906
rect 1514 2896 1516 2904
rect 1524 2896 1526 2904
rect 874 2696 876 2704
rect 884 2696 886 2704
rect 874 2694 886 2696
rect 970 2704 982 2706
rect 970 2696 972 2704
rect 980 2696 982 2704
rect 906 2584 918 2586
rect 906 2576 908 2584
rect 916 2576 918 2584
rect 170 2436 172 2444
rect 180 2436 182 2444
rect 170 2434 182 2436
rect 266 2544 278 2546
rect 266 2536 268 2544
rect 276 2536 278 2544
rect 138 2136 140 2144
rect 148 2136 150 2144
rect 138 2134 150 2136
rect 106 1956 108 1964
rect 116 1956 118 1964
rect 106 1954 118 1956
rect 266 1864 278 2536
rect 874 2284 886 2286
rect 874 2276 876 2284
rect 884 2276 886 2284
rect 874 2244 886 2276
rect 906 2284 918 2576
rect 906 2276 908 2284
rect 916 2276 918 2284
rect 906 2274 918 2276
rect 874 2236 876 2244
rect 884 2236 886 2244
rect 874 2234 886 2236
rect 650 2204 662 2206
rect 650 2196 652 2204
rect 660 2196 662 2204
rect 266 1856 268 1864
rect 276 1856 278 1864
rect 266 1854 278 1856
rect 298 2124 310 2126
rect 298 2116 300 2124
rect 308 2116 310 2124
rect 298 1804 310 2116
rect 650 1984 662 2196
rect 970 2144 982 2696
rect 1418 2324 1430 2326
rect 1418 2316 1420 2324
rect 1428 2316 1430 2324
rect 970 2136 972 2144
rect 980 2136 982 2144
rect 970 2134 982 2136
rect 1034 2304 1046 2306
rect 1034 2296 1036 2304
rect 1044 2296 1046 2304
rect 650 1976 652 1984
rect 660 1976 662 1984
rect 650 1974 662 1976
rect 298 1796 300 1804
rect 308 1796 310 1804
rect 298 1794 310 1796
rect 330 1944 342 1946
rect 330 1936 332 1944
rect 340 1936 342 1944
rect 138 1724 150 1726
rect 138 1716 140 1724
rect 148 1716 150 1724
rect 42 1504 54 1506
rect 42 1496 44 1504
rect 52 1496 54 1504
rect 42 1184 54 1496
rect 42 1176 44 1184
rect 52 1176 54 1184
rect 42 1174 54 1176
rect 106 1484 118 1486
rect 106 1476 108 1484
rect 116 1476 118 1484
rect 42 1144 54 1146
rect 42 1136 44 1144
rect 52 1136 54 1144
rect 42 944 54 1136
rect 106 1124 118 1476
rect 138 1484 150 1716
rect 138 1476 140 1484
rect 148 1476 150 1484
rect 138 1474 150 1476
rect 170 1524 182 1526
rect 170 1516 172 1524
rect 180 1516 182 1524
rect 106 1116 108 1124
rect 116 1116 118 1124
rect 106 1114 118 1116
rect 42 936 44 944
rect 52 936 54 944
rect 42 934 54 936
rect 74 1084 86 1086
rect 74 1076 76 1084
rect 84 1076 86 1084
rect 74 864 86 1076
rect 170 1084 182 1516
rect 330 1484 342 1936
rect 906 1864 918 1866
rect 906 1856 908 1864
rect 916 1856 918 1864
rect 842 1824 854 1826
rect 842 1816 844 1824
rect 852 1816 854 1824
rect 714 1784 726 1786
rect 714 1776 716 1784
rect 724 1776 726 1784
rect 714 1524 726 1776
rect 714 1516 716 1524
rect 724 1516 726 1524
rect 714 1514 726 1516
rect 778 1744 790 1746
rect 778 1736 780 1744
rect 788 1736 790 1744
rect 330 1476 332 1484
rect 340 1476 342 1484
rect 330 1474 342 1476
rect 618 1504 630 1506
rect 618 1496 620 1504
rect 628 1496 630 1504
rect 618 1424 630 1496
rect 618 1416 620 1424
rect 628 1416 630 1424
rect 618 1414 630 1416
rect 714 1484 726 1486
rect 714 1476 716 1484
rect 724 1476 726 1484
rect 586 1384 598 1386
rect 586 1376 588 1384
rect 596 1376 598 1384
rect 458 1344 470 1346
rect 458 1336 460 1344
rect 468 1336 470 1344
rect 170 1076 172 1084
rect 180 1076 182 1084
rect 170 1074 182 1076
rect 266 1084 278 1086
rect 266 1076 268 1084
rect 276 1076 278 1084
rect 74 856 76 864
rect 84 856 86 864
rect 74 854 86 856
rect 266 864 278 1076
rect 266 856 268 864
rect 276 856 278 864
rect 266 854 278 856
rect 362 804 374 806
rect 362 796 364 804
rect 372 796 374 804
rect 106 704 118 706
rect 106 696 108 704
rect 116 696 118 704
rect 10 684 22 686
rect 10 676 12 684
rect 20 676 22 684
rect 10 504 22 676
rect 10 496 12 504
rect 20 496 22 504
rect 10 494 22 496
rect 106 244 118 696
rect 362 384 374 796
rect 458 724 470 1336
rect 586 1104 598 1376
rect 586 1096 588 1104
rect 596 1096 598 1104
rect 586 1094 598 1096
rect 714 804 726 1476
rect 778 1364 790 1736
rect 842 1484 854 1816
rect 842 1476 844 1484
rect 852 1476 854 1484
rect 842 1474 854 1476
rect 778 1356 780 1364
rect 788 1356 790 1364
rect 778 1354 790 1356
rect 906 1304 918 1856
rect 1034 1744 1046 2296
rect 1034 1736 1036 1744
rect 1044 1736 1046 1744
rect 1034 1734 1046 1736
rect 1130 2144 1142 2146
rect 1130 2136 1132 2144
rect 1140 2136 1142 2144
rect 1130 1484 1142 2136
rect 1386 1924 1398 1926
rect 1386 1916 1388 1924
rect 1396 1916 1398 1924
rect 1130 1476 1132 1484
rect 1140 1476 1142 1484
rect 1130 1474 1142 1476
rect 1194 1884 1206 1886
rect 1194 1876 1196 1884
rect 1204 1876 1206 1884
rect 1194 1344 1206 1876
rect 1290 1824 1302 1826
rect 1290 1816 1292 1824
rect 1300 1816 1302 1824
rect 1290 1424 1302 1816
rect 1290 1416 1292 1424
rect 1300 1416 1302 1424
rect 1290 1414 1302 1416
rect 1194 1336 1196 1344
rect 1204 1336 1206 1344
rect 1194 1334 1206 1336
rect 1386 1364 1398 1916
rect 1418 1924 1430 2316
rect 1514 2284 1526 2896
rect 1514 2276 1516 2284
rect 1524 2276 1526 2284
rect 1418 1916 1420 1924
rect 1428 1916 1430 1924
rect 1418 1914 1430 1916
rect 1450 2184 1462 2186
rect 1450 2176 1452 2184
rect 1460 2176 1462 2184
rect 1386 1356 1388 1364
rect 1396 1356 1398 1364
rect 906 1296 908 1304
rect 916 1296 918 1304
rect 906 1294 918 1296
rect 1290 1284 1302 1286
rect 1290 1276 1292 1284
rect 1300 1276 1302 1284
rect 1130 1204 1142 1206
rect 1130 1196 1132 1204
rect 1140 1196 1142 1204
rect 1066 1024 1078 1026
rect 1066 1016 1068 1024
rect 1076 1016 1078 1024
rect 714 796 716 804
rect 724 796 726 804
rect 714 794 726 796
rect 970 1004 982 1006
rect 970 996 972 1004
rect 980 996 982 1004
rect 970 804 982 996
rect 970 796 972 804
rect 980 796 982 804
rect 970 794 982 796
rect 458 716 460 724
rect 468 716 470 724
rect 458 564 470 716
rect 810 744 822 746
rect 810 736 812 744
rect 820 736 822 744
rect 650 684 662 686
rect 650 676 652 684
rect 660 676 662 684
rect 458 556 460 564
rect 468 556 470 564
rect 458 554 470 556
rect 522 564 534 566
rect 522 556 524 564
rect 532 556 534 564
rect 362 376 364 384
rect 372 376 374 384
rect 362 374 374 376
rect 522 384 534 556
rect 650 504 662 676
rect 650 496 652 504
rect 660 496 662 504
rect 650 494 662 496
rect 682 604 694 606
rect 682 596 684 604
rect 692 596 694 604
rect 522 376 524 384
rect 532 376 534 384
rect 362 344 374 346
rect 362 336 364 344
rect 372 336 374 344
rect 362 284 374 336
rect 522 324 534 376
rect 586 444 598 446
rect 586 436 588 444
rect 596 436 598 444
rect 522 316 524 324
rect 532 316 534 324
rect 522 314 534 316
rect 554 324 566 326
rect 554 316 556 324
rect 564 316 566 324
rect 554 286 566 316
rect 362 276 364 284
rect 372 276 374 284
rect 362 274 374 276
rect 490 274 566 286
rect 106 236 108 244
rect 116 236 118 244
rect 106 234 118 236
rect 490 184 502 274
rect 490 176 492 184
rect 500 176 502 184
rect 490 174 502 176
rect 586 84 598 436
rect 682 424 694 596
rect 810 484 822 736
rect 1066 724 1078 1016
rect 1066 716 1068 724
rect 1076 716 1078 724
rect 1066 714 1078 716
rect 1130 524 1142 1196
rect 1258 1164 1270 1166
rect 1258 1156 1260 1164
rect 1268 1156 1270 1164
rect 1130 516 1132 524
rect 1140 516 1142 524
rect 1130 514 1142 516
rect 1194 804 1206 806
rect 1194 796 1196 804
rect 1204 796 1206 804
rect 1194 524 1206 796
rect 1258 704 1270 1156
rect 1290 1084 1302 1276
rect 1386 1104 1398 1356
rect 1450 1344 1462 2176
rect 1514 2004 1526 2276
rect 1768 2814 1816 3206
rect 2026 3664 2038 3666
rect 2026 3656 2028 3664
rect 2036 3656 2038 3664
rect 2026 3564 2038 3656
rect 2026 3556 2028 3564
rect 2036 3556 2038 3564
rect 2026 3104 2038 3556
rect 2058 3304 2070 3836
rect 2314 3744 2326 3746
rect 2314 3736 2316 3744
rect 2324 3736 2326 3744
rect 2314 3404 2326 3736
rect 2314 3396 2316 3404
rect 2324 3396 2326 3404
rect 2314 3394 2326 3396
rect 2058 3296 2060 3304
rect 2068 3296 2070 3304
rect 2058 3294 2070 3296
rect 2474 3304 2486 3306
rect 2474 3296 2476 3304
rect 2484 3296 2486 3304
rect 2026 3096 2028 3104
rect 2036 3096 2038 3104
rect 1768 2806 1772 2814
rect 1780 2806 1788 2814
rect 1796 2806 1804 2814
rect 1812 2806 1816 2814
rect 1768 2414 1816 2806
rect 1768 2406 1772 2414
rect 1780 2406 1788 2414
rect 1796 2406 1804 2414
rect 1812 2406 1816 2414
rect 1514 1996 1516 2004
rect 1524 1996 1526 2004
rect 1514 1994 1526 1996
rect 1738 2224 1750 2226
rect 1738 2216 1740 2224
rect 1748 2216 1750 2224
rect 1450 1336 1452 1344
rect 1460 1336 1462 1344
rect 1450 1334 1462 1336
rect 1482 1664 1494 1666
rect 1482 1656 1484 1664
rect 1492 1656 1494 1664
rect 1482 1304 1494 1656
rect 1738 1604 1750 2216
rect 1738 1596 1740 1604
rect 1748 1596 1750 1604
rect 1738 1594 1750 1596
rect 1768 2014 1816 2406
rect 1768 2006 1772 2014
rect 1780 2006 1788 2014
rect 1796 2006 1804 2014
rect 1812 2006 1816 2014
rect 1768 1614 1816 2006
rect 1994 2984 2006 2986
rect 1994 2976 1996 2984
rect 2004 2976 2006 2984
rect 1994 1924 2006 2976
rect 2026 2864 2038 3096
rect 2474 2924 2486 3296
rect 2506 3104 2518 4036
rect 2666 4004 2678 4536
rect 3018 4504 3030 4716
rect 3146 4604 3158 4756
rect 3146 4596 3148 4604
rect 3156 4596 3158 4604
rect 3146 4594 3158 4596
rect 3304 4614 3352 4840
rect 4824 4814 4872 4840
rect 4824 4806 4828 4814
rect 4836 4806 4844 4814
rect 4852 4806 4860 4814
rect 4868 4806 4872 4814
rect 3304 4606 3308 4614
rect 3316 4606 3324 4614
rect 3332 4606 3340 4614
rect 3348 4606 3352 4614
rect 3018 4496 3020 4504
rect 3028 4496 3030 4504
rect 3018 4494 3030 4496
rect 2858 4344 2870 4346
rect 2858 4336 2860 4344
rect 2868 4336 2870 4344
rect 2666 3996 2668 4004
rect 2676 3996 2678 4004
rect 2602 3824 2614 3826
rect 2602 3816 2604 3824
rect 2612 3816 2614 3824
rect 2602 3164 2614 3816
rect 2602 3156 2604 3164
rect 2612 3156 2614 3164
rect 2602 3154 2614 3156
rect 2666 3304 2678 3996
rect 2666 3296 2668 3304
rect 2676 3296 2678 3304
rect 2506 3096 2508 3104
rect 2516 3096 2518 3104
rect 2506 3094 2518 3096
rect 2474 2916 2476 2924
rect 2484 2916 2486 2924
rect 2474 2914 2486 2916
rect 2666 2884 2678 3296
rect 2666 2876 2668 2884
rect 2676 2876 2678 2884
rect 2666 2874 2678 2876
rect 2698 4304 2710 4306
rect 2698 4296 2700 4304
rect 2708 4296 2710 4304
rect 2026 2856 2028 2864
rect 2036 2856 2038 2864
rect 2026 2854 2038 2856
rect 2346 2844 2358 2846
rect 2346 2836 2348 2844
rect 2356 2836 2358 2844
rect 2154 2804 2166 2806
rect 2154 2796 2156 2804
rect 2164 2796 2166 2804
rect 2090 2764 2102 2766
rect 2090 2756 2092 2764
rect 2100 2756 2102 2764
rect 2090 2484 2102 2756
rect 2090 2476 2092 2484
rect 2100 2476 2102 2484
rect 2090 2474 2102 2476
rect 2154 2324 2166 2796
rect 2154 2316 2156 2324
rect 2164 2316 2166 2324
rect 2154 2314 2166 2316
rect 2218 2564 2230 2566
rect 2218 2556 2220 2564
rect 2228 2556 2230 2564
rect 2218 1944 2230 2556
rect 2218 1936 2220 1944
rect 2228 1936 2230 1944
rect 2218 1934 2230 1936
rect 1994 1916 1996 1924
rect 2004 1916 2006 1924
rect 1994 1914 2006 1916
rect 2346 1924 2358 2836
rect 2698 2804 2710 4296
rect 2858 4164 2870 4336
rect 3210 4324 3222 4326
rect 3210 4316 3212 4324
rect 3220 4316 3222 4324
rect 2858 4156 2860 4164
rect 2868 4156 2870 4164
rect 2858 4154 2870 4156
rect 2986 4184 2998 4186
rect 2986 4176 2988 4184
rect 2996 4176 2998 4184
rect 2858 4004 2870 4006
rect 2858 3996 2860 4004
rect 2868 3996 2870 4004
rect 2858 3704 2870 3996
rect 2858 3696 2860 3704
rect 2868 3696 2870 3704
rect 2858 3694 2870 3696
rect 2890 3784 2902 3786
rect 2890 3776 2892 3784
rect 2900 3776 2902 3784
rect 2730 3584 2742 3586
rect 2730 3576 2732 3584
rect 2740 3576 2742 3584
rect 2730 3144 2742 3576
rect 2890 3544 2902 3776
rect 2890 3536 2892 3544
rect 2900 3536 2902 3544
rect 2890 3534 2902 3536
rect 2826 3464 2838 3466
rect 2826 3456 2828 3464
rect 2836 3456 2838 3464
rect 2730 3136 2732 3144
rect 2740 3136 2742 3144
rect 2730 3134 2742 3136
rect 2762 3164 2774 3166
rect 2762 3156 2764 3164
rect 2772 3156 2774 3164
rect 2762 2964 2774 3156
rect 2762 2956 2764 2964
rect 2772 2956 2774 2964
rect 2762 2954 2774 2956
rect 2698 2796 2700 2804
rect 2708 2796 2710 2804
rect 2698 2794 2710 2796
rect 2794 2804 2806 2806
rect 2794 2796 2796 2804
rect 2804 2796 2806 2804
rect 2730 2704 2742 2706
rect 2730 2696 2732 2704
rect 2740 2696 2742 2704
rect 2730 2664 2742 2696
rect 2730 2656 2732 2664
rect 2740 2656 2742 2664
rect 2730 2654 2742 2656
rect 2410 2644 2422 2646
rect 2410 2636 2412 2644
rect 2420 2636 2422 2644
rect 2410 2584 2422 2636
rect 2410 2576 2412 2584
rect 2420 2576 2422 2584
rect 2410 2574 2422 2576
rect 2698 2424 2710 2426
rect 2698 2416 2700 2424
rect 2708 2416 2710 2424
rect 2378 2204 2390 2206
rect 2378 2196 2380 2204
rect 2388 2196 2390 2204
rect 2378 1984 2390 2196
rect 2698 2164 2710 2416
rect 2698 2156 2700 2164
rect 2708 2156 2710 2164
rect 2698 2154 2710 2156
rect 2378 1976 2380 1984
rect 2388 1976 2390 1984
rect 2378 1974 2390 1976
rect 2794 1964 2806 2796
rect 2826 2384 2838 3456
rect 2954 3124 2966 3126
rect 2954 3116 2956 3124
rect 2964 3116 2966 3124
rect 2954 3064 2966 3116
rect 2954 3056 2956 3064
rect 2964 3056 2966 3064
rect 2954 3054 2966 3056
rect 2986 3024 2998 4176
rect 3210 4104 3222 4316
rect 3210 4096 3212 4104
rect 3220 4096 3222 4104
rect 3210 4094 3222 4096
rect 3304 4214 3352 4606
rect 3786 4724 3798 4726
rect 3786 4716 3788 4724
rect 3796 4716 3798 4724
rect 3304 4206 3308 4214
rect 3316 4206 3324 4214
rect 3332 4206 3340 4214
rect 3348 4206 3352 4214
rect 3658 4424 3670 4426
rect 3658 4416 3660 4424
rect 3668 4416 3670 4424
rect 3304 3814 3352 4206
rect 3562 4204 3574 4206
rect 3562 4196 3564 4204
rect 3572 4196 3574 4204
rect 3562 4164 3574 4196
rect 3562 4156 3564 4164
rect 3572 4156 3574 4164
rect 3562 4154 3574 4156
rect 3304 3806 3308 3814
rect 3316 3806 3324 3814
rect 3332 3806 3340 3814
rect 3348 3806 3352 3814
rect 2986 3016 2988 3024
rect 2996 3016 2998 3024
rect 2986 3014 2998 3016
rect 3082 3504 3094 3506
rect 3082 3496 3084 3504
rect 3092 3496 3094 3504
rect 3050 2744 3062 2746
rect 3050 2736 3052 2744
rect 3060 2736 3062 2744
rect 3050 2524 3062 2736
rect 3050 2516 3052 2524
rect 3060 2516 3062 2524
rect 3050 2514 3062 2516
rect 2826 2376 2828 2384
rect 2836 2376 2838 2384
rect 2826 2374 2838 2376
rect 2794 1956 2796 1964
rect 2804 1956 2806 1964
rect 2794 1954 2806 1956
rect 2922 2204 2934 2206
rect 2922 2196 2924 2204
rect 2932 2196 2934 2204
rect 2346 1916 2348 1924
rect 2356 1916 2358 1924
rect 2346 1914 2358 1916
rect 2922 1884 2934 2196
rect 3082 2124 3094 3496
rect 3304 3414 3352 3806
rect 3626 3864 3638 3866
rect 3626 3856 3628 3864
rect 3636 3856 3638 3864
rect 3626 3784 3638 3856
rect 3626 3776 3628 3784
rect 3636 3776 3638 3784
rect 3626 3774 3638 3776
rect 3658 3744 3670 4416
rect 3786 4424 3798 4716
rect 4650 4564 4662 4566
rect 4650 4556 4652 4564
rect 4660 4556 4662 4564
rect 4650 4484 4662 4556
rect 4650 4476 4652 4484
rect 4660 4476 4662 4484
rect 4650 4474 4662 4476
rect 3786 4416 3788 4424
rect 3796 4416 3798 4424
rect 3786 4414 3798 4416
rect 4746 4464 4758 4466
rect 4746 4456 4748 4464
rect 4756 4456 4758 4464
rect 4106 4384 4118 4386
rect 4106 4376 4108 4384
rect 4116 4376 4118 4384
rect 3946 4324 3958 4326
rect 3946 4316 3948 4324
rect 3956 4316 3958 4324
rect 3946 4284 3958 4316
rect 3946 4276 3948 4284
rect 3956 4276 3958 4284
rect 3946 4274 3958 4276
rect 4074 4264 4086 4266
rect 4074 4256 4076 4264
rect 4084 4256 4086 4264
rect 3658 3736 3660 3744
rect 3668 3736 3670 3744
rect 3658 3734 3670 3736
rect 3818 3904 3830 3906
rect 3818 3896 3820 3904
rect 3828 3896 3830 3904
rect 3818 3664 3830 3896
rect 3818 3656 3820 3664
rect 3828 3656 3830 3664
rect 3304 3406 3308 3414
rect 3316 3406 3324 3414
rect 3332 3406 3340 3414
rect 3348 3406 3352 3414
rect 3304 3014 3352 3406
rect 3658 3524 3670 3526
rect 3658 3516 3660 3524
rect 3668 3516 3670 3524
rect 3658 3384 3670 3516
rect 3658 3376 3660 3384
rect 3668 3376 3670 3384
rect 3658 3374 3670 3376
rect 3722 3224 3734 3226
rect 3722 3216 3724 3224
rect 3732 3216 3734 3224
rect 3722 3124 3734 3216
rect 3722 3116 3724 3124
rect 3732 3116 3734 3124
rect 3722 3114 3734 3116
rect 3304 3006 3308 3014
rect 3316 3006 3324 3014
rect 3332 3006 3340 3014
rect 3348 3006 3352 3014
rect 3304 2614 3352 3006
rect 3818 2884 3830 3656
rect 4074 3584 4086 4256
rect 4106 3884 4118 4376
rect 4106 3876 4108 3884
rect 4116 3876 4118 3884
rect 4106 3874 4118 3876
rect 4362 4304 4374 4306
rect 4362 4296 4364 4304
rect 4372 4296 4374 4304
rect 4362 3764 4374 4296
rect 4714 4284 4726 4286
rect 4714 4276 4716 4284
rect 4724 4276 4726 4284
rect 4362 3756 4364 3764
rect 4372 3756 4374 3764
rect 4362 3754 4374 3756
rect 4458 4124 4470 4126
rect 4458 4116 4460 4124
rect 4468 4116 4470 4124
rect 4074 3576 4076 3584
rect 4084 3576 4086 3584
rect 4074 3574 4086 3576
rect 4106 3704 4118 3706
rect 4106 3696 4108 3704
rect 4116 3696 4118 3704
rect 3882 3424 3894 3426
rect 3882 3416 3884 3424
rect 3892 3416 3894 3424
rect 3882 3124 3894 3416
rect 4042 3404 4054 3406
rect 4042 3396 4044 3404
rect 4052 3396 4054 3404
rect 4042 3184 4054 3396
rect 4042 3176 4044 3184
rect 4052 3176 4054 3184
rect 4042 3174 4054 3176
rect 3882 3116 3884 3124
rect 3892 3116 3894 3124
rect 3882 3114 3894 3116
rect 4010 3124 4022 3126
rect 4010 3116 4012 3124
rect 4020 3116 4022 3124
rect 4010 3004 4022 3116
rect 4010 2996 4012 3004
rect 4020 2996 4022 3004
rect 4010 2994 4022 2996
rect 4074 3104 4086 3106
rect 4074 3096 4076 3104
rect 4084 3096 4086 3104
rect 4074 2984 4086 3096
rect 4074 2976 4076 2984
rect 4084 2976 4086 2984
rect 4074 2974 4086 2976
rect 3818 2876 3820 2884
rect 3828 2876 3830 2884
rect 3818 2874 3830 2876
rect 4106 2864 4118 3696
rect 4458 3544 4470 4116
rect 4714 3964 4726 4276
rect 4746 4184 4758 4456
rect 4746 4176 4748 4184
rect 4756 4176 4758 4184
rect 4746 4174 4758 4176
rect 4824 4414 4872 4806
rect 6570 4764 6582 4766
rect 6570 4756 6572 4764
rect 6580 4756 6582 4764
rect 6314 4744 6326 4746
rect 6314 4736 6316 4744
rect 6324 4736 6326 4744
rect 5162 4724 5174 4726
rect 5162 4716 5164 4724
rect 5172 4716 5174 4724
rect 5162 4424 5174 4716
rect 5866 4684 5878 4686
rect 5866 4676 5868 4684
rect 5876 4676 5878 4684
rect 5866 4644 5878 4676
rect 6154 4684 6166 4686
rect 6154 4676 6156 4684
rect 6164 4676 6166 4684
rect 5866 4636 5868 4644
rect 5876 4636 5878 4644
rect 5866 4634 5878 4636
rect 6026 4664 6038 4666
rect 6026 4656 6028 4664
rect 6036 4656 6038 4664
rect 5866 4604 5878 4606
rect 5866 4596 5868 4604
rect 5876 4596 5878 4604
rect 5514 4584 5526 4586
rect 5514 4576 5516 4584
rect 5524 4576 5526 4584
rect 5162 4416 5164 4424
rect 5172 4416 5174 4424
rect 5162 4414 5174 4416
rect 5386 4564 5398 4566
rect 5386 4556 5388 4564
rect 5396 4556 5398 4564
rect 4824 4406 4828 4414
rect 4836 4406 4844 4414
rect 4852 4406 4860 4414
rect 4868 4406 4872 4414
rect 4714 3956 4716 3964
rect 4724 3956 4726 3964
rect 4714 3954 4726 3956
rect 4824 4014 4872 4406
rect 5130 4224 5142 4226
rect 5130 4216 5132 4224
rect 5140 4216 5142 4224
rect 5066 4164 5078 4166
rect 5066 4156 5068 4164
rect 5076 4156 5078 4164
rect 4824 4006 4828 4014
rect 4836 4006 4844 4014
rect 4852 4006 4860 4014
rect 4868 4006 4872 4014
rect 4458 3536 4460 3544
rect 4468 3536 4470 3544
rect 4458 3534 4470 3536
rect 4824 3614 4872 4006
rect 5002 4064 5014 4066
rect 5002 4056 5004 4064
rect 5012 4056 5014 4064
rect 5002 3864 5014 4056
rect 5002 3856 5004 3864
rect 5012 3856 5014 3864
rect 5002 3854 5014 3856
rect 5034 4004 5046 4006
rect 5034 3996 5036 4004
rect 5044 3996 5046 4004
rect 4824 3606 4828 3614
rect 4836 3606 4844 3614
rect 4852 3606 4860 3614
rect 4868 3606 4872 3614
rect 4234 3424 4246 3426
rect 4234 3416 4236 3424
rect 4244 3416 4246 3424
rect 4106 2856 4108 2864
rect 4116 2856 4118 2864
rect 4106 2854 4118 2856
rect 4170 3104 4182 3106
rect 4170 3096 4172 3104
rect 4180 3096 4182 3104
rect 4170 2864 4182 3096
rect 4234 2924 4246 3416
rect 4266 3364 4278 3366
rect 4266 3356 4268 3364
rect 4276 3356 4278 3364
rect 4266 3104 4278 3356
rect 4618 3304 4630 3306
rect 4618 3296 4620 3304
rect 4628 3296 4630 3304
rect 4618 3164 4630 3296
rect 4618 3156 4620 3164
rect 4628 3156 4630 3164
rect 4618 3154 4630 3156
rect 4824 3214 4872 3606
rect 4824 3206 4828 3214
rect 4836 3206 4844 3214
rect 4852 3206 4860 3214
rect 4868 3206 4872 3214
rect 4266 3096 4268 3104
rect 4276 3096 4278 3104
rect 4266 3094 4278 3096
rect 4330 3144 4342 3146
rect 4330 3136 4332 3144
rect 4340 3136 4342 3144
rect 4234 2916 4236 2924
rect 4244 2916 4246 2924
rect 4234 2914 4246 2916
rect 4298 3024 4310 3026
rect 4298 3016 4300 3024
rect 4308 3016 4310 3024
rect 4298 2904 4310 3016
rect 4330 2944 4342 3136
rect 4490 3084 4502 3086
rect 4490 3076 4492 3084
rect 4500 3076 4502 3084
rect 4490 3046 4502 3076
rect 4490 3044 4534 3046
rect 4490 3036 4524 3044
rect 4532 3036 4534 3044
rect 4490 3034 4534 3036
rect 4618 2964 4630 2966
rect 4618 2956 4620 2964
rect 4628 2956 4630 2964
rect 4330 2936 4332 2944
rect 4340 2936 4342 2944
rect 4330 2934 4342 2936
rect 4490 2944 4502 2946
rect 4490 2936 4492 2944
rect 4500 2936 4502 2944
rect 4298 2896 4300 2904
rect 4308 2896 4310 2904
rect 4298 2894 4310 2896
rect 4170 2856 4172 2864
rect 4180 2856 4182 2864
rect 4170 2854 4182 2856
rect 4490 2784 4502 2936
rect 4618 2844 4630 2956
rect 4714 2944 4726 2946
rect 4714 2936 4716 2944
rect 4724 2936 4726 2944
rect 4714 2884 4726 2936
rect 4714 2876 4716 2884
rect 4724 2876 4726 2884
rect 4714 2874 4726 2876
rect 4746 2924 4758 2926
rect 4746 2916 4748 2924
rect 4756 2916 4758 2924
rect 4746 2846 4758 2916
rect 4618 2836 4620 2844
rect 4628 2836 4630 2844
rect 4618 2834 4630 2836
rect 4714 2844 4758 2846
rect 4714 2836 4716 2844
rect 4724 2836 4758 2844
rect 4714 2834 4758 2836
rect 4490 2776 4492 2784
rect 4500 2776 4502 2784
rect 4490 2774 4502 2776
rect 4824 2814 4872 3206
rect 4906 3804 4918 3806
rect 4906 3796 4908 3804
rect 4916 3796 4918 3804
rect 4906 3204 4918 3796
rect 5034 3744 5046 3996
rect 5034 3736 5036 3744
rect 5044 3736 5046 3744
rect 5034 3734 5046 3736
rect 4970 3604 4982 3606
rect 4970 3596 4972 3604
rect 4980 3596 4982 3604
rect 4970 3384 4982 3596
rect 4970 3376 4972 3384
rect 4980 3376 4982 3384
rect 4970 3374 4982 3376
rect 4906 3196 4908 3204
rect 4916 3196 4918 3204
rect 4906 3194 4918 3196
rect 4938 3244 4950 3246
rect 4938 3236 4940 3244
rect 4948 3236 4950 3244
rect 4938 3184 4950 3236
rect 4938 3176 4940 3184
rect 4948 3176 4950 3184
rect 4938 3174 4950 3176
rect 5066 3084 5078 4156
rect 5098 3824 5110 3826
rect 5098 3816 5100 3824
rect 5108 3816 5110 3824
rect 5098 3704 5110 3816
rect 5098 3696 5100 3704
rect 5108 3696 5110 3704
rect 5098 3664 5110 3696
rect 5130 3784 5142 4216
rect 5194 3924 5222 3926
rect 5194 3916 5212 3924
rect 5220 3916 5222 3924
rect 5194 3914 5222 3916
rect 5194 3904 5206 3914
rect 5194 3896 5196 3904
rect 5204 3896 5206 3904
rect 5194 3894 5206 3896
rect 5130 3776 5132 3784
rect 5140 3776 5142 3784
rect 5130 3704 5142 3776
rect 5130 3696 5132 3704
rect 5140 3696 5142 3704
rect 5130 3694 5142 3696
rect 5354 3784 5366 3786
rect 5354 3776 5356 3784
rect 5364 3776 5366 3784
rect 5098 3656 5100 3664
rect 5108 3656 5110 3664
rect 5098 3654 5110 3656
rect 5354 3644 5366 3776
rect 5386 3704 5398 4556
rect 5514 3744 5526 4576
rect 5514 3736 5516 3744
rect 5524 3736 5526 3744
rect 5514 3734 5526 3736
rect 5578 4484 5590 4486
rect 5578 4476 5580 4484
rect 5588 4476 5590 4484
rect 5386 3696 5388 3704
rect 5396 3696 5398 3704
rect 5386 3694 5398 3696
rect 5354 3636 5356 3644
rect 5364 3636 5366 3644
rect 5354 3634 5366 3636
rect 5418 3684 5430 3686
rect 5418 3676 5420 3684
rect 5428 3676 5430 3684
rect 5418 3264 5430 3676
rect 5578 3464 5590 4476
rect 5770 4464 5782 4466
rect 5770 4456 5772 4464
rect 5780 4456 5782 4464
rect 5770 4164 5782 4456
rect 5770 4156 5772 4164
rect 5780 4156 5782 4164
rect 5770 4154 5782 4156
rect 5802 4364 5814 4366
rect 5802 4356 5804 4364
rect 5812 4356 5814 4364
rect 5770 4004 5782 4006
rect 5770 3996 5772 4004
rect 5780 3996 5782 4004
rect 5706 3724 5750 3726
rect 5706 3716 5708 3724
rect 5716 3716 5750 3724
rect 5706 3714 5750 3716
rect 5738 3704 5750 3714
rect 5738 3696 5740 3704
rect 5748 3696 5750 3704
rect 5738 3694 5750 3696
rect 5578 3456 5580 3464
rect 5588 3456 5590 3464
rect 5578 3454 5590 3456
rect 5610 3484 5622 3486
rect 5610 3476 5612 3484
rect 5620 3476 5622 3484
rect 5418 3256 5420 3264
rect 5428 3256 5430 3264
rect 5418 3254 5430 3256
rect 5066 3076 5068 3084
rect 5076 3076 5078 3084
rect 5066 3074 5078 3076
rect 5354 3124 5366 3126
rect 5354 3116 5356 3124
rect 5364 3116 5366 3124
rect 4824 2806 4828 2814
rect 4836 2806 4844 2814
rect 4852 2806 4860 2814
rect 4868 2806 4872 2814
rect 4266 2744 4278 2746
rect 4266 2736 4268 2744
rect 4276 2736 4278 2744
rect 3304 2606 3308 2614
rect 3316 2606 3324 2614
rect 3332 2606 3340 2614
rect 3348 2606 3352 2614
rect 3274 2264 3286 2266
rect 3274 2256 3276 2264
rect 3284 2256 3286 2264
rect 3274 2144 3286 2256
rect 3274 2136 3276 2144
rect 3284 2136 3286 2144
rect 3274 2134 3286 2136
rect 3304 2214 3352 2606
rect 4202 2664 4214 2666
rect 4202 2656 4204 2664
rect 4212 2656 4214 2664
rect 4106 2584 4118 2586
rect 4106 2576 4108 2584
rect 4116 2576 4118 2584
rect 3914 2564 3926 2566
rect 3914 2556 3916 2564
rect 3924 2556 3926 2564
rect 3304 2206 3308 2214
rect 3316 2206 3324 2214
rect 3332 2206 3340 2214
rect 3348 2206 3352 2214
rect 3082 2116 3084 2124
rect 3092 2116 3094 2124
rect 3082 2114 3094 2116
rect 2922 1876 2924 1884
rect 2932 1876 2934 1884
rect 2922 1874 2934 1876
rect 1768 1606 1772 1614
rect 1780 1606 1788 1614
rect 1796 1606 1804 1614
rect 1812 1606 1816 1614
rect 1514 1524 1526 1526
rect 1514 1516 1516 1524
rect 1524 1516 1526 1524
rect 1514 1324 1526 1516
rect 1514 1316 1516 1324
rect 1524 1316 1526 1324
rect 1514 1314 1526 1316
rect 1578 1424 1590 1426
rect 1578 1416 1580 1424
rect 1588 1416 1590 1424
rect 1482 1296 1484 1304
rect 1492 1296 1494 1304
rect 1482 1294 1494 1296
rect 1578 1304 1590 1416
rect 1578 1296 1580 1304
rect 1588 1296 1590 1304
rect 1578 1244 1590 1296
rect 1674 1424 1686 1426
rect 1674 1416 1676 1424
rect 1684 1416 1686 1424
rect 1674 1304 1686 1416
rect 1674 1296 1676 1304
rect 1684 1296 1686 1304
rect 1674 1294 1686 1296
rect 1578 1236 1580 1244
rect 1588 1236 1590 1244
rect 1578 1234 1590 1236
rect 1768 1214 1816 1606
rect 3304 1814 3352 2206
rect 3530 2264 3542 2266
rect 3530 2256 3532 2264
rect 3540 2256 3542 2264
rect 3304 1806 3308 1814
rect 3316 1806 3324 1814
rect 3332 1806 3340 1814
rect 3348 1806 3352 1814
rect 1930 1524 1942 1526
rect 1930 1516 1932 1524
rect 1940 1516 1942 1524
rect 1930 1304 1942 1516
rect 2986 1484 2998 1486
rect 2986 1476 2988 1484
rect 2996 1476 2998 1484
rect 2986 1344 2998 1476
rect 2986 1336 2988 1344
rect 2996 1336 2998 1344
rect 2986 1334 2998 1336
rect 3304 1414 3352 1806
rect 3402 2164 3414 2166
rect 3402 2156 3404 2164
rect 3412 2156 3414 2164
rect 3402 1544 3414 2156
rect 3530 1604 3542 2256
rect 3914 1764 3926 2556
rect 4106 2504 4118 2576
rect 4106 2496 4108 2504
rect 4116 2496 4118 2504
rect 4106 2494 4118 2496
rect 4202 2504 4214 2656
rect 4202 2496 4204 2504
rect 4212 2496 4214 2504
rect 4202 2494 4214 2496
rect 3914 1756 3916 1764
rect 3924 1756 3926 1764
rect 3914 1754 3926 1756
rect 3946 1824 3958 1826
rect 3946 1816 3948 1824
rect 3956 1816 3958 1824
rect 3530 1596 3532 1604
rect 3540 1596 3542 1604
rect 3530 1594 3542 1596
rect 3402 1536 3404 1544
rect 3412 1536 3414 1544
rect 3402 1534 3414 1536
rect 3946 1524 3958 1816
rect 3946 1516 3948 1524
rect 3956 1516 3958 1524
rect 3946 1514 3958 1516
rect 4042 1524 4054 1526
rect 4042 1516 4044 1524
rect 4052 1516 4054 1524
rect 3304 1406 3308 1414
rect 3316 1406 3324 1414
rect 3332 1406 3340 1414
rect 3348 1406 3352 1414
rect 1930 1296 1932 1304
rect 1940 1296 1942 1304
rect 1930 1294 1942 1296
rect 1768 1206 1772 1214
rect 1780 1206 1788 1214
rect 1796 1206 1804 1214
rect 1812 1206 1816 1214
rect 1386 1096 1388 1104
rect 1396 1096 1398 1104
rect 1386 1094 1398 1096
rect 1706 1104 1718 1106
rect 1706 1096 1708 1104
rect 1716 1096 1718 1104
rect 1290 1076 1292 1084
rect 1300 1076 1302 1084
rect 1290 1074 1302 1076
rect 1290 1044 1302 1046
rect 1290 1036 1292 1044
rect 1300 1036 1302 1044
rect 1290 724 1302 1036
rect 1290 716 1292 724
rect 1300 716 1302 724
rect 1290 714 1302 716
rect 1482 1044 1494 1046
rect 1482 1036 1484 1044
rect 1492 1036 1494 1044
rect 1258 696 1260 704
rect 1268 696 1270 704
rect 1258 694 1270 696
rect 1194 516 1196 524
rect 1204 516 1206 524
rect 1194 514 1206 516
rect 1482 544 1494 1036
rect 1706 884 1718 1096
rect 1706 876 1708 884
rect 1716 876 1718 884
rect 1706 874 1718 876
rect 1482 536 1484 544
rect 1492 536 1494 544
rect 810 476 812 484
rect 820 476 822 484
rect 810 474 822 476
rect 682 416 684 424
rect 692 416 694 424
rect 682 414 694 416
rect 746 394 822 406
rect 746 366 758 394
rect 810 384 822 394
rect 810 376 812 384
rect 820 376 822 384
rect 810 374 822 376
rect 874 404 886 406
rect 874 396 876 404
rect 884 396 886 404
rect 618 354 758 366
rect 778 364 790 366
rect 778 356 780 364
rect 788 356 790 364
rect 618 104 630 354
rect 666 324 694 326
rect 666 316 668 324
rect 676 316 694 324
rect 666 314 694 316
rect 682 246 694 314
rect 778 284 790 356
rect 778 276 780 284
rect 788 276 790 284
rect 778 274 790 276
rect 874 284 886 396
rect 1482 344 1494 536
rect 1768 814 1816 1206
rect 3242 1204 3254 1206
rect 3242 1196 3244 1204
rect 3252 1196 3254 1204
rect 2090 1124 2102 1126
rect 2090 1116 2092 1124
rect 2100 1116 2102 1124
rect 1768 806 1772 814
rect 1780 806 1788 814
rect 1796 806 1804 814
rect 1812 806 1816 814
rect 1482 336 1484 344
rect 1492 336 1494 344
rect 1482 334 1494 336
rect 1674 444 1686 446
rect 1674 436 1676 444
rect 1684 436 1686 444
rect 874 276 876 284
rect 884 276 886 284
rect 874 274 886 276
rect 938 304 950 306
rect 938 296 940 304
rect 948 296 950 304
rect 938 246 950 296
rect 682 234 950 246
rect 1258 284 1270 286
rect 1258 276 1260 284
rect 1268 276 1270 284
rect 842 164 854 166
rect 842 156 844 164
rect 852 156 854 164
rect 714 144 726 146
rect 714 136 716 144
rect 724 136 726 144
rect 714 126 726 136
rect 778 144 790 146
rect 778 136 780 144
rect 788 136 790 144
rect 778 126 790 136
rect 842 126 854 156
rect 1258 164 1270 276
rect 1258 156 1260 164
rect 1268 156 1270 164
rect 1258 154 1270 156
rect 714 114 854 126
rect 938 144 950 146
rect 938 136 940 144
rect 948 136 950 144
rect 618 96 620 104
rect 628 96 630 104
rect 618 94 630 96
rect 586 76 588 84
rect 596 76 598 84
rect 586 74 598 76
rect 938 84 950 136
rect 1578 144 1590 146
rect 1578 136 1580 144
rect 1588 136 1590 144
rect 938 76 940 84
rect 948 76 950 84
rect 938 74 950 76
rect 1514 124 1526 126
rect 1514 116 1516 124
rect 1524 116 1526 124
rect 1514 86 1526 116
rect 1578 86 1590 136
rect 1514 74 1590 86
rect 1674 64 1686 436
rect 1674 56 1676 64
rect 1684 56 1686 64
rect 1674 54 1686 56
rect 1768 414 1816 806
rect 2026 1064 2038 1066
rect 2026 1056 2028 1064
rect 2036 1056 2038 1064
rect 2026 604 2038 1056
rect 2090 684 2102 1116
rect 2698 824 2710 826
rect 2698 816 2700 824
rect 2708 816 2710 824
rect 2090 676 2092 684
rect 2100 676 2102 684
rect 2090 674 2102 676
rect 2538 804 2550 806
rect 2538 796 2540 804
rect 2548 796 2550 804
rect 2538 764 2550 796
rect 2538 756 2540 764
rect 2548 756 2550 764
rect 2538 664 2550 756
rect 2698 684 2710 816
rect 2698 676 2700 684
rect 2708 676 2710 684
rect 2698 674 2710 676
rect 2538 656 2540 664
rect 2548 656 2550 664
rect 2538 654 2550 656
rect 2026 596 2028 604
rect 2036 596 2038 604
rect 2026 594 2038 596
rect 2058 624 2070 626
rect 2058 616 2060 624
rect 2068 616 2070 624
rect 1768 406 1772 414
rect 1780 406 1788 414
rect 1796 406 1804 414
rect 1812 406 1816 414
rect 1866 444 1878 446
rect 1866 436 1868 444
rect 1876 436 1878 444
rect 1768 14 1816 406
rect 1834 404 1846 406
rect 1834 396 1836 404
rect 1844 396 1846 404
rect 1834 264 1846 396
rect 1834 256 1836 264
rect 1844 256 1846 264
rect 1834 254 1846 256
rect 1866 264 1878 436
rect 1866 256 1868 264
rect 1876 256 1878 264
rect 1866 254 1878 256
rect 2026 404 2038 406
rect 2026 396 2028 404
rect 2036 396 2038 404
rect 2026 206 2038 396
rect 2058 404 2070 616
rect 2090 624 2102 626
rect 2090 616 2092 624
rect 2100 616 2102 624
rect 2090 464 2102 616
rect 2090 456 2092 464
rect 2100 456 2102 464
rect 2090 454 2102 456
rect 2378 504 2390 506
rect 2378 496 2380 504
rect 2388 496 2390 504
rect 2058 396 2060 404
rect 2068 396 2070 404
rect 2058 394 2070 396
rect 2378 244 2390 496
rect 2474 384 2486 386
rect 2474 376 2476 384
rect 2484 376 2486 384
rect 2474 304 2486 376
rect 3146 324 3158 326
rect 3146 316 3148 324
rect 3156 316 3158 324
rect 2474 296 2476 304
rect 2484 296 2486 304
rect 2474 294 2486 296
rect 2570 304 2582 306
rect 2570 296 2572 304
rect 2580 296 2582 304
rect 2570 286 2582 296
rect 3146 286 3158 316
rect 2570 274 2614 286
rect 3130 284 3158 286
rect 3130 276 3132 284
rect 3140 276 3158 284
rect 3130 274 3158 276
rect 2602 264 2614 274
rect 2602 256 2604 264
rect 2612 256 2614 264
rect 2602 254 2614 256
rect 3050 264 3062 266
rect 3050 256 3052 264
rect 3060 256 3062 264
rect 2378 236 2380 244
rect 2388 236 2390 244
rect 2378 234 2390 236
rect 3050 224 3062 256
rect 3050 216 3052 224
rect 3060 216 3062 224
rect 3050 214 3062 216
rect 3242 224 3254 1196
rect 3304 1014 3352 1406
rect 3658 1484 3670 1486
rect 3658 1476 3660 1484
rect 3668 1476 3670 1484
rect 3304 1006 3308 1014
rect 3316 1006 3324 1014
rect 3332 1006 3340 1014
rect 3348 1006 3352 1014
rect 3274 864 3286 866
rect 3274 856 3276 864
rect 3284 856 3286 864
rect 3274 564 3286 856
rect 3274 556 3276 564
rect 3284 556 3286 564
rect 3274 554 3286 556
rect 3304 614 3352 1006
rect 3562 1324 3574 1326
rect 3562 1316 3564 1324
rect 3572 1316 3574 1324
rect 3562 824 3574 1316
rect 3658 1284 3670 1476
rect 3818 1344 3830 1346
rect 3818 1336 3820 1344
rect 3828 1336 3830 1344
rect 3818 1326 3830 1336
rect 4042 1344 4054 1516
rect 4042 1336 4044 1344
rect 4052 1336 4054 1344
rect 4042 1334 4054 1336
rect 3818 1324 3846 1326
rect 3818 1316 3836 1324
rect 3844 1316 3846 1324
rect 3818 1314 3846 1316
rect 3882 1324 3894 1326
rect 3882 1316 3884 1324
rect 3892 1316 3894 1324
rect 3658 1276 3660 1284
rect 3668 1276 3670 1284
rect 3658 1274 3670 1276
rect 3882 1264 3894 1316
rect 3882 1256 3884 1264
rect 3892 1256 3894 1264
rect 3882 1254 3894 1256
rect 3914 1084 3926 1086
rect 3914 1076 3916 1084
rect 3924 1076 3926 1084
rect 3914 844 3926 1076
rect 3914 836 3916 844
rect 3924 836 3926 844
rect 3914 834 3926 836
rect 3562 816 3564 824
rect 3572 816 3574 824
rect 3562 814 3574 816
rect 3304 606 3308 614
rect 3316 606 3324 614
rect 3332 606 3340 614
rect 3348 606 3352 614
rect 3242 216 3244 224
rect 3252 216 3254 224
rect 3242 214 3254 216
rect 3304 214 3352 606
rect 3498 664 3510 666
rect 3498 656 3500 664
rect 3508 656 3510 664
rect 3498 504 3510 656
rect 3498 496 3500 504
rect 3508 496 3510 504
rect 3498 494 3510 496
rect 3882 504 3894 506
rect 3882 496 3884 504
rect 3892 496 3894 504
rect 3882 486 3894 496
rect 3882 484 3926 486
rect 3882 476 3916 484
rect 3924 476 3926 484
rect 3882 474 3926 476
rect 3402 384 3414 386
rect 3402 376 3404 384
rect 3412 376 3414 384
rect 3304 206 3308 214
rect 3316 206 3324 214
rect 3332 206 3340 214
rect 3348 206 3352 214
rect 2026 204 2054 206
rect 2026 196 2044 204
rect 2052 196 2054 204
rect 2026 194 2054 196
rect 3082 204 3094 206
rect 3082 196 3084 204
rect 3092 196 3094 204
rect 2922 184 2934 186
rect 2922 176 2924 184
rect 2932 176 2934 184
rect 2922 166 2934 176
rect 3082 166 3094 196
rect 2874 164 2998 166
rect 2874 156 2876 164
rect 2884 156 2988 164
rect 2996 156 2998 164
rect 2874 154 2998 156
rect 3018 164 3030 166
rect 3018 156 3020 164
rect 3028 156 3030 164
rect 3018 126 3030 156
rect 1898 124 1910 126
rect 1898 116 1900 124
rect 1908 116 1910 124
rect 1898 86 1910 116
rect 2922 114 3030 126
rect 3050 154 3094 166
rect 3274 184 3286 186
rect 3274 176 3276 184
rect 3284 176 3286 184
rect 1898 84 1958 86
rect 1898 76 1948 84
rect 1956 76 1958 84
rect 1898 74 1958 76
rect 2474 84 2502 86
rect 2474 76 2492 84
rect 2500 76 2502 84
rect 2474 74 2502 76
rect 2474 64 2486 74
rect 2474 56 2476 64
rect 2484 56 2486 64
rect 2474 54 2486 56
rect 2858 64 2870 66
rect 2858 56 2860 64
rect 2868 56 2870 64
rect 2858 46 2870 56
rect 2922 64 2934 114
rect 3050 86 3062 154
rect 2922 56 2924 64
rect 2932 56 2934 64
rect 2922 54 2934 56
rect 3018 74 3062 86
rect 2794 44 2870 46
rect 2794 36 2796 44
rect 2804 36 2870 44
rect 2794 34 2870 36
rect 3018 24 3030 74
rect 3018 16 3020 24
rect 3028 16 3030 24
rect 3018 14 3030 16
rect 3274 24 3286 176
rect 3274 16 3276 24
rect 3284 16 3286 24
rect 3274 14 3286 16
rect 1768 6 1772 14
rect 1780 6 1788 14
rect 1796 6 1804 14
rect 1812 6 1816 14
rect 1768 -40 1816 6
rect 3304 -40 3352 206
rect 3370 224 3382 226
rect 3370 216 3372 224
rect 3380 216 3382 224
rect 3370 84 3382 216
rect 3402 204 3414 376
rect 3402 196 3404 204
rect 3412 196 3414 204
rect 3402 194 3414 196
rect 3434 344 3446 346
rect 3434 336 3436 344
rect 3444 336 3446 344
rect 3434 144 3446 336
rect 3818 324 3830 326
rect 3818 316 3820 324
rect 3828 316 3830 324
rect 3818 204 3830 316
rect 4266 264 4278 2736
rect 4746 2684 4758 2686
rect 4746 2676 4748 2684
rect 4756 2676 4758 2684
rect 4586 2524 4598 2526
rect 4586 2516 4588 2524
rect 4596 2516 4598 2524
rect 4362 2404 4374 2406
rect 4362 2396 4364 2404
rect 4372 2396 4374 2404
rect 4362 1204 4374 2396
rect 4522 2284 4534 2286
rect 4522 2276 4524 2284
rect 4532 2276 4534 2284
rect 4522 1824 4534 2276
rect 4586 2244 4598 2516
rect 4746 2404 4758 2676
rect 4746 2396 4748 2404
rect 4756 2396 4758 2404
rect 4746 2394 4758 2396
rect 4824 2414 4872 2806
rect 5002 2584 5014 2586
rect 5002 2576 5004 2584
rect 5012 2576 5014 2584
rect 4824 2406 4828 2414
rect 4836 2406 4844 2414
rect 4852 2406 4860 2414
rect 4868 2406 4872 2414
rect 4586 2236 4588 2244
rect 4596 2236 4598 2244
rect 4586 2234 4598 2236
rect 4682 2224 4694 2226
rect 4682 2216 4684 2224
rect 4692 2216 4694 2224
rect 4586 2124 4598 2126
rect 4586 2116 4588 2124
rect 4596 2116 4598 2124
rect 4586 2004 4598 2116
rect 4586 1996 4588 2004
rect 4596 1996 4598 2004
rect 4586 1994 4598 1996
rect 4522 1816 4524 1824
rect 4532 1816 4534 1824
rect 4522 1814 4534 1816
rect 4682 1684 4694 2216
rect 4682 1676 4684 1684
rect 4692 1676 4694 1684
rect 4682 1674 4694 1676
rect 4824 2014 4872 2406
rect 4938 2544 4950 2546
rect 4938 2536 4940 2544
rect 4948 2536 4950 2544
rect 4938 2324 4950 2536
rect 5002 2544 5014 2576
rect 5002 2536 5004 2544
rect 5012 2536 5014 2544
rect 5002 2534 5014 2536
rect 5130 2564 5142 2566
rect 5130 2556 5132 2564
rect 5140 2556 5142 2564
rect 5130 2444 5142 2556
rect 5130 2436 5132 2444
rect 5140 2436 5142 2444
rect 5130 2434 5142 2436
rect 4938 2316 4940 2324
rect 4948 2316 4950 2324
rect 4938 2084 4950 2316
rect 4938 2076 4940 2084
rect 4948 2076 4950 2084
rect 4938 2074 4950 2076
rect 5066 2284 5078 2286
rect 5066 2276 5068 2284
rect 5076 2276 5078 2284
rect 5066 2064 5078 2276
rect 5066 2056 5068 2064
rect 5076 2056 5078 2064
rect 5066 2054 5078 2056
rect 4824 2006 4828 2014
rect 4836 2006 4844 2014
rect 4852 2006 4860 2014
rect 4868 2006 4872 2014
rect 4824 1614 4872 2006
rect 5354 1964 5366 3116
rect 5610 3044 5622 3476
rect 5770 3444 5782 3996
rect 5802 3744 5814 4356
rect 5866 4064 5878 4596
rect 6026 4544 6038 4656
rect 6026 4536 6028 4544
rect 6036 4536 6038 4544
rect 6026 4534 6038 4536
rect 6058 4584 6070 4586
rect 6058 4576 6060 4584
rect 6068 4576 6070 4584
rect 6026 4304 6038 4306
rect 6026 4296 6028 4304
rect 6036 4296 6038 4304
rect 5866 4056 5868 4064
rect 5876 4056 5878 4064
rect 5866 4054 5878 4056
rect 5930 4244 5942 4246
rect 5930 4236 5932 4244
rect 5940 4236 5942 4244
rect 5802 3736 5804 3744
rect 5812 3736 5814 3744
rect 5802 3544 5814 3736
rect 5802 3536 5804 3544
rect 5812 3536 5814 3544
rect 5802 3534 5814 3536
rect 5770 3436 5772 3444
rect 5780 3436 5782 3444
rect 5770 3434 5782 3436
rect 5834 3444 5846 3446
rect 5834 3436 5836 3444
rect 5844 3436 5846 3444
rect 5770 3404 5782 3406
rect 5770 3396 5772 3404
rect 5780 3396 5782 3404
rect 5706 3324 5718 3326
rect 5706 3316 5708 3324
rect 5716 3316 5718 3324
rect 5610 3036 5612 3044
rect 5620 3036 5622 3044
rect 5610 3034 5622 3036
rect 5642 3064 5654 3066
rect 5642 3056 5644 3064
rect 5652 3056 5654 3064
rect 5642 2964 5654 3056
rect 5642 2956 5644 2964
rect 5652 2956 5654 2964
rect 5642 2954 5654 2956
rect 5546 2944 5558 2946
rect 5546 2936 5548 2944
rect 5556 2936 5558 2944
rect 5546 2864 5558 2936
rect 5546 2856 5548 2864
rect 5556 2856 5558 2864
rect 5546 2854 5558 2856
rect 5578 2504 5590 2506
rect 5578 2496 5580 2504
rect 5588 2496 5590 2504
rect 5482 2484 5494 2486
rect 5482 2476 5484 2484
rect 5492 2476 5494 2484
rect 5354 1956 5356 1964
rect 5364 1956 5366 1964
rect 5354 1954 5366 1956
rect 5386 1964 5398 1966
rect 5386 1956 5388 1964
rect 5396 1956 5398 1964
rect 5258 1914 5366 1926
rect 5258 1904 5270 1914
rect 5258 1896 5260 1904
rect 5268 1896 5270 1904
rect 5258 1894 5270 1896
rect 5354 1904 5366 1914
rect 5354 1896 5356 1904
rect 5364 1896 5366 1904
rect 5354 1894 5366 1896
rect 4824 1606 4828 1614
rect 4836 1606 4844 1614
rect 4852 1606 4860 1614
rect 4868 1606 4872 1614
rect 4522 1604 4534 1606
rect 4522 1596 4524 1604
rect 4532 1596 4534 1604
rect 4522 1526 4534 1596
rect 4522 1514 4566 1526
rect 4554 1484 4566 1514
rect 4554 1476 4556 1484
rect 4564 1476 4566 1484
rect 4554 1474 4566 1476
rect 4362 1196 4364 1204
rect 4372 1196 4374 1204
rect 4362 1194 4374 1196
rect 4778 1384 4790 1386
rect 4778 1376 4780 1384
rect 4788 1376 4790 1384
rect 4554 744 4566 746
rect 4554 736 4556 744
rect 4564 736 4566 744
rect 4266 256 4268 264
rect 4276 256 4278 264
rect 4266 254 4278 256
rect 4522 604 4534 606
rect 4522 596 4524 604
rect 4532 596 4534 604
rect 3818 196 3820 204
rect 3828 196 3830 204
rect 3818 194 3830 196
rect 3434 136 3436 144
rect 3444 136 3446 144
rect 3434 134 3446 136
rect 4522 124 4534 596
rect 4554 564 4566 736
rect 4618 744 4630 746
rect 4618 736 4620 744
rect 4628 736 4630 744
rect 4618 624 4630 736
rect 4618 616 4620 624
rect 4628 616 4630 624
rect 4618 614 4630 616
rect 4554 556 4556 564
rect 4564 556 4566 564
rect 4554 554 4566 556
rect 4586 564 4598 566
rect 4586 556 4588 564
rect 4596 556 4598 564
rect 4586 524 4598 556
rect 4778 564 4790 1376
rect 4778 556 4780 564
rect 4788 556 4790 564
rect 4778 554 4790 556
rect 4824 1214 4872 1606
rect 4938 1884 4950 1886
rect 4938 1876 4940 1884
rect 4948 1876 4950 1884
rect 4938 1584 4950 1876
rect 4938 1576 4940 1584
rect 4948 1576 4950 1584
rect 4938 1574 4950 1576
rect 5034 1884 5046 1886
rect 5034 1876 5036 1884
rect 5044 1876 5046 1884
rect 5034 1744 5046 1876
rect 5194 1864 5206 1866
rect 5194 1856 5196 1864
rect 5204 1856 5206 1864
rect 5034 1736 5036 1744
rect 5044 1736 5046 1744
rect 4938 1364 4950 1366
rect 4938 1356 4940 1364
rect 4948 1356 4950 1364
rect 4938 1324 4950 1356
rect 4938 1316 4940 1324
rect 4948 1316 4950 1324
rect 4938 1314 4950 1316
rect 5034 1344 5046 1736
rect 5130 1804 5142 1806
rect 5130 1796 5132 1804
rect 5140 1796 5142 1804
rect 5034 1336 5036 1344
rect 5044 1336 5046 1344
rect 4824 1206 4828 1214
rect 4836 1206 4844 1214
rect 4852 1206 4860 1214
rect 4868 1206 4872 1214
rect 4824 814 4872 1206
rect 4824 806 4828 814
rect 4836 806 4844 814
rect 4852 806 4860 814
rect 4868 806 4872 814
rect 4586 516 4588 524
rect 4596 516 4598 524
rect 4586 514 4598 516
rect 4522 116 4524 124
rect 4532 116 4534 124
rect 4522 114 4534 116
rect 4824 414 4872 806
rect 5034 704 5046 1336
rect 5098 1644 5110 1646
rect 5098 1636 5100 1644
rect 5108 1636 5110 1644
rect 5066 1224 5078 1226
rect 5066 1216 5068 1224
rect 5076 1216 5078 1224
rect 5066 1004 5078 1216
rect 5066 996 5068 1004
rect 5076 996 5078 1004
rect 5066 994 5078 996
rect 5098 844 5110 1636
rect 5130 1244 5142 1796
rect 5130 1236 5132 1244
rect 5140 1236 5142 1244
rect 5130 1234 5142 1236
rect 5162 1364 5174 1366
rect 5162 1356 5164 1364
rect 5172 1356 5174 1364
rect 5098 836 5100 844
rect 5108 836 5110 844
rect 5098 834 5110 836
rect 5034 696 5036 704
rect 5044 696 5046 704
rect 5034 694 5046 696
rect 5162 564 5174 1356
rect 5162 556 5164 564
rect 5172 556 5174 564
rect 5162 554 5174 556
rect 5194 524 5206 1856
rect 5322 1504 5334 1506
rect 5322 1496 5324 1504
rect 5332 1496 5334 1504
rect 5322 1324 5334 1496
rect 5322 1316 5324 1324
rect 5332 1316 5334 1324
rect 5258 1164 5270 1166
rect 5258 1156 5260 1164
rect 5268 1156 5270 1164
rect 5258 1044 5270 1156
rect 5258 1036 5260 1044
rect 5268 1036 5270 1044
rect 5258 1034 5270 1036
rect 5322 864 5334 1316
rect 5322 856 5324 864
rect 5332 856 5334 864
rect 5322 854 5334 856
rect 5386 604 5398 1956
rect 5418 1864 5430 1866
rect 5418 1856 5420 1864
rect 5428 1856 5430 1864
rect 5418 1704 5430 1856
rect 5418 1696 5420 1704
rect 5428 1696 5430 1704
rect 5418 1694 5430 1696
rect 5482 1644 5494 2476
rect 5482 1636 5484 1644
rect 5492 1636 5494 1644
rect 5482 1634 5494 1636
rect 5514 2004 5526 2006
rect 5514 1996 5516 2004
rect 5524 1996 5526 2004
rect 5514 1664 5526 1996
rect 5514 1656 5516 1664
rect 5524 1656 5526 1664
rect 5450 1524 5462 1526
rect 5450 1516 5452 1524
rect 5460 1516 5462 1524
rect 5450 1384 5462 1516
rect 5450 1376 5452 1384
rect 5460 1376 5462 1384
rect 5450 1374 5462 1376
rect 5514 1364 5526 1656
rect 5578 1664 5590 2496
rect 5674 2504 5686 2506
rect 5674 2496 5676 2504
rect 5684 2496 5686 2504
rect 5642 2364 5654 2366
rect 5642 2356 5644 2364
rect 5652 2356 5654 2364
rect 5578 1656 5580 1664
rect 5588 1656 5590 1664
rect 5578 1654 5590 1656
rect 5610 2184 5622 2186
rect 5610 2176 5612 2184
rect 5620 2176 5622 2184
rect 5514 1356 5516 1364
rect 5524 1356 5526 1364
rect 5514 1354 5526 1356
rect 5418 1184 5430 1186
rect 5418 1176 5420 1184
rect 5428 1176 5430 1184
rect 5418 764 5430 1176
rect 5418 756 5420 764
rect 5428 756 5430 764
rect 5418 754 5430 756
rect 5386 596 5388 604
rect 5396 596 5398 604
rect 5386 594 5398 596
rect 5610 604 5622 2176
rect 5642 1264 5654 2356
rect 5674 1824 5686 2496
rect 5674 1816 5676 1824
rect 5684 1816 5686 1824
rect 5674 1814 5686 1816
rect 5642 1256 5644 1264
rect 5652 1256 5654 1264
rect 5642 1254 5654 1256
rect 5674 1604 5686 1606
rect 5674 1596 5676 1604
rect 5684 1596 5686 1604
rect 5610 596 5612 604
rect 5620 596 5622 604
rect 5610 594 5622 596
rect 5674 724 5686 1596
rect 5706 1204 5718 3316
rect 5738 3324 5750 3326
rect 5738 3316 5740 3324
rect 5748 3316 5750 3324
rect 5738 3084 5750 3316
rect 5738 3076 5740 3084
rect 5748 3076 5750 3084
rect 5738 3074 5750 3076
rect 5706 1196 5708 1204
rect 5716 1196 5718 1204
rect 5706 1194 5718 1196
rect 5738 1964 5750 1966
rect 5738 1956 5740 1964
rect 5748 1956 5750 1964
rect 5738 1104 5750 1956
rect 5770 1824 5782 3396
rect 5802 3004 5814 3006
rect 5802 2996 5804 3004
rect 5812 2996 5814 3004
rect 5802 2864 5814 2996
rect 5802 2856 5804 2864
rect 5812 2856 5814 2864
rect 5802 2854 5814 2856
rect 5770 1816 5772 1824
rect 5780 1816 5782 1824
rect 5770 1814 5782 1816
rect 5802 2524 5814 2526
rect 5802 2516 5804 2524
rect 5812 2516 5814 2524
rect 5802 1804 5814 2516
rect 5834 2184 5846 3436
rect 5898 3064 5910 3066
rect 5898 3056 5900 3064
rect 5908 3056 5910 3064
rect 5834 2176 5836 2184
rect 5844 2176 5846 2184
rect 5834 2174 5846 2176
rect 5866 2644 5878 2646
rect 5866 2636 5868 2644
rect 5876 2636 5878 2644
rect 5802 1796 5804 1804
rect 5812 1796 5814 1804
rect 5802 1794 5814 1796
rect 5802 1744 5814 1746
rect 5802 1736 5804 1744
rect 5812 1736 5814 1744
rect 5770 1504 5782 1506
rect 5770 1496 5772 1504
rect 5780 1496 5782 1504
rect 5770 1364 5782 1496
rect 5802 1444 5814 1736
rect 5802 1436 5804 1444
rect 5812 1436 5814 1444
rect 5802 1434 5814 1436
rect 5834 1444 5846 1446
rect 5834 1436 5836 1444
rect 5844 1436 5846 1444
rect 5770 1356 5772 1364
rect 5780 1356 5782 1364
rect 5770 1354 5782 1356
rect 5738 1096 5740 1104
rect 5748 1096 5750 1104
rect 5738 1094 5750 1096
rect 5770 1064 5782 1066
rect 5770 1056 5772 1064
rect 5780 1056 5782 1064
rect 5770 844 5782 1056
rect 5834 1064 5846 1436
rect 5866 1444 5878 2636
rect 5898 2384 5910 3056
rect 5930 2904 5942 4236
rect 5994 4204 6006 4206
rect 5994 4196 5996 4204
rect 6004 4196 6006 4204
rect 5994 3904 6006 4196
rect 6026 4084 6038 4296
rect 6026 4076 6028 4084
rect 6036 4076 6038 4084
rect 6026 4074 6038 4076
rect 5994 3896 5996 3904
rect 6004 3896 6006 3904
rect 5994 3894 6006 3896
rect 6058 3844 6070 4576
rect 6090 4144 6102 4146
rect 6090 4136 6092 4144
rect 6100 4136 6102 4144
rect 6090 4104 6102 4136
rect 6090 4096 6092 4104
rect 6100 4096 6102 4104
rect 6090 4094 6102 4096
rect 6058 3836 6060 3844
rect 6068 3836 6070 3844
rect 6058 3834 6070 3836
rect 6090 3904 6102 3906
rect 6090 3896 6092 3904
rect 6100 3896 6102 3904
rect 6090 3804 6102 3896
rect 6090 3796 6092 3804
rect 6100 3796 6102 3804
rect 5994 3744 6006 3746
rect 5994 3736 5996 3744
rect 6004 3736 6006 3744
rect 5962 3684 5974 3686
rect 5962 3676 5964 3684
rect 5972 3676 5974 3684
rect 5962 3424 5974 3676
rect 5994 3464 6006 3736
rect 6058 3744 6070 3746
rect 6058 3736 6060 3744
rect 6068 3736 6070 3744
rect 5994 3456 5996 3464
rect 6004 3456 6006 3464
rect 5994 3454 6006 3456
rect 6026 3464 6038 3466
rect 6026 3456 6028 3464
rect 6036 3456 6038 3464
rect 5962 3416 5964 3424
rect 5972 3416 5974 3424
rect 5962 3414 5974 3416
rect 5930 2896 5932 2904
rect 5940 2896 5942 2904
rect 5930 2894 5942 2896
rect 5962 3324 5974 3326
rect 5962 3316 5964 3324
rect 5972 3316 5974 3324
rect 5898 2376 5900 2384
rect 5908 2376 5910 2384
rect 5898 2374 5910 2376
rect 5962 2084 5974 3316
rect 6026 3184 6038 3456
rect 6026 3176 6028 3184
rect 6036 3176 6038 3184
rect 6026 3174 6038 3176
rect 5994 3124 6006 3126
rect 5994 3116 5996 3124
rect 6004 3116 6006 3124
rect 5994 2924 6006 3116
rect 6058 3124 6070 3736
rect 6090 3564 6102 3796
rect 6090 3556 6092 3564
rect 6100 3556 6102 3564
rect 6090 3554 6102 3556
rect 6122 3744 6134 3746
rect 6122 3736 6124 3744
rect 6132 3736 6134 3744
rect 6122 3464 6134 3736
rect 6122 3456 6124 3464
rect 6132 3456 6134 3464
rect 6122 3454 6134 3456
rect 6154 3364 6166 4676
rect 6282 4324 6294 4326
rect 6282 4316 6284 4324
rect 6292 4316 6294 4324
rect 6186 4144 6198 4146
rect 6186 4136 6188 4144
rect 6196 4136 6198 4144
rect 6186 3704 6198 4136
rect 6186 3696 6188 3704
rect 6196 3696 6198 3704
rect 6186 3694 6198 3696
rect 6218 4044 6230 4046
rect 6218 4036 6220 4044
rect 6228 4036 6230 4044
rect 6218 3624 6230 4036
rect 6218 3616 6220 3624
rect 6228 3616 6230 3624
rect 6218 3614 6230 3616
rect 6186 3604 6198 3606
rect 6186 3596 6188 3604
rect 6196 3596 6198 3604
rect 6186 3524 6198 3596
rect 6186 3516 6188 3524
rect 6196 3516 6198 3524
rect 6186 3514 6198 3516
rect 6218 3524 6230 3526
rect 6218 3516 6220 3524
rect 6228 3516 6230 3524
rect 6154 3356 6156 3364
rect 6164 3356 6166 3364
rect 6154 3354 6166 3356
rect 6186 3424 6198 3426
rect 6186 3416 6188 3424
rect 6196 3416 6198 3424
rect 6058 3116 6060 3124
rect 6068 3116 6070 3124
rect 6058 3114 6070 3116
rect 6122 3224 6134 3226
rect 6122 3216 6124 3224
rect 6132 3216 6134 3224
rect 5994 2916 5996 2924
rect 6004 2916 6006 2924
rect 5994 2914 6006 2916
rect 6122 2764 6134 3216
rect 6186 3124 6198 3416
rect 6186 3116 6188 3124
rect 6196 3116 6198 3124
rect 6186 3114 6198 3116
rect 6122 2756 6124 2764
rect 6132 2756 6134 2764
rect 6122 2754 6134 2756
rect 5962 2076 5964 2084
rect 5972 2076 5974 2084
rect 5962 2074 5974 2076
rect 5994 2664 6006 2666
rect 5994 2656 5996 2664
rect 6004 2656 6006 2664
rect 5962 1904 5974 1906
rect 5962 1896 5964 1904
rect 5972 1896 5974 1904
rect 5962 1886 5974 1896
rect 5898 1874 5974 1886
rect 5898 1864 5910 1874
rect 5898 1856 5900 1864
rect 5908 1856 5910 1864
rect 5898 1854 5910 1856
rect 5962 1624 5974 1626
rect 5962 1616 5964 1624
rect 5972 1616 5974 1624
rect 5866 1436 5868 1444
rect 5876 1436 5878 1444
rect 5866 1434 5878 1436
rect 5898 1604 5910 1606
rect 5898 1596 5900 1604
rect 5908 1596 5910 1604
rect 5866 1404 5878 1406
rect 5866 1396 5868 1404
rect 5876 1396 5878 1404
rect 5866 1344 5878 1396
rect 5866 1336 5868 1344
rect 5876 1336 5878 1344
rect 5866 1334 5878 1336
rect 5834 1056 5836 1064
rect 5844 1056 5846 1064
rect 5834 1054 5846 1056
rect 5770 836 5772 844
rect 5780 836 5782 844
rect 5770 834 5782 836
rect 5674 716 5676 724
rect 5684 716 5686 724
rect 5354 584 5366 586
rect 5354 576 5356 584
rect 5364 576 5366 584
rect 5354 566 5366 576
rect 5674 584 5686 716
rect 5674 576 5676 584
rect 5684 576 5686 584
rect 5674 574 5686 576
rect 5322 564 5366 566
rect 5322 556 5324 564
rect 5332 556 5366 564
rect 5322 554 5366 556
rect 5194 516 5196 524
rect 5204 516 5206 524
rect 5194 514 5206 516
rect 5898 444 5910 1596
rect 5898 436 5900 444
rect 5908 436 5910 444
rect 5898 434 5910 436
rect 5930 1244 5942 1246
rect 5930 1236 5932 1244
rect 5940 1236 5942 1244
rect 4824 406 4828 414
rect 4836 406 4844 414
rect 4852 406 4860 414
rect 4868 406 4872 414
rect 3370 76 3372 84
rect 3380 76 3382 84
rect 3370 74 3382 76
rect 4824 14 4872 406
rect 5322 324 5334 326
rect 5322 316 5324 324
rect 5332 316 5334 324
rect 5322 124 5334 316
rect 5930 204 5942 1236
rect 5962 924 5974 1616
rect 5994 1604 6006 2656
rect 6154 2644 6166 2646
rect 6154 2636 6156 2644
rect 6164 2636 6166 2644
rect 6122 2344 6134 2346
rect 6122 2336 6124 2344
rect 6132 2336 6134 2344
rect 5994 1596 5996 1604
rect 6004 1596 6006 1604
rect 5994 1594 6006 1596
rect 6026 1664 6038 1666
rect 6026 1656 6028 1664
rect 6036 1656 6038 1664
rect 5962 916 5964 924
rect 5972 916 5974 924
rect 5962 914 5974 916
rect 5994 984 6006 986
rect 5994 976 5996 984
rect 6004 976 6006 984
rect 5930 196 5932 204
rect 5940 196 5942 204
rect 5930 194 5942 196
rect 5962 844 5974 846
rect 5962 836 5964 844
rect 5972 836 5974 844
rect 5962 184 5974 836
rect 5994 844 6006 976
rect 5994 836 5996 844
rect 6004 836 6006 844
rect 5994 834 6006 836
rect 5962 176 5964 184
rect 5972 176 5974 184
rect 5962 174 5974 176
rect 6026 164 6038 1656
rect 6090 1564 6102 1566
rect 6090 1556 6092 1564
rect 6100 1556 6102 1564
rect 6058 1504 6070 1506
rect 6058 1496 6060 1504
rect 6068 1496 6070 1504
rect 6058 884 6070 1496
rect 6090 924 6102 1556
rect 6122 1304 6134 2336
rect 6154 1464 6166 2636
rect 6218 2224 6230 3516
rect 6218 2216 6220 2224
rect 6228 2216 6230 2224
rect 6218 2214 6230 2216
rect 6250 2244 6262 2246
rect 6250 2236 6252 2244
rect 6260 2236 6262 2244
rect 6218 2024 6230 2026
rect 6218 2016 6220 2024
rect 6228 2016 6230 2024
rect 6154 1456 6156 1464
rect 6164 1456 6166 1464
rect 6154 1454 6166 1456
rect 6186 2004 6198 2006
rect 6186 1996 6188 2004
rect 6196 1996 6198 2004
rect 6122 1296 6124 1304
rect 6132 1296 6134 1304
rect 6122 1294 6134 1296
rect 6154 1364 6166 1366
rect 6154 1356 6156 1364
rect 6164 1356 6166 1364
rect 6090 916 6092 924
rect 6100 916 6102 924
rect 6090 914 6102 916
rect 6122 1264 6134 1266
rect 6122 1256 6124 1264
rect 6132 1256 6134 1264
rect 6058 876 6060 884
rect 6068 876 6070 884
rect 6058 874 6070 876
rect 6026 156 6028 164
rect 6036 156 6038 164
rect 6026 154 6038 156
rect 6058 744 6070 746
rect 6058 736 6060 744
rect 6068 736 6070 744
rect 5322 116 5324 124
rect 5332 116 5334 124
rect 5322 114 5334 116
rect 6058 84 6070 736
rect 6122 144 6134 1256
rect 6154 1104 6166 1356
rect 6154 1096 6156 1104
rect 6164 1096 6166 1104
rect 6154 1064 6166 1096
rect 6154 1056 6156 1064
rect 6164 1056 6166 1064
rect 6154 1054 6166 1056
rect 6186 1024 6198 1996
rect 6218 1064 6230 2016
rect 6218 1056 6220 1064
rect 6228 1056 6230 1064
rect 6218 1054 6230 1056
rect 6186 1016 6188 1024
rect 6196 1016 6198 1024
rect 6186 1014 6198 1016
rect 6154 1004 6166 1006
rect 6154 996 6156 1004
rect 6164 996 6166 1004
rect 6154 204 6166 996
rect 6250 704 6262 2236
rect 6282 1744 6294 4316
rect 6314 4304 6326 4736
rect 6538 4724 6550 4726
rect 6538 4716 6540 4724
rect 6548 4716 6550 4724
rect 6474 4704 6486 4706
rect 6474 4696 6476 4704
rect 6484 4696 6486 4704
rect 6442 4624 6454 4626
rect 6442 4616 6444 4624
rect 6452 4616 6454 4624
rect 6314 4296 6316 4304
rect 6324 4296 6326 4304
rect 6314 4294 6326 4296
rect 6410 4444 6422 4446
rect 6410 4436 6412 4444
rect 6420 4436 6422 4444
rect 6378 4164 6390 4166
rect 6378 4156 6380 4164
rect 6388 4156 6390 4164
rect 6346 4144 6358 4146
rect 6346 4136 6348 4144
rect 6356 4136 6358 4144
rect 6346 4024 6358 4136
rect 6346 4016 6348 4024
rect 6356 4016 6358 4024
rect 6346 4014 6358 4016
rect 6314 3944 6326 3946
rect 6314 3936 6316 3944
rect 6324 3936 6326 3944
rect 6314 3884 6326 3936
rect 6314 3876 6316 3884
rect 6324 3876 6326 3884
rect 6314 3804 6326 3876
rect 6314 3796 6316 3804
rect 6324 3796 6326 3804
rect 6314 3794 6326 3796
rect 6346 3804 6358 3806
rect 6346 3796 6348 3804
rect 6356 3796 6358 3804
rect 6314 3624 6326 3626
rect 6314 3616 6316 3624
rect 6324 3616 6326 3624
rect 6314 3204 6326 3616
rect 6314 3196 6316 3204
rect 6324 3196 6326 3204
rect 6314 3194 6326 3196
rect 6346 3104 6358 3796
rect 6346 3096 6348 3104
rect 6356 3096 6358 3104
rect 6346 3094 6358 3096
rect 6346 2204 6358 2206
rect 6346 2196 6348 2204
rect 6356 2196 6358 2204
rect 6346 1784 6358 2196
rect 6346 1776 6348 1784
rect 6356 1776 6358 1784
rect 6346 1774 6358 1776
rect 6282 1736 6284 1744
rect 6292 1736 6294 1744
rect 6282 1734 6294 1736
rect 6346 1684 6358 1686
rect 6346 1676 6348 1684
rect 6356 1676 6358 1684
rect 6282 1564 6294 1566
rect 6282 1556 6284 1564
rect 6292 1556 6294 1564
rect 6282 1144 6294 1556
rect 6346 1324 6358 1676
rect 6346 1316 6348 1324
rect 6356 1316 6358 1324
rect 6346 1314 6358 1316
rect 6346 1284 6358 1286
rect 6346 1276 6348 1284
rect 6356 1276 6358 1284
rect 6282 1136 6284 1144
rect 6292 1136 6294 1144
rect 6282 1134 6294 1136
rect 6314 1244 6326 1246
rect 6314 1236 6316 1244
rect 6324 1236 6326 1244
rect 6314 984 6326 1236
rect 6346 1104 6358 1276
rect 6346 1096 6348 1104
rect 6356 1096 6358 1104
rect 6346 1094 6358 1096
rect 6314 976 6316 984
rect 6324 976 6326 984
rect 6250 696 6252 704
rect 6260 696 6262 704
rect 6250 694 6262 696
rect 6282 964 6294 966
rect 6282 956 6284 964
rect 6292 956 6294 964
rect 6250 664 6262 666
rect 6250 656 6252 664
rect 6260 656 6262 664
rect 6250 544 6262 656
rect 6250 536 6252 544
rect 6260 536 6262 544
rect 6250 534 6262 536
rect 6154 196 6156 204
rect 6164 196 6166 204
rect 6154 194 6166 196
rect 6186 464 6198 466
rect 6186 456 6188 464
rect 6196 456 6198 464
rect 6122 136 6124 144
rect 6132 136 6134 144
rect 6122 134 6134 136
rect 6058 76 6060 84
rect 6068 76 6070 84
rect 6058 74 6070 76
rect 6186 84 6198 456
rect 6250 324 6262 326
rect 6250 316 6252 324
rect 6260 316 6262 324
rect 6250 244 6262 316
rect 6250 236 6252 244
rect 6260 236 6262 244
rect 6250 234 6262 236
rect 6282 144 6294 956
rect 6282 136 6284 144
rect 6292 136 6294 144
rect 6282 134 6294 136
rect 6314 104 6326 976
rect 6346 1044 6358 1046
rect 6346 1036 6348 1044
rect 6356 1036 6358 1044
rect 6346 224 6358 1036
rect 6346 216 6348 224
rect 6356 216 6358 224
rect 6346 214 6358 216
rect 6378 124 6390 4156
rect 6410 2204 6422 4436
rect 6442 4284 6454 4616
rect 6442 4276 6444 4284
rect 6452 4276 6454 4284
rect 6442 4274 6454 4276
rect 6442 4184 6454 4186
rect 6442 4176 6444 4184
rect 6452 4176 6454 4184
rect 6442 4024 6454 4176
rect 6442 4016 6444 4024
rect 6452 4016 6454 4024
rect 6442 4014 6454 4016
rect 6442 3884 6454 3886
rect 6442 3876 6444 3884
rect 6452 3876 6454 3884
rect 6442 3804 6454 3876
rect 6442 3796 6444 3804
rect 6452 3796 6454 3804
rect 6442 3794 6454 3796
rect 6442 3764 6454 3766
rect 6442 3756 6444 3764
rect 6452 3756 6454 3764
rect 6442 3644 6454 3756
rect 6442 3636 6444 3644
rect 6452 3636 6454 3644
rect 6442 3634 6454 3636
rect 6442 3404 6454 3406
rect 6442 3396 6444 3404
rect 6452 3396 6454 3404
rect 6442 3224 6454 3396
rect 6442 3216 6444 3224
rect 6452 3216 6454 3224
rect 6442 3214 6454 3216
rect 6410 2196 6412 2204
rect 6420 2196 6422 2204
rect 6410 2194 6422 2196
rect 6442 3144 6454 3146
rect 6442 3136 6444 3144
rect 6452 3136 6454 3144
rect 6442 1504 6454 3136
rect 6474 2444 6486 4696
rect 6506 3804 6518 3806
rect 6506 3796 6508 3804
rect 6516 3796 6518 3804
rect 6506 3764 6518 3796
rect 6506 3756 6508 3764
rect 6516 3756 6518 3764
rect 6506 3754 6518 3756
rect 6506 3544 6518 3546
rect 6506 3536 6508 3544
rect 6516 3536 6518 3544
rect 6506 2724 6518 3536
rect 6506 2716 6508 2724
rect 6516 2716 6518 2724
rect 6506 2714 6518 2716
rect 6474 2436 6476 2444
rect 6484 2436 6486 2444
rect 6474 2434 6486 2436
rect 6506 2144 6518 2146
rect 6506 2136 6508 2144
rect 6516 2136 6518 2144
rect 6474 1824 6486 1826
rect 6474 1816 6476 1824
rect 6484 1816 6486 1824
rect 6474 1644 6486 1816
rect 6506 1824 6518 2136
rect 6538 2084 6550 4716
rect 6570 4264 6582 4756
rect 6602 4664 6614 4666
rect 6602 4656 6604 4664
rect 6612 4656 6614 4664
rect 6602 4584 6614 4656
rect 6602 4576 6604 4584
rect 6612 4576 6614 4584
rect 6602 4574 6614 4576
rect 6634 4584 6646 4586
rect 6634 4576 6636 4584
rect 6644 4576 6646 4584
rect 6570 4256 6572 4264
rect 6580 4256 6582 4264
rect 6570 4254 6582 4256
rect 6602 4544 6614 4546
rect 6602 4536 6604 4544
rect 6612 4536 6614 4544
rect 6602 3944 6614 4536
rect 6602 3936 6604 3944
rect 6612 3936 6614 3944
rect 6602 3934 6614 3936
rect 6602 3904 6614 3906
rect 6602 3896 6604 3904
rect 6612 3896 6614 3904
rect 6570 3804 6582 3806
rect 6570 3796 6572 3804
rect 6580 3796 6582 3804
rect 6570 3584 6582 3796
rect 6602 3744 6614 3896
rect 6602 3736 6604 3744
rect 6612 3736 6614 3744
rect 6602 3734 6614 3736
rect 6570 3576 6572 3584
rect 6580 3576 6582 3584
rect 6570 3574 6582 3576
rect 6570 3504 6582 3506
rect 6570 3496 6572 3504
rect 6580 3496 6582 3504
rect 6570 3404 6582 3496
rect 6570 3396 6572 3404
rect 6580 3396 6582 3404
rect 6570 3394 6582 3396
rect 6602 3344 6614 3346
rect 6602 3336 6604 3344
rect 6612 3336 6614 3344
rect 6538 2076 6540 2084
rect 6548 2076 6550 2084
rect 6538 2074 6550 2076
rect 6570 3324 6582 3326
rect 6570 3316 6572 3324
rect 6580 3316 6582 3324
rect 6506 1816 6508 1824
rect 6516 1816 6518 1824
rect 6506 1814 6518 1816
rect 6474 1636 6476 1644
rect 6484 1636 6486 1644
rect 6474 1634 6486 1636
rect 6506 1744 6518 1746
rect 6506 1736 6508 1744
rect 6516 1736 6518 1744
rect 6442 1496 6444 1504
rect 6452 1496 6454 1504
rect 6442 1494 6454 1496
rect 6474 1604 6486 1606
rect 6474 1596 6476 1604
rect 6484 1596 6486 1604
rect 6410 1284 6422 1286
rect 6410 1276 6412 1284
rect 6420 1276 6422 1284
rect 6410 284 6422 1276
rect 6442 1144 6454 1146
rect 6442 1136 6444 1144
rect 6452 1136 6454 1144
rect 6442 964 6454 1136
rect 6442 956 6444 964
rect 6452 956 6454 964
rect 6442 904 6454 956
rect 6442 896 6444 904
rect 6452 896 6454 904
rect 6442 894 6454 896
rect 6442 864 6454 866
rect 6442 856 6444 864
rect 6452 856 6454 864
rect 6442 384 6454 856
rect 6442 376 6444 384
rect 6452 376 6454 384
rect 6442 374 6454 376
rect 6410 276 6412 284
rect 6420 276 6422 284
rect 6410 274 6422 276
rect 6378 116 6380 124
rect 6388 116 6390 124
rect 6378 114 6390 116
rect 6410 144 6422 146
rect 6410 136 6412 144
rect 6420 136 6422 144
rect 6314 96 6316 104
rect 6324 96 6326 104
rect 6314 94 6326 96
rect 6186 76 6188 84
rect 6196 76 6198 84
rect 6186 74 6198 76
rect 6410 44 6422 136
rect 6474 144 6486 1596
rect 6506 164 6518 1736
rect 6506 156 6508 164
rect 6516 156 6518 164
rect 6506 154 6518 156
rect 6538 1644 6550 1646
rect 6538 1636 6540 1644
rect 6548 1636 6550 1644
rect 6474 136 6476 144
rect 6484 136 6486 144
rect 6474 134 6486 136
rect 6538 104 6550 1636
rect 6570 1024 6582 3316
rect 6602 3184 6614 3336
rect 6602 3176 6604 3184
rect 6612 3176 6614 3184
rect 6602 3174 6614 3176
rect 6570 1016 6572 1024
rect 6580 1016 6582 1024
rect 6570 1014 6582 1016
rect 6602 3144 6614 3146
rect 6602 3136 6604 3144
rect 6612 3136 6614 3144
rect 6570 944 6582 946
rect 6570 936 6572 944
rect 6580 936 6582 944
rect 6570 844 6582 936
rect 6602 924 6614 3136
rect 6602 916 6604 924
rect 6612 916 6614 924
rect 6602 914 6614 916
rect 6570 836 6572 844
rect 6580 836 6582 844
rect 6570 834 6582 836
rect 6602 844 6614 846
rect 6602 836 6604 844
rect 6612 836 6614 844
rect 6570 604 6582 606
rect 6570 596 6572 604
rect 6580 596 6582 604
rect 6570 484 6582 596
rect 6570 476 6572 484
rect 6580 476 6582 484
rect 6570 474 6582 476
rect 6538 96 6540 104
rect 6548 96 6550 104
rect 6538 94 6550 96
rect 6570 444 6582 446
rect 6570 436 6572 444
rect 6580 436 6582 444
rect 6410 36 6412 44
rect 6420 36 6422 44
rect 6410 34 6422 36
rect 6570 24 6582 436
rect 6602 284 6614 836
rect 6634 424 6646 4576
rect 6634 416 6636 424
rect 6644 416 6646 424
rect 6634 414 6646 416
rect 6602 276 6604 284
rect 6612 276 6614 284
rect 6602 274 6614 276
rect 6634 284 6646 286
rect 6634 276 6636 284
rect 6644 276 6646 284
rect 6602 184 6614 186
rect 6602 176 6604 184
rect 6612 176 6614 184
rect 6602 64 6614 176
rect 6634 84 6646 276
rect 6634 76 6636 84
rect 6644 76 6646 84
rect 6634 74 6646 76
rect 6602 56 6604 64
rect 6612 56 6614 64
rect 6602 54 6614 56
rect 6570 16 6572 24
rect 6580 16 6582 24
rect 6570 14 6582 16
rect 4824 6 4828 14
rect 4836 6 4844 14
rect 4852 6 4860 14
rect 4868 6 4872 14
rect 4824 -40 4872 6
use NAND3X1  NAND3X1_165
timestamp 1742918108
transform -1 0 184 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_268
timestamp 1742918108
transform -1 0 120 0 1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_95
timestamp 1742918108
transform -1 0 72 0 1 210
box -4 -6 68 206
use XOR2X1  XOR2X1_14
timestamp 1742918108
transform 1 0 88 0 -1 210
box -4 -6 116 206
use NAND2X1  NAND2X1_269
timestamp 1742918108
transform 1 0 40 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_223
timestamp 1742918108
transform 1 0 8 0 -1 210
box -4 -6 36 206
use NAND3X1  NAND3X1_131
timestamp 1742918108
transform -1 0 312 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_126
timestamp 1742918108
transform -1 0 248 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_87
timestamp 1742918108
transform 1 0 200 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_125
timestamp 1742918108
transform 1 0 312 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_162
timestamp 1742918108
transform -1 0 392 0 -1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_86
timestamp 1742918108
transform -1 0 328 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_128
timestamp 1742918108
transform -1 0 504 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_122
timestamp 1742918108
transform -1 0 440 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_93
timestamp 1742918108
transform 1 0 392 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_124
timestamp 1742918108
transform -1 0 568 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_251
timestamp 1742918108
transform -1 0 568 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_267
timestamp 1742918108
transform 1 0 456 0 -1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_121
timestamp 1742918108
transform -1 0 632 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_250
timestamp 1742918108
transform -1 0 632 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_161
timestamp 1742918108
transform -1 0 696 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_247
timestamp 1742918108
transform -1 0 696 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_117
timestamp 1742918108
transform 1 0 696 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_252
timestamp 1742918108
transform -1 0 760 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_123
timestamp 1742918108
transform 1 0 760 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_253
timestamp 1742918108
transform -1 0 824 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_266
timestamp 1742918108
transform -1 0 936 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_266
timestamp 1742918108
transform -1 0 872 0 1 210
box -4 -6 52 206
use INVX1  INVX1_271
timestamp 1742918108
transform 1 0 888 0 -1 210
box -4 -6 36 206
use AOI21X1  AOI21X1_126
timestamp 1742918108
transform 1 0 824 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_164
timestamp 1742918108
transform -1 0 1000 0 1 210
box -4 -6 68 206
use AOI22X1  AOI22X1_36
timestamp 1742918108
transform -1 0 1064 0 -1 210
box -4 -6 84 206
use NAND3X1  NAND3X1_254
timestamp 1742918108
transform -1 0 984 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_268
timestamp 1742918108
transform -1 0 1096 0 1 210
box -4 -6 68 206
use INVX1  INVX1_222
timestamp 1742918108
transform -1 0 1032 0 1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_354
timestamp 1742918108
transform -1 0 1112 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_264
timestamp 1742918108
transform -1 0 1256 0 1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_92
timestamp 1742918108
transform -1 0 1208 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_247
timestamp 1742918108
transform -1 0 1144 0 1 210
box -4 -6 52 206
use NOR3X1  NOR3X1_10
timestamp 1742918108
transform -1 0 1304 0 -1 210
box -4 -6 132 206
use OR2X2  OR2X2_26
timestamp 1742918108
transform -1 0 1176 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_246
timestamp 1742918108
transform -1 0 1368 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_340
timestamp 1742918108
transform -1 0 1304 0 1 210
box -4 -6 52 206
use NOR3X1  NOR3X1_11
timestamp 1742918108
transform -1 0 1432 0 -1 210
box -4 -6 132 206
use OAI21X1  OAI21X1_316
timestamp 1742918108
transform -1 0 1496 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_248
timestamp 1742918108
transform 1 0 1368 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_328
timestamp 1742918108
transform -1 0 1496 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_262
timestamp 1742918108
transform 1 0 1496 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_322
timestamp 1742918108
transform 1 0 1496 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_217
timestamp 1742918108
transform -1 0 1656 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_125
timestamp 1742918108
transform -1 0 1592 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_132
timestamp 1742918108
transform 1 0 1560 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_222
timestamp 1742918108
transform -1 0 1720 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_327
timestamp 1742918108
transform 1 0 1624 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_223
timestamp 1742918108
transform 1 0 1720 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_261
timestamp 1742918108
transform 1 0 1688 0 -1 210
box -4 -6 68 206
use FILL  FILL_1_0_1
timestamp 1742918108
transform -1 0 1816 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_0
timestamp 1742918108
transform -1 0 1800 0 1 210
box -4 -6 20 206
use NAND3X1  NAND3X1_260
timestamp 1742918108
transform 1 0 1800 0 -1 210
box -4 -6 68 206
use FILL  FILL_0_0_2
timestamp 1742918108
transform 1 0 1784 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1742918108
transform 1 0 1768 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_0
timestamp 1742918108
transform 1 0 1752 0 -1 210
box -4 -6 20 206
use XOR2X1  XOR2X1_19
timestamp 1742918108
transform 1 0 1896 0 1 210
box -4 -6 116 206
use NAND3X1  NAND3X1_220
timestamp 1742918108
transform -1 0 1896 0 1 210
box -4 -6 68 206
use FILL  FILL_1_0_2
timestamp 1742918108
transform -1 0 1832 0 1 210
box -4 -6 20 206
use AOI21X1  AOI21X1_128
timestamp 1742918108
transform 1 0 1928 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_255
timestamp 1742918108
transform -1 0 1928 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_336
timestamp 1742918108
transform -1 0 2056 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_325
timestamp 1742918108
transform 1 0 2024 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_270
timestamp 1742918108
transform -1 0 2024 0 -1 210
box -4 -6 36 206
use AOI21X1  AOI21X1_112
timestamp 1742918108
transform 1 0 2120 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_224
timestamp 1742918108
transform -1 0 2120 0 1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_45
timestamp 1742918108
transform 1 0 2152 0 -1 210
box -4 -6 116 206
use NAND3X1  NAND3X1_256
timestamp 1742918108
transform 1 0 2088 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_357
timestamp 1742918108
transform -1 0 2328 0 1 210
box -4 -6 52 206
use AND2X2  AND2X2_42
timestamp 1742918108
transform -1 0 2280 0 1 210
box -4 -6 68 206
use INVX1  INVX1_263
timestamp 1742918108
transform -1 0 2216 0 1 210
box -4 -6 36 206
use NAND3X1  NAND3X1_264
timestamp 1742918108
transform -1 0 2328 0 -1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_44
timestamp 1742918108
transform 1 0 2328 0 1 210
box -4 -6 116 206
use NAND3X1  NAND3X1_265
timestamp 1742918108
transform -1 0 2456 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_262
timestamp 1742918108
transform -1 0 2392 0 -1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_113
timestamp 1742918108
transform 1 0 2504 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_221
timestamp 1742918108
transform -1 0 2504 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_130
timestamp 1742918108
transform -1 0 2584 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_257
timestamp 1742918108
transform -1 0 2520 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_323
timestamp 1742918108
transform -1 0 2632 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_313
timestamp 1742918108
transform 1 0 2616 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_247
timestamp 1742918108
transform -1 0 2616 0 -1 210
box -4 -6 36 206
use NAND3X1  NAND3X1_225
timestamp 1742918108
transform -1 0 2760 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_131
timestamp 1742918108
transform -1 0 2696 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_235
timestamp 1742918108
transform -1 0 2744 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_228
timestamp 1742918108
transform 1 0 2760 0 1 210
box -4 -6 68 206
use AOI22X1  AOI22X1_41
timestamp 1742918108
transform 1 0 2744 0 -1 210
box -4 -6 84 206
use OAI21X1  OAI21X1_311
timestamp 1742918108
transform -1 0 2888 0 1 210
box -4 -6 68 206
use AOI22X1  AOI22X1_37
timestamp 1742918108
transform 1 0 2824 0 -1 210
box -4 -6 84 206
use OAI21X1  OAI21X1_312
timestamp 1742918108
transform 1 0 2888 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_326
timestamp 1742918108
transform -1 0 3000 0 1 210
box -4 -6 52 206
use AOI22X1  AOI22X1_40
timestamp 1742918108
transform 1 0 2904 0 -1 210
box -4 -6 84 206
use NAND3X1  NAND3X1_227
timestamp 1742918108
transform -1 0 3128 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_117
timestamp 1742918108
transform 1 0 3000 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_332
timestamp 1742918108
transform 1 0 3064 0 -1 210
box -4 -6 68 206
use AOI22X1  AOI22X1_38
timestamp 1742918108
transform 1 0 2984 0 -1 210
box -4 -6 84 206
use NAND3X1  NAND3X1_231
timestamp 1742918108
transform 1 0 3128 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_330
timestamp 1742918108
transform 1 0 3128 0 -1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_129
timestamp 1742918108
transform -1 0 3256 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_263
timestamp 1742918108
transform -1 0 3304 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_360
timestamp 1742918108
transform 1 0 3192 0 -1 210
box -4 -6 52 206
use FILL  FILL_1_1_0
timestamp 1742918108
transform 1 0 3320 0 1 210
box -4 -6 20 206
use NAND3X1  NAND3X1_229
timestamp 1742918108
transform -1 0 3320 0 1 210
box -4 -6 68 206
use FILL  FILL_0_1_1
timestamp 1742918108
transform 1 0 3320 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_0
timestamp 1742918108
transform 1 0 3304 0 -1 210
box -4 -6 20 206
use NAND3X1  NAND3X1_232
timestamp 1742918108
transform 1 0 3368 0 1 210
box -4 -6 68 206
use FILL  FILL_1_1_2
timestamp 1742918108
transform 1 0 3352 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_1
timestamp 1742918108
transform 1 0 3336 0 1 210
box -4 -6 20 206
use NAND3X1  NAND3X1_266
timestamp 1742918108
transform 1 0 3352 0 -1 210
box -4 -6 68 206
use FILL  FILL_0_1_2
timestamp 1742918108
transform 1 0 3336 0 -1 210
box -4 -6 20 206
use NAND3X1  NAND3X1_230
timestamp 1742918108
transform -1 0 3496 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_240
timestamp 1742918108
transform -1 0 3528 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_359
timestamp 1742918108
transform 1 0 3416 0 -1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_236
timestamp 1742918108
transform 1 0 3496 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_237
timestamp 1742918108
transform -1 0 3592 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_233
timestamp 1742918108
transform -1 0 3624 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_241
timestamp 1742918108
transform -1 0 3656 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_246
timestamp 1742918108
transform -1 0 3704 0 1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_318
timestamp 1742918108
transform -1 0 3672 0 1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_115
timestamp 1742918108
transform 1 0 3656 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_329
timestamp 1742918108
transform 1 0 3704 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_116
timestamp 1742918108
transform -1 0 3784 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_188
timestamp 1742918108
transform 1 0 3816 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_358
timestamp 1742918108
transform 1 0 3768 0 1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_133
timestamp 1742918108
transform 1 0 3816 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_265
timestamp 1742918108
transform -1 0 3816 0 -1 210
box -4 -6 36 206
use NAND3X1  NAND3X1_239
timestamp 1742918108
transform 1 0 3864 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_238
timestamp 1742918108
transform -1 0 3944 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_234
timestamp 1742918108
transform 1 0 3928 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_331
timestamp 1742918108
transform -1 0 4008 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_188
timestamp 1742918108
transform 1 0 4136 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_317
timestamp 1742918108
transform 1 0 4088 0 1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_114
timestamp 1742918108
transform -1 0 4088 0 1 210
box -4 -6 68 206
use INVX1  INVX1_264
timestamp 1742918108
transform 1 0 3992 0 1 210
box -4 -6 36 206
use XNOR2X1  XNOR2X1_41
timestamp 1742918108
transform 1 0 4056 0 -1 210
box -4 -6 116 206
use NAND2X1  NAND2X1_338
timestamp 1742918108
transform 1 0 4008 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_312
timestamp 1742918108
transform 1 0 4328 0 1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_195
timestamp 1742918108
transform 1 0 4264 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_190
timestamp 1742918108
transform -1 0 4264 0 1 210
box -4 -6 68 206
use BUFX2  BUFX2_18
timestamp 1742918108
transform -1 0 4264 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_17
timestamp 1742918108
transform -1 0 4216 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_122
timestamp 1742918108
transform -1 0 4456 0 -1 210
box -4 -6 196 206
use BUFX2  BUFX2_19
timestamp 1742918108
transform -1 0 4504 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_123
timestamp 1742918108
transform -1 0 4696 0 -1 210
box -4 -6 196 206
use NAND3X1  NAND3X1_193
timestamp 1742918108
transform -1 0 4440 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_108
timestamp 1742918108
transform 1 0 4440 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_314
timestamp 1742918108
transform 1 0 4504 0 1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_196
timestamp 1742918108
transform 1 0 4552 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_316
timestamp 1742918108
transform -1 0 4664 0 1 210
box -4 -6 52 206
use AOI22X1  AOI22X1_39
timestamp 1742918108
transform -1 0 4744 0 1 210
box -4 -6 84 206
use FILL  FILL_1_2_2
timestamp 1742918108
transform -1 0 4840 0 1 210
box -4 -6 20 206
use FILL  FILL_1_2_1
timestamp 1742918108
transform -1 0 4824 0 1 210
box -4 -6 20 206
use FILL  FILL_1_2_0
timestamp 1742918108
transform -1 0 4808 0 1 210
box -4 -6 20 206
use NAND2X1  NAND2X1_315
timestamp 1742918108
transform 1 0 4744 0 1 210
box -4 -6 52 206
use FILL  FILL_0_2_2
timestamp 1742918108
transform 1 0 4872 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_2_1
timestamp 1742918108
transform 1 0 4856 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_2_0
timestamp 1742918108
transform 1 0 4840 0 -1 210
box -4 -6 20 206
use INVX1  INVX1_138
timestamp 1742918108
transform -1 0 4840 0 -1 210
box -4 -6 36 206
use XNOR2X1  XNOR2X1_18
timestamp 1742918108
transform 1 0 4696 0 -1 210
box -4 -6 116 206
use NAND2X1  NAND2X1_116
timestamp 1742918108
transform -1 0 5080 0 1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_14
timestamp 1742918108
transform 1 0 5032 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_126
timestamp 1742918108
transform -1 0 5032 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_124
timestamp 1742918108
transform -1 0 4984 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_125
timestamp 1742918108
transform 1 0 4888 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_121
timestamp 1742918108
transform -1 0 5032 0 1 210
box -4 -6 196 206
use OAI21X1  OAI21X1_163
timestamp 1742918108
transform 1 0 5224 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_123
timestamp 1742918108
transform -1 0 5224 0 1 210
box -4 -6 52 206
use OR2X2  OR2X2_8
timestamp 1742918108
transform -1 0 5176 0 1 210
box -4 -6 68 206
use INVX1  INVX1_135
timestamp 1742918108
transform 1 0 5080 0 1 210
box -4 -6 36 206
use BUFX2  BUFX2_20
timestamp 1742918108
transform 1 0 5096 0 -1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_41
timestamp 1742918108
transform -1 0 5400 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_118
timestamp 1742918108
transform -1 0 5336 0 1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_129
timestamp 1742918108
transform 1 0 5400 0 1 210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_125
timestamp 1742918108
transform 1 0 5336 0 -1 210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_124
timestamp 1742918108
transform -1 0 5336 0 -1 210
box -4 -6 196 206
use BUFX2  BUFX2_21
timestamp 1742918108
transform 1 0 5528 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_25
timestamp 1742918108
transform 1 0 5576 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_131
timestamp 1742918108
transform -1 0 5672 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_22
timestamp 1742918108
transform -1 0 5720 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_126
timestamp 1742918108
transform -1 0 5912 0 -1 210
box -4 -6 196 206
use INVX1  INVX1_137
timestamp 1742918108
transform 1 0 5592 0 1 210
box -4 -6 36 206
use OR2X2  OR2X2_9
timestamp 1742918108
transform -1 0 5688 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_109
timestamp 1742918108
transform 1 0 5688 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_127
timestamp 1742918108
transform -1 0 5784 0 1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_42
timestamp 1742918108
transform 1 0 5848 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_15
timestamp 1742918108
transform 1 0 5784 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_33
timestamp 1742918108
transform 1 0 5992 0 1 210
box -4 -6 68 206
use INVX1  INVX1_140
timestamp 1742918108
transform 1 0 5960 0 1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_108
timestamp 1742918108
transform 1 0 5912 0 1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_22
timestamp 1742918108
transform -1 0 6024 0 -1 210
box -4 -6 116 206
use NAND2X1  NAND2X1_149
timestamp 1742918108
transform -1 0 6168 0 1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_69
timestamp 1742918108
transform -1 0 6120 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_53
timestamp 1742918108
transform -1 0 6200 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_33
timestamp 1742918108
transform 1 0 6088 0 -1 210
box -4 -6 52 206
use OR2X2  OR2X2_7
timestamp 1742918108
transform 1 0 6024 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_26
timestamp 1742918108
transform 1 0 6200 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_29
timestamp 1742918108
transform 1 0 6248 0 -1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_283
timestamp 1742918108
transform 1 0 6296 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_2
timestamp 1742918108
transform -1 0 6408 0 -1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_46
timestamp 1742918108
transform -1 0 6472 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_398
timestamp 1742918108
transform -1 0 6520 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_130
timestamp 1742918108
transform -1 0 6360 0 1 210
box -4 -6 196 206
use BUFX2  BUFX2_23
timestamp 1742918108
transform -1 0 6408 0 1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_128
timestamp 1742918108
transform -1 0 6600 0 1 210
box -4 -6 196 206
use XNOR2X1  XNOR2X1_30
timestamp 1742918108
transform -1 0 6632 0 -1 210
box -4 -6 116 206
use FILL  FILL_1_1
timestamp 1742918108
transform -1 0 6648 0 -1 210
box -4 -6 20 206
use INVX1  INVX1_133
timestamp 1742918108
transform -1 0 6632 0 1 210
box -4 -6 36 206
use FILL  FILL_2_1
timestamp 1742918108
transform 1 0 6632 0 1 210
box -4 -6 20 206
use XNOR2X1  XNOR2X1_37
timestamp 1742918108
transform 1 0 8 0 -1 610
box -4 -6 116 206
use NAND2X1  NAND2X1_270
timestamp 1742918108
transform -1 0 168 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_225
timestamp 1742918108
transform -1 0 200 0 -1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_272
timestamp 1742918108
transform 1 0 200 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_216
timestamp 1742918108
transform 1 0 248 0 -1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_81
timestamp 1742918108
transform 1 0 280 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_129
timestamp 1742918108
transform 1 0 344 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_127
timestamp 1742918108
transform -1 0 472 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_132
timestamp 1742918108
transform -1 0 536 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_80
timestamp 1742918108
transform -1 0 600 0 -1 610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_34
timestamp 1742918108
transform -1 0 712 0 -1 610
box -4 -6 116 206
use NAND3X1  NAND3X1_119
timestamp 1742918108
transform -1 0 776 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_114
timestamp 1742918108
transform 1 0 776 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_118
timestamp 1742918108
transform 1 0 840 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_111
timestamp 1742918108
transform -1 0 968 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_248
timestamp 1742918108
transform 1 0 968 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_252
timestamp 1742918108
transform -1 0 1080 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_251
timestamp 1742918108
transform -1 0 1144 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_163
timestamp 1742918108
transform -1 0 1208 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_215
timestamp 1742918108
transform -1 0 1240 0 -1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_116
timestamp 1742918108
transform 1 0 1240 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_249
timestamp 1742918108
transform -1 0 1368 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_244
timestamp 1742918108
transform 1 0 1368 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_119
timestamp 1742918108
transform 1 0 1432 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_213
timestamp 1742918108
transform 1 0 1496 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_218
timestamp 1742918108
transform -1 0 1624 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_124
timestamp 1742918108
transform -1 0 1688 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_216
timestamp 1742918108
transform 1 0 1688 0 -1 610
box -4 -6 68 206
use FILL  FILL_2_0_0
timestamp 1742918108
transform -1 0 1768 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1742918108
transform -1 0 1784 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1742918108
transform -1 0 1800 0 -1 610
box -4 -6 20 206
use NAND3X1  NAND3X1_219
timestamp 1742918108
transform -1 0 1864 0 -1 610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_39
timestamp 1742918108
transform 1 0 1864 0 -1 610
box -4 -6 116 206
use INVX1  INVX1_256
timestamp 1742918108
transform -1 0 2008 0 -1 610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_43
timestamp 1742918108
transform 1 0 2008 0 -1 610
box -4 -6 116 206
use XNOR2X1  XNOR2X1_42
timestamp 1742918108
transform 1 0 2120 0 -1 610
box -4 -6 116 206
use INVX1  INVX1_267
timestamp 1742918108
transform -1 0 2264 0 -1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_356
timestamp 1742918108
transform 1 0 2264 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_339
timestamp 1742918108
transform -1 0 2360 0 -1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_259
timestamp 1742918108
transform 1 0 2360 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_355
timestamp 1742918108
transform -1 0 2472 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_326
timestamp 1742918108
transform -1 0 2536 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_258
timestamp 1742918108
transform 1 0 2536 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_249
timestamp 1742918108
transform 1 0 2600 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_324
timestamp 1742918108
transform -1 0 2696 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_310
timestamp 1742918108
transform -1 0 2760 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_337
timestamp 1742918108
transform -1 0 2808 0 -1 610
box -4 -6 52 206
use AOI21X1  AOI21X1_127
timestamp 1742918108
transform -1 0 2872 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_254
timestamp 1742918108
transform -1 0 2904 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_303
timestamp 1742918108
transform -1 0 2968 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_200
timestamp 1742918108
transform 1 0 2968 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_226
timestamp 1742918108
transform 1 0 3032 0 -1 610
box -4 -6 68 206
use OR2X2  OR2X2_24
timestamp 1742918108
transform -1 0 3160 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_194
timestamp 1742918108
transform 1 0 3160 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_248
timestamp 1742918108
transform -1 0 3240 0 -1 610
box -4 -6 36 206
use INVX1  INVX1_245
timestamp 1742918108
transform -1 0 3272 0 -1 610
box -4 -6 36 206
use FILL  FILL_2_1_0
timestamp 1742918108
transform 1 0 3272 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1742918108
transform 1 0 3288 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1742918108
transform 1 0 3304 0 -1 610
box -4 -6 20 206
use AOI22X1  AOI22X1_31
timestamp 1742918108
transform 1 0 3320 0 -1 610
box -4 -6 84 206
use AOI22X1  AOI22X1_30
timestamp 1742918108
transform -1 0 3480 0 -1 610
box -4 -6 84 206
use AOI22X1  AOI22X1_29
timestamp 1742918108
transform 1 0 3480 0 -1 610
box -4 -6 84 206
use AOI22X1  AOI22X1_32
timestamp 1742918108
transform 1 0 3560 0 -1 610
box -4 -6 84 206
use OAI21X1  OAI21X1_298
timestamp 1742918108
transform -1 0 3704 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_294
timestamp 1742918108
transform 1 0 3704 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_296
timestamp 1742918108
transform 1 0 3768 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_293
timestamp 1742918108
transform 1 0 3832 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_295
timestamp 1742918108
transform 1 0 3896 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_192
timestamp 1742918108
transform -1 0 4024 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_189
timestamp 1742918108
transform -1 0 4088 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_191
timestamp 1742918108
transform -1 0 4152 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_292
timestamp 1742918108
transform 1 0 4152 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_235
timestamp 1742918108
transform 1 0 4200 0 -1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_183
timestamp 1742918108
transform -1 0 4296 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_102
timestamp 1742918108
transform -1 0 4360 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_107
timestamp 1742918108
transform -1 0 4424 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_194
timestamp 1742918108
transform 1 0 4424 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_297
timestamp 1742918108
transform -1 0 4552 0 -1 610
box -4 -6 68 206
use XOR2X1  XOR2X1_18
timestamp 1742918108
transform 1 0 4552 0 -1 610
box -4 -6 116 206
use NOR2X1  NOR2X1_102
timestamp 1742918108
transform -1 0 4712 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_103
timestamp 1742918108
transform 1 0 4760 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_187
timestamp 1742918108
transform 1 0 4712 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_104
timestamp 1742918108
transform 1 0 4808 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_162
timestamp 1742918108
transform 1 0 4904 0 -1 610
box -4 -6 68 206
use FILL  FILL_2_2_2
timestamp 1742918108
transform 1 0 4888 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_2_1
timestamp 1742918108
transform 1 0 4872 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_2_0
timestamp 1742918108
transform 1 0 4856 0 -1 610
box -4 -6 20 206
use INVX1  INVX1_134
timestamp 1742918108
transform 1 0 4968 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_165
timestamp 1742918108
transform -1 0 5112 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_105
timestamp 1742918108
transform -1 0 5048 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_164
timestamp 1742918108
transform 1 0 5112 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_168
timestamp 1742918108
transform -1 0 5240 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_119
timestamp 1742918108
transform -1 0 5288 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_136
timestamp 1742918108
transform 1 0 5288 0 -1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_120
timestamp 1742918108
transform -1 0 5368 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_201
timestamp 1742918108
transform 1 0 5368 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_132
timestamp 1742918108
transform 1 0 5416 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_143
timestamp 1742918108
transform -1 0 5496 0 -1 610
box -4 -6 36 206
use OR2X2  OR2X2_11
timestamp 1742918108
transform 1 0 5496 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_16
timestamp 1742918108
transform -1 0 5624 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_17
timestamp 1742918108
transform -1 0 5688 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_43
timestamp 1742918108
transform 1 0 5688 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_174
timestamp 1742918108
transform -1 0 5816 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_185
timestamp 1742918108
transform 1 0 5816 0 -1 610
box -4 -6 68 206
use AOI22X1  AOI22X1_6
timestamp 1742918108
transform -1 0 5960 0 -1 610
box -4 -6 84 206
use OAI21X1  OAI21X1_186
timestamp 1742918108
transform 1 0 5960 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_32
timestamp 1742918108
transform -1 0 6088 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_160
timestamp 1742918108
transform -1 0 6120 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_184
timestamp 1742918108
transform -1 0 6184 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_67
timestamp 1742918108
transform 1 0 6184 0 -1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_127
timestamp 1742918108
transform 1 0 6248 0 -1 610
box -4 -6 196 206
use XNOR2X1  XNOR2X1_24
timestamp 1742918108
transform -1 0 6552 0 -1 610
box -4 -6 116 206
use BUFX2  BUFX2_31
timestamp 1742918108
transform 1 0 6552 0 -1 610
box -4 -6 52 206
use FILL  FILL_3_1
timestamp 1742918108
transform -1 0 6616 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_2
timestamp 1742918108
transform -1 0 6632 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_3
timestamp 1742918108
transform -1 0 6648 0 -1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_272
timestamp 1742918108
transform 1 0 8 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_166
timestamp 1742918108
transform -1 0 136 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_271
timestamp 1742918108
transform 1 0 136 0 1 610
box -4 -6 68 206
use INVX1  INVX1_224
timestamp 1742918108
transform -1 0 232 0 1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_168
timestamp 1742918108
transform 1 0 232 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_271
timestamp 1742918108
transform -1 0 344 0 1 610
box -4 -6 52 206
use AOI21X1  AOI21X1_94
timestamp 1742918108
transform 1 0 344 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_130
timestamp 1742918108
transform -1 0 472 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_136
timestamp 1742918108
transform -1 0 536 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_137
timestamp 1742918108
transform 1 0 536 0 1 610
box -4 -6 68 206
use INVX1  INVX1_217
timestamp 1742918108
transform 1 0 600 0 1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_133
timestamp 1742918108
transform 1 0 632 0 1 610
box -4 -6 68 206
use INVX1  INVX1_212
timestamp 1742918108
transform 1 0 696 0 1 610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_32
timestamp 1742918108
transform -1 0 840 0 1 610
box -4 -6 116 206
use XNOR2X1  XNOR2X1_33
timestamp 1742918108
transform 1 0 840 0 1 610
box -4 -6 116 206
use AOI21X1  AOI21X1_91
timestamp 1742918108
transform 1 0 952 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_265
timestamp 1742918108
transform 1 0 1016 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_265
timestamp 1742918108
transform -1 0 1128 0 1 610
box -4 -6 52 206
use AND2X2  AND2X2_32
timestamp 1742918108
transform 1 0 1128 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_120
timestamp 1742918108
transform 1 0 1192 0 1 610
box -4 -6 68 206
use INVX1  INVX1_214
timestamp 1742918108
transform 1 0 1256 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_259
timestamp 1742918108
transform 1 0 1288 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_159
timestamp 1742918108
transform -1 0 1416 0 1 610
box -4 -6 68 206
use INVX1  INVX1_221
timestamp 1742918108
transform 1 0 1416 0 1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_158
timestamp 1742918108
transform 1 0 1448 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_156
timestamp 1742918108
transform 1 0 1512 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_243
timestamp 1742918108
transform 1 0 1576 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_352
timestamp 1742918108
transform 1 0 1640 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_353
timestamp 1742918108
transform -1 0 1736 0 1 610
box -4 -6 52 206
use FILL  FILL_3_0_0
timestamp 1742918108
transform -1 0 1752 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1742918108
transform -1 0 1768 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1742918108
transform -1 0 1784 0 1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_321
timestamp 1742918108
transform -1 0 1848 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_123
timestamp 1742918108
transform -1 0 1912 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_210
timestamp 1742918108
transform 1 0 1912 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_203
timestamp 1742918108
transform 1 0 1976 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_309
timestamp 1742918108
transform -1 0 2104 0 1 610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_40
timestamp 1742918108
transform -1 0 2216 0 1 610
box -4 -6 116 206
use NAND2X1  NAND2X1_335
timestamp 1742918108
transform 1 0 2216 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_193
timestamp 1742918108
transform -1 0 2312 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_191
timestamp 1742918108
transform 1 0 2312 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_321
timestamp 1742918108
transform -1 0 2408 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_314
timestamp 1742918108
transform 1 0 2408 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_190
timestamp 1742918108
transform -1 0 2520 0 1 610
box -4 -6 52 206
use INVX1  INVX1_266
timestamp 1742918108
transform 1 0 2520 0 1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_118
timestamp 1742918108
transform -1 0 2616 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_315
timestamp 1742918108
transform -1 0 2680 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_300
timestamp 1742918108
transform 1 0 2680 0 1 610
box -4 -6 68 206
use NOR3X1  NOR3X1_8
timestamp 1742918108
transform 1 0 2744 0 1 610
box -4 -6 132 206
use OAI21X1  OAI21X1_301
timestamp 1742918108
transform -1 0 2936 0 1 610
box -4 -6 68 206
use INVX1  INVX1_252
timestamp 1742918108
transform -1 0 2968 0 1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_110
timestamp 1742918108
transform 1 0 2968 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_198
timestamp 1742918108
transform 1 0 3032 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_109
timestamp 1742918108
transform -1 0 3160 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_199
timestamp 1742918108
transform 1 0 3160 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_304
timestamp 1742918108
transform -1 0 3288 0 1 610
box -4 -6 68 206
use FILL  FILL_3_1_0
timestamp 1742918108
transform 1 0 3288 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1742918108
transform 1 0 3304 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1742918108
transform 1 0 3320 0 1 610
box -4 -6 20 206
use NOR3X1  NOR3X1_9
timestamp 1742918108
transform 1 0 3336 0 1 610
box -4 -6 132 206
use NAND2X1  NAND2X1_308
timestamp 1742918108
transform -1 0 3512 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_311
timestamp 1742918108
transform 1 0 3512 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_299
timestamp 1742918108
transform 1 0 3560 0 1 610
box -4 -6 68 206
use INVX2  INVX2_32
timestamp 1742918108
transform -1 0 3656 0 1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_298
timestamp 1742918108
transform 1 0 3656 0 1 610
box -4 -6 52 206
use OR2X2  OR2X2_23
timestamp 1742918108
transform 1 0 3704 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_299
timestamp 1742918108
transform 1 0 3768 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_309
timestamp 1742918108
transform -1 0 3864 0 1 610
box -4 -6 52 206
use INVX1  INVX1_236
timestamp 1742918108
transform -1 0 3896 0 1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_300
timestamp 1742918108
transform 1 0 3896 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_310
timestamp 1742918108
transform -1 0 3992 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_301
timestamp 1742918108
transform 1 0 3992 0 1 610
box -4 -6 52 206
use INVX1  INVX1_239
timestamp 1742918108
transform -1 0 4072 0 1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_179
timestamp 1742918108
transform 1 0 4072 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_289
timestamp 1742918108
transform 1 0 4120 0 1 610
box -4 -6 52 206
use INVX1  INVX1_234
timestamp 1742918108
transform 1 0 4168 0 1 610
box -4 -6 36 206
use AND2X2  AND2X2_35
timestamp 1742918108
transform 1 0 4200 0 1 610
box -4 -6 68 206
use INVX1  INVX1_244
timestamp 1742918108
transform 1 0 4264 0 1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_106
timestamp 1742918108
transform -1 0 4360 0 1 610
box -4 -6 68 206
use AND2X2  AND2X2_34
timestamp 1742918108
transform 1 0 4360 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_291
timestamp 1742918108
transform 1 0 4424 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_286
timestamp 1742918108
transform -1 0 4536 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_294
timestamp 1742918108
transform -1 0 4584 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_285
timestamp 1742918108
transform 1 0 4584 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_295
timestamp 1742918108
transform -1 0 4696 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_290
timestamp 1742918108
transform 1 0 4696 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_293
timestamp 1742918108
transform 1 0 4744 0 1 610
box -4 -6 52 206
use AOI21X1  AOI21X1_103
timestamp 1742918108
transform -1 0 4856 0 1 610
box -4 -6 68 206
use FILL  FILL_3_2_0
timestamp 1742918108
transform 1 0 4856 0 1 610
box -4 -6 20 206
use FILL  FILL_3_2_1
timestamp 1742918108
transform 1 0 4872 0 1 610
box -4 -6 20 206
use FILL  FILL_3_2_2
timestamp 1742918108
transform 1 0 4888 0 1 610
box -4 -6 20 206
use NAND3X1  NAND3X1_182
timestamp 1742918108
transform 1 0 4904 0 1 610
box -4 -6 68 206
use INVX1  INVX1_230
timestamp 1742918108
transform -1 0 5000 0 1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_184
timestamp 1742918108
transform 1 0 5000 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_313
timestamp 1742918108
transform -1 0 5112 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_101
timestamp 1742918108
transform 1 0 5112 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_121
timestamp 1742918108
transform -1 0 5208 0 1 610
box -4 -6 52 206
use INVX2  INVX2_8
timestamp 1742918108
transform -1 0 5240 0 1 610
box -4 -6 36 206
use INVX2  INVX2_9
timestamp 1742918108
transform -1 0 5272 0 1 610
box -4 -6 36 206
use INVX1  INVX1_142
timestamp 1742918108
transform 1 0 5272 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_171
timestamp 1742918108
transform 1 0 5304 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_111
timestamp 1742918108
transform -1 0 5416 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_172
timestamp 1742918108
transform 1 0 5416 0 1 610
box -4 -6 68 206
use AND2X2  AND2X2_19
timestamp 1742918108
transform 1 0 5480 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_117
timestamp 1742918108
transform 1 0 5544 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_173
timestamp 1742918108
transform 1 0 5592 0 1 610
box -4 -6 68 206
use OR2X2  OR2X2_10
timestamp 1742918108
transform 1 0 5656 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_133
timestamp 1742918108
transform -1 0 5768 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_134
timestamp 1742918108
transform -1 0 5816 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_112
timestamp 1742918108
transform -1 0 5864 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_117
timestamp 1742918108
transform 1 0 5864 0 1 610
box -4 -6 52 206
use INVX2  INVX2_11
timestamp 1742918108
transform -1 0 5944 0 1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_31
timestamp 1742918108
transform -1 0 6008 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_51
timestamp 1742918108
transform -1 0 6072 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_30
timestamp 1742918108
transform -1 0 6136 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_52
timestamp 1742918108
transform -1 0 6200 0 1 610
box -4 -6 68 206
use NOR3X1  NOR3X1_6
timestamp 1742918108
transform 1 0 6200 0 1 610
box -4 -6 132 206
use OAI21X1  OAI21X1_215
timestamp 1742918108
transform 1 0 6328 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_68
timestamp 1742918108
transform -1 0 6456 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_51
timestamp 1742918108
transform 1 0 6456 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_189
timestamp 1742918108
transform 1 0 6520 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_168
timestamp 1742918108
transform -1 0 6616 0 1 610
box -4 -6 52 206
use FILL  FILL_4_1
timestamp 1742918108
transform 1 0 6616 0 1 610
box -4 -6 20 206
use FILL  FILL_4_2
timestamp 1742918108
transform 1 0 6632 0 1 610
box -4 -6 20 206
use AOI21X1  AOI21X1_99
timestamp 1742918108
transform 1 0 8 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_85
timestamp 1742918108
transform -1 0 136 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_134
timestamp 1742918108
transform -1 0 200 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_140
timestamp 1742918108
transform -1 0 264 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_270
timestamp 1742918108
transform -1 0 328 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_255
timestamp 1742918108
transform -1 0 392 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_138
timestamp 1742918108
transform 1 0 392 0 -1 1010
box -4 -6 68 206
use INVX2  INVX2_26
timestamp 1742918108
transform -1 0 488 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_249
timestamp 1742918108
transform 1 0 488 0 -1 1010
box -4 -6 68 206
use OAI22X1  OAI22X1_18
timestamp 1742918108
transform 1 0 552 0 -1 1010
box -4 -6 84 206
use AOI22X1  AOI22X1_25
timestamp 1742918108
transform 1 0 632 0 -1 1010
box -4 -6 84 206
use NAND3X1  NAND3X1_113
timestamp 1742918108
transform 1 0 712 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_110
timestamp 1742918108
transform -1 0 840 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_112
timestamp 1742918108
transform 1 0 840 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_107
timestamp 1742918108
transform 1 0 904 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_262
timestamp 1742918108
transform 1 0 968 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_160
timestamp 1742918108
transform 1 0 1032 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_158
timestamp 1742918108
transform -1 0 1144 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_244
timestamp 1742918108
transform -1 0 1192 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_263
timestamp 1742918108
transform 1 0 1192 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_262
timestamp 1742918108
transform -1 0 1288 0 -1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_157
timestamp 1742918108
transform -1 0 1352 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_261
timestamp 1742918108
transform -1 0 1416 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_263
timestamp 1742918108
transform -1 0 1480 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_157
timestamp 1742918108
transform -1 0 1528 0 -1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_245
timestamp 1742918108
transform -1 0 1592 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_209
timestamp 1742918108
transform 1 0 1592 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_214
timestamp 1742918108
transform -1 0 1720 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_212
timestamp 1742918108
transform 1 0 1720 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_0_0
timestamp 1742918108
transform 1 0 1784 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_1
timestamp 1742918108
transform 1 0 1800 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_2
timestamp 1742918108
transform 1 0 1816 0 -1 1010
box -4 -6 20 206
use NAND3X1  NAND3X1_215
timestamp 1742918108
transform 1 0 1832 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_259
timestamp 1742918108
transform 1 0 1896 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_206
timestamp 1742918108
transform -1 0 1992 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_211
timestamp 1742918108
transform 1 0 1992 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_205
timestamp 1742918108
transform -1 0 2120 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_202
timestamp 1742918108
transform -1 0 2184 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_257
timestamp 1742918108
transform 1 0 2184 0 -1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_192
timestamp 1742918108
transform 1 0 2216 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_253
timestamp 1742918108
transform -1 0 2296 0 -1 1010
box -4 -6 36 206
use AOI22X1  AOI22X1_33
timestamp 1742918108
transform 1 0 2296 0 -1 1010
box -4 -6 84 206
use OAI21X1  OAI21X1_302
timestamp 1742918108
transform -1 0 2440 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_325
timestamp 1742918108
transform 1 0 2440 0 -1 1010
box -4 -6 52 206
use AOI22X1  AOI22X1_34
timestamp 1742918108
transform -1 0 2568 0 -1 1010
box -4 -6 84 206
use OR2X2  OR2X2_25
timestamp 1742918108
transform -1 0 2632 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_189
timestamp 1742918108
transform 1 0 2632 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_251
timestamp 1742918108
transform 1 0 2680 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_197
timestamp 1742918108
transform 1 0 2712 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_324
timestamp 1742918108
transform 1 0 2776 0 -1 1010
box -4 -6 52 206
use AND2X2  AND2X2_36
timestamp 1742918108
transform 1 0 2824 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_322
timestamp 1742918108
transform -1 0 2936 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_288
timestamp 1742918108
transform 1 0 2936 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_105
timestamp 1742918108
transform -1 0 3064 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_296
timestamp 1742918108
transform 1 0 3064 0 -1 1010
box -4 -6 52 206
use INVX2  INVX2_34
timestamp 1742918108
transform -1 0 3144 0 -1 1010
box -4 -6 36 206
use INVX1  INVX1_237
timestamp 1742918108
transform 1 0 3144 0 -1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_168
timestamp 1742918108
transform -1 0 3224 0 -1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_177
timestamp 1742918108
transform -1 0 3288 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_1_0
timestamp 1742918108
transform -1 0 3304 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_1
timestamp 1742918108
transform -1 0 3320 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_2
timestamp 1742918108
transform -1 0 3336 0 -1 1010
box -4 -6 20 206
use NAND3X1  NAND3X1_187
timestamp 1742918108
transform -1 0 3400 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_228
timestamp 1742918108
transform -1 0 3432 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_186
timestamp 1742918108
transform -1 0 3496 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_240
timestamp 1742918108
transform -1 0 3528 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_287
timestamp 1742918108
transform -1 0 3592 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_178
timestamp 1742918108
transform -1 0 3640 0 -1 1010
box -4 -6 52 206
use XOR2X1  XOR2X1_17
timestamp 1742918108
transform -1 0 3752 0 -1 1010
box -4 -6 116 206
use INVX1  INVX1_233
timestamp 1742918108
transform 1 0 3752 0 -1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_288
timestamp 1742918108
transform 1 0 3784 0 -1 1010
box -4 -6 52 206
use OR2X2  OR2X2_22
timestamp 1742918108
transform 1 0 3832 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_282
timestamp 1742918108
transform -1 0 3960 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_283
timestamp 1742918108
transform 1 0 3960 0 -1 1010
box -4 -6 52 206
use OR2X2  OR2X2_21
timestamp 1742918108
transform 1 0 4008 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_179
timestamp 1742918108
transform -1 0 4136 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_101
timestamp 1742918108
transform 1 0 4136 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_173
timestamp 1742918108
transform 1 0 4200 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_174
timestamp 1742918108
transform -1 0 4296 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_284
timestamp 1742918108
transform 1 0 4296 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_175
timestamp 1742918108
transform 1 0 4344 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_231
timestamp 1742918108
transform -1 0 4424 0 -1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_197
timestamp 1742918108
transform 1 0 4424 0 -1 1010
box -4 -6 52 206
use AND2X2  AND2X2_25
timestamp 1742918108
transform -1 0 4536 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_104
timestamp 1742918108
transform -1 0 4600 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_361
timestamp 1742918108
transform -1 0 4648 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_198
timestamp 1742918108
transform -1 0 4696 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_185
timestamp 1742918108
transform -1 0 4744 0 -1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_58
timestamp 1742918108
transform -1 0 4808 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_182
timestamp 1742918108
transform 1 0 4808 0 -1 1010
box -4 -6 36 206
use FILL  FILL_4_2_0
timestamp 1742918108
transform 1 0 4840 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_2_1
timestamp 1742918108
transform 1 0 4856 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_2_2
timestamp 1742918108
transform 1 0 4872 0 -1 1010
box -4 -6 20 206
use NAND3X1  NAND3X1_57
timestamp 1742918108
transform 1 0 4888 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_207
timestamp 1742918108
transform -1 0 5016 0 -1 1010
box -4 -6 68 206
use OAI22X1  OAI22X1_16
timestamp 1742918108
transform -1 0 5096 0 -1 1010
box -4 -6 84 206
use NOR2X1  NOR2X1_127
timestamp 1742918108
transform -1 0 5144 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_205
timestamp 1742918108
transform -1 0 5208 0 -1 1010
box -4 -6 68 206
use OAI22X1  OAI22X1_17
timestamp 1742918108
transform -1 0 5288 0 -1 1010
box -4 -6 84 206
use NOR2X1  NOR2X1_123
timestamp 1742918108
transform 1 0 5288 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_203
timestamp 1742918108
transform -1 0 5400 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_144
timestamp 1742918108
transform -1 0 5432 0 -1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_119
timestamp 1742918108
transform 1 0 5432 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_191
timestamp 1742918108
transform 1 0 5480 0 -1 1010
box -4 -6 68 206
use AOI22X1  AOI22X1_8
timestamp 1742918108
transform 1 0 5544 0 -1 1010
box -4 -6 84 206
use NAND2X1  NAND2X1_160
timestamp 1742918108
transform -1 0 5672 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_192
timestamp 1742918108
transform -1 0 5736 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_164
timestamp 1742918108
transform 1 0 5736 0 -1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_155
timestamp 1742918108
transform 1 0 5768 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_27
timestamp 1742918108
transform 1 0 5816 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_159
timestamp 1742918108
transform -1 0 5896 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_27
timestamp 1742918108
transform -1 0 5960 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_29
timestamp 1742918108
transform 1 0 5960 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_24
timestamp 1742918108
transform 1 0 6024 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_28
timestamp 1742918108
transform 1 0 6088 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_150
timestamp 1742918108
transform 1 0 6152 0 -1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_72
timestamp 1742918108
transform -1 0 6264 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_74
timestamp 1742918108
transform -1 0 6328 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_75
timestamp 1742918108
transform -1 0 6392 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_216
timestamp 1742918108
transform -1 0 6456 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_185
timestamp 1742918108
transform -1 0 6488 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_73
timestamp 1742918108
transform 1 0 6488 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_60
timestamp 1742918108
transform -1 0 6616 0 -1 1010
box -4 -6 68 206
use FILL  FILL_5_1
timestamp 1742918108
transform -1 0 6632 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_2
timestamp 1742918108
transform -1 0 6648 0 -1 1010
box -4 -6 20 206
use NAND3X1  NAND3X1_167
timestamp 1742918108
transform -1 0 72 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_256
timestamp 1742918108
transform -1 0 136 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_172
timestamp 1742918108
transform 1 0 136 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_169
timestamp 1742918108
transform 1 0 200 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_139
timestamp 1742918108
transform 1 0 264 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_143
timestamp 1742918108
transform 1 0 328 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_238
timestamp 1742918108
transform 1 0 392 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_269
timestamp 1742918108
transform -1 0 504 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_251
timestamp 1742918108
transform 1 0 504 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_254
timestamp 1742918108
transform -1 0 616 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_247
timestamp 1742918108
transform 1 0 616 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_205
timestamp 1742918108
transform -1 0 712 0 1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_242
timestamp 1742918108
transform -1 0 760 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_218
timestamp 1742918108
transform -1 0 808 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_241
timestamp 1742918108
transform -1 0 856 0 1 1010
box -4 -6 52 206
use AOI22X1  AOI22X1_24
timestamp 1742918108
transform -1 0 936 0 1 1010
box -4 -6 84 206
use NAND2X1  NAND2X1_243
timestamp 1742918108
transform -1 0 984 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_240
timestamp 1742918108
transform -1 0 1032 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_250
timestamp 1742918108
transform -1 0 1080 0 1 1010
box -4 -6 52 206
use AND2X2  AND2X2_31
timestamp 1742918108
transform -1 0 1144 0 1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_89
timestamp 1742918108
transform 1 0 1144 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_159
timestamp 1742918108
transform 1 0 1208 0 1 1010
box -4 -6 52 206
use AND2X2  AND2X2_30
timestamp 1742918108
transform -1 0 1320 0 1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_79
timestamp 1742918108
transform -1 0 1384 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_261
timestamp 1742918108
transform 1 0 1384 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_259
timestamp 1742918108
transform 1 0 1432 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_260
timestamp 1742918108
transform -1 0 1528 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_258
timestamp 1742918108
transform -1 0 1576 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_257
timestamp 1742918108
transform -1 0 1624 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_256
timestamp 1742918108
transform -1 0 1672 0 1 1010
box -4 -6 52 206
use AOI21X1  AOI21X1_88
timestamp 1742918108
transform 1 0 1672 0 1 1010
box -4 -6 68 206
use FILL  FILL_5_0_0
timestamp 1742918108
transform -1 0 1752 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_1
timestamp 1742918108
transform -1 0 1768 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_2
timestamp 1742918108
transform -1 0 1784 0 1 1010
box -4 -6 20 206
use AND2X2  AND2X2_41
timestamp 1742918108
transform -1 0 1848 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_345
timestamp 1742918108
transform -1 0 1896 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_242
timestamp 1742918108
transform -1 0 1960 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_268
timestamp 1742918108
transform -1 0 1992 0 1 1010
box -4 -6 36 206
use AND2X2  AND2X2_39
timestamp 1742918108
transform -1 0 2056 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_333
timestamp 1742918108
transform -1 0 2104 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_201
timestamp 1742918108
transform 1 0 2104 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_204
timestamp 1742918108
transform 1 0 2168 0 1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_122
timestamp 1742918108
transform 1 0 2232 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_332
timestamp 1742918108
transform -1 0 2344 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_195
timestamp 1742918108
transform -1 0 2392 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_334
timestamp 1742918108
transform -1 0 2440 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_329
timestamp 1742918108
transform 1 0 2440 0 1 1010
box -4 -6 52 206
use OAI22X1  OAI22X1_20
timestamp 1742918108
transform -1 0 2568 0 1 1010
box -4 -6 84 206
use OAI21X1  OAI21X1_305
timestamp 1742918108
transform 1 0 2568 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_255
timestamp 1742918108
transform -1 0 2664 0 1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_320
timestamp 1742918108
transform -1 0 2712 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_319
timestamp 1742918108
transform 1 0 2712 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_323
timestamp 1742918108
transform 1 0 2760 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_250
timestamp 1742918108
transform -1 0 2840 0 1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_327
timestamp 1742918108
transform -1 0 2888 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_306
timestamp 1742918108
transform 1 0 2888 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_185
timestamp 1742918108
transform 1 0 2936 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_184
timestamp 1742918108
transform 1 0 3000 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_292
timestamp 1742918108
transform -1 0 3112 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_304
timestamp 1742918108
transform -1 0 3160 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_181
timestamp 1742918108
transform 1 0 3160 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_238
timestamp 1742918108
transform -1 0 3240 0 1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_182
timestamp 1742918108
transform -1 0 3288 0 1 1010
box -4 -6 52 206
use FILL  FILL_5_1_0
timestamp 1742918108
transform -1 0 3304 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_1
timestamp 1742918108
transform -1 0 3320 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_2
timestamp 1742918108
transform -1 0 3336 0 1 1010
box -4 -6 20 206
use NOR2X1  NOR2X1_180
timestamp 1742918108
transform -1 0 3384 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_297
timestamp 1742918108
transform -1 0 3432 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_307
timestamp 1742918108
transform 1 0 3432 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_302
timestamp 1742918108
transform 1 0 3480 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_181
timestamp 1742918108
transform -1 0 3592 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_286
timestamp 1742918108
transform 1 0 3592 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_287
timestamp 1742918108
transform 1 0 3640 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_284
timestamp 1742918108
transform -1 0 3752 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_177
timestamp 1742918108
transform 1 0 3752 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_232
timestamp 1742918108
transform -1 0 3832 0 1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_167
timestamp 1742918108
transform 1 0 3832 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_282
timestamp 1742918108
transform 1 0 3880 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_279
timestamp 1742918108
transform 1 0 3928 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_278
timestamp 1742918108
transform -1 0 4040 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_227
timestamp 1742918108
transform -1 0 4072 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_276
timestamp 1742918108
transform 1 0 4072 0 1 1010
box -4 -6 68 206
use INVX2  INVX2_31
timestamp 1742918108
transform -1 0 4168 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_277
timestamp 1742918108
transform -1 0 4232 0 1 1010
box -4 -6 68 206
use AND2X2  AND2X2_33
timestamp 1742918108
transform 1 0 4232 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_226
timestamp 1742918108
transform -1 0 4328 0 1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_176
timestamp 1742918108
transform -1 0 4392 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_172
timestamp 1742918108
transform 1 0 4392 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_59
timestamp 1742918108
transform -1 0 4504 0 1 1010
box -4 -6 68 206
use AOI22X1  AOI22X1_14
timestamp 1742918108
transform -1 0 4584 0 1 1010
box -4 -6 84 206
use NAND2X1  NAND2X1_186
timestamp 1742918108
transform -1 0 4632 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_61
timestamp 1742918108
transform 1 0 4632 0 1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_63
timestamp 1742918108
transform 1 0 4696 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_130
timestamp 1742918108
transform -1 0 4808 0 1 1010
box -4 -6 52 206
use FILL  FILL_5_2_0
timestamp 1742918108
transform -1 0 4824 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_2_1
timestamp 1742918108
transform -1 0 4840 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_2_2
timestamp 1742918108
transform -1 0 4856 0 1 1010
box -4 -6 20 206
use XOR2X1  XOR2X1_11
timestamp 1742918108
transform -1 0 4968 0 1 1010
box -4 -6 116 206
use INVX1  INVX1_163
timestamp 1742918108
transform -1 0 5000 0 1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_124
timestamp 1742918108
transform -1 0 5048 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_181
timestamp 1742918108
transform 1 0 5048 0 1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_128
timestamp 1742918108
transform -1 0 5128 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_126
timestamp 1742918108
transform 1 0 5128 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_129
timestamp 1742918108
transform -1 0 5224 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_206
timestamp 1742918108
transform 1 0 5224 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_204
timestamp 1742918108
transform -1 0 5352 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_180
timestamp 1742918108
transform -1 0 5384 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_189
timestamp 1742918108
transform 1 0 5384 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_159
timestamp 1742918108
transform 1 0 5448 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_157
timestamp 1742918108
transform 1 0 5496 0 1 1010
box -4 -6 52 206
use AOI22X1  AOI22X1_7
timestamp 1742918108
transform 1 0 5544 0 1 1010
box -4 -6 84 206
use OAI21X1  OAI21X1_190
timestamp 1742918108
transform -1 0 5688 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_120
timestamp 1742918108
transform 1 0 5688 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_158
timestamp 1742918108
transform -1 0 5784 0 1 1010
box -4 -6 52 206
use AND2X2  AND2X2_22
timestamp 1742918108
transform -1 0 5848 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_118
timestamp 1742918108
transform 1 0 5848 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_154
timestamp 1742918108
transform -1 0 5944 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_66
timestamp 1742918108
transform -1 0 6008 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_67
timestamp 1742918108
transform 1 0 6008 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_212
timestamp 1742918108
transform -1 0 6136 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_213
timestamp 1742918108
transform -1 0 6200 0 1 1010
box -4 -6 68 206
use AOI22X1  AOI22X1_15
timestamp 1742918108
transform 1 0 6200 0 1 1010
box -4 -6 84 206
use NAND2X1  NAND2X1_188
timestamp 1742918108
transform -1 0 6328 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_70
timestamp 1742918108
transform 1 0 6328 0 1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_66
timestamp 1742918108
transform 1 0 6392 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_214
timestamp 1742918108
transform 1 0 6456 0 1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_59
timestamp 1742918108
transform -1 0 6584 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_32
timestamp 1742918108
transform 1 0 6584 0 1 1010
box -4 -6 52 206
use FILL  FILL_6_1
timestamp 1742918108
transform 1 0 6632 0 1 1010
box -4 -6 20 206
use NAND3X1  NAND3X1_173
timestamp 1742918108
transform -1 0 72 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_98
timestamp 1742918108
transform 1 0 72 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_275
timestamp 1742918108
transform -1 0 184 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_273
timestamp 1742918108
transform -1 0 232 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_144
timestamp 1742918108
transform 1 0 232 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_141
timestamp 1742918108
transform -1 0 360 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_96
timestamp 1742918108
transform 1 0 360 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_106
timestamp 1742918108
transform -1 0 488 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_135
timestamp 1742918108
transform -1 0 552 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_211
timestamp 1742918108
transform -1 0 584 0 -1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_105
timestamp 1742918108
transform 1 0 584 0 -1 1410
box -4 -6 68 206
use INVX2  INVX2_24
timestamp 1742918108
transform -1 0 680 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_248
timestamp 1742918108
transform -1 0 744 0 -1 1410
box -4 -6 68 206
use NOR3X1  NOR3X1_7
timestamp 1742918108
transform 1 0 744 0 -1 1410
box -4 -6 132 206
use NAND2X1  NAND2X1_216
timestamp 1742918108
transform -1 0 920 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_109
timestamp 1742918108
transform 1 0 920 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_108
timestamp 1742918108
transform 1 0 984 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_213
timestamp 1742918108
transform 1 0 1048 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_250
timestamp 1742918108
transform -1 0 1144 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_253
timestamp 1742918108
transform 1 0 1144 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_245
timestamp 1742918108
transform 1 0 1208 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_115
timestamp 1742918108
transform -1 0 1320 0 -1 1410
box -4 -6 68 206
use AND2X2  AND2X2_29
timestamp 1742918108
transform 1 0 1320 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_249
timestamp 1742918108
transform -1 0 1432 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_154
timestamp 1742918108
transform -1 0 1496 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_155
timestamp 1742918108
transform -1 0 1560 0 -1 1410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_36
timestamp 1742918108
transform 1 0 1560 0 -1 1410
box -4 -6 116 206
use NAND2X1  NAND2X1_351
timestamp 1742918108
transform -1 0 1720 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_346
timestamp 1742918108
transform -1 0 1768 0 -1 1410
box -4 -6 52 206
use FILL  FILL_6_0_0
timestamp 1742918108
transform -1 0 1784 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_1
timestamp 1742918108
transform -1 0 1800 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_2
timestamp 1742918108
transform -1 0 1816 0 -1 1410
box -4 -6 20 206
use NAND2X1  NAND2X1_350
timestamp 1742918108
transform -1 0 1864 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_344
timestamp 1742918108
transform -1 0 1912 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_269
timestamp 1742918108
transform -1 0 1944 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_319
timestamp 1742918108
transform -1 0 2008 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_121
timestamp 1742918108
transform -1 0 2072 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_208
timestamp 1742918108
transform -1 0 2136 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_260
timestamp 1742918108
transform -1 0 2168 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_330
timestamp 1742918108
transform -1 0 2216 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_261
timestamp 1742918108
transform 1 0 2216 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_308
timestamp 1742918108
transform 1 0 2248 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_317
timestamp 1742918108
transform -1 0 2376 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_307
timestamp 1742918108
transform -1 0 2440 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_306
timestamp 1742918108
transform 1 0 2440 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_331
timestamp 1742918108
transform -1 0 2552 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_207
timestamp 1742918108
transform -1 0 2616 0 -1 1410
box -4 -6 68 206
use AOI22X1  AOI22X1_35
timestamp 1742918108
transform -1 0 2696 0 -1 1410
box -4 -6 84 206
use INVX1  INVX1_243
timestamp 1742918108
transform 1 0 2696 0 -1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_186
timestamp 1742918108
transform 1 0 2728 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_290
timestamp 1742918108
transform 1 0 2776 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_291
timestamp 1742918108
transform -1 0 2904 0 -1 1410
box -4 -6 68 206
use INVX2  INVX2_33
timestamp 1742918108
transform -1 0 2936 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_303
timestamp 1742918108
transform 1 0 2936 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_241
timestamp 1742918108
transform 1 0 2984 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_289
timestamp 1742918108
transform -1 0 3080 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_183
timestamp 1742918108
transform -1 0 3128 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_176
timestamp 1742918108
transform -1 0 3176 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_180
timestamp 1742918108
transform -1 0 3240 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_283
timestamp 1742918108
transform -1 0 3304 0 -1 1410
box -4 -6 68 206
use FILL  FILL_6_1_0
timestamp 1742918108
transform -1 0 3320 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_1
timestamp 1742918108
transform -1 0 3336 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_2
timestamp 1742918108
transform -1 0 3352 0 -1 1410
box -4 -6 20 206
use NOR2X1  NOR2X1_171
timestamp 1742918108
transform -1 0 3400 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_279
timestamp 1742918108
transform 1 0 3400 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_172
timestamp 1742918108
transform -1 0 3512 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_169
timestamp 1742918108
transform 1 0 3512 0 -1 1410
box -4 -6 52 206
use AOI22X1  AOI22X1_28
timestamp 1742918108
transform 1 0 3560 0 -1 1410
box -4 -6 84 206
use OAI21X1  OAI21X1_280
timestamp 1742918108
transform 1 0 3640 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_280
timestamp 1742918108
transform -1 0 3752 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_229
timestamp 1742918108
transform 1 0 3752 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_281
timestamp 1742918108
transform 1 0 3784 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_178
timestamp 1742918108
transform 1 0 3832 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_281
timestamp 1742918108
transform -1 0 3960 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_170
timestamp 1742918108
transform 1 0 3960 0 -1 1410
box -4 -6 52 206
use INVX2  INVX2_30
timestamp 1742918108
transform 1 0 4008 0 -1 1410
box -4 -6 36 206
use AOI22X1  AOI22X1_11
timestamp 1742918108
transform 1 0 4040 0 -1 1410
box -4 -6 84 206
use NAND2X1  NAND2X1_177
timestamp 1742918108
transform 1 0 4120 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_177
timestamp 1742918108
transform -1 0 4200 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_180
timestamp 1742918108
transform -1 0 4248 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_176
timestamp 1742918108
transform -1 0 4296 0 -1 1410
box -4 -6 52 206
use XOR2X1  XOR2X1_10
timestamp 1742918108
transform 1 0 4296 0 -1 1410
box -4 -6 116 206
use OAI21X1  OAI21X1_202
timestamp 1742918108
transform 1 0 4408 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_208
timestamp 1742918108
transform 1 0 4472 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_56
timestamp 1742918108
transform 1 0 4536 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_60
timestamp 1742918108
transform 1 0 4600 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_122
timestamp 1742918108
transform -1 0 4712 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_164
timestamp 1742918108
transform -1 0 4760 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_165
timestamp 1742918108
transform -1 0 4808 0 -1 1410
box -4 -6 52 206
use FILL  FILL_6_2_0
timestamp 1742918108
transform 1 0 4808 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_2_1
timestamp 1742918108
transform 1 0 4824 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_2_2
timestamp 1742918108
transform 1 0 4840 0 -1 1410
box -4 -6 20 206
use OAI21X1  OAI21X1_199
timestamp 1742918108
transform 1 0 4856 0 -1 1410
box -4 -6 68 206
use AND2X2  AND2X2_23
timestamp 1742918108
transform -1 0 4984 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_167
timestamp 1742918108
transform -1 0 5032 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_166
timestamp 1742918108
transform -1 0 5080 0 -1 1410
box -4 -6 52 206
use OR2X2  OR2X2_13
timestamp 1742918108
transform -1 0 5144 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_125
timestamp 1742918108
transform 1 0 5144 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_168
timestamp 1742918108
transform 1 0 5192 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_156
timestamp 1742918108
transform -1 0 5272 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_110
timestamp 1742918108
transform 1 0 5272 0 -1 1410
box -4 -6 52 206
use AOI22X1  AOI22X1_9
timestamp 1742918108
transform 1 0 5320 0 -1 1410
box -4 -6 84 206
use INVX1  INVX1_166
timestamp 1742918108
transform -1 0 5432 0 -1 1410
box -4 -6 36 206
use INVX1  INVX1_165
timestamp 1742918108
transform 1 0 5432 0 -1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_34
timestamp 1742918108
transform 1 0 5464 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_167
timestamp 1742918108
transform -1 0 5560 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_193
timestamp 1742918108
transform 1 0 5560 0 -1 1410
box -4 -6 68 206
use NOR3X1  NOR3X1_2
timestamp 1742918108
transform 1 0 5624 0 -1 1410
box -4 -6 132 206
use OAI21X1  OAI21X1_209
timestamp 1742918108
transform 1 0 5752 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_53
timestamp 1742918108
transform -1 0 5880 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_211
timestamp 1742918108
transform 1 0 5880 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_184
timestamp 1742918108
transform 1 0 5944 0 -1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_62
timestamp 1742918108
transform -1 0 6040 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_183
timestamp 1742918108
transform -1 0 6072 0 -1 1410
box -4 -6 36 206
use AOI21X1  AOI21X1_64
timestamp 1742918108
transform -1 0 6136 0 -1 1410
box -4 -6 68 206
use NOR3X1  NOR3X1_5
timestamp 1742918108
transform 1 0 6136 0 -1 1410
box -4 -6 132 206
use NAND3X1  NAND3X1_71
timestamp 1742918108
transform 1 0 6264 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_47
timestamp 1742918108
transform 1 0 6328 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_52
timestamp 1742918108
transform -1 0 6456 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_24
timestamp 1742918108
transform -1 0 6504 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_175
timestamp 1742918108
transform -1 0 6536 0 -1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_50
timestamp 1742918108
transform 1 0 6536 0 -1 1410
box -4 -6 68 206
use FILL  FILL_7_1
timestamp 1742918108
transform -1 0 6616 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_2
timestamp 1742918108
transform -1 0 6632 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_3
timestamp 1742918108
transform -1 0 6648 0 -1 1410
box -4 -6 20 206
use NAND3X1  NAND3X1_147
timestamp 1742918108
transform -1 0 72 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_209
timestamp 1742918108
transform 1 0 72 0 1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_142
timestamp 1742918108
transform -1 0 168 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_148
timestamp 1742918108
transform 1 0 168 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_145
timestamp 1742918108
transform -1 0 296 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_97
timestamp 1742918108
transform 1 0 296 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_218
timestamp 1742918108
transform -1 0 392 0 1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_156
timestamp 1742918108
transform 1 0 392 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_239
timestamp 1742918108
transform 1 0 440 0 1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_88
timestamp 1742918108
transform -1 0 552 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_78
timestamp 1742918108
transform -1 0 616 0 1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_149
timestamp 1742918108
transform -1 0 664 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_235
timestamp 1742918108
transform 1 0 664 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_203
timestamp 1742918108
transform -1 0 760 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_258
timestamp 1742918108
transform -1 0 824 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_257
timestamp 1742918108
transform -1 0 888 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_101
timestamp 1742918108
transform -1 0 952 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_245
timestamp 1742918108
transform 1 0 952 0 1 1410
box -4 -6 68 206
use AOI22X1  AOI22X1_23
timestamp 1742918108
transform -1 0 1096 0 1 1410
box -4 -6 84 206
use AOI21X1  AOI21X1_90
timestamp 1742918108
transform -1 0 1160 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_236
timestamp 1742918108
transform -1 0 1208 0 1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_104
timestamp 1742918108
transform -1 0 1272 0 1 1410
box -4 -6 68 206
use AOI22X1  AOI22X1_22
timestamp 1742918108
transform -1 0 1352 0 1 1410
box -4 -6 84 206
use NAND2X1  NAND2X1_235
timestamp 1742918108
transform -1 0 1400 0 1 1410
box -4 -6 52 206
use INVX2  INVX2_25
timestamp 1742918108
transform -1 0 1432 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_246
timestamp 1742918108
transform -1 0 1496 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_244
timestamp 1742918108
transform 1 0 1496 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_246
timestamp 1742918108
transform 1 0 1560 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_260
timestamp 1742918108
transform 1 0 1608 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_253
timestamp 1742918108
transform -1 0 1720 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_348
timestamp 1742918108
transform 1 0 1720 0 1 1410
box -4 -6 52 206
use FILL  FILL_7_0_0
timestamp 1742918108
transform 1 0 1768 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_1
timestamp 1742918108
transform 1 0 1784 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_2
timestamp 1742918108
transform 1 0 1800 0 1 1410
box -4 -6 20 206
use XOR2X1  XOR2X1_15
timestamp 1742918108
transform 1 0 1816 0 1 1410
box -4 -6 116 206
use NAND2X1  NAND2X1_349
timestamp 1742918108
transform 1 0 1928 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_347
timestamp 1742918108
transform -1 0 2024 0 1 1410
box -4 -6 52 206
use AND2X2  AND2X2_40
timestamp 1742918108
transform -1 0 2088 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_343
timestamp 1742918108
transform -1 0 2136 0 1 1410
box -4 -6 52 206
use AOI21X1  AOI21X1_120
timestamp 1742918108
transform -1 0 2200 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_320
timestamp 1742918108
transform -1 0 2264 0 1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_196
timestamp 1742918108
transform -1 0 2312 0 1 1410
box -4 -6 52 206
use AND2X2  AND2X2_37
timestamp 1742918108
transform -1 0 2376 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_258
timestamp 1742918108
transform 1 0 2376 0 1 1410
box -4 -6 36 206
use OR2X2  OR2X2_27
timestamp 1742918108
transform -1 0 2472 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_342
timestamp 1742918108
transform -1 0 2520 0 1 1410
box -4 -6 52 206
use AND2X2  AND2X2_38
timestamp 1742918108
transform -1 0 2584 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_328
timestamp 1742918108
transform -1 0 2632 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_318
timestamp 1742918108
transform -1 0 2696 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_305
timestamp 1742918108
transform 1 0 2696 0 1 1410
box -4 -6 52 206
use AOI21X1  AOI21X1_111
timestamp 1742918108
transform -1 0 2808 0 1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_185
timestamp 1742918108
transform 1 0 2808 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_242
timestamp 1742918108
transform -1 0 2888 0 1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_341
timestamp 1742918108
transform -1 0 2936 0 1 1410
box -4 -6 52 206
use INVX2  INVX2_28
timestamp 1742918108
transform 1 0 2936 0 1 1410
box -4 -6 36 206
use INVX1  INVX1_131
timestamp 1742918108
transform 1 0 2968 0 1 1410
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_4
timestamp 1742918108
transform 1 0 3000 0 1 1410
box -4 -6 196 206
use NAND2X1  NAND2X1_285
timestamp 1742918108
transform -1 0 3240 0 1 1410
box -4 -6 52 206
use INVX2  INVX2_29
timestamp 1742918108
transform -1 0 3272 0 1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_163
timestamp 1742918108
transform -1 0 3320 0 1 1410
box -4 -6 52 206
use FILL  FILL_7_1_0
timestamp 1742918108
transform 1 0 3320 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_1
timestamp 1742918108
transform 1 0 3336 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_2
timestamp 1742918108
transform 1 0 3352 0 1 1410
box -4 -6 20 206
use INVX2  INVX2_27
timestamp 1742918108
transform 1 0 3368 0 1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_278
timestamp 1742918108
transform 1 0 3400 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_166
timestamp 1742918108
transform -1 0 3496 0 1 1410
box -4 -6 52 206
use XNOR2X1  XNOR2X1_38
timestamp 1742918108
transform -1 0 3608 0 1 1410
box -4 -6 116 206
use INVX1  INVX1_176
timestamp 1742918108
transform -1 0 3640 0 1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_178
timestamp 1742918108
transform 1 0 3640 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_174
timestamp 1742918108
transform 1 0 3688 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_179
timestamp 1742918108
transform 1 0 3736 0 1 1410
box -4 -6 52 206
use AOI22X1  AOI22X1_12
timestamp 1742918108
transform 1 0 3784 0 1 1410
box -4 -6 84 206
use NAND2X1  NAND2X1_173
timestamp 1742918108
transform 1 0 3864 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_181
timestamp 1742918108
transform -1 0 3960 0 1 1410
box -4 -6 52 206
use XNOR2X1  XNOR2X1_29
timestamp 1742918108
transform 1 0 3960 0 1 1410
box -4 -6 116 206
use NAND2X1  NAND2X1_183
timestamp 1742918108
transform 1 0 4072 0 1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_55
timestamp 1742918108
transform 1 0 4120 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_179
timestamp 1742918108
transform 1 0 4184 0 1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_184
timestamp 1742918108
transform -1 0 4264 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_178
timestamp 1742918108
transform 1 0 4264 0 1 1410
box -4 -6 36 206
use AOI21X1  AOI21X1_62
timestamp 1742918108
transform -1 0 4360 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_39
timestamp 1742918108
transform -1 0 4424 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_169
timestamp 1742918108
transform 1 0 4424 0 1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_36
timestamp 1742918108
transform -1 0 4536 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_40
timestamp 1742918108
transform -1 0 4600 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_38
timestamp 1742918108
transform 1 0 4600 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_161
timestamp 1742918108
transform 1 0 4664 0 1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_19
timestamp 1742918108
transform 1 0 4712 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_54
timestamp 1742918108
transform 1 0 4776 0 1 1410
box -4 -6 68 206
use FILL  FILL_7_2_0
timestamp 1742918108
transform -1 0 4856 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_2_1
timestamp 1742918108
transform -1 0 4872 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_2_2
timestamp 1742918108
transform -1 0 4888 0 1 1410
box -4 -6 20 206
use NAND3X1  NAND3X1_65
timestamp 1742918108
transform -1 0 4952 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_57
timestamp 1742918108
transform 1 0 4952 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_173
timestamp 1742918108
transform 1 0 5016 0 1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_64
timestamp 1742918108
transform -1 0 5112 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_55
timestamp 1742918108
transform -1 0 5176 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_122
timestamp 1742918108
transform 1 0 5176 0 1 1410
box -4 -6 52 206
use AOI21X1  AOI21X1_58
timestamp 1742918108
transform 1 0 5224 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_170
timestamp 1742918108
transform -1 0 5352 0 1 1410
box -4 -6 68 206
use AOI22X1  AOI22X1_13
timestamp 1742918108
transform 1 0 5352 0 1 1410
box -4 -6 84 206
use NAND3X1  NAND3X1_63
timestamp 1742918108
transform -1 0 5496 0 1 1410
box -4 -6 68 206
use NOR3X1  NOR3X1_4
timestamp 1742918108
transform -1 0 5624 0 1 1410
box -4 -6 132 206
use OAI21X1  OAI21X1_210
timestamp 1742918108
transform 1 0 5624 0 1 1410
box -4 -6 68 206
use NOR3X1  NOR3X1_3
timestamp 1742918108
transform -1 0 5816 0 1 1410
box -4 -6 132 206
use INVX2  INVX2_15
timestamp 1742918108
transform -1 0 5848 0 1 1410
box -4 -6 36 206
use AOI21X1  AOI21X1_56
timestamp 1742918108
transform 1 0 5848 0 1 1410
box -4 -6 68 206
use OAI22X1  OAI22X1_12
timestamp 1742918108
transform -1 0 5992 0 1 1410
box -4 -6 84 206
use OAI22X1  OAI22X1_15
timestamp 1742918108
transform -1 0 6072 0 1 1410
box -4 -6 84 206
use OAI22X1  OAI22X1_14
timestamp 1742918108
transform 1 0 6072 0 1 1410
box -4 -6 84 206
use OAI22X1  OAI22X1_13
timestamp 1742918108
transform -1 0 6232 0 1 1410
box -4 -6 84 206
use NAND3X1  NAND3X1_41
timestamp 1742918108
transform -1 0 6296 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_44
timestamp 1742918108
transform -1 0 6360 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_45
timestamp 1742918108
transform 1 0 6360 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_65
timestamp 1742918108
transform 1 0 6424 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_42
timestamp 1742918108
transform 1 0 6488 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_49
timestamp 1742918108
transform 1 0 6552 0 1 1410
box -4 -6 68 206
use FILL  FILL_8_1
timestamp 1742918108
transform 1 0 6616 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_2
timestamp 1742918108
transform 1 0 6632 0 1 1410
box -4 -6 20 206
use NAND2X1  NAND2X1_274
timestamp 1742918108
transform 1 0 8 0 -1 1810
box -4 -6 52 206
use AOI21X1  AOI21X1_100
timestamp 1742918108
transform 1 0 56 0 -1 1810
box -4 -6 68 206
use OAI22X1  OAI22X1_19
timestamp 1742918108
transform 1 0 120 0 -1 1810
box -4 -6 84 206
use OAI21X1  OAI21X1_275
timestamp 1742918108
transform 1 0 200 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_160
timestamp 1742918108
transform -1 0 312 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_229
timestamp 1742918108
transform -1 0 360 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_208
timestamp 1742918108
transform -1 0 392 0 -1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_153
timestamp 1742918108
transform -1 0 440 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_242
timestamp 1742918108
transform -1 0 504 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_231
timestamp 1742918108
transform -1 0 552 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_223
timestamp 1742918108
transform 1 0 552 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_220
timestamp 1742918108
transform -1 0 648 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_221
timestamp 1742918108
transform -1 0 696 0 -1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_89
timestamp 1742918108
transform 1 0 696 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_202
timestamp 1742918108
transform -1 0 792 0 -1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_87
timestamp 1742918108
transform -1 0 856 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_232
timestamp 1742918108
transform -1 0 920 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_217
timestamp 1742918108
transform 1 0 920 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_148
timestamp 1742918108
transform -1 0 1016 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_198
timestamp 1742918108
transform -1 0 1064 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_264
timestamp 1742918108
transform 1 0 1064 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_100
timestamp 1742918108
transform 1 0 1128 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_210
timestamp 1742918108
transform -1 0 1224 0 -1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_103
timestamp 1742918108
transform -1 0 1288 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_237
timestamp 1742918108
transform -1 0 1336 0 -1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_99
timestamp 1742918108
transform -1 0 1400 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_102
timestamp 1742918108
transform 1 0 1400 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_154
timestamp 1742918108
transform 1 0 1464 0 -1 1810
box -4 -6 52 206
use OR2X2  OR2X2_19
timestamp 1742918108
transform 1 0 1512 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_267
timestamp 1742918108
transform -1 0 1640 0 -1 1810
box -4 -6 68 206
use XOR2X1  XOR2X1_16
timestamp 1742918108
transform 1 0 1640 0 -1 1810
box -4 -6 116 206
use FILL  FILL_8_0_0
timestamp 1742918108
transform -1 0 1768 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_1
timestamp 1742918108
transform -1 0 1784 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_2
timestamp 1742918108
transform -1 0 1800 0 -1 1810
box -4 -6 20 206
use NAND2X1  NAND2X1_255
timestamp 1742918108
transform -1 0 1848 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_12
timestamp 1742918108
transform -1 0 2040 0 -1 1810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_7
timestamp 1742918108
transform 1 0 2040 0 -1 1810
box -4 -6 196 206
use CLKBUF1  CLKBUF1_5
timestamp 1742918108
transform -1 0 2376 0 -1 1810
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_6
timestamp 1742918108
transform -1 0 2568 0 -1 1810
box -4 -6 196 206
use NAND2X1  NAND2X1_114
timestamp 1742918108
transform 1 0 2568 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_157
timestamp 1742918108
transform -1 0 2680 0 -1 1810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_3
timestamp 1742918108
transform -1 0 2872 0 -1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_152
timestamp 1742918108
transform -1 0 2936 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_110
timestamp 1742918108
transform -1 0 2984 0 -1 1810
box -4 -6 52 206
use AOI22X1  AOI22X1_4
timestamp 1742918108
transform 1 0 2984 0 -1 1810
box -4 -6 84 206
use OR2X2  OR2X2_5
timestamp 1742918108
transform -1 0 3128 0 -1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_35
timestamp 1742918108
transform 1 0 3128 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_84
timestamp 1742918108
transform 1 0 3192 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_124
timestamp 1742918108
transform 1 0 3240 0 -1 1810
box -4 -6 68 206
use FILL  FILL_8_1_0
timestamp 1742918108
transform 1 0 3304 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_1
timestamp 1742918108
transform 1 0 3320 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_2
timestamp 1742918108
transform 1 0 3336 0 -1 1810
box -4 -6 20 206
use INVX1  INVX1_120
timestamp 1742918108
transform 1 0 3352 0 -1 1810
box -4 -6 36 206
use AOI21X1  AOI21X1_21
timestamp 1742918108
transform 1 0 3384 0 -1 1810
box -4 -6 68 206
use AOI22X1  AOI22X1_2
timestamp 1742918108
transform -1 0 3528 0 -1 1810
box -4 -6 84 206
use INVX1  INVX1_119
timestamp 1742918108
transform -1 0 3560 0 -1 1810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_28
timestamp 1742918108
transform 1 0 3560 0 -1 1810
box -4 -6 196 206
use CLKBUF1  CLKBUF1_9
timestamp 1742918108
transform -1 0 3896 0 -1 1810
box -4 -6 148 206
use XNOR2X1  XNOR2X1_27
timestamp 1742918108
transform 1 0 3896 0 -1 1810
box -4 -6 116 206
use XOR2X1  XOR2X1_8
timestamp 1742918108
transform 1 0 4008 0 -1 1810
box -4 -6 116 206
use NAND2X1  NAND2X1_182
timestamp 1742918108
transform -1 0 4168 0 -1 1810
box -4 -6 52 206
use OR2X2  OR2X2_14
timestamp 1742918108
transform -1 0 4232 0 -1 1810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_28
timestamp 1742918108
transform -1 0 4344 0 -1 1810
box -4 -6 116 206
use XNOR2X1  XNOR2X1_26
timestamp 1742918108
transform -1 0 4456 0 -1 1810
box -4 -6 116 206
use INVX2  INVX2_13
timestamp 1742918108
transform -1 0 4488 0 -1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_128
timestamp 1742918108
transform 1 0 4488 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_198
timestamp 1742918108
transform -1 0 4600 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_200
timestamp 1742918108
transform 1 0 4600 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_169
timestamp 1742918108
transform -1 0 4696 0 -1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_37
timestamp 1742918108
transform 1 0 4696 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_35
timestamp 1742918108
transform -1 0 4824 0 -1 1810
box -4 -6 68 206
use FILL  FILL_8_2_0
timestamp 1742918108
transform -1 0 4840 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_2_1
timestamp 1742918108
transform -1 0 4856 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_2_2
timestamp 1742918108
transform -1 0 4872 0 -1 1810
box -4 -6 20 206
use INVX1  INVX1_171
timestamp 1742918108
transform -1 0 4904 0 -1 1810
box -4 -6 36 206
use XNOR2X1  XNOR2X1_19
timestamp 1742918108
transform -1 0 5016 0 -1 1810
box -4 -6 116 206
use INVX1  INVX1_172
timestamp 1742918108
transform 1 0 5016 0 -1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_13
timestamp 1742918108
transform -1 0 5112 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_107
timestamp 1742918108
transform 1 0 5112 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_167
timestamp 1742918108
transform -1 0 5224 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_169
timestamp 1742918108
transform -1 0 5288 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_131
timestamp 1742918108
transform 1 0 5288 0 -1 1810
box -4 -6 52 206
use AND2X2  AND2X2_20
timestamp 1742918108
transform 1 0 5336 0 -1 1810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_20
timestamp 1742918108
transform 1 0 5400 0 -1 1810
box -4 -6 116 206
use NAND2X1  NAND2X1_140
timestamp 1742918108
transform 1 0 5512 0 -1 1810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_21
timestamp 1742918108
transform 1 0 5560 0 -1 1810
box -4 -6 116 206
use OR2X2  OR2X2_12
timestamp 1742918108
transform 1 0 5672 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_135
timestamp 1742918108
transform 1 0 5736 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_113
timestamp 1742918108
transform 1 0 5784 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_175
timestamp 1742918108
transform 1 0 5832 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_157
timestamp 1742918108
transform 1 0 5896 0 -1 1810
box -4 -6 36 206
use INVX1  INVX1_158
timestamp 1742918108
transform 1 0 5928 0 -1 1810
box -4 -6 36 206
use AOI21X1  AOI21X1_50
timestamp 1742918108
transform 1 0 5960 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_26
timestamp 1742918108
transform 1 0 6024 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_23
timestamp 1742918108
transform -1 0 6152 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_22
timestamp 1742918108
transform 1 0 6152 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_25
timestamp 1742918108
transform 1 0 6216 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_153
timestamp 1742918108
transform -1 0 6328 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_162
timestamp 1742918108
transform -1 0 6360 0 -1 1810
box -4 -6 36 206
use INVX1  INVX1_174
timestamp 1742918108
transform 1 0 6360 0 -1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_69
timestamp 1742918108
transform -1 0 6456 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_187
timestamp 1742918108
transform -1 0 6504 0 -1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_43
timestamp 1742918108
transform -1 0 6568 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_161
timestamp 1742918108
transform -1 0 6600 0 -1 1810
box -4 -6 36 206
use FILL  FILL_9_1
timestamp 1742918108
transform -1 0 6616 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_2
timestamp 1742918108
transform -1 0 6632 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_3
timestamp 1742918108
transform -1 0 6648 0 -1 1810
box -4 -6 20 206
use NAND3X1  NAND3X1_152
timestamp 1742918108
transform 1 0 8 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_149
timestamp 1742918108
transform -1 0 136 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_151
timestamp 1742918108
transform 1 0 136 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_146
timestamp 1742918108
transform 1 0 200 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_170
timestamp 1742918108
transform -1 0 328 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_174
timestamp 1742918108
transform 1 0 328 0 1 1810
box -4 -6 68 206
use OR2X2  OR2X2_20
timestamp 1742918108
transform -1 0 456 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_273
timestamp 1742918108
transform -1 0 520 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_230
timestamp 1742918108
transform -1 0 568 0 1 1810
box -4 -6 52 206
use AOI22X1  AOI22X1_19
timestamp 1742918108
transform -1 0 648 0 1 1810
box -4 -6 84 206
use AOI22X1  AOI22X1_17
timestamp 1742918108
transform -1 0 728 0 1 1810
box -4 -6 84 206
use INVX1  INVX1_207
timestamp 1742918108
transform -1 0 760 0 1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_219
timestamp 1742918108
transform 1 0 760 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_241
timestamp 1742918108
transform -1 0 872 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_145
timestamp 1742918108
transform 1 0 872 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_201
timestamp 1742918108
transform -1 0 952 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_243
timestamp 1742918108
transform -1 0 1016 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_233
timestamp 1742918108
transform -1 0 1080 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_151
timestamp 1742918108
transform 1 0 1080 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_234
timestamp 1742918108
transform -1 0 1192 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_155
timestamp 1742918108
transform -1 0 1240 0 1 1810
box -4 -6 52 206
use INVX2  INVX2_21
timestamp 1742918108
transform 1 0 1240 0 1 1810
box -4 -6 36 206
use INVX1  INVX1_189
timestamp 1742918108
transform -1 0 1304 0 1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_215
timestamp 1742918108
transform -1 0 1352 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_192
timestamp 1742918108
transform 1 0 1352 0 1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_81
timestamp 1742918108
transform 1 0 1384 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_150
timestamp 1742918108
transform 1 0 1448 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_204
timestamp 1742918108
transform -1 0 1528 0 1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_233
timestamp 1742918108
transform -1 0 1576 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_211
timestamp 1742918108
transform 1 0 1576 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_232
timestamp 1742918108
transform -1 0 1672 0 1 1810
box -4 -6 52 206
use AOI22X1  AOI22X1_21
timestamp 1742918108
transform -1 0 1752 0 1 1810
box -4 -6 84 206
use FILL  FILL_9_0_0
timestamp 1742918108
transform 1 0 1752 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_1
timestamp 1742918108
transform 1 0 1768 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_2
timestamp 1742918108
transform 1 0 1784 0 1 1810
box -4 -6 20 206
use NAND2X1  NAND2X1_234
timestamp 1742918108
transform 1 0 1800 0 1 1810
box -4 -6 52 206
use AND2X2  AND2X2_28
timestamp 1742918108
transform -1 0 1912 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_254
timestamp 1742918108
transform -1 0 1960 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_104
timestamp 1742918108
transform 1 0 1960 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_102
timestamp 1742918108
transform 1 0 1992 0 1 1810
box -4 -6 68 206
use OR2X2  OR2X2_6
timestamp 1742918108
transform 1 0 2056 0 1 1810
box -4 -6 68 206
use AND2X2  AND2X2_18
timestamp 1742918108
transform -1 0 2184 0 1 1810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_1
timestamp 1742918108
transform 1 0 2184 0 1 1810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_75
timestamp 1742918108
transform 1 0 2376 0 1 1810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_76
timestamp 1742918108
transform -1 0 2760 0 1 1810
box -4 -6 196 206
use NOR2X1  NOR2X1_80
timestamp 1742918108
transform 1 0 2760 0 1 1810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_16
timestamp 1742918108
transform 1 0 2808 0 1 1810
box -4 -6 116 206
use INVX1  INVX1_85
timestamp 1742918108
transform 1 0 2920 0 1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_51
timestamp 1742918108
transform -1 0 3000 0 1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_82
timestamp 1742918108
transform -1 0 3048 0 1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_83
timestamp 1742918108
transform -1 0 3096 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_125
timestamp 1742918108
transform 1 0 3096 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_126
timestamp 1742918108
transform -1 0 3224 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_81
timestamp 1742918108
transform -1 0 3272 0 1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_79
timestamp 1742918108
transform -1 0 3320 0 1 1810
box -4 -6 52 206
use FILL  FILL_9_1_0
timestamp 1742918108
transform -1 0 3336 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_1
timestamp 1742918108
transform -1 0 3352 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_2
timestamp 1742918108
transform -1 0 3368 0 1 1810
box -4 -6 20 206
use INVX1  INVX1_56
timestamp 1742918108
transform -1 0 3400 0 1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_36
timestamp 1742918108
transform -1 0 3448 0 1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_60
timestamp 1742918108
transform -1 0 3640 0 1 1810
box -4 -6 196 206
use OAI21X1  OAI21X1_122
timestamp 1742918108
transform 1 0 3640 0 1 1810
box -4 -6 68 206
use AND2X2  AND2X2_14
timestamp 1742918108
transform 1 0 3704 0 1 1810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_77
timestamp 1742918108
transform 1 0 3768 0 1 1810
box -4 -6 196 206
use NOR2X1  NOR2X1_52
timestamp 1742918108
transform 1 0 3960 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_86
timestamp 1742918108
transform -1 0 4040 0 1 1810
box -4 -6 36 206
use XOR2X1  XOR2X1_9
timestamp 1742918108
transform -1 0 4152 0 1 1810
box -4 -6 116 206
use OAI21X1  OAI21X1_123
timestamp 1742918108
transform 1 0 4152 0 1 1810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_27
timestamp 1742918108
transform 1 0 4216 0 1 1810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_107
timestamp 1742918108
transform 1 0 4408 0 1 1810
box -4 -6 196 206
use AND2X2  AND2X2_24
timestamp 1742918108
transform -1 0 4664 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_201
timestamp 1742918108
transform 1 0 4664 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_61
timestamp 1742918108
transform -1 0 4792 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_163
timestamp 1742918108
transform -1 0 4840 0 1 1810
box -4 -6 52 206
use FILL  FILL_9_2_0
timestamp 1742918108
transform -1 0 4856 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_2_1
timestamp 1742918108
transform -1 0 4872 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_2_2
timestamp 1742918108
transform -1 0 4888 0 1 1810
box -4 -6 20 206
use NOR2X1  NOR2X1_121
timestamp 1742918108
transform -1 0 4936 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_196
timestamp 1742918108
transform -1 0 5000 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_195
timestamp 1742918108
transform 1 0 5000 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_129
timestamp 1742918108
transform -1 0 5112 0 1 1810
box -4 -6 52 206
use XOR2X1  XOR2X1_6
timestamp 1742918108
transform 1 0 5112 0 1 1810
box -4 -6 116 206
use INVX1  INVX1_150
timestamp 1742918108
transform 1 0 5224 0 1 1810
box -4 -6 36 206
use INVX1  INVX1_141
timestamp 1742918108
transform 1 0 5256 0 1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_106
timestamp 1742918108
transform 1 0 5288 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_180
timestamp 1742918108
transform 1 0 5336 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_130
timestamp 1742918108
transform -1 0 5448 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_181
timestamp 1742918108
transform 1 0 5448 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_194
timestamp 1742918108
transform -1 0 5576 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_148
timestamp 1742918108
transform 1 0 5576 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_146
timestamp 1742918108
transform -1 0 5672 0 1 1810
box -4 -6 52 206
use INVX1  INVX1_154
timestamp 1742918108
transform 1 0 5672 0 1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_144
timestamp 1742918108
transform 1 0 5704 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_147
timestamp 1742918108
transform 1 0 5752 0 1 1810
box -4 -6 52 206
use AOI21X1  AOI21X1_49
timestamp 1742918108
transform 1 0 5800 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_46
timestamp 1742918108
transform 1 0 5864 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_155
timestamp 1742918108
transform 1 0 5928 0 1 1810
box -4 -6 36 206
use AOI21X1  AOI21X1_48
timestamp 1742918108
transform -1 0 6024 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_45
timestamp 1742918108
transform 1 0 6024 0 1 1810
box -4 -6 68 206
use OAI22X1  OAI22X1_10
timestamp 1742918108
transform -1 0 6168 0 1 1810
box -4 -6 84 206
use INVX1  INVX1_149
timestamp 1742918108
transform -1 0 6200 0 1 1810
box -4 -6 36 206
use OAI22X1  OAI22X1_7
timestamp 1742918108
transform 1 0 6200 0 1 1810
box -4 -6 84 206
use OAI22X1  OAI22X1_9
timestamp 1742918108
transform -1 0 6360 0 1 1810
box -4 -6 84 206
use OAI22X1  OAI22X1_8
timestamp 1742918108
transform -1 0 6440 0 1 1810
box -4 -6 84 206
use NAND3X1  NAND3X1_68
timestamp 1742918108
transform 1 0 6440 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_151
timestamp 1742918108
transform 1 0 6504 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_152
timestamp 1742918108
transform 1 0 6552 0 1 1810
box -4 -6 52 206
use FILL  FILL_10_1
timestamp 1742918108
transform 1 0 6600 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_2
timestamp 1742918108
transform 1 0 6616 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_3
timestamp 1742918108
transform 1 0 6632 0 1 1810
box -4 -6 20 206
use NAND3X1  NAND3X1_153
timestamp 1742918108
transform -1 0 72 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_83
timestamp 1742918108
transform 1 0 72 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_84
timestamp 1742918108
transform 1 0 136 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_171
timestamp 1742918108
transform 1 0 200 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_175
timestamp 1742918108
transform 1 0 264 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_276
timestamp 1742918108
transform 1 0 328 0 -1 2210
box -4 -6 52 206
use AOI22X1  AOI22X1_20
timestamp 1742918108
transform -1 0 456 0 -1 2210
box -4 -6 84 206
use AOI22X1  AOI22X1_18
timestamp 1742918108
transform 1 0 456 0 -1 2210
box -4 -6 84 206
use OR2X2  OR2X2_18
timestamp 1742918108
transform -1 0 600 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_222
timestamp 1742918108
transform -1 0 648 0 -1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_214
timestamp 1742918108
transform -1 0 696 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_199
timestamp 1742918108
transform -1 0 728 0 -1 2210
box -4 -6 36 206
use NAND3X1  NAND3X1_86
timestamp 1742918108
transform 1 0 728 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_213
timestamp 1742918108
transform -1 0 840 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_147
timestamp 1742918108
transform 1 0 840 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_146
timestamp 1742918108
transform -1 0 936 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_200
timestamp 1742918108
transform -1 0 968 0 -1 2210
box -4 -6 36 206
use AOI21X1  AOI21X1_74
timestamp 1742918108
transform 1 0 968 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_231
timestamp 1742918108
transform -1 0 1096 0 -1 2210
box -4 -6 68 206
use INVX2  INVX2_23
timestamp 1742918108
transform 1 0 1096 0 -1 2210
box -4 -6 36 206
use NOR2X1  NOR2X1_139
timestamp 1742918108
transform 1 0 1128 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_230
timestamp 1742918108
transform 1 0 1176 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_224
timestamp 1742918108
transform 1 0 1240 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_82
timestamp 1742918108
transform 1 0 1304 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_200
timestamp 1742918108
transform 1 0 1368 0 -1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_199
timestamp 1742918108
transform -1 0 1464 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_14
timestamp 1742918108
transform -1 0 1656 0 -1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_13
timestamp 1742918108
transform -1 0 1848 0 -1 2210
box -4 -6 196 206
use FILL  FILL_10_0_0
timestamp 1742918108
transform -1 0 1864 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_0_1
timestamp 1742918108
transform -1 0 1880 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_0_2
timestamp 1742918108
transform -1 0 1896 0 -1 2210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_16
timestamp 1742918108
transform -1 0 2088 0 -1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_19
timestamp 1742918108
transform -1 0 2280 0 -1 2210
box -4 -6 196 206
use NAND2X1  NAND2X1_97
timestamp 1742918108
transform 1 0 2280 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_137
timestamp 1742918108
transform -1 0 2392 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_2
timestamp 1742918108
transform 1 0 2392 0 -1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_59
timestamp 1742918108
transform 1 0 2584 0 -1 2210
box -4 -6 196 206
use NOR2X1  NOR2X1_35
timestamp 1742918108
transform 1 0 2776 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_55
timestamp 1742918108
transform 1 0 2824 0 -1 2210
box -4 -6 36 206
use NOR2X1  NOR2X1_50
timestamp 1742918108
transform 1 0 2856 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_76
timestamp 1742918108
transform 1 0 2904 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_84
timestamp 1742918108
transform 1 0 2952 0 -1 2210
box -4 -6 36 206
use NOR2X1  NOR2X1_77
timestamp 1742918108
transform 1 0 2984 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_78
timestamp 1742918108
transform 1 0 3032 0 -1 2210
box -4 -6 52 206
use AOI21X1  AOI21X1_34
timestamp 1742918108
transform 1 0 3080 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_36
timestamp 1742918108
transform -1 0 3208 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_113
timestamp 1742918108
transform -1 0 3256 0 -1 2210
box -4 -6 52 206
use AOI21X1  AOI21X1_22
timestamp 1742918108
transform -1 0 3320 0 -1 2210
box -4 -6 68 206
use FILL  FILL_10_1_0
timestamp 1742918108
transform 1 0 3320 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_1_1
timestamp 1742918108
transform 1 0 3336 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_1_2
timestamp 1742918108
transform 1 0 3352 0 -1 2210
box -4 -6 20 206
use NOR2X1  NOR2X1_85
timestamp 1742918108
transform 1 0 3368 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_5
timestamp 1742918108
transform -1 0 3608 0 -1 2210
box -4 -6 196 206
use NAND2X1  NAND2X1_112
timestamp 1742918108
transform 1 0 3608 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_155
timestamp 1742918108
transform -1 0 3720 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_154
timestamp 1742918108
transform -1 0 3784 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_61
timestamp 1742918108
transform 1 0 3784 0 -1 2210
box -4 -6 196 206
use NAND2X1  NAND2X1_115
timestamp 1742918108
transform 1 0 3976 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_156
timestamp 1742918108
transform 1 0 4024 0 -1 2210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_17
timestamp 1742918108
transform 1 0 4088 0 -1 2210
box -4 -6 116 206
use NAND2X1  NAND2X1_86
timestamp 1742918108
transform -1 0 4248 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_98
timestamp 1742918108
transform 1 0 4248 0 -1 2210
box -4 -6 52 206
use INVX2  INVX2_6
timestamp 1742918108
transform 1 0 4296 0 -1 2210
box -4 -6 36 206
use XNOR2X1  XNOR2X1_14
timestamp 1742918108
transform -1 0 4440 0 -1 2210
box -4 -6 116 206
use OAI21X1  OAI21X1_130
timestamp 1742918108
transform 1 0 4440 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_90
timestamp 1742918108
transform -1 0 4552 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_30
timestamp 1742918108
transform 1 0 4552 0 -1 2210
box -4 -6 196 206
use NAND2X1  NAND2X1_175
timestamp 1742918108
transform -1 0 4792 0 -1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_162
timestamp 1742918108
transform -1 0 4840 0 -1 2210
box -4 -6 52 206
use FILL  FILL_10_2_0
timestamp 1742918108
transform -1 0 4856 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_2_1
timestamp 1742918108
transform -1 0 4872 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_2_2
timestamp 1742918108
transform -1 0 4888 0 -1 2210
box -4 -6 20 206
use INVX2  INVX2_16
timestamp 1742918108
transform -1 0 4920 0 -1 2210
box -4 -6 36 206
use XOR2X1  XOR2X1_7
timestamp 1742918108
transform -1 0 5032 0 -1 2210
box -4 -6 116 206
use XNOR2X1  XNOR2X1_23
timestamp 1742918108
transform -1 0 5144 0 -1 2210
box -4 -6 116 206
use OAI22X1  OAI22X1_11
timestamp 1742918108
transform -1 0 5224 0 -1 2210
box -4 -6 84 206
use INVX1  INVX1_170
timestamp 1742918108
transform 1 0 5224 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_197
timestamp 1742918108
transform -1 0 5320 0 -1 2210
box -4 -6 68 206
use INVX1  INVX1_139
timestamp 1742918108
transform -1 0 5352 0 -1 2210
box -4 -6 36 206
use INVX1  INVX1_153
timestamp 1742918108
transform -1 0 5384 0 -1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_141
timestamp 1742918108
transform -1 0 5432 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_166
timestamp 1742918108
transform 1 0 5432 0 -1 2210
box -4 -6 68 206
use INVX2  INVX2_10
timestamp 1742918108
transform 1 0 5496 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_183
timestamp 1742918108
transform 1 0 5528 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_145
timestamp 1742918108
transform 1 0 5592 0 -1 2210
box -4 -6 52 206
use AND2X2  AND2X2_21
timestamp 1742918108
transform 1 0 5640 0 -1 2210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_6
timestamp 1742918108
transform 1 0 5704 0 -1 2210
box -4 -6 148 206
use OAI21X1  OAI21X1_176
timestamp 1742918108
transform 1 0 5848 0 -1 2210
box -4 -6 68 206
use INVX2  INVX2_12
timestamp 1742918108
transform 1 0 5912 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_188
timestamp 1742918108
transform 1 0 5944 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_137
timestamp 1742918108
transform -1 0 6056 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_146
timestamp 1742918108
transform 1 0 6056 0 -1 2210
box -4 -6 36 206
use NOR2X1  NOR2X1_115
timestamp 1742918108
transform -1 0 6136 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_145
timestamp 1742918108
transform -1 0 6168 0 -1 2210
box -4 -6 36 206
use NAND3X1  NAND3X1_18
timestamp 1742918108
transform 1 0 6168 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_44
timestamp 1742918108
transform -1 0 6296 0 -1 2210
box -4 -6 68 206
use INVX1  INVX1_156
timestamp 1742918108
transform 1 0 6296 0 -1 2210
box -4 -6 36 206
use AOI21X1  AOI21X1_47
timestamp 1742918108
transform 1 0 6328 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_21
timestamp 1742918108
transform 1 0 6392 0 -1 2210
box -4 -6 68 206
use NOR2X1  NOR2X1_114
timestamp 1742918108
transform -1 0 6504 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_187
timestamp 1742918108
transform 1 0 6504 0 -1 2210
box -4 -6 68 206
use INVX2  INVX2_14
timestamp 1742918108
transform 1 0 6568 0 -1 2210
box -4 -6 36 206
use FILL  FILL_11_1
timestamp 1742918108
transform -1 0 6616 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_2
timestamp 1742918108
transform -1 0 6632 0 -1 2210
box -4 -6 20 206
use FILL  FILL_11_3
timestamp 1742918108
transform -1 0 6648 0 -1 2210
box -4 -6 20 206
use NAND2X1  NAND2X1_228
timestamp 1742918108
transform -1 0 56 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_219
timestamp 1742918108
transform 1 0 56 0 1 2210
box -4 -6 36 206
use AOI21X1  AOI21X1_82
timestamp 1742918108
transform -1 0 152 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_90
timestamp 1742918108
transform 1 0 152 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_93
timestamp 1742918108
transform -1 0 280 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_91
timestamp 1742918108
transform 1 0 280 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_94
timestamp 1742918108
transform 1 0 344 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_237
timestamp 1742918108
transform -1 0 472 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_239
timestamp 1742918108
transform 1 0 472 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_236
timestamp 1742918108
transform -1 0 600 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_238
timestamp 1742918108
transform -1 0 664 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_196
timestamp 1742918108
transform 1 0 664 0 1 2210
box -4 -6 36 206
use INVX1  INVX1_195
timestamp 1742918108
transform -1 0 728 0 1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_203
timestamp 1742918108
transform -1 0 776 0 1 2210
box -4 -6 52 206
use OR2X2  OR2X2_17
timestamp 1742918108
transform -1 0 840 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_212
timestamp 1742918108
transform -1 0 888 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_202
timestamp 1742918108
transform 1 0 888 0 1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_144
timestamp 1742918108
transform 1 0 936 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_210
timestamp 1742918108
transform 1 0 984 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_194
timestamp 1742918108
transform -1 0 1064 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_220
timestamp 1742918108
transform 1 0 1064 0 1 2210
box -4 -6 68 206
use INVX2  INVX2_19
timestamp 1742918108
transform 1 0 1128 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_227
timestamp 1742918108
transform 1 0 1160 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_201
timestamp 1742918108
transform -1 0 1272 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_226
timestamp 1742918108
transform -1 0 1336 0 1 2210
box -4 -6 68 206
use NOR2X1  NOR2X1_142
timestamp 1742918108
transform -1 0 1384 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_225
timestamp 1742918108
transform 1 0 1384 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_193
timestamp 1742918108
transform -1 0 1480 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_104
timestamp 1742918108
transform 1 0 1576 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_106
timestamp 1742918108
transform 1 0 1544 0 1 2210
box -4 -6 36 206
use INVX2  INVX2_18
timestamp 1742918108
transform -1 0 1544 0 1 2210
box -4 -6 36 206
use INVX2  INVX2_17
timestamp 1742918108
transform -1 0 1512 0 1 2210
box -4 -6 36 206
use FILL  FILL_11_0_2
timestamp 1742918108
transform -1 0 1784 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_0_1
timestamp 1742918108
transform -1 0 1768 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_0_0
timestamp 1742918108
transform -1 0 1752 0 1 2210
box -4 -6 20 206
use OAI21X1  OAI21X1_103
timestamp 1742918108
transform 1 0 1672 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_105
timestamp 1742918108
transform 1 0 1640 0 1 2210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_15
timestamp 1742918108
transform -1 0 1976 0 1 2210
box -4 -6 196 206
use INVX1  INVX1_107
timestamp 1742918108
transform 1 0 1976 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_105
timestamp 1742918108
transform 1 0 2008 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_108
timestamp 1742918108
transform 1 0 2072 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_106
timestamp 1742918108
transform 1 0 2104 0 1 2210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_10
timestamp 1742918108
transform -1 0 2360 0 1 2210
box -4 -6 196 206
use INVX1  INVX1_102
timestamp 1742918108
transform 1 0 2360 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_100
timestamp 1742918108
transform 1 0 2392 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_150
timestamp 1742918108
transform 1 0 2456 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_109
timestamp 1742918108
transform -1 0 2568 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_107
timestamp 1742918108
transform 1 0 2568 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_149
timestamp 1742918108
transform -1 0 2680 0 1 2210
box -4 -6 68 206
use NOR2X1  NOR2X1_96
timestamp 1742918108
transform -1 0 2728 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_148
timestamp 1742918108
transform -1 0 2792 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_130
timestamp 1742918108
transform -1 0 2824 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_151
timestamp 1742918108
transform 1 0 2824 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_117
timestamp 1742918108
transform 1 0 2888 0 1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_111
timestamp 1742918108
transform -1 0 2968 0 1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_97
timestamp 1742918108
transform 1 0 2968 0 1 2210
box -4 -6 52 206
use AOI21X1  AOI21X1_37
timestamp 1742918108
transform 1 0 3016 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_153
timestamp 1742918108
transform 1 0 3080 0 1 2210
box -4 -6 68 206
use NOR2X1  NOR2X1_75
timestamp 1742918108
transform -1 0 3192 0 1 2210
box -4 -6 52 206
use AOI21X1  AOI21X1_20
timestamp 1742918108
transform 1 0 3192 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_89
timestamp 1742918108
transform 1 0 3256 0 1 2210
box -4 -6 52 206
use FILL  FILL_11_1_0
timestamp 1742918108
transform 1 0 3304 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_1_1
timestamp 1742918108
transform 1 0 3320 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_1_2
timestamp 1742918108
transform 1 0 3336 0 1 2210
box -4 -6 20 206
use OAI21X1  OAI21X1_127
timestamp 1742918108
transform 1 0 3352 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_121
timestamp 1742918108
transform 1 0 3416 0 1 2210
box -4 -6 36 206
use INVX1  INVX1_122
timestamp 1742918108
transform 1 0 3448 0 1 2210
box -4 -6 36 206
use AOI21X1  AOI21X1_23
timestamp 1742918108
transform 1 0 3480 0 1 2210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_8
timestamp 1742918108
transform -1 0 3736 0 1 2210
box -4 -6 196 206
use AND2X2  AND2X2_16
timestamp 1742918108
transform -1 0 3800 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_132
timestamp 1742918108
transform 1 0 3800 0 1 2210
box -4 -6 36 206
use NOR2X1  NOR2X1_37
timestamp 1742918108
transform 1 0 3832 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_57
timestamp 1742918108
transform -1 0 3912 0 1 2210
box -4 -6 36 206
use NOR2X1  NOR2X1_86
timestamp 1742918108
transform -1 0 3960 0 1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_87
timestamp 1742918108
transform 1 0 3960 0 1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_88
timestamp 1742918108
transform -1 0 4056 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_92
timestamp 1742918108
transform 1 0 4056 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_125
timestamp 1742918108
transform 1 0 4104 0 1 2210
box -4 -6 36 206
use AOI21X1  AOI21X1_26
timestamp 1742918108
transform 1 0 4136 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_126
timestamp 1742918108
transform -1 0 4232 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_131
timestamp 1742918108
transform 1 0 4232 0 1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_25
timestamp 1742918108
transform 1 0 4296 0 1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_24
timestamp 1742918108
transform -1 0 4424 0 1 2210
box -4 -6 68 206
use NOR2X1  NOR2X1_89
timestamp 1742918108
transform -1 0 4472 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_123
timestamp 1742918108
transform 1 0 4472 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_128
timestamp 1742918108
transform 1 0 4504 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_129
timestamp 1742918108
transform 1 0 4568 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_88
timestamp 1742918108
transform -1 0 4680 0 1 2210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_29
timestamp 1742918108
transform 1 0 4680 0 1 2210
box -4 -6 196 206
use FILL  FILL_11_2_0
timestamp 1742918108
transform 1 0 4872 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_2_1
timestamp 1742918108
transform 1 0 4888 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_2_2
timestamp 1742918108
transform 1 0 4904 0 1 2210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_31
timestamp 1742918108
transform 1 0 4920 0 1 2210
box -4 -6 196 206
use NAND2X1  NAND2X1_139
timestamp 1742918108
transform 1 0 5112 0 1 2210
box -4 -6 52 206
use AOI22X1  AOI22X1_10
timestamp 1742918108
transform -1 0 5240 0 1 2210
box -4 -6 84 206
use INVX1  INVX1_152
timestamp 1742918108
transform 1 0 5240 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_182
timestamp 1742918108
transform 1 0 5272 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_142
timestamp 1742918108
transform -1 0 5384 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_151
timestamp 1742918108
transform 1 0 5384 0 1 2210
box -4 -6 36 206
use NAND3X1  NAND3X1_20
timestamp 1742918108
transform -1 0 5480 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_143
timestamp 1742918108
transform 1 0 5480 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_3
timestamp 1742918108
transform 1 0 5528 0 1 2210
box -4 -6 52 206
use CLKBUF1  CLKBUF1_11
timestamp 1742918108
transform 1 0 5576 0 1 2210
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_109
timestamp 1742918108
transform 1 0 5720 0 1 2210
box -4 -6 196 206
use NAND2X1  NAND2X1_136
timestamp 1742918108
transform 1 0 5912 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_178
timestamp 1742918108
transform 1 0 5960 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_148
timestamp 1742918108
transform 1 0 6024 0 1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_138
timestamp 1742918108
transform 1 0 6056 0 1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_116
timestamp 1742918108
transform -1 0 6152 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_179
timestamp 1742918108
transform -1 0 6216 0 1 2210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_136
timestamp 1742918108
transform 1 0 6216 0 1 2210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_133
timestamp 1742918108
transform 1 0 6408 0 1 2210
box -4 -6 196 206
use FILL  FILL_12_1
timestamp 1742918108
transform 1 0 6600 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_2
timestamp 1742918108
transform 1 0 6616 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_3
timestamp 1742918108
transform 1 0 6632 0 1 2210
box -4 -6 20 206
use NAND2X1  NAND2X1_252
timestamp 1742918108
transform 1 0 8 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_220
timestamp 1742918108
transform -1 0 88 0 -1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_150
timestamp 1742918108
transform 1 0 88 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_274
timestamp 1742918108
transform -1 0 216 0 -1 2610
box -4 -6 68 206
use AOI22X1  AOI22X1_27
timestamp 1742918108
transform -1 0 296 0 -1 2610
box -4 -6 84 206
use NAND2X1  NAND2X1_225
timestamp 1742918108
transform 1 0 296 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_206
timestamp 1742918108
transform -1 0 376 0 -1 2610
box -4 -6 36 206
use AOI21X1  AOI21X1_75
timestamp 1742918108
transform -1 0 440 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_206
timestamp 1742918108
transform 1 0 440 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_229
timestamp 1742918108
transform -1 0 552 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_208
timestamp 1742918108
transform 1 0 552 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_207
timestamp 1742918108
transform -1 0 648 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_209
timestamp 1742918108
transform 1 0 648 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_204
timestamp 1742918108
transform -1 0 744 0 -1 2610
box -4 -6 52 206
use OR2X2  OR2X2_16
timestamp 1742918108
transform -1 0 808 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_205
timestamp 1742918108
transform 1 0 808 0 -1 2610
box -4 -6 52 206
use XOR2X1  XOR2X1_12
timestamp 1742918108
transform -1 0 968 0 -1 2610
box -4 -6 116 206
use AOI22X1  AOI22X1_16
timestamp 1742918108
transform 1 0 968 0 -1 2610
box -4 -6 84 206
use NOR2X1  NOR2X1_140
timestamp 1742918108
transform -1 0 1096 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_192
timestamp 1742918108
transform -1 0 1144 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_137
timestamp 1742918108
transform -1 0 1192 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_136
timestamp 1742918108
transform 1 0 1192 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_143
timestamp 1742918108
transform -1 0 1288 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_135
timestamp 1742918108
transform -1 0 1336 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_190
timestamp 1742918108
transform 1 0 1336 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_132
timestamp 1742918108
transform 1 0 1384 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_9
timestamp 1742918108
transform -1 0 1624 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_24
timestamp 1742918108
transform -1 0 1816 0 -1 2610
box -4 -6 196 206
use FILL  FILL_12_0_0
timestamp 1742918108
transform -1 0 1832 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_0_1
timestamp 1742918108
transform -1 0 1848 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_0_2
timestamp 1742918108
transform -1 0 1864 0 -1 2610
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_74
timestamp 1742918108
transform -1 0 2056 0 -1 2610
box -4 -6 196 206
use BUFX4  BUFX4_13
timestamp 1742918108
transform 1 0 2056 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_61
timestamp 1742918108
transform 1 0 2120 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_71
timestamp 1742918108
transform -1 0 2200 0 -1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_95
timestamp 1742918108
transform 1 0 2200 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_58
timestamp 1742918108
transform 1 0 2248 0 -1 2610
box -4 -6 196 206
use NAND2X1  NAND2X1_100
timestamp 1742918108
transform 1 0 2440 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_49
timestamp 1742918108
transform 1 0 2488 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_34
timestamp 1742918108
transform 1 0 2536 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_54
timestamp 1742918108
transform 1 0 2584 0 -1 2610
box -4 -6 36 206
use INVX1  INVX1_83
timestamp 1742918108
transform 1 0 2616 0 -1 2610
box -4 -6 36 206
use NOR2X1  NOR2X1_72
timestamp 1742918108
transform -1 0 2696 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_73
timestamp 1742918108
transform 1 0 2696 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_87
timestamp 1742918108
transform 1 0 2744 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_74
timestamp 1742918108
transform 1 0 2792 0 -1 2610
box -4 -6 52 206
use AOI21X1  AOI21X1_33
timestamp 1742918108
transform -1 0 2904 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_121
timestamp 1742918108
transform -1 0 2968 0 -1 2610
box -4 -6 68 206
use INVX2  INVX2_5
timestamp 1742918108
transform -1 0 3000 0 -1 2610
box -4 -6 36 206
use BUFX4  BUFX4_11
timestamp 1742918108
transform -1 0 3064 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_70
timestamp 1742918108
transform 1 0 3064 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_116
timestamp 1742918108
transform 1 0 3112 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_117
timestamp 1742918108
transform 1 0 3176 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_78
timestamp 1742918108
transform -1 0 3288 0 -1 2610
box -4 -6 52 206
use FILL  FILL_12_1_0
timestamp 1742918108
transform 1 0 3288 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_1_1
timestamp 1742918108
transform 1 0 3304 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_1_2
timestamp 1742918108
transform 1 0 3320 0 -1 2610
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_25
timestamp 1742918108
transform 1 0 3336 0 -1 2610
box -4 -6 196 206
use NAND2X1  NAND2X1_84
timestamp 1742918108
transform -1 0 3576 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_92
timestamp 1742918108
transform -1 0 3640 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_94
timestamp 1742918108
transform -1 0 3672 0 -1 2610
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_34
timestamp 1742918108
transform 1 0 3672 0 -1 2610
box -4 -6 196 206
use AOI22X1  AOI22X1_5
timestamp 1742918108
transform 1 0 3864 0 -1 2610
box -4 -6 84 206
use OAI21X1  OAI21X1_160
timestamp 1742918108
transform -1 0 4008 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_161
timestamp 1742918108
transform -1 0 4072 0 -1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_40
timestamp 1742918108
transform -1 0 4136 0 -1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_39
timestamp 1742918108
transform -1 0 4200 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_99
timestamp 1742918108
transform -1 0 4248 0 -1 2610
box -4 -6 52 206
use AND2X2  AND2X2_17
timestamp 1742918108
transform -1 0 4312 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_128
timestamp 1742918108
transform -1 0 4344 0 -1 2610
box -4 -6 36 206
use AOI21X1  AOI21X1_27
timestamp 1742918108
transform -1 0 4408 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_94
timestamp 1742918108
transform 1 0 4408 0 -1 2610
box -4 -6 52 206
use AOI21X1  AOI21X1_28
timestamp 1742918108
transform 1 0 4456 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_132
timestamp 1742918108
transform 1 0 4520 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_159
timestamp 1742918108
transform 1 0 4584 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_158
timestamp 1742918108
transform -1 0 4712 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_92
timestamp 1742918108
transform -1 0 4760 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_133
timestamp 1742918108
transform 1 0 4760 0 -1 2610
box -4 -6 68 206
use FILL  FILL_12_2_0
timestamp 1742918108
transform -1 0 4840 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_2_1
timestamp 1742918108
transform -1 0 4856 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_2_2
timestamp 1742918108
transform -1 0 4872 0 -1 2610
box -4 -6 20 206
use NAND2X1  NAND2X1_91
timestamp 1742918108
transform -1 0 4920 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_171
timestamp 1742918108
transform -1 0 4968 0 -1 2610
box -4 -6 52 206
use XNOR2X1  XNOR2X1_25
timestamp 1742918108
transform -1 0 5080 0 -1 2610
box -4 -6 116 206
use NAND2X1  NAND2X1_170
timestamp 1742918108
transform -1 0 5128 0 -1 2610
box -4 -6 52 206
use AOI21X1  AOI21X1_38
timestamp 1742918108
transform -1 0 5192 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_91
timestamp 1742918108
transform 1 0 5192 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_87
timestamp 1742918108
transform -1 0 5272 0 -1 2610
box -4 -6 36 206
use NOR2X1  NOR2X1_53
timestamp 1742918108
transform -1 0 5320 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_78
timestamp 1742918108
transform -1 0 5512 0 -1 2610
box -4 -6 196 206
use CLKBUF1  CLKBUF1_3
timestamp 1742918108
transform 1 0 5512 0 -1 2610
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_110
timestamp 1742918108
transform 1 0 5656 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_108
timestamp 1742918108
transform 1 0 5848 0 -1 2610
box -4 -6 196 206
use INVX1  INVX1_147
timestamp 1742918108
transform -1 0 6072 0 -1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_177
timestamp 1742918108
transform -1 0 6136 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_164
timestamp 1742918108
transform -1 0 6184 0 -1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_165
timestamp 1742918108
transform 1 0 6184 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_106
timestamp 1742918108
transform 1 0 6232 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_105
timestamp 1742918108
transform 1 0 6424 0 -1 2610
box -4 -6 196 206
use FILL  FILL_13_1
timestamp 1742918108
transform -1 0 6632 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_2
timestamp 1742918108
transform -1 0 6648 0 -1 2610
box -4 -6 20 206
use XNOR2X1  XNOR2X1_35
timestamp 1742918108
transform 1 0 8 0 1 2610
box -4 -6 116 206
use NAND2X1  NAND2X1_227
timestamp 1742918108
transform -1 0 168 0 1 2610
box -4 -6 52 206
use AOI22X1  AOI22X1_26
timestamp 1742918108
transform -1 0 248 0 1 2610
box -4 -6 84 206
use NAND2X1  NAND2X1_226
timestamp 1742918108
transform -1 0 296 0 1 2610
box -4 -6 52 206
use AOI21X1  AOI21X1_77
timestamp 1742918108
transform 1 0 296 0 1 2610
box -4 -6 68 206
use AND2X2  AND2X2_27
timestamp 1742918108
transform -1 0 424 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_152
timestamp 1742918108
transform 1 0 424 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_228
timestamp 1742918108
transform 1 0 472 0 1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_71
timestamp 1742918108
transform -1 0 600 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_84
timestamp 1742918108
transform -1 0 664 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_197
timestamp 1742918108
transform -1 0 696 0 1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_83
timestamp 1742918108
transform 1 0 696 0 1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_72
timestamp 1742918108
transform 1 0 760 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_77
timestamp 1742918108
transform -1 0 888 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_191
timestamp 1742918108
transform 1 0 888 0 1 2610
box -4 -6 52 206
use AND2X2  AND2X2_26
timestamp 1742918108
transform -1 0 1000 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_187
timestamp 1742918108
transform 1 0 1000 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_217
timestamp 1742918108
transform -1 0 1096 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_219
timestamp 1742918108
transform 1 0 1096 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_188
timestamp 1742918108
transform 1 0 1160 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_221
timestamp 1742918108
transform 1 0 1192 0 1 2610
box -4 -6 68 206
use INVX2  INVX2_22
timestamp 1742918108
transform -1 0 1288 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_218
timestamp 1742918108
transform -1 0 1352 0 1 2610
box -4 -6 68 206
use INVX2  INVX2_20
timestamp 1742918108
transform -1 0 1384 0 1 2610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_31
timestamp 1742918108
transform -1 0 1496 0 1 2610
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_11
timestamp 1742918108
transform -1 0 1688 0 1 2610
box -4 -6 196 206
use INVX1  INVX1_103
timestamp 1742918108
transform 1 0 1688 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_101
timestamp 1742918108
transform 1 0 1720 0 1 2610
box -4 -6 68 206
use FILL  FILL_13_0_0
timestamp 1742918108
transform 1 0 1784 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_0_1
timestamp 1742918108
transform 1 0 1800 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_0_2
timestamp 1742918108
transform 1 0 1816 0 1 2610
box -4 -6 20 206
use INVX1  INVX1_129
timestamp 1742918108
transform 1 0 1832 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_142
timestamp 1742918108
transform 1 0 1864 0 1 2610
box -4 -6 68 206
use BUFX4  BUFX4_4
timestamp 1742918108
transform -1 0 1992 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_101
timestamp 1742918108
transform 1 0 1992 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_99
timestamp 1742918108
transform 1 0 2024 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_133
timestamp 1742918108
transform -1 0 2136 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_56
timestamp 1742918108
transform 1 0 2136 0 1 2610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_88
timestamp 1742918108
transform -1 0 2392 0 1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_22
timestamp 1742918108
transform -1 0 2584 0 1 2610
box -4 -6 196 206
use OAI21X1  OAI21X1_140
timestamp 1742918108
transform -1 0 2648 0 1 2610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_15
timestamp 1742918108
transform 1 0 2648 0 1 2610
box -4 -6 116 206
use AOI21X1  AOI21X1_32
timestamp 1742918108
transform 1 0 2760 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_69
timestamp 1742918108
transform -1 0 2872 0 1 2610
box -4 -6 52 206
use BUFX4  BUFX4_9
timestamp 1742918108
transform -1 0 2936 0 1 2610
box -4 -6 68 206
use BUFX4  BUFX4_5
timestamp 1742918108
transform 1 0 2936 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_118
timestamp 1742918108
transform -1 0 3064 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_119
timestamp 1742918108
transform 1 0 3064 0 1 2610
box -4 -6 68 206
use AND2X2  AND2X2_13
timestamp 1742918108
transform 1 0 3128 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_120
timestamp 1742918108
transform 1 0 3192 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_50
timestamp 1742918108
transform -1 0 3320 0 1 2610
box -4 -6 68 206
use FILL  FILL_13_1_0
timestamp 1742918108
transform -1 0 3336 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_1_1
timestamp 1742918108
transform -1 0 3352 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_1_2
timestamp 1742918108
transform -1 0 3368 0 1 2610
box -4 -6 20 206
use INVX1  INVX1_65
timestamp 1742918108
transform -1 0 3400 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_55
timestamp 1742918108
transform 1 0 3400 0 1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_82
timestamp 1742918108
transform -1 0 3640 0 1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_26
timestamp 1742918108
transform 1 0 3640 0 1 2610
box -4 -6 196 206
use BUFX4  BUFX4_10
timestamp 1742918108
transform 1 0 3832 0 1 2610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_63
timestamp 1742918108
transform 1 0 3896 0 1 2610
box -4 -6 196 206
use INVX1  INVX1_59
timestamp 1742918108
transform 1 0 4088 0 1 2610
box -4 -6 36 206
use NOR2X1  NOR2X1_100
timestamp 1742918108
transform -1 0 4168 0 1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_39
timestamp 1742918108
transform 1 0 4168 0 1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_93
timestamp 1742918108
transform -1 0 4264 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_93
timestamp 1742918108
transform 1 0 4264 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_124
timestamp 1742918108
transform 1 0 4312 0 1 2610
box -4 -6 36 206
use AND2X2  AND2X2_15
timestamp 1742918108
transform 1 0 4344 0 1 2610
box -4 -6 68 206
use INVX2  INVX2_7
timestamp 1742918108
transform 1 0 4408 0 1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_134
timestamp 1742918108
transform -1 0 4504 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_94
timestamp 1742918108
transform 1 0 4504 0 1 2610
box -4 -6 52 206
use AOI22X1  AOI22X1_3
timestamp 1742918108
transform -1 0 4632 0 1 2610
box -4 -6 84 206
use INVX1  INVX1_127
timestamp 1742918108
transform -1 0 4664 0 1 2610
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_32
timestamp 1742918108
transform 1 0 4664 0 1 2610
box -4 -6 196 206
use FILL  FILL_13_2_0
timestamp 1742918108
transform 1 0 4856 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_2_1
timestamp 1742918108
transform 1 0 4872 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_2_2
timestamp 1742918108
transform 1 0 4888 0 1 2610
box -4 -6 20 206
use NOR2X1  NOR2X1_134
timestamp 1742918108
transform 1 0 4904 0 1 2610
box -4 -6 52 206
use NOR2X1  NOR2X1_90
timestamp 1742918108
transform -1 0 5000 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_58
timestamp 1742918108
transform -1 0 5032 0 1 2610
box -4 -6 36 206
use NOR2X1  NOR2X1_38
timestamp 1742918108
transform -1 0 5080 0 1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_62
timestamp 1742918108
transform 1 0 5080 0 1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_113
timestamp 1742918108
transform 1 0 5272 0 1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_112
timestamp 1742918108
transform 1 0 5464 0 1 2610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_131
timestamp 1742918108
transform 1 0 5656 0 1 2610
box -4 -6 196 206
use BUFX2  BUFX2_6
timestamp 1742918108
transform 1 0 5848 0 1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_111
timestamp 1742918108
transform 1 0 5896 0 1 2610
box -4 -6 196 206
use BUFX2  BUFX2_4
timestamp 1742918108
transform 1 0 6088 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_9
timestamp 1742918108
transform 1 0 6136 0 1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_114
timestamp 1742918108
transform 1 0 6184 0 1 2610
box -4 -6 196 206
use BUFX2  BUFX2_7
timestamp 1742918108
transform 1 0 6376 0 1 2610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_135
timestamp 1742918108
transform 1 0 6424 0 1 2610
box -4 -6 196 206
use FILL  FILL_14_1
timestamp 1742918108
transform 1 0 6616 0 1 2610
box -4 -6 20 206
use FILL  FILL_14_2
timestamp 1742918108
transform 1 0 6632 0 1 2610
box -4 -6 20 206
use NAND3X1  NAND3X1_97
timestamp 1742918108
transform -1 0 72 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_98
timestamp 1742918108
transform -1 0 136 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_92
timestamp 1742918108
transform -1 0 200 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_224
timestamp 1742918108
transform 1 0 200 0 -1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_96
timestamp 1742918108
transform 1 0 248 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_95
timestamp 1742918108
transform 1 0 312 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_76
timestamp 1742918108
transform -1 0 440 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_240
timestamp 1742918108
transform -1 0 504 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_198
timestamp 1742918108
transform -1 0 536 0 -1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_277
timestamp 1742918108
transform -1 0 584 0 -1 3010
box -4 -6 52 206
use AOI21X1  AOI21X1_73
timestamp 1742918108
transform 1 0 584 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_85
timestamp 1742918108
transform -1 0 712 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_80
timestamp 1742918108
transform -1 0 776 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_70
timestamp 1742918108
transform -1 0 840 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_197
timestamp 1742918108
transform -1 0 888 0 -1 3010
box -4 -6 52 206
use INVX1  INVX1_190
timestamp 1742918108
transform -1 0 920 0 -1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_79
timestamp 1742918108
transform 1 0 920 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_196
timestamp 1742918108
transform 1 0 984 0 -1 3010
box -4 -6 52 206
use OR2X2  OR2X2_15
timestamp 1742918108
transform -1 0 1096 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_223
timestamp 1742918108
transform 1 0 1096 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_78
timestamp 1742918108
transform -1 0 1224 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_193
timestamp 1742918108
transform -1 0 1272 0 -1 3010
box -4 -6 52 206
use INVX1  INVX1_186
timestamp 1742918108
transform -1 0 1304 0 -1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_76
timestamp 1742918108
transform -1 0 1368 0 -1 3010
box -4 -6 68 206
use CLKBUF1  CLKBUF1_10
timestamp 1742918108
transform -1 0 1512 0 -1 3010
box -4 -6 148 206
use NAND2X1  NAND2X1_80
timestamp 1742918108
transform -1 0 1560 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_111
timestamp 1742918108
transform 1 0 1560 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_115
timestamp 1742918108
transform 1 0 1624 0 -1 3010
box -4 -6 196 206
use FILL  FILL_14_0_0
timestamp 1742918108
transform -1 0 1832 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_0_1
timestamp 1742918108
transform -1 0 1848 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_0_2
timestamp 1742918108
transform -1 0 1864 0 -1 3010
box -4 -6 20 206
use NOR2X1  NOR2X1_71
timestamp 1742918108
transform -1 0 1912 0 -1 3010
box -4 -6 52 206
use AOI21X1  AOI21X1_19
timestamp 1742918108
transform 1 0 1912 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_115
timestamp 1742918108
transform 1 0 1976 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_118
timestamp 1742918108
transform -1 0 2072 0 -1 3010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_17
timestamp 1742918108
transform -1 0 2264 0 -1 3010
box -4 -6 196 206
use OAI21X1  OAI21X1_135
timestamp 1742918108
transform -1 0 2328 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_49
timestamp 1742918108
transform -1 0 2392 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_63
timestamp 1742918108
transform -1 0 2424 0 -1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_54
timestamp 1742918108
transform -1 0 2472 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_101
timestamp 1742918108
transform 1 0 2472 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_23
timestamp 1742918108
transform -1 0 2712 0 -1 3010
box -4 -6 196 206
use OAI21X1  OAI21X1_141
timestamp 1742918108
transform -1 0 2776 0 -1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_68
timestamp 1742918108
transform 1 0 2776 0 -1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_67
timestamp 1742918108
transform 1 0 2824 0 -1 3010
box -4 -6 52 206
use INVX1  INVX1_82
timestamp 1742918108
transform -1 0 2904 0 -1 3010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_73
timestamp 1742918108
transform -1 0 3096 0 -1 3010
box -4 -6 196 206
use INVX1  INVX1_67
timestamp 1742918108
transform 1 0 3096 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_52
timestamp 1742918108
transform 1 0 3128 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_84
timestamp 1742918108
transform 1 0 3192 0 -1 3010
box -4 -6 196 206
use FILL  FILL_14_1_0
timestamp 1742918108
transform 1 0 3384 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_1_1
timestamp 1742918108
transform 1 0 3400 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_1_2
timestamp 1742918108
transform 1 0 3416 0 -1 3010
box -4 -6 20 206
use BUFX2  BUFX2_11
timestamp 1742918108
transform 1 0 3432 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_98
timestamp 1742918108
transform -1 0 3544 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_100
timestamp 1742918108
transform -1 0 3576 0 -1 3010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_40
timestamp 1742918108
transform 1 0 3576 0 -1 3010
box -4 -6 196 206
use OAI21X1  OAI21X1_91
timestamp 1742918108
transform -1 0 3832 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_33
timestamp 1742918108
transform 1 0 3832 0 -1 3010
box -4 -6 196 206
use NAND2X1  NAND2X1_426
timestamp 1742918108
transform -1 0 4072 0 -1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_54
timestamp 1742918108
transform 1 0 4072 0 -1 3010
box -4 -6 52 206
use INVX1  INVX1_88
timestamp 1742918108
transform -1 0 4152 0 -1 3010
box -4 -6 36 206
use XNOR2X1  XNOR2X1_51
timestamp 1742918108
transform -1 0 4264 0 -1 3010
box -4 -6 116 206
use XOR2X1  XOR2X1_23
timestamp 1742918108
transform -1 0 4376 0 -1 3010
box -4 -6 116 206
use NAND3X1  NAND3X1_347
timestamp 1742918108
transform -1 0 4440 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_155
timestamp 1742918108
transform 1 0 4440 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_381
timestamp 1742918108
transform 1 0 4504 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_383
timestamp 1742918108
transform 1 0 4568 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_307
timestamp 1742918108
transform -1 0 4664 0 -1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_349
timestamp 1742918108
transform 1 0 4664 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_348
timestamp 1742918108
transform 1 0 4728 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_351
timestamp 1742918108
transform 1 0 4792 0 -1 3010
box -4 -6 68 206
use FILL  FILL_14_2_0
timestamp 1742918108
transform 1 0 4856 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_2_1
timestamp 1742918108
transform 1 0 4872 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_2_2
timestamp 1742918108
transform 1 0 4888 0 -1 3010
box -4 -6 20 206
use NAND3X1  NAND3X1_352
timestamp 1742918108
transform 1 0 4904 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_427
timestamp 1742918108
transform 1 0 4968 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_429
timestamp 1742918108
transform 1 0 5016 0 -1 3010
box -4 -6 52 206
use XOR2X1  XOR2X1_24
timestamp 1742918108
transform 1 0 5064 0 -1 3010
box -4 -6 116 206
use NAND3X1  NAND3X1_354
timestamp 1742918108
transform -1 0 5240 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_158
timestamp 1742918108
transform -1 0 5304 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_436
timestamp 1742918108
transform -1 0 5352 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_430
timestamp 1742918108
transform 1 0 5352 0 -1 3010
box -4 -6 52 206
use OR2X2  OR2X2_33
timestamp 1742918108
transform 1 0 5400 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_159
timestamp 1742918108
transform 1 0 5464 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_353
timestamp 1742918108
transform 1 0 5528 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_385
timestamp 1742918108
transform 1 0 5592 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_308
timestamp 1742918108
transform 1 0 5656 0 -1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_355
timestamp 1742918108
transform 1 0 5688 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_437
timestamp 1742918108
transform -1 0 5800 0 -1 3010
box -4 -6 52 206
use AOI21X1  AOI21X1_161
timestamp 1742918108
transform 1 0 5800 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_356
timestamp 1742918108
transform 1 0 5864 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_310
timestamp 1742918108
transform 1 0 5928 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_388
timestamp 1742918108
transform 1 0 5960 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_164
timestamp 1742918108
transform -1 0 6088 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_364
timestamp 1742918108
transform 1 0 6088 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_444
timestamp 1742918108
transform -1 0 6200 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_120
timestamp 1742918108
transform 1 0 6200 0 -1 3010
box -4 -6 196 206
use BUFX2  BUFX2_10
timestamp 1742918108
transform 1 0 6392 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_16
timestamp 1742918108
transform 1 0 6440 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_28
timestamp 1742918108
transform 1 0 6488 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_8
timestamp 1742918108
transform 1 0 6536 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_30
timestamp 1742918108
transform 1 0 6584 0 -1 3010
box -4 -6 52 206
use FILL  FILL_15_1
timestamp 1742918108
transform -1 0 6648 0 -1 3010
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_119
timestamp 1742918108
transform 1 0 8 0 1 3010
box -4 -6 196 206
use XOR2X1  XOR2X1_13
timestamp 1742918108
transform 1 0 200 0 1 3010
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_118
timestamp 1742918108
transform 1 0 312 0 1 3010
box -4 -6 196 206
use NOR2X1  NOR2X1_161
timestamp 1742918108
transform -1 0 552 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_162
timestamp 1742918108
transform -1 0 600 0 1 3010
box -4 -6 52 206
use INVX1  INVX1_191
timestamp 1742918108
transform -1 0 632 0 1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_11
timestamp 1742918108
transform 1 0 632 0 1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_141
timestamp 1742918108
transform -1 0 744 0 1 3010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_116
timestamp 1742918108
transform 1 0 744 0 1 3010
box -4 -6 196 206
use NAND2X1  NAND2X1_195
timestamp 1742918108
transform 1 0 936 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_222
timestamp 1742918108
transform -1 0 1048 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_194
timestamp 1742918108
transform -1 0 1096 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_138
timestamp 1742918108
transform -1 0 1144 0 1 3010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_12
timestamp 1742918108
transform 1 0 1144 0 1 3010
box -4 -6 116 206
use INVX1  INVX1_114
timestamp 1742918108
transform 1 0 1256 0 1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_81
timestamp 1742918108
transform 1 0 1288 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_110
timestamp 1742918108
transform 1 0 1336 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_113
timestamp 1742918108
transform 1 0 1400 0 1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_82
timestamp 1742918108
transform -1 0 1480 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_112
timestamp 1742918108
transform 1 0 1480 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_72
timestamp 1742918108
transform 1 0 1544 0 1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_8
timestamp 1742918108
transform 1 0 1592 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_114
timestamp 1742918108
transform 1 0 1656 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_18
timestamp 1742918108
transform 1 0 1720 0 1 3010
box -4 -6 68 206
use FILL  FILL_15_0_0
timestamp 1742918108
transform 1 0 1784 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_0_1
timestamp 1742918108
transform 1 0 1800 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_0_2
timestamp 1742918108
transform 1 0 1816 0 1 3010
box -4 -6 20 206
use CLKBUF1  CLKBUF1_8
timestamp 1742918108
transform 1 0 1832 0 1 3010
box -4 -6 148 206
use BUFX4  BUFX4_12
timestamp 1742918108
transform 1 0 1976 0 1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_81
timestamp 1742918108
transform 1 0 2040 0 1 3010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_57
timestamp 1742918108
transform 1 0 2232 0 1 3010
box -4 -6 196 206
use NAND2X1  NAND2X1_56
timestamp 1742918108
transform -1 0 2472 0 1 3010
box -4 -6 52 206
use INVX1  INVX1_52
timestamp 1742918108
transform 1 0 2472 0 1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_60
timestamp 1742918108
transform 1 0 2504 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_97
timestamp 1742918108
transform -1 0 2616 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_99
timestamp 1742918108
transform -1 0 2648 0 1 3010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_39
timestamp 1742918108
transform 1 0 2648 0 1 3010
box -4 -6 196 206
use AOI21X1  AOI21X1_12
timestamp 1742918108
transform 1 0 2840 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_85
timestamp 1742918108
transform 1 0 2904 0 1 3010
box -4 -6 52 206
use BUFX4  BUFX4_7
timestamp 1742918108
transform 1 0 2952 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_57
timestamp 1742918108
transform 1 0 3016 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_94
timestamp 1742918108
transform -1 0 3128 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_96
timestamp 1742918108
transform -1 0 3192 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_98
timestamp 1742918108
transform -1 0 3224 0 1 3010
box -4 -6 36 206
use FILL  FILL_15_1_0
timestamp 1742918108
transform 1 0 3224 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_1_1
timestamp 1742918108
transform 1 0 3240 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_1_2
timestamp 1742918108
transform 1 0 3256 0 1 3010
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_38
timestamp 1742918108
transform 1 0 3272 0 1 3010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_79
timestamp 1742918108
transform 1 0 3464 0 1 3010
box -4 -6 196 206
use NAND2X1  NAND2X1_425
timestamp 1742918108
transform 1 0 3656 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_419
timestamp 1742918108
transform 1 0 3704 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_420
timestamp 1742918108
transform 1 0 3752 0 1 3010
box -4 -6 52 206
use INVX1  INVX1_93
timestamp 1742918108
transform -1 0 3832 0 1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_433
timestamp 1742918108
transform 1 0 3832 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_225
timestamp 1742918108
transform 1 0 3880 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_434
timestamp 1742918108
transform 1 0 3928 0 1 3010
box -4 -6 52 206
use AOI22X1  AOI22X1_52
timestamp 1742918108
transform 1 0 3976 0 1 3010
box -4 -6 84 206
use NAND3X1  NAND3X1_299
timestamp 1742918108
transform -1 0 4120 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_376
timestamp 1742918108
transform 1 0 4120 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_428
timestamp 1742918108
transform 1 0 4184 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_224
timestamp 1742918108
transform 1 0 4232 0 1 3010
box -4 -6 52 206
use AOI21X1  AOI21X1_153
timestamp 1742918108
transform -1 0 4344 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_303
timestamp 1742918108
transform -1 0 4408 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_156
timestamp 1742918108
transform 1 0 4408 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_157
timestamp 1742918108
transform -1 0 4536 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_305
timestamp 1742918108
transform -1 0 4600 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_310
timestamp 1742918108
transform -1 0 4664 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_312
timestamp 1742918108
transform -1 0 4728 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_315
timestamp 1742918108
transform -1 0 4792 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_308
timestamp 1742918108
transform 1 0 4792 0 1 3010
box -4 -6 68 206
use FILL  FILL_15_2_0
timestamp 1742918108
transform 1 0 4856 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_2_1
timestamp 1742918108
transform 1 0 4872 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_2_2
timestamp 1742918108
transform 1 0 4888 0 1 3010
box -4 -6 20 206
use NAND3X1  NAND3X1_314
timestamp 1742918108
transform 1 0 4904 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_375
timestamp 1742918108
transform 1 0 4968 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_319
timestamp 1742918108
transform 1 0 5032 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_316
timestamp 1742918108
transform -1 0 5160 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_150
timestamp 1742918108
transform 1 0 5160 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_151
timestamp 1742918108
transform 1 0 5224 0 1 3010
box -4 -6 68 206
use XOR2X1  XOR2X1_22
timestamp 1742918108
transform -1 0 5400 0 1 3010
box -4 -6 116 206
use BUFX2  BUFX2_12
timestamp 1742918108
transform 1 0 5400 0 1 3010
box -4 -6 52 206
use INVX1  INVX1_309
timestamp 1742918108
transform 1 0 5448 0 1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_438
timestamp 1742918108
transform 1 0 5480 0 1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_359
timestamp 1742918108
transform -1 0 5592 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_357
timestamp 1742918108
transform 1 0 5592 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_363
timestamp 1742918108
transform -1 0 5720 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_165
timestamp 1742918108
transform 1 0 5720 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_389
timestamp 1742918108
transform -1 0 5848 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_358
timestamp 1742918108
transform 1 0 5848 0 1 3010
box -4 -6 68 206
use OAI22X1  OAI22X1_22
timestamp 1742918108
transform 1 0 5912 0 1 3010
box -4 -6 84 206
use NAND3X1  NAND3X1_365
timestamp 1742918108
transform -1 0 6056 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_361
timestamp 1742918108
transform 1 0 6056 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_362
timestamp 1742918108
transform -1 0 6184 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_445
timestamp 1742918108
transform 1 0 6184 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_14
timestamp 1742918108
transform 1 0 6232 0 1 3010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_132
timestamp 1742918108
transform 1 0 6280 0 1 3010
box -4 -6 196 206
use BUFX2  BUFX2_5
timestamp 1742918108
transform 1 0 6472 0 1 3010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_50
timestamp 1742918108
transform -1 0 6632 0 1 3010
box -4 -6 116 206
use FILL  FILL_16_1
timestamp 1742918108
transform 1 0 6632 0 1 3010
box -4 -6 20 206
use CLKBUF1  CLKBUF1_2
timestamp 1742918108
transform 1 0 8 0 -1 3410
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_68
timestamp 1742918108
transform 1 0 152 0 -1 3410
box -4 -6 196 206
use INVX1  INVX1_111
timestamp 1742918108
transform 1 0 344 0 -1 3410
box -4 -6 36 206
use NOR2X1  NOR2X1_65
timestamp 1742918108
transform 1 0 376 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_108
timestamp 1742918108
transform -1 0 488 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_66
timestamp 1742918108
transform -1 0 536 0 -1 3410
box -4 -6 52 206
use INVX1  INVX1_109
timestamp 1742918108
transform -1 0 568 0 -1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_109
timestamp 1742918108
transform -1 0 632 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_68
timestamp 1742918108
transform 1 0 632 0 -1 3410
box -4 -6 52 206
use BUFX4  BUFX4_16
timestamp 1742918108
transform -1 0 744 0 -1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_17
timestamp 1742918108
transform -1 0 808 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_10
timestamp 1742918108
transform -1 0 872 0 -1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_95
timestamp 1742918108
transform -1 0 920 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_37
timestamp 1742918108
transform -1 0 968 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_37
timestamp 1742918108
transform 1 0 968 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_23
timestamp 1742918108
transform -1 0 1080 0 -1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_54
timestamp 1742918108
transform 1 0 1080 0 -1 3410
box -4 -6 196 206
use NAND2X1  NAND2X1_106
timestamp 1742918108
transform 1 0 1272 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_145
timestamp 1742918108
transform -1 0 1384 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_147
timestamp 1742918108
transform 1 0 1384 0 -1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_31
timestamp 1742918108
transform 1 0 1448 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_12
timestamp 1742918108
transform -1 0 1576 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_115
timestamp 1742918108
transform -1 0 1608 0 -1 3410
box -4 -6 36 206
use NOR2X1  NOR2X1_66
timestamp 1742918108
transform -1 0 1656 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_79
timestamp 1742918108
transform -1 0 1704 0 -1 3410
box -4 -6 52 206
use AND2X2  AND2X2_12
timestamp 1742918108
transform 1 0 1704 0 -1 3410
box -4 -6 68 206
use FILL  FILL_16_0_0
timestamp 1742918108
transform -1 0 1784 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_0_1
timestamp 1742918108
transform -1 0 1800 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_0_2
timestamp 1742918108
transform -1 0 1816 0 -1 3410
box -4 -6 20 206
use OAI21X1  OAI21X1_146
timestamp 1742918108
transform -1 0 1880 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_83
timestamp 1742918108
transform -1 0 1928 0 -1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_18
timestamp 1742918108
transform -1 0 2120 0 -1 3410
box -4 -6 196 206
use NAND2X1  NAND2X1_96
timestamp 1742918108
transform 1 0 2120 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_136
timestamp 1742918108
transform -1 0 2232 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_83
timestamp 1742918108
transform 1 0 2232 0 -1 3410
box -4 -6 196 206
use INVX1  INVX1_66
timestamp 1742918108
transform 1 0 2424 0 -1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_51
timestamp 1742918108
transform 1 0 2456 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_98
timestamp 1742918108
transform 1 0 2520 0 -1 3410
box -4 -6 52 206
use INVX1  INVX1_70
timestamp 1742918108
transform 1 0 2568 0 -1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_55
timestamp 1742918108
transform 1 0 2600 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_87
timestamp 1742918108
transform -1 0 2856 0 -1 3410
box -4 -6 196 206
use OAI21X1  OAI21X1_93
timestamp 1742918108
transform -1 0 2920 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_95
timestamp 1742918108
transform -1 0 2952 0 -1 3410
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_35
timestamp 1742918108
transform -1 0 3144 0 -1 3410
box -4 -6 196 206
use INVX1  INVX1_96
timestamp 1742918108
transform -1 0 3176 0 -1 3410
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_36
timestamp 1742918108
transform 1 0 3176 0 -1 3410
box -4 -6 196 206
use FILL  FILL_16_1_0
timestamp 1742918108
transform 1 0 3368 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_1_1
timestamp 1742918108
transform 1 0 3384 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_1_2
timestamp 1742918108
transform 1 0 3400 0 -1 3410
box -4 -6 20 206
use CLKBUF1  CLKBUF1_4
timestamp 1742918108
transform 1 0 3416 0 -1 3410
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_117
timestamp 1742918108
transform 1 0 3560 0 -1 3410
box -4 -6 196 206
use NAND3X1  NAND3X1_307
timestamp 1742918108
transform -1 0 3816 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_311
timestamp 1742918108
transform -1 0 3880 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_300
timestamp 1742918108
transform -1 0 3912 0 -1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_367
timestamp 1742918108
transform -1 0 3976 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_368
timestamp 1742918108
transform 1 0 3976 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_379
timestamp 1742918108
transform -1 0 4104 0 -1 3410
box -4 -6 68 206
use BUFX2  BUFX2_13
timestamp 1742918108
transform 1 0 4104 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_416
timestamp 1742918108
transform -1 0 4200 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_418
timestamp 1742918108
transform 1 0 4200 0 -1 3410
box -4 -6 52 206
use NAND3X1  NAND3X1_300
timestamp 1742918108
transform -1 0 4312 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_366
timestamp 1742918108
transform -1 0 4376 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_298
timestamp 1742918108
transform -1 0 4440 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_304
timestamp 1742918108
transform 1 0 4440 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_301
timestamp 1742918108
transform -1 0 4568 0 -1 3410
box -4 -6 68 206
use INVX2  INVX2_44
timestamp 1742918108
transform 1 0 4568 0 -1 3410
box -4 -6 36 206
use NAND3X1  NAND3X1_309
timestamp 1742918108
transform -1 0 4664 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_302
timestamp 1742918108
transform 1 0 4664 0 -1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_152
timestamp 1742918108
transform 1 0 4728 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_313
timestamp 1742918108
transform -1 0 4856 0 -1 3410
box -4 -6 68 206
use FILL  FILL_16_2_0
timestamp 1742918108
transform -1 0 4872 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_2_1
timestamp 1742918108
transform -1 0 4888 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_2_2
timestamp 1742918108
transform -1 0 4904 0 -1 3410
box -4 -6 20 206
use NAND3X1  NAND3X1_318
timestamp 1742918108
transform -1 0 4968 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_323
timestamp 1742918108
transform -1 0 5032 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_320
timestamp 1742918108
transform -1 0 5096 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_302
timestamp 1742918108
transform 1 0 5096 0 -1 3410
box -4 -6 36 206
use NAND3X1  NAND3X1_322
timestamp 1742918108
transform 1 0 5128 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_317
timestamp 1742918108
transform -1 0 5256 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_321
timestamp 1742918108
transform -1 0 5320 0 -1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_145
timestamp 1742918108
transform 1 0 5320 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_327
timestamp 1742918108
transform -1 0 5448 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_387
timestamp 1742918108
transform 1 0 5448 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_440
timestamp 1742918108
transform -1 0 5560 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_441
timestamp 1742918108
transform -1 0 5608 0 -1 3410
box -4 -6 52 206
use AOI21X1  AOI21X1_144
timestamp 1742918108
transform -1 0 5672 0 -1 3410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_52
timestamp 1742918108
transform -1 0 5784 0 -1 3410
box -4 -6 116 206
use NAND2X1  NAND2X1_439
timestamp 1742918108
transform -1 0 5832 0 -1 3410
box -4 -6 52 206
use INVX1  INVX1_311
timestamp 1742918108
transform 1 0 5832 0 -1 3410
box -4 -6 36 206
use NAND3X1  NAND3X1_360
timestamp 1742918108
transform -1 0 5928 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_442
timestamp 1742918108
transform 1 0 5928 0 -1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_226
timestamp 1742918108
transform -1 0 6024 0 -1 3410
box -4 -6 52 206
use OR2X2  OR2X2_34
timestamp 1742918108
transform 1 0 6024 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_294
timestamp 1742918108
transform -1 0 6120 0 -1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_392
timestamp 1742918108
transform -1 0 6184 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_366
timestamp 1742918108
transform -1 0 6248 0 -1 3410
box -4 -6 68 206
use DFFSR  DFFSR_1
timestamp 1742918108
transform -1 0 6600 0 -1 3410
box -4 -6 356 206
use FILL  FILL_17_1
timestamp 1742918108
transform -1 0 6616 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_2
timestamp 1742918108
transform -1 0 6632 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_3
timestamp 1742918108
transform -1 0 6648 0 -1 3410
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_91
timestamp 1742918108
transform 1 0 8 0 1 3410
box -4 -6 196 206
use INVX1  INVX1_89
timestamp 1742918108
transform -1 0 232 0 1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_5
timestamp 1742918108
transform 1 0 232 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_6
timestamp 1742918108
transform -1 0 344 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_34
timestamp 1742918108
transform -1 0 392 0 1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_89
timestamp 1742918108
transform -1 0 200 0 -1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_7
timestamp 1742918108
transform 1 0 200 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_9
timestamp 1742918108
transform -1 0 312 0 -1 3810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_92
timestamp 1742918108
transform -1 0 504 0 -1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_61
timestamp 1742918108
transform -1 0 456 0 1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_67
timestamp 1742918108
transform 1 0 456 0 1 3410
box -4 -6 196 206
use NAND2X1  NAND2X1_67
timestamp 1742918108
transform -1 0 696 0 1 3410
box -4 -6 52 206
use BUFX4  BUFX4_15
timestamp 1742918108
transform -1 0 760 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_62
timestamp 1742918108
transform 1 0 504 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_35
timestamp 1742918108
transform -1 0 616 0 -1 3810
box -4 -6 52 206
use INVX1  INVX1_112
timestamp 1742918108
transform 1 0 616 0 -1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_17
timestamp 1742918108
transform 1 0 648 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_31
timestamp 1742918108
transform -1 0 760 0 -1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_16
timestamp 1742918108
transform -1 0 952 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_63
timestamp 1742918108
transform 1 0 840 0 1 3410
box -4 -6 52 206
use INVX1  INVX1_110
timestamp 1742918108
transform 1 0 808 0 1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_64
timestamp 1742918108
transform 1 0 760 0 1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_103
timestamp 1742918108
transform 1 0 1048 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_104
timestamp 1742918108
transform 1 0 1000 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_22
timestamp 1742918108
transform -1 0 1000 0 -1 3810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_13
timestamp 1742918108
transform -1 0 1176 0 1 3410
box -4 -6 116 206
use OAI21X1  OAI21X1_144
timestamp 1742918108
transform 1 0 1000 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_65
timestamp 1742918108
transform -1 0 1000 0 1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_51
timestamp 1742918108
transform -1 0 952 0 -1 3810
box -4 -6 196 206
use AOI21X1  AOI21X1_29
timestamp 1742918108
transform 1 0 1176 0 1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_70
timestamp 1742918108
transform -1 0 1432 0 1 3410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_53
timestamp 1742918108
transform 1 0 1432 0 1 3410
box -4 -6 196 206
use OAI21X1  OAI21X1_143
timestamp 1742918108
transform -1 0 1160 0 -1 3810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_11
timestamp 1742918108
transform -1 0 1272 0 -1 3810
box -4 -6 116 206
use OAI21X1  OAI21X1_65
timestamp 1742918108
transform -1 0 1336 0 -1 3810
box -4 -6 68 206
use AND2X2  AND2X2_3
timestamp 1742918108
transform 1 0 1336 0 -1 3810
box -4 -6 68 206
use OAI22X1  OAI22X1_3
timestamp 1742918108
transform -1 0 1480 0 -1 3810
box -4 -6 84 206
use NAND2X1  NAND2X1_105
timestamp 1742918108
transform -1 0 1672 0 1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_69
timestamp 1742918108
transform -1 0 1720 0 1 3410
box -4 -6 52 206
use INVX1  INVX1_75
timestamp 1742918108
transform -1 0 1704 0 -1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_71
timestamp 1742918108
transform 1 0 1720 0 1 3410
box -4 -6 52 206
use INVX1  INVX1_41
timestamp 1742918108
transform 1 0 1704 0 -1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_70
timestamp 1742918108
transform 1 0 1736 0 -1 3810
box -4 -6 52 206
use FILL  FILL_17_0_0
timestamp 1742918108
transform 1 0 1768 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_0_1
timestamp 1742918108
transform 1 0 1784 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_0_0
timestamp 1742918108
transform -1 0 1800 0 -1 3810
box -4 -6 20 206
use FILL  FILL_17_0_2
timestamp 1742918108
transform 1 0 1800 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_0_1
timestamp 1742918108
transform -1 0 1816 0 -1 3810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_69
timestamp 1742918108
transform 1 0 1480 0 -1 3810
box -4 -6 196 206
use FILL  FILL_18_0_2
timestamp 1742918108
transform -1 0 1832 0 -1 3810
box -4 -6 20 206
use XOR2X1  XOR2X1_4
timestamp 1742918108
transform 1 0 1880 0 1 3410
box -4 -6 116 206
use AOI21X1  AOI21X1_30
timestamp 1742918108
transform 1 0 1816 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_78
timestamp 1742918108
transform -1 0 2200 0 -1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_9
timestamp 1742918108
transform 1 0 2104 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_47
timestamp 1742918108
transform 1 0 2072 0 -1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_73
timestamp 1742918108
transform -1 0 2072 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_77
timestamp 1742918108
transform -1 0 2200 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_113
timestamp 1742918108
transform -1 0 2152 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_74
timestamp 1742918108
transform -1 0 2088 0 1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_75
timestamp 1742918108
transform 1 0 1992 0 1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_55
timestamp 1742918108
transform -1 0 2024 0 -1 3810
box -4 -6 196 206
use INVX1  INVX1_116
timestamp 1742918108
transform -1 0 2232 0 1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_108
timestamp 1742918108
transform -1 0 2280 0 1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_76
timestamp 1742918108
transform 1 0 2280 0 1 3410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_20
timestamp 1742918108
transform -1 0 2520 0 1 3410
box -4 -6 196 206
use OAI21X1  OAI21X1_138
timestamp 1742918108
transform -1 0 2584 0 1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_56
timestamp 1742918108
transform -1 0 2392 0 -1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_40
timestamp 1742918108
transform 1 0 2392 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_30
timestamp 1742918108
transform 1 0 2456 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_15
timestamp 1742918108
transform 1 0 2504 0 -1 3810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_21
timestamp 1742918108
transform -1 0 2776 0 1 3410
box -4 -6 196 206
use NAND2X1  NAND2X1_59
timestamp 1742918108
transform 1 0 2776 0 1 3410
box -4 -6 52 206
use BUFX4  BUFX4_1
timestamp 1742918108
transform 1 0 2824 0 1 3410
box -4 -6 68 206
use BUFX4  BUFX4_6
timestamp 1742918108
transform 1 0 2888 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_99
timestamp 1742918108
transform 1 0 2552 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_139
timestamp 1742918108
transform -1 0 2664 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_86
timestamp 1742918108
transform 1 0 2664 0 -1 3810
box -4 -6 196 206
use INVX1  INVX1_69
timestamp 1742918108
transform 1 0 2856 0 -1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_54
timestamp 1742918108
transform -1 0 2952 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_58
timestamp 1742918108
transform -1 0 3000 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_19
timestamp 1742918108
transform 1 0 3000 0 1 3410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_99
timestamp 1742918108
transform 1 0 3064 0 1 3410
box -4 -6 196 206
use BUFX4  BUFX4_14
timestamp 1742918108
transform 1 0 2952 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_20
timestamp 1742918108
transform 1 0 3016 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_100
timestamp 1742918108
transform 1 0 3080 0 -1 3810
box -4 -6 196 206
use INVX2  INVX2_3
timestamp 1742918108
transform 1 0 3256 0 1 3410
box -4 -6 36 206
use FILL  FILL_17_1_0
timestamp 1742918108
transform -1 0 3304 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_1_1
timestamp 1742918108
transform -1 0 3320 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_1_2
timestamp 1742918108
transform -1 0 3336 0 1 3410
box -4 -6 20 206
use INVX1  INVX1_27
timestamp 1742918108
transform 1 0 3272 0 -1 3810
box -4 -6 36 206
use FILL  FILL_18_1_0
timestamp 1742918108
transform -1 0 3320 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_1_1
timestamp 1742918108
transform -1 0 3336 0 -1 3810
box -4 -6 20 206
use OAI21X1  OAI21X1_24
timestamp 1742918108
transform -1 0 3400 0 1 3410
box -4 -6 68 206
use FILL  FILL_18_1_2
timestamp 1742918108
transform -1 0 3352 0 -1 3810
box -4 -6 20 206
use NOR2X1  NOR2X1_61
timestamp 1742918108
transform -1 0 3400 0 -1 3810
box -4 -6 52 206
use INVX1  INVX1_30
timestamp 1742918108
transform -1 0 3432 0 1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_53
timestamp 1742918108
transform -1 0 3480 0 1 3410
box -4 -6 52 206
use AOI21X1  AOI21X1_14
timestamp 1742918108
transform -1 0 3464 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_89
timestamp 1742918108
transform -1 0 3640 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_88
timestamp 1742918108
transform -1 0 3576 0 -1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_59
timestamp 1742918108
transform 1 0 3464 0 -1 3810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_104
timestamp 1742918108
transform 1 0 3480 0 1 3410
box -4 -6 196 206
use OAI21X1  OAI21X1_95
timestamp 1742918108
transform -1 0 3736 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_97
timestamp 1742918108
transform -1 0 3768 0 1 3410
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_37
timestamp 1742918108
transform 1 0 3768 0 1 3410
box -4 -6 196 206
use INVX1  INVX1_301
timestamp 1742918108
transform 1 0 3960 0 1 3410
box -4 -6 36 206
use INVX1  INVX1_92
timestamp 1742918108
transform -1 0 3672 0 -1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_90
timestamp 1742918108
transform -1 0 3736 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_48
timestamp 1742918108
transform 1 0 3736 0 -1 3810
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_41
timestamp 1742918108
transform 1 0 3928 0 -1 3810
box -4 -6 196 206
use NAND3X1  NAND3X1_306
timestamp 1742918108
transform -1 0 4056 0 1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_143
timestamp 1742918108
transform -1 0 4120 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_421
timestamp 1742918108
transform -1 0 4232 0 -1 3810
box -4 -6 52 206
use NAND3X1  NAND3X1_346
timestamp 1742918108
transform 1 0 4120 0 -1 3810
box -4 -6 68 206
use AND2X2  AND2X2_46
timestamp 1742918108
transform -1 0 4248 0 1 3410
box -4 -6 68 206
use AND2X2  AND2X2_47
timestamp 1742918108
transform -1 0 4184 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_422
timestamp 1742918108
transform -1 0 4280 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_417
timestamp 1742918108
transform 1 0 4248 0 1 3410
box -4 -6 52 206
use AND2X2  AND2X2_48
timestamp 1742918108
transform 1 0 4328 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_412
timestamp 1742918108
transform 1 0 4280 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_369
timestamp 1742918108
transform 1 0 4328 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_299
timestamp 1742918108
transform 1 0 4296 0 1 3410
box -4 -6 36 206
use OAI22X1  OAI22X1_21
timestamp 1742918108
transform 1 0 4392 0 -1 3810
box -4 -6 84 206
use OAI21X1  OAI21X1_380
timestamp 1742918108
transform 1 0 4392 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_350
timestamp 1742918108
transform -1 0 4536 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_291
timestamp 1742918108
transform 1 0 4504 0 1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_415
timestamp 1742918108
transform -1 0 4504 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_365
timestamp 1742918108
transform 1 0 4536 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_378
timestamp 1742918108
transform 1 0 4536 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_290
timestamp 1742918108
transform 1 0 4664 0 -1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_345
timestamp 1742918108
transform -1 0 4664 0 -1 3810
box -4 -6 68 206
use AOI22X1  AOI22X1_51
timestamp 1742918108
transform 1 0 4648 0 1 3410
box -4 -6 84 206
use NAND2X1  NAND2X1_431
timestamp 1742918108
transform 1 0 4600 0 1 3410
box -4 -6 52 206
use FILL  FILL_18_2_0
timestamp 1742918108
transform 1 0 4808 0 -1 3810
box -4 -6 20 206
use NOR2X1  NOR2X1_218
timestamp 1742918108
transform 1 0 4760 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_336
timestamp 1742918108
transform 1 0 4696 0 -1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_217
timestamp 1742918108
transform -1 0 4840 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_382
timestamp 1742918108
transform 1 0 4728 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_207
timestamp 1742918108
transform 1 0 4920 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_349
timestamp 1742918108
transform 1 0 4856 0 -1 3810
box -4 -6 68 206
use FILL  FILL_18_2_2
timestamp 1742918108
transform 1 0 4840 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_2_1
timestamp 1742918108
transform 1 0 4824 0 -1 3810
box -4 -6 20 206
use NAND2X1  NAND2X1_435
timestamp 1742918108
transform 1 0 4888 0 1 3410
box -4 -6 52 206
use FILL  FILL_17_2_2
timestamp 1742918108
transform 1 0 4872 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_2_1
timestamp 1742918108
transform 1 0 4856 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_2_0
timestamp 1742918108
transform 1 0 4840 0 1 3410
box -4 -6 20 206
use NAND2X1  NAND2X1_364
timestamp 1742918108
transform -1 0 5096 0 -1 3810
box -4 -6 52 206
use AOI22X1  AOI22X1_42
timestamp 1742918108
transform 1 0 4968 0 -1 3810
box -4 -6 84 206
use INVX1  INVX1_298
timestamp 1742918108
transform -1 0 5080 0 1 3410
box -4 -6 36 206
use XNOR2X1  XNOR2X1_49
timestamp 1742918108
transform -1 0 5048 0 1 3410
box -4 -6 116 206
use INVX2  INVX2_38
timestamp 1742918108
transform 1 0 5144 0 -1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_411
timestamp 1742918108
transform 1 0 5096 0 -1 3810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_47
timestamp 1742918108
transform -1 0 5192 0 1 3410
box -4 -6 116 206
use XNOR2X1  XNOR2X1_46
timestamp 1742918108
transform -1 0 5400 0 -1 3810
box -4 -6 116 206
use NAND2X1  NAND2X1_362
timestamp 1742918108
transform 1 0 5240 0 -1 3810
box -4 -6 52 206
use NAND3X1  NAND3X1_267
timestamp 1742918108
transform -1 0 5240 0 -1 3810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_48
timestamp 1742918108
transform -1 0 5304 0 1 3410
box -4 -6 116 206
use NAND3X1  NAND3X1_331
timestamp 1742918108
transform -1 0 5464 0 -1 3810
box -4 -6 68 206
use INVX2  INVX2_35
timestamp 1742918108
transform 1 0 5384 0 1 3410
box -4 -6 36 206
use NOR2X1  NOR2X1_200
timestamp 1742918108
transform -1 0 5384 0 1 3410
box -4 -6 52 206
use INVX2  INVX2_36
timestamp 1742918108
transform -1 0 5336 0 1 3410
box -4 -6 36 206
use NAND3X1  NAND3X1_325
timestamp 1742918108
transform -1 0 5528 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_329
timestamp 1742918108
transform 1 0 5464 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_199
timestamp 1742918108
transform -1 0 5464 0 1 3410
box -4 -6 52 206
use AOI21X1  AOI21X1_149
timestamp 1742918108
transform 1 0 5528 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_328
timestamp 1742918108
transform 1 0 5560 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_303
timestamp 1742918108
transform 1 0 5528 0 1 3410
box -4 -6 36 206
use NAND3X1  NAND3X1_330
timestamp 1742918108
transform -1 0 5656 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_324
timestamp 1742918108
transform 1 0 5624 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_334
timestamp 1742918108
transform 1 0 5656 0 -1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_160
timestamp 1742918108
transform 1 0 5688 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_372
timestamp 1742918108
transform -1 0 5784 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_371
timestamp 1742918108
transform 1 0 5752 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_338
timestamp 1742918108
transform -1 0 5896 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_401
timestamp 1742918108
transform 1 0 5784 0 -1 3810
box -4 -6 52 206
use NAND3X1  NAND3X1_332
timestamp 1742918108
transform -1 0 5880 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_333
timestamp 1742918108
transform -1 0 5960 0 -1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_162
timestamp 1742918108
transform -1 0 5944 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_337
timestamp 1742918108
transform -1 0 6056 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_295
timestamp 1742918108
transform 1 0 5960 0 -1 3810
box -4 -6 36 206
use AOI21X1  AOI21X1_163
timestamp 1742918108
transform -1 0 6008 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_342
timestamp 1742918108
transform -1 0 6120 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_335
timestamp 1742918108
transform -1 0 6072 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_340
timestamp 1742918108
transform 1 0 6120 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_339
timestamp 1742918108
transform 1 0 6136 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_336
timestamp 1742918108
transform 1 0 6072 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_343
timestamp 1742918108
transform -1 0 6248 0 -1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_166
timestamp 1742918108
transform -1 0 6264 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_341
timestamp 1742918108
transform -1 0 6312 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_443
timestamp 1742918108
transform -1 0 6312 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_391
timestamp 1742918108
transform -1 0 6376 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_344
timestamp 1742918108
transform -1 0 6376 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_227
timestamp 1742918108
transform 1 0 6408 0 -1 3810
box -4 -6 52 206
use INVX1  INVX1_306
timestamp 1742918108
transform 1 0 6376 0 -1 3810
box -4 -6 36 206
use AOI21X1  AOI21X1_147
timestamp 1742918108
transform 1 0 6376 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_228
timestamp 1742918108
transform -1 0 6504 0 -1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_148
timestamp 1742918108
transform -1 0 6504 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_424
timestamp 1742918108
transform 1 0 6504 0 1 3410
box -4 -6 52 206
use NAND3X1  NAND3X1_54
timestamp 1742918108
transform 1 0 6552 0 1 3410
box -4 -6 68 206
use FILL  FILL_18_1
timestamp 1742918108
transform 1 0 6616 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_2
timestamp 1742918108
transform 1 0 6632 0 1 3410
box -4 -6 20 206
use XOR2X1  XOR2X1_21
timestamp 1742918108
transform -1 0 6616 0 -1 3810
box -4 -6 116 206
use FILL  FILL_19_1
timestamp 1742918108
transform -1 0 6632 0 -1 3810
box -4 -6 20 206
use FILL  FILL_19_2
timestamp 1742918108
transform -1 0 6648 0 -1 3810
box -4 -6 20 206
use NOR2X1  NOR2X1_55
timestamp 1742918108
transform -1 0 56 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_1
timestamp 1742918108
transform 1 0 56 0 1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_2
timestamp 1742918108
transform 1 0 88 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_39
timestamp 1742918108
transform -1 0 200 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_57
timestamp 1742918108
transform -1 0 264 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_56
timestamp 1742918108
transform -1 0 312 0 1 3810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_65
timestamp 1742918108
transform 1 0 312 0 1 3810
box -4 -6 196 206
use INVX1  INVX1_72
timestamp 1742918108
transform 1 0 504 0 1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_102
timestamp 1742918108
transform -1 0 584 0 1 3810
box -4 -6 52 206
use NOR2X1  NOR2X1_63
timestamp 1742918108
transform -1 0 632 0 1 3810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_49
timestamp 1742918108
transform -1 0 824 0 1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_33
timestamp 1742918108
transform 1 0 824 0 1 3810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_52
timestamp 1742918108
transform 1 0 888 0 1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_107
timestamp 1742918108
transform 1 0 1080 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_64
timestamp 1742918108
transform 1 0 1144 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_40
timestamp 1742918108
transform -1 0 1240 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_12
timestamp 1742918108
transform -1 0 1272 0 1 3810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_93
timestamp 1742918108
transform -1 0 1464 0 1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_35
timestamp 1742918108
transform -1 0 1528 0 1 3810
box -4 -6 68 206
use OAI22X1  OAI22X1_1
timestamp 1742918108
transform 1 0 1528 0 1 3810
box -4 -6 84 206
use OAI22X1  OAI22X1_5
timestamp 1742918108
transform 1 0 1608 0 1 3810
box -4 -6 84 206
use FILL  FILL_19_0_0
timestamp 1742918108
transform 1 0 1688 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_0_1
timestamp 1742918108
transform 1 0 1704 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_0_2
timestamp 1742918108
transform 1 0 1720 0 1 3810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_94
timestamp 1742918108
transform 1 0 1736 0 1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_11
timestamp 1742918108
transform 1 0 1928 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_10
timestamp 1742918108
transform -1 0 2040 0 1 3810
box -4 -6 52 206
use OR2X2  OR2X2_3
timestamp 1742918108
transform 1 0 2040 0 1 3810
box -4 -6 68 206
use INVX8  INVX8_1
timestamp 1742918108
transform 1 0 2104 0 1 3810
box -4 -6 84 206
use DFFPOSX1  DFFPOSX1_71
timestamp 1742918108
transform -1 0 2376 0 1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_70
timestamp 1742918108
transform 1 0 2376 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_80
timestamp 1742918108
transform -1 0 2472 0 1 3810
box -4 -6 36 206
use AOI22X1  AOI22X1_1
timestamp 1742918108
transform 1 0 2472 0 1 3810
box -4 -6 84 206
use DFFPOSX1  DFFPOSX1_72
timestamp 1742918108
transform -1 0 2744 0 1 3810
box -4 -6 196 206
use CLKBUF1  CLKBUF1_1
timestamp 1742918108
transform -1 0 2888 0 1 3810
box -4 -6 148 206
use BUFX4  BUFX4_8
timestamp 1742918108
transform -1 0 2952 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_68
timestamp 1742918108
transform 1 0 2952 0 1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_53
timestamp 1742918108
transform 1 0 2984 0 1 3810
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_85
timestamp 1742918108
transform -1 0 3240 0 1 3810
box -4 -6 196 206
use OAI21X1  OAI21X1_18
timestamp 1742918108
transform 1 0 3240 0 1 3810
box -4 -6 68 206
use FILL  FILL_19_1_0
timestamp 1742918108
transform 1 0 3304 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_1_1
timestamp 1742918108
transform 1 0 3320 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_1_2
timestamp 1742918108
transform 1 0 3336 0 1 3810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_98
timestamp 1742918108
transform 1 0 3352 0 1 3810
box -4 -6 196 206
use INVX2  INVX2_2
timestamp 1742918108
transform -1 0 3576 0 1 3810
box -4 -6 36 206
use AND2X2  AND2X2_10
timestamp 1742918108
transform -1 0 3640 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_44
timestamp 1742918108
transform 1 0 3640 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_78
timestamp 1742918108
transform 1 0 3688 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_79
timestamp 1742918108
transform 1 0 3752 0 1 3810
box -4 -6 68 206
use BUFX4  BUFX4_17
timestamp 1742918108
transform 1 0 3816 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_46
timestamp 1742918108
transform -1 0 3928 0 1 3810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_43
timestamp 1742918108
transform 1 0 3928 0 1 3810
box -4 -6 196 206
use XOR2X1  XOR2X1_5
timestamp 1742918108
transform -1 0 4232 0 1 3810
box -4 -6 116 206
use NAND2X1  NAND2X1_432
timestamp 1742918108
transform -1 0 4280 0 1 3810
box -4 -6 52 206
use AOI22X1  AOI22X1_50
timestamp 1742918108
transform 1 0 4280 0 1 3810
box -4 -6 84 206
use NAND2X1  NAND2X1_390
timestamp 1742918108
transform -1 0 4408 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_388
timestamp 1742918108
transform 1 0 4408 0 1 3810
box -4 -6 52 206
use XOR2X1  XOR2X1_25
timestamp 1742918108
transform -1 0 4568 0 1 3810
box -4 -6 116 206
use NAND2X1  NAND2X1_413
timestamp 1742918108
transform 1 0 4568 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_414
timestamp 1742918108
transform -1 0 4664 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_370
timestamp 1742918108
transform -1 0 4712 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_275
timestamp 1742918108
transform 1 0 4712 0 1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_340
timestamp 1742918108
transform 1 0 4744 0 1 3810
box -4 -6 68 206
use INVX2  INVX2_37
timestamp 1742918108
transform 1 0 4808 0 1 3810
box -4 -6 36 206
use FILL  FILL_19_2_0
timestamp 1742918108
transform 1 0 4840 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_2_1
timestamp 1742918108
transform 1 0 4856 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_2_2
timestamp 1742918108
transform 1 0 4872 0 1 3810
box -4 -6 20 206
use OAI21X1  OAI21X1_350
timestamp 1742918108
transform 1 0 4888 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_206
timestamp 1742918108
transform -1 0 5000 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_337
timestamp 1742918108
transform 1 0 5000 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_274
timestamp 1742918108
transform -1 0 5096 0 1 3810
box -4 -6 36 206
use NOR2X1  NOR2X1_202
timestamp 1742918108
transform -1 0 5144 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_365
timestamp 1742918108
transform 1 0 5144 0 1 3810
box -4 -6 52 206
use NAND3X1  NAND3X1_269
timestamp 1742918108
transform 1 0 5192 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_205
timestamp 1742918108
transform 1 0 5256 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_335
timestamp 1742918108
transform -1 0 5368 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_273
timestamp 1742918108
transform 1 0 5368 0 1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_333
timestamp 1742918108
transform 1 0 5400 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_338
timestamp 1742918108
transform 1 0 5464 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_334
timestamp 1742918108
transform 1 0 5528 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_366
timestamp 1742918108
transform -1 0 5640 0 1 3810
box -4 -6 52 206
use AND2X2  AND2X2_43
timestamp 1742918108
transform 1 0 5640 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_367
timestamp 1742918108
transform 1 0 5704 0 1 3810
box -4 -6 52 206
use OR2X2  OR2X2_28
timestamp 1742918108
transform 1 0 5752 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_368
timestamp 1742918108
transform 1 0 5816 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_369
timestamp 1742918108
transform -1 0 5912 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_276
timestamp 1742918108
transform -1 0 5944 0 1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_270
timestamp 1742918108
transform 1 0 5944 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_390
timestamp 1742918108
transform 1 0 6008 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_220
timestamp 1742918108
transform 1 0 6072 0 1 3810
box -4 -6 52 206
use NAND3X1  NAND3X1_271
timestamp 1742918108
transform -1 0 6184 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_272
timestamp 1742918108
transform 1 0 6184 0 1 3810
box -4 -6 36 206
use AOI21X1  AOI21X1_134
timestamp 1742918108
transform -1 0 6280 0 1 3810
box -4 -6 68 206
use AOI22X1  AOI22X1_54
timestamp 1742918108
transform -1 0 6360 0 1 3810
box -4 -6 84 206
use NOR2X1  NOR2X1_208
timestamp 1742918108
transform 1 0 6360 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_277
timestamp 1742918108
transform -1 0 6440 0 1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_446
timestamp 1742918108
transform -1 0 6488 0 1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_137
timestamp 1742918108
transform -1 0 6552 0 1 3810
box -4 -6 68 206
use AOI22X1  AOI22X1_53
timestamp 1742918108
transform -1 0 6632 0 1 3810
box -4 -6 84 206
use FILL  FILL_20_1
timestamp 1742918108
transform 1 0 6632 0 1 3810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_90
timestamp 1742918108
transform -1 0 200 0 -1 4210
box -4 -6 196 206
use XNOR2X1  XNOR2X1_3
timestamp 1742918108
transform 1 0 200 0 -1 4210
box -4 -6 116 206
use INVX1  INVX1_9
timestamp 1742918108
transform 1 0 312 0 -1 4210
box -4 -6 36 206
use AOI21X1  AOI21X1_1
timestamp 1742918108
transform -1 0 408 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_8
timestamp 1742918108
transform -1 0 440 0 -1 4210
box -4 -6 36 206
use XNOR2X1  XNOR2X1_2
timestamp 1742918108
transform -1 0 552 0 -1 4210
box -4 -6 116 206
use AOI21X1  AOI21X1_2
timestamp 1742918108
transform -1 0 616 0 -1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_6
timestamp 1742918108
transform -1 0 664 0 -1 4210
box -4 -6 52 206
use XOR2X1  XOR2X1_2
timestamp 1742918108
transform -1 0 776 0 -1 4210
box -4 -6 116 206
use INVX1  INVX1_31
timestamp 1742918108
transform 1 0 776 0 -1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_26
timestamp 1742918108
transform 1 0 808 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_4
timestamp 1742918108
transform -1 0 920 0 -1 4210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_50
timestamp 1742918108
transform 1 0 920 0 -1 4210
box -4 -6 196 206
use OR2X2  OR2X2_1
timestamp 1742918108
transform -1 0 1176 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_29
timestamp 1742918108
transform -1 0 1240 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_16
timestamp 1742918108
transform -1 0 1288 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_62
timestamp 1742918108
transform 1 0 1288 0 -1 4210
box -4 -6 52 206
use INVX1  INVX1_73
timestamp 1742918108
transform -1 0 1368 0 -1 4210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_66
timestamp 1742918108
transform -1 0 1560 0 -1 4210
box -4 -6 196 206
use OAI21X1  OAI21X1_9
timestamp 1742918108
transform -1 0 1624 0 -1 4210
box -4 -6 68 206
use AND2X2  AND2X2_1
timestamp 1742918108
transform -1 0 1688 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_76
timestamp 1742918108
transform -1 0 1720 0 -1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_36
timestamp 1742918108
transform -1 0 1768 0 -1 4210
box -4 -6 52 206
use FILL  FILL_20_0_0
timestamp 1742918108
transform -1 0 1784 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_0_1
timestamp 1742918108
transform -1 0 1800 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_0_2
timestamp 1742918108
transform -1 0 1816 0 -1 4210
box -4 -6 20 206
use OAI21X1  OAI21X1_63
timestamp 1742918108
transform -1 0 1880 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_15
timestamp 1742918108
transform -1 0 1912 0 -1 4210
box -4 -6 36 206
use XNOR2X1  XNOR2X1_4
timestamp 1742918108
transform -1 0 2024 0 -1 4210
box -4 -6 116 206
use NAND2X1  NAND2X1_11
timestamp 1742918108
transform 1 0 2024 0 -1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_5
timestamp 1742918108
transform 1 0 2072 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_10
timestamp 1742918108
transform 1 0 2120 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_17
timestamp 1742918108
transform -1 0 2216 0 -1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_12
timestamp 1742918108
transform 1 0 2216 0 -1 4210
box -4 -6 68 206
use OAI22X1  OAI22X1_4
timestamp 1742918108
transform -1 0 2360 0 -1 4210
box -4 -6 84 206
use NAND2X1  NAND2X1_28
timestamp 1742918108
transform -1 0 2408 0 -1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_6
timestamp 1742918108
transform 1 0 2408 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_53
timestamp 1742918108
transform 1 0 2472 0 -1 4210
box -4 -6 36 206
use OR2X2  OR2X2_2
timestamp 1742918108
transform 1 0 2504 0 -1 4210
box -4 -6 68 206
use BUFX4  BUFX4_3
timestamp 1742918108
transform -1 0 2632 0 -1 4210
box -4 -6 68 206
use OAI22X1  OAI22X1_6
timestamp 1742918108
transform 1 0 2632 0 -1 4210
box -4 -6 84 206
use OAI21X1  OAI21X1_72
timestamp 1742918108
transform -1 0 2776 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_12
timestamp 1742918108
transform -1 0 2824 0 -1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_13
timestamp 1742918108
transform -1 0 2872 0 -1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_48
timestamp 1742918108
transform 1 0 2872 0 -1 4210
box -4 -6 52 206
use OAI22X1  OAI22X1_2
timestamp 1742918108
transform -1 0 3000 0 -1 4210
box -4 -6 84 206
use INVX1  INVX1_20
timestamp 1742918108
transform -1 0 3032 0 -1 4210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_95
timestamp 1742918108
transform -1 0 3224 0 -1 4210
box -4 -6 196 206
use INVX1  INVX1_29
timestamp 1742918108
transform -1 0 3256 0 -1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_23
timestamp 1742918108
transform 1 0 3256 0 -1 4210
box -4 -6 68 206
use FILL  FILL_20_1_0
timestamp 1742918108
transform 1 0 3320 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_1_1
timestamp 1742918108
transform 1 0 3336 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_1_2
timestamp 1742918108
transform 1 0 3352 0 -1 4210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_103
timestamp 1742918108
transform 1 0 3368 0 -1 4210
box -4 -6 196 206
use INVX1  INVX1_24
timestamp 1742918108
transform -1 0 3592 0 -1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_48
timestamp 1742918108
transform -1 0 3640 0 -1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_60
timestamp 1742918108
transform 1 0 3640 0 -1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_58
timestamp 1742918108
transform -1 0 3736 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_80
timestamp 1742918108
transform 1 0 3736 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_76
timestamp 1742918108
transform -1 0 3864 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_45
timestamp 1742918108
transform 1 0 3864 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_74
timestamp 1742918108
transform 1 0 3912 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_75
timestamp 1742918108
transform 1 0 3976 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_42
timestamp 1742918108
transform -1 0 4088 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_43
timestamp 1742918108
transform -1 0 4136 0 -1 4210
box -4 -6 52 206
use OR2X2  OR2X2_4
timestamp 1742918108
transform 1 0 4136 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_87
timestamp 1742918108
transform 1 0 4200 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_52
timestamp 1742918108
transform -1 0 4312 0 -1 4210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_47
timestamp 1742918108
transform 1 0 4312 0 -1 4210
box -4 -6 196 206
use AND2X2  AND2X2_45
timestamp 1742918108
transform -1 0 4568 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_406
timestamp 1742918108
transform -1 0 4616 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_384
timestamp 1742918108
transform -1 0 4680 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_377
timestamp 1742918108
transform -1 0 4744 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_348
timestamp 1742918108
transform 1 0 4744 0 -1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_215
timestamp 1742918108
transform -1 0 4856 0 -1 4210
box -4 -6 52 206
use FILL  FILL_20_2_0
timestamp 1742918108
transform 1 0 4856 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_2_1
timestamp 1742918108
transform 1 0 4872 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_2_2
timestamp 1742918108
transform 1 0 4888 0 -1 4210
box -4 -6 20 206
use INVX1  INVX1_278
timestamp 1742918108
transform 1 0 4904 0 -1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_272
timestamp 1742918108
transform -1 0 5000 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_278
timestamp 1742918108
transform -1 0 5064 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_391
timestamp 1742918108
transform -1 0 5112 0 -1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_204
timestamp 1742918108
transform 1 0 5112 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_371
timestamp 1742918108
transform 1 0 5160 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_341
timestamp 1742918108
transform -1 0 5272 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_273
timestamp 1742918108
transform 1 0 5272 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_387
timestamp 1742918108
transform 1 0 5336 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_372
timestamp 1742918108
transform 1 0 5384 0 -1 4210
box -4 -6 52 206
use INVX2  INVX2_40
timestamp 1742918108
transform 1 0 5432 0 -1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_363
timestamp 1742918108
transform -1 0 5512 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_357
timestamp 1742918108
transform 1 0 5512 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_339
timestamp 1742918108
transform 1 0 5576 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_377
timestamp 1742918108
transform 1 0 5640 0 -1 4210
box -4 -6 52 206
use OR2X2  OR2X2_29
timestamp 1742918108
transform 1 0 5688 0 -1 4210
box -4 -6 68 206
use XOR2X1  XOR2X1_20
timestamp 1742918108
transform -1 0 5864 0 -1 4210
box -4 -6 116 206
use INVX1  INVX1_293
timestamp 1742918108
transform 1 0 5864 0 -1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_381
timestamp 1742918108
transform 1 0 5896 0 -1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_274
timestamp 1742918108
transform -1 0 6008 0 -1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_136
timestamp 1742918108
transform 1 0 6008 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_283
timestamp 1742918108
transform 1 0 6072 0 -1 4210
box -4 -6 36 206
use AOI21X1  AOI21X1_135
timestamp 1742918108
transform 1 0 6104 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_275
timestamp 1742918108
transform 1 0 6168 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_356
timestamp 1742918108
transform 1 0 6232 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_276
timestamp 1742918108
transform 1 0 6296 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_284
timestamp 1742918108
transform 1 0 6360 0 -1 4210
box -4 -6 36 206
use AOI21X1  AOI21X1_140
timestamp 1742918108
transform 1 0 6392 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_344
timestamp 1742918108
transform 1 0 6456 0 -1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_219
timestamp 1742918108
transform -1 0 6568 0 -1 4210
box -4 -6 52 206
use AND2X2  AND2X2_44
timestamp 1742918108
transform 1 0 6568 0 -1 4210
box -4 -6 68 206
use FILL  FILL_21_1
timestamp 1742918108
transform -1 0 6648 0 -1 4210
box -4 -6 20 206
use INVX1  INVX1_4
timestamp 1742918108
transform 1 0 8 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_4
timestamp 1742918108
transform -1 0 104 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_10
timestamp 1742918108
transform 1 0 104 0 1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_7
timestamp 1742918108
transform 1 0 136 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_11
timestamp 1742918108
transform -1 0 216 0 1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_43
timestamp 1742918108
transform -1 0 264 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_6
timestamp 1742918108
transform -1 0 312 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_8
timestamp 1742918108
transform -1 0 360 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_16
timestamp 1742918108
transform 1 0 360 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_8
timestamp 1742918108
transform -1 0 456 0 1 4210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_10
timestamp 1742918108
transform -1 0 568 0 1 4210
box -4 -6 116 206
use AOI21X1  AOI21X1_10
timestamp 1742918108
transform -1 0 632 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_5
timestamp 1742918108
transform -1 0 696 0 1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_9
timestamp 1742918108
transform 1 0 696 0 1 4210
box -4 -6 68 206
use AND2X2  AND2X2_8
timestamp 1742918108
transform 1 0 760 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_3
timestamp 1742918108
transform 1 0 824 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_6
timestamp 1742918108
transform 1 0 872 0 1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_42
timestamp 1742918108
transform -1 0 952 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_2
timestamp 1742918108
transform -1 0 1000 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_7
timestamp 1742918108
transform -1 0 1032 0 1 4210
box -4 -6 36 206
use INVX1  INVX1_32
timestamp 1742918108
transform 1 0 1032 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_25
timestamp 1742918108
transform 1 0 1064 0 1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_18
timestamp 1742918108
transform 1 0 1128 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_15
timestamp 1742918108
transform 1 0 1176 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_28
timestamp 1742918108
transform 1 0 1224 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_33
timestamp 1742918108
transform -1 0 1320 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_59
timestamp 1742918108
transform -1 0 1384 0 1 4210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_8
timestamp 1742918108
transform 1 0 1384 0 1 4210
box -4 -6 116 206
use INVX1  INVX1_45
timestamp 1742918108
transform -1 0 1528 0 1 4210
box -4 -6 36 206
use BUFX4  BUFX4_2
timestamp 1742918108
transform -1 0 1592 0 1 4210
box -4 -6 68 206
use XOR2X1  XOR2X1_3
timestamp 1742918108
transform 1 0 1592 0 1 4210
box -4 -6 116 206
use OAI21X1  OAI21X1_64
timestamp 1742918108
transform -1 0 1768 0 1 4210
box -4 -6 68 206
use FILL  FILL_21_0_0
timestamp 1742918108
transform -1 0 1784 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_0_1
timestamp 1742918108
transform -1 0 1800 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_0_2
timestamp 1742918108
transform -1 0 1816 0 1 4210
box -4 -6 20 206
use INVX1  INVX1_77
timestamp 1742918108
transform -1 0 1848 0 1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_45
timestamp 1742918108
transform -1 0 1896 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_68
timestamp 1742918108
transform -1 0 1960 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_14
timestamp 1742918108
transform 1 0 1960 0 1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_44
timestamp 1742918108
transform 1 0 1992 0 1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_3
timestamp 1742918108
transform 1 0 2040 0 1 4210
box -4 -6 52 206
use AOI21X1  AOI21X1_3
timestamp 1742918108
transform 1 0 2088 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_13
timestamp 1742918108
transform -1 0 2184 0 1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_4
timestamp 1742918108
transform -1 0 2232 0 1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_46
timestamp 1742918108
transform -1 0 2280 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_69
timestamp 1742918108
transform 1 0 2280 0 1 4210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_9
timestamp 1742918108
transform 1 0 2344 0 1 4210
box -4 -6 116 206
use NAND2X1  NAND2X1_38
timestamp 1742918108
transform -1 0 2504 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_79
timestamp 1742918108
transform -1 0 2536 0 1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_33
timestamp 1742918108
transform -1 0 2584 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_71
timestamp 1742918108
transform 1 0 2584 0 1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_47
timestamp 1742918108
transform -1 0 2696 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_81
timestamp 1742918108
transform 1 0 2696 0 1 4210
box -4 -6 36 206
use AOI21X1  AOI21X1_11
timestamp 1742918108
transform 1 0 2728 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_25
timestamp 1742918108
transform 1 0 2792 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_16
timestamp 1742918108
transform 1 0 2824 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_13
timestamp 1742918108
transform -1 0 2936 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_22
timestamp 1742918108
transform 1 0 2936 0 1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_57
timestamp 1742918108
transform -1 0 3048 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_51
timestamp 1742918108
transform 1 0 3048 0 1 4210
box -4 -6 52 206
use INVX2  INVX2_4
timestamp 1742918108
transform -1 0 3128 0 1 4210
box -4 -6 36 206
use AOI21X1  AOI21X1_15
timestamp 1742918108
transform -1 0 3192 0 1 4210
box -4 -6 68 206
use NOR3X1  NOR3X1_1
timestamp 1742918108
transform -1 0 3320 0 1 4210
box -4 -6 132 206
use FILL  FILL_21_1_0
timestamp 1742918108
transform 1 0 3320 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_1_1
timestamp 1742918108
transform 1 0 3336 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_1_2
timestamp 1742918108
transform 1 0 3352 0 1 4210
box -4 -6 20 206
use OAI21X1  OAI21X1_17
timestamp 1742918108
transform 1 0 3368 0 1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_13
timestamp 1742918108
transform 1 0 3432 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_41
timestamp 1742918108
transform 1 0 3496 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_91
timestamp 1742918108
transform -1 0 3576 0 1 4210
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_97
timestamp 1742918108
transform 1 0 3576 0 1 4210
box -4 -6 196 206
use OAI21X1  OAI21X1_81
timestamp 1742918108
transform 1 0 3768 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_47
timestamp 1742918108
transform -1 0 3880 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_77
timestamp 1742918108
transform 1 0 3880 0 1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_42
timestamp 1742918108
transform 1 0 3944 0 1 4210
box -4 -6 196 206
use AND2X2  AND2X2_6
timestamp 1742918108
transform 1 0 4136 0 1 4210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_64
timestamp 1742918108
transform -1 0 4392 0 1 4210
box -4 -6 196 206
use NAND2X1  NAND2X1_383
timestamp 1742918108
transform -1 0 4440 0 1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_290
timestamp 1742918108
transform -1 0 4504 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_293
timestamp 1742918108
transform -1 0 4568 0 1 4210
box -4 -6 68 206
use INVX2  INVX2_43
timestamp 1742918108
transform 1 0 4568 0 1 4210
box -4 -6 36 206
use AOI21X1  AOI21X1_154
timestamp 1742918108
transform 1 0 4600 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_362
timestamp 1742918108
transform -1 0 4728 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_373
timestamp 1742918108
transform 1 0 4728 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_289
timestamp 1742918108
transform 1 0 4792 0 1 4210
box -4 -6 36 206
use FILL  FILL_21_2_0
timestamp 1742918108
transform 1 0 4824 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_2_1
timestamp 1742918108
transform 1 0 4840 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_2_2
timestamp 1742918108
transform 1 0 4856 0 1 4210
box -4 -6 20 206
use OAI21X1  OAI21X1_374
timestamp 1742918108
transform 1 0 4872 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_287
timestamp 1742918108
transform 1 0 4936 0 1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_216
timestamp 1742918108
transform 1 0 4968 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_351
timestamp 1742918108
transform 1 0 5016 0 1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_210
timestamp 1742918108
transform -1 0 5128 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_342
timestamp 1742918108
transform -1 0 5192 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_373
timestamp 1742918108
transform 1 0 5192 0 1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_209
timestamp 1742918108
transform -1 0 5288 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_343
timestamp 1742918108
transform -1 0 5352 0 1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_203
timestamp 1742918108
transform -1 0 5400 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_280
timestamp 1742918108
transform 1 0 5400 0 1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_268
timestamp 1742918108
transform -1 0 5496 0 1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_212
timestamp 1742918108
transform 1 0 5496 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_374
timestamp 1742918108
transform 1 0 5544 0 1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_211
timestamp 1742918108
transform -1 0 5640 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_375
timestamp 1742918108
transform 1 0 5640 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_378
timestamp 1742918108
transform 1 0 5688 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_345
timestamp 1742918108
transform 1 0 5736 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_292
timestamp 1742918108
transform 1 0 5800 0 1 4210
box -4 -6 36 206
use AOI21X1  AOI21X1_139
timestamp 1742918108
transform -1 0 5896 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_282
timestamp 1742918108
transform -1 0 5928 0 1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_376
timestamp 1742918108
transform 1 0 5928 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_379
timestamp 1742918108
transform 1 0 5976 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_380
timestamp 1742918108
transform 1 0 6024 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_281
timestamp 1742918108
transform 1 0 6072 0 1 4210
box -4 -6 36 206
use INVX1  INVX1_305
timestamp 1742918108
transform 1 0 6104 0 1 4210
box -4 -6 36 206
use AOI21X1  AOI21X1_146
timestamp 1742918108
transform -1 0 6200 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_400
timestamp 1742918108
transform 1 0 6200 0 1 4210
box -4 -6 52 206
use AOI21X1  AOI21X1_141
timestamp 1742918108
transform -1 0 6312 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_397
timestamp 1742918108
transform -1 0 6360 0 1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_288
timestamp 1742918108
transform -1 0 6424 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_286
timestamp 1742918108
transform 1 0 6424 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_289
timestamp 1742918108
transform -1 0 6552 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_399
timestamp 1742918108
transform -1 0 6600 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_396
timestamp 1742918108
transform -1 0 6648 0 1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_1
timestamp 1742918108
transform -1 0 72 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_1
timestamp 1742918108
transform -1 0 120 0 -1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_1
timestamp 1742918108
transform 1 0 120 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_3
timestamp 1742918108
transform -1 0 248 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_3
timestamp 1742918108
transform 1 0 248 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_58
timestamp 1742918108
transform 1 0 312 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_5
timestamp 1742918108
transform -1 0 440 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_74
timestamp 1742918108
transform 1 0 440 0 -1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_60
timestamp 1742918108
transform 1 0 472 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_4
timestamp 1742918108
transform -1 0 600 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_21
timestamp 1742918108
transform -1 0 648 0 -1 4610
box -4 -6 52 206
use XNOR2X1  XNOR2X1_6
timestamp 1742918108
transform 1 0 648 0 -1 4610
box -4 -6 116 206
use NAND2X1  NAND2X1_18
timestamp 1742918108
transform 1 0 760 0 -1 4610
box -4 -6 52 206
use XNOR2X1  XNOR2X1_7
timestamp 1742918108
transform 1 0 808 0 -1 4610
box -4 -6 116 206
use INVX1  INVX1_40
timestamp 1742918108
transform -1 0 952 0 -1 4610
box -4 -6 36 206
use AND2X2  AND2X2_2
timestamp 1742918108
transform 1 0 952 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_4
timestamp 1742918108
transform 1 0 1016 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_35
timestamp 1742918108
transform 1 0 1080 0 -1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_30
timestamp 1742918108
transform 1 0 1112 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_27
timestamp 1742918108
transform -1 0 1240 0 -1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_19
timestamp 1742918108
transform 1 0 1240 0 -1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_32
timestamp 1742918108
transform -1 0 1336 0 -1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_20
timestamp 1742918108
transform -1 0 1384 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_34
timestamp 1742918108
transform -1 0 1416 0 -1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_36
timestamp 1742918108
transform -1 0 1480 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_46
timestamp 1742918108
transform -1 0 1512 0 -1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_27
timestamp 1742918108
transform 1 0 1512 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_60
timestamp 1742918108
transform 1 0 1560 0 -1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_24
timestamp 1742918108
transform -1 0 1640 0 -1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_38
timestamp 1742918108
transform 1 0 1640 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_5
timestamp 1742918108
transform 1 0 1704 0 -1 4610
box -4 -6 68 206
use FILL  FILL_22_0_0
timestamp 1742918108
transform 1 0 1768 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_0_1
timestamp 1742918108
transform 1 0 1784 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_0_2
timestamp 1742918108
transform 1 0 1800 0 -1 4610
box -4 -6 20 206
use INVX1  INVX1_19
timestamp 1742918108
transform 1 0 1816 0 -1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_7
timestamp 1742918108
transform 1 0 1848 0 -1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_9
timestamp 1742918108
transform 1 0 1896 0 -1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_66
timestamp 1742918108
transform 1 0 1944 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_67
timestamp 1742918108
transform -1 0 2072 0 -1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_8
timestamp 1742918108
transform -1 0 2120 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_18
timestamp 1742918108
transform -1 0 2152 0 -1 4610
box -4 -6 36 206
use INVX1  INVX1_50
timestamp 1742918108
transform 1 0 2152 0 -1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_27
timestamp 1742918108
transform -1 0 2232 0 -1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_30
timestamp 1742918108
transform 1 0 2232 0 -1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_39
timestamp 1742918108
transform 1 0 2280 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_41
timestamp 1742918108
transform 1 0 2344 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_51
timestamp 1742918108
transform 1 0 2408 0 -1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_32
timestamp 1742918108
transform 1 0 2440 0 -1 4610
box -4 -6 52 206
use INVX2  INVX2_1
timestamp 1742918108
transform 1 0 2488 0 -1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_10
timestamp 1742918108
transform 1 0 2520 0 -1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_12
timestamp 1742918108
transform 1 0 2568 0 -1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_11
timestamp 1742918108
transform -1 0 2664 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_21
timestamp 1742918108
transform -1 0 2696 0 -1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_13
timestamp 1742918108
transform 1 0 2696 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_23
timestamp 1742918108
transform 1 0 2760 0 -1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_14
timestamp 1742918108
transform 1 0 2792 0 -1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_73
timestamp 1742918108
transform 1 0 2840 0 -1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_15
timestamp 1742918108
transform -1 0 2952 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_22
timestamp 1742918108
transform 1 0 2952 0 -1 4610
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_102
timestamp 1742918108
transform 1 0 2984 0 -1 4610
box -4 -6 196 206
use NOR2X1  NOR2X1_62
timestamp 1742918108
transform 1 0 3176 0 -1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_84
timestamp 1742918108
transform -1 0 3288 0 -1 4610
box -4 -6 68 206
use FILL  FILL_22_1_0
timestamp 1742918108
transform -1 0 3304 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_1_1
timestamp 1742918108
transform -1 0 3320 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_1_2
timestamp 1742918108
transform -1 0 3336 0 -1 4610
box -4 -6 20 206
use OAI21X1  OAI21X1_85
timestamp 1742918108
transform -1 0 3400 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_28
timestamp 1742918108
transform 1 0 3400 0 -1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_21
timestamp 1742918108
transform -1 0 3496 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_7
timestamp 1742918108
transform 1 0 3496 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_86
timestamp 1742918108
transform 1 0 3560 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_50
timestamp 1742918108
transform -1 0 3672 0 -1 4610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_46
timestamp 1742918108
transform 1 0 3672 0 -1 4610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_44
timestamp 1742918108
transform 1 0 3864 0 -1 4610
box -4 -6 196 206
use AND2X2  AND2X2_9
timestamp 1742918108
transform 1 0 4056 0 -1 4610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_7
timestamp 1742918108
transform 1 0 4120 0 -1 4610
box -4 -6 148 206
use NAND2X1  NAND2X1_404
timestamp 1742918108
transform 1 0 4264 0 -1 4610
box -4 -6 52 206
use AOI22X1  AOI22X1_47
timestamp 1742918108
transform 1 0 4312 0 -1 4610
box -4 -6 84 206
use OAI21X1  OAI21X1_360
timestamp 1742918108
transform 1 0 4392 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_295
timestamp 1742918108
transform 1 0 4456 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_294
timestamp 1742918108
transform 1 0 4520 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_296
timestamp 1742918108
transform -1 0 4616 0 -1 4610
box -4 -6 36 206
use NAND3X1  NAND3X1_291
timestamp 1742918108
transform 1 0 4616 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_408
timestamp 1742918108
transform -1 0 4728 0 -1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_361
timestamp 1742918108
transform 1 0 4728 0 -1 4610
box -4 -6 68 206
use AOI22X1  AOI22X1_49
timestamp 1742918108
transform 1 0 4792 0 -1 4610
box -4 -6 84 206
use FILL  FILL_22_2_0
timestamp 1742918108
transform 1 0 4872 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_2_1
timestamp 1742918108
transform 1 0 4888 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_2_2
timestamp 1742918108
transform 1 0 4904 0 -1 4610
box -4 -6 20 206
use NAND3X1  NAND3X1_292
timestamp 1742918108
transform 1 0 4920 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_389
timestamp 1742918108
transform -1 0 5032 0 -1 4610
box -4 -6 52 206
use INVX2  INVX2_42
timestamp 1742918108
transform 1 0 5032 0 -1 4610
box -4 -6 36 206
use NAND3X1  NAND3X1_296
timestamp 1742918108
transform -1 0 5128 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_142
timestamp 1742918108
transform 1 0 5128 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_386
timestamp 1742918108
transform 1 0 5192 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_279
timestamp 1742918108
transform -1 0 5288 0 -1 4610
box -4 -6 36 206
use INVX2  INVX2_41
timestamp 1742918108
transform -1 0 5320 0 -1 4610
box -4 -6 36 206
use INVX2  INVX2_39
timestamp 1742918108
transform -1 0 5352 0 -1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_346
timestamp 1742918108
transform -1 0 5416 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_347
timestamp 1742918108
transform 1 0 5416 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_138
timestamp 1742918108
transform -1 0 5544 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_286
timestamp 1742918108
transform 1 0 5544 0 -1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_213
timestamp 1742918108
transform -1 0 5624 0 -1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_214
timestamp 1742918108
transform -1 0 5672 0 -1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_280
timestamp 1742918108
transform -1 0 5736 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_392
timestamp 1742918108
transform 1 0 5736 0 -1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_223
timestamp 1742918108
transform 1 0 5784 0 -1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_279
timestamp 1742918108
transform -1 0 5896 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_393
timestamp 1742918108
transform -1 0 5944 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_288
timestamp 1742918108
transform 1 0 5944 0 -1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_395
timestamp 1742918108
transform 1 0 5976 0 -1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_352
timestamp 1742918108
transform 1 0 6024 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_354
timestamp 1742918108
transform 1 0 6088 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_353
timestamp 1742918108
transform -1 0 6216 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_355
timestamp 1742918108
transform 1 0 6216 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_285
timestamp 1742918108
transform 1 0 6280 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_282
timestamp 1742918108
transform -1 0 6408 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_284
timestamp 1742918108
transform 1 0 6408 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_281
timestamp 1742918108
transform 1 0 6472 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_287
timestamp 1742918108
transform 1 0 6536 0 -1 4610
box -4 -6 68 206
use FILL  FILL_23_1
timestamp 1742918108
transform -1 0 6616 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_2
timestamp 1742918108
transform -1 0 6632 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_3
timestamp 1742918108
transform -1 0 6648 0 -1 4610
box -4 -6 20 206
use XOR2X1  XOR2X1_1
timestamp 1742918108
transform 1 0 8 0 1 4610
box -4 -6 116 206
use NOR2X1  NOR2X1_1
timestamp 1742918108
transform 1 0 120 0 1 4610
box -4 -6 52 206
use INVX1  INVX1_2
timestamp 1742918108
transform -1 0 200 0 1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_2
timestamp 1742918108
transform 1 0 200 0 1 4610
box -4 -6 52 206
use INVX1  INVX1_3
timestamp 1742918108
transform 1 0 248 0 1 4610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_1
timestamp 1742918108
transform 1 0 280 0 1 4610
box -4 -6 116 206
use INVX1  INVX1_5
timestamp 1742918108
transform 1 0 392 0 1 4610
box -4 -6 36 206
use INVX1  INVX1_38
timestamp 1742918108
transform 1 0 424 0 1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_20
timestamp 1742918108
transform 1 0 456 0 1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_41
timestamp 1742918108
transform -1 0 552 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_19
timestamp 1742918108
transform 1 0 552 0 1 4610
box -4 -6 52 206
use INVX1  INVX1_39
timestamp 1742918108
transform -1 0 632 0 1 4610
box -4 -6 36 206
use AOI21X1  AOI21X1_7
timestamp 1742918108
transform -1 0 696 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_36
timestamp 1742918108
transform 1 0 696 0 1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_40
timestamp 1742918108
transform -1 0 776 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_32
timestamp 1742918108
transform -1 0 840 0 1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_23
timestamp 1742918108
transform 1 0 840 0 1 4610
box -4 -6 52 206
use INVX1  INVX1_37
timestamp 1742918108
transform -1 0 920 0 1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_22
timestamp 1742918108
transform 1 0 920 0 1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_24
timestamp 1742918108
transform -1 0 1016 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_34
timestamp 1742918108
transform -1 0 1080 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_42
timestamp 1742918108
transform -1 0 1112 0 1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_42
timestamp 1742918108
transform 1 0 1112 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_43
timestamp 1742918108
transform -1 0 1240 0 1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_21
timestamp 1742918108
transform 1 0 1240 0 1 4610
box -4 -6 52 206
use AOI21X1  AOI21X1_6
timestamp 1742918108
transform 1 0 1288 0 1 4610
box -4 -6 68 206
use AND2X2  AND2X2_7
timestamp 1742918108
transform 1 0 1352 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_62
timestamp 1742918108
transform -1 0 1448 0 1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_45
timestamp 1742918108
transform 1 0 1448 0 1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_25
timestamp 1742918108
transform 1 0 1512 0 1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_2
timestamp 1742918108
transform -1 0 1624 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_43
timestamp 1742918108
transform 1 0 1624 0 1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_26
timestamp 1742918108
transform 1 0 1656 0 1 4610
box -4 -6 52 206
use INVX1  INVX1_44
timestamp 1742918108
transform -1 0 1736 0 1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_29
timestamp 1742918108
transform -1 0 1784 0 1 4610
box -4 -6 52 206
use FILL  FILL_23_0_0
timestamp 1742918108
transform 1 0 1784 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_0_1
timestamp 1742918108
transform 1 0 1800 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_0_2
timestamp 1742918108
transform 1 0 1816 0 1 4610
box -4 -6 20 206
use NOR2X1  NOR2X1_28
timestamp 1742918108
transform 1 0 1832 0 1 4610
box -4 -6 52 206
use AND2X2  AND2X2_4
timestamp 1742918108
transform -1 0 1944 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_61
timestamp 1742918108
transform 1 0 1944 0 1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_44
timestamp 1742918108
transform 1 0 1976 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_46
timestamp 1742918108
transform 1 0 2040 0 1 4610
box -4 -6 68 206
use AND2X2  AND2X2_5
timestamp 1742918108
transform -1 0 2168 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_26
timestamp 1742918108
transform 1 0 2168 0 1 4610
box -4 -6 52 206
use INVX1  INVX1_48
timestamp 1742918108
transform 1 0 2216 0 1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_25
timestamp 1742918108
transform -1 0 2296 0 1 4610
box -4 -6 52 206
use INVX1  INVX1_49
timestamp 1742918108
transform -1 0 2328 0 1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_31
timestamp 1742918108
transform 1 0 2328 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_47
timestamp 1742918108
transform 1 0 2376 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_48
timestamp 1742918108
transform -1 0 2504 0 1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_31
timestamp 1742918108
transform 1 0 2504 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_29
timestamp 1742918108
transform -1 0 2600 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_33
timestamp 1742918108
transform -1 0 2648 0 1 4610
box -4 -6 52 206
use AOI21X1  AOI21X1_8
timestamp 1742918108
transform -1 0 2712 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_64
timestamp 1742918108
transform -1 0 2744 0 1 4610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_5
timestamp 1742918108
transform 1 0 2744 0 1 4610
box -4 -6 116 206
use NOR2X1  NOR2X1_16
timestamp 1742918108
transform 1 0 2856 0 1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_17
timestamp 1742918108
transform 1 0 2904 0 1 4610
box -4 -6 52 206
use INVX1  INVX1_26
timestamp 1742918108
transform 1 0 2952 0 1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_15
timestamp 1742918108
transform 1 0 2984 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_14
timestamp 1742918108
transform 1 0 3048 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_14
timestamp 1742918108
transform -1 0 3160 0 1 4610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_96
timestamp 1742918108
transform 1 0 3160 0 1 4610
box -4 -6 196 206
use FILL  FILL_23_1_0
timestamp 1742918108
transform 1 0 3352 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_1_1
timestamp 1742918108
transform 1 0 3368 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_1_2
timestamp 1742918108
transform 1 0 3384 0 1 4610
box -4 -6 20 206
use INVX1  INVX1_90
timestamp 1742918108
transform 1 0 3400 0 1 4610
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_101
timestamp 1742918108
transform 1 0 3432 0 1 4610
box -4 -6 196 206
use OAI21X1  OAI21X1_82
timestamp 1742918108
transform -1 0 3688 0 1 4610
box -4 -6 68 206
use AND2X2  AND2X2_11
timestamp 1742918108
transform 1 0 3688 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_83
timestamp 1742918108
transform 1 0 3752 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_49
timestamp 1742918108
transform -1 0 3864 0 1 4610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_45
timestamp 1742918108
transform 1 0 3864 0 1 4610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_80
timestamp 1742918108
transform 1 0 4056 0 1 4610
box -4 -6 196 206
use NAND2X1  NAND2X1_405
timestamp 1742918108
transform 1 0 4248 0 1 4610
box -4 -6 52 206
use OR2X2  OR2X2_32
timestamp 1742918108
transform 1 0 4296 0 1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_221
timestamp 1742918108
transform -1 0 4408 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_409
timestamp 1742918108
transform 1 0 4408 0 1 4610
box -4 -6 52 206
use AOI22X1  AOI22X1_48
timestamp 1742918108
transform -1 0 4536 0 1 4610
box -4 -6 84 206
use NAND2X1  NAND2X1_407
timestamp 1742918108
transform 1 0 4536 0 1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_222
timestamp 1742918108
transform 1 0 4584 0 1 4610
box -4 -6 52 206
use NOR3X1  NOR3X1_12
timestamp 1742918108
transform -1 0 4760 0 1 4610
box -4 -6 132 206
use OAI21X1  OAI21X1_364
timestamp 1742918108
transform 1 0 4760 0 1 4610
box -4 -6 68 206
use FILL  FILL_23_2_0
timestamp 1742918108
transform 1 0 4824 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_2_1
timestamp 1742918108
transform 1 0 4840 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_2_2
timestamp 1742918108
transform 1 0 4856 0 1 4610
box -4 -6 20 206
use OAI21X1  OAI21X1_370
timestamp 1742918108
transform 1 0 4872 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_363
timestamp 1742918108
transform 1 0 4936 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_297
timestamp 1742918108
transform 1 0 5000 0 1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_410
timestamp 1742918108
transform -1 0 5080 0 1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_297
timestamp 1742918108
transform 1 0 5080 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_326
timestamp 1742918108
transform -1 0 5208 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_423
timestamp 1742918108
transform 1 0 5208 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_359
timestamp 1742918108
transform 1 0 5256 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_382
timestamp 1742918108
transform -1 0 5368 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_384
timestamp 1742918108
transform -1 0 5416 0 1 4610
box -4 -6 52 206
use OR2X2  OR2X2_30
timestamp 1742918108
transform 1 0 5416 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_385
timestamp 1742918108
transform 1 0 5480 0 1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_277
timestamp 1742918108
transform -1 0 5592 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_285
timestamp 1742918108
transform 1 0 5592 0 1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_386
timestamp 1742918108
transform 1 0 5624 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_394
timestamp 1742918108
transform 1 0 5672 0 1 4610
box -4 -6 52 206
use OR2X2  OR2X2_31
timestamp 1742918108
transform 1 0 5720 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_304
timestamp 1742918108
transform -1 0 5816 0 1 4610
box -4 -6 36 206
use AOI22X1  AOI22X1_45
timestamp 1742918108
transform -1 0 5896 0 1 4610
box -4 -6 84 206
use AOI22X1  AOI22X1_43
timestamp 1742918108
transform -1 0 5976 0 1 4610
box -4 -6 84 206
use AOI22X1  AOI22X1_44
timestamp 1742918108
transform -1 0 6056 0 1 4610
box -4 -6 84 206
use AOI22X1  AOI22X1_46
timestamp 1742918108
transform 1 0 6056 0 1 4610
box -4 -6 84 206
use NAND2X1  NAND2X1_403
timestamp 1742918108
transform -1 0 6184 0 1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_358
timestamp 1742918108
transform -1 0 6248 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_402
timestamp 1742918108
transform -1 0 6296 0 1 4610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_134
timestamp 1742918108
transform 1 0 6296 0 1 4610
box -4 -6 196 206
use NAND3X1  NAND3X1_48
timestamp 1742918108
transform 1 0 6488 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_1
timestamp 1742918108
transform 1 0 6552 0 1 4610
box -4 -6 52 206
use FILL  FILL_24_1
timestamp 1742918108
transform 1 0 6600 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_2
timestamp 1742918108
transform 1 0 6616 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_3
timestamp 1742918108
transform 1 0 6632 0 1 4610
box -4 -6 20 206
<< labels >>
flabel metal4 s 1768 -40 1816 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 3304 -40 3352 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -19 4497 -13 4503 7 FreeSans 24 0 0 0 clk
port 2 nsew
flabel metal3 s 6669 3777 6675 3783 6 FreeSans 24 0 0 0 reset
port 3 nsew
flabel metal2 s 2989 4837 2995 4843 3 FreeSans 24 90 0 0 start
port 4 nsew
flabel metal3 s -19 4537 -13 4543 7 FreeSans 24 0 0 0 x0[0]
port 5 nsew
flabel metal3 s -19 4577 -13 4583 7 FreeSans 24 0 0 0 x0[1]
port 6 nsew
flabel metal3 s -19 4617 -13 4623 7 FreeSans 24 0 0 0 x0[2]
port 7 nsew
flabel metal3 s -19 4657 -13 4663 7 FreeSans 24 0 0 0 x0[3]
port 8 nsew
flabel metal3 s -19 4697 -13 4703 7 FreeSans 24 0 0 0 x0[4]
port 9 nsew
flabel metal3 s -19 4737 -13 4743 7 FreeSans 24 0 0 0 x0[5]
port 10 nsew
flabel metal3 s -19 4777 -13 4783 7 FreeSans 24 0 0 0 x0[6]
port 11 nsew
flabel metal3 s -19 4817 -13 4823 7 FreeSans 24 90 0 0 x0[7]
port 12 nsew
flabel metal3 s -19 4177 -13 4183 7 FreeSans 24 0 0 0 x1[0]
port 13 nsew
flabel metal3 s -19 4217 -13 4223 7 FreeSans 24 0 0 0 x1[1]
port 14 nsew
flabel metal3 s -19 4257 -13 4263 7 FreeSans 24 0 0 0 x1[2]
port 15 nsew
flabel metal3 s -19 4297 -13 4303 7 FreeSans 24 0 0 0 x1[3]
port 16 nsew
flabel metal3 s -19 4337 -13 4343 7 FreeSans 24 0 0 0 x1[4]
port 17 nsew
flabel metal3 s -19 4377 -13 4383 7 FreeSans 24 0 0 0 x1[5]
port 18 nsew
flabel metal3 s -19 4417 -13 4423 7 FreeSans 24 0 0 0 x1[6]
port 19 nsew
flabel metal3 s -19 4457 -13 4463 7 FreeSans 24 0 0 0 x1[7]
port 20 nsew
flabel metal2 s 3021 4837 3027 4843 3 FreeSans 24 90 0 0 x2[0]
port 21 nsew
flabel metal2 s 3053 4837 3059 4843 3 FreeSans 24 90 0 0 x2[1]
port 22 nsew
flabel metal2 s 3085 4837 3091 4843 3 FreeSans 24 90 0 0 x2[2]
port 23 nsew
flabel metal2 s 3117 4837 3123 4843 3 FreeSans 24 90 0 0 x2[3]
port 24 nsew
flabel metal2 s 3149 4837 3155 4843 3 FreeSans 24 90 0 0 x2[4]
port 25 nsew
flabel metal2 s 3181 4837 3187 4843 3 FreeSans 24 90 0 0 x2[5]
port 26 nsew
flabel metal2 s 3213 4837 3219 4843 3 FreeSans 24 90 0 0 x2[6]
port 27 nsew
flabel metal2 s 3245 4837 3251 4843 3 FreeSans 24 90 0 0 x2[7]
port 28 nsew
flabel metal2 s 205 4837 211 4843 3 FreeSans 24 90 0 0 x3[0]
port 29 nsew
flabel metal2 s 253 4837 259 4843 3 FreeSans 24 90 0 0 x3[1]
port 30 nsew
flabel metal2 s 989 4837 995 4843 3 FreeSans 24 90 0 0 x3[2]
port 31 nsew
flabel metal2 s 1021 4837 1027 4843 3 FreeSans 24 90 0 0 x3[3]
port 32 nsew
flabel metal2 s 2205 4837 2211 4843 3 FreeSans 24 90 0 0 x3[4]
port 33 nsew
flabel metal2 s 2237 4837 2243 4843 3 FreeSans 24 90 0 0 x3[5]
port 34 nsew
flabel metal2 s 2653 4837 2659 4843 3 FreeSans 24 90 0 0 x3[6]
port 35 nsew
flabel metal2 s 2957 4837 2963 4843 3 FreeSans 24 90 0 0 x3[7]
port 36 nsew
flabel metal3 s 6669 4537 6675 4543 6 FreeSans 24 0 0 0 X0_mag[0]
port 37 nsew
flabel metal3 s 6669 4577 6675 4583 6 FreeSans 24 0 0 0 X0_mag[1]
port 38 nsew
flabel metal3 s 6669 4617 6675 4623 6 FreeSans 24 0 0 0 X0_mag[2]
port 39 nsew
flabel metal3 s 6669 4657 6675 4663 6 FreeSans 24 0 0 0 X0_mag[3]
port 40 nsew
flabel metal3 s 6669 4697 6675 4703 6 FreeSans 24 0 0 0 X0_mag[4]
port 41 nsew
flabel metal3 s 6669 4737 6675 4743 6 FreeSans 24 0 0 0 X0_mag[5]
port 42 nsew
flabel metal3 s 6669 4777 6675 4783 6 FreeSans 24 0 0 0 X0_mag[6]
port 43 nsew
flabel metal3 s 6669 4817 6675 4823 3 FreeSans 24 90 0 0 X0_mag[7]
port 44 nsew
flabel metal3 s 6669 2697 6675 2703 6 FreeSans 24 0 0 0 X1_mag[0]
port 45 nsew
flabel metal3 s 6669 2897 6675 2903 6 FreeSans 24 0 0 0 X1_mag[1]
port 46 nsew
flabel metal3 s 6669 2937 6675 2943 6 FreeSans 24 0 0 0 X1_mag[2]
port 47 nsew
flabel metal3 s 6669 3097 6675 3103 6 FreeSans 24 0 0 0 X1_mag[3]
port 48 nsew
flabel metal3 s 6669 3297 6675 3303 6 FreeSans 24 0 0 0 X1_mag[4]
port 49 nsew
flabel metal3 s 6669 3337 6675 3343 6 FreeSans 24 0 0 0 X1_mag[5]
port 50 nsew
flabel metal3 s 6669 3697 6675 3703 6 FreeSans 24 0 0 0 X1_mag[6]
port 51 nsew
flabel metal3 s 6669 3737 6675 3743 6 FreeSans 24 0 0 0 X1_mag[7]
port 52 nsew
flabel metal2 s 4189 -23 4195 -17 7 FreeSans 24 270 0 0 X2_mag[0]
port 53 nsew
flabel metal2 s 4237 -23 4243 -17 7 FreeSans 24 270 0 0 X2_mag[1]
port 54 nsew
flabel metal2 s 4477 -23 4483 -17 7 FreeSans 24 270 0 0 X2_mag[2]
port 55 nsew
flabel metal2 s 5117 -23 5123 -17 7 FreeSans 24 270 0 0 X2_mag[3]
port 56 nsew
flabel metal2 s 5549 -23 5555 -17 7 FreeSans 24 270 0 0 X2_mag[4]
port 57 nsew
flabel metal2 s 5693 -23 5699 -17 7 FreeSans 24 270 0 0 X2_mag[5]
port 58 nsew
flabel metal2 s 6269 -23 6275 -17 7 FreeSans 24 270 0 0 X2_mag[6]
port 59 nsew
flabel metal2 s 6301 -23 6307 -17 7 FreeSans 24 270 0 0 X2_mag[7]
port 60 nsew
flabel metal2 s 6333 -23 6339 -17 7 FreeSans 24 270 0 0 X3_mag[0]
port 61 nsew
flabel metal2 s 6365 -23 6371 -17 7 FreeSans 24 270 0 0 X3_mag[1]
port 62 nsew
flabel metal2 s 6397 -23 6403 -17 7 FreeSans 24 270 0 0 X3_mag[2]
port 63 nsew
flabel metal2 s 6461 -23 6467 -17 7 FreeSans 24 270 0 0 X3_mag[3]
port 64 nsew
flabel metal2 s 6493 -23 6499 -17 7 FreeSans 24 270 0 0 X3_mag[4]
port 65 nsew
flabel metal2 s 6541 -23 6547 -17 7 FreeSans 24 270 0 0 X3_mag[5]
port 66 nsew
flabel metal2 s 6573 -23 6579 -17 7 FreeSans 24 270 0 0 X3_mag[6]
port 67 nsew
flabel metal2 s 6605 -23 6611 -17 7 FreeSans 24 270 0 0 X3_mag[7]
port 68 nsew
flabel metal2 s 6637 -23 6643 -17 7 FreeSans 24 270 0 0 done
port 69 nsew
<< end >>

magic
tech scmos
magscale 1 2
timestamp 1739819275
<< checkpaint >>
rect -70 -66 116 270
<< nwell >>
rect -10 96 56 210
<< ntransistor >>
rect 14 12 18 32
rect 30 12 34 52
<< ptransistor >>
rect 14 148 18 188
rect 30 108 34 188
<< ndiffusion >>
rect 20 51 30 52
rect 4 31 14 32
rect 12 13 14 31
rect 4 12 14 13
rect 18 13 20 32
rect 28 13 30 51
rect 18 12 30 13
rect 34 51 44 52
rect 34 13 36 51
rect 34 12 44 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 149 14 187
rect 4 148 14 149
rect 18 148 20 188
rect 28 120 30 188
rect 20 108 30 120
rect 34 187 44 188
rect 34 109 36 187
rect 34 108 44 109
<< ndcontact >>
rect 4 13 12 31
rect 20 13 28 51
rect 36 13 44 51
<< pdcontact >>
rect 4 149 12 187
rect 20 120 28 188
rect 36 109 44 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 14 114 18 148
rect 12 110 18 114
rect 12 82 16 110
rect 30 102 34 108
rect 32 94 34 102
rect 12 78 18 82
rect 14 32 18 78
rect 30 52 34 94
rect 14 8 18 12
rect 30 8 34 12
<< polycontact >>
rect 4 78 12 86
rect 24 94 32 102
<< metal1 >>
rect -4 204 52 206
rect 4 196 28 204
rect 36 196 52 204
rect -4 194 52 196
rect 20 188 28 194
rect 4 187 12 188
rect 4 114 12 149
rect 36 187 44 188
rect 4 108 26 114
rect 36 108 44 109
rect 20 102 26 108
rect 20 94 24 102
rect 4 86 12 94
rect 20 64 26 94
rect 38 86 44 108
rect 4 58 26 64
rect 4 31 12 58
rect 4 12 12 13
rect 20 51 28 52
rect 20 6 28 13
rect 36 51 44 86
rect 36 12 44 13
rect -4 4 52 6
rect 4 -4 28 4
rect 36 -4 52 4
rect -4 -6 52 -4
<< m1p >>
rect 4 86 12 94
rect 36 66 44 74
<< labels >>
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 90 8 90 4 A
rlabel metal1 40 70 40 70 4 Y
<< end >>

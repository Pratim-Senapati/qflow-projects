magic
tech scmos
magscale 1 2
timestamp 1740382396
<< nwell >>
rect -10 96 168 210
<< ntransistor >>
rect 14 12 18 52
rect 24 12 28 52
rect 56 12 60 32
rect 72 12 76 52
rect 88 12 92 52
rect 104 12 108 52
rect 136 12 140 32
<< ptransistor >>
rect 14 148 18 188
rect 30 148 34 188
rect 62 148 66 188
rect 78 148 82 188
rect 94 108 98 188
rect 104 108 108 188
rect 136 148 140 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 12 24 52
rect 28 51 38 52
rect 28 13 30 51
rect 66 50 72 52
rect 28 12 38 13
rect 46 31 56 32
rect 54 13 56 31
rect 46 12 56 13
rect 60 12 62 32
rect 70 12 72 50
rect 76 51 88 52
rect 76 13 78 51
rect 86 13 88 51
rect 76 12 88 13
rect 92 24 94 52
rect 102 24 104 52
rect 92 12 104 24
rect 108 48 114 52
rect 108 44 118 48
rect 108 16 110 44
rect 108 12 118 16
rect 126 31 136 32
rect 134 13 136 31
rect 126 12 136 13
rect 140 31 150 32
rect 140 13 142 31
rect 140 12 150 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 149 14 187
rect 4 148 14 149
rect 18 184 30 188
rect 18 156 20 184
rect 28 156 30 184
rect 18 148 30 156
rect 34 187 44 188
rect 34 149 36 187
rect 34 148 44 149
rect 52 187 62 188
rect 60 149 62 187
rect 52 148 62 149
rect 66 187 78 188
rect 66 149 68 187
rect 76 149 78 187
rect 66 148 78 149
rect 82 187 94 188
rect 82 148 84 187
rect 92 109 94 187
rect 84 108 94 109
rect 98 108 104 188
rect 108 187 118 188
rect 108 109 110 187
rect 126 187 136 188
rect 134 149 136 187
rect 126 148 136 149
rect 140 187 150 188
rect 140 149 142 187
rect 140 148 150 149
rect 108 108 118 109
<< ndcontact >>
rect 4 13 12 51
rect 30 13 38 51
rect 46 13 54 31
rect 62 12 70 50
rect 78 13 86 51
rect 94 24 102 52
rect 110 16 118 44
rect 126 13 134 31
rect 142 13 150 31
<< pdcontact >>
rect 4 149 12 187
rect 20 156 28 184
rect 36 149 44 187
rect 52 149 60 187
rect 68 149 76 187
rect 84 109 92 187
rect 110 109 118 187
rect 126 149 134 187
rect 142 149 150 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
rect 92 -4 100 4
rect 124 -4 132 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
rect 92 196 100 204
rect 124 196 132 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 62 188 66 192
rect 78 188 82 192
rect 94 188 98 192
rect 104 188 108 192
rect 136 188 140 192
rect 14 146 18 148
rect 12 142 18 146
rect 12 66 16 142
rect 30 80 34 148
rect 32 72 34 80
rect 16 58 18 64
rect 30 58 34 72
rect 62 146 66 148
rect 78 146 82 148
rect 62 142 82 146
rect 62 58 66 142
rect 136 146 140 148
rect 126 142 140 146
rect 94 104 98 108
rect 88 100 98 104
rect 88 86 92 100
rect 14 52 18 58
rect 24 54 34 58
rect 56 54 76 58
rect 24 52 28 54
rect 56 32 60 54
rect 72 52 76 54
rect 88 52 92 78
rect 104 74 108 108
rect 104 52 108 66
rect 126 38 130 142
rect 126 34 140 38
rect 136 32 140 34
rect 14 8 18 12
rect 24 8 28 12
rect 56 8 60 12
rect 72 8 76 12
rect 88 8 92 12
rect 104 8 108 12
rect 136 8 140 12
<< polycontact >>
rect 24 72 32 80
rect 8 58 16 66
rect 84 78 92 86
rect 48 46 56 54
rect 100 66 108 74
rect 118 54 126 62
<< metal1 >>
rect -4 204 164 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 92 204
rect 100 196 124 204
rect 132 196 164 204
rect -4 194 164 196
rect 4 187 12 188
rect 20 184 28 194
rect 20 152 28 156
rect 36 187 44 188
rect 4 148 12 149
rect 6 146 12 148
rect 36 146 44 149
rect 6 140 44 146
rect 20 86 28 94
rect 38 92 44 140
rect 52 187 60 188
rect 52 92 60 149
rect 68 187 76 194
rect 68 148 76 149
rect 84 187 92 188
rect 84 108 92 109
rect 110 187 118 194
rect 126 187 134 194
rect 126 148 134 149
rect 142 187 150 188
rect 142 148 150 149
rect 144 142 150 148
rect 134 136 150 142
rect 134 114 140 136
rect 110 108 118 109
rect 86 102 92 108
rect 132 106 140 114
rect 86 96 120 102
rect 22 80 30 86
rect 4 66 12 74
rect 72 78 84 84
rect 32 72 78 78
rect 84 66 100 72
rect 4 60 8 66
rect 16 60 90 66
rect 114 62 120 96
rect 114 60 118 62
rect 96 54 118 60
rect 4 51 12 52
rect 4 6 12 13
rect 30 51 38 52
rect 46 46 48 54
rect 96 52 102 54
rect 78 51 86 52
rect 30 12 38 13
rect 46 31 54 32
rect 46 12 54 13
rect 110 44 118 48
rect 86 16 110 18
rect 134 46 140 106
rect 134 40 150 46
rect 144 32 150 40
rect 86 13 118 16
rect 78 12 118 13
rect 126 31 134 32
rect 62 6 70 12
rect 126 6 134 13
rect 142 31 150 32
rect 142 12 150 13
rect -4 4 164 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 92 4
rect 100 -4 124 4
rect 132 -4 164 4
rect -4 -6 164 -4
<< m2contact >>
rect 38 84 46 92
rect 52 84 60 92
rect 38 46 46 54
rect 46 32 54 40
<< metal2 >>
rect 38 54 44 84
rect 54 32 60 84
<< m1p >>
rect 52 106 60 114
rect 132 106 140 114
rect 20 86 28 94
rect 4 66 12 74
<< labels >>
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 56 110 56 110 4 YC
rlabel metal1 8 70 8 70 4 A
rlabel metal1 24 90 24 90 4 B
rlabel metal1 136 110 136 110 4 YS
<< end >>

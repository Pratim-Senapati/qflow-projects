magic
tech scmos
magscale 1 2
timestamp 1742223327
<< metal1 >>
rect 520 606 526 614
rect 534 606 540 614
rect 548 606 554 614
rect 562 606 568 614
rect 509 543 515 563
rect 573 557 648 563
rect 477 537 515 543
rect 29 517 76 523
rect 541 517 563 523
rect 684 517 707 523
rect 684 512 692 517
rect 676 497 691 503
rect 628 437 643 443
rect 152 406 158 414
rect 166 406 172 414
rect 180 406 186 414
rect 194 406 200 414
rect 100 357 115 363
rect 13 337 35 343
rect 45 297 92 303
rect 430 297 460 303
rect 717 297 732 303
rect 717 277 723 297
rect 797 262 819 263
rect 804 257 819 262
rect 660 236 664 244
rect 520 206 526 214
rect 534 206 540 214
rect 548 206 554 214
rect 562 206 568 214
rect 765 177 780 183
rect 429 157 460 163
rect 356 137 419 143
rect 152 6 158 14
rect 166 6 172 14
rect 180 6 186 14
rect 194 6 200 14
<< m2contact >>
rect 526 606 534 614
rect 540 606 548 614
rect 554 606 562 614
rect 732 576 740 584
rect 252 556 260 564
rect 492 556 500 564
rect 12 536 20 544
rect 220 536 228 544
rect 460 536 468 544
rect 524 536 532 544
rect 780 536 788 544
rect 76 516 84 524
rect 124 516 132 524
rect 444 516 452 524
rect 668 516 676 524
rect 748 516 756 524
rect 796 516 804 524
rect 124 496 132 504
rect 668 496 676 504
rect 412 476 420 484
rect 652 476 660 484
rect 828 476 836 484
rect 124 436 132 444
rect 620 436 628 444
rect 158 406 166 414
rect 172 406 180 414
rect 186 406 194 414
rect 140 376 148 384
rect 92 356 100 364
rect 140 316 148 324
rect 92 296 100 304
rect 140 296 148 304
rect 460 296 468 304
rect 236 276 244 284
rect 460 276 468 284
rect 556 276 564 284
rect 620 276 628 284
rect 732 296 740 304
rect 780 296 788 304
rect 764 276 772 284
rect 268 256 276 264
rect 796 254 804 262
rect 508 236 516 244
rect 652 236 660 244
rect 526 206 534 214
rect 540 206 548 214
rect 554 206 562 214
rect 332 176 340 184
rect 780 176 788 184
rect 812 176 820 184
rect 172 156 180 164
rect 460 156 468 164
rect 652 156 660 164
rect 140 136 148 144
rect 348 136 356 144
rect 620 136 628 144
rect 76 116 84 124
rect 252 116 260 124
rect 524 116 532 124
rect 44 96 52 104
rect 524 96 532 104
rect 44 36 52 44
rect 524 36 532 44
rect 158 6 166 14
rect 172 6 180 14
rect 186 6 194 14
<< metal2 >>
rect 520 606 526 614
rect 534 606 540 614
rect 548 606 554 614
rect 562 606 568 614
rect 13 504 19 536
rect 77 304 83 516
rect 125 444 131 496
rect 253 443 259 556
rect 461 524 467 536
rect 445 504 451 516
rect 253 437 275 443
rect 152 406 158 414
rect 166 406 172 414
rect 180 406 186 414
rect 194 406 200 414
rect 93 324 99 356
rect 141 324 147 376
rect 93 304 99 316
rect 77 124 83 296
rect 173 264 179 356
rect 173 164 179 256
rect 237 244 243 276
rect 269 264 275 437
rect 445 283 451 496
rect 461 304 467 516
rect 493 484 499 556
rect 557 284 563 516
rect 797 484 803 516
rect 829 484 835 496
rect 621 284 627 436
rect 445 277 460 283
rect 269 164 275 256
rect 461 184 467 276
rect 520 206 526 214
rect 534 206 540 214
rect 548 206 554 214
rect 562 206 568 214
rect 653 184 659 236
rect 733 184 739 296
rect 765 284 771 296
rect 781 184 787 296
rect 797 262 803 316
rect 461 164 467 176
rect 621 144 627 176
rect 45 44 51 96
rect 525 44 531 96
rect 152 6 158 14
rect 166 6 172 14
rect 180 6 186 14
rect 194 6 200 14
<< m3contact >>
rect 526 606 534 614
rect 540 606 548 614
rect 554 606 562 614
rect 732 576 740 584
rect 220 536 228 544
rect 76 516 84 524
rect 124 516 132 524
rect 12 496 20 504
rect 460 516 468 524
rect 444 496 452 504
rect 412 476 420 484
rect 158 406 166 414
rect 172 406 180 414
rect 186 406 194 414
rect 172 356 180 364
rect 92 316 100 324
rect 76 296 84 304
rect 140 296 148 304
rect 172 256 180 264
rect 524 536 532 544
rect 780 536 788 544
rect 556 516 564 524
rect 668 516 676 524
rect 748 516 756 524
rect 492 476 500 484
rect 668 496 676 504
rect 828 496 836 504
rect 652 476 660 484
rect 796 476 804 484
rect 796 316 804 324
rect 764 296 772 304
rect 268 256 276 264
rect 236 236 244 244
rect 508 236 516 244
rect 526 206 534 214
rect 540 206 548 214
rect 554 206 562 214
rect 332 176 340 184
rect 460 176 468 184
rect 620 176 628 184
rect 652 176 660 184
rect 732 176 740 184
rect 812 176 820 184
rect 268 156 276 164
rect 652 156 660 164
rect 140 136 148 144
rect 348 136 356 144
rect 252 116 260 124
rect 524 116 532 124
rect 158 6 166 14
rect 172 6 180 14
rect 186 6 194 14
<< metal3 >>
rect 520 614 568 616
rect 520 606 524 614
rect 534 606 540 614
rect 548 606 554 614
rect 564 606 568 614
rect 520 604 568 606
rect 740 577 867 583
rect 228 537 524 543
rect 788 537 867 543
rect 84 517 124 523
rect 468 517 556 523
rect 564 517 668 523
rect 676 517 748 523
rect -19 497 12 503
rect 452 497 668 503
rect 836 497 867 503
rect 420 477 492 483
rect 500 477 652 483
rect 660 477 796 483
rect 152 414 200 416
rect 152 406 156 414
rect 166 406 172 414
rect 180 406 186 414
rect 196 406 200 414
rect 152 404 200 406
rect -19 357 172 363
rect -19 317 92 323
rect 804 317 867 323
rect 84 297 140 303
rect 772 297 867 303
rect 180 257 268 263
rect 244 237 508 243
rect 520 214 568 216
rect 520 206 524 214
rect 534 206 540 214
rect 548 206 554 214
rect 564 206 568 214
rect 520 204 568 206
rect 340 177 460 183
rect 628 177 652 183
rect 740 177 812 183
rect 276 157 652 163
rect 148 137 348 143
rect 260 117 524 123
rect 152 14 200 16
rect 152 6 156 14
rect 166 6 172 14
rect 180 6 186 14
rect 196 6 200 14
rect 152 4 200 6
<< m4contact >>
rect 524 606 526 614
rect 526 606 532 614
rect 540 606 548 614
rect 556 606 562 614
rect 562 606 564 614
rect 156 406 158 414
rect 158 406 164 414
rect 172 406 180 414
rect 188 406 194 414
rect 194 406 196 414
rect 524 206 526 214
rect 526 206 532 214
rect 540 206 548 214
rect 556 206 562 214
rect 562 206 564 214
rect 156 6 158 14
rect 158 6 164 14
rect 172 6 180 14
rect 188 6 194 14
rect 194 6 196 14
<< metal4 >>
rect 152 414 200 620
rect 152 406 156 414
rect 164 406 172 414
rect 180 406 188 414
rect 196 406 200 414
rect 152 14 200 406
rect 152 6 156 14
rect 164 6 172 14
rect 180 6 188 14
rect 196 6 200 14
rect 152 0 200 6
rect 520 614 568 620
rect 520 606 524 614
rect 532 606 540 614
rect 548 606 556 614
rect 564 606 568 614
rect 520 214 568 606
rect 520 206 524 214
rect 532 206 540 214
rect 548 206 556 214
rect 564 206 568 214
rect 520 0 568 206
use DFFSR  DFFSR_1
timestamp 1742223327
transform 1 0 8 0 -1 210
box -4 -6 356 206
use FILL  FILL_0_0_0
timestamp 1742223327
transform -1 0 376 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_6
timestamp 1742223327
transform -1 0 56 0 1 210
box -4 -6 52 206
use FILL  FILL_1_0_0
timestamp 1742223327
transform 1 0 56 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1742223327
transform 1 0 72 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_2
timestamp 1742223327
transform 1 0 88 0 1 210
box -4 -6 20 206
use DFFSR  DFFSR_2
timestamp 1742223327
transform 1 0 104 0 1 210
box -4 -6 356 206
use XOR2X1  XOR2X1_1
timestamp 1742223327
transform 1 0 456 0 1 210
box -4 -6 116 206
use FILL  FILL_0_1_2
timestamp 1742223327
transform 1 0 472 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1742223327
transform 1 0 456 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_0
timestamp 1742223327
transform 1 0 440 0 -1 210
box -4 -6 20 206
use INVX1  INVX1_1
timestamp 1742223327
transform -1 0 440 0 -1 210
box -4 -6 36 206
use FILL  FILL_0_0_2
timestamp 1742223327
transform -1 0 408 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1742223327
transform -1 0 392 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_4
timestamp 1742223327
transform 1 0 728 0 1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_1
timestamp 1742223327
transform 1 0 616 0 1 210
box -4 -6 116 206
use FILL  FILL_1_1_2
timestamp 1742223327
transform 1 0 600 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_1
timestamp 1742223327
transform 1 0 584 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_0
timestamp 1742223327
transform 1 0 568 0 1 210
box -4 -6 20 206
use DFFSR  DFFSR_4
timestamp 1742223327
transform 1 0 488 0 -1 210
box -4 -6 356 206
use BUFX2  BUFX2_5
timestamp 1742223327
transform 1 0 776 0 1 210
box -4 -6 52 206
use FILL  FILL_2_1
timestamp 1742223327
transform 1 0 824 0 1 210
box -4 -6 20 206
use INVX2  INVX2_1
timestamp 1742223327
transform 1 0 8 0 -1 610
box -4 -6 36 206
use FILL  FILL_2_0_0
timestamp 1742223327
transform 1 0 40 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1742223327
transform 1 0 56 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1742223327
transform 1 0 72 0 -1 610
box -4 -6 20 206
use DFFSR  DFFSR_3
timestamp 1742223327
transform 1 0 88 0 -1 610
box -4 -6 356 206
use AOI21X1  AOI21X1_1
timestamp 1742223327
transform 1 0 440 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_1
timestamp 1742223327
transform 1 0 504 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_2
timestamp 1742223327
transform -1 0 584 0 -1 610
box -4 -6 36 206
use FILL  FILL_2_1_0
timestamp 1742223327
transform -1 0 600 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1742223327
transform -1 0 616 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1742223327
transform -1 0 632 0 -1 610
box -4 -6 20 206
use NAND3X1  NAND3X1_1
timestamp 1742223327
transform -1 0 696 0 -1 610
box -4 -6 68 206
use BUFX2  BUFX2_1
timestamp 1742223327
transform 1 0 696 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_2
timestamp 1742223327
transform 1 0 744 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_3
timestamp 1742223327
transform 1 0 792 0 -1 610
box -4 -6 52 206
<< labels >>
flabel metal3 s -16 320 -16 320 7 FreeSans 24 0 0 0 vdd
port 0 nsew
flabel metal3 s 864 320 864 320 3 FreeSans 24 0 0 0 gnd
port 1 nsew
flabel metal3 s -19 357 -13 363 7 FreeSans 24 0 0 0 clk
port 2 nsew
flabel metal3 s -19 497 -13 503 7 FreeSans 24 0 0 0 rst
port 3 nsew
flabel metal3 s 861 577 867 583 3 FreeSans 24 90 0 0 count[0]
port 4 nsew
flabel metal3 s 861 537 867 543 3 FreeSans 24 0 0 0 count[1]
port 5 nsew
flabel metal3 s 861 497 867 503 3 FreeSans 24 0 0 0 count[2]
port 6 nsew
flabel metal3 s 861 297 867 303 3 FreeSans 24 0 0 0 count[3]
port 7 nsew
<< end >>

magic
tech scmos
timestamp 1740169866
<< metal1 >>
rect 30 1497 420 1500
rect 3 1010 447 1497
rect 0 521 450 1010
rect 3 489 447 521
rect 0 9 450 489
rect 0 0 171 9
rect 174 0 274 4
rect 278 0 450 9
<< metal2 >>
rect 30 1497 420 1500
rect 3 1010 447 1497
rect 0 648 450 1010
rect 3 626 447 648
rect 0 521 450 626
rect 3 489 447 521
rect 0 384 450 489
rect 3 383 448 384
rect 3 362 447 383
rect 0 0 450 362
<< metal3 >>
rect 3 3 447 1497
<< metal4 >>
rect 3 1495 178 1497
rect 265 1495 447 1497
rect 3 1358 447 1495
rect 3 1265 178 1358
rect 187 1274 256 1349
rect 265 1265 447 1358
rect 3 3 447 1265
<< labels >>
rlabel metal4 s 187 1274 256 1349 6 YPAD
port 1 nsew default output
rlabel metal1 s 174 0 274 4 6 gnd
port 2 nsew ground bidirectional
<< properties >>
string LEFsite IO
string LEFclass PAD
string FIXED_BBOX 0 0 450 1500
string LEFsymmetry R90
string LEFview TRUE
<< end >>

magic
tech scmos
magscale 1 2
timestamp 1740717622
<< nwell >>
rect -10 96 252 210
rect 46 92 200 96
rect 130 78 200 92
<< ntransistor >>
rect 14 12 18 52
rect 30 12 34 52
rect 46 12 50 52
rect 62 12 66 52
rect 72 12 76 52
rect 88 12 92 52
rect 104 12 108 52
rect 120 12 124 52
rect 136 12 140 52
rect 154 12 158 52
rect 164 12 168 52
rect 174 12 178 52
rect 190 12 194 32
rect 222 12 226 32
<< ptransistor >>
rect 14 108 18 188
rect 30 108 34 188
rect 46 108 50 188
rect 62 108 66 188
rect 72 108 76 188
rect 88 108 92 188
rect 104 116 108 188
rect 120 116 124 188
rect 136 116 140 188
rect 154 92 158 188
rect 164 92 168 188
rect 174 92 178 188
rect 190 148 194 188
rect 222 148 226 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 40 30 52
rect 18 12 20 40
rect 28 12 30 40
rect 34 51 46 52
rect 34 13 36 51
rect 44 13 46 51
rect 34 12 46 13
rect 50 42 62 52
rect 50 14 52 42
rect 60 14 62 42
rect 50 12 62 14
rect 66 12 72 52
rect 76 44 88 52
rect 76 16 78 44
rect 86 16 88 44
rect 76 12 88 16
rect 92 50 104 52
rect 92 12 94 50
rect 102 12 104 50
rect 108 34 120 52
rect 108 16 110 34
rect 118 16 120 34
rect 108 12 120 16
rect 124 50 136 52
rect 124 12 126 50
rect 134 12 136 50
rect 140 41 154 52
rect 140 13 143 41
rect 151 13 154 41
rect 140 12 154 13
rect 158 12 164 52
rect 168 12 174 52
rect 178 50 188 52
rect 178 12 180 50
rect 188 12 190 32
rect 194 31 204 32
rect 194 13 196 31
rect 194 12 204 13
rect 212 31 222 32
rect 220 13 222 31
rect 212 12 222 13
rect 226 31 236 32
rect 226 13 228 31
rect 226 12 236 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 109 14 187
rect 4 108 14 109
rect 18 120 20 188
rect 28 120 30 188
rect 18 108 30 120
rect 34 187 46 188
rect 34 109 36 187
rect 44 109 46 187
rect 34 108 46 109
rect 50 186 62 188
rect 50 118 52 186
rect 60 118 62 186
rect 50 108 62 118
rect 66 108 72 188
rect 76 187 88 188
rect 76 109 78 187
rect 86 109 88 187
rect 76 108 88 109
rect 92 187 104 188
rect 92 109 94 187
rect 102 116 104 187
rect 108 187 120 188
rect 108 129 110 187
rect 118 129 120 187
rect 108 116 120 129
rect 124 186 136 188
rect 124 118 126 186
rect 134 118 136 186
rect 124 116 136 118
rect 140 184 154 188
rect 140 116 143 184
rect 92 108 102 109
rect 142 106 143 116
rect 151 106 154 184
rect 142 102 154 106
rect 144 94 154 102
rect 148 92 154 94
rect 158 92 164 188
rect 168 92 174 188
rect 178 184 190 188
rect 178 96 180 184
rect 188 148 190 184
rect 194 187 204 188
rect 194 149 196 187
rect 194 148 204 149
rect 212 187 222 188
rect 220 149 222 187
rect 212 148 222 149
rect 226 187 236 188
rect 226 149 228 187
rect 226 148 236 149
rect 178 92 188 96
<< ndcontact >>
rect 4 13 12 51
rect 20 12 28 40
rect 36 13 44 51
rect 52 14 60 42
rect 78 16 86 44
rect 94 12 102 50
rect 110 16 118 34
rect 126 12 134 50
rect 143 13 151 41
rect 180 12 188 50
rect 196 13 204 31
rect 212 13 220 31
rect 228 13 236 31
<< pdcontact >>
rect 4 109 12 187
rect 20 120 28 188
rect 36 109 44 187
rect 52 118 60 186
rect 78 109 86 187
rect 94 109 102 187
rect 110 129 118 187
rect 126 118 134 186
rect 143 106 151 184
rect 180 96 188 184
rect 196 149 204 187
rect 212 149 220 187
rect 228 149 236 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
rect 92 -4 100 4
rect 124 -4 132 4
rect 156 -4 164 4
rect 188 -4 196 4
rect 220 -4 228 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
rect 92 196 100 204
rect 124 196 132 204
rect 156 196 164 204
rect 188 196 196 204
rect 220 196 228 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 46 188 50 192
rect 62 188 66 192
rect 72 188 76 192
rect 88 188 92 192
rect 104 188 108 192
rect 120 188 124 192
rect 136 188 140 192
rect 154 188 158 192
rect 164 188 168 192
rect 174 188 178 192
rect 190 188 194 192
rect 222 188 226 192
rect 14 66 18 108
rect 30 78 34 108
rect 46 94 50 108
rect 14 52 18 58
rect 30 52 34 70
rect 46 52 50 86
rect 62 78 66 108
rect 72 106 76 108
rect 88 106 92 108
rect 104 106 108 116
rect 120 114 124 116
rect 136 114 140 116
rect 72 102 92 106
rect 98 102 108 106
rect 114 110 124 114
rect 132 110 140 114
rect 62 52 66 70
rect 74 64 78 102
rect 98 76 102 102
rect 114 90 118 110
rect 132 102 136 110
rect 102 68 108 72
rect 72 56 74 58
rect 82 56 92 58
rect 72 54 92 56
rect 72 52 76 54
rect 88 52 92 54
rect 104 52 108 68
rect 114 58 118 82
rect 132 58 136 94
rect 190 146 194 148
rect 190 142 198 146
rect 154 88 158 92
rect 152 84 158 88
rect 148 58 152 80
rect 164 76 168 92
rect 174 88 178 92
rect 174 84 182 88
rect 114 54 124 58
rect 132 54 140 58
rect 148 54 158 58
rect 120 52 124 54
rect 136 52 140 54
rect 154 52 158 54
rect 164 52 168 68
rect 178 76 182 84
rect 194 78 198 142
rect 222 114 226 148
rect 224 106 226 114
rect 178 60 182 68
rect 174 56 182 60
rect 174 52 178 56
rect 194 50 198 70
rect 190 46 198 50
rect 190 32 194 46
rect 222 32 226 106
rect 14 8 18 12
rect 30 8 34 12
rect 46 8 50 12
rect 62 8 66 12
rect 72 8 76 12
rect 88 8 92 12
rect 104 8 108 12
rect 120 8 124 12
rect 136 8 140 12
rect 154 8 158 12
rect 164 8 168 12
rect 174 8 178 12
rect 190 8 194 12
rect 222 8 226 12
<< polycontact >>
rect 44 86 52 94
rect 28 70 36 78
rect 12 58 20 66
rect 58 70 66 78
rect 128 94 136 102
rect 110 82 118 90
rect 94 68 102 76
rect 74 56 82 64
rect 144 80 152 88
rect 160 68 168 76
rect 216 106 224 114
rect 178 68 186 76
rect 194 70 202 78
<< metal1 >>
rect -4 204 244 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 92 204
rect 100 196 124 204
rect 132 196 156 204
rect 164 196 188 204
rect 196 196 220 204
rect 228 196 244 204
rect -4 194 244 196
rect 20 188 28 194
rect 4 187 12 188
rect 36 187 44 188
rect 12 109 36 114
rect 4 108 44 109
rect 52 186 60 188
rect 52 116 60 118
rect 78 187 86 194
rect 78 108 86 109
rect 94 187 102 188
rect 110 187 118 194
rect 110 128 118 129
rect 126 186 134 188
rect 102 118 126 122
rect 102 116 134 118
rect 142 184 152 188
rect 94 108 102 109
rect 142 106 143 184
rect 151 106 152 184
rect 142 102 152 106
rect 180 184 188 194
rect 196 187 204 188
rect 20 86 28 94
rect 36 86 44 94
rect 180 92 188 96
rect 194 149 196 154
rect 194 148 204 149
rect 212 187 220 194
rect 212 148 220 149
rect 228 187 236 188
rect 228 148 236 149
rect 194 98 200 148
rect 194 92 214 98
rect 52 86 110 92
rect 4 66 12 74
rect 22 72 28 86
rect 104 82 110 86
rect 118 82 144 88
rect 36 70 58 76
rect 66 70 94 76
rect 102 68 160 74
rect 6 60 12 66
rect 20 58 74 64
rect 178 62 184 68
rect 82 56 184 62
rect 208 54 214 92
rect 230 74 236 148
rect 228 66 236 74
rect 4 51 44 52
rect 12 46 36 51
rect 4 12 12 13
rect 36 12 44 13
rect 52 42 60 44
rect 52 12 60 14
rect 78 44 86 48
rect 20 6 28 12
rect 78 6 86 16
rect 102 44 126 50
rect 110 34 118 38
rect 110 6 118 16
rect 142 41 152 42
rect 142 13 143 41
rect 151 13 152 41
rect 142 12 152 13
rect 208 46 220 54
rect 208 44 214 46
rect 198 38 214 44
rect 198 32 204 38
rect 230 32 236 66
rect 196 31 204 32
rect 196 12 204 13
rect 212 31 220 32
rect 180 6 188 12
rect 212 6 220 13
rect 228 31 236 32
rect 228 12 236 13
rect -4 4 244 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 92 4
rect 100 -4 124 4
rect 132 -4 156 4
rect 164 -4 188 4
rect 196 -4 220 4
rect 228 -4 244 4
rect -4 -6 244 -4
<< m2contact >>
rect 52 108 60 116
rect 120 96 128 104
rect 144 94 152 102
rect 208 106 216 114
rect 194 78 202 86
rect 52 44 60 52
rect 144 42 152 50
<< metal2 >>
rect 60 108 208 114
rect 54 52 60 108
rect 120 104 128 108
rect 146 84 152 94
rect 146 78 194 84
rect 146 50 152 78
<< m1p >>
rect 20 86 28 94
rect 36 86 44 94
rect 4 66 12 74
rect 228 66 236 74
rect 212 46 220 54
<< labels >>
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 70 8 70 4 A
rlabel metal1 24 90 24 90 4 B
rlabel metal1 40 90 40 90 4 C
rlabel metal1 232 70 232 70 4 YC
rlabel metal1 216 50 216 50 4 YS
<< end >>

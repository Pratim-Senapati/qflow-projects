magic
tech scmos
magscale 1 2
timestamp 1740382396
<< nwell >>
rect -16 96 288 210
<< ntransistor >>
rect 14 12 18 52
rect 30 12 34 52
rect 46 12 50 52
rect 62 12 66 52
rect 78 12 82 52
rect 94 12 98 52
rect 110 12 114 52
rect 126 12 130 52
rect 142 12 146 52
rect 158 12 162 52
rect 174 12 178 52
rect 190 12 194 52
rect 206 12 210 52
rect 222 12 226 52
rect 238 12 242 52
rect 254 12 258 52
<< ptransistor >>
rect 14 108 18 188
rect 30 108 34 188
rect 46 108 50 188
rect 62 108 66 188
rect 78 108 82 188
rect 94 108 98 188
rect 110 108 114 188
rect 126 108 130 188
rect 142 108 146 188
rect 158 108 162 188
rect 174 108 178 188
rect 190 108 194 188
rect 206 108 210 188
rect 222 108 226 188
rect 238 108 242 188
rect 254 108 258 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 51 30 52
rect 18 13 20 51
rect 28 13 30 51
rect 18 12 30 13
rect 34 51 46 52
rect 34 13 36 51
rect 44 13 46 51
rect 34 12 46 13
rect 50 51 62 52
rect 50 13 52 51
rect 60 13 62 51
rect 50 12 62 13
rect 66 51 78 52
rect 66 13 68 51
rect 76 13 78 51
rect 66 12 78 13
rect 82 51 94 52
rect 82 13 84 51
rect 92 13 94 51
rect 82 12 94 13
rect 98 51 110 52
rect 98 13 100 51
rect 108 13 110 51
rect 98 12 110 13
rect 114 51 126 52
rect 114 13 116 51
rect 124 13 126 51
rect 114 12 126 13
rect 130 51 142 52
rect 130 13 132 51
rect 140 13 142 51
rect 130 12 142 13
rect 146 51 158 52
rect 146 13 148 51
rect 156 13 158 51
rect 146 12 158 13
rect 162 51 174 52
rect 162 13 164 51
rect 172 13 174 51
rect 162 12 174 13
rect 178 51 190 52
rect 178 13 180 51
rect 188 13 190 51
rect 178 12 190 13
rect 194 51 206 52
rect 194 13 196 51
rect 204 13 206 51
rect 194 12 206 13
rect 210 51 222 52
rect 210 13 212 51
rect 220 13 222 51
rect 210 12 222 13
rect 226 51 238 52
rect 226 13 228 51
rect 236 13 238 51
rect 226 12 238 13
rect 242 51 254 52
rect 242 13 244 51
rect 252 13 254 51
rect 242 12 254 13
rect 258 51 268 52
rect 258 13 260 51
rect 258 12 268 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 109 14 187
rect 4 108 14 109
rect 18 187 30 188
rect 18 109 20 187
rect 28 109 30 187
rect 18 108 30 109
rect 34 187 46 188
rect 34 109 36 187
rect 44 109 46 187
rect 34 108 46 109
rect 50 187 62 188
rect 50 109 52 187
rect 60 109 62 187
rect 50 108 62 109
rect 66 187 78 188
rect 66 109 68 187
rect 76 109 78 187
rect 66 108 78 109
rect 82 187 94 188
rect 82 109 84 187
rect 92 109 94 187
rect 82 108 94 109
rect 98 187 110 188
rect 98 109 100 187
rect 108 109 110 187
rect 98 108 110 109
rect 114 187 126 188
rect 114 109 116 187
rect 124 109 126 187
rect 114 108 126 109
rect 130 187 142 188
rect 130 109 132 187
rect 140 109 142 187
rect 130 108 142 109
rect 146 187 158 188
rect 146 109 148 187
rect 156 109 158 187
rect 146 108 158 109
rect 162 187 174 188
rect 162 109 164 187
rect 172 109 174 187
rect 162 108 174 109
rect 178 187 190 188
rect 178 109 180 187
rect 188 109 190 187
rect 178 108 190 109
rect 194 187 206 188
rect 194 109 196 187
rect 204 109 206 187
rect 194 108 206 109
rect 210 187 222 188
rect 210 109 212 187
rect 220 109 222 187
rect 210 108 222 109
rect 226 187 238 188
rect 226 109 228 187
rect 236 109 238 187
rect 226 108 238 109
rect 242 187 254 188
rect 242 109 244 187
rect 252 109 254 187
rect 242 108 254 109
rect 258 187 268 188
rect 258 109 260 187
rect 258 108 268 109
<< ndcontact >>
rect 4 13 12 51
rect 20 13 28 51
rect 36 13 44 51
rect 52 13 60 51
rect 68 13 76 51
rect 84 13 92 51
rect 100 13 108 51
rect 116 13 124 51
rect 132 13 140 51
rect 148 13 156 51
rect 164 13 172 51
rect 180 13 188 51
rect 196 13 204 51
rect 212 13 220 51
rect 228 13 236 51
rect 244 13 252 51
rect 260 13 268 51
<< pdcontact >>
rect 4 109 12 187
rect 20 109 28 187
rect 36 109 44 187
rect 52 109 60 187
rect 68 109 76 187
rect 84 109 92 187
rect 100 109 108 187
rect 116 109 124 187
rect 132 109 140 187
rect 148 109 156 187
rect 164 109 172 187
rect 180 109 188 187
rect 196 109 204 187
rect 212 109 220 187
rect 228 109 236 187
rect 244 109 252 187
rect 260 109 268 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
rect 92 -4 100 4
rect 124 -4 132 4
rect 156 -4 164 4
rect 188 -4 196 4
rect 220 -4 228 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
rect 92 196 100 204
rect 124 196 132 204
rect 156 196 164 204
rect 188 196 196 204
rect 220 196 228 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 46 188 50 192
rect 62 188 66 192
rect 78 188 82 192
rect 94 188 98 192
rect 110 188 114 192
rect 126 188 130 192
rect 142 188 146 192
rect 158 188 162 192
rect 174 188 178 192
rect 190 188 194 192
rect 206 188 210 192
rect 222 188 226 192
rect 238 188 242 192
rect 254 188 258 192
rect 14 80 18 108
rect 30 80 34 108
rect 22 72 34 80
rect 14 52 18 72
rect 30 52 34 72
rect 46 80 50 108
rect 62 80 66 108
rect 46 72 48 80
rect 56 72 66 80
rect 46 52 50 72
rect 62 52 66 72
rect 78 52 82 108
rect 94 80 98 108
rect 110 80 114 108
rect 126 80 130 108
rect 90 72 98 80
rect 108 72 116 80
rect 124 72 130 80
rect 94 52 98 72
rect 110 52 114 72
rect 126 52 130 72
rect 142 80 146 108
rect 158 80 162 108
rect 150 72 162 80
rect 142 52 146 72
rect 158 52 162 72
rect 174 80 178 108
rect 190 80 194 108
rect 174 72 176 80
rect 184 72 194 80
rect 174 52 178 72
rect 190 52 194 72
rect 206 52 210 108
rect 222 80 226 108
rect 238 80 242 108
rect 254 80 258 108
rect 218 72 226 80
rect 236 72 244 80
rect 252 72 258 80
rect 222 52 226 72
rect 238 52 242 72
rect 254 52 258 72
rect 14 8 18 12
rect 30 8 34 12
rect 46 8 50 12
rect 62 8 66 12
rect 78 8 82 12
rect 94 8 98 12
rect 110 8 114 12
rect 126 8 130 12
rect 142 8 146 12
rect 158 8 162 12
rect 174 8 178 12
rect 190 8 194 12
rect 206 8 210 12
rect 222 8 226 12
rect 238 8 242 12
rect 254 8 258 12
<< polycontact >>
rect 14 72 22 80
rect 48 72 56 80
rect 82 72 90 80
rect 116 72 124 80
rect 142 72 150 80
rect 176 72 184 80
rect 210 72 218 80
rect 244 72 252 80
<< metal1 >>
rect -4 204 276 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 92 204
rect 100 196 124 204
rect 132 196 156 204
rect 164 196 188 204
rect 196 196 220 204
rect 228 196 276 204
rect -4 194 276 196
rect 4 187 12 194
rect 4 108 12 109
rect 20 187 28 188
rect 20 102 28 109
rect 36 187 44 194
rect 36 108 44 109
rect 52 187 60 188
rect 52 102 60 109
rect 68 187 76 194
rect 68 108 76 109
rect 84 187 92 188
rect 84 102 92 109
rect 100 187 108 194
rect 100 108 108 109
rect 116 187 124 188
rect 116 102 124 109
rect 132 187 140 194
rect 132 108 140 109
rect 148 187 156 188
rect 148 102 156 109
rect 164 187 172 194
rect 164 108 172 109
rect 180 187 188 188
rect 180 102 188 109
rect 196 187 204 194
rect 196 108 204 109
rect 212 187 220 188
rect 212 102 220 109
rect 228 187 236 194
rect 228 108 236 109
rect 244 187 252 188
rect 244 102 252 109
rect 260 187 268 194
rect 260 108 268 109
rect 20 94 38 102
rect 52 94 74 102
rect 84 94 106 102
rect 116 94 140 102
rect 148 94 166 102
rect 180 94 202 102
rect 212 94 234 102
rect 244 94 268 102
rect 30 80 38 94
rect 66 80 74 94
rect 98 80 106 94
rect 132 80 140 94
rect 158 80 166 94
rect 194 80 202 94
rect 226 80 234 94
rect 4 72 14 80
rect 30 72 48 80
rect 66 72 82 80
rect 98 72 116 80
rect 132 72 142 80
rect 158 72 176 80
rect 194 72 210 80
rect 226 72 244 80
rect 4 66 12 72
rect 30 66 38 72
rect 66 66 74 72
rect 98 66 106 72
rect 132 66 140 72
rect 158 66 166 72
rect 194 66 202 72
rect 226 66 234 72
rect 260 66 268 94
rect 20 58 38 66
rect 52 58 74 66
rect 84 58 106 66
rect 116 58 140 66
rect 148 58 166 66
rect 180 58 202 66
rect 212 58 234 66
rect 244 58 268 66
rect 4 51 12 52
rect 4 6 12 13
rect 20 51 28 58
rect 20 12 28 13
rect 36 51 44 52
rect 36 6 44 13
rect 52 51 60 58
rect 52 12 60 13
rect 68 51 76 52
rect 68 6 76 13
rect 84 51 92 58
rect 84 12 92 13
rect 100 51 108 52
rect 100 6 108 13
rect 116 51 124 58
rect 116 12 124 13
rect 132 51 140 52
rect 132 6 140 13
rect 148 51 156 58
rect 148 12 156 13
rect 164 51 172 52
rect 164 6 172 13
rect 180 51 188 58
rect 180 12 188 13
rect 196 51 204 52
rect 196 6 204 13
rect 212 51 220 58
rect 212 12 220 13
rect 228 51 236 52
rect 228 6 236 13
rect 244 51 252 58
rect 244 12 252 13
rect 260 51 268 52
rect 260 6 268 13
rect -4 4 276 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 92 4
rect 100 -4 124 4
rect 132 -4 156 4
rect 164 -4 188 4
rect 196 -4 220 4
rect 228 -4 276 4
rect -4 -6 276 -4
<< m1p >>
rect 260 86 268 94
rect 4 66 12 74
<< labels >>
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 70 8 70 4 A
rlabel metal1 264 90 264 90 4 Y
<< end >>

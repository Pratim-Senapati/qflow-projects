* NGSPICE file created from map9v3.ext - technology: scmos

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

.subckt map9v3 vdd gnd clock reset start N[0] N[1] N[2] N[3] N[4] N[5] N[6] N[7] N[8]
+ dp[0] dp[1] dp[2] dp[3] dp[4] dp[5] dp[6] dp[7] dp[8] done counter[0] counter[1]
+ counter[2] counter[3] counter[4] counter[5] counter[6] counter[7] sr[0] sr[1] sr[2]
+ sr[3] sr[4] sr[5] sr[6] sr[7]
XDFFSR_9 BUFX2_2/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_9/D gnd vdd DFFSR
XOAI21X1_19 BUFX2_3/A INVX1_24/A BUFX2_4/A gnd AND2X2_2/A vdd OAI21X1
XFILL_3_2_0 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XAOI22X1_1 INVX4_1/A AOI22X1_1/B AOI22X1_1/C AOI22X1_1/D gnd DFFSR_13/D vdd AOI22X1
XFILL_10_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XAOI22X1_2 INVX8_1/A AOI22X1_2/B BUFX2_7/A AOI22X1_2/D gnd AOI22X1_2/Y vdd AOI22X1
XFILL_10_2 gnd vdd FILL
XINVX8_1 INVX8_1/A gnd BUFX4_4/A vdd INVX8
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_1_3_0 gnd vdd FILL
XFILL_6_2_0 gnd vdd FILL
XNOR3X1_1 BUFX2_6/A BUFX2_5/A BUFX2_7/A gnd NOR3X1_1/Y vdd NOR3X1
XFILL_10_3 gnd vdd FILL
XINVX8_2 reset gnd BUFX4_5/A vdd INVX8
XFILL_3_0_0 gnd vdd FILL
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XCLKBUF1_1 clock gnd DFFSR_5/CLK vdd CLKBUF1
XCLKBUF1_2 clock gnd CLKBUF1_2/Y vdd CLKBUF1
XMUX2X1_1 INVX1_5/Y INVX1_6/Y MUX2X1_2/S gnd DFFSR_26/D vdd MUX2X1
XFILL_4_3_0 gnd vdd FILL
XFILL_9_2_0 gnd vdd FILL
XFILL_7_1 gnd vdd FILL
XNAND3X1_1 NOR2X1_1/Y NOR2X1_2/Y NOR3X1_1/Y gnd NAND3X1_1/Y vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XXOR2X1_1 INVX1_24/A BUFX2_3/A gnd XOR2X1_1/Y vdd XOR2X1
XCLKBUF1_3 clock gnd DFFSR_9/CLK vdd CLKBUF1
XFILL_6_0_0 gnd vdd FILL
XMUX2X1_2 INVX1_7/Y INVX1_8/Y MUX2X1_2/S gnd MUX2X1_2/Y vdd MUX2X1
XFILL_7_2 gnd vdd FILL
XNAND3X1_2 DFFSR_3/Q INVX4_1/Y BUFX4_2/Y gnd MUX2X1_2/S vdd NAND3X1
XMUX2X1_3 INVX1_9/Y MUX2X1_3/B MUX2X1_2/S gnd DFFSR_28/D vdd MUX2X1
XCLKBUF1_4 clock gnd DFFSR_3/CLK vdd CLKBUF1
XFILL_7_3 gnd vdd FILL
XNAND3X1_3 DFFSR_5/Q BUFX4_2/Y INVX1_21/Y gnd NAND3X1_3/Y vdd NAND3X1
XMUX2X1_4 INVX1_11/Y INVX1_12/Y MUX2X1_2/S gnd DFFSR_29/D vdd MUX2X1
XFILL_7_3_0 gnd vdd FILL
XCLKBUF1_5 clock gnd DFFSR_8/CLK vdd CLKBUF1
XBUFX4_1 BUFX4_4/A gnd BUFX4_1/Y vdd BUFX4
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XFILL_4_1_0 gnd vdd FILL
XFILL_9_0_0 gnd vdd FILL
XNAND3X1_4 INVX4_1/A NAND2X1_5/Y NAND3X1_4/C gnd NAND3X1_4/Y vdd NAND3X1
XOAI21X1_1 BUFX2_8/A NAND3X1_1/Y INVX8_1/A gnd OAI21X1_1/Y vdd OAI21X1
XMUX2X1_5 INVX1_13/Y INVX1_14/Y MUX2X1_2/S gnd DFFSR_30/D vdd MUX2X1
XBUFX4_2 BUFX4_4/A gnd BUFX4_2/Y vdd BUFX4
XNAND3X1_5 INVX8_1/A NOR2X1_1/Y NOR2X1_2/Y gnd AND2X2_2/B vdd NAND3X1
XOAI21X1_2 INVX1_1/Y NOR2X1_3/Y INVX1_2/Y gnd DFFSR_2/D vdd OAI21X1
XMUX2X1_6 MUX2X1_6/A MUX2X1_6/B MUX2X1_2/S gnd MUX2X1_6/Y vdd MUX2X1
XBUFX4_3 BUFX4_4/A gnd BUFX4_3/Y vdd BUFX4
XNAND3X1_6 INVX2_1/A NOR2X1_10/Y NOR2X1_13/Y gnd INVX1_30/A vdd NAND3X1
XMUX2X1_7 MUX2X1_7/A MUX2X1_7/B MUX2X1_2/S gnd MUX2X1_7/Y vdd MUX2X1
XOAI21X1_3 XNOR2X1_1/Y XNOR2X1_2/Y INVX8_1/A gnd OAI21X1_3/Y vdd OAI21X1
XFILL_2_2_0 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XBUFX2_1 BUFX2_1/A gnd counter[0] vdd BUFX2
XBUFX4_4 BUFX4_4/A gnd BUFX4_4/Y vdd BUFX4
XNAND3X1_7 INVX1_28/Y INVX1_26/Y INVX1_32/Y gnd NOR2X1_14/A vdd NAND3X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XOAI21X1_4 INVX8_1/A BUFX2_19/A INVX4_1/Y gnd NOR2X1_6/A vdd OAI21X1
XFILL_3_1 gnd vdd FILL
XAOI21X1_1 INVX1_4/Y MUX2X1_2/S NOR2X1_4/Y gnd DFFSR_25/D vdd AOI21X1
XBUFX4_5 BUFX4_5/A gnd DFFSR_9/R vdd BUFX4
XAOI21X1_2 INVX1_19/Y MUX2X1_2/S NOR2X1_5/Y gnd DFFSR_24/D vdd AOI21X1
XBUFX2_2 BUFX2_2/A gnd counter[1] vdd BUFX2
XNAND3X1_8 INVX1_28/Y INVX1_26/Y INVX1_27/Y gnd AOI22X1_2/D vdd NAND3X1
XBUFX2_20 INVX1_6/A gnd sr[1] vdd BUFX2
XAOI21X1_10 BUFX4_2/Y INVX1_6/Y AOI21X1_10/C gnd DFFSR_17/D vdd AOI21X1
XOAI21X1_5 INVX1_6/A BUFX4_1/Y INVX4_1/Y gnd AOI21X1_4/C vdd OAI21X1
XBUFX2_3 BUFX2_3/A gnd counter[2] vdd BUFX2
XBUFX4_6 BUFX4_5/A gnd BUFX4_6/Y vdd BUFX4
XNAND3X1_9 INVX1_29/Y N[8] INVX1_30/Y gnd NAND3X1_9/Y vdd NAND3X1
XFILL_0_3_0 gnd vdd FILL
XBUFX2_10 BUFX2_10/A gnd dp[0] vdd BUFX2
XNOR2X1_1 BUFX2_4/A BUFX2_3/A gnd NOR2X1_1/Y vdd NOR2X1
XFILL_5_2_0 gnd vdd FILL
XAOI21X1_3 XNOR2X1_1/Y XNOR2X1_2/Y OAI21X1_3/Y gnd NOR2X1_6/B vdd AOI21X1
XOAI21X1_6 INVX1_8/A BUFX4_1/Y INVX4_1/Y gnd OAI21X1_6/Y vdd OAI21X1
XBUFX2_21 INVX1_8/A gnd sr[2] vdd BUFX2
XAOI21X1_11 NAND3X1_3/Y INVX1_20/Y INVX4_1/A gnd DFFSR_33/D vdd AOI21X1
XFILL_2_0_0 gnd vdd FILL
XBUFX4_7 BUFX4_5/A gnd BUFX4_7/Y vdd BUFX4
XNOR2X1_2 BUFX2_2/A BUFX2_1/A gnd NOR2X1_2/Y vdd NOR2X1
XBUFX2_4 BUFX2_4/A gnd counter[3] vdd BUFX2
XBUFX2_22 BUFX2_22/A gnd sr[3] vdd BUFX2
XAOI21X1_4 BUFX4_1/Y INVX1_8/Y AOI21X1_4/C gnd DFFSR_18/D vdd AOI21X1
XBUFX2_11 INVX1_4/A gnd dp[1] vdd BUFX2
XAOI21X1_12 INVX2_1/Y N[3] INVX4_1/Y gnd OAI21X1_16/C vdd AOI21X1
XOAI21X1_7 BUFX2_22/A BUFX4_2/Y INVX4_1/Y gnd OAI21X1_7/Y vdd OAI21X1
XFILL_1_1 gnd vdd FILL
XBUFX4_8 BUFX4_5/A gnd DFFSR_3/R vdd BUFX4
XAOI21X1_13 NOR2X1_10/Y INVX2_1/A INVX1_25/Y gnd OAI21X1_23/A vdd AOI21X1
XBUFX2_5 BUFX2_5/A gnd counter[4] vdd BUFX2
XBUFX2_23 BUFX2_23/A gnd sr[4] vdd BUFX2
XOAI21X1_8 BUFX2_23/A BUFX4_3/Y INVX4_1/Y gnd AOI21X1_7/C vdd OAI21X1
XNOR2X1_3 DFFSR_7/Q INVX1_3/Y gnd NOR2X1_3/Y vdd NOR2X1
XBUFX2_12 INVX1_5/A gnd dp[2] vdd BUFX2
XAOI21X1_5 BUFX4_1/Y MUX2X1_3/B OAI21X1_6/Y gnd DFFSR_19/D vdd AOI21X1
XFILL_1_2 gnd vdd FILL
XBUFX4_9 BUFX4_5/A gnd BUFX4_9/Y vdd BUFX4
XFILL_3_3_0 gnd vdd FILL
XBUFX2_24 INVX1_14/A gnd sr[5] vdd BUFX2
XFILL_8_2_0 gnd vdd FILL
XAOI21X1_6 BUFX4_3/Y INVX1_12/Y OAI21X1_7/Y gnd DFFSR_20/D vdd AOI21X1
XBUFX2_6 BUFX2_6/A gnd counter[5] vdd BUFX2
XFILL_0_1_0 gnd vdd FILL
XBUFX2_13 INVX1_7/A gnd dp[3] vdd BUFX2
XNAND2X1_1 INVX4_1/Y OAI21X1_1/Y gnd DFFSR_4/D vdd NAND2X1
XOAI21X1_9 INVX1_14/A BUFX4_3/Y INVX4_1/Y gnd OAI21X1_9/Y vdd OAI21X1
XAOI21X1_14 NOR2X1_12/Y INVX1_28/Y INVX4_1/A gnd AOI22X1_1/D vdd AOI21X1
XNOR2X1_4 BUFX2_19/A MUX2X1_2/S gnd NOR2X1_4/Y vdd NOR2X1
XFILL_5_0_0 gnd vdd FILL
XNOR2X1_5 N[0] MUX2X1_2/S gnd NOR2X1_5/Y vdd NOR2X1
XNAND2X1_2 N[1] N[2] gnd INVX2_1/A vdd NAND2X1
XBUFX2_25 BUFX2_25/A gnd sr[6] vdd BUFX2
XAOI21X1_7 BUFX4_3/Y INVX1_14/Y AOI21X1_7/C gnd DFFSR_21/D vdd AOI21X1
XBUFX2_14 INVX1_9/A gnd dp[4] vdd BUFX2
XBUFX2_7 BUFX2_7/A gnd counter[6] vdd BUFX2
XNAND2X1_3 INVX1_23/Y NOR2X1_9/B gnd INVX1_24/A vdd NAND2X1
XAOI21X1_8 BUFX4_3/Y MUX2X1_6/B OAI21X1_9/Y gnd DFFSR_22/D vdd AOI21X1
XBUFX2_8 BUFX2_8/A gnd counter[7] vdd BUFX2
XBUFX2_26 BUFX2_26/A gnd sr[7] vdd BUFX2
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XBUFX2_15 DFFSR_29/Q gnd dp[5] vdd BUFX2
XFILL_6_3_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XNAND2X1_4 NAND2X1_4/A NAND2X1_4/B gnd DFFSR_9/D vdd NAND2X1
XAOI21X1_9 BUFX4_4/Y MUX2X1_7/B AOI21X1_9/C gnd DFFSR_23/D vdd AOI21X1
XNOR2X1_7 BUFX2_1/A BUFX4_4/Y gnd NOR2X1_9/B vdd NOR2X1
XBUFX2_16 BUFX2_16/A gnd dp[6] vdd BUFX2
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XBUFX2_9 BUFX2_9/A gnd done vdd BUFX2
XFILL_8_0_0 gnd vdd FILL
XNAND2X1_5 INVX2_1/A NOR2X1_10/Y gnd NAND2X1_5/Y vdd NAND2X1
XNOR2X1_8 N[1] N[2] gnd NOR2X1_8/Y vdd NOR2X1
XBUFX2_17 INVX1_15/A gnd dp[7] vdd BUFX2
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XINVX1_20 BUFX2_9/A gnd INVX1_20/Y vdd INVX1
XBUFX2_18 INVX1_17/A gnd dp[8] vdd BUFX2
XNOR2X1_9 INVX1_23/Y NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XNAND2X1_6 INVX1_30/A NAND2X1_6/B gnd AOI22X1_1/B vdd NAND2X1
XINVX1_32 BUFX2_7/A gnd INVX1_32/Y vdd INVX1
XINVX1_10 BUFX2_22/A gnd MUX2X1_3/B vdd INVX1
XINVX1_21 DFFSR_3/Q gnd INVX1_21/Y vdd INVX1
XFILL_9_3_0 gnd vdd FILL
XFILL_8_1 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XDFFSR_30 BUFX2_16/A CLKBUF1_2/Y BUFX4_7/Y vdd DFFSR_30/D gnd vdd DFFSR
XFILL_6_1_0 gnd vdd FILL
XNAND2X1_7 NOR2X1_1/Y NOR2X1_2/Y gnd NOR2X1_14/B vdd NAND2X1
XINVX1_22 N[1] gnd INVX1_22/Y vdd INVX1
XBUFX2_19 BUFX2_19/A gnd sr[0] vdd BUFX2
XINVX1_11 DFFSR_29/Q gnd INVX1_11/Y vdd INVX1
XINVX1_33 N[8] gnd INVX1_33/Y vdd INVX1
XDFFSR_31 INVX1_15/A DFFSR_9/CLK DFFSR_9/R vdd MUX2X1_6/Y gnd vdd DFFSR
XDFFSR_20 BUFX2_23/A CLKBUF1_2/Y DFFSR_9/R vdd DFFSR_20/D gnd vdd DFFSR
XINVX1_23 BUFX2_2/A gnd INVX1_23/Y vdd INVX1
XINVX1_12 BUFX2_23/A gnd INVX1_12/Y vdd INVX1
XINVX1_34 BUFX2_8/A gnd INVX1_34/Y vdd INVX1
XDFFSR_32 INVX1_17/A DFFSR_9/CLK DFFSR_9/R vdd MUX2X1_7/Y gnd vdd DFFSR
XDFFSR_21 INVX1_14/A DFFSR_9/CLK BUFX4_6/Y vdd DFFSR_21/D gnd vdd DFFSR
XDFFSR_10 BUFX2_3/A DFFSR_8/CLK BUFX4_6/Y vdd DFFSR_10/D gnd vdd DFFSR
XNOR2X1_10 N[3] N[4] gnd NOR2X1_10/Y vdd NOR2X1
XNAND3X1_10 INVX4_1/A OAI21X1_29/Y NAND3X1_9/Y gnd AND2X2_3/B vdd NAND3X1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XINVX1_13 BUFX2_16/A gnd INVX1_13/Y vdd INVX1
XINVX1_35 INVX1_35/A gnd DFFSR_3/D vdd INVX1
XFILL_6_1 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XOAI21X1_30 BUFX4_2/Y NAND3X1_1/Y BUFX2_8/A gnd NAND3X1_12/B vdd OAI21X1
XFILL_9_1_0 gnd vdd FILL
XDFFSR_22 BUFX2_25/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_22/D gnd vdd DFFSR
XDFFSR_11 BUFX2_4/A DFFSR_8/CLK BUFX4_6/Y vdd DFFSR_11/D gnd vdd DFFSR
XFILL_1_0_0 gnd vdd FILL
XDFFSR_33 BUFX2_9/A DFFSR_5/CLK BUFX4_9/Y vdd DFFSR_33/D gnd vdd DFFSR
XINVX1_25 N[5] gnd INVX1_25/Y vdd INVX1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XNOR2X1_11 INVX1_26/Y INVX1_27/Y gnd NOR2X1_11/Y vdd NOR2X1
XNAND3X1_11 INVX8_1/A INVX1_34/Y AOI22X1_2/B gnd INVX1_35/A vdd NAND3X1
XOAI21X1_20 INVX4_1/A AND2X2_2/Y NAND3X1_4/Y gnd DFFSR_11/D vdd OAI21X1
XDFFSR_23 BUFX2_26/A DFFSR_9/CLK BUFX4_6/Y vdd DFFSR_23/D gnd vdd DFFSR
XDFFSR_12 BUFX2_5/A DFFSR_8/CLK BUFX4_6/Y vdd DFFSR_12/D gnd vdd DFFSR
XFILL_6_2 gnd vdd FILL
XNOR2X1_12 BUFX2_5/A AND2X2_2/B gnd NOR2X1_12/Y vdd NOR2X1
XNAND3X1_12 INVX4_1/Y NAND3X1_12/B INVX1_35/A gnd AND2X2_3/A vdd NAND3X1
XINVX1_15 INVX1_15/A gnd MUX2X1_6/A vdd INVX1
XINVX1_26 BUFX2_5/A gnd INVX1_26/Y vdd INVX1
XOAI21X1_21 N[5] NAND2X1_5/Y INVX4_1/A gnd OAI21X1_21/Y vdd OAI21X1
XOAI21X1_10 BUFX2_25/A BUFX4_4/Y INVX4_1/Y gnd AOI21X1_9/C vdd OAI21X1
XDFFSR_24 BUFX2_10/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_24/D gnd vdd DFFSR
XDFFSR_13 BUFX2_6/A DFFSR_8/CLK BUFX4_6/Y vdd DFFSR_13/D gnd vdd DFFSR
XFILL_2_3_0 gnd vdd FILL
XNOR2X1_13 N[5] N[6] gnd NOR2X1_13/Y vdd NOR2X1
XINVX1_16 BUFX2_25/A gnd MUX2X1_6/B vdd INVX1
XINVX1_27 AND2X2_2/B gnd INVX1_27/Y vdd INVX1
XDFFSR_1 INVX4_1/A DFFSR_5/CLK vdd BUFX4_9/Y DFFSR_1/D gnd vdd DFFSR
XFILL_7_2_0 gnd vdd FILL
XOAI21X1_22 NOR2X1_12/Y NOR2X1_11/Y INVX4_1/Y gnd OAI21X1_22/Y vdd OAI21X1
XOAI21X1_11 BUFX2_19/A BUFX4_1/Y INVX4_1/Y gnd AOI21X1_10/C vdd OAI21X1
XFILL_4_0_0 gnd vdd FILL
XDFFSR_14 BUFX2_7/A DFFSR_5/CLK BUFX4_9/Y vdd DFFSR_14/D gnd vdd DFFSR
XDFFSR_25 INVX1_4/A CLKBUF1_2/Y BUFX4_7/Y vdd DFFSR_25/D gnd vdd DFFSR
XFILL_4_1 gnd vdd FILL
XINVX1_17 INVX1_17/A gnd MUX2X1_7/A vdd INVX1
XINVX1_28 BUFX2_6/A gnd INVX1_28/Y vdd INVX1
XNOR2X1_14 NOR2X1_14/A NOR2X1_14/B gnd AOI22X1_2/B vdd NOR2X1
XDFFSR_2 DFFSR_2/Q DFFSR_5/CLK BUFX4_9/Y vdd DFFSR_2/D gnd vdd DFFSR
XOAI21X1_12 NOR2X1_9/B AND2X2_1/Y INVX4_1/Y gnd OAI21X1_13/C vdd OAI21X1
XOAI21X1_23 OAI21X1_23/A OAI21X1_21/Y OAI21X1_22/Y gnd DFFSR_12/D vdd OAI21X1
XDFFSR_15 BUFX2_8/A DFFSR_8/CLK BUFX4_7/Y vdd AND2X2_3/Y gnd vdd DFFSR
XDFFSR_26 INVX1_5/A DFFSR_3/CLK DFFSR_3/R vdd DFFSR_26/D gnd vdd DFFSR
XFILL_4_2 gnd vdd FILL
XDFFSR_3 DFFSR_3/Q DFFSR_3/CLK DFFSR_3/R vdd DFFSR_3/D gnd vdd DFFSR
XINVX1_18 BUFX2_26/A gnd MUX2X1_7/B vdd INVX1
XINVX1_29 N[7] gnd INVX1_29/Y vdd INVX1
XOAI21X1_24 N[5] NAND2X1_5/Y N[6] gnd NAND2X1_6/B vdd OAI21X1
XOAI21X1_13 INVX4_1/Y INVX1_22/Y OAI21X1_13/C gnd DFFSR_8/D vdd OAI21X1
XDFFSR_16 BUFX2_19/A CLKBUF1_2/Y DFFSR_9/R vdd NOR2X1_6/Y gnd vdd DFFSR
XDFFSR_27 INVX1_7/A DFFSR_3/CLK DFFSR_3/R vdd MUX2X1_2/Y gnd vdd DFFSR
XFILL_5_3_0 gnd vdd FILL
XFILL_4_3 gnd vdd FILL
XINVX1_19 BUFX2_10/A gnd INVX1_19/Y vdd INVX1
XFILL_2_1_0 gnd vdd FILL
XDFFSR_4 INVX8_1/A CLKBUF1_2/Y BUFX4_7/Y vdd DFFSR_4/D gnd vdd DFFSR
XOAI21X1_14 NOR2X1_8/Y INVX2_1/Y INVX4_1/A gnd NAND2X1_4/A vdd OAI21X1
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_25 BUFX2_5/A AND2X2_2/B BUFX2_6/A gnd AOI22X1_1/C vdd OAI21X1
XXNOR2X1_1 INVX1_14/A BUFX2_26/A gnd XNOR2X1_1/Y vdd XNOR2X1
XINVX1_1 DFFSR_2/Q gnd INVX1_1/Y vdd INVX1
XDFFSR_28 INVX1_9/A DFFSR_3/CLK DFFSR_3/R vdd DFFSR_28/D gnd vdd DFFSR
XDFFSR_17 INVX1_6/A CLKBUF1_2/Y BUFX4_7/Y vdd DFFSR_17/D gnd vdd DFFSR
XAND2X2_1 BUFX4_4/Y BUFX2_1/A gnd AND2X2_1/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XDFFSR_5 DFFSR_5/Q DFFSR_5/CLK BUFX4_7/Y vdd DFFSR_3/Q gnd vdd DFFSR
XOAI21X1_15 NOR2X1_9/Y INVX1_24/Y INVX4_1/Y gnd NAND2X1_4/B vdd OAI21X1
XDFFSR_29 DFFSR_29/Q CLKBUF1_2/Y BUFX4_7/Y vdd DFFSR_29/D gnd vdd DFFSR
XOAI21X1_26 N[7] INVX1_30/A INVX4_1/A gnd INVX1_31/A vdd OAI21X1
XDFFSR_18 INVX1_8/A DFFSR_3/CLK DFFSR_3/R vdd DFFSR_18/D gnd vdd DFFSR
XAND2X2_2 AND2X2_2/A AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XXNOR2X1_2 BUFX2_22/A BUFX2_23/A gnd XNOR2X1_2/Y vdd XNOR2X1
XINVX1_2 DFFSR_5/Q gnd INVX1_2/Y vdd INVX1
XDFFSR_6 DFFSR_6/Q DFFSR_5/CLK BUFX4_9/Y vdd start gnd vdd DFFSR
XOAI21X1_16 N[3] INVX2_1/Y OAI21X1_16/C gnd OAI21X1_16/Y vdd OAI21X1
XOAI21X1_27 INVX1_29/Y INVX1_30/Y INVX1_31/Y gnd OAI21X1_27/Y vdd OAI21X1
XFILL_8_3_0 gnd vdd FILL
XINVX1_3 DFFSR_6/Q gnd INVX1_3/Y vdd INVX1
XFILL_0_2_0 gnd vdd FILL
XDFFSR_19 BUFX2_22/A DFFSR_3/CLK DFFSR_3/R vdd DFFSR_19/D gnd vdd DFFSR
XFILL_5_1_0 gnd vdd FILL
XAND2X2_3 AND2X2_3/A AND2X2_3/B gnd AND2X2_3/Y vdd AND2X2
XDFFSR_7 DFFSR_7/Q DFFSR_5/CLK BUFX4_9/Y vdd DFFSR_6/Q gnd vdd DFFSR
XOAI21X1_17 INVX4_1/A XOR2X1_1/Y OAI21X1_16/Y gnd DFFSR_10/D vdd OAI21X1
XOAI21X1_28 INVX4_1/A AOI22X1_2/Y OAI21X1_27/Y gnd DFFSR_14/D vdd OAI21X1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XDFFSR_8 BUFX2_1/A DFFSR_8/CLK BUFX4_6/Y vdd DFFSR_8/D gnd vdd DFFSR
XAND2X2_4 NOR2X1_3/Y DFFSR_2/Q gnd DFFSR_1/D vdd AND2X2
XOAI21X1_18 N[3] INVX2_1/Y N[4] gnd NAND3X1_4/C vdd OAI21X1
XOAI21X1_29 N[7] INVX1_30/A INVX1_33/Y gnd OAI21X1_29/Y vdd OAI21X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
.ends


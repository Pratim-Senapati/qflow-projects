VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO noc_top
  CLASS BLOCK ;
  FOREIGN noc_top ;
  ORIGIN 1.900 4.000 ;
  SIZE 618.200 BY 568.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.400 560.400 614.000 561.600 ;
        RECT 2.800 555.800 3.600 560.400 ;
        RECT 4.400 555.800 5.200 560.400 ;
        RECT 7.600 555.800 8.400 560.400 ;
        RECT 10.800 555.800 11.600 560.400 ;
        RECT 17.200 555.800 18.000 560.400 ;
        RECT 20.400 555.800 21.200 560.400 ;
        RECT 28.400 555.800 29.200 560.400 ;
        RECT 31.600 555.800 32.400 560.400 ;
        RECT 34.800 555.800 35.600 560.400 ;
        RECT 38.000 555.800 38.800 560.400 ;
        RECT 41.200 553.000 42.000 560.400 ;
        RECT 44.400 555.800 45.200 560.400 ;
        RECT 47.600 555.800 48.400 560.400 ;
        RECT 50.800 555.800 51.600 560.400 ;
        RECT 7.600 551.800 8.400 552.400 ;
        RECT 11.000 551.800 11.800 552.000 ;
        RECT 52.400 551.800 53.200 560.400 ;
        RECT 56.600 555.800 57.400 560.400 ;
        RECT 58.800 551.800 59.600 560.400 ;
        RECT 63.000 555.800 63.800 560.400 ;
        RECT 65.200 555.800 66.000 560.400 ;
        RECT 68.400 555.800 69.200 560.400 ;
        RECT 71.600 555.800 72.400 560.400 ;
        RECT 74.800 555.800 75.600 560.400 ;
        RECT 82.800 555.800 83.600 560.400 ;
        RECT 86.000 555.800 86.800 560.400 ;
        RECT 92.400 555.800 93.200 560.400 ;
        RECT 95.600 555.800 96.400 560.400 ;
        RECT 98.800 555.800 99.600 560.400 ;
        RECT 92.200 551.800 93.000 552.000 ;
        RECT 95.600 551.800 96.400 552.400 ;
        RECT 102.000 552.000 102.800 560.400 ;
        RECT 107.600 555.800 108.400 560.400 ;
        RECT 110.800 555.800 111.600 560.400 ;
        RECT 116.400 551.800 117.200 560.400 ;
        RECT 121.200 552.000 122.000 560.400 ;
        RECT 126.800 555.800 127.600 560.400 ;
        RECT 130.000 555.800 130.800 560.400 ;
        RECT 135.600 551.800 136.400 560.400 ;
        RECT 143.600 555.800 144.400 560.400 ;
        RECT 146.800 555.800 147.600 560.400 ;
        RECT 150.000 555.800 150.800 560.400 ;
        RECT 156.400 555.800 157.200 560.400 ;
        RECT 159.600 555.800 160.400 560.400 ;
        RECT 167.600 555.800 168.400 560.400 ;
        RECT 170.800 555.800 171.600 560.400 ;
        RECT 174.000 555.800 174.800 560.400 ;
        RECT 177.200 555.800 178.000 560.400 ;
        RECT 180.400 553.000 181.200 560.400 ;
        RECT 183.600 555.800 184.400 560.400 ;
        RECT 187.400 555.800 188.200 560.400 ;
        RECT 146.800 551.800 147.600 552.400 ;
        RECT 150.200 551.800 151.000 552.000 ;
        RECT 191.600 551.800 192.400 560.400 ;
        RECT 193.200 555.800 194.000 560.400 ;
        RECT 196.400 555.800 197.200 560.400 ;
        RECT 199.600 553.000 200.400 560.400 ;
        RECT 202.800 555.800 203.600 560.400 ;
        RECT 206.000 555.800 206.800 560.400 ;
        RECT 209.200 555.800 210.000 560.400 ;
        RECT 215.600 555.800 216.400 560.400 ;
        RECT 218.800 555.800 219.600 560.400 ;
        RECT 226.800 555.800 227.600 560.400 ;
        RECT 230.000 555.800 230.800 560.400 ;
        RECT 233.200 555.800 234.000 560.400 ;
        RECT 236.400 555.800 237.200 560.400 ;
        RECT 238.000 555.800 238.800 560.400 ;
        RECT 206.000 551.800 206.800 552.400 ;
        RECT 209.400 551.800 210.200 552.000 ;
        RECT 241.200 551.800 242.000 560.400 ;
        RECT 245.400 555.800 246.200 560.400 ;
        RECT 247.600 555.800 248.400 560.400 ;
        RECT 250.800 555.800 251.600 560.400 ;
        RECT 254.000 553.000 254.800 560.400 ;
        RECT 257.200 555.800 258.000 560.400 ;
        RECT 260.400 555.800 261.200 560.400 ;
        RECT 263.600 555.800 264.400 560.400 ;
        RECT 270.000 555.800 270.800 560.400 ;
        RECT 273.200 555.800 274.000 560.400 ;
        RECT 281.200 555.800 282.000 560.400 ;
        RECT 284.400 555.800 285.200 560.400 ;
        RECT 287.600 555.800 288.400 560.400 ;
        RECT 290.800 555.800 291.600 560.400 ;
        RECT 294.000 553.000 294.800 560.400 ;
        RECT 302.000 555.800 302.800 560.400 ;
        RECT 305.200 555.800 306.000 560.400 ;
        RECT 308.400 555.800 309.200 560.400 ;
        RECT 311.600 555.800 312.400 560.400 ;
        RECT 319.600 555.800 320.400 560.400 ;
        RECT 322.800 555.800 323.600 560.400 ;
        RECT 329.200 555.800 330.000 560.400 ;
        RECT 332.400 555.800 333.200 560.400 ;
        RECT 335.600 555.800 336.400 560.400 ;
        RECT 337.200 555.800 338.000 560.400 ;
        RECT 260.400 551.800 261.200 552.400 ;
        RECT 263.800 551.800 264.600 552.000 ;
        RECT 329.000 551.800 329.800 552.000 ;
        RECT 332.400 551.800 333.200 552.400 ;
        RECT 340.400 551.800 341.200 560.400 ;
        RECT 344.600 555.800 345.400 560.400 ;
        RECT 347.400 555.800 348.200 560.400 ;
        RECT 351.600 551.800 352.400 560.400 ;
        RECT 353.200 555.800 354.000 560.400 ;
        RECT 356.400 551.800 357.200 560.400 ;
        RECT 360.600 555.800 361.400 560.400 ;
        RECT 362.800 551.800 363.600 560.400 ;
        RECT 367.000 555.800 367.800 560.400 ;
        RECT 369.200 555.800 370.000 560.400 ;
        RECT 372.400 555.800 373.200 560.400 ;
        RECT 375.600 555.800 376.400 560.400 ;
        RECT 378.800 555.800 379.600 560.400 ;
        RECT 386.800 555.800 387.600 560.400 ;
        RECT 390.000 555.800 390.800 560.400 ;
        RECT 396.400 555.800 397.200 560.400 ;
        RECT 399.600 555.800 400.400 560.400 ;
        RECT 402.800 555.800 403.600 560.400 ;
        RECT 396.200 551.800 397.200 552.000 ;
        RECT 399.600 551.800 400.400 552.400 ;
        RECT 404.400 551.800 405.200 560.400 ;
        RECT 407.600 551.800 408.400 560.400 ;
        RECT 410.800 551.800 411.600 560.400 ;
        RECT 414.000 551.800 414.800 560.400 ;
        RECT 417.200 551.800 418.000 560.400 ;
        RECT 420.400 551.800 421.200 560.400 ;
        RECT 426.000 555.800 426.800 560.400 ;
        RECT 429.200 555.800 430.000 560.400 ;
        RECT 434.800 552.000 435.600 560.400 ;
        RECT 438.000 551.800 438.800 560.400 ;
        RECT 442.200 555.800 443.000 560.400 ;
        RECT 445.000 555.800 445.800 560.400 ;
        RECT 449.200 551.800 450.000 560.400 ;
        RECT 453.000 551.800 453.800 560.400 ;
        RECT 463.600 551.800 464.400 560.400 ;
        RECT 469.200 555.800 470.000 560.400 ;
        RECT 472.400 555.800 473.200 560.400 ;
        RECT 478.000 552.000 478.800 560.400 ;
        RECT 481.200 551.800 482.000 560.400 ;
        RECT 485.400 555.800 486.200 560.400 ;
        RECT 488.200 555.800 489.000 560.400 ;
        RECT 492.400 551.800 493.200 560.400 ;
        RECT 495.600 551.800 496.400 560.400 ;
        RECT 501.200 555.800 502.000 560.400 ;
        RECT 504.400 555.800 505.200 560.400 ;
        RECT 510.000 552.000 510.800 560.400 ;
        RECT 513.200 551.800 514.000 560.400 ;
        RECT 517.400 555.800 518.200 560.400 ;
        RECT 521.200 552.200 522.000 560.400 ;
        RECT 526.400 551.800 527.200 560.400 ;
        RECT 529.800 555.800 530.600 560.400 ;
        RECT 534.000 551.800 534.800 560.400 ;
        RECT 535.600 555.800 536.400 560.400 ;
        RECT 540.400 551.800 541.200 560.400 ;
        RECT 546.000 555.800 546.800 560.400 ;
        RECT 549.200 555.800 550.000 560.400 ;
        RECT 554.800 552.000 555.600 560.400 ;
        RECT 558.000 555.800 558.800 560.400 ;
        RECT 561.200 555.800 562.000 560.400 ;
        RECT 564.400 555.800 565.200 560.400 ;
        RECT 567.600 555.800 568.400 560.400 ;
        RECT 575.600 555.800 576.400 560.400 ;
        RECT 578.800 555.800 579.600 560.400 ;
        RECT 585.200 555.800 586.000 560.400 ;
        RECT 588.400 555.800 589.200 560.400 ;
        RECT 591.600 555.800 592.400 560.400 ;
        RECT 594.800 555.800 595.600 560.400 ;
        RECT 585.000 551.800 586.000 552.000 ;
        RECT 588.400 551.800 589.200 552.400 ;
        RECT 596.400 551.800 597.200 560.400 ;
        RECT 599.600 551.800 600.400 560.400 ;
        RECT 602.800 551.800 603.600 560.400 ;
        RECT 606.000 551.800 606.800 560.400 ;
        RECT 609.200 551.800 610.000 560.400 ;
        RECT 7.600 551.200 34.600 551.800 ;
        RECT 33.800 551.000 34.600 551.200 ;
        RECT 69.400 551.200 96.400 551.800 ;
        RECT 146.800 551.200 173.800 551.800 ;
        RECT 206.000 551.200 233.000 551.800 ;
        RECT 260.400 551.200 287.400 551.800 ;
        RECT 69.400 551.000 70.200 551.200 ;
        RECT 173.000 551.000 173.800 551.200 ;
        RECT 232.200 551.000 233.000 551.200 ;
        RECT 286.600 551.000 287.400 551.200 ;
        RECT 306.200 551.200 333.200 551.800 ;
        RECT 373.400 551.200 400.400 551.800 ;
        RECT 562.200 551.200 589.200 551.800 ;
        RECT 306.200 551.000 307.000 551.200 ;
        RECT 373.400 551.000 374.200 551.200 ;
        RECT 562.200 551.000 563.000 551.200 ;
        RECT 30.600 530.800 31.400 531.000 ;
        RECT 4.400 530.200 31.400 530.800 ;
        RECT 67.800 530.800 68.600 531.000 ;
        RECT 144.600 530.800 145.400 531.000 ;
        RECT 205.000 530.800 205.800 531.000 ;
        RECT 67.800 530.200 94.800 530.800 ;
        RECT 144.600 530.200 171.600 530.800 ;
        RECT 4.400 529.600 5.200 530.200 ;
        RECT 7.600 530.000 8.600 530.200 ;
        RECT 1.200 521.600 2.000 526.200 ;
        RECT 4.400 521.600 5.200 526.200 ;
        RECT 7.600 521.600 8.400 526.200 ;
        RECT 14.000 521.600 14.800 526.200 ;
        RECT 17.200 521.600 18.000 526.200 ;
        RECT 25.200 521.600 26.000 526.200 ;
        RECT 28.400 521.600 29.200 526.200 ;
        RECT 31.600 521.600 32.400 526.200 ;
        RECT 34.800 521.600 35.600 526.200 ;
        RECT 37.000 521.600 37.800 526.200 ;
        RECT 41.200 521.600 42.000 530.200 ;
        RECT 42.800 521.600 43.600 526.200 ;
        RECT 46.000 521.600 46.800 526.200 ;
        RECT 47.600 521.600 48.400 526.200 ;
        RECT 50.800 521.600 51.600 530.200 ;
        RECT 55.000 521.600 55.800 526.200 ;
        RECT 57.200 521.600 58.000 530.200 ;
        RECT 90.600 530.000 91.400 530.200 ;
        RECT 94.000 529.600 94.800 530.200 ;
        RECT 61.400 521.600 62.200 526.200 ;
        RECT 63.600 521.600 64.400 526.200 ;
        RECT 66.800 521.600 67.600 526.200 ;
        RECT 70.000 521.600 70.800 526.200 ;
        RECT 73.200 521.600 74.000 526.200 ;
        RECT 81.200 521.600 82.000 526.200 ;
        RECT 84.400 521.600 85.200 526.200 ;
        RECT 90.800 521.600 91.600 526.200 ;
        RECT 94.000 521.600 94.800 526.200 ;
        RECT 97.200 521.600 98.000 526.200 ;
        RECT 98.800 521.600 99.600 530.200 ;
        RECT 103.000 521.600 103.800 526.200 ;
        RECT 105.200 521.600 106.000 530.200 ;
        RECT 109.400 521.600 110.200 526.200 ;
        RECT 111.600 521.600 112.400 530.200 ;
        RECT 115.800 521.600 116.600 526.200 ;
        RECT 118.600 521.600 119.400 526.200 ;
        RECT 122.800 521.600 123.600 530.200 ;
        RECT 167.400 530.000 168.200 530.200 ;
        RECT 170.800 529.600 171.600 530.200 ;
        RECT 178.800 530.200 205.800 530.800 ;
        RECT 229.400 530.800 230.200 531.000 ;
        RECT 289.800 530.800 290.600 531.000 ;
        RECT 229.400 530.200 256.400 530.800 ;
        RECT 178.800 529.600 179.600 530.200 ;
        RECT 182.000 530.000 183.000 530.200 ;
        RECT 126.000 522.200 127.000 528.800 ;
        RECT 126.200 521.600 127.000 522.200 ;
        RECT 132.200 521.600 133.200 528.800 ;
        RECT 140.400 521.600 141.200 526.200 ;
        RECT 143.600 521.600 144.400 526.200 ;
        RECT 146.800 521.600 147.600 526.200 ;
        RECT 150.000 521.600 150.800 526.200 ;
        RECT 158.000 521.600 158.800 526.200 ;
        RECT 161.200 521.600 162.000 526.200 ;
        RECT 167.600 521.600 168.400 526.200 ;
        RECT 170.800 521.600 171.600 526.200 ;
        RECT 174.000 521.600 174.800 526.200 ;
        RECT 175.600 521.600 176.400 526.200 ;
        RECT 178.800 521.600 179.600 526.200 ;
        RECT 182.000 521.600 182.800 526.200 ;
        RECT 188.400 521.600 189.200 526.200 ;
        RECT 191.600 521.600 192.400 526.200 ;
        RECT 199.600 521.600 200.400 526.200 ;
        RECT 202.800 521.600 203.600 526.200 ;
        RECT 206.000 521.600 206.800 526.200 ;
        RECT 209.200 521.600 210.000 526.200 ;
        RECT 210.800 521.600 211.600 526.200 ;
        RECT 214.000 521.600 214.800 530.200 ;
        RECT 252.200 530.000 253.000 530.200 ;
        RECT 255.600 529.600 256.400 530.200 ;
        RECT 263.600 530.200 290.600 530.800 ;
        RECT 319.000 530.800 319.800 531.000 ;
        RECT 386.200 530.800 387.000 531.000 ;
        RECT 547.800 530.800 548.600 531.000 ;
        RECT 319.000 530.200 346.000 530.800 ;
        RECT 386.200 530.200 413.200 530.800 ;
        RECT 547.800 530.200 574.800 530.800 ;
        RECT 263.600 529.600 264.400 530.200 ;
        RECT 267.000 530.000 267.800 530.200 ;
        RECT 218.200 521.600 219.000 526.200 ;
        RECT 220.400 521.600 221.200 526.200 ;
        RECT 223.600 521.600 224.400 526.200 ;
        RECT 225.200 521.600 226.000 526.200 ;
        RECT 228.400 521.600 229.200 526.200 ;
        RECT 231.600 521.600 232.400 526.200 ;
        RECT 234.800 521.600 235.600 526.200 ;
        RECT 242.800 521.600 243.600 526.200 ;
        RECT 246.000 521.600 246.800 526.200 ;
        RECT 252.400 521.600 253.200 526.200 ;
        RECT 255.600 521.600 256.400 526.200 ;
        RECT 258.800 521.600 259.600 526.200 ;
        RECT 260.400 521.600 261.200 526.200 ;
        RECT 263.600 521.600 264.400 526.200 ;
        RECT 266.800 521.600 267.600 526.200 ;
        RECT 273.200 521.600 274.000 526.200 ;
        RECT 276.400 521.600 277.200 526.200 ;
        RECT 284.400 521.600 285.200 526.200 ;
        RECT 287.600 521.600 288.400 526.200 ;
        RECT 290.800 521.600 291.600 526.200 ;
        RECT 294.000 521.600 294.800 526.200 ;
        RECT 295.600 521.600 296.400 526.200 ;
        RECT 298.800 521.600 299.600 530.200 ;
        RECT 341.800 530.000 342.800 530.200 ;
        RECT 345.200 529.600 346.000 530.200 ;
        RECT 303.000 521.600 303.800 526.200 ;
        RECT 310.000 521.600 310.800 526.200 ;
        RECT 313.200 521.600 314.000 526.200 ;
        RECT 314.800 521.600 315.600 526.200 ;
        RECT 318.000 521.600 318.800 526.200 ;
        RECT 321.200 521.600 322.000 526.200 ;
        RECT 324.400 521.600 325.200 526.200 ;
        RECT 332.400 521.600 333.200 526.200 ;
        RECT 335.600 521.600 336.400 526.200 ;
        RECT 342.000 521.600 342.800 526.200 ;
        RECT 345.200 521.600 346.000 526.200 ;
        RECT 348.400 521.600 349.200 526.200 ;
        RECT 350.600 521.600 351.400 526.200 ;
        RECT 354.800 521.600 355.600 530.200 ;
        RECT 358.000 521.600 358.800 526.200 ;
        RECT 360.200 521.600 361.000 526.200 ;
        RECT 364.400 521.600 365.200 530.200 ;
        RECT 366.000 521.600 366.800 530.200 ;
        RECT 370.200 521.600 371.000 526.200 ;
        RECT 372.400 521.600 373.200 526.200 ;
        RECT 375.600 521.600 376.400 530.200 ;
        RECT 409.000 530.000 410.000 530.200 ;
        RECT 412.400 529.600 413.200 530.200 ;
        RECT 379.800 521.600 380.600 526.200 ;
        RECT 382.000 521.600 382.800 526.200 ;
        RECT 385.200 521.600 386.000 526.200 ;
        RECT 388.400 521.600 389.200 526.200 ;
        RECT 391.600 521.600 392.400 526.200 ;
        RECT 399.600 521.600 400.400 526.200 ;
        RECT 402.800 521.600 403.600 526.200 ;
        RECT 409.200 521.600 410.000 526.200 ;
        RECT 412.400 521.600 413.200 526.200 ;
        RECT 415.600 521.600 416.400 526.200 ;
        RECT 417.200 521.600 418.000 530.200 ;
        RECT 420.400 521.600 421.200 530.200 ;
        RECT 423.600 521.600 424.400 530.200 ;
        RECT 426.800 521.600 427.600 530.200 ;
        RECT 430.000 521.600 430.800 530.200 ;
        RECT 433.200 521.600 434.000 530.200 ;
        RECT 438.800 521.600 439.600 526.200 ;
        RECT 442.000 521.600 442.800 526.200 ;
        RECT 447.600 521.600 448.400 530.000 ;
        RECT 450.800 521.600 451.600 530.200 ;
        RECT 455.000 521.600 455.800 526.200 ;
        RECT 462.600 521.600 463.400 526.200 ;
        RECT 466.800 521.600 467.600 530.200 ;
        RECT 470.000 521.600 470.800 529.000 ;
        RECT 473.200 521.600 474.000 530.200 ;
        RECT 474.800 521.600 475.600 530.200 ;
        RECT 479.000 521.600 479.800 526.200 ;
        RECT 481.800 521.600 482.600 526.200 ;
        RECT 486.000 521.600 486.800 530.200 ;
        RECT 487.600 521.600 488.400 530.200 ;
        RECT 491.800 521.600 492.600 526.200 ;
        RECT 494.600 521.600 495.400 526.200 ;
        RECT 498.800 521.600 499.600 530.200 ;
        RECT 502.000 521.600 502.800 530.000 ;
        RECT 507.600 521.600 508.400 526.200 ;
        RECT 510.800 521.600 511.600 526.200 ;
        RECT 516.400 521.600 517.200 530.200 ;
        RECT 519.600 521.600 520.400 526.200 ;
        RECT 522.800 521.600 523.600 526.200 ;
        RECT 526.000 521.600 526.800 529.000 ;
        RECT 529.200 521.600 530.000 530.200 ;
        RECT 532.400 521.600 533.200 529.000 ;
        RECT 535.600 521.600 536.400 530.200 ;
        RECT 537.200 521.600 538.000 530.200 ;
        RECT 570.600 530.000 571.400 530.200 ;
        RECT 574.000 529.600 574.800 530.200 ;
        RECT 541.400 521.600 542.200 526.200 ;
        RECT 543.600 521.600 544.400 526.200 ;
        RECT 546.800 521.600 547.600 526.200 ;
        RECT 550.000 521.600 550.800 526.200 ;
        RECT 553.200 521.600 554.000 526.200 ;
        RECT 561.200 521.600 562.000 526.200 ;
        RECT 564.400 521.600 565.200 526.200 ;
        RECT 570.800 521.600 571.600 526.200 ;
        RECT 574.000 521.600 574.800 526.200 ;
        RECT 577.200 521.600 578.000 526.200 ;
        RECT 578.800 521.600 579.600 530.200 ;
        RECT 583.000 521.600 583.800 526.200 ;
        RECT 585.200 521.600 586.000 530.200 ;
        RECT 588.400 521.600 589.200 530.200 ;
        RECT 591.600 521.600 592.400 530.200 ;
        RECT 594.800 521.600 595.600 530.200 ;
        RECT 598.000 521.600 598.800 530.200 ;
        RECT 600.200 521.600 601.000 526.200 ;
        RECT 604.400 521.600 605.200 530.200 ;
        RECT 607.600 521.600 608.400 526.200 ;
        RECT 0.400 520.400 614.000 521.600 ;
        RECT 2.800 512.000 3.600 520.400 ;
        RECT 8.400 515.800 9.200 520.400 ;
        RECT 11.600 515.800 12.400 520.400 ;
        RECT 17.200 511.800 18.000 520.400 ;
        RECT 22.000 512.000 22.800 520.400 ;
        RECT 27.600 515.800 28.400 520.400 ;
        RECT 30.800 515.800 31.600 520.400 ;
        RECT 36.400 511.800 37.200 520.400 ;
        RECT 39.600 511.800 40.400 520.400 ;
        RECT 43.800 515.800 44.600 520.400 ;
        RECT 47.600 512.200 48.400 520.400 ;
        RECT 52.800 511.800 53.600 520.400 ;
        RECT 56.200 515.800 57.000 520.400 ;
        RECT 60.400 511.800 61.200 520.400 ;
        RECT 62.000 511.800 62.800 520.400 ;
        RECT 66.200 515.800 67.000 520.400 ;
        RECT 69.000 515.800 69.800 520.400 ;
        RECT 73.200 511.800 74.000 520.400 ;
        RECT 76.400 512.000 77.200 520.400 ;
        RECT 82.000 515.800 82.800 520.400 ;
        RECT 85.200 515.800 86.000 520.400 ;
        RECT 90.800 511.800 91.600 520.400 ;
        RECT 95.600 512.000 96.400 520.400 ;
        RECT 101.200 515.800 102.000 520.400 ;
        RECT 104.400 515.800 105.200 520.400 ;
        RECT 110.000 511.800 110.800 520.400 ;
        RECT 114.800 515.800 115.600 520.400 ;
        RECT 116.400 515.800 117.200 520.400 ;
        RECT 120.800 511.800 121.600 520.400 ;
        RECT 126.000 512.200 126.800 520.400 ;
        RECT 130.800 512.200 131.600 520.400 ;
        RECT 136.000 511.800 136.800 520.400 ;
        RECT 138.800 511.800 139.600 520.400 ;
        RECT 143.600 515.800 144.400 520.400 ;
        RECT 151.600 511.800 152.400 520.400 ;
        RECT 154.800 511.800 155.600 520.400 ;
        RECT 158.000 511.800 158.800 520.400 ;
        RECT 161.200 511.800 162.000 520.400 ;
        RECT 164.400 511.800 165.200 520.400 ;
        RECT 166.000 515.800 166.800 520.400 ;
        RECT 169.200 511.800 170.000 520.400 ;
        RECT 175.600 513.200 176.600 520.400 ;
        RECT 181.800 519.800 182.600 520.400 ;
        RECT 181.800 513.200 182.800 519.800 ;
        RECT 185.200 511.800 186.000 520.400 ;
        RECT 188.400 511.800 189.200 520.400 ;
        RECT 191.600 511.800 192.400 520.400 ;
        RECT 194.800 511.800 195.600 520.400 ;
        RECT 198.000 511.800 198.800 520.400 ;
        RECT 199.600 515.800 200.400 520.400 ;
        RECT 202.800 515.800 203.600 520.400 ;
        RECT 206.000 515.800 206.800 520.400 ;
        RECT 212.400 515.800 213.200 520.400 ;
        RECT 215.600 515.800 216.400 520.400 ;
        RECT 223.600 515.800 224.400 520.400 ;
        RECT 226.800 515.800 227.600 520.400 ;
        RECT 230.000 515.800 230.800 520.400 ;
        RECT 233.200 515.800 234.000 520.400 ;
        RECT 235.400 515.800 236.200 520.400 ;
        RECT 202.800 511.800 203.600 512.400 ;
        RECT 206.200 511.800 207.000 512.000 ;
        RECT 239.600 511.800 240.400 520.400 ;
        RECT 241.200 515.800 242.000 520.400 ;
        RECT 244.400 515.800 245.200 520.400 ;
        RECT 246.000 515.800 246.800 520.400 ;
        RECT 249.200 515.800 250.000 520.400 ;
        RECT 252.400 515.800 253.200 520.400 ;
        RECT 255.600 515.800 256.400 520.400 ;
        RECT 262.000 515.800 262.800 520.400 ;
        RECT 265.200 515.800 266.000 520.400 ;
        RECT 273.200 515.800 274.000 520.400 ;
        RECT 276.400 515.800 277.200 520.400 ;
        RECT 279.600 515.800 280.400 520.400 ;
        RECT 282.800 515.800 283.600 520.400 ;
        RECT 284.400 515.800 285.200 520.400 ;
        RECT 287.600 515.800 288.400 520.400 ;
        RECT 290.800 515.800 291.600 520.400 ;
        RECT 297.200 515.800 298.000 520.400 ;
        RECT 300.400 515.800 301.200 520.400 ;
        RECT 308.400 515.800 309.200 520.400 ;
        RECT 311.600 515.800 312.400 520.400 ;
        RECT 314.800 515.800 315.600 520.400 ;
        RECT 318.000 515.800 318.800 520.400 ;
        RECT 324.400 515.800 325.200 520.400 ;
        RECT 327.600 515.800 328.400 520.400 ;
        RECT 329.200 515.800 330.000 520.400 ;
        RECT 332.400 515.800 333.200 520.400 ;
        RECT 252.400 511.800 253.200 512.400 ;
        RECT 255.600 511.800 256.600 512.000 ;
        RECT 287.600 511.800 288.400 512.400 ;
        RECT 335.600 512.000 336.400 520.400 ;
        RECT 341.200 515.800 342.000 520.400 ;
        RECT 344.400 515.800 345.200 520.400 ;
        RECT 291.000 511.800 291.800 512.000 ;
        RECT 350.000 511.800 350.800 520.400 ;
        RECT 353.200 515.800 354.000 520.400 ;
        RECT 356.400 515.800 357.200 520.400 ;
        RECT 359.600 512.000 360.400 520.400 ;
        RECT 365.200 515.800 366.000 520.400 ;
        RECT 368.400 515.800 369.200 520.400 ;
        RECT 374.000 511.800 374.800 520.400 ;
        RECT 378.800 512.200 379.600 520.400 ;
        RECT 384.000 511.800 384.800 520.400 ;
        RECT 386.800 511.800 387.600 520.400 ;
        RECT 391.000 515.800 391.800 520.400 ;
        RECT 393.200 515.800 394.000 520.400 ;
        RECT 396.400 515.800 397.200 520.400 ;
        RECT 398.600 515.800 399.400 520.400 ;
        RECT 402.800 511.800 403.600 520.400 ;
        RECT 404.400 511.800 405.200 520.400 ;
        RECT 407.600 513.000 408.400 520.400 ;
        RECT 410.800 515.800 411.600 520.400 ;
        RECT 415.200 511.800 416.000 520.400 ;
        RECT 420.400 512.200 421.200 520.400 ;
        RECT 423.600 511.800 424.400 520.400 ;
        RECT 427.800 515.800 428.600 520.400 ;
        RECT 430.000 511.800 430.800 520.400 ;
        RECT 433.200 513.000 434.000 520.400 ;
        RECT 436.400 515.800 437.200 520.400 ;
        RECT 439.600 515.800 440.400 520.400 ;
        RECT 442.800 513.000 443.600 520.400 ;
        RECT 446.000 511.800 446.800 520.400 ;
        RECT 448.800 511.800 449.600 520.400 ;
        RECT 454.000 512.200 454.800 520.400 ;
        RECT 463.600 515.800 464.400 520.400 ;
        RECT 465.200 515.800 466.000 520.400 ;
        RECT 468.400 515.800 469.200 520.400 ;
        RECT 471.600 512.200 472.400 520.400 ;
        RECT 476.800 511.800 477.600 520.400 ;
        RECT 479.600 515.800 480.400 520.400 ;
        RECT 482.800 515.800 483.600 520.400 ;
        RECT 485.600 511.800 486.400 520.400 ;
        RECT 490.800 512.200 491.600 520.400 ;
        RECT 494.000 511.800 494.800 520.400 ;
        RECT 497.200 513.000 498.000 520.400 ;
        RECT 500.400 515.800 501.200 520.400 ;
        RECT 503.600 515.800 504.400 520.400 ;
        RECT 506.800 513.000 507.600 520.400 ;
        RECT 510.000 511.800 510.800 520.400 ;
        RECT 511.600 511.800 512.400 520.400 ;
        RECT 515.800 515.800 516.600 520.400 ;
        RECT 519.600 515.800 520.400 520.400 ;
        RECT 522.800 512.200 523.600 520.400 ;
        RECT 528.000 511.800 528.800 520.400 ;
        RECT 530.800 511.800 531.600 520.400 ;
        RECT 535.000 515.800 535.800 520.400 ;
        RECT 537.200 511.800 538.000 520.400 ;
        RECT 541.400 515.800 542.200 520.400 ;
        RECT 543.600 511.800 544.400 520.400 ;
        RECT 547.800 515.800 548.600 520.400 ;
        RECT 551.600 511.800 552.400 520.400 ;
        RECT 557.200 515.800 558.000 520.400 ;
        RECT 560.400 515.800 561.200 520.400 ;
        RECT 566.000 512.000 566.800 520.400 ;
        RECT 569.200 515.800 570.000 520.400 ;
        RECT 572.400 515.800 573.200 520.400 ;
        RECT 574.000 515.800 574.800 520.400 ;
        RECT 577.200 515.800 578.000 520.400 ;
        RECT 580.400 515.800 581.200 520.400 ;
        RECT 583.600 515.800 584.400 520.400 ;
        RECT 591.600 515.800 592.400 520.400 ;
        RECT 594.800 515.800 595.600 520.400 ;
        RECT 601.200 515.800 602.000 520.400 ;
        RECT 604.400 515.800 605.200 520.400 ;
        RECT 607.600 515.800 608.400 520.400 ;
        RECT 601.000 511.800 602.000 512.000 ;
        RECT 604.400 511.800 605.200 512.400 ;
        RECT 202.800 511.200 229.800 511.800 ;
        RECT 252.400 511.200 279.400 511.800 ;
        RECT 287.600 511.200 314.600 511.800 ;
        RECT 229.000 511.000 229.800 511.200 ;
        RECT 278.600 511.000 279.400 511.200 ;
        RECT 313.800 511.000 314.600 511.200 ;
        RECT 578.200 511.200 605.200 511.800 ;
        RECT 578.200 511.000 579.000 511.200 ;
        RECT 133.400 490.800 134.200 491.000 ;
        RECT 178.200 490.800 179.000 491.000 ;
        RECT 213.400 490.800 214.200 491.000 ;
        RECT 581.400 490.800 582.200 491.000 ;
        RECT 133.400 490.200 160.400 490.800 ;
        RECT 178.200 490.200 205.200 490.800 ;
        RECT 213.400 490.200 240.400 490.800 ;
        RECT 581.400 490.200 608.400 490.800 ;
        RECT 1.800 481.600 2.600 486.200 ;
        RECT 6.000 481.600 6.800 490.200 ;
        RECT 8.800 481.600 9.600 490.200 ;
        RECT 14.000 481.600 14.800 489.800 ;
        RECT 17.800 481.600 18.600 486.200 ;
        RECT 22.000 481.600 22.800 490.200 ;
        RECT 25.200 481.600 26.000 490.000 ;
        RECT 30.800 481.600 31.600 486.200 ;
        RECT 34.000 481.600 34.800 486.200 ;
        RECT 39.600 481.600 40.400 490.200 ;
        RECT 42.800 481.600 43.600 490.200 ;
        RECT 47.000 481.600 47.800 486.200 ;
        RECT 50.400 481.600 51.200 490.200 ;
        RECT 55.600 481.600 56.400 489.800 ;
        RECT 59.400 481.600 60.200 486.200 ;
        RECT 63.600 481.600 64.400 490.200 ;
        RECT 66.800 481.600 67.600 489.800 ;
        RECT 72.000 481.600 72.800 490.200 ;
        RECT 74.800 481.600 75.600 486.200 ;
        RECT 78.000 481.600 78.800 486.200 ;
        RECT 79.600 481.600 80.400 486.200 ;
        RECT 82.800 481.600 83.600 486.200 ;
        RECT 84.400 481.600 85.200 486.200 ;
        RECT 87.600 481.600 88.400 490.200 ;
        RECT 91.800 481.600 92.600 486.200 ;
        RECT 94.600 481.600 95.400 486.200 ;
        RECT 98.800 481.600 99.600 490.200 ;
        RECT 101.000 481.600 101.800 486.200 ;
        RECT 105.200 481.600 106.000 490.200 ;
        RECT 106.800 481.600 107.600 486.200 ;
        RECT 110.000 481.600 110.800 485.800 ;
        RECT 113.800 481.600 114.600 486.200 ;
        RECT 118.000 481.600 118.800 490.200 ;
        RECT 119.600 481.600 120.400 486.200 ;
        RECT 122.800 481.600 123.600 486.200 ;
        RECT 127.600 481.600 128.400 490.200 ;
        RECT 156.200 490.000 157.000 490.200 ;
        RECT 159.600 489.600 160.400 490.200 ;
        RECT 129.200 481.600 130.000 486.200 ;
        RECT 132.400 481.600 133.200 486.200 ;
        RECT 135.600 481.600 136.400 486.200 ;
        RECT 138.800 481.600 139.600 486.200 ;
        RECT 146.800 481.600 147.600 486.200 ;
        RECT 150.000 481.600 150.800 486.200 ;
        RECT 156.400 481.600 157.200 486.200 ;
        RECT 159.600 481.600 160.400 486.200 ;
        RECT 162.800 481.600 163.600 486.200 ;
        RECT 172.400 481.600 173.200 490.200 ;
        RECT 201.000 490.000 201.800 490.200 ;
        RECT 204.400 489.600 205.200 490.200 ;
        RECT 236.200 490.000 237.000 490.200 ;
        RECT 239.600 489.600 240.400 490.200 ;
        RECT 174.000 481.600 174.800 486.200 ;
        RECT 177.200 481.600 178.000 486.200 ;
        RECT 180.400 481.600 181.200 486.200 ;
        RECT 183.600 481.600 184.400 486.200 ;
        RECT 191.600 481.600 192.400 486.200 ;
        RECT 194.800 481.600 195.600 486.200 ;
        RECT 201.200 481.600 202.000 486.200 ;
        RECT 204.400 481.600 205.200 486.200 ;
        RECT 207.600 481.600 208.400 486.200 ;
        RECT 209.200 481.600 210.000 486.200 ;
        RECT 212.400 481.600 213.200 486.200 ;
        RECT 215.600 481.600 216.400 486.200 ;
        RECT 218.800 481.600 219.600 486.200 ;
        RECT 226.800 481.600 227.600 486.200 ;
        RECT 230.000 481.600 230.800 486.200 ;
        RECT 236.400 481.600 237.200 486.200 ;
        RECT 239.600 481.600 240.400 486.200 ;
        RECT 242.800 481.600 243.600 486.200 ;
        RECT 246.000 481.600 246.800 489.000 ;
        RECT 249.200 481.600 250.000 490.200 ;
        RECT 250.800 481.600 251.600 490.200 ;
        RECT 254.000 481.600 254.800 490.200 ;
        RECT 257.200 481.600 258.000 490.200 ;
        RECT 260.400 481.600 261.200 490.200 ;
        RECT 263.600 481.600 264.400 490.200 ;
        RECT 265.200 481.600 266.000 490.200 ;
        RECT 268.400 481.600 269.200 490.200 ;
        RECT 271.600 481.600 272.400 490.200 ;
        RECT 274.800 481.600 275.600 490.200 ;
        RECT 278.000 481.600 278.800 490.200 ;
        RECT 280.200 481.600 281.000 486.200 ;
        RECT 284.400 481.600 285.200 490.200 ;
        RECT 286.000 481.600 286.800 486.200 ;
        RECT 289.200 481.600 290.000 486.200 ;
        RECT 290.800 481.600 291.600 490.200 ;
        RECT 295.000 481.600 295.800 486.200 ;
        RECT 297.200 481.600 298.000 490.200 ;
        RECT 301.400 481.600 302.200 486.200 ;
        RECT 309.600 481.600 310.400 490.200 ;
        RECT 314.800 481.600 315.600 489.800 ;
        RECT 318.000 481.600 318.800 490.200 ;
        RECT 321.200 481.600 322.000 489.000 ;
        RECT 324.400 481.600 325.200 490.200 ;
        RECT 328.600 481.600 329.400 486.200 ;
        RECT 330.800 481.600 331.600 490.200 ;
        RECT 337.200 481.600 338.000 489.000 ;
        RECT 340.400 481.600 341.200 490.200 ;
        RECT 342.600 481.600 343.400 486.200 ;
        RECT 346.800 481.600 347.600 490.200 ;
        RECT 349.600 481.600 350.400 490.200 ;
        RECT 354.800 481.600 355.600 489.800 ;
        RECT 358.000 481.600 358.800 490.200 ;
        RECT 362.200 481.600 363.000 486.200 ;
        RECT 365.000 481.600 365.800 486.200 ;
        RECT 369.200 481.600 370.000 490.200 ;
        RECT 372.000 481.600 372.800 490.200 ;
        RECT 377.200 481.600 378.000 489.800 ;
        RECT 382.000 481.600 382.800 490.200 ;
        RECT 387.600 481.600 388.400 486.200 ;
        RECT 390.800 481.600 391.600 486.200 ;
        RECT 396.400 481.600 397.200 490.000 ;
        RECT 399.600 481.600 400.400 490.200 ;
        RECT 403.800 481.600 404.600 486.200 ;
        RECT 406.600 481.600 407.400 486.200 ;
        RECT 410.800 481.600 411.600 490.200 ;
        RECT 414.000 481.600 414.800 490.000 ;
        RECT 419.600 481.600 420.400 486.200 ;
        RECT 422.800 481.600 423.600 486.200 ;
        RECT 428.400 481.600 429.200 490.200 ;
        RECT 432.800 481.600 433.600 490.200 ;
        RECT 438.000 481.600 438.800 489.800 ;
        RECT 441.200 481.600 442.000 490.200 ;
        RECT 445.400 481.600 446.200 486.200 ;
        RECT 448.200 481.600 449.000 486.200 ;
        RECT 452.400 481.600 453.200 490.200 ;
        RECT 454.000 481.600 454.800 490.200 ;
        RECT 458.200 481.600 459.000 486.200 ;
        RECT 465.200 481.600 466.000 490.200 ;
        RECT 469.400 481.600 470.200 486.200 ;
        RECT 472.200 481.600 473.000 486.200 ;
        RECT 476.400 481.600 477.200 490.200 ;
        RECT 479.600 481.600 480.400 490.200 ;
        RECT 485.200 481.600 486.000 486.200 ;
        RECT 488.400 481.600 489.200 486.200 ;
        RECT 494.000 481.600 494.800 490.000 ;
        RECT 498.800 481.600 499.600 489.800 ;
        RECT 504.000 481.600 504.800 490.200 ;
        RECT 506.800 481.600 507.600 490.200 ;
        RECT 511.000 481.600 511.800 486.200 ;
        RECT 513.800 481.600 514.600 486.200 ;
        RECT 518.000 481.600 518.800 490.200 ;
        RECT 521.200 481.600 522.000 490.200 ;
        RECT 526.800 481.600 527.600 486.200 ;
        RECT 530.000 481.600 530.800 486.200 ;
        RECT 535.600 481.600 536.400 490.000 ;
        RECT 538.800 481.600 539.600 490.200 ;
        RECT 543.000 481.600 543.800 486.200 ;
        RECT 545.200 481.600 546.000 490.200 ;
        RECT 549.400 481.600 550.200 486.200 ;
        RECT 553.200 481.600 554.000 490.200 ;
        RECT 558.800 481.600 559.600 486.200 ;
        RECT 562.000 481.600 562.800 486.200 ;
        RECT 567.600 481.600 568.400 490.000 ;
        RECT 571.400 481.600 572.200 486.200 ;
        RECT 575.600 481.600 576.400 490.200 ;
        RECT 604.200 490.000 605.200 490.200 ;
        RECT 607.600 489.600 608.400 490.200 ;
        RECT 577.200 481.600 578.000 486.200 ;
        RECT 580.400 481.600 581.200 486.200 ;
        RECT 583.600 481.600 584.400 486.200 ;
        RECT 586.800 481.600 587.600 486.200 ;
        RECT 594.800 481.600 595.600 486.200 ;
        RECT 598.000 481.600 598.800 486.200 ;
        RECT 604.400 481.600 605.200 486.200 ;
        RECT 607.600 481.600 608.400 486.200 ;
        RECT 610.800 481.600 611.600 486.200 ;
        RECT 0.400 480.400 614.000 481.600 ;
        RECT 2.800 472.000 3.600 480.400 ;
        RECT 8.400 475.800 9.200 480.400 ;
        RECT 11.600 475.800 12.400 480.400 ;
        RECT 17.200 471.800 18.000 480.400 ;
        RECT 20.400 471.800 21.200 480.400 ;
        RECT 24.600 475.800 25.400 480.400 ;
        RECT 27.400 475.800 28.200 480.400 ;
        RECT 31.600 471.800 32.400 480.400 ;
        RECT 34.800 472.000 35.600 480.400 ;
        RECT 40.400 475.800 41.200 480.400 ;
        RECT 43.600 475.800 44.400 480.400 ;
        RECT 49.200 471.800 50.000 480.400 ;
        RECT 52.400 471.800 53.200 480.400 ;
        RECT 56.600 475.800 57.400 480.400 ;
        RECT 59.400 475.800 60.200 480.400 ;
        RECT 63.600 471.800 64.400 480.400 ;
        RECT 66.400 471.800 67.200 480.400 ;
        RECT 71.600 472.200 72.400 480.400 ;
        RECT 74.800 475.800 75.600 480.400 ;
        RECT 78.000 475.800 78.800 480.400 ;
        RECT 80.800 471.800 81.600 480.400 ;
        RECT 86.000 472.200 86.800 480.400 ;
        RECT 89.200 471.800 90.000 480.400 ;
        RECT 92.400 473.000 93.200 480.400 ;
        RECT 96.800 471.800 97.600 480.400 ;
        RECT 102.000 472.200 102.800 480.400 ;
        RECT 105.200 471.800 106.000 480.400 ;
        RECT 108.400 473.000 109.200 480.400 ;
        RECT 111.600 475.800 112.400 480.400 ;
        RECT 114.800 475.800 115.600 480.400 ;
        RECT 118.000 476.200 118.800 480.400 ;
        RECT 121.800 475.800 122.600 480.400 ;
        RECT 126.000 471.800 126.800 480.400 ;
        RECT 128.200 475.800 129.000 480.400 ;
        RECT 132.400 471.800 133.200 480.400 ;
        RECT 134.000 471.800 134.800 480.400 ;
        RECT 138.200 475.800 139.000 480.400 ;
        RECT 140.400 471.800 141.200 480.400 ;
        RECT 145.200 471.800 146.000 480.400 ;
        RECT 149.400 475.800 150.200 480.400 ;
        RECT 158.000 473.000 158.800 480.400 ;
        RECT 161.200 471.800 162.000 480.400 ;
        RECT 164.000 471.800 164.800 480.400 ;
        RECT 169.200 472.200 170.000 480.400 ;
        RECT 172.400 471.800 173.200 480.400 ;
        RECT 176.600 475.800 177.400 480.400 ;
        RECT 178.800 471.800 179.600 480.400 ;
        RECT 183.000 475.800 183.800 480.400 ;
        RECT 186.800 471.800 187.600 480.400 ;
        RECT 192.400 475.800 193.200 480.400 ;
        RECT 195.600 475.800 196.400 480.400 ;
        RECT 201.200 472.000 202.000 480.400 ;
        RECT 204.400 475.800 205.200 480.400 ;
        RECT 207.600 475.800 208.400 480.400 ;
        RECT 209.200 471.800 210.000 480.400 ;
        RECT 212.400 471.800 213.200 480.400 ;
        RECT 216.600 475.800 217.400 480.400 ;
        RECT 219.400 475.800 220.200 480.400 ;
        RECT 223.600 471.800 224.400 480.400 ;
        RECT 226.800 473.200 227.800 480.400 ;
        RECT 233.000 479.800 233.800 480.400 ;
        RECT 233.000 473.200 234.000 479.800 ;
        RECT 237.000 475.800 237.800 480.400 ;
        RECT 241.200 471.800 242.000 480.400 ;
        RECT 246.000 471.800 246.800 480.400 ;
        RECT 249.200 473.000 250.000 480.400 ;
        RECT 252.400 471.800 253.200 480.400 ;
        RECT 254.000 475.800 254.800 480.400 ;
        RECT 257.200 475.800 258.000 480.400 ;
        RECT 260.400 475.800 261.200 480.400 ;
        RECT 266.800 475.600 267.600 480.400 ;
        RECT 270.000 475.800 270.800 480.400 ;
        RECT 278.000 475.800 278.800 480.400 ;
        RECT 281.200 475.800 282.000 480.400 ;
        RECT 284.400 475.800 285.200 480.400 ;
        RECT 287.600 475.800 288.400 480.400 ;
        RECT 289.200 475.800 290.000 480.400 ;
        RECT 292.400 475.800 293.200 480.400 ;
        RECT 297.200 471.800 298.000 480.400 ;
        RECT 298.800 471.800 299.600 480.400 ;
        RECT 302.000 473.000 302.800 480.400 ;
        RECT 311.600 472.000 312.400 480.400 ;
        RECT 317.200 475.800 318.000 480.400 ;
        RECT 320.400 475.800 321.200 480.400 ;
        RECT 326.000 471.800 326.800 480.400 ;
        RECT 329.800 475.800 330.600 480.400 ;
        RECT 334.000 471.800 334.800 480.400 ;
        RECT 335.600 471.800 336.400 480.400 ;
        RECT 339.800 475.800 340.600 480.400 ;
        RECT 343.600 475.800 344.400 480.400 ;
        RECT 345.200 471.800 346.000 480.400 ;
        RECT 349.400 475.800 350.200 480.400 ;
        RECT 352.200 475.800 353.000 480.400 ;
        RECT 356.400 471.800 357.200 480.400 ;
        RECT 359.200 471.800 360.000 480.400 ;
        RECT 364.400 472.200 365.200 480.400 ;
        RECT 369.200 472.000 370.000 480.400 ;
        RECT 374.800 475.800 375.600 480.400 ;
        RECT 378.000 475.800 378.800 480.400 ;
        RECT 383.600 471.800 384.400 480.400 ;
        RECT 386.800 471.800 387.600 480.400 ;
        RECT 390.000 473.000 390.800 480.400 ;
        RECT 393.800 475.800 394.600 480.400 ;
        RECT 398.000 471.800 398.800 480.400 ;
        RECT 399.600 475.800 400.400 480.400 ;
        RECT 404.400 472.000 405.200 480.400 ;
        RECT 410.000 475.800 410.800 480.400 ;
        RECT 413.200 475.800 414.000 480.400 ;
        RECT 418.800 471.800 419.600 480.400 ;
        RECT 422.000 475.800 422.800 480.400 ;
        RECT 425.200 475.800 426.000 480.400 ;
        RECT 426.800 475.800 427.600 480.400 ;
        RECT 430.000 475.800 430.800 480.400 ;
        RECT 431.600 471.800 432.400 480.400 ;
        RECT 435.800 475.800 436.600 480.400 ;
        RECT 438.600 475.800 439.400 480.400 ;
        RECT 442.800 471.800 443.600 480.400 ;
        RECT 446.000 472.200 446.800 480.400 ;
        RECT 451.200 471.800 452.000 480.400 ;
        RECT 460.000 471.800 460.800 480.400 ;
        RECT 465.200 472.200 466.000 480.400 ;
        RECT 468.400 475.800 469.200 480.400 ;
        RECT 471.600 475.800 472.400 480.400 ;
        RECT 473.200 471.800 474.000 480.400 ;
        RECT 477.400 475.800 478.200 480.400 ;
        RECT 479.600 471.800 480.400 480.400 ;
        RECT 482.800 473.000 483.600 480.400 ;
        RECT 487.600 472.200 488.400 480.400 ;
        RECT 492.800 471.800 493.600 480.400 ;
        RECT 495.600 475.800 496.400 480.400 ;
        RECT 498.800 471.800 499.600 480.400 ;
        RECT 503.000 475.800 503.800 480.400 ;
        RECT 505.200 475.800 506.000 480.400 ;
        RECT 508.400 475.800 509.200 480.400 ;
        RECT 513.200 471.800 514.000 480.400 ;
        RECT 514.800 471.800 515.600 480.400 ;
        RECT 521.200 472.200 522.000 480.400 ;
        RECT 526.400 471.800 527.200 480.400 ;
        RECT 532.400 471.800 533.200 480.400 ;
        RECT 535.600 475.800 536.400 480.400 ;
        RECT 538.800 473.200 539.800 480.400 ;
        RECT 545.000 479.800 545.800 480.400 ;
        RECT 545.000 473.200 546.000 479.800 ;
        RECT 551.600 471.800 552.400 480.400 ;
        RECT 554.800 475.800 555.600 480.400 ;
        RECT 558.200 479.800 559.000 480.400 ;
        RECT 558.000 473.200 559.000 479.800 ;
        RECT 564.200 473.200 565.200 480.400 ;
        RECT 569.400 479.800 570.200 480.400 ;
        RECT 569.200 473.200 570.200 479.800 ;
        RECT 575.400 473.200 576.400 480.400 ;
        RECT 578.800 475.800 579.600 480.400 ;
        RECT 582.000 475.800 582.800 480.400 ;
        RECT 585.200 475.800 586.000 480.400 ;
        RECT 588.400 475.800 589.200 480.400 ;
        RECT 596.400 475.800 597.200 480.400 ;
        RECT 599.600 475.800 600.400 480.400 ;
        RECT 606.000 475.800 606.800 480.400 ;
        RECT 609.200 475.800 610.000 480.400 ;
        RECT 612.400 475.800 613.200 480.400 ;
        RECT 605.800 471.800 606.600 472.000 ;
        RECT 609.200 471.800 610.000 472.400 ;
        RECT 583.000 471.200 610.000 471.800 ;
        RECT 583.000 471.000 583.800 471.200 ;
        RECT 255.400 470.000 278.800 470.600 ;
        RECT 255.400 469.800 256.200 470.000 ;
        RECT 260.400 469.600 261.200 470.000 ;
        RECT 266.800 469.600 267.600 470.000 ;
        RECT 278.000 469.400 278.800 470.000 ;
        RECT 240.600 450.800 241.400 451.000 ;
        RECT 299.800 450.800 300.600 451.000 ;
        RECT 543.000 450.800 543.800 451.000 ;
        RECT 578.200 450.800 579.000 451.000 ;
        RECT 240.600 450.200 267.600 450.800 ;
        RECT 299.800 450.200 326.800 450.800 ;
        RECT 543.000 450.200 570.000 450.800 ;
        RECT 578.200 450.200 605.200 450.800 ;
        RECT 2.800 441.600 3.600 450.200 ;
        RECT 8.400 441.600 9.200 446.200 ;
        RECT 11.600 441.600 12.400 446.200 ;
        RECT 17.200 441.600 18.000 450.000 ;
        RECT 20.400 441.600 21.200 450.200 ;
        RECT 24.600 441.600 25.400 446.200 ;
        RECT 28.000 441.600 28.800 450.200 ;
        RECT 33.200 441.600 34.000 449.800 ;
        RECT 36.400 441.600 37.200 446.200 ;
        RECT 39.600 441.600 40.400 450.200 ;
        RECT 42.800 441.600 43.600 449.000 ;
        RECT 46.600 441.600 47.400 446.200 ;
        RECT 50.800 441.600 51.600 450.200 ;
        RECT 54.000 441.600 54.800 450.000 ;
        RECT 59.600 441.600 60.400 446.200 ;
        RECT 62.800 441.600 63.600 446.200 ;
        RECT 68.400 441.600 69.200 450.200 ;
        RECT 73.200 441.600 74.000 449.800 ;
        RECT 78.400 441.600 79.200 450.200 ;
        RECT 81.200 441.600 82.000 450.200 ;
        RECT 85.400 441.600 86.200 446.200 ;
        RECT 88.200 441.600 89.000 446.200 ;
        RECT 92.400 441.600 93.200 450.200 ;
        RECT 94.000 441.600 94.800 450.200 ;
        RECT 97.200 441.600 98.000 449.000 ;
        RECT 100.400 441.600 101.200 450.200 ;
        RECT 104.600 441.600 105.400 446.200 ;
        RECT 106.800 441.600 107.600 446.200 ;
        RECT 110.000 441.600 110.800 445.800 ;
        RECT 113.200 441.600 114.000 446.200 ;
        RECT 116.400 441.600 117.200 445.800 ;
        RECT 120.800 441.600 121.600 450.200 ;
        RECT 126.000 441.600 126.800 449.800 ;
        RECT 129.200 441.600 130.000 446.200 ;
        RECT 132.400 441.600 133.200 450.200 ;
        RECT 136.600 441.600 137.400 446.200 ;
        RECT 138.800 441.600 139.600 450.200 ;
        RECT 143.000 441.600 143.800 446.200 ;
        RECT 145.200 441.600 146.000 446.200 ;
        RECT 148.400 441.600 149.200 446.200 ;
        RECT 156.000 441.600 156.800 450.200 ;
        RECT 161.200 441.600 162.000 449.800 ;
        RECT 166.000 441.600 166.800 445.800 ;
        RECT 169.200 441.600 170.000 446.200 ;
        RECT 170.800 441.600 171.600 450.200 ;
        RECT 175.000 441.600 175.800 446.200 ;
        RECT 178.800 441.600 179.600 450.200 ;
        RECT 184.400 441.600 185.200 446.200 ;
        RECT 187.600 441.600 188.400 446.200 ;
        RECT 193.200 441.600 194.000 450.000 ;
        RECT 196.400 441.600 197.200 446.200 ;
        RECT 199.600 441.600 200.400 445.800 ;
        RECT 202.800 441.600 203.600 446.200 ;
        RECT 206.000 441.600 206.800 446.200 ;
        RECT 209.200 441.600 210.000 446.200 ;
        RECT 210.800 441.600 211.600 450.200 ;
        RECT 214.000 441.600 214.800 450.200 ;
        RECT 217.200 441.600 218.000 450.200 ;
        RECT 220.400 441.600 221.200 450.200 ;
        RECT 223.600 441.600 224.400 450.200 ;
        RECT 225.200 441.600 226.000 446.200 ;
        RECT 228.400 441.600 229.200 446.200 ;
        RECT 231.600 441.600 232.400 449.000 ;
        RECT 234.800 441.600 235.600 450.200 ;
        RECT 263.400 450.000 264.200 450.200 ;
        RECT 266.800 449.600 267.600 450.200 ;
        RECT 236.400 441.600 237.200 446.200 ;
        RECT 239.600 441.600 240.400 446.200 ;
        RECT 242.800 441.600 243.600 446.200 ;
        RECT 246.000 441.600 246.800 446.200 ;
        RECT 254.000 441.600 254.800 446.200 ;
        RECT 257.200 441.600 258.000 446.200 ;
        RECT 263.600 441.600 264.400 446.200 ;
        RECT 266.800 441.600 267.600 446.200 ;
        RECT 270.000 441.600 270.800 446.200 ;
        RECT 273.800 441.600 274.600 450.200 ;
        RECT 279.600 441.600 280.400 449.000 ;
        RECT 282.800 441.600 283.600 450.200 ;
        RECT 284.400 441.600 285.200 450.200 ;
        RECT 322.600 450.000 323.400 450.200 ;
        RECT 326.000 449.600 326.800 450.200 ;
        RECT 288.600 441.600 289.400 446.200 ;
        RECT 295.600 441.600 296.400 446.200 ;
        RECT 298.800 441.600 299.600 446.200 ;
        RECT 302.000 441.600 302.800 446.200 ;
        RECT 305.200 441.600 306.000 446.200 ;
        RECT 313.200 441.600 314.000 446.200 ;
        RECT 316.400 441.600 317.200 446.200 ;
        RECT 322.800 441.600 323.600 446.200 ;
        RECT 326.000 441.600 326.800 446.200 ;
        RECT 329.200 441.600 330.000 446.200 ;
        RECT 332.400 441.600 333.200 450.200 ;
        RECT 338.000 441.600 338.800 446.200 ;
        RECT 341.200 441.600 342.000 446.200 ;
        RECT 346.800 441.600 347.600 450.000 ;
        RECT 350.000 441.600 350.800 446.200 ;
        RECT 354.800 441.600 355.600 449.000 ;
        RECT 358.000 441.600 358.800 450.200 ;
        RECT 359.600 441.600 360.400 450.200 ;
        RECT 363.800 441.600 364.600 446.200 ;
        RECT 367.600 441.600 368.400 449.800 ;
        RECT 372.800 441.600 373.600 450.200 ;
        RECT 377.200 441.600 378.000 449.800 ;
        RECT 382.400 441.600 383.200 450.200 ;
        RECT 385.200 441.600 386.000 450.200 ;
        RECT 389.400 441.600 390.200 446.200 ;
        RECT 393.200 441.600 394.000 450.000 ;
        RECT 398.800 441.600 399.600 446.200 ;
        RECT 402.000 441.600 402.800 446.200 ;
        RECT 407.600 441.600 408.400 450.200 ;
        RECT 411.400 441.600 412.200 446.200 ;
        RECT 415.600 441.600 416.400 450.200 ;
        RECT 417.800 441.600 418.600 446.200 ;
        RECT 422.000 441.600 422.800 450.200 ;
        RECT 424.200 441.600 425.000 446.200 ;
        RECT 428.400 441.600 429.200 450.200 ;
        RECT 430.000 441.600 430.800 450.200 ;
        RECT 434.200 441.600 435.000 446.200 ;
        RECT 436.400 441.600 437.200 450.200 ;
        RECT 440.600 441.600 441.400 446.200 ;
        RECT 442.800 441.600 443.600 446.200 ;
        RECT 446.000 441.600 446.800 445.800 ;
        RECT 449.200 441.600 450.000 446.200 ;
        RECT 452.400 441.600 453.200 445.800 ;
        RECT 455.600 441.600 456.400 446.200 ;
        RECT 463.600 441.600 464.400 450.200 ;
        RECT 467.800 441.600 468.600 446.200 ;
        RECT 470.000 441.600 470.800 450.200 ;
        RECT 474.200 441.600 475.000 446.200 ;
        RECT 477.000 441.600 477.800 446.200 ;
        RECT 481.200 441.600 482.000 450.200 ;
        RECT 484.400 441.600 485.200 449.800 ;
        RECT 489.600 441.600 490.400 450.200 ;
        RECT 493.000 441.600 493.800 446.200 ;
        RECT 497.200 441.600 498.000 450.200 ;
        RECT 498.800 441.600 499.600 450.200 ;
        RECT 503.000 441.600 503.800 446.200 ;
        RECT 508.400 441.600 509.200 450.200 ;
        RECT 511.600 441.600 512.400 445.800 ;
        RECT 514.800 441.600 515.600 446.200 ;
        RECT 517.000 441.600 517.800 446.200 ;
        RECT 521.200 441.600 522.000 450.200 ;
        RECT 522.800 441.600 523.600 446.200 ;
        RECT 526.600 441.600 527.400 446.200 ;
        RECT 530.800 441.600 531.600 450.200 ;
        RECT 534.000 441.600 534.800 449.000 ;
        RECT 537.200 441.600 538.000 450.200 ;
        RECT 565.800 450.000 566.600 450.200 ;
        RECT 569.200 449.600 570.000 450.200 ;
        RECT 601.000 450.000 602.000 450.200 ;
        RECT 604.400 449.600 605.200 450.200 ;
        RECT 538.800 441.600 539.600 446.200 ;
        RECT 542.000 441.600 542.800 446.200 ;
        RECT 545.200 441.600 546.000 446.200 ;
        RECT 548.400 441.600 549.200 446.200 ;
        RECT 556.400 441.600 557.200 446.200 ;
        RECT 559.600 441.600 560.400 446.200 ;
        RECT 566.000 441.600 566.800 446.200 ;
        RECT 569.200 441.600 570.000 446.200 ;
        RECT 572.400 441.600 573.200 446.200 ;
        RECT 574.000 441.600 574.800 446.200 ;
        RECT 577.200 441.600 578.000 446.200 ;
        RECT 580.400 441.600 581.200 446.200 ;
        RECT 583.600 441.600 584.400 446.200 ;
        RECT 591.600 441.600 592.400 446.200 ;
        RECT 594.800 441.600 595.600 446.200 ;
        RECT 601.200 441.600 602.000 446.200 ;
        RECT 604.400 441.600 605.200 446.200 ;
        RECT 607.600 441.600 608.400 446.200 ;
        RECT 0.400 440.400 614.000 441.600 ;
        RECT 1.200 435.800 2.000 440.400 ;
        RECT 4.400 431.800 5.200 440.400 ;
        RECT 8.600 435.800 9.400 440.400 ;
        RECT 10.800 431.800 11.600 440.400 ;
        RECT 14.000 431.800 14.800 440.400 ;
        RECT 17.200 431.800 18.000 440.400 ;
        RECT 20.400 431.800 21.200 440.400 ;
        RECT 23.600 431.800 24.400 440.400 ;
        RECT 25.800 435.800 26.600 440.400 ;
        RECT 30.000 431.800 30.800 440.400 ;
        RECT 34.200 431.800 35.000 440.400 ;
        RECT 38.000 431.800 38.800 440.400 ;
        RECT 41.200 431.800 42.000 440.400 ;
        RECT 44.400 431.800 45.200 440.400 ;
        RECT 47.600 431.800 48.400 440.400 ;
        RECT 50.800 431.800 51.600 440.400 ;
        RECT 54.000 432.000 54.800 440.400 ;
        RECT 59.600 435.800 60.400 440.400 ;
        RECT 62.800 435.800 63.600 440.400 ;
        RECT 68.400 431.800 69.200 440.400 ;
        RECT 73.200 432.200 74.000 440.400 ;
        RECT 78.400 431.800 79.200 440.400 ;
        RECT 81.200 431.800 82.000 440.400 ;
        RECT 85.400 435.800 86.200 440.400 ;
        RECT 88.200 435.800 89.000 440.400 ;
        RECT 92.400 431.800 93.200 440.400 ;
        RECT 94.000 435.800 94.800 440.400 ;
        RECT 97.200 435.800 98.000 440.400 ;
        RECT 100.400 432.200 101.200 440.400 ;
        RECT 105.600 431.800 106.400 440.400 ;
        RECT 108.400 431.800 109.200 440.400 ;
        RECT 112.600 435.800 113.400 440.400 ;
        RECT 115.400 435.800 116.200 440.400 ;
        RECT 119.600 431.800 120.400 440.400 ;
        RECT 121.200 435.800 122.000 440.400 ;
        RECT 124.400 431.800 125.200 440.400 ;
        RECT 128.600 435.800 129.400 440.400 ;
        RECT 130.800 435.800 131.600 440.400 ;
        RECT 135.600 431.800 136.400 440.400 ;
        RECT 141.200 435.800 142.000 440.400 ;
        RECT 144.400 435.800 145.200 440.400 ;
        RECT 150.000 432.000 150.800 440.400 ;
        RECT 158.000 431.800 158.800 440.400 ;
        RECT 162.200 435.800 163.000 440.400 ;
        RECT 165.000 435.800 165.800 440.400 ;
        RECT 169.200 431.800 170.000 440.400 ;
        RECT 170.800 431.800 171.600 440.400 ;
        RECT 175.000 435.800 175.800 440.400 ;
        RECT 177.800 435.800 178.600 440.400 ;
        RECT 182.000 431.800 182.800 440.400 ;
        RECT 185.200 431.800 186.000 440.400 ;
        RECT 190.800 435.800 191.600 440.400 ;
        RECT 194.000 435.800 194.800 440.400 ;
        RECT 199.600 432.000 200.400 440.400 ;
        RECT 202.800 431.800 203.600 440.400 ;
        RECT 207.000 435.800 207.800 440.400 ;
        RECT 209.200 431.800 210.000 440.400 ;
        RECT 213.400 435.800 214.200 440.400 ;
        RECT 215.600 435.800 216.400 440.400 ;
        RECT 218.800 435.800 219.600 440.400 ;
        RECT 221.000 435.800 221.800 440.400 ;
        RECT 225.200 431.800 226.000 440.400 ;
        RECT 228.400 432.200 229.200 440.400 ;
        RECT 231.600 435.800 232.400 440.400 ;
        RECT 233.200 435.800 234.000 440.400 ;
        RECT 236.400 435.800 237.200 440.400 ;
        RECT 238.000 435.800 238.800 440.400 ;
        RECT 241.200 435.800 242.000 440.400 ;
        RECT 243.400 435.800 244.200 440.400 ;
        RECT 247.600 431.800 248.400 440.400 ;
        RECT 250.800 435.800 251.600 440.400 ;
        RECT 253.000 435.800 253.800 440.400 ;
        RECT 257.200 431.800 258.000 440.400 ;
        RECT 260.400 432.200 261.200 440.400 ;
        RECT 265.600 431.800 266.400 440.400 ;
        RECT 270.000 432.200 270.800 440.400 ;
        RECT 275.200 431.800 276.000 440.400 ;
        RECT 278.000 435.800 278.800 440.400 ;
        RECT 281.200 435.800 282.000 440.400 ;
        RECT 282.800 435.800 283.600 440.400 ;
        RECT 286.000 435.800 286.800 440.400 ;
        RECT 289.200 435.800 290.000 440.400 ;
        RECT 292.400 435.800 293.200 440.400 ;
        RECT 295.600 435.800 296.400 440.400 ;
        RECT 303.600 435.800 304.400 440.400 ;
        RECT 306.800 435.800 307.600 440.400 ;
        RECT 313.200 435.800 314.000 440.400 ;
        RECT 316.400 435.800 317.200 440.400 ;
        RECT 319.600 435.800 320.400 440.400 ;
        RECT 326.000 435.800 326.800 440.400 ;
        RECT 313.000 431.800 313.800 432.000 ;
        RECT 316.400 431.800 317.200 432.400 ;
        RECT 330.800 432.000 331.600 440.400 ;
        RECT 336.400 435.800 337.200 440.400 ;
        RECT 339.600 435.800 340.400 440.400 ;
        RECT 345.200 431.800 346.000 440.400 ;
        RECT 350.000 432.200 350.800 440.400 ;
        RECT 355.200 431.800 356.000 440.400 ;
        RECT 358.000 431.800 358.800 440.400 ;
        RECT 362.200 435.800 363.000 440.400 ;
        RECT 365.000 435.800 365.800 440.400 ;
        RECT 369.200 431.800 370.000 440.400 ;
        RECT 372.000 431.800 372.800 440.400 ;
        RECT 377.200 432.200 378.000 440.400 ;
        RECT 380.400 431.800 381.200 440.400 ;
        RECT 384.600 435.800 385.400 440.400 ;
        RECT 388.000 431.800 388.800 440.400 ;
        RECT 393.200 432.200 394.000 440.400 ;
        RECT 396.400 435.800 397.200 440.400 ;
        RECT 400.800 431.800 401.600 440.400 ;
        RECT 406.000 432.200 406.800 440.400 ;
        RECT 409.200 431.800 410.000 440.400 ;
        RECT 413.400 435.800 414.200 440.400 ;
        RECT 417.200 431.800 418.000 440.400 ;
        RECT 422.800 435.800 423.600 440.400 ;
        RECT 426.000 435.800 426.800 440.400 ;
        RECT 431.600 432.000 432.400 440.400 ;
        RECT 434.800 435.800 435.600 440.400 ;
        RECT 438.000 431.800 438.800 440.400 ;
        RECT 442.200 435.800 443.000 440.400 ;
        RECT 446.000 432.000 446.800 440.400 ;
        RECT 451.600 435.800 452.400 440.400 ;
        RECT 454.800 435.800 455.600 440.400 ;
        RECT 460.400 431.800 461.200 440.400 ;
        RECT 470.000 436.200 470.800 440.400 ;
        RECT 473.200 435.800 474.000 440.400 ;
        RECT 474.800 435.800 475.600 440.400 ;
        RECT 478.000 435.800 478.800 440.400 ;
        RECT 481.200 435.800 482.000 440.400 ;
        RECT 484.400 435.800 485.200 440.400 ;
        RECT 492.400 435.800 493.200 440.400 ;
        RECT 495.600 435.800 496.400 440.400 ;
        RECT 502.000 435.800 502.800 440.400 ;
        RECT 505.200 435.800 506.000 440.400 ;
        RECT 508.400 435.800 509.200 440.400 ;
        RECT 510.000 435.800 510.800 440.400 ;
        RECT 513.200 435.800 514.000 440.400 ;
        RECT 516.400 435.800 517.200 440.400 ;
        RECT 519.600 435.800 520.400 440.400 ;
        RECT 527.600 435.800 528.400 440.400 ;
        RECT 530.800 435.800 531.600 440.400 ;
        RECT 537.200 435.800 538.000 440.400 ;
        RECT 540.400 435.800 541.200 440.400 ;
        RECT 543.600 435.800 544.400 440.400 ;
        RECT 501.800 431.800 502.800 432.000 ;
        RECT 505.200 431.800 506.000 432.400 ;
        RECT 537.000 431.800 537.800 432.000 ;
        RECT 540.400 431.800 541.200 432.400 ;
        RECT 546.800 432.200 547.600 440.400 ;
        RECT 552.000 431.800 552.800 440.400 ;
        RECT 556.400 432.200 557.200 440.400 ;
        RECT 561.600 431.800 562.400 440.400 ;
        RECT 564.400 435.800 565.200 440.400 ;
        RECT 567.600 435.800 568.400 440.400 ;
        RECT 570.800 435.800 571.600 440.400 ;
        RECT 574.000 435.800 574.800 440.400 ;
        RECT 582.000 435.800 582.800 440.400 ;
        RECT 585.200 435.800 586.000 440.400 ;
        RECT 591.600 435.800 592.400 440.400 ;
        RECT 594.800 435.800 595.600 440.400 ;
        RECT 598.000 435.800 598.800 440.400 ;
        RECT 591.400 431.800 592.200 432.000 ;
        RECT 594.800 431.800 595.600 432.400 ;
        RECT 599.600 431.800 600.400 440.400 ;
        RECT 602.800 431.800 603.600 440.400 ;
        RECT 606.000 431.800 606.800 440.400 ;
        RECT 609.200 431.800 610.000 440.400 ;
        RECT 612.400 431.800 613.200 440.400 ;
        RECT 290.200 431.200 317.200 431.800 ;
        RECT 479.000 431.200 506.000 431.800 ;
        RECT 514.200 431.200 541.200 431.800 ;
        RECT 568.600 431.200 595.600 431.800 ;
        RECT 290.200 431.000 291.000 431.200 ;
        RECT 479.000 431.000 479.800 431.200 ;
        RECT 514.200 431.000 515.000 431.200 ;
        RECT 568.600 431.000 569.400 431.200 ;
        RECT 30.600 410.800 31.400 411.000 ;
        RECT 211.400 410.800 212.200 411.000 ;
        RECT 329.800 410.800 330.600 411.000 ;
        RECT 605.000 410.800 605.800 411.000 ;
        RECT 4.400 410.200 31.400 410.800 ;
        RECT 185.200 410.200 212.200 410.800 ;
        RECT 303.600 410.200 330.600 410.800 ;
        RECT 578.800 410.200 605.800 410.800 ;
        RECT 4.400 409.600 5.200 410.200 ;
        RECT 7.800 410.000 8.600 410.200 ;
        RECT 1.200 401.600 2.000 406.200 ;
        RECT 4.400 401.600 5.200 406.200 ;
        RECT 7.600 401.600 8.400 406.200 ;
        RECT 14.000 401.600 14.800 406.200 ;
        RECT 17.200 401.600 18.000 406.200 ;
        RECT 25.200 401.600 26.000 406.200 ;
        RECT 28.400 401.600 29.200 406.200 ;
        RECT 31.600 401.600 32.400 406.200 ;
        RECT 34.800 401.600 35.600 406.200 ;
        RECT 37.000 401.600 37.800 406.200 ;
        RECT 41.200 401.600 42.000 410.200 ;
        RECT 42.800 401.600 43.600 410.200 ;
        RECT 47.000 401.600 47.800 406.200 ;
        RECT 50.800 401.600 51.600 409.800 ;
        RECT 56.000 401.600 56.800 410.200 ;
        RECT 59.400 401.600 60.200 406.200 ;
        RECT 63.600 401.600 64.400 410.200 ;
        RECT 66.800 401.600 67.600 410.000 ;
        RECT 72.400 401.600 73.200 406.200 ;
        RECT 75.600 401.600 76.400 406.200 ;
        RECT 81.200 401.600 82.000 410.200 ;
        RECT 84.400 401.600 85.200 410.200 ;
        RECT 88.600 401.600 89.400 406.200 ;
        RECT 91.400 401.600 92.200 406.200 ;
        RECT 95.600 401.600 96.400 410.200 ;
        RECT 97.200 401.600 98.000 406.200 ;
        RECT 100.400 401.600 101.200 406.200 ;
        RECT 102.000 401.600 102.800 410.200 ;
        RECT 106.200 401.600 107.000 406.200 ;
        RECT 108.400 401.600 109.200 410.200 ;
        RECT 111.600 401.600 112.400 409.000 ;
        RECT 114.800 401.600 115.600 410.200 ;
        RECT 118.000 401.600 118.800 409.000 ;
        RECT 122.800 401.600 123.600 409.000 ;
        RECT 126.000 401.600 126.800 410.200 ;
        RECT 127.600 401.600 128.400 406.200 ;
        RECT 130.800 401.600 131.600 410.200 ;
        RECT 135.000 401.600 135.800 406.200 ;
        RECT 138.800 401.600 139.600 409.800 ;
        RECT 144.000 401.600 144.800 410.200 ;
        RECT 146.800 401.600 147.600 406.200 ;
        RECT 150.000 401.600 150.800 406.200 ;
        RECT 156.400 401.600 157.200 410.200 ;
        RECT 160.600 401.600 161.400 406.200 ;
        RECT 162.800 401.600 163.600 410.200 ;
        RECT 167.000 401.600 167.800 406.200 ;
        RECT 170.800 401.600 171.600 409.000 ;
        RECT 174.000 401.600 174.800 410.200 ;
        RECT 175.600 401.600 176.400 410.200 ;
        RECT 185.200 409.600 186.000 410.200 ;
        RECT 188.400 410.000 189.400 410.200 ;
        RECT 179.800 401.600 180.600 406.200 ;
        RECT 182.000 401.600 182.800 406.200 ;
        RECT 185.200 401.600 186.000 406.200 ;
        RECT 188.400 401.600 189.200 406.200 ;
        RECT 194.800 401.600 195.600 406.200 ;
        RECT 198.000 401.600 198.800 406.200 ;
        RECT 206.000 401.600 206.800 406.200 ;
        RECT 209.200 401.600 210.000 406.200 ;
        RECT 212.400 401.600 213.200 406.200 ;
        RECT 215.600 401.600 216.400 406.200 ;
        RECT 217.200 401.600 218.000 406.200 ;
        RECT 220.400 401.600 221.200 410.200 ;
        RECT 228.400 401.600 229.200 409.000 ;
        RECT 233.200 401.600 234.000 405.800 ;
        RECT 236.400 401.600 237.200 406.200 ;
        RECT 240.600 401.600 241.400 410.200 ;
        RECT 247.600 401.600 248.400 410.200 ;
        RECT 250.800 402.200 251.800 408.800 ;
        RECT 251.000 401.600 251.800 402.200 ;
        RECT 257.000 401.600 258.000 408.800 ;
        RECT 261.000 401.600 261.800 406.200 ;
        RECT 265.200 401.600 266.000 410.200 ;
        RECT 268.400 402.200 269.400 408.800 ;
        RECT 268.600 401.600 269.400 402.200 ;
        RECT 274.600 401.600 275.600 408.800 ;
        RECT 278.000 401.600 278.800 410.200 ;
        RECT 282.200 401.600 283.000 406.200 ;
        RECT 284.400 401.600 285.200 410.200 ;
        RECT 303.600 409.600 304.400 410.200 ;
        RECT 306.800 410.000 307.800 410.200 ;
        RECT 288.600 401.600 289.400 406.200 ;
        RECT 290.800 401.600 291.600 406.200 ;
        RECT 294.000 401.600 294.800 406.200 ;
        RECT 300.400 401.600 301.200 406.200 ;
        RECT 303.600 401.600 304.400 406.200 ;
        RECT 306.800 401.600 307.600 406.200 ;
        RECT 313.200 401.600 314.000 406.200 ;
        RECT 316.400 401.600 317.200 406.200 ;
        RECT 324.400 401.600 325.200 406.200 ;
        RECT 327.600 401.600 328.400 406.200 ;
        RECT 330.800 401.600 331.600 406.200 ;
        RECT 334.000 401.600 334.800 406.200 ;
        RECT 337.200 401.600 338.000 410.000 ;
        RECT 342.800 401.600 343.600 406.200 ;
        RECT 346.000 401.600 346.800 406.200 ;
        RECT 351.600 401.600 352.400 410.200 ;
        RECT 354.800 401.600 355.600 410.200 ;
        RECT 359.000 401.600 359.800 406.200 ;
        RECT 361.800 401.600 362.600 406.200 ;
        RECT 366.000 401.600 366.800 410.200 ;
        RECT 367.600 401.600 368.400 406.200 ;
        RECT 370.800 401.600 371.600 410.200 ;
        RECT 375.000 401.600 375.800 406.200 ;
        RECT 377.800 401.600 378.600 406.200 ;
        RECT 382.000 401.600 382.800 410.200 ;
        RECT 383.600 401.600 384.400 406.200 ;
        RECT 386.800 401.600 387.600 410.200 ;
        RECT 391.000 401.600 391.800 406.200 ;
        RECT 393.200 401.600 394.000 406.200 ;
        RECT 396.400 401.600 397.200 405.800 ;
        RECT 399.600 401.600 400.400 406.200 ;
        RECT 402.800 401.600 403.600 405.800 ;
        RECT 406.000 401.600 406.800 410.200 ;
        RECT 410.200 401.600 411.000 406.200 ;
        RECT 412.400 401.600 413.200 406.200 ;
        RECT 415.600 401.600 416.400 410.200 ;
        RECT 419.800 401.600 420.600 406.200 ;
        RECT 422.000 401.600 422.800 410.200 ;
        RECT 426.200 401.600 427.000 406.200 ;
        RECT 428.400 401.600 429.200 410.200 ;
        RECT 432.600 401.600 433.400 406.200 ;
        RECT 434.800 401.600 435.600 406.200 ;
        RECT 438.000 401.600 438.800 406.200 ;
        RECT 441.200 401.600 442.000 406.200 ;
        RECT 442.800 401.600 443.600 410.200 ;
        RECT 447.000 401.600 447.800 406.200 ;
        RECT 449.200 401.600 450.000 406.200 ;
        RECT 452.400 401.600 453.200 406.200 ;
        RECT 454.000 401.600 454.800 410.200 ;
        RECT 462.600 401.600 463.400 406.200 ;
        RECT 466.800 401.600 467.600 410.200 ;
        RECT 469.000 401.600 469.800 406.200 ;
        RECT 473.200 401.600 474.000 410.200 ;
        RECT 476.400 401.600 477.400 408.800 ;
        RECT 482.600 402.200 483.600 408.800 ;
        RECT 482.600 401.600 483.400 402.200 ;
        RECT 486.600 401.600 487.400 406.200 ;
        RECT 490.800 401.600 491.600 410.200 ;
        RECT 494.000 401.600 494.800 409.800 ;
        RECT 497.200 401.600 498.000 406.200 ;
        RECT 502.000 401.600 502.800 409.000 ;
        RECT 505.200 401.600 506.000 406.200 ;
        RECT 508.400 401.600 509.200 406.200 ;
        RECT 510.000 401.600 510.800 406.200 ;
        RECT 513.200 401.600 514.000 406.200 ;
        RECT 514.800 401.600 515.600 406.200 ;
        RECT 518.000 401.600 518.800 405.800 ;
        RECT 521.200 401.600 522.000 406.200 ;
        RECT 524.400 401.600 525.200 410.200 ;
        RECT 531.400 401.600 532.200 410.200 ;
        RECT 537.200 402.200 538.200 408.800 ;
        RECT 537.400 401.600 538.200 402.200 ;
        RECT 543.400 401.600 544.400 408.800 ;
        RECT 546.800 401.600 547.600 410.200 ;
        RECT 551.000 401.600 551.800 406.200 ;
        RECT 553.200 401.600 554.000 410.200 ;
        RECT 578.800 409.600 579.600 410.200 ;
        RECT 582.000 410.000 583.000 410.200 ;
        RECT 557.400 401.600 558.200 406.200 ;
        RECT 561.200 402.200 562.200 408.800 ;
        RECT 561.400 401.600 562.200 402.200 ;
        RECT 567.400 401.600 568.400 408.800 ;
        RECT 570.800 401.600 571.600 406.200 ;
        RECT 574.000 401.600 574.800 406.200 ;
        RECT 575.600 401.600 576.400 406.200 ;
        RECT 578.800 401.600 579.600 406.200 ;
        RECT 582.000 401.600 582.800 406.200 ;
        RECT 588.400 401.600 589.200 406.200 ;
        RECT 591.600 401.600 592.400 406.200 ;
        RECT 599.600 401.600 600.400 406.200 ;
        RECT 602.800 401.600 603.600 406.200 ;
        RECT 606.000 401.600 606.800 406.200 ;
        RECT 609.200 401.600 610.000 406.200 ;
        RECT 0.400 400.400 614.000 401.600 ;
        RECT 1.200 395.800 2.000 400.400 ;
        RECT 4.400 395.800 5.200 400.400 ;
        RECT 7.600 395.800 8.400 400.400 ;
        RECT 14.000 395.800 14.800 400.400 ;
        RECT 17.200 395.800 18.000 400.400 ;
        RECT 25.200 395.800 26.000 400.400 ;
        RECT 28.400 395.800 29.200 400.400 ;
        RECT 31.600 395.800 32.400 400.400 ;
        RECT 34.800 395.800 35.600 400.400 ;
        RECT 36.400 395.800 37.200 400.400 ;
        RECT 39.600 395.800 40.400 400.400 ;
        RECT 4.400 391.800 5.200 392.400 ;
        RECT 7.800 391.800 8.600 392.000 ;
        RECT 41.200 391.800 42.000 400.400 ;
        RECT 44.400 393.000 45.200 400.400 ;
        RECT 49.200 392.000 50.000 400.400 ;
        RECT 54.800 395.800 55.600 400.400 ;
        RECT 58.000 395.800 58.800 400.400 ;
        RECT 63.600 391.800 64.400 400.400 ;
        RECT 68.400 393.000 69.200 400.400 ;
        RECT 71.600 391.800 72.400 400.400 ;
        RECT 73.800 395.800 74.600 400.400 ;
        RECT 78.000 391.800 78.800 400.400 ;
        RECT 80.800 391.800 81.600 400.400 ;
        RECT 86.000 392.200 86.800 400.400 ;
        RECT 90.400 391.800 91.200 400.400 ;
        RECT 95.600 392.200 96.400 400.400 ;
        RECT 100.400 395.800 101.200 400.400 ;
        RECT 102.000 391.800 102.800 400.400 ;
        RECT 105.200 393.000 106.000 400.400 ;
        RECT 111.600 391.800 112.400 400.400 ;
        RECT 114.800 392.000 115.600 400.400 ;
        RECT 120.400 395.800 121.200 400.400 ;
        RECT 123.600 395.800 124.400 400.400 ;
        RECT 129.200 391.800 130.000 400.400 ;
        RECT 132.400 391.800 133.200 400.400 ;
        RECT 136.600 395.800 137.400 400.400 ;
        RECT 139.400 395.800 140.200 400.400 ;
        RECT 143.600 391.800 144.400 400.400 ;
        RECT 145.200 391.800 146.000 400.400 ;
        RECT 148.400 393.000 149.200 400.400 ;
        RECT 156.400 395.800 157.200 400.400 ;
        RECT 159.600 391.800 160.400 400.400 ;
        RECT 162.800 393.000 163.600 400.400 ;
        RECT 166.000 395.800 166.800 400.400 ;
        RECT 169.200 395.800 170.000 400.400 ;
        RECT 172.400 395.800 173.200 400.400 ;
        RECT 175.600 395.800 176.400 400.400 ;
        RECT 183.600 395.800 184.400 400.400 ;
        RECT 186.800 395.800 187.600 400.400 ;
        RECT 193.200 395.800 194.000 400.400 ;
        RECT 196.400 395.800 197.200 400.400 ;
        RECT 199.600 395.800 200.400 400.400 ;
        RECT 201.200 395.800 202.000 400.400 ;
        RECT 204.400 395.800 205.200 400.400 ;
        RECT 207.600 395.800 208.400 400.400 ;
        RECT 209.200 395.800 210.000 400.400 ;
        RECT 212.400 395.800 213.200 400.400 ;
        RECT 214.000 395.800 214.800 400.400 ;
        RECT 217.200 395.800 218.000 400.400 ;
        RECT 220.400 395.800 221.200 400.400 ;
        RECT 226.800 395.800 227.600 400.400 ;
        RECT 230.000 395.800 230.800 400.400 ;
        RECT 238.000 395.800 238.800 400.400 ;
        RECT 241.200 395.800 242.000 400.400 ;
        RECT 244.400 395.800 245.200 400.400 ;
        RECT 247.600 395.800 248.400 400.400 ;
        RECT 249.200 395.800 250.000 400.400 ;
        RECT 252.400 395.800 253.200 400.400 ;
        RECT 254.600 395.800 255.400 400.400 ;
        RECT 193.000 391.800 193.800 392.000 ;
        RECT 196.400 391.800 197.200 392.400 ;
        RECT 4.400 391.200 31.400 391.800 ;
        RECT 30.600 391.000 31.400 391.200 ;
        RECT 170.200 391.200 197.200 391.800 ;
        RECT 217.200 391.800 218.000 392.400 ;
        RECT 220.400 391.800 221.400 392.000 ;
        RECT 258.800 391.800 259.600 400.400 ;
        RECT 262.000 393.000 262.800 400.400 ;
        RECT 265.200 395.800 266.000 400.400 ;
        RECT 268.400 395.800 269.200 400.400 ;
        RECT 271.600 395.800 272.400 400.400 ;
        RECT 278.000 395.800 278.800 400.400 ;
        RECT 281.200 395.800 282.000 400.400 ;
        RECT 289.200 395.800 290.000 400.400 ;
        RECT 292.400 395.800 293.200 400.400 ;
        RECT 295.600 395.800 296.400 400.400 ;
        RECT 298.800 395.800 299.600 400.400 ;
        RECT 305.200 395.800 306.000 400.400 ;
        RECT 308.400 395.800 309.200 400.400 ;
        RECT 311.600 395.800 312.400 400.400 ;
        RECT 318.000 395.800 318.800 400.400 ;
        RECT 321.200 395.800 322.000 400.400 ;
        RECT 329.200 395.800 330.000 400.400 ;
        RECT 332.400 395.800 333.200 400.400 ;
        RECT 335.600 395.800 336.400 400.400 ;
        RECT 338.800 395.800 339.600 400.400 ;
        RECT 340.400 395.800 341.200 400.400 ;
        RECT 343.600 395.800 344.400 400.400 ;
        RECT 346.800 395.800 347.600 400.400 ;
        RECT 350.000 395.800 350.800 400.400 ;
        RECT 358.000 395.800 358.800 400.400 ;
        RECT 361.200 395.800 362.000 400.400 ;
        RECT 367.600 395.800 368.400 400.400 ;
        RECT 370.800 395.800 371.600 400.400 ;
        RECT 374.000 395.800 374.800 400.400 ;
        RECT 268.400 391.800 269.200 392.400 ;
        RECT 271.800 391.800 272.600 392.000 ;
        RECT 308.400 391.800 309.200 392.400 ;
        RECT 311.800 391.800 312.600 392.000 ;
        RECT 367.400 391.800 368.200 392.000 ;
        RECT 370.800 391.800 371.600 392.400 ;
        RECT 377.200 392.000 378.000 400.400 ;
        RECT 382.800 395.800 383.600 400.400 ;
        RECT 386.000 395.800 386.800 400.400 ;
        RECT 391.600 391.800 392.400 400.400 ;
        RECT 394.800 395.800 395.600 400.400 ;
        RECT 398.000 395.800 398.800 400.400 ;
        RECT 402.800 393.000 403.600 400.400 ;
        RECT 406.000 391.800 406.800 400.400 ;
        RECT 407.600 395.800 408.400 400.400 ;
        RECT 410.800 395.800 411.600 400.400 ;
        RECT 414.000 395.800 414.800 400.400 ;
        RECT 417.200 395.800 418.000 400.400 ;
        RECT 425.200 395.800 426.000 400.400 ;
        RECT 428.400 395.800 429.200 400.400 ;
        RECT 434.800 395.800 435.600 400.400 ;
        RECT 438.000 395.800 438.800 400.400 ;
        RECT 441.200 395.800 442.000 400.400 ;
        RECT 442.800 395.800 443.600 400.400 ;
        RECT 446.000 395.800 446.800 400.400 ;
        RECT 448.200 395.800 449.000 400.400 ;
        RECT 434.600 391.800 435.400 392.000 ;
        RECT 438.000 391.800 438.800 392.400 ;
        RECT 452.400 391.800 453.200 400.400 ;
        RECT 458.800 395.800 459.600 400.400 ;
        RECT 462.000 395.800 462.800 400.400 ;
        RECT 465.200 395.800 466.000 400.400 ;
        RECT 471.600 395.800 472.400 400.400 ;
        RECT 474.800 395.800 475.600 400.400 ;
        RECT 482.800 395.800 483.600 400.400 ;
        RECT 486.000 395.800 486.800 400.400 ;
        RECT 489.200 395.800 490.000 400.400 ;
        RECT 492.400 395.800 493.200 400.400 ;
        RECT 462.000 391.800 462.800 392.400 ;
        RECT 465.400 391.800 466.200 392.000 ;
        RECT 494.000 391.800 494.800 400.400 ;
        RECT 497.200 391.800 498.000 400.400 ;
        RECT 500.400 391.800 501.200 400.400 ;
        RECT 503.600 391.800 504.400 400.400 ;
        RECT 506.800 391.800 507.600 400.400 ;
        RECT 511.600 391.800 512.400 400.400 ;
        RECT 513.200 395.800 514.000 400.400 ;
        RECT 516.400 395.800 517.200 400.400 ;
        RECT 518.000 395.800 518.800 400.400 ;
        RECT 521.200 395.800 522.000 400.400 ;
        RECT 524.400 395.800 525.200 400.400 ;
        RECT 530.800 395.800 531.600 400.400 ;
        RECT 534.000 395.800 534.800 400.400 ;
        RECT 542.000 395.800 542.800 400.400 ;
        RECT 545.200 395.800 546.000 400.400 ;
        RECT 548.400 395.800 549.200 400.400 ;
        RECT 551.600 395.800 552.400 400.400 ;
        RECT 521.200 391.800 522.000 392.400 ;
        RECT 524.600 391.800 525.400 392.000 ;
        RECT 556.400 391.800 557.200 400.400 ;
        RECT 558.600 395.800 559.400 400.400 ;
        RECT 562.800 391.800 563.600 400.400 ;
        RECT 566.000 395.800 566.800 400.400 ;
        RECT 569.800 391.800 570.600 400.400 ;
        RECT 574.000 395.800 574.800 400.400 ;
        RECT 577.200 395.800 578.000 400.400 ;
        RECT 580.400 395.800 581.200 400.400 ;
        RECT 586.800 395.800 587.600 400.400 ;
        RECT 590.000 395.800 590.800 400.400 ;
        RECT 598.000 395.800 598.800 400.400 ;
        RECT 601.200 395.800 602.000 400.400 ;
        RECT 604.400 395.800 605.200 400.400 ;
        RECT 607.600 395.800 608.400 400.400 ;
        RECT 577.200 391.800 578.000 392.400 ;
        RECT 580.600 391.800 581.400 392.000 ;
        RECT 217.200 391.200 244.200 391.800 ;
        RECT 268.400 391.200 295.400 391.800 ;
        RECT 308.400 391.200 335.400 391.800 ;
        RECT 170.200 391.000 171.000 391.200 ;
        RECT 243.400 391.000 244.200 391.200 ;
        RECT 294.600 391.000 295.400 391.200 ;
        RECT 334.600 391.000 335.400 391.200 ;
        RECT 344.600 391.200 371.600 391.800 ;
        RECT 411.800 391.200 438.800 391.800 ;
        RECT 462.000 391.200 489.000 391.800 ;
        RECT 521.200 391.200 548.200 391.800 ;
        RECT 577.200 391.200 604.200 391.800 ;
        RECT 344.600 391.000 345.400 391.200 ;
        RECT 411.800 391.000 412.600 391.200 ;
        RECT 488.200 391.000 489.000 391.200 ;
        RECT 547.400 391.000 548.200 391.200 ;
        RECT 603.400 391.000 604.200 391.200 ;
        RECT 529.200 372.000 530.000 372.600 ;
        RECT 546.800 372.000 547.600 372.400 ;
        RECT 551.800 372.000 552.600 372.200 ;
        RECT 529.200 371.400 552.600 372.000 ;
        RECT 203.400 370.800 204.200 371.000 ;
        RECT 177.200 370.200 204.200 370.800 ;
        RECT 237.400 370.800 238.200 371.000 ;
        RECT 373.000 370.800 373.800 371.000 ;
        RECT 237.400 370.200 264.400 370.800 ;
        RECT 346.800 370.200 373.800 370.800 ;
        RECT 383.000 370.800 383.800 371.000 ;
        RECT 451.800 370.800 452.600 371.000 ;
        RECT 576.600 370.800 577.400 371.000 ;
        RECT 383.000 370.200 410.000 370.800 ;
        RECT 451.800 370.200 478.800 370.800 ;
        RECT 576.600 370.200 603.600 370.800 ;
        RECT 1.200 361.600 2.000 366.200 ;
        RECT 4.400 361.600 5.200 366.200 ;
        RECT 7.600 361.600 8.400 370.200 ;
        RECT 11.800 361.600 12.600 366.200 ;
        RECT 14.000 361.600 14.800 370.200 ;
        RECT 18.200 361.600 19.000 366.200 ;
        RECT 21.000 361.600 21.800 366.200 ;
        RECT 25.200 361.600 26.000 370.200 ;
        RECT 26.800 361.600 27.600 370.200 ;
        RECT 31.000 361.600 31.800 366.200 ;
        RECT 33.800 361.600 34.600 366.200 ;
        RECT 38.000 361.600 38.800 370.200 ;
        RECT 40.200 361.600 41.000 366.200 ;
        RECT 44.400 361.600 45.200 370.200 ;
        RECT 46.000 361.600 46.800 366.200 ;
        RECT 49.200 361.600 50.000 366.200 ;
        RECT 51.400 361.600 52.200 366.200 ;
        RECT 55.600 361.600 56.400 370.200 ;
        RECT 58.800 361.600 59.600 369.800 ;
        RECT 64.000 361.600 64.800 370.200 ;
        RECT 66.800 361.600 67.600 370.200 ;
        RECT 71.000 361.600 71.800 366.200 ;
        RECT 73.800 361.600 74.600 366.200 ;
        RECT 78.000 361.600 78.800 370.200 ;
        RECT 79.600 361.600 80.400 370.200 ;
        RECT 83.800 361.600 84.600 366.200 ;
        RECT 86.600 361.600 87.400 366.200 ;
        RECT 90.800 361.600 91.600 370.200 ;
        RECT 94.000 361.600 94.800 370.200 ;
        RECT 99.600 361.600 100.400 366.200 ;
        RECT 102.800 361.600 103.600 366.200 ;
        RECT 108.400 361.600 109.200 370.000 ;
        RECT 111.600 361.600 112.400 366.200 ;
        RECT 115.400 361.600 116.200 366.200 ;
        RECT 119.600 361.600 120.400 370.200 ;
        RECT 121.200 361.600 122.000 370.200 ;
        RECT 125.400 361.600 126.200 366.200 ;
        RECT 129.200 361.600 130.000 369.800 ;
        RECT 134.400 361.600 135.200 370.200 ;
        RECT 137.200 361.600 138.000 370.200 ;
        RECT 141.400 361.600 142.200 366.200 ;
        RECT 143.600 361.600 144.400 370.200 ;
        RECT 147.800 361.600 148.600 366.200 ;
        RECT 156.400 361.600 157.200 370.000 ;
        RECT 162.000 361.600 162.800 366.200 ;
        RECT 165.200 361.600 166.000 366.200 ;
        RECT 170.800 361.600 171.600 370.200 ;
        RECT 177.200 369.600 178.000 370.200 ;
        RECT 180.400 370.000 181.400 370.200 ;
        RECT 174.000 361.600 174.800 366.200 ;
        RECT 177.200 361.600 178.000 366.200 ;
        RECT 180.400 361.600 181.200 366.200 ;
        RECT 186.800 361.600 187.600 366.200 ;
        RECT 190.000 361.600 190.800 366.200 ;
        RECT 198.000 361.600 198.800 366.200 ;
        RECT 201.200 361.600 202.000 366.200 ;
        RECT 204.400 361.600 205.200 366.200 ;
        RECT 207.600 361.600 208.400 366.200 ;
        RECT 209.200 361.600 210.000 366.200 ;
        RECT 212.400 361.600 213.200 366.200 ;
        RECT 214.600 361.600 215.400 366.200 ;
        RECT 218.800 361.600 219.600 370.200 ;
        RECT 221.000 361.600 221.800 366.200 ;
        RECT 225.200 361.600 226.000 370.200 ;
        RECT 226.800 361.600 227.600 370.200 ;
        RECT 260.200 370.000 261.000 370.200 ;
        RECT 263.600 369.600 264.400 370.200 ;
        RECT 231.000 361.600 231.800 366.200 ;
        RECT 233.200 361.600 234.000 366.200 ;
        RECT 236.400 361.600 237.200 366.200 ;
        RECT 239.600 361.600 240.400 366.200 ;
        RECT 242.800 361.600 243.600 366.200 ;
        RECT 250.800 361.600 251.600 366.200 ;
        RECT 254.000 361.600 254.800 366.200 ;
        RECT 260.400 361.600 261.200 366.200 ;
        RECT 263.600 361.600 264.400 366.200 ;
        RECT 266.800 361.600 267.600 366.200 ;
        RECT 268.400 361.600 269.200 370.200 ;
        RECT 271.600 361.600 272.400 369.000 ;
        RECT 274.800 361.600 275.600 370.200 ;
        RECT 278.000 361.600 278.800 370.200 ;
        RECT 281.200 361.600 282.000 370.200 ;
        RECT 284.400 361.600 285.200 370.200 ;
        RECT 287.600 361.600 288.400 370.200 ;
        RECT 289.200 361.600 290.000 370.200 ;
        RECT 292.400 361.600 293.200 370.200 ;
        RECT 295.600 361.600 296.400 370.200 ;
        RECT 298.800 361.600 299.600 370.200 ;
        RECT 302.000 361.600 302.800 370.200 ;
        RECT 310.000 361.600 310.800 369.800 ;
        RECT 315.200 361.600 316.000 370.200 ;
        RECT 319.600 361.600 320.400 366.200 ;
        RECT 321.800 361.600 322.600 366.200 ;
        RECT 326.000 361.600 326.800 370.200 ;
        RECT 329.200 361.600 330.000 366.200 ;
        RECT 332.400 361.600 333.200 369.800 ;
        RECT 337.600 361.600 338.400 370.200 ;
        RECT 346.800 369.600 347.600 370.200 ;
        RECT 350.000 370.000 351.000 370.200 ;
        RECT 405.800 370.000 406.800 370.200 ;
        RECT 409.200 369.600 410.000 370.200 ;
        RECT 342.000 361.600 342.800 366.200 ;
        RECT 343.600 361.600 344.400 366.200 ;
        RECT 346.800 361.600 347.600 366.200 ;
        RECT 350.000 361.600 350.800 366.200 ;
        RECT 356.400 361.600 357.200 366.200 ;
        RECT 359.600 361.600 360.400 366.200 ;
        RECT 367.600 361.600 368.400 366.200 ;
        RECT 370.800 361.600 371.600 366.200 ;
        RECT 374.000 361.600 374.800 366.200 ;
        RECT 377.200 361.600 378.000 366.200 ;
        RECT 378.800 361.600 379.600 366.200 ;
        RECT 382.000 361.600 382.800 366.200 ;
        RECT 385.200 361.600 386.000 366.200 ;
        RECT 388.400 361.600 389.200 366.200 ;
        RECT 396.400 361.600 397.200 366.200 ;
        RECT 399.600 361.600 400.400 366.200 ;
        RECT 406.000 361.600 406.800 366.200 ;
        RECT 409.200 361.600 410.000 366.200 ;
        RECT 412.400 361.600 413.200 366.200 ;
        RECT 415.600 361.600 416.400 369.000 ;
        RECT 418.800 361.600 419.600 370.200 ;
        RECT 420.400 361.600 421.200 366.200 ;
        RECT 423.600 361.600 424.400 366.200 ;
        RECT 425.800 361.600 426.600 366.200 ;
        RECT 430.000 361.600 430.800 370.200 ;
        RECT 431.600 361.600 432.400 370.200 ;
        RECT 474.600 370.000 475.600 370.200 ;
        RECT 478.000 369.600 478.800 370.200 ;
        RECT 435.800 361.600 436.600 366.200 ;
        RECT 438.000 361.600 438.800 366.200 ;
        RECT 441.200 361.600 442.000 366.200 ;
        RECT 447.600 361.600 448.400 366.200 ;
        RECT 450.800 361.600 451.600 366.200 ;
        RECT 454.000 361.600 454.800 366.200 ;
        RECT 457.200 361.600 458.000 366.200 ;
        RECT 465.200 361.600 466.000 366.200 ;
        RECT 468.400 361.600 469.200 366.200 ;
        RECT 474.800 361.600 475.600 366.200 ;
        RECT 478.000 361.600 478.800 366.200 ;
        RECT 481.200 361.600 482.000 366.200 ;
        RECT 484.400 361.600 485.200 366.200 ;
        RECT 486.000 361.600 486.800 370.200 ;
        RECT 489.200 361.600 490.000 370.200 ;
        RECT 492.400 361.600 493.200 370.200 ;
        RECT 495.600 361.600 496.400 370.200 ;
        RECT 498.800 361.600 499.600 370.200 ;
        RECT 500.400 361.600 501.200 370.200 ;
        RECT 503.600 361.600 504.400 369.000 ;
        RECT 506.800 361.600 507.600 370.200 ;
        RECT 510.000 361.600 510.800 369.000 ;
        RECT 513.200 361.600 514.000 370.200 ;
        RECT 516.400 361.600 517.200 369.000 ;
        RECT 519.600 361.600 520.400 366.200 ;
        RECT 522.800 361.600 523.600 366.200 ;
        RECT 526.000 361.600 526.800 366.200 ;
        RECT 529.200 361.600 530.000 366.200 ;
        RECT 537.200 361.600 538.000 366.200 ;
        RECT 540.400 361.600 541.200 366.200 ;
        RECT 546.800 361.600 547.600 366.200 ;
        RECT 550.000 361.600 550.800 366.200 ;
        RECT 553.200 361.600 554.000 366.200 ;
        RECT 556.400 361.600 557.200 369.000 ;
        RECT 559.600 361.600 560.400 370.200 ;
        RECT 561.200 361.600 562.000 366.200 ;
        RECT 564.400 361.600 565.200 366.200 ;
        RECT 566.000 361.600 566.800 370.200 ;
        RECT 599.400 370.000 600.200 370.200 ;
        RECT 602.800 369.600 603.600 370.200 ;
        RECT 570.200 361.600 571.000 366.200 ;
        RECT 572.400 361.600 573.200 366.200 ;
        RECT 575.600 361.600 576.400 366.200 ;
        RECT 578.800 361.600 579.600 366.200 ;
        RECT 582.000 361.600 582.800 366.200 ;
        RECT 590.000 361.600 590.800 366.200 ;
        RECT 593.200 361.600 594.000 366.200 ;
        RECT 599.600 361.600 600.400 366.200 ;
        RECT 602.800 361.600 603.600 366.200 ;
        RECT 606.000 361.600 606.800 366.200 ;
        RECT 609.200 361.600 610.000 369.000 ;
        RECT 0.400 360.400 614.000 361.600 ;
        RECT 1.200 355.800 2.000 360.400 ;
        RECT 4.400 351.800 5.200 360.400 ;
        RECT 8.600 355.800 9.400 360.400 ;
        RECT 10.800 355.800 11.600 360.400 ;
        RECT 14.000 355.800 14.800 360.400 ;
        RECT 17.200 355.800 18.000 360.400 ;
        RECT 23.600 355.800 24.400 360.400 ;
        RECT 26.800 355.800 27.600 360.400 ;
        RECT 34.800 355.800 35.600 360.400 ;
        RECT 38.000 355.800 38.800 360.400 ;
        RECT 41.200 355.800 42.000 360.400 ;
        RECT 44.400 355.800 45.200 360.400 ;
        RECT 46.000 355.800 46.800 360.400 ;
        RECT 50.800 355.800 51.600 360.400 ;
        RECT 52.400 355.800 53.200 360.400 ;
        RECT 55.600 355.800 56.400 360.400 ;
        RECT 58.800 355.800 59.600 360.400 ;
        RECT 14.000 351.800 14.800 352.400 ;
        RECT 62.000 352.000 62.800 360.400 ;
        RECT 67.600 355.800 68.400 360.400 ;
        RECT 70.800 355.800 71.600 360.400 ;
        RECT 17.400 351.800 18.200 352.000 ;
        RECT 76.400 351.800 77.200 360.400 ;
        RECT 81.200 355.800 82.000 360.400 ;
        RECT 82.800 355.800 83.600 360.400 ;
        RECT 86.000 355.800 86.800 360.400 ;
        RECT 88.200 355.800 89.000 360.400 ;
        RECT 92.400 351.800 93.200 360.400 ;
        RECT 94.600 355.800 95.400 360.400 ;
        RECT 98.800 351.800 99.600 360.400 ;
        RECT 102.000 355.800 102.800 360.400 ;
        RECT 105.200 352.200 106.000 360.400 ;
        RECT 110.400 351.800 111.200 360.400 ;
        RECT 113.200 351.800 114.000 360.400 ;
        RECT 117.400 355.800 118.200 360.400 ;
        RECT 120.200 355.800 121.000 360.400 ;
        RECT 124.400 351.800 125.200 360.400 ;
        RECT 126.600 355.800 127.400 360.400 ;
        RECT 130.800 351.800 131.600 360.400 ;
        RECT 134.000 352.200 134.800 360.400 ;
        RECT 139.200 351.800 140.000 360.400 ;
        RECT 142.000 351.800 142.800 360.400 ;
        RECT 145.200 351.800 146.000 360.400 ;
        RECT 148.400 351.800 149.200 360.400 ;
        RECT 151.600 351.800 152.400 360.400 ;
        RECT 154.800 351.800 155.600 360.400 ;
        RECT 161.200 355.800 162.000 360.400 ;
        RECT 165.600 351.800 166.400 360.400 ;
        RECT 170.800 352.200 171.600 360.400 ;
        RECT 175.600 353.000 176.400 360.400 ;
        RECT 178.800 355.800 179.600 360.400 ;
        RECT 182.000 355.800 182.800 360.400 ;
        RECT 185.200 355.800 186.000 360.400 ;
        RECT 191.600 355.800 192.400 360.400 ;
        RECT 194.800 355.800 195.600 360.400 ;
        RECT 202.800 355.800 203.600 360.400 ;
        RECT 206.000 355.800 206.800 360.400 ;
        RECT 209.200 355.800 210.000 360.400 ;
        RECT 212.400 355.800 213.200 360.400 ;
        RECT 182.000 351.800 182.800 352.400 ;
        RECT 185.400 351.800 186.200 352.000 ;
        RECT 214.000 351.800 214.800 360.400 ;
        RECT 217.200 353.000 218.000 360.400 ;
        RECT 220.400 351.800 221.200 360.400 ;
        RECT 223.600 351.800 224.400 360.400 ;
        RECT 226.800 351.800 227.600 360.400 ;
        RECT 230.000 353.000 230.800 360.400 ;
        RECT 233.200 351.800 234.000 360.400 ;
        RECT 234.800 355.800 235.600 360.400 ;
        RECT 238.000 355.800 238.800 360.400 ;
        RECT 241.200 355.800 242.000 360.400 ;
        RECT 247.600 355.800 248.400 360.400 ;
        RECT 250.800 355.800 251.600 360.400 ;
        RECT 258.800 355.800 259.600 360.400 ;
        RECT 262.000 355.800 262.800 360.400 ;
        RECT 265.200 355.800 266.000 360.400 ;
        RECT 268.400 355.800 269.200 360.400 ;
        RECT 238.000 351.800 238.800 352.400 ;
        RECT 271.600 352.200 272.400 360.400 ;
        RECT 241.400 351.800 242.200 352.000 ;
        RECT 276.800 351.800 277.600 360.400 ;
        RECT 281.200 355.800 282.000 360.400 ;
        RECT 282.800 355.800 283.600 360.400 ;
        RECT 286.000 355.800 286.800 360.400 ;
        RECT 289.200 355.800 290.000 360.400 ;
        RECT 292.400 355.800 293.200 360.400 ;
        RECT 298.800 355.800 299.600 360.400 ;
        RECT 302.000 355.800 302.800 360.400 ;
        RECT 310.000 355.800 310.800 360.400 ;
        RECT 313.200 355.800 314.000 360.400 ;
        RECT 316.400 355.800 317.200 360.400 ;
        RECT 319.600 355.800 320.400 360.400 ;
        RECT 289.200 351.800 290.000 352.400 ;
        RECT 327.600 352.200 328.400 360.400 ;
        RECT 292.400 351.800 293.400 352.000 ;
        RECT 332.800 351.800 333.600 360.400 ;
        RECT 337.200 355.800 338.000 360.400 ;
        RECT 338.800 355.800 339.600 360.400 ;
        RECT 342.000 355.800 342.800 360.400 ;
        RECT 345.200 355.800 346.000 360.400 ;
        RECT 351.600 355.800 352.400 360.400 ;
        RECT 354.800 355.800 355.600 360.400 ;
        RECT 362.800 355.800 363.600 360.400 ;
        RECT 366.000 355.800 366.800 360.400 ;
        RECT 369.200 355.800 370.000 360.400 ;
        RECT 372.400 355.800 373.200 360.400 ;
        RECT 374.000 355.800 374.800 360.400 ;
        RECT 377.200 355.800 378.000 360.400 ;
        RECT 380.400 355.800 381.200 360.400 ;
        RECT 342.000 351.800 342.800 352.400 ;
        RECT 345.400 351.800 346.200 352.000 ;
        RECT 383.200 351.800 384.000 360.400 ;
        RECT 388.400 352.200 389.200 360.400 ;
        RECT 392.800 351.800 393.600 360.400 ;
        RECT 398.000 352.200 398.800 360.400 ;
        RECT 401.200 355.800 402.000 360.400 ;
        RECT 404.400 355.800 405.200 360.400 ;
        RECT 407.600 355.800 408.400 360.400 ;
        RECT 409.200 355.800 410.000 360.400 ;
        RECT 412.400 355.800 413.200 360.400 ;
        RECT 414.000 355.800 414.800 360.400 ;
        RECT 417.200 355.800 418.000 360.400 ;
        RECT 420.400 355.800 421.200 360.400 ;
        RECT 423.600 355.800 424.400 360.400 ;
        RECT 431.600 355.800 432.400 360.400 ;
        RECT 434.800 355.800 435.600 360.400 ;
        RECT 441.200 355.800 442.000 360.400 ;
        RECT 444.400 355.800 445.200 360.400 ;
        RECT 447.600 355.800 448.400 360.400 ;
        RECT 441.000 351.800 441.800 352.000 ;
        RECT 444.400 351.800 445.200 352.400 ;
        RECT 449.200 351.800 450.000 360.400 ;
        RECT 458.800 355.800 459.600 360.400 ;
        RECT 462.000 355.800 462.800 360.400 ;
        RECT 465.200 355.800 466.000 360.400 ;
        RECT 468.400 355.800 469.200 360.400 ;
        RECT 476.400 355.800 477.200 360.400 ;
        RECT 479.600 355.800 480.400 360.400 ;
        RECT 486.000 355.800 486.800 360.400 ;
        RECT 489.200 355.800 490.000 360.400 ;
        RECT 492.400 355.800 493.200 360.400 ;
        RECT 494.000 355.800 494.800 360.400 ;
        RECT 497.200 355.800 498.000 360.400 ;
        RECT 500.400 355.800 501.200 360.400 ;
        RECT 506.800 355.800 507.600 360.400 ;
        RECT 510.000 355.800 510.800 360.400 ;
        RECT 518.000 355.800 518.800 360.400 ;
        RECT 521.200 355.800 522.000 360.400 ;
        RECT 524.400 355.800 525.200 360.400 ;
        RECT 527.600 355.800 528.400 360.400 ;
        RECT 529.200 355.800 530.000 360.400 ;
        RECT 532.400 355.800 533.200 360.400 ;
        RECT 485.800 351.800 486.800 352.000 ;
        RECT 489.200 351.800 490.000 352.400 ;
        RECT 14.000 351.200 41.000 351.800 ;
        RECT 182.000 351.200 209.000 351.800 ;
        RECT 238.000 351.200 265.000 351.800 ;
        RECT 289.200 351.200 316.200 351.800 ;
        RECT 342.000 351.200 369.000 351.800 ;
        RECT 40.200 351.000 41.000 351.200 ;
        RECT 208.200 351.000 209.000 351.200 ;
        RECT 264.200 351.000 265.000 351.200 ;
        RECT 315.400 351.000 316.200 351.200 ;
        RECT 368.200 351.000 369.000 351.200 ;
        RECT 418.200 351.200 445.200 351.800 ;
        RECT 463.000 351.200 490.000 351.800 ;
        RECT 497.200 351.800 498.000 352.400 ;
        RECT 500.400 351.800 501.400 352.000 ;
        RECT 534.000 351.800 534.800 360.400 ;
        RECT 537.200 353.000 538.000 360.400 ;
        RECT 542.000 353.000 542.800 360.400 ;
        RECT 545.200 351.800 546.000 360.400 ;
        RECT 546.800 351.800 547.600 360.400 ;
        RECT 550.000 351.800 550.800 360.400 ;
        RECT 553.200 351.800 554.000 360.400 ;
        RECT 554.800 355.800 555.600 360.400 ;
        RECT 558.000 355.800 558.800 360.400 ;
        RECT 559.600 351.800 560.400 360.400 ;
        RECT 563.800 355.800 564.600 360.400 ;
        RECT 566.000 355.800 566.800 360.400 ;
        RECT 569.200 355.800 570.000 360.400 ;
        RECT 572.400 355.800 573.200 360.400 ;
        RECT 578.800 355.800 579.600 360.400 ;
        RECT 582.000 355.800 582.800 360.400 ;
        RECT 590.000 355.800 590.800 360.400 ;
        RECT 593.200 355.800 594.000 360.400 ;
        RECT 596.400 355.800 597.200 360.400 ;
        RECT 599.600 355.800 600.400 360.400 ;
        RECT 601.200 355.800 602.000 360.400 ;
        RECT 604.400 355.800 605.200 360.400 ;
        RECT 607.600 353.000 608.400 360.400 ;
        RECT 569.200 351.800 570.000 352.400 ;
        RECT 572.600 351.800 573.400 352.000 ;
        RECT 497.200 351.200 524.200 351.800 ;
        RECT 569.200 351.200 596.200 351.800 ;
        RECT 418.200 351.000 419.000 351.200 ;
        RECT 463.000 351.000 463.800 351.200 ;
        RECT 523.400 351.000 524.200 351.200 ;
        RECT 595.400 351.000 596.200 351.200 ;
        RECT 30.600 330.800 31.400 331.000 ;
        RECT 4.400 330.200 31.400 330.800 ;
        RECT 63.000 330.800 63.800 331.000 ;
        RECT 157.400 330.800 158.200 331.000 ;
        RECT 224.200 330.800 225.000 331.000 ;
        RECT 270.600 330.800 271.400 331.000 ;
        RECT 63.000 330.200 90.000 330.800 ;
        RECT 157.400 330.200 184.400 330.800 ;
        RECT 198.000 330.200 225.000 330.800 ;
        RECT 244.400 330.200 271.400 330.800 ;
        RECT 339.800 330.800 340.600 331.000 ;
        RECT 400.600 330.800 401.400 331.000 ;
        RECT 509.400 330.800 510.200 331.000 ;
        RECT 569.800 330.800 570.600 331.000 ;
        RECT 339.800 330.200 366.800 330.800 ;
        RECT 400.600 330.200 427.600 330.800 ;
        RECT 509.400 330.200 536.400 330.800 ;
        RECT 4.400 329.600 5.200 330.200 ;
        RECT 7.800 330.000 8.600 330.200 ;
        RECT 1.200 321.600 2.000 326.200 ;
        RECT 4.400 321.600 5.200 326.200 ;
        RECT 7.600 321.600 8.400 326.200 ;
        RECT 14.000 321.600 14.800 326.200 ;
        RECT 17.200 321.600 18.000 326.200 ;
        RECT 25.200 321.600 26.000 326.200 ;
        RECT 28.400 321.600 29.200 326.200 ;
        RECT 31.600 321.600 32.400 326.200 ;
        RECT 34.800 321.600 35.600 326.200 ;
        RECT 36.400 321.600 37.200 330.200 ;
        RECT 39.600 321.600 40.400 329.000 ;
        RECT 44.400 321.600 45.200 326.200 ;
        RECT 47.200 321.600 48.000 330.200 ;
        RECT 85.800 330.000 86.600 330.200 ;
        RECT 52.400 321.600 53.200 329.800 ;
        RECT 89.200 329.600 90.000 330.200 ;
        RECT 55.600 321.600 56.400 326.200 ;
        RECT 58.800 321.600 59.600 326.200 ;
        RECT 62.000 321.600 62.800 326.200 ;
        RECT 65.200 321.600 66.000 326.200 ;
        RECT 68.400 321.600 69.200 326.200 ;
        RECT 76.400 321.600 77.200 326.200 ;
        RECT 79.600 321.600 80.400 326.200 ;
        RECT 86.000 321.600 86.800 326.200 ;
        RECT 89.200 321.600 90.000 326.200 ;
        RECT 92.400 321.600 93.200 326.200 ;
        RECT 94.000 321.600 94.800 326.200 ;
        RECT 98.400 321.600 99.200 330.200 ;
        RECT 103.600 321.600 104.400 329.800 ;
        RECT 108.400 321.600 109.200 330.000 ;
        RECT 114.000 321.600 114.800 326.200 ;
        RECT 117.200 321.600 118.000 326.200 ;
        RECT 122.800 321.600 123.600 330.200 ;
        RECT 127.600 321.600 128.400 330.000 ;
        RECT 133.200 321.600 134.000 326.200 ;
        RECT 136.400 321.600 137.200 326.200 ;
        RECT 142.000 321.600 142.800 330.200 ;
        RECT 180.200 330.000 181.000 330.200 ;
        RECT 183.600 329.600 184.400 330.200 ;
        RECT 146.800 321.600 147.600 326.200 ;
        RECT 153.200 321.600 154.000 326.200 ;
        RECT 156.400 321.600 157.200 326.200 ;
        RECT 159.600 321.600 160.400 326.200 ;
        RECT 162.800 321.600 163.600 326.200 ;
        RECT 170.800 321.600 171.600 326.200 ;
        RECT 174.000 321.600 174.800 326.200 ;
        RECT 180.400 321.600 181.200 326.200 ;
        RECT 183.600 321.600 184.400 326.200 ;
        RECT 186.800 321.600 187.600 326.200 ;
        RECT 190.000 321.600 190.800 329.000 ;
        RECT 193.200 321.600 194.000 330.200 ;
        RECT 198.000 329.600 198.800 330.200 ;
        RECT 201.200 330.000 202.200 330.200 ;
        RECT 194.800 321.600 195.600 326.200 ;
        RECT 198.000 321.600 198.800 326.200 ;
        RECT 201.200 321.600 202.000 326.200 ;
        RECT 207.600 321.600 208.400 326.200 ;
        RECT 210.800 321.600 211.600 326.200 ;
        RECT 218.800 321.600 219.600 326.200 ;
        RECT 222.000 321.600 222.800 326.200 ;
        RECT 225.200 321.600 226.000 326.200 ;
        RECT 228.400 321.600 229.200 326.200 ;
        RECT 230.000 321.600 230.800 330.200 ;
        RECT 233.200 321.600 234.000 330.200 ;
        RECT 236.400 321.600 237.200 330.200 ;
        RECT 244.400 329.600 245.200 330.200 ;
        RECT 247.600 330.000 248.600 330.200 ;
        RECT 238.000 321.600 238.800 326.200 ;
        RECT 241.200 321.600 242.000 326.200 ;
        RECT 244.400 321.600 245.200 326.200 ;
        RECT 247.600 321.600 248.400 326.200 ;
        RECT 254.000 321.600 254.800 326.200 ;
        RECT 257.200 321.600 258.000 326.200 ;
        RECT 265.200 321.600 266.000 326.200 ;
        RECT 268.400 321.600 269.200 326.200 ;
        RECT 271.600 321.600 272.400 326.200 ;
        RECT 274.800 321.600 275.600 326.200 ;
        RECT 278.000 321.600 278.800 326.200 ;
        RECT 281.200 321.600 282.000 325.800 ;
        RECT 284.400 321.600 285.200 326.200 ;
        RECT 287.600 321.600 288.400 325.800 ;
        RECT 290.800 321.600 291.600 326.200 ;
        RECT 294.000 321.600 294.800 325.800 ;
        RECT 297.200 321.600 298.000 326.200 ;
        RECT 300.400 321.600 301.200 325.800 ;
        RECT 303.600 321.600 304.400 326.200 ;
        RECT 310.000 321.600 310.800 330.200 ;
        RECT 313.200 321.600 314.000 329.000 ;
        RECT 316.400 321.600 317.200 326.200 ;
        RECT 319.600 321.600 320.400 326.200 ;
        RECT 321.200 321.600 322.000 330.200 ;
        RECT 327.600 321.600 328.400 330.200 ;
        RECT 329.800 321.600 330.600 326.200 ;
        RECT 334.000 321.600 334.800 330.200 ;
        RECT 362.600 330.000 363.400 330.200 ;
        RECT 366.000 329.600 366.800 330.200 ;
        RECT 335.600 321.600 336.400 326.200 ;
        RECT 338.800 321.600 339.600 326.200 ;
        RECT 342.000 321.600 342.800 326.200 ;
        RECT 345.200 321.600 346.000 326.200 ;
        RECT 353.200 321.600 354.000 326.200 ;
        RECT 356.400 321.600 357.200 326.200 ;
        RECT 362.800 321.600 363.600 326.200 ;
        RECT 366.000 321.600 366.800 326.200 ;
        RECT 369.200 321.600 370.000 326.200 ;
        RECT 371.400 321.600 372.200 326.200 ;
        RECT 375.600 321.600 376.400 330.200 ;
        RECT 377.200 321.600 378.000 330.200 ;
        RECT 383.600 321.600 384.400 330.200 ;
        RECT 385.200 321.600 386.000 326.200 ;
        RECT 388.400 321.600 389.200 326.200 ;
        RECT 390.000 321.600 390.800 330.200 ;
        RECT 423.400 330.000 424.200 330.200 ;
        RECT 426.800 329.600 427.600 330.200 ;
        RECT 393.200 321.600 394.000 329.000 ;
        RECT 396.400 321.600 397.200 326.200 ;
        RECT 399.600 321.600 400.400 326.200 ;
        RECT 402.800 321.600 403.600 326.200 ;
        RECT 406.000 321.600 406.800 326.200 ;
        RECT 414.000 321.600 414.800 326.200 ;
        RECT 417.200 321.600 418.000 326.200 ;
        RECT 423.600 321.600 424.400 326.200 ;
        RECT 426.800 321.600 427.600 326.200 ;
        RECT 430.000 321.600 430.800 326.200 ;
        RECT 431.600 321.600 432.400 326.200 ;
        RECT 434.800 321.600 435.600 326.200 ;
        RECT 436.400 321.600 437.200 326.200 ;
        RECT 439.600 321.600 440.400 330.200 ;
        RECT 443.800 321.600 444.600 326.200 ;
        RECT 446.000 321.600 446.800 330.200 ;
        RECT 450.200 321.600 451.000 326.200 ;
        RECT 452.400 321.600 453.200 326.200 ;
        RECT 455.600 321.600 456.400 326.200 ;
        RECT 463.600 321.600 464.400 329.000 ;
        RECT 468.400 321.600 469.200 330.200 ;
        RECT 476.400 321.600 477.200 330.200 ;
        RECT 478.600 321.600 479.400 326.200 ;
        RECT 482.800 321.600 483.600 330.200 ;
        RECT 484.400 321.600 485.200 326.200 ;
        RECT 487.600 321.600 488.400 326.200 ;
        RECT 489.200 321.600 490.000 330.200 ;
        RECT 492.400 321.600 493.200 330.200 ;
        RECT 494.000 321.600 494.800 326.200 ;
        RECT 497.200 321.600 498.000 325.800 ;
        RECT 503.600 321.600 504.400 330.200 ;
        RECT 532.200 330.000 533.200 330.200 ;
        RECT 535.600 329.600 536.400 330.200 ;
        RECT 543.600 330.200 570.600 330.800 ;
        RECT 543.600 329.600 544.400 330.200 ;
        RECT 547.000 330.000 547.800 330.200 ;
        RECT 505.200 321.600 506.000 326.200 ;
        RECT 508.400 321.600 509.200 326.200 ;
        RECT 511.600 321.600 512.400 326.200 ;
        RECT 514.800 321.600 515.600 326.200 ;
        RECT 522.800 321.600 523.600 326.200 ;
        RECT 526.000 321.600 526.800 326.200 ;
        RECT 532.400 321.600 533.200 326.200 ;
        RECT 535.600 321.600 536.400 326.200 ;
        RECT 538.800 321.600 539.600 326.200 ;
        RECT 540.400 321.600 541.200 326.200 ;
        RECT 543.600 321.600 544.400 326.200 ;
        RECT 546.800 321.600 547.600 326.200 ;
        RECT 553.200 321.600 554.000 326.200 ;
        RECT 556.400 321.600 557.200 326.200 ;
        RECT 564.400 321.600 565.200 326.200 ;
        RECT 567.600 321.600 568.400 326.200 ;
        RECT 570.800 321.600 571.600 326.200 ;
        RECT 574.000 321.600 574.800 326.200 ;
        RECT 575.600 321.600 576.400 326.200 ;
        RECT 578.800 321.600 579.600 326.200 ;
        RECT 581.000 321.600 581.800 326.200 ;
        RECT 585.200 321.600 586.000 330.200 ;
        RECT 588.400 321.600 589.200 326.200 ;
        RECT 590.000 321.600 590.800 326.200 ;
        RECT 593.200 321.600 594.000 326.200 ;
        RECT 595.400 321.600 596.200 326.200 ;
        RECT 599.600 321.600 600.400 330.200 ;
        RECT 602.800 321.600 603.600 326.200 ;
        RECT 604.400 321.600 605.200 330.200 ;
        RECT 607.600 321.600 608.400 330.200 ;
        RECT 610.800 321.600 611.600 330.200 ;
        RECT 0.400 320.400 614.000 321.600 ;
        RECT 1.200 311.800 2.000 320.400 ;
        RECT 4.400 311.800 5.200 320.400 ;
        RECT 7.600 311.800 8.400 320.400 ;
        RECT 10.800 311.800 11.600 320.400 ;
        RECT 14.000 311.800 14.800 320.400 ;
        RECT 15.600 315.800 16.400 320.400 ;
        RECT 18.800 315.800 19.600 320.400 ;
        RECT 22.000 315.800 22.800 320.400 ;
        RECT 28.400 315.800 29.200 320.400 ;
        RECT 31.600 315.800 32.400 320.400 ;
        RECT 39.600 315.800 40.400 320.400 ;
        RECT 42.800 315.800 43.600 320.400 ;
        RECT 46.000 315.800 46.800 320.400 ;
        RECT 49.200 315.800 50.000 320.400 ;
        RECT 50.800 315.800 51.600 320.400 ;
        RECT 54.000 315.800 54.800 320.400 ;
        RECT 57.200 315.800 58.000 320.400 ;
        RECT 60.400 315.800 61.200 320.400 ;
        RECT 68.400 315.800 69.200 320.400 ;
        RECT 71.600 315.800 72.400 320.400 ;
        RECT 78.000 315.800 78.800 320.400 ;
        RECT 81.200 315.800 82.000 320.400 ;
        RECT 84.400 315.800 85.200 320.400 ;
        RECT 18.800 311.800 19.600 312.400 ;
        RECT 22.200 311.800 23.000 312.000 ;
        RECT 77.800 311.800 78.600 312.000 ;
        RECT 81.200 311.800 82.000 312.400 ;
        RECT 87.200 311.800 88.000 320.400 ;
        RECT 92.400 312.200 93.200 320.400 ;
        RECT 97.200 312.200 98.000 320.400 ;
        RECT 102.400 311.800 103.200 320.400 ;
        RECT 106.800 315.800 107.600 320.400 ;
        RECT 108.400 315.800 109.200 320.400 ;
        RECT 111.600 315.800 112.400 320.400 ;
        RECT 114.800 315.800 115.600 320.400 ;
        RECT 118.000 315.800 118.800 320.400 ;
        RECT 126.000 315.800 126.800 320.400 ;
        RECT 129.200 315.800 130.000 320.400 ;
        RECT 135.600 315.800 136.400 320.400 ;
        RECT 138.800 315.800 139.600 320.400 ;
        RECT 142.000 315.800 142.800 320.400 ;
        RECT 135.400 311.800 136.200 312.000 ;
        RECT 138.800 311.800 139.600 312.400 ;
        RECT 143.600 311.800 144.400 320.400 ;
        RECT 156.400 313.000 157.200 320.400 ;
        RECT 159.600 315.800 160.400 320.400 ;
        RECT 162.800 315.800 163.600 320.400 ;
        RECT 166.000 315.800 166.800 320.400 ;
        RECT 169.200 315.800 170.000 320.400 ;
        RECT 177.200 315.800 178.000 320.400 ;
        RECT 180.400 315.800 181.200 320.400 ;
        RECT 186.800 315.800 187.600 320.400 ;
        RECT 190.000 315.800 190.800 320.400 ;
        RECT 193.200 315.800 194.000 320.400 ;
        RECT 194.800 315.800 195.600 320.400 ;
        RECT 198.000 316.200 198.800 320.400 ;
        RECT 201.200 315.800 202.000 320.400 ;
        RECT 204.400 315.800 205.200 320.400 ;
        RECT 207.600 315.800 208.400 320.400 ;
        RECT 214.000 315.800 214.800 320.400 ;
        RECT 217.200 315.800 218.000 320.400 ;
        RECT 225.200 315.800 226.000 320.400 ;
        RECT 228.400 315.800 229.200 320.400 ;
        RECT 231.600 315.800 232.400 320.400 ;
        RECT 234.800 315.800 235.600 320.400 ;
        RECT 186.600 311.800 187.600 312.000 ;
        RECT 190.000 311.800 190.800 312.400 ;
        RECT 18.800 311.200 45.800 311.800 ;
        RECT 45.000 311.000 45.800 311.200 ;
        RECT 55.000 311.200 82.000 311.800 ;
        RECT 112.600 311.200 139.600 311.800 ;
        RECT 163.800 311.200 190.800 311.800 ;
        RECT 204.400 311.800 205.200 312.400 ;
        RECT 207.600 311.800 208.600 312.000 ;
        RECT 238.000 311.800 238.800 320.400 ;
        RECT 239.600 315.800 240.400 320.400 ;
        RECT 242.800 315.800 243.600 320.400 ;
        RECT 244.400 315.800 245.200 320.400 ;
        RECT 247.600 315.800 248.400 320.400 ;
        RECT 250.800 313.000 251.600 320.400 ;
        RECT 254.000 311.800 254.800 320.400 ;
        RECT 256.800 311.800 257.600 320.400 ;
        RECT 262.000 312.200 262.800 320.400 ;
        RECT 266.800 312.200 267.600 320.400 ;
        RECT 272.000 311.800 272.800 320.400 ;
        RECT 275.400 315.800 276.200 320.400 ;
        RECT 279.600 311.800 280.400 320.400 ;
        RECT 281.200 315.800 282.000 320.400 ;
        RECT 284.400 315.800 285.200 320.400 ;
        RECT 287.600 311.800 288.400 320.400 ;
        RECT 290.800 311.800 291.600 320.400 ;
        RECT 297.200 315.800 298.000 320.400 ;
        RECT 300.400 315.800 301.200 320.400 ;
        RECT 303.600 315.800 304.400 320.400 ;
        RECT 306.800 315.800 307.600 320.400 ;
        RECT 314.800 315.800 315.600 320.400 ;
        RECT 318.000 315.800 318.800 320.400 ;
        RECT 324.400 315.800 325.200 320.400 ;
        RECT 327.600 315.800 328.400 320.400 ;
        RECT 330.800 315.800 331.600 320.400 ;
        RECT 332.400 315.800 333.200 320.400 ;
        RECT 335.600 315.800 336.400 320.400 ;
        RECT 337.200 315.800 338.000 320.400 ;
        RECT 340.400 315.800 341.200 320.400 ;
        RECT 342.600 315.800 343.400 320.400 ;
        RECT 324.200 311.800 325.200 312.000 ;
        RECT 327.600 311.800 328.400 312.400 ;
        RECT 346.800 311.800 347.600 320.400 ;
        RECT 349.000 315.800 349.800 320.400 ;
        RECT 353.200 311.800 354.000 320.400 ;
        RECT 356.400 315.800 357.200 320.400 ;
        RECT 358.000 315.800 358.800 320.400 ;
        RECT 361.200 316.200 362.000 320.400 ;
        RECT 364.400 311.800 365.200 320.400 ;
        RECT 367.600 311.800 368.400 320.400 ;
        RECT 369.200 315.800 370.000 320.400 ;
        RECT 372.400 316.200 373.200 320.400 ;
        RECT 380.400 313.000 381.200 320.400 ;
        RECT 383.600 315.800 384.400 320.400 ;
        RECT 386.800 315.800 387.600 320.400 ;
        RECT 390.000 313.000 390.800 320.400 ;
        RECT 396.400 311.800 397.200 320.400 ;
        RECT 400.600 315.800 401.400 320.400 ;
        RECT 402.800 311.800 403.600 320.400 ;
        RECT 407.000 315.800 407.800 320.400 ;
        RECT 410.800 315.800 411.600 320.400 ;
        RECT 413.000 315.800 413.800 320.400 ;
        RECT 417.200 311.800 418.000 320.400 ;
        RECT 418.800 311.800 419.600 320.400 ;
        RECT 423.000 315.800 423.800 320.400 ;
        RECT 425.200 315.800 426.000 320.400 ;
        RECT 428.400 315.800 429.200 320.400 ;
        RECT 431.600 315.800 432.400 320.400 ;
        RECT 438.000 315.800 438.800 320.400 ;
        RECT 441.200 315.800 442.000 320.400 ;
        RECT 449.200 315.800 450.000 320.400 ;
        RECT 452.400 315.800 453.200 320.400 ;
        RECT 455.600 315.800 456.400 320.400 ;
        RECT 458.800 315.800 459.600 320.400 ;
        RECT 428.400 311.800 429.200 312.400 ;
        RECT 431.800 311.800 432.600 312.000 ;
        RECT 465.200 311.800 466.000 320.400 ;
        RECT 469.400 315.800 470.200 320.400 ;
        RECT 471.600 315.800 472.400 320.400 ;
        RECT 474.800 311.800 475.600 320.400 ;
        RECT 479.000 315.800 479.800 320.400 ;
        RECT 481.800 315.800 482.600 320.400 ;
        RECT 486.000 311.800 486.800 320.400 ;
        RECT 488.200 315.800 489.000 320.400 ;
        RECT 492.400 311.800 493.200 320.400 ;
        RECT 497.200 313.000 498.000 320.400 ;
        RECT 500.400 311.800 501.200 320.400 ;
        RECT 504.600 315.800 505.400 320.400 ;
        RECT 506.800 311.800 507.600 320.400 ;
        RECT 511.000 315.800 511.800 320.400 ;
        RECT 513.200 315.800 514.000 320.400 ;
        RECT 516.400 315.800 517.200 320.400 ;
        RECT 518.000 315.800 518.800 320.400 ;
        RECT 521.200 315.800 522.000 320.400 ;
        RECT 523.400 315.800 524.200 320.400 ;
        RECT 527.600 311.800 528.400 320.400 ;
        RECT 530.800 313.000 531.600 320.400 ;
        RECT 534.000 315.800 534.800 320.400 ;
        RECT 537.200 315.800 538.000 320.400 ;
        RECT 540.400 313.000 541.200 320.400 ;
        RECT 543.600 311.800 544.400 320.400 ;
        RECT 545.200 311.800 546.000 320.400 ;
        RECT 548.400 311.800 549.200 320.400 ;
        RECT 550.000 315.800 550.800 320.400 ;
        RECT 553.200 315.800 554.000 320.400 ;
        RECT 556.400 315.800 557.200 320.400 ;
        RECT 562.800 315.800 563.600 320.400 ;
        RECT 566.000 315.800 566.800 320.400 ;
        RECT 574.000 315.800 574.800 320.400 ;
        RECT 577.200 315.800 578.000 320.400 ;
        RECT 580.400 315.800 581.200 320.400 ;
        RECT 583.600 315.800 584.400 320.400 ;
        RECT 585.800 315.800 586.600 320.400 ;
        RECT 553.200 311.800 554.000 312.400 ;
        RECT 556.600 311.800 557.400 312.000 ;
        RECT 590.000 311.800 590.800 320.400 ;
        RECT 593.200 315.800 594.000 320.400 ;
        RECT 595.400 315.800 596.200 320.400 ;
        RECT 599.600 311.800 600.400 320.400 ;
        RECT 602.800 315.800 603.600 320.400 ;
        RECT 606.000 313.000 606.800 320.400 ;
        RECT 204.400 311.200 231.400 311.800 ;
        RECT 55.000 311.000 55.800 311.200 ;
        RECT 112.600 311.000 113.400 311.200 ;
        RECT 163.800 311.000 164.600 311.200 ;
        RECT 230.600 311.000 231.400 311.200 ;
        RECT 301.400 311.200 328.400 311.800 ;
        RECT 428.400 311.200 455.400 311.800 ;
        RECT 553.200 311.200 580.200 311.800 ;
        RECT 301.400 311.000 302.200 311.200 ;
        RECT 454.600 311.000 455.400 311.200 ;
        RECT 579.400 311.000 580.200 311.200 ;
        RECT 45.000 290.800 45.800 291.000 ;
        RECT 91.400 290.800 92.200 291.000 ;
        RECT 18.800 290.200 45.800 290.800 ;
        RECT 65.200 290.200 92.200 290.800 ;
        RECT 125.400 290.800 126.200 291.000 ;
        RECT 200.200 290.800 201.000 291.000 ;
        RECT 248.200 290.800 249.000 291.000 ;
        RECT 296.200 290.800 297.000 291.000 ;
        RECT 125.400 290.200 152.400 290.800 ;
        RECT 174.000 290.200 201.000 290.800 ;
        RECT 222.000 290.200 249.000 290.800 ;
        RECT 270.000 290.200 297.000 290.800 ;
        RECT 402.200 290.800 403.000 291.000 ;
        RECT 541.400 290.800 542.200 291.000 ;
        RECT 606.600 290.800 607.400 291.000 ;
        RECT 402.200 290.200 429.200 290.800 ;
        RECT 541.400 290.200 568.400 290.800 ;
        RECT 1.200 281.600 2.000 290.200 ;
        RECT 4.400 281.600 5.200 290.200 ;
        RECT 7.600 281.600 8.400 290.200 ;
        RECT 10.800 281.600 11.600 290.200 ;
        RECT 14.000 281.600 14.800 290.200 ;
        RECT 18.800 289.600 19.600 290.200 ;
        RECT 22.200 290.000 23.000 290.200 ;
        RECT 15.600 281.600 16.400 286.200 ;
        RECT 18.800 281.600 19.600 286.200 ;
        RECT 22.000 281.600 22.800 286.200 ;
        RECT 28.400 281.600 29.200 286.200 ;
        RECT 31.600 281.600 32.400 286.200 ;
        RECT 39.600 281.600 40.400 286.200 ;
        RECT 42.800 281.600 43.600 286.200 ;
        RECT 46.000 281.600 46.800 286.200 ;
        RECT 49.200 281.600 50.000 286.200 ;
        RECT 50.800 281.600 51.600 290.200 ;
        RECT 65.200 289.600 66.000 290.200 ;
        RECT 68.600 290.000 69.400 290.200 ;
        RECT 58.800 281.600 59.600 289.000 ;
        RECT 62.000 281.600 62.800 286.200 ;
        RECT 65.200 281.600 66.000 286.200 ;
        RECT 68.400 281.600 69.200 286.200 ;
        RECT 74.800 281.600 75.600 286.200 ;
        RECT 78.000 281.600 78.800 286.200 ;
        RECT 86.000 281.600 86.800 286.200 ;
        RECT 89.200 281.600 90.000 286.200 ;
        RECT 92.400 281.600 93.200 286.200 ;
        RECT 95.600 281.600 96.400 286.200 ;
        RECT 97.200 281.600 98.000 290.200 ;
        RECT 105.200 281.600 106.000 289.000 ;
        RECT 108.400 281.600 109.200 286.200 ;
        RECT 113.200 281.600 114.000 289.800 ;
        RECT 118.400 281.600 119.200 290.200 ;
        RECT 148.200 290.000 149.200 290.200 ;
        RECT 151.600 289.600 152.400 290.200 ;
        RECT 121.200 281.600 122.000 286.200 ;
        RECT 124.400 281.600 125.200 286.200 ;
        RECT 127.600 281.600 128.400 286.200 ;
        RECT 130.800 281.600 131.600 286.200 ;
        RECT 138.800 281.600 139.600 286.200 ;
        RECT 142.000 281.600 142.800 286.200 ;
        RECT 148.400 281.600 149.200 286.200 ;
        RECT 151.600 281.600 152.400 286.200 ;
        RECT 154.800 281.600 155.600 286.200 ;
        RECT 161.200 281.600 162.000 286.200 ;
        RECT 164.400 281.600 165.200 290.200 ;
        RECT 174.000 289.600 174.800 290.200 ;
        RECT 177.200 290.000 178.200 290.200 ;
        RECT 168.600 281.600 169.400 286.200 ;
        RECT 170.800 281.600 171.600 286.200 ;
        RECT 174.000 281.600 174.800 286.200 ;
        RECT 177.200 281.600 178.000 286.200 ;
        RECT 183.600 281.600 184.400 286.200 ;
        RECT 186.800 281.600 187.600 286.200 ;
        RECT 194.800 281.600 195.600 286.200 ;
        RECT 198.000 281.600 198.800 286.200 ;
        RECT 201.200 281.600 202.000 286.200 ;
        RECT 204.400 281.600 205.200 286.200 ;
        RECT 206.000 281.600 206.800 290.200 ;
        RECT 222.000 289.600 222.800 290.200 ;
        RECT 225.400 290.000 226.200 290.200 ;
        RECT 209.200 281.600 210.000 286.200 ;
        RECT 212.400 281.600 213.200 286.200 ;
        RECT 214.000 281.600 214.800 286.200 ;
        RECT 217.200 281.600 218.000 286.200 ;
        RECT 218.800 281.600 219.600 286.200 ;
        RECT 222.000 281.600 222.800 286.200 ;
        RECT 225.200 281.600 226.000 286.200 ;
        RECT 231.600 281.600 232.400 286.200 ;
        RECT 234.800 281.600 235.600 286.200 ;
        RECT 242.800 281.600 243.600 286.200 ;
        RECT 246.000 281.600 246.800 286.200 ;
        RECT 249.200 281.600 250.000 286.200 ;
        RECT 252.400 281.600 253.200 286.200 ;
        RECT 254.000 281.600 254.800 286.200 ;
        RECT 258.400 281.600 259.200 290.200 ;
        RECT 263.600 281.600 264.400 289.800 ;
        RECT 270.000 289.600 270.800 290.200 ;
        RECT 273.400 290.000 274.200 290.200 ;
        RECT 266.800 281.600 267.600 286.200 ;
        RECT 270.000 281.600 270.800 286.200 ;
        RECT 273.200 281.600 274.000 286.200 ;
        RECT 279.600 281.600 280.400 286.200 ;
        RECT 282.800 281.600 283.600 286.200 ;
        RECT 290.800 281.600 291.600 286.200 ;
        RECT 294.000 281.600 294.800 286.200 ;
        RECT 297.200 281.600 298.000 286.200 ;
        RECT 300.400 281.600 301.200 286.200 ;
        RECT 302.000 281.600 302.800 286.200 ;
        RECT 305.200 281.600 306.000 286.200 ;
        RECT 311.600 281.600 312.400 286.200 ;
        RECT 314.800 281.600 315.600 286.200 ;
        RECT 316.400 281.600 317.200 286.200 ;
        RECT 319.600 281.600 320.400 286.200 ;
        RECT 321.200 281.600 322.000 290.200 ;
        RECT 325.400 281.600 326.200 286.200 ;
        RECT 327.600 281.600 328.400 290.200 ;
        RECT 331.800 281.600 332.600 286.200 ;
        RECT 334.000 281.600 334.800 286.200 ;
        RECT 337.200 281.600 338.000 286.200 ;
        RECT 338.800 281.600 339.600 290.200 ;
        RECT 345.200 281.600 346.000 286.200 ;
        RECT 346.800 281.600 347.600 286.200 ;
        RECT 350.000 281.600 350.800 285.800 ;
        RECT 353.200 281.600 354.000 286.200 ;
        RECT 356.400 281.600 357.200 285.800 ;
        RECT 361.200 281.600 362.000 289.800 ;
        RECT 366.400 281.600 367.200 290.200 ;
        RECT 369.200 281.600 370.000 286.200 ;
        RECT 372.400 281.600 373.200 286.200 ;
        RECT 374.000 281.600 374.800 286.200 ;
        RECT 377.200 281.600 378.000 285.800 ;
        RECT 380.400 281.600 381.200 290.200 ;
        RECT 383.600 281.600 384.400 290.200 ;
        RECT 425.000 290.000 425.800 290.200 ;
        RECT 428.400 289.600 429.200 290.200 ;
        RECT 390.000 281.600 390.800 289.000 ;
        RECT 393.200 281.600 394.000 286.200 ;
        RECT 396.400 281.600 397.200 286.200 ;
        RECT 398.000 281.600 398.800 286.200 ;
        RECT 401.200 281.600 402.000 286.200 ;
        RECT 404.400 281.600 405.200 286.200 ;
        RECT 407.600 281.600 408.400 286.200 ;
        RECT 415.600 281.600 416.400 286.200 ;
        RECT 418.800 281.600 419.600 286.200 ;
        RECT 425.200 281.600 426.000 286.200 ;
        RECT 428.400 281.600 429.200 286.200 ;
        RECT 431.600 281.600 432.400 286.200 ;
        RECT 438.000 281.600 438.800 289.000 ;
        RECT 446.000 281.600 446.800 289.000 ;
        RECT 450.800 281.600 451.600 286.200 ;
        RECT 454.000 281.600 454.800 286.200 ;
        RECT 460.400 281.600 461.200 286.200 ;
        RECT 463.600 281.600 464.400 285.800 ;
        RECT 466.800 281.600 467.600 286.200 ;
        RECT 470.000 281.600 470.800 285.800 ;
        RECT 474.800 281.600 475.600 289.000 ;
        RECT 479.600 281.600 480.400 286.200 ;
        RECT 482.800 281.600 483.600 286.200 ;
        RECT 486.000 281.600 486.800 289.000 ;
        RECT 490.800 281.600 491.600 290.200 ;
        RECT 495.600 281.600 496.400 286.200 ;
        RECT 498.800 281.600 499.600 286.200 ;
        RECT 501.000 281.600 501.800 286.200 ;
        RECT 505.200 281.600 506.000 290.200 ;
        RECT 506.800 281.600 507.600 290.200 ;
        RECT 511.000 281.600 511.800 286.200 ;
        RECT 513.200 281.600 514.000 286.200 ;
        RECT 516.400 281.600 517.200 286.200 ;
        RECT 521.200 281.600 522.000 290.200 ;
        RECT 522.800 281.600 523.600 290.200 ;
        RECT 527.600 281.600 528.400 290.200 ;
        RECT 531.400 281.600 532.200 286.200 ;
        RECT 535.600 281.600 536.400 290.200 ;
        RECT 564.200 290.000 565.200 290.200 ;
        RECT 567.600 289.600 568.400 290.200 ;
        RECT 580.400 290.200 607.400 290.800 ;
        RECT 580.400 289.600 581.200 290.200 ;
        RECT 583.800 290.000 584.600 290.200 ;
        RECT 537.200 281.600 538.000 286.200 ;
        RECT 540.400 281.600 541.200 286.200 ;
        RECT 543.600 281.600 544.400 286.200 ;
        RECT 546.800 281.600 547.600 286.200 ;
        RECT 554.800 281.600 555.600 286.200 ;
        RECT 558.000 281.600 558.800 286.200 ;
        RECT 564.400 281.600 565.200 286.200 ;
        RECT 567.600 281.600 568.400 286.200 ;
        RECT 570.800 281.600 571.600 286.200 ;
        RECT 572.400 281.600 573.200 286.200 ;
        RECT 575.600 281.600 576.400 286.200 ;
        RECT 577.200 281.600 578.000 286.200 ;
        RECT 580.400 281.600 581.200 286.200 ;
        RECT 583.600 281.600 584.400 286.200 ;
        RECT 590.000 281.600 590.800 286.200 ;
        RECT 593.200 281.600 594.000 286.200 ;
        RECT 601.200 281.600 602.000 286.200 ;
        RECT 604.400 281.600 605.200 286.200 ;
        RECT 607.600 281.600 608.400 286.200 ;
        RECT 610.800 281.600 611.600 286.200 ;
        RECT 0.400 280.400 614.000 281.600 ;
        RECT 1.200 275.800 2.000 280.400 ;
        RECT 4.400 275.800 5.200 280.400 ;
        RECT 7.600 275.800 8.400 280.400 ;
        RECT 14.000 275.800 14.800 280.400 ;
        RECT 17.200 275.800 18.000 280.400 ;
        RECT 25.200 275.800 26.000 280.400 ;
        RECT 28.400 275.800 29.200 280.400 ;
        RECT 31.600 275.800 32.400 280.400 ;
        RECT 34.800 275.800 35.600 280.400 ;
        RECT 36.400 275.800 37.200 280.400 ;
        RECT 39.600 275.800 40.400 280.400 ;
        RECT 42.800 275.800 43.600 280.400 ;
        RECT 46.000 275.800 46.800 280.400 ;
        RECT 54.000 275.800 54.800 280.400 ;
        RECT 57.200 275.800 58.000 280.400 ;
        RECT 63.600 275.800 64.400 280.400 ;
        RECT 66.800 275.800 67.600 280.400 ;
        RECT 70.000 275.800 70.800 280.400 ;
        RECT 4.400 271.800 5.200 272.400 ;
        RECT 7.800 271.800 8.600 272.000 ;
        RECT 63.400 271.800 64.200 272.000 ;
        RECT 66.800 271.800 67.600 272.400 ;
        RECT 71.600 271.800 72.400 280.400 ;
        RECT 79.600 273.000 80.400 280.400 ;
        RECT 82.800 275.800 83.600 280.400 ;
        RECT 86.000 275.800 86.800 280.400 ;
        RECT 89.200 275.800 90.000 280.400 ;
        RECT 92.400 275.800 93.200 280.400 ;
        RECT 100.400 275.800 101.200 280.400 ;
        RECT 103.600 275.800 104.400 280.400 ;
        RECT 110.000 275.800 110.800 280.400 ;
        RECT 113.200 275.800 114.000 280.400 ;
        RECT 116.400 275.800 117.200 280.400 ;
        RECT 121.200 273.000 122.000 280.400 ;
        RECT 109.800 271.800 110.600 272.000 ;
        RECT 113.200 271.800 114.000 272.400 ;
        RECT 124.400 271.800 125.200 280.400 ;
        RECT 127.600 271.800 128.400 280.400 ;
        RECT 130.800 271.800 131.600 280.400 ;
        RECT 134.000 271.800 134.800 280.400 ;
        RECT 137.200 271.800 138.000 280.400 ;
        RECT 138.800 271.800 139.600 280.400 ;
        RECT 142.000 271.800 142.800 280.400 ;
        RECT 145.200 271.800 146.000 280.400 ;
        RECT 148.400 271.800 149.200 280.400 ;
        RECT 151.600 271.800 152.400 280.400 ;
        RECT 159.600 273.000 160.400 280.400 ;
        RECT 162.800 271.800 163.600 280.400 ;
        RECT 167.600 271.800 168.400 280.400 ;
        RECT 171.400 271.800 172.200 280.400 ;
        RECT 175.600 275.800 176.400 280.400 ;
        RECT 178.800 275.800 179.600 280.400 ;
        RECT 182.000 275.800 182.800 280.400 ;
        RECT 188.400 275.800 189.200 280.400 ;
        RECT 191.600 275.800 192.400 280.400 ;
        RECT 199.600 275.800 200.400 280.400 ;
        RECT 202.800 275.800 203.600 280.400 ;
        RECT 206.000 275.800 206.800 280.400 ;
        RECT 209.200 275.800 210.000 280.400 ;
        RECT 178.800 271.800 179.600 272.400 ;
        RECT 182.200 271.800 183.000 272.000 ;
        RECT 212.400 271.800 213.200 280.400 ;
        RECT 214.000 275.800 214.800 280.400 ;
        RECT 217.200 275.800 218.000 280.400 ;
        RECT 218.800 275.800 219.600 280.400 ;
        RECT 222.000 275.800 222.800 280.400 ;
        RECT 223.600 271.800 224.400 280.400 ;
        RECT 226.800 271.800 227.600 280.400 ;
        RECT 230.000 271.800 230.800 280.400 ;
        RECT 231.600 275.800 232.400 280.400 ;
        RECT 234.800 275.800 235.600 280.400 ;
        RECT 238.000 275.800 238.800 280.400 ;
        RECT 244.400 275.800 245.200 280.400 ;
        RECT 247.600 275.800 248.400 280.400 ;
        RECT 255.600 275.800 256.400 280.400 ;
        RECT 258.800 275.800 259.600 280.400 ;
        RECT 262.000 275.800 262.800 280.400 ;
        RECT 265.200 275.800 266.000 280.400 ;
        RECT 234.800 271.800 235.600 272.400 ;
        RECT 268.400 272.200 269.200 280.400 ;
        RECT 238.200 271.800 239.000 272.000 ;
        RECT 273.600 271.800 274.400 280.400 ;
        RECT 278.000 275.800 278.800 280.400 ;
        RECT 280.200 275.800 281.000 280.400 ;
        RECT 284.400 271.800 285.200 280.400 ;
        RECT 286.000 271.800 286.800 280.400 ;
        RECT 290.200 275.800 291.000 280.400 ;
        RECT 292.400 275.800 293.200 280.400 ;
        RECT 297.200 272.200 298.000 280.400 ;
        RECT 302.400 271.800 303.200 280.400 ;
        RECT 310.000 275.800 310.800 280.400 ;
        RECT 313.200 275.800 314.000 280.400 ;
        RECT 316.400 275.800 317.200 280.400 ;
        RECT 322.800 275.800 323.600 280.400 ;
        RECT 326.000 275.800 326.800 280.400 ;
        RECT 334.000 275.800 334.800 280.400 ;
        RECT 337.200 275.800 338.000 280.400 ;
        RECT 340.400 275.800 341.200 280.400 ;
        RECT 343.600 275.800 344.400 280.400 ;
        RECT 346.800 275.800 347.600 280.400 ;
        RECT 349.000 275.800 349.800 280.400 ;
        RECT 313.200 271.800 314.000 272.400 ;
        RECT 316.400 271.800 317.400 272.000 ;
        RECT 353.200 271.800 354.000 280.400 ;
        RECT 354.800 271.800 355.600 280.400 ;
        RECT 359.000 275.800 359.800 280.400 ;
        RECT 362.800 275.800 363.600 280.400 ;
        RECT 364.400 275.800 365.200 280.400 ;
        RECT 367.600 275.800 368.400 280.400 ;
        RECT 369.200 275.800 370.000 280.400 ;
        RECT 372.400 276.200 373.200 280.400 ;
        RECT 375.600 275.800 376.400 280.400 ;
        RECT 378.800 276.200 379.600 280.400 ;
        RECT 382.000 275.800 382.800 280.400 ;
        RECT 385.200 276.200 386.000 280.400 ;
        RECT 388.400 275.800 389.200 280.400 ;
        RECT 391.600 276.200 392.400 280.400 ;
        RECT 396.400 273.000 397.200 280.400 ;
        RECT 404.400 273.000 405.200 280.400 ;
        RECT 410.800 275.800 411.600 280.400 ;
        RECT 414.000 275.800 414.800 280.400 ;
        RECT 420.400 273.000 421.200 280.400 ;
        RECT 428.400 273.000 429.200 280.400 ;
        RECT 431.600 275.800 432.400 280.400 ;
        RECT 434.800 276.200 435.600 280.400 ;
        RECT 439.600 276.200 440.400 280.400 ;
        RECT 442.800 275.800 443.600 280.400 ;
        RECT 449.200 273.000 450.000 280.400 ;
        RECT 454.000 276.200 454.800 280.400 ;
        RECT 457.200 275.800 458.000 280.400 ;
        RECT 463.600 275.800 464.400 280.400 ;
        RECT 466.800 276.200 467.600 280.400 ;
        RECT 470.000 275.800 470.800 280.400 ;
        RECT 473.200 276.200 474.000 280.400 ;
        RECT 476.400 275.800 477.200 280.400 ;
        RECT 479.600 276.200 480.400 280.400 ;
        RECT 486.000 271.800 486.800 280.400 ;
        RECT 487.600 271.800 488.400 280.400 ;
        RECT 494.000 271.800 494.800 280.400 ;
        RECT 497.200 273.000 498.000 280.400 ;
        RECT 502.000 271.800 502.800 280.400 ;
        RECT 507.400 275.800 508.200 280.400 ;
        RECT 511.600 271.800 512.400 280.400 ;
        RECT 513.200 271.800 514.000 280.400 ;
        RECT 521.200 271.800 522.000 280.400 ;
        RECT 522.800 271.800 523.600 280.400 ;
        RECT 527.000 275.800 527.800 280.400 ;
        RECT 529.200 271.800 530.000 280.400 ;
        RECT 535.600 271.800 536.400 280.400 ;
        RECT 537.200 275.800 538.000 280.400 ;
        RECT 540.400 275.800 541.200 280.400 ;
        RECT 543.600 275.800 544.400 280.400 ;
        RECT 545.200 275.800 546.000 280.400 ;
        RECT 548.400 275.800 549.200 280.400 ;
        RECT 550.000 275.800 550.800 280.400 ;
        RECT 553.200 275.800 554.000 280.400 ;
        RECT 554.800 271.800 555.600 280.400 ;
        RECT 559.000 275.800 559.800 280.400 ;
        RECT 561.200 275.800 562.000 280.400 ;
        RECT 564.400 275.800 565.200 280.400 ;
        RECT 566.000 271.800 566.800 280.400 ;
        RECT 570.200 275.800 571.000 280.400 ;
        RECT 572.400 275.800 573.200 280.400 ;
        RECT 575.600 275.800 576.400 280.400 ;
        RECT 577.200 275.800 578.000 280.400 ;
        RECT 580.400 275.800 581.200 280.400 ;
        RECT 583.600 275.800 584.400 280.400 ;
        RECT 586.800 275.800 587.600 280.400 ;
        RECT 594.800 275.800 595.600 280.400 ;
        RECT 598.000 275.800 598.800 280.400 ;
        RECT 604.400 275.800 605.200 280.400 ;
        RECT 607.600 275.800 608.400 280.400 ;
        RECT 610.800 275.800 611.600 280.400 ;
        RECT 604.200 271.800 605.200 272.000 ;
        RECT 607.600 271.800 608.400 272.400 ;
        RECT 4.400 271.200 31.400 271.800 ;
        RECT 30.600 271.000 31.400 271.200 ;
        RECT 40.600 271.200 67.600 271.800 ;
        RECT 87.000 271.200 114.000 271.800 ;
        RECT 178.800 271.200 205.800 271.800 ;
        RECT 234.800 271.200 261.800 271.800 ;
        RECT 313.200 271.200 340.200 271.800 ;
        RECT 40.600 271.000 41.400 271.200 ;
        RECT 87.000 271.000 87.800 271.200 ;
        RECT 205.000 271.000 205.800 271.200 ;
        RECT 261.000 271.000 261.800 271.200 ;
        RECT 339.400 271.000 340.200 271.200 ;
        RECT 581.400 271.200 608.400 271.800 ;
        RECT 581.400 271.000 582.200 271.200 ;
        RECT 30.600 250.800 31.400 251.000 ;
        RECT 69.000 250.800 69.800 251.000 ;
        RECT 4.400 250.200 31.400 250.800 ;
        RECT 42.800 250.200 69.800 250.800 ;
        RECT 98.200 250.800 99.000 251.000 ;
        RECT 147.800 250.800 148.600 251.000 ;
        RECT 224.200 250.800 225.000 251.000 ;
        RECT 98.200 250.200 125.200 250.800 ;
        RECT 147.800 250.200 174.800 250.800 ;
        RECT 198.000 250.200 225.000 250.800 ;
        RECT 253.400 250.800 254.200 251.000 ;
        RECT 381.000 250.800 381.800 251.000 ;
        RECT 253.400 250.200 280.400 250.800 ;
        RECT 354.800 250.200 381.800 250.800 ;
        RECT 573.400 250.800 574.200 251.000 ;
        RECT 573.400 250.200 600.400 250.800 ;
        RECT 4.400 249.600 5.200 250.200 ;
        RECT 7.800 250.000 8.600 250.200 ;
        RECT 42.800 249.600 43.600 250.200 ;
        RECT 46.000 250.000 47.000 250.200 ;
        RECT 1.200 241.600 2.000 246.200 ;
        RECT 4.400 241.600 5.200 246.200 ;
        RECT 7.600 241.600 8.400 246.200 ;
        RECT 14.000 241.600 14.800 246.200 ;
        RECT 17.200 241.600 18.000 246.200 ;
        RECT 25.200 241.600 26.000 246.200 ;
        RECT 28.400 241.600 29.200 246.200 ;
        RECT 31.600 241.600 32.400 246.200 ;
        RECT 34.800 241.600 35.600 246.200 ;
        RECT 38.000 241.600 38.800 246.200 ;
        RECT 39.600 241.600 40.400 246.200 ;
        RECT 42.800 241.600 43.600 246.200 ;
        RECT 46.000 241.600 46.800 246.200 ;
        RECT 52.400 241.600 53.200 246.200 ;
        RECT 55.600 241.600 56.400 246.200 ;
        RECT 63.600 241.600 64.400 246.200 ;
        RECT 66.800 241.600 67.600 246.200 ;
        RECT 70.000 241.600 70.800 246.200 ;
        RECT 73.200 241.600 74.000 246.200 ;
        RECT 74.800 241.600 75.600 250.200 ;
        RECT 82.800 241.600 83.600 249.000 ;
        RECT 87.600 241.600 88.400 246.200 ;
        RECT 92.400 241.600 93.200 250.200 ;
        RECT 121.000 250.000 122.000 250.200 ;
        RECT 124.400 249.600 125.200 250.200 ;
        RECT 94.000 241.600 94.800 246.200 ;
        RECT 97.200 241.600 98.000 246.200 ;
        RECT 100.400 241.600 101.200 246.200 ;
        RECT 103.600 241.600 104.400 246.200 ;
        RECT 111.600 241.600 112.400 246.200 ;
        RECT 114.800 241.600 115.600 246.200 ;
        RECT 121.200 241.600 122.000 246.200 ;
        RECT 124.400 241.600 125.200 246.200 ;
        RECT 127.600 241.600 128.400 246.200 ;
        RECT 130.800 241.600 131.600 246.200 ;
        RECT 132.400 241.600 133.200 250.200 ;
        RECT 170.600 250.000 171.600 250.200 ;
        RECT 174.000 249.600 174.800 250.200 ;
        RECT 135.600 241.600 136.400 249.000 ;
        RECT 143.600 241.600 144.400 246.200 ;
        RECT 146.800 241.600 147.600 246.200 ;
        RECT 150.000 241.600 150.800 246.200 ;
        RECT 153.200 241.600 154.000 246.200 ;
        RECT 161.200 241.600 162.000 246.200 ;
        RECT 164.400 241.600 165.200 246.200 ;
        RECT 170.800 241.600 171.600 246.200 ;
        RECT 174.000 241.600 174.800 246.200 ;
        RECT 177.200 241.600 178.000 246.200 ;
        RECT 178.800 241.600 179.600 246.200 ;
        RECT 182.000 241.600 182.800 246.200 ;
        RECT 184.200 241.600 185.000 246.200 ;
        RECT 188.400 241.600 189.200 250.200 ;
        RECT 190.000 241.600 190.800 250.200 ;
        RECT 193.200 241.600 194.000 250.200 ;
        RECT 198.000 249.600 198.800 250.200 ;
        RECT 201.200 250.000 202.200 250.200 ;
        RECT 194.800 241.600 195.600 246.200 ;
        RECT 198.000 241.600 198.800 246.200 ;
        RECT 201.200 241.600 202.000 246.200 ;
        RECT 207.600 241.600 208.400 246.200 ;
        RECT 210.800 241.600 211.600 246.200 ;
        RECT 218.800 241.600 219.600 246.200 ;
        RECT 222.000 241.600 222.800 246.200 ;
        RECT 225.200 241.600 226.000 246.200 ;
        RECT 228.400 241.600 229.200 246.200 ;
        RECT 230.000 241.600 230.800 246.200 ;
        RECT 234.400 241.600 235.200 250.200 ;
        RECT 239.600 241.600 240.400 249.800 ;
        RECT 242.800 241.600 243.600 250.200 ;
        RECT 276.200 250.000 277.000 250.200 ;
        RECT 279.600 249.600 280.400 250.200 ;
        RECT 246.000 241.600 246.800 249.000 ;
        RECT 249.200 241.600 250.000 246.200 ;
        RECT 252.400 241.600 253.200 246.200 ;
        RECT 255.600 241.600 256.400 246.200 ;
        RECT 258.800 241.600 259.600 246.200 ;
        RECT 266.800 241.600 267.600 246.200 ;
        RECT 270.000 241.600 270.800 246.200 ;
        RECT 276.400 241.600 277.200 246.200 ;
        RECT 279.600 241.600 280.400 246.200 ;
        RECT 282.800 241.600 283.600 246.200 ;
        RECT 284.400 241.600 285.200 250.200 ;
        RECT 290.800 241.600 291.600 250.200 ;
        RECT 293.000 241.600 293.800 246.200 ;
        RECT 297.200 241.600 298.000 250.200 ;
        RECT 298.800 241.600 299.600 246.200 ;
        RECT 302.000 241.600 302.800 246.200 ;
        RECT 311.000 241.600 311.800 250.200 ;
        RECT 314.800 241.600 315.600 250.200 ;
        RECT 318.000 241.600 318.800 249.000 ;
        RECT 321.800 241.600 322.600 246.200 ;
        RECT 326.000 241.600 326.800 250.200 ;
        RECT 327.600 241.600 328.400 250.200 ;
        RECT 334.000 241.600 334.800 250.200 ;
        RECT 354.800 249.600 355.600 250.200 ;
        RECT 358.000 250.000 359.000 250.200 ;
        RECT 335.600 241.600 336.400 246.200 ;
        RECT 338.800 241.600 339.600 246.200 ;
        RECT 340.400 241.600 341.200 246.200 ;
        RECT 343.600 241.600 344.400 245.800 ;
        RECT 348.400 241.600 349.200 249.000 ;
        RECT 351.600 241.600 352.400 246.200 ;
        RECT 354.800 241.600 355.600 246.200 ;
        RECT 358.000 241.600 358.800 246.200 ;
        RECT 364.400 241.600 365.200 246.200 ;
        RECT 367.600 241.600 368.400 246.200 ;
        RECT 375.600 241.600 376.400 246.200 ;
        RECT 378.800 241.600 379.600 246.200 ;
        RECT 382.000 241.600 382.800 246.200 ;
        RECT 385.200 241.600 386.000 246.200 ;
        RECT 388.400 241.600 389.200 246.200 ;
        RECT 390.000 241.600 390.800 246.200 ;
        RECT 393.200 241.600 394.000 245.800 ;
        RECT 401.200 241.600 402.000 249.000 ;
        RECT 409.200 241.600 410.000 249.000 ;
        RECT 412.400 241.600 413.200 246.200 ;
        RECT 415.600 241.600 416.400 246.200 ;
        RECT 417.200 241.600 418.000 246.200 ;
        RECT 420.400 241.600 421.200 245.800 ;
        RECT 423.600 241.600 424.400 246.200 ;
        RECT 426.800 241.600 427.600 246.200 ;
        RECT 430.000 241.600 430.800 249.000 ;
        RECT 436.400 241.600 437.200 246.200 ;
        RECT 439.600 241.600 440.400 246.200 ;
        RECT 441.200 241.600 442.000 246.200 ;
        RECT 444.400 241.600 445.200 246.200 ;
        RECT 446.000 241.600 446.800 246.200 ;
        RECT 449.200 241.600 450.000 245.800 ;
        RECT 457.200 241.600 458.000 249.000 ;
        RECT 470.000 241.600 470.800 249.000 ;
        RECT 473.200 241.600 474.000 246.200 ;
        RECT 476.400 241.600 477.200 245.800 ;
        RECT 479.600 241.600 480.400 250.200 ;
        RECT 487.600 241.600 488.400 250.200 ;
        RECT 490.800 241.600 491.600 246.200 ;
        RECT 494.000 241.600 494.800 246.200 ;
        RECT 497.200 241.600 498.000 249.000 ;
        RECT 502.000 241.600 502.800 246.200 ;
        RECT 505.200 241.600 506.000 246.200 ;
        RECT 508.400 241.600 509.200 245.800 ;
        RECT 511.600 241.600 512.400 246.200 ;
        RECT 516.400 241.600 517.200 250.200 ;
        RECT 518.000 241.600 518.800 250.200 ;
        RECT 524.400 241.600 525.200 250.200 ;
        RECT 526.000 241.600 526.800 250.200 ;
        RECT 532.400 241.600 533.200 250.200 ;
        RECT 534.000 241.600 534.800 246.200 ;
        RECT 537.200 241.600 538.000 250.200 ;
        RECT 543.600 241.600 544.400 250.200 ;
        RECT 545.200 241.600 546.000 250.200 ;
        RECT 548.400 241.600 549.200 250.200 ;
        RECT 552.600 241.600 553.400 246.200 ;
        RECT 554.800 241.600 555.600 250.200 ;
        RECT 558.000 241.600 558.800 250.200 ;
        RECT 561.200 241.600 562.000 250.200 ;
        RECT 564.400 241.600 565.200 250.200 ;
        RECT 567.600 241.600 568.400 250.200 ;
        RECT 596.200 250.000 597.200 250.200 ;
        RECT 599.600 249.600 600.400 250.200 ;
        RECT 569.200 241.600 570.000 246.200 ;
        RECT 572.400 241.600 573.200 246.200 ;
        RECT 575.600 241.600 576.400 246.200 ;
        RECT 578.800 241.600 579.600 246.200 ;
        RECT 586.800 241.600 587.600 246.200 ;
        RECT 590.000 241.600 590.800 246.200 ;
        RECT 596.400 241.600 597.200 246.200 ;
        RECT 599.600 241.600 600.400 246.200 ;
        RECT 602.800 241.600 603.600 246.200 ;
        RECT 606.000 241.600 606.800 249.000 ;
        RECT 0.400 240.400 614.000 241.600 ;
        RECT 1.200 235.800 2.000 240.400 ;
        RECT 4.400 235.800 5.200 240.400 ;
        RECT 7.600 231.800 8.400 240.400 ;
        RECT 11.800 235.800 12.600 240.400 ;
        RECT 14.000 231.800 14.800 240.400 ;
        RECT 18.200 235.800 19.000 240.400 ;
        RECT 20.400 231.800 21.200 240.400 ;
        RECT 24.600 235.800 25.400 240.400 ;
        RECT 26.800 235.800 27.600 240.400 ;
        RECT 30.000 235.800 30.800 240.400 ;
        RECT 31.600 231.800 32.400 240.400 ;
        RECT 35.800 235.800 36.600 240.400 ;
        RECT 39.600 235.800 40.400 240.400 ;
        RECT 41.200 235.800 42.000 240.400 ;
        RECT 44.400 235.800 45.200 240.400 ;
        RECT 47.600 235.800 48.400 240.400 ;
        RECT 50.800 235.800 51.600 240.400 ;
        RECT 57.200 235.800 58.000 240.400 ;
        RECT 60.400 235.800 61.200 240.400 ;
        RECT 68.400 235.800 69.200 240.400 ;
        RECT 71.600 235.800 72.400 240.400 ;
        RECT 74.800 235.800 75.600 240.400 ;
        RECT 78.000 235.800 78.800 240.400 ;
        RECT 79.600 235.800 80.400 240.400 ;
        RECT 82.800 235.800 83.600 240.400 ;
        RECT 47.600 231.800 48.400 232.400 ;
        RECT 51.000 231.800 51.800 232.000 ;
        RECT 84.400 231.800 85.200 240.400 ;
        RECT 87.600 231.800 88.400 240.400 ;
        RECT 90.800 231.800 91.600 240.400 ;
        RECT 94.000 231.800 94.800 240.400 ;
        RECT 97.200 231.800 98.000 240.400 ;
        RECT 100.400 233.000 101.200 240.400 ;
        RECT 103.600 231.800 104.400 240.400 ;
        RECT 106.800 232.000 107.600 240.400 ;
        RECT 112.400 235.800 113.200 240.400 ;
        RECT 115.600 235.800 116.400 240.400 ;
        RECT 121.200 231.800 122.000 240.400 ;
        RECT 125.000 235.800 125.800 240.400 ;
        RECT 129.200 231.800 130.000 240.400 ;
        RECT 134.000 231.800 134.800 240.400 ;
        RECT 135.600 231.800 136.400 240.400 ;
        RECT 139.800 235.800 140.600 240.400 ;
        RECT 143.600 235.800 144.400 240.400 ;
        RECT 150.000 235.800 150.800 240.400 ;
        RECT 153.200 235.800 154.000 240.400 ;
        RECT 156.400 235.800 157.200 240.400 ;
        RECT 162.800 235.800 163.600 240.400 ;
        RECT 166.000 235.800 166.800 240.400 ;
        RECT 174.000 235.800 174.800 240.400 ;
        RECT 177.200 235.800 178.000 240.400 ;
        RECT 180.400 235.800 181.200 240.400 ;
        RECT 183.600 235.800 184.400 240.400 ;
        RECT 185.200 235.800 186.000 240.400 ;
        RECT 188.400 235.800 189.200 240.400 ;
        RECT 191.600 235.800 192.400 240.400 ;
        RECT 194.800 235.800 195.600 240.400 ;
        RECT 201.200 235.800 202.000 240.400 ;
        RECT 204.400 235.800 205.200 240.400 ;
        RECT 212.400 235.800 213.200 240.400 ;
        RECT 215.600 235.800 216.400 240.400 ;
        RECT 218.800 235.800 219.600 240.400 ;
        RECT 222.000 235.800 222.800 240.400 ;
        RECT 153.200 231.800 154.000 232.400 ;
        RECT 156.400 231.800 157.400 232.000 ;
        RECT 191.600 231.800 192.400 232.400 ;
        RECT 195.000 231.800 195.800 232.000 ;
        RECT 223.600 231.800 224.400 240.400 ;
        RECT 226.800 231.800 227.600 240.400 ;
        RECT 230.000 231.800 230.800 240.400 ;
        RECT 231.600 235.800 232.400 240.400 ;
        RECT 234.800 235.800 235.600 240.400 ;
        RECT 238.000 235.800 238.800 240.400 ;
        RECT 244.400 235.800 245.200 240.400 ;
        RECT 247.600 235.800 248.400 240.400 ;
        RECT 255.600 235.800 256.400 240.400 ;
        RECT 258.800 235.800 259.600 240.400 ;
        RECT 262.000 235.800 262.800 240.400 ;
        RECT 265.200 235.800 266.000 240.400 ;
        RECT 266.800 235.800 267.600 240.400 ;
        RECT 270.000 235.800 270.800 240.400 ;
        RECT 271.600 235.800 272.400 240.400 ;
        RECT 274.800 235.800 275.600 240.400 ;
        RECT 234.800 231.800 235.600 232.400 ;
        RECT 238.200 231.800 239.000 232.000 ;
        RECT 276.400 231.800 277.200 240.400 ;
        RECT 280.200 235.800 281.000 240.400 ;
        RECT 284.400 231.800 285.200 240.400 ;
        RECT 287.600 235.800 288.400 240.400 ;
        RECT 289.800 235.800 290.600 240.400 ;
        RECT 294.000 231.800 294.800 240.400 ;
        RECT 295.600 231.800 296.400 240.400 ;
        RECT 299.800 235.800 300.600 240.400 ;
        RECT 302.000 235.800 302.800 240.400 ;
        RECT 305.200 235.800 306.000 240.400 ;
        RECT 311.600 231.800 312.400 240.400 ;
        RECT 315.800 235.800 316.600 240.400 ;
        RECT 318.000 235.800 318.800 240.400 ;
        RECT 321.200 236.200 322.000 240.400 ;
        RECT 324.400 231.800 325.200 240.400 ;
        RECT 327.600 231.800 328.400 240.400 ;
        RECT 330.800 231.800 331.600 240.400 ;
        RECT 334.000 231.800 334.800 240.400 ;
        RECT 337.200 231.800 338.000 240.400 ;
        RECT 338.800 235.800 339.600 240.400 ;
        RECT 342.000 236.200 342.800 240.400 ;
        RECT 345.200 235.800 346.000 240.400 ;
        RECT 348.400 236.200 349.200 240.400 ;
        RECT 351.600 235.800 352.400 240.400 ;
        RECT 354.800 236.200 355.600 240.400 ;
        RECT 359.600 232.200 360.400 240.400 ;
        RECT 364.800 231.800 365.600 240.400 ;
        RECT 367.600 235.800 368.400 240.400 ;
        RECT 370.800 235.800 371.600 240.400 ;
        RECT 374.000 235.800 374.800 240.400 ;
        RECT 380.400 235.800 381.200 240.400 ;
        RECT 383.600 235.800 384.400 240.400 ;
        RECT 391.600 235.800 392.400 240.400 ;
        RECT 394.800 235.800 395.600 240.400 ;
        RECT 398.000 235.800 398.800 240.400 ;
        RECT 401.200 235.800 402.000 240.400 ;
        RECT 404.400 235.800 405.200 240.400 ;
        RECT 406.000 235.800 406.800 240.400 ;
        RECT 409.200 235.800 410.000 240.400 ;
        RECT 412.400 233.000 413.200 240.400 ;
        RECT 370.800 231.800 371.600 232.400 ;
        RECT 374.000 231.800 375.000 232.000 ;
        RECT 415.600 231.800 416.400 240.400 ;
        RECT 417.200 231.800 418.000 240.400 ;
        RECT 420.400 231.800 421.200 240.400 ;
        RECT 423.600 231.800 424.400 240.400 ;
        RECT 426.800 231.800 427.600 240.400 ;
        RECT 430.000 231.800 430.800 240.400 ;
        RECT 431.600 231.800 432.400 240.400 ;
        RECT 434.800 231.800 435.600 240.400 ;
        RECT 438.000 231.800 438.800 240.400 ;
        RECT 441.200 231.800 442.000 240.400 ;
        RECT 444.400 231.800 445.200 240.400 ;
        RECT 447.600 233.000 448.400 240.400 ;
        RECT 458.800 233.000 459.600 240.400 ;
        RECT 466.800 235.800 467.600 240.400 ;
        RECT 470.000 235.800 470.800 240.400 ;
        RECT 471.600 235.800 472.400 240.400 ;
        RECT 474.800 236.200 475.600 240.400 ;
        RECT 478.000 235.800 478.800 240.400 ;
        RECT 481.200 235.800 482.000 240.400 ;
        RECT 484.400 233.000 485.200 240.400 ;
        RECT 492.400 236.200 493.200 240.400 ;
        RECT 495.600 235.800 496.400 240.400 ;
        RECT 500.400 233.000 501.200 240.400 ;
        RECT 505.200 236.200 506.000 240.400 ;
        RECT 508.400 235.800 509.200 240.400 ;
        RECT 511.600 236.200 512.400 240.400 ;
        RECT 514.800 235.800 515.600 240.400 ;
        RECT 516.400 235.800 517.200 240.400 ;
        RECT 519.600 236.200 520.400 240.400 ;
        RECT 522.800 235.800 523.600 240.400 ;
        RECT 526.000 236.200 526.800 240.400 ;
        RECT 529.200 235.800 530.000 240.400 ;
        RECT 532.400 236.200 533.200 240.400 ;
        RECT 537.200 236.200 538.000 240.400 ;
        RECT 540.400 235.800 541.200 240.400 ;
        RECT 543.600 236.200 544.400 240.400 ;
        RECT 546.800 235.800 547.600 240.400 ;
        RECT 548.400 235.800 549.200 240.400 ;
        RECT 551.600 235.800 552.400 240.400 ;
        RECT 553.200 231.800 554.000 240.400 ;
        RECT 556.400 235.800 557.200 240.400 ;
        RECT 559.600 236.200 560.400 240.400 ;
        RECT 562.800 235.800 563.600 240.400 ;
        RECT 566.000 235.800 566.800 240.400 ;
        RECT 567.600 235.800 568.400 240.400 ;
        RECT 570.800 235.800 571.600 240.400 ;
        RECT 574.000 235.800 574.800 240.400 ;
        RECT 577.200 235.800 578.000 240.400 ;
        RECT 585.200 235.800 586.000 240.400 ;
        RECT 588.400 235.800 589.200 240.400 ;
        RECT 594.800 235.800 595.600 240.400 ;
        RECT 598.000 235.800 598.800 240.400 ;
        RECT 601.200 235.800 602.000 240.400 ;
        RECT 594.600 231.800 595.400 232.000 ;
        RECT 598.000 231.800 598.800 232.400 ;
        RECT 602.800 231.800 603.600 240.400 ;
        RECT 607.000 235.800 607.800 240.400 ;
        RECT 47.600 231.200 74.600 231.800 ;
        RECT 153.200 231.200 180.200 231.800 ;
        RECT 191.600 231.200 218.600 231.800 ;
        RECT 234.800 231.200 261.800 231.800 ;
        RECT 370.800 231.200 397.800 231.800 ;
        RECT 73.800 231.000 74.600 231.200 ;
        RECT 179.400 231.000 180.200 231.200 ;
        RECT 217.800 231.000 218.600 231.200 ;
        RECT 261.000 231.000 261.800 231.200 ;
        RECT 397.000 231.000 397.800 231.200 ;
        RECT 571.800 231.200 598.800 231.800 ;
        RECT 571.800 231.000 572.600 231.200 ;
        RECT 181.400 210.800 182.200 211.000 ;
        RECT 241.800 210.800 242.600 211.000 ;
        RECT 280.200 210.800 281.000 211.000 ;
        RECT 181.400 210.200 208.400 210.800 ;
        RECT 1.200 201.600 2.000 206.200 ;
        RECT 4.400 201.600 5.200 210.200 ;
        RECT 8.600 201.600 9.400 206.200 ;
        RECT 13.000 201.600 13.800 210.200 ;
        RECT 17.200 201.600 18.000 210.200 ;
        RECT 21.400 201.600 22.200 206.200 ;
        RECT 23.600 201.600 24.400 206.200 ;
        RECT 26.800 201.600 27.600 206.200 ;
        RECT 29.000 201.600 29.800 206.200 ;
        RECT 33.200 201.600 34.000 210.200 ;
        RECT 35.400 201.600 36.200 206.200 ;
        RECT 39.600 201.600 40.400 210.200 ;
        RECT 41.200 201.600 42.000 210.200 ;
        RECT 44.400 201.600 45.200 210.200 ;
        RECT 47.600 201.600 48.400 210.200 ;
        RECT 50.800 201.600 51.600 210.200 ;
        RECT 54.000 201.600 54.800 210.200 ;
        RECT 55.600 201.600 56.400 210.200 ;
        RECT 58.800 201.600 59.600 210.200 ;
        RECT 62.000 201.600 62.800 210.200 ;
        RECT 65.200 201.600 66.000 210.200 ;
        RECT 68.400 201.600 69.200 210.200 ;
        RECT 71.200 201.600 72.000 210.200 ;
        RECT 76.400 201.600 77.200 209.800 ;
        RECT 81.200 201.600 82.000 210.200 ;
        RECT 86.800 201.600 87.600 206.200 ;
        RECT 90.000 201.600 90.800 206.200 ;
        RECT 95.600 201.600 96.400 210.000 ;
        RECT 98.800 201.600 99.600 210.200 ;
        RECT 103.000 201.600 103.800 206.200 ;
        RECT 105.800 201.600 106.600 206.200 ;
        RECT 110.000 201.600 110.800 210.200 ;
        RECT 111.600 201.600 112.400 210.200 ;
        RECT 115.800 201.600 116.600 206.200 ;
        RECT 118.600 201.600 119.400 206.200 ;
        RECT 122.800 201.600 123.600 210.200 ;
        RECT 124.400 201.600 125.200 210.200 ;
        RECT 128.600 201.600 129.400 206.200 ;
        RECT 131.400 201.600 132.200 206.200 ;
        RECT 135.600 201.600 136.400 210.200 ;
        RECT 138.800 201.600 139.600 210.200 ;
        RECT 144.400 201.600 145.200 206.200 ;
        RECT 147.600 201.600 148.400 206.200 ;
        RECT 153.200 201.600 154.000 210.000 ;
        RECT 161.200 201.600 162.000 210.200 ;
        RECT 204.200 210.000 205.000 210.200 ;
        RECT 207.600 209.600 208.400 210.200 ;
        RECT 215.600 210.200 242.600 210.800 ;
        RECT 254.000 210.200 281.000 210.800 ;
        RECT 312.600 210.800 313.400 211.000 ;
        RECT 354.200 210.800 355.000 211.000 ;
        RECT 429.400 210.800 430.200 211.000 ;
        RECT 517.000 210.800 517.800 211.000 ;
        RECT 312.600 210.200 339.600 210.800 ;
        RECT 354.200 210.200 381.200 210.800 ;
        RECT 429.400 210.200 456.400 210.800 ;
        RECT 215.600 209.600 216.400 210.200 ;
        RECT 219.000 210.000 219.800 210.200 ;
        RECT 254.000 209.600 254.800 210.200 ;
        RECT 257.200 210.000 258.200 210.200 ;
        RECT 167.600 201.600 168.600 208.800 ;
        RECT 173.800 202.200 174.800 208.800 ;
        RECT 173.800 201.600 174.600 202.200 ;
        RECT 177.200 201.600 178.000 206.200 ;
        RECT 180.400 201.600 181.200 206.200 ;
        RECT 183.600 201.600 184.400 206.200 ;
        RECT 186.800 201.600 187.600 206.200 ;
        RECT 194.800 201.600 195.600 206.200 ;
        RECT 198.000 201.600 198.800 206.200 ;
        RECT 204.400 201.600 205.200 206.200 ;
        RECT 207.600 201.600 208.400 206.200 ;
        RECT 210.800 201.600 211.600 206.200 ;
        RECT 212.400 201.600 213.200 206.200 ;
        RECT 215.600 201.600 216.400 206.200 ;
        RECT 218.800 201.600 219.600 206.200 ;
        RECT 225.200 201.600 226.000 206.200 ;
        RECT 228.400 201.600 229.200 206.200 ;
        RECT 236.400 201.600 237.200 206.200 ;
        RECT 239.600 201.600 240.400 206.200 ;
        RECT 242.800 201.600 243.600 206.200 ;
        RECT 246.000 201.600 246.800 206.200 ;
        RECT 247.600 201.600 248.400 206.200 ;
        RECT 250.800 201.600 251.600 206.200 ;
        RECT 254.000 201.600 254.800 206.200 ;
        RECT 257.200 201.600 258.000 206.200 ;
        RECT 263.600 201.600 264.400 206.200 ;
        RECT 266.800 201.600 267.600 206.200 ;
        RECT 274.800 201.600 275.600 206.200 ;
        RECT 278.000 201.600 278.800 206.200 ;
        RECT 281.200 201.600 282.000 206.200 ;
        RECT 284.400 201.600 285.200 206.200 ;
        RECT 287.600 201.600 288.400 206.200 ;
        RECT 289.200 201.600 290.000 210.200 ;
        RECT 292.400 201.600 293.200 210.200 ;
        RECT 295.600 201.600 296.400 210.200 ;
        RECT 298.800 201.600 299.600 210.200 ;
        RECT 302.000 201.600 302.800 210.200 ;
        RECT 335.400 210.000 336.200 210.200 ;
        RECT 338.800 209.600 339.600 210.200 ;
        RECT 308.400 201.600 309.200 206.200 ;
        RECT 311.600 201.600 312.400 206.200 ;
        RECT 314.800 201.600 315.600 206.200 ;
        RECT 318.000 201.600 318.800 206.200 ;
        RECT 326.000 201.600 326.800 206.200 ;
        RECT 329.200 201.600 330.000 206.200 ;
        RECT 335.600 201.600 336.400 206.200 ;
        RECT 338.800 201.600 339.600 206.200 ;
        RECT 342.000 201.600 342.800 206.200 ;
        RECT 343.600 201.600 344.400 210.200 ;
        RECT 377.000 210.000 378.000 210.200 ;
        RECT 380.400 209.600 381.200 210.200 ;
        RECT 347.800 201.600 348.600 206.200 ;
        RECT 350.000 201.600 350.800 206.200 ;
        RECT 353.200 201.600 354.000 206.200 ;
        RECT 356.400 201.600 357.200 206.200 ;
        RECT 359.600 201.600 360.400 206.200 ;
        RECT 367.600 201.600 368.400 206.200 ;
        RECT 370.800 201.600 371.600 206.200 ;
        RECT 377.200 201.600 378.000 206.200 ;
        RECT 380.400 201.600 381.200 206.200 ;
        RECT 383.600 201.600 384.400 206.200 ;
        RECT 385.200 201.600 386.000 206.200 ;
        RECT 388.400 201.600 389.200 206.200 ;
        RECT 390.000 201.600 390.800 210.200 ;
        RECT 393.200 201.600 394.000 210.200 ;
        RECT 396.400 201.600 397.200 210.200 ;
        RECT 399.600 201.600 400.400 209.000 ;
        RECT 402.800 201.600 403.600 210.200 ;
        RECT 404.400 201.600 405.200 210.200 ;
        RECT 408.600 201.600 409.400 206.200 ;
        RECT 410.800 201.600 411.600 206.200 ;
        RECT 415.600 201.600 416.400 209.000 ;
        RECT 418.800 201.600 419.600 210.200 ;
        RECT 452.200 210.000 453.200 210.200 ;
        RECT 455.600 209.600 456.400 210.200 ;
        RECT 490.800 210.200 517.800 210.800 ;
        RECT 541.400 210.800 542.200 211.000 ;
        RECT 541.400 210.200 568.400 210.800 ;
        RECT 420.400 201.600 421.200 206.200 ;
        RECT 423.600 201.600 424.400 206.200 ;
        RECT 425.200 201.600 426.000 206.200 ;
        RECT 428.400 201.600 429.200 206.200 ;
        RECT 431.600 201.600 432.400 206.200 ;
        RECT 434.800 201.600 435.600 206.200 ;
        RECT 442.800 201.600 443.600 206.200 ;
        RECT 446.000 201.600 446.800 206.200 ;
        RECT 452.400 201.600 453.200 206.200 ;
        RECT 455.600 201.600 456.400 206.200 ;
        RECT 458.800 201.600 459.600 206.200 ;
        RECT 465.200 201.600 466.000 206.200 ;
        RECT 468.400 201.600 469.200 206.200 ;
        RECT 471.600 201.600 472.400 206.200 ;
        RECT 474.800 201.600 475.600 206.200 ;
        RECT 478.000 201.600 478.800 206.200 ;
        RECT 482.800 201.600 483.600 209.800 ;
        RECT 490.800 209.600 491.600 210.200 ;
        RECT 494.000 210.000 495.000 210.200 ;
        RECT 486.000 201.600 486.800 206.200 ;
        RECT 487.600 201.600 488.400 206.200 ;
        RECT 490.800 201.600 491.600 206.200 ;
        RECT 494.000 201.600 494.800 206.200 ;
        RECT 500.400 201.600 501.200 206.200 ;
        RECT 503.600 201.600 504.400 206.200 ;
        RECT 511.600 201.600 512.400 206.200 ;
        RECT 514.800 201.600 515.600 206.200 ;
        RECT 518.000 201.600 518.800 206.200 ;
        RECT 521.200 201.600 522.000 206.200 ;
        RECT 522.800 201.600 523.600 206.200 ;
        RECT 526.000 201.600 526.800 210.200 ;
        RECT 564.200 210.000 565.200 210.200 ;
        RECT 567.600 209.600 568.400 210.200 ;
        RECT 530.200 201.600 531.000 206.200 ;
        RECT 532.400 201.600 533.200 206.200 ;
        RECT 535.600 201.600 536.400 206.200 ;
        RECT 537.200 201.600 538.000 206.200 ;
        RECT 540.400 201.600 541.200 206.200 ;
        RECT 543.600 201.600 544.400 206.200 ;
        RECT 546.800 201.600 547.600 206.200 ;
        RECT 554.800 201.600 555.600 206.200 ;
        RECT 558.000 201.600 558.800 206.200 ;
        RECT 564.400 201.600 565.200 206.200 ;
        RECT 567.600 201.600 568.400 206.200 ;
        RECT 570.800 201.600 571.600 206.200 ;
        RECT 572.400 201.600 573.200 210.200 ;
        RECT 576.600 201.600 577.400 206.200 ;
        RECT 578.800 201.600 579.600 210.200 ;
        RECT 582.000 201.600 582.800 210.200 ;
        RECT 585.200 201.600 586.000 210.200 ;
        RECT 588.400 201.600 589.200 210.200 ;
        RECT 591.600 201.600 592.400 210.200 ;
        RECT 593.200 201.600 594.000 210.200 ;
        RECT 596.400 201.600 597.200 210.200 ;
        RECT 599.600 201.600 600.400 210.200 ;
        RECT 602.800 201.600 603.600 210.200 ;
        RECT 606.000 201.600 606.800 210.200 ;
        RECT 0.400 200.400 614.000 201.600 ;
        RECT 1.200 195.800 2.000 200.400 ;
        RECT 4.400 195.800 5.200 200.400 ;
        RECT 7.600 195.800 8.400 200.400 ;
        RECT 14.000 195.800 14.800 200.400 ;
        RECT 17.200 195.800 18.000 200.400 ;
        RECT 25.200 195.800 26.000 200.400 ;
        RECT 28.400 195.800 29.200 200.400 ;
        RECT 31.600 195.800 32.400 200.400 ;
        RECT 34.800 195.800 35.600 200.400 ;
        RECT 38.000 195.800 38.800 200.400 ;
        RECT 4.400 191.800 5.200 192.400 ;
        RECT 41.200 192.000 42.000 200.400 ;
        RECT 46.800 195.800 47.600 200.400 ;
        RECT 50.000 195.800 50.800 200.400 ;
        RECT 7.800 191.800 8.600 192.000 ;
        RECT 55.600 191.800 56.400 200.400 ;
        RECT 59.400 195.800 60.200 200.400 ;
        RECT 63.600 191.800 64.400 200.400 ;
        RECT 65.200 191.800 66.000 200.400 ;
        RECT 69.400 195.800 70.200 200.400 ;
        RECT 72.800 191.800 73.600 200.400 ;
        RECT 78.000 192.200 78.800 200.400 ;
        RECT 81.200 191.800 82.000 200.400 ;
        RECT 84.400 193.000 85.200 200.400 ;
        RECT 89.200 192.000 90.000 200.400 ;
        RECT 94.800 195.800 95.600 200.400 ;
        RECT 98.000 195.800 98.800 200.400 ;
        RECT 103.600 191.800 104.400 200.400 ;
        RECT 106.800 191.800 107.600 200.400 ;
        RECT 111.000 195.800 111.800 200.400 ;
        RECT 114.800 192.200 115.600 200.400 ;
        RECT 120.000 191.800 120.800 200.400 ;
        RECT 123.400 195.800 124.200 200.400 ;
        RECT 127.600 191.800 128.400 200.400 ;
        RECT 130.800 192.200 131.600 200.400 ;
        RECT 136.000 191.800 136.800 200.400 ;
        RECT 140.400 193.000 141.200 200.400 ;
        RECT 143.600 191.800 144.400 200.400 ;
        RECT 146.800 195.800 147.600 200.400 ;
        RECT 148.400 191.800 149.200 200.400 ;
        RECT 159.600 195.800 160.400 200.400 ;
        RECT 163.000 199.800 163.800 200.400 ;
        RECT 162.800 193.200 163.800 199.800 ;
        RECT 169.000 193.200 170.000 200.400 ;
        RECT 172.400 195.800 173.200 200.400 ;
        RECT 175.600 195.800 176.400 200.400 ;
        RECT 178.800 195.800 179.600 200.400 ;
        RECT 182.000 195.800 182.800 200.400 ;
        RECT 190.000 195.800 190.800 200.400 ;
        RECT 193.200 195.800 194.000 200.400 ;
        RECT 199.600 195.800 200.400 200.400 ;
        RECT 202.800 195.800 203.600 200.400 ;
        RECT 206.000 195.800 206.800 200.400 ;
        RECT 207.600 195.800 208.400 200.400 ;
        RECT 210.800 195.800 211.600 200.400 ;
        RECT 199.400 191.800 200.200 192.000 ;
        RECT 202.800 191.800 203.600 192.400 ;
        RECT 212.400 191.800 213.200 200.400 ;
        RECT 216.600 195.800 217.400 200.400 ;
        RECT 220.400 193.000 221.200 200.400 ;
        RECT 223.600 191.800 224.400 200.400 ;
        RECT 226.800 191.800 227.600 200.400 ;
        RECT 230.000 191.800 230.800 200.400 ;
        RECT 231.600 191.800 232.400 200.400 ;
        RECT 235.800 195.800 236.600 200.400 ;
        RECT 238.000 191.800 238.800 200.400 ;
        RECT 242.200 195.800 243.000 200.400 ;
        RECT 244.400 195.800 245.200 200.400 ;
        RECT 247.600 195.800 248.400 200.400 ;
        RECT 249.200 191.800 250.000 200.400 ;
        RECT 252.400 193.000 253.200 200.400 ;
        RECT 255.600 195.800 256.400 200.400 ;
        RECT 258.800 195.800 259.600 200.400 ;
        RECT 262.000 195.800 262.800 200.400 ;
        RECT 268.400 195.800 269.200 200.400 ;
        RECT 271.600 195.800 272.400 200.400 ;
        RECT 279.600 195.800 280.400 200.400 ;
        RECT 282.800 195.800 283.600 200.400 ;
        RECT 286.000 195.800 286.800 200.400 ;
        RECT 289.200 195.800 290.000 200.400 ;
        RECT 291.400 195.800 292.200 200.400 ;
        RECT 258.800 191.800 259.600 192.400 ;
        RECT 262.200 191.800 263.000 192.000 ;
        RECT 295.600 191.800 296.400 200.400 ;
        RECT 298.800 193.000 299.600 200.400 ;
        RECT 302.000 191.800 302.800 200.400 ;
        RECT 308.400 195.800 309.200 200.400 ;
        RECT 311.600 191.800 312.400 200.400 ;
        RECT 316.400 191.800 317.200 200.400 ;
        RECT 320.600 195.800 321.400 200.400 ;
        RECT 322.800 195.800 323.600 200.400 ;
        RECT 326.000 195.800 326.800 200.400 ;
        RECT 329.200 195.800 330.000 200.400 ;
        RECT 332.400 195.800 333.200 200.400 ;
        RECT 340.400 195.800 341.200 200.400 ;
        RECT 343.600 195.800 344.400 200.400 ;
        RECT 350.000 195.800 350.800 200.400 ;
        RECT 353.200 195.800 354.000 200.400 ;
        RECT 356.400 195.800 357.200 200.400 ;
        RECT 358.600 195.800 359.400 200.400 ;
        RECT 349.800 191.800 350.800 192.000 ;
        RECT 353.200 191.800 354.000 192.400 ;
        RECT 362.800 191.800 363.600 200.400 ;
        RECT 364.400 195.800 365.200 200.400 ;
        RECT 367.600 195.800 368.400 200.400 ;
        RECT 370.800 195.800 371.600 200.400 ;
        RECT 374.000 195.800 374.800 200.400 ;
        RECT 382.000 195.800 382.800 200.400 ;
        RECT 385.200 195.800 386.000 200.400 ;
        RECT 391.600 195.800 392.400 200.400 ;
        RECT 394.800 195.800 395.600 200.400 ;
        RECT 398.000 195.800 398.800 200.400 ;
        RECT 399.600 195.800 400.400 200.400 ;
        RECT 402.800 195.800 403.600 200.400 ;
        RECT 406.000 195.800 406.800 200.400 ;
        RECT 412.400 195.800 413.200 200.400 ;
        RECT 415.600 195.800 416.400 200.400 ;
        RECT 423.600 195.800 424.400 200.400 ;
        RECT 426.800 195.800 427.600 200.400 ;
        RECT 430.000 195.800 430.800 200.400 ;
        RECT 433.200 195.800 434.000 200.400 ;
        RECT 434.800 195.800 435.600 200.400 ;
        RECT 438.000 195.800 438.800 200.400 ;
        RECT 441.200 195.800 442.000 200.400 ;
        RECT 447.600 195.800 448.400 200.400 ;
        RECT 450.800 195.800 451.600 200.400 ;
        RECT 458.800 195.800 459.600 200.400 ;
        RECT 462.000 195.800 462.800 200.400 ;
        RECT 465.200 195.800 466.000 200.400 ;
        RECT 468.400 195.800 469.200 200.400 ;
        RECT 391.400 191.800 392.200 192.000 ;
        RECT 394.800 191.800 395.600 192.400 ;
        RECT 4.400 191.200 31.400 191.800 ;
        RECT 30.600 191.000 31.400 191.200 ;
        RECT 176.600 191.200 203.600 191.800 ;
        RECT 258.800 191.200 285.800 191.800 ;
        RECT 176.600 191.000 177.400 191.200 ;
        RECT 285.000 191.000 285.800 191.200 ;
        RECT 327.000 191.200 354.000 191.800 ;
        RECT 368.600 191.200 395.600 191.800 ;
        RECT 402.800 191.800 403.600 192.400 ;
        RECT 406.000 191.800 407.000 192.000 ;
        RECT 438.000 191.800 438.800 192.400 ;
        RECT 476.400 192.000 477.200 200.400 ;
        RECT 482.000 195.800 482.800 200.400 ;
        RECT 485.200 195.800 486.000 200.400 ;
        RECT 441.400 191.800 442.200 192.000 ;
        RECT 490.800 191.800 491.600 200.400 ;
        RECT 494.000 191.800 494.800 200.400 ;
        RECT 498.200 195.800 499.000 200.400 ;
        RECT 500.400 195.800 501.200 200.400 ;
        RECT 503.600 195.800 504.400 200.400 ;
        RECT 505.200 191.800 506.000 200.400 ;
        RECT 508.400 191.800 509.200 200.400 ;
        RECT 511.600 191.800 512.400 200.400 ;
        RECT 516.400 191.800 517.200 200.400 ;
        RECT 518.600 195.800 519.400 200.400 ;
        RECT 522.800 191.800 523.600 200.400 ;
        RECT 526.000 195.800 526.800 200.400 ;
        RECT 527.600 195.800 528.400 200.400 ;
        RECT 530.800 195.800 531.600 200.400 ;
        RECT 534.000 195.800 534.800 200.400 ;
        RECT 537.200 195.800 538.000 200.400 ;
        RECT 545.200 195.800 546.000 200.400 ;
        RECT 548.400 195.800 549.200 200.400 ;
        RECT 554.800 195.800 555.600 200.400 ;
        RECT 558.000 195.800 558.800 200.400 ;
        RECT 561.200 195.800 562.000 200.400 ;
        RECT 562.800 195.800 563.600 200.400 ;
        RECT 566.000 195.800 566.800 200.400 ;
        RECT 569.200 195.800 570.000 200.400 ;
        RECT 575.600 195.800 576.400 200.400 ;
        RECT 578.800 195.800 579.600 200.400 ;
        RECT 586.800 195.800 587.600 200.400 ;
        RECT 590.000 195.800 590.800 200.400 ;
        RECT 593.200 195.800 594.000 200.400 ;
        RECT 596.400 195.800 597.200 200.400 ;
        RECT 598.600 195.800 599.400 200.400 ;
        RECT 554.600 191.800 555.400 192.000 ;
        RECT 558.000 191.800 558.800 192.400 ;
        RECT 402.800 191.200 429.800 191.800 ;
        RECT 438.000 191.200 465.000 191.800 ;
        RECT 327.000 191.000 327.800 191.200 ;
        RECT 368.600 191.000 369.400 191.200 ;
        RECT 429.000 191.000 429.800 191.200 ;
        RECT 464.200 191.000 465.000 191.200 ;
        RECT 531.800 191.200 558.800 191.800 ;
        RECT 566.000 191.800 566.800 192.400 ;
        RECT 569.200 191.800 570.200 192.000 ;
        RECT 602.800 191.800 603.600 200.400 ;
        RECT 606.000 193.000 606.800 200.400 ;
        RECT 566.000 191.200 593.000 191.800 ;
        RECT 531.800 191.000 532.600 191.200 ;
        RECT 592.200 191.000 593.000 191.200 ;
        RECT 154.200 170.800 155.000 171.000 ;
        RECT 211.800 170.800 212.600 171.000 ;
        RECT 272.200 170.800 273.000 171.000 ;
        RECT 331.400 170.800 332.200 171.000 ;
        RECT 154.200 170.200 181.200 170.800 ;
        RECT 211.800 170.200 238.800 170.800 ;
        RECT 2.800 161.600 3.600 170.000 ;
        RECT 8.400 161.600 9.200 166.200 ;
        RECT 11.600 161.600 12.400 166.200 ;
        RECT 17.200 161.600 18.000 170.200 ;
        RECT 21.000 161.600 21.800 166.200 ;
        RECT 25.200 161.600 26.000 170.200 ;
        RECT 28.400 161.600 29.200 169.800 ;
        RECT 33.600 161.600 34.400 170.200 ;
        RECT 36.400 161.600 37.200 170.200 ;
        RECT 39.600 161.600 40.400 169.000 ;
        RECT 43.400 161.600 44.200 166.200 ;
        RECT 47.600 161.600 48.400 170.200 ;
        RECT 50.800 161.600 51.600 166.200 ;
        RECT 54.000 161.600 54.800 170.200 ;
        RECT 59.600 161.600 60.400 166.200 ;
        RECT 62.800 161.600 63.600 166.200 ;
        RECT 68.400 161.600 69.200 170.000 ;
        RECT 72.800 161.600 73.600 170.200 ;
        RECT 78.000 161.600 78.800 169.800 ;
        RECT 81.200 161.600 82.000 170.200 ;
        RECT 85.400 161.600 86.200 166.200 ;
        RECT 88.200 161.600 89.000 166.200 ;
        RECT 92.400 161.600 93.200 170.200 ;
        RECT 94.000 161.600 94.800 166.200 ;
        RECT 98.400 161.600 99.200 170.200 ;
        RECT 103.600 161.600 104.400 169.800 ;
        RECT 106.800 161.600 107.600 166.200 ;
        RECT 110.000 161.600 110.800 166.200 ;
        RECT 113.200 161.600 114.000 166.200 ;
        RECT 114.800 161.600 115.600 166.200 ;
        RECT 118.000 161.600 118.800 166.200 ;
        RECT 121.200 161.600 122.000 166.200 ;
        RECT 124.400 161.600 125.200 166.200 ;
        RECT 126.000 161.600 126.800 170.200 ;
        RECT 130.800 161.600 131.600 170.200 ;
        RECT 134.000 161.600 134.800 169.000 ;
        RECT 137.200 161.600 138.000 166.200 ;
        RECT 143.600 161.600 144.400 170.200 ;
        RECT 177.000 170.000 177.800 170.200 ;
        RECT 180.400 169.600 181.200 170.200 ;
        RECT 150.000 161.600 150.800 166.200 ;
        RECT 153.200 161.600 154.000 166.200 ;
        RECT 156.400 161.600 157.200 166.200 ;
        RECT 159.600 161.600 160.400 166.200 ;
        RECT 167.600 161.600 168.400 166.200 ;
        RECT 170.800 161.600 171.600 166.200 ;
        RECT 177.200 161.600 178.000 166.200 ;
        RECT 180.400 161.600 181.200 166.200 ;
        RECT 183.600 161.600 184.400 166.200 ;
        RECT 185.200 161.600 186.000 170.200 ;
        RECT 188.400 161.600 189.200 169.000 ;
        RECT 191.600 161.600 192.400 166.200 ;
        RECT 194.800 161.600 195.600 166.200 ;
        RECT 196.400 161.600 197.200 166.200 ;
        RECT 199.600 161.600 200.400 166.200 ;
        RECT 201.800 161.600 202.600 166.200 ;
        RECT 206.000 161.600 206.800 170.200 ;
        RECT 234.600 170.000 235.600 170.200 ;
        RECT 238.000 169.600 238.800 170.200 ;
        RECT 246.000 170.200 273.000 170.800 ;
        RECT 305.200 170.200 332.200 170.800 ;
        RECT 568.600 170.800 569.400 171.000 ;
        RECT 568.600 170.200 595.600 170.800 ;
        RECT 246.000 169.600 246.800 170.200 ;
        RECT 249.400 170.000 250.200 170.200 ;
        RECT 207.600 161.600 208.400 166.200 ;
        RECT 210.800 161.600 211.600 166.200 ;
        RECT 214.000 161.600 214.800 166.200 ;
        RECT 217.200 161.600 218.000 166.200 ;
        RECT 225.200 161.600 226.000 166.200 ;
        RECT 228.400 161.600 229.200 166.200 ;
        RECT 234.800 161.600 235.600 166.200 ;
        RECT 238.000 161.600 238.800 166.200 ;
        RECT 241.200 161.600 242.000 166.200 ;
        RECT 242.800 161.600 243.600 166.200 ;
        RECT 246.000 161.600 246.800 166.200 ;
        RECT 249.200 161.600 250.000 166.200 ;
        RECT 255.600 161.600 256.400 166.200 ;
        RECT 258.800 161.600 259.600 166.200 ;
        RECT 266.800 161.600 267.600 166.200 ;
        RECT 270.000 161.600 270.800 166.200 ;
        RECT 273.200 161.600 274.000 166.200 ;
        RECT 276.400 161.600 277.200 166.200 ;
        RECT 278.000 161.600 278.800 166.200 ;
        RECT 281.200 161.600 282.000 166.200 ;
        RECT 282.800 161.600 283.600 170.200 ;
        RECT 286.000 161.600 286.800 170.200 ;
        RECT 289.200 161.600 290.000 170.200 ;
        RECT 292.400 161.600 293.200 170.200 ;
        RECT 295.600 161.600 296.400 170.200 ;
        RECT 305.200 169.600 306.000 170.200 ;
        RECT 308.400 170.000 309.400 170.200 ;
        RECT 302.000 161.600 302.800 166.200 ;
        RECT 305.200 161.600 306.000 166.200 ;
        RECT 308.400 161.600 309.200 166.200 ;
        RECT 314.800 161.600 315.600 166.200 ;
        RECT 318.000 161.600 318.800 166.200 ;
        RECT 326.000 161.600 326.800 166.200 ;
        RECT 329.200 161.600 330.000 166.200 ;
        RECT 332.400 161.600 333.200 166.200 ;
        RECT 335.600 161.600 336.400 166.200 ;
        RECT 337.200 161.600 338.000 166.200 ;
        RECT 340.400 161.600 341.200 166.200 ;
        RECT 342.600 161.600 343.400 166.200 ;
        RECT 346.800 161.600 347.600 170.200 ;
        RECT 348.400 161.600 349.200 166.200 ;
        RECT 351.600 161.600 352.400 166.200 ;
        RECT 354.800 161.600 355.600 169.000 ;
        RECT 358.000 161.600 358.800 170.200 ;
        RECT 359.600 161.600 360.400 166.200 ;
        RECT 362.800 161.600 363.600 166.200 ;
        RECT 364.400 161.600 365.200 170.200 ;
        RECT 368.600 161.600 369.400 166.200 ;
        RECT 372.400 161.600 373.200 169.000 ;
        RECT 375.600 161.600 376.400 170.200 ;
        RECT 377.200 161.600 378.000 166.200 ;
        RECT 380.400 161.600 381.200 166.200 ;
        RECT 383.600 161.600 384.400 166.200 ;
        RECT 386.800 161.600 387.600 170.200 ;
        RECT 392.400 161.600 393.200 166.200 ;
        RECT 395.600 161.600 396.400 166.200 ;
        RECT 401.200 161.600 402.000 170.000 ;
        RECT 404.400 161.600 405.200 170.200 ;
        RECT 408.600 161.600 409.400 166.200 ;
        RECT 411.400 161.600 412.200 166.200 ;
        RECT 415.600 161.600 416.400 170.200 ;
        RECT 418.400 161.600 419.200 170.200 ;
        RECT 423.600 161.600 424.400 169.800 ;
        RECT 428.400 161.600 429.200 170.000 ;
        RECT 434.000 161.600 434.800 166.200 ;
        RECT 437.200 161.600 438.000 166.200 ;
        RECT 442.800 161.600 443.600 170.200 ;
        RECT 446.000 161.600 446.800 170.200 ;
        RECT 450.200 161.600 451.000 166.200 ;
        RECT 453.000 161.600 453.800 166.200 ;
        RECT 457.200 161.600 458.000 170.200 ;
        RECT 463.600 161.600 464.400 170.200 ;
        RECT 467.800 161.600 468.600 166.200 ;
        RECT 470.000 161.600 470.800 170.200 ;
        RECT 474.200 161.600 475.000 166.200 ;
        RECT 477.600 161.600 478.400 170.200 ;
        RECT 482.800 161.600 483.600 169.800 ;
        RECT 487.600 161.600 488.400 170.200 ;
        RECT 493.200 161.600 494.000 166.200 ;
        RECT 496.400 161.600 497.200 166.200 ;
        RECT 502.000 161.600 502.800 170.000 ;
        RECT 505.200 161.600 506.000 170.200 ;
        RECT 509.400 161.600 510.200 166.200 ;
        RECT 512.200 161.600 513.000 166.200 ;
        RECT 516.400 161.600 517.200 170.200 ;
        RECT 519.600 161.600 520.400 169.800 ;
        RECT 524.800 161.600 525.600 170.200 ;
        RECT 529.200 161.600 530.000 169.800 ;
        RECT 534.400 161.600 535.200 170.200 ;
        RECT 537.200 161.600 538.000 170.200 ;
        RECT 541.400 161.600 542.200 166.200 ;
        RECT 543.600 161.600 544.400 170.200 ;
        RECT 547.800 161.600 548.600 166.200 ;
        RECT 551.600 161.600 552.400 166.200 ;
        RECT 553.200 161.600 554.000 166.200 ;
        RECT 556.400 161.600 557.200 166.200 ;
        RECT 558.000 161.600 558.800 170.200 ;
        RECT 591.400 170.000 592.400 170.200 ;
        RECT 594.800 169.600 595.600 170.200 ;
        RECT 562.200 161.600 563.000 166.200 ;
        RECT 564.400 161.600 565.200 166.200 ;
        RECT 567.600 161.600 568.400 166.200 ;
        RECT 570.800 161.600 571.600 166.200 ;
        RECT 574.000 161.600 574.800 166.200 ;
        RECT 582.000 161.600 582.800 166.200 ;
        RECT 585.200 161.600 586.000 166.200 ;
        RECT 591.600 161.600 592.400 166.200 ;
        RECT 594.800 161.600 595.600 166.200 ;
        RECT 598.000 161.600 598.800 166.200 ;
        RECT 600.200 161.600 601.000 166.200 ;
        RECT 604.400 161.600 605.200 170.200 ;
        RECT 607.600 161.600 608.400 166.200 ;
        RECT 0.400 160.400 614.000 161.600 ;
        RECT 2.800 152.000 3.600 160.400 ;
        RECT 8.400 155.800 9.200 160.400 ;
        RECT 11.600 155.800 12.400 160.400 ;
        RECT 17.200 151.800 18.000 160.400 ;
        RECT 21.000 155.800 21.800 160.400 ;
        RECT 25.200 151.800 26.000 160.400 ;
        RECT 26.800 151.800 27.600 160.400 ;
        RECT 31.000 155.800 31.800 160.400 ;
        RECT 33.800 155.800 34.600 160.400 ;
        RECT 38.000 151.800 38.800 160.400 ;
        RECT 40.800 151.800 41.600 160.400 ;
        RECT 46.000 152.200 46.800 160.400 ;
        RECT 50.400 151.800 51.200 160.400 ;
        RECT 55.600 152.200 56.400 160.400 ;
        RECT 58.800 151.800 59.600 160.400 ;
        RECT 63.000 155.800 63.800 160.400 ;
        RECT 65.800 155.800 66.600 160.400 ;
        RECT 70.000 151.800 70.800 160.400 ;
        RECT 73.200 152.000 74.000 160.400 ;
        RECT 78.800 155.800 79.600 160.400 ;
        RECT 82.000 155.800 82.800 160.400 ;
        RECT 87.600 151.800 88.400 160.400 ;
        RECT 90.800 155.800 91.600 160.400 ;
        RECT 94.000 156.200 94.800 160.400 ;
        RECT 97.200 151.800 98.000 160.400 ;
        RECT 101.400 155.800 102.200 160.400 ;
        RECT 103.600 155.800 104.400 160.400 ;
        RECT 106.800 156.200 107.600 160.400 ;
        RECT 110.000 151.800 110.800 160.400 ;
        RECT 114.200 155.800 115.000 160.400 ;
        RECT 117.000 155.800 117.800 160.400 ;
        RECT 121.200 151.800 122.000 160.400 ;
        RECT 122.800 151.800 123.600 160.400 ;
        RECT 127.000 155.800 127.800 160.400 ;
        RECT 129.200 151.800 130.000 160.400 ;
        RECT 133.400 155.800 134.200 160.400 ;
        RECT 135.600 151.800 136.400 160.400 ;
        RECT 139.800 155.800 140.600 160.400 ;
        RECT 142.000 151.800 142.800 160.400 ;
        RECT 146.800 153.200 147.800 160.400 ;
        RECT 153.000 159.800 153.800 160.400 ;
        RECT 153.000 153.200 154.000 159.800 ;
        RECT 161.200 155.800 162.000 160.400 ;
        RECT 164.400 155.800 165.200 160.400 ;
        RECT 167.600 155.800 168.400 160.400 ;
        RECT 174.000 155.800 174.800 160.400 ;
        RECT 177.200 155.800 178.000 160.400 ;
        RECT 185.200 155.800 186.000 160.400 ;
        RECT 188.400 155.800 189.200 160.400 ;
        RECT 191.600 155.800 192.400 160.400 ;
        RECT 194.800 155.800 195.600 160.400 ;
        RECT 197.000 155.800 197.800 160.400 ;
        RECT 164.400 151.800 165.200 152.400 ;
        RECT 167.600 151.800 168.600 152.000 ;
        RECT 201.200 151.800 202.000 160.400 ;
        RECT 202.800 151.800 203.600 160.400 ;
        RECT 206.000 153.000 206.800 160.400 ;
        RECT 212.400 151.800 213.200 160.400 ;
        RECT 214.000 155.800 214.800 160.400 ;
        RECT 217.200 155.800 218.000 160.400 ;
        RECT 218.800 151.800 219.600 160.400 ;
        RECT 223.000 155.800 223.800 160.400 ;
        RECT 225.200 155.800 226.000 160.400 ;
        RECT 228.400 155.800 229.200 160.400 ;
        RECT 231.600 155.800 232.400 160.400 ;
        RECT 238.000 155.800 238.800 160.400 ;
        RECT 241.200 155.800 242.000 160.400 ;
        RECT 249.200 155.800 250.000 160.400 ;
        RECT 252.400 155.800 253.200 160.400 ;
        RECT 255.600 155.800 256.400 160.400 ;
        RECT 258.800 155.800 259.600 160.400 ;
        RECT 260.400 155.800 261.200 160.400 ;
        RECT 263.600 155.800 264.400 160.400 ;
        RECT 265.200 155.800 266.000 160.400 ;
        RECT 268.400 155.800 269.200 160.400 ;
        RECT 271.600 155.800 272.400 160.400 ;
        RECT 278.000 155.800 278.800 160.400 ;
        RECT 281.200 155.800 282.000 160.400 ;
        RECT 289.200 155.800 290.000 160.400 ;
        RECT 292.400 155.800 293.200 160.400 ;
        RECT 295.600 155.800 296.400 160.400 ;
        RECT 298.800 155.800 299.600 160.400 ;
        RECT 302.000 155.800 302.800 160.400 ;
        RECT 228.400 151.800 229.200 152.400 ;
        RECT 231.600 151.800 232.600 152.000 ;
        RECT 268.400 151.800 269.200 152.400 ;
        RECT 271.800 151.800 272.600 152.000 ;
        RECT 308.400 151.800 309.200 160.400 ;
        RECT 312.600 155.800 313.400 160.400 ;
        RECT 314.800 155.800 315.600 160.400 ;
        RECT 318.000 155.800 318.800 160.400 ;
        RECT 319.600 155.800 320.400 160.400 ;
        RECT 322.800 155.800 323.600 160.400 ;
        RECT 326.000 155.800 326.800 160.400 ;
        RECT 332.400 155.800 333.200 160.400 ;
        RECT 335.600 155.800 336.400 160.400 ;
        RECT 343.600 155.800 344.400 160.400 ;
        RECT 346.800 155.800 347.600 160.400 ;
        RECT 350.000 155.800 350.800 160.400 ;
        RECT 353.200 155.800 354.000 160.400 ;
        RECT 354.800 155.800 355.600 160.400 ;
        RECT 358.000 155.800 358.800 160.400 ;
        RECT 360.200 155.800 361.000 160.400 ;
        RECT 322.800 151.800 323.600 152.400 ;
        RECT 326.000 151.800 327.000 152.000 ;
        RECT 364.400 151.800 365.200 160.400 ;
        RECT 366.000 155.800 366.800 160.400 ;
        RECT 369.200 155.800 370.000 160.400 ;
        RECT 371.400 155.800 372.200 160.400 ;
        RECT 375.600 151.800 376.400 160.400 ;
        RECT 377.800 155.800 378.600 160.400 ;
        RECT 382.000 151.800 382.800 160.400 ;
        RECT 383.600 151.800 384.400 160.400 ;
        RECT 387.800 155.800 388.600 160.400 ;
        RECT 390.600 155.800 391.400 160.400 ;
        RECT 394.800 151.800 395.600 160.400 ;
        RECT 398.000 156.200 398.800 160.400 ;
        RECT 401.200 155.800 402.000 160.400 ;
        RECT 404.400 156.200 405.200 160.400 ;
        RECT 407.600 155.800 408.400 160.400 ;
        RECT 409.200 151.800 410.000 160.400 ;
        RECT 413.400 155.800 414.200 160.400 ;
        RECT 416.200 155.800 417.000 160.400 ;
        RECT 420.400 151.800 421.200 160.400 ;
        RECT 423.200 151.800 424.000 160.400 ;
        RECT 428.400 152.200 429.200 160.400 ;
        RECT 432.200 155.800 433.000 160.400 ;
        RECT 436.400 151.800 437.200 160.400 ;
        RECT 439.600 155.800 440.400 160.400 ;
        RECT 442.800 152.200 443.600 160.400 ;
        RECT 448.000 151.800 448.800 160.400 ;
        RECT 450.800 155.800 451.600 160.400 ;
        RECT 454.000 155.800 454.800 160.400 ;
        RECT 462.000 151.800 462.800 160.400 ;
        RECT 467.600 155.800 468.400 160.400 ;
        RECT 470.800 155.800 471.600 160.400 ;
        RECT 476.400 152.000 477.200 160.400 ;
        RECT 481.200 155.800 482.000 160.400 ;
        RECT 484.400 152.200 485.200 160.400 ;
        RECT 489.600 151.800 490.400 160.400 ;
        RECT 492.400 155.800 493.200 160.400 ;
        RECT 495.600 155.800 496.400 160.400 ;
        RECT 497.800 155.800 498.600 160.400 ;
        RECT 502.000 151.800 502.800 160.400 ;
        RECT 503.600 151.800 504.400 160.400 ;
        RECT 507.800 155.800 508.600 160.400 ;
        RECT 510.600 155.800 511.400 160.400 ;
        RECT 514.800 151.800 515.600 160.400 ;
        RECT 518.000 151.800 518.800 160.400 ;
        RECT 523.600 155.800 524.400 160.400 ;
        RECT 526.800 155.800 527.600 160.400 ;
        RECT 532.400 152.000 533.200 160.400 ;
        RECT 535.600 151.800 536.400 160.400 ;
        RECT 539.800 155.800 540.600 160.400 ;
        RECT 543.600 151.800 544.400 160.400 ;
        RECT 549.200 155.800 550.000 160.400 ;
        RECT 552.400 155.800 553.200 160.400 ;
        RECT 558.000 152.000 558.800 160.400 ;
        RECT 563.800 151.800 564.600 160.400 ;
        RECT 567.600 155.800 568.400 160.400 ;
        RECT 570.800 155.800 571.600 160.400 ;
        RECT 574.000 155.800 574.800 160.400 ;
        RECT 577.200 155.800 578.000 160.400 ;
        RECT 585.200 155.800 586.000 160.400 ;
        RECT 588.400 155.800 589.200 160.400 ;
        RECT 594.800 155.800 595.600 160.400 ;
        RECT 598.000 155.800 598.800 160.400 ;
        RECT 601.200 155.800 602.000 160.400 ;
        RECT 604.400 155.800 605.200 160.400 ;
        RECT 607.600 153.000 608.400 160.400 ;
        RECT 594.600 151.800 595.400 152.000 ;
        RECT 598.000 151.800 598.800 152.400 ;
        RECT 164.400 151.200 191.400 151.800 ;
        RECT 228.400 151.200 255.400 151.800 ;
        RECT 268.400 151.200 295.400 151.800 ;
        RECT 322.800 151.200 349.800 151.800 ;
        RECT 190.600 151.000 191.400 151.200 ;
        RECT 254.600 151.000 255.400 151.200 ;
        RECT 294.600 151.000 295.400 151.200 ;
        RECT 349.000 151.000 349.800 151.200 ;
        RECT 571.800 151.200 598.800 151.800 ;
        RECT 571.800 151.000 572.600 151.200 ;
        RECT 5.400 130.800 6.200 131.000 ;
        RECT 167.000 130.800 167.800 131.000 ;
        RECT 213.400 130.800 214.200 131.000 ;
        RECT 271.000 130.800 271.800 131.000 ;
        RECT 350.600 130.800 351.400 131.000 ;
        RECT 408.200 130.800 409.000 131.000 ;
        RECT 5.400 130.200 32.400 130.800 ;
        RECT 167.000 130.200 194.000 130.800 ;
        RECT 213.400 130.200 240.400 130.800 ;
        RECT 271.000 130.200 298.000 130.800 ;
        RECT 324.400 130.200 351.400 130.800 ;
        RECT 382.000 130.200 409.000 130.800 ;
        RECT 28.200 130.000 29.000 130.200 ;
        RECT 31.600 129.600 32.400 130.200 ;
        RECT 1.200 121.600 2.000 126.200 ;
        RECT 4.400 121.600 5.200 126.200 ;
        RECT 7.600 121.600 8.400 126.200 ;
        RECT 10.800 121.600 11.600 126.200 ;
        RECT 18.800 121.600 19.600 126.200 ;
        RECT 22.000 121.600 22.800 126.200 ;
        RECT 28.400 121.600 29.200 126.200 ;
        RECT 31.600 121.600 32.400 126.200 ;
        RECT 34.800 121.600 35.600 126.200 ;
        RECT 36.400 121.600 37.200 126.200 ;
        RECT 39.600 121.600 40.400 126.200 ;
        RECT 41.800 121.600 42.600 126.200 ;
        RECT 46.000 121.600 46.800 130.200 ;
        RECT 48.800 121.600 49.600 130.200 ;
        RECT 54.000 121.600 54.800 129.800 ;
        RECT 57.200 121.600 58.000 130.200 ;
        RECT 61.400 121.600 62.200 126.200 ;
        RECT 64.200 121.600 65.000 126.200 ;
        RECT 68.400 121.600 69.200 130.200 ;
        RECT 71.600 121.600 72.400 130.000 ;
        RECT 77.200 121.600 78.000 126.200 ;
        RECT 80.400 121.600 81.200 126.200 ;
        RECT 86.000 121.600 86.800 130.200 ;
        RECT 89.200 121.600 90.000 130.200 ;
        RECT 92.400 121.600 93.200 129.000 ;
        RECT 96.200 121.600 97.000 126.200 ;
        RECT 100.400 121.600 101.200 130.200 ;
        RECT 103.600 121.600 104.400 130.000 ;
        RECT 109.200 121.600 110.000 126.200 ;
        RECT 112.400 121.600 113.200 126.200 ;
        RECT 118.000 121.600 118.800 130.200 ;
        RECT 121.200 121.600 122.000 126.200 ;
        RECT 124.400 121.600 125.200 126.200 ;
        RECT 126.000 121.600 126.800 126.200 ;
        RECT 129.200 121.600 130.000 126.200 ;
        RECT 132.400 121.600 133.200 126.200 ;
        RECT 134.000 121.600 134.800 130.200 ;
        RECT 138.200 121.600 139.000 126.200 ;
        RECT 140.400 121.600 141.200 130.200 ;
        RECT 144.600 121.600 145.400 126.200 ;
        RECT 146.800 121.600 147.600 126.200 ;
        RECT 150.000 121.600 150.800 126.200 ;
        RECT 156.400 121.600 157.200 130.200 ;
        RECT 189.800 130.000 190.800 130.200 ;
        RECT 193.200 129.600 194.000 130.200 ;
        RECT 160.600 121.600 161.400 126.200 ;
        RECT 162.800 121.600 163.600 126.200 ;
        RECT 166.000 121.600 166.800 126.200 ;
        RECT 169.200 121.600 170.000 126.200 ;
        RECT 172.400 121.600 173.200 126.200 ;
        RECT 180.400 121.600 181.200 126.200 ;
        RECT 183.600 121.600 184.400 126.200 ;
        RECT 190.000 121.600 190.800 126.200 ;
        RECT 193.200 121.600 194.000 126.200 ;
        RECT 196.400 121.600 197.200 126.200 ;
        RECT 198.000 121.600 198.800 126.200 ;
        RECT 201.200 121.600 202.000 126.200 ;
        RECT 202.800 121.600 203.600 130.200 ;
        RECT 236.200 130.000 237.000 130.200 ;
        RECT 239.600 129.600 240.400 130.200 ;
        RECT 206.000 121.600 206.800 129.000 ;
        RECT 209.200 121.600 210.000 126.200 ;
        RECT 212.400 121.600 213.200 126.200 ;
        RECT 215.600 121.600 216.400 126.200 ;
        RECT 218.800 121.600 219.600 126.200 ;
        RECT 226.800 121.600 227.600 126.200 ;
        RECT 230.000 121.600 230.800 126.200 ;
        RECT 236.400 121.600 237.200 126.200 ;
        RECT 239.600 121.600 240.400 126.200 ;
        RECT 242.800 121.600 243.600 126.200 ;
        RECT 247.600 121.600 248.400 130.200 ;
        RECT 249.200 121.600 250.000 130.200 ;
        RECT 255.600 121.600 256.400 129.000 ;
        RECT 258.800 121.600 259.600 130.200 ;
        RECT 260.400 121.600 261.200 130.200 ;
        RECT 293.800 130.000 294.800 130.200 ;
        RECT 297.200 129.600 298.000 130.200 ;
        RECT 264.600 121.600 265.400 126.200 ;
        RECT 266.800 121.600 267.600 126.200 ;
        RECT 270.000 121.600 270.800 126.200 ;
        RECT 273.200 121.600 274.000 126.200 ;
        RECT 276.400 121.600 277.200 126.200 ;
        RECT 284.400 121.600 285.200 126.200 ;
        RECT 287.600 121.600 288.400 126.200 ;
        RECT 294.000 121.600 294.800 126.200 ;
        RECT 297.200 121.600 298.000 126.200 ;
        RECT 300.400 121.600 301.200 126.200 ;
        RECT 306.800 121.600 307.600 130.200 ;
        RECT 310.000 121.600 310.800 130.200 ;
        RECT 313.200 121.600 314.000 130.200 ;
        RECT 316.400 121.600 317.200 130.200 ;
        RECT 319.600 121.600 320.400 130.200 ;
        RECT 324.400 129.600 325.200 130.200 ;
        RECT 327.800 130.000 328.600 130.200 ;
        RECT 321.200 121.600 322.000 126.200 ;
        RECT 324.400 121.600 325.200 126.200 ;
        RECT 327.600 121.600 328.400 126.200 ;
        RECT 334.000 121.600 334.800 126.200 ;
        RECT 337.200 121.600 338.000 126.200 ;
        RECT 345.200 121.600 346.000 126.200 ;
        RECT 348.400 121.600 349.200 126.200 ;
        RECT 351.600 121.600 352.400 126.200 ;
        RECT 354.800 121.600 355.600 126.200 ;
        RECT 358.000 121.600 358.800 129.000 ;
        RECT 361.200 121.600 362.000 130.200 ;
        RECT 364.400 121.600 365.200 129.000 ;
        RECT 367.600 121.600 368.400 130.200 ;
        RECT 382.000 129.600 382.800 130.200 ;
        RECT 385.200 130.000 386.200 130.200 ;
        RECT 371.800 121.600 372.600 126.200 ;
        RECT 374.000 121.600 374.800 126.200 ;
        RECT 377.200 121.600 378.000 126.200 ;
        RECT 378.800 121.600 379.600 126.200 ;
        RECT 382.000 121.600 382.800 126.200 ;
        RECT 385.200 121.600 386.000 126.200 ;
        RECT 391.600 121.600 392.400 126.200 ;
        RECT 394.800 121.600 395.600 126.200 ;
        RECT 402.800 121.600 403.600 126.200 ;
        RECT 406.000 121.600 406.800 126.200 ;
        RECT 409.200 121.600 410.000 126.200 ;
        RECT 412.400 121.600 413.200 126.200 ;
        RECT 414.000 121.600 414.800 130.200 ;
        RECT 417.200 121.600 418.000 130.200 ;
        RECT 420.400 121.600 421.200 130.200 ;
        RECT 423.600 121.600 424.400 130.200 ;
        RECT 426.800 121.600 427.600 130.200 ;
        RECT 429.000 121.600 429.800 126.200 ;
        RECT 433.200 121.600 434.000 130.200 ;
        RECT 436.400 121.600 437.200 129.000 ;
        RECT 439.600 121.600 440.400 130.200 ;
        RECT 442.800 121.600 443.600 125.800 ;
        RECT 446.000 121.600 446.800 126.200 ;
        RECT 447.600 121.600 448.400 130.200 ;
        RECT 454.000 122.200 455.000 128.800 ;
        RECT 454.200 121.600 455.000 122.200 ;
        RECT 460.200 121.600 461.200 128.800 ;
        RECT 470.000 121.600 470.800 126.200 ;
        RECT 471.600 121.600 472.400 130.200 ;
        RECT 476.400 121.600 477.200 130.200 ;
        RECT 480.600 121.600 481.400 126.200 ;
        RECT 482.800 121.600 483.600 130.200 ;
        RECT 486.000 121.600 486.800 129.000 ;
        RECT 489.800 121.600 490.600 126.200 ;
        RECT 494.000 121.600 494.800 130.200 ;
        RECT 496.800 121.600 497.600 130.200 ;
        RECT 502.000 121.600 502.800 129.800 ;
        RECT 505.200 121.600 506.000 130.200 ;
        RECT 508.400 121.600 509.200 129.000 ;
        RECT 511.600 121.600 512.400 130.200 ;
        RECT 515.800 121.600 516.600 126.200 ;
        RECT 519.600 121.600 520.400 130.200 ;
        RECT 525.200 121.600 526.000 126.200 ;
        RECT 528.400 121.600 529.200 126.200 ;
        RECT 534.000 121.600 534.800 130.000 ;
        RECT 537.200 121.600 538.000 130.200 ;
        RECT 541.400 121.600 542.200 126.200 ;
        RECT 545.200 121.600 546.000 126.200 ;
        RECT 548.400 121.600 549.200 129.000 ;
        RECT 551.600 121.600 552.400 130.200 ;
        RECT 554.800 121.600 555.600 129.000 ;
        RECT 558.000 121.600 558.800 130.200 ;
        RECT 561.200 121.600 562.000 126.200 ;
        RECT 562.800 121.600 563.600 130.200 ;
        RECT 567.000 121.600 567.800 126.200 ;
        RECT 570.800 121.600 571.600 129.800 ;
        RECT 576.000 121.600 576.800 130.200 ;
        RECT 578.800 121.600 579.600 130.200 ;
        RECT 583.000 121.600 583.800 126.200 ;
        RECT 585.200 121.600 586.000 126.200 ;
        RECT 588.400 121.600 589.200 126.200 ;
        RECT 591.600 121.600 592.400 130.000 ;
        RECT 597.200 121.600 598.000 126.200 ;
        RECT 600.400 121.600 601.200 126.200 ;
        RECT 606.000 121.600 606.800 130.200 ;
        RECT 0.400 120.400 614.000 121.600 ;
        RECT 2.800 112.000 3.600 120.400 ;
        RECT 8.400 115.800 9.200 120.400 ;
        RECT 11.600 115.800 12.400 120.400 ;
        RECT 17.200 111.800 18.000 120.400 ;
        RECT 21.000 115.800 21.800 120.400 ;
        RECT 25.200 111.800 26.000 120.400 ;
        RECT 27.400 115.800 28.200 120.400 ;
        RECT 31.600 111.800 32.400 120.400 ;
        RECT 33.200 111.800 34.000 120.400 ;
        RECT 36.400 113.000 37.200 120.400 ;
        RECT 40.800 111.800 41.600 120.400 ;
        RECT 46.000 112.200 46.800 120.400 ;
        RECT 49.200 111.800 50.000 120.400 ;
        RECT 53.400 115.800 54.200 120.400 ;
        RECT 56.200 115.800 57.000 120.400 ;
        RECT 60.400 111.800 61.200 120.400 ;
        RECT 63.200 111.800 64.000 120.400 ;
        RECT 68.400 112.200 69.200 120.400 ;
        RECT 71.600 111.800 72.400 120.400 ;
        RECT 74.800 113.000 75.600 120.400 ;
        RECT 78.000 111.800 78.800 120.400 ;
        RECT 81.200 113.000 82.000 120.400 ;
        RECT 84.400 115.800 85.200 120.400 ;
        RECT 87.600 115.800 88.400 120.400 ;
        RECT 89.200 115.800 90.000 120.400 ;
        RECT 92.400 116.200 93.200 120.400 ;
        RECT 96.200 115.800 97.000 120.400 ;
        RECT 100.400 111.800 101.200 120.400 ;
        RECT 102.000 111.800 102.800 120.400 ;
        RECT 106.200 115.800 107.000 120.400 ;
        RECT 108.400 111.800 109.200 120.400 ;
        RECT 112.600 115.800 113.400 120.400 ;
        RECT 114.800 111.800 115.600 120.400 ;
        RECT 119.000 115.800 119.800 120.400 ;
        RECT 122.800 113.000 123.600 120.400 ;
        RECT 126.000 111.800 126.800 120.400 ;
        RECT 127.600 115.800 128.400 120.400 ;
        RECT 130.800 115.800 131.600 120.400 ;
        RECT 132.400 115.800 133.200 120.400 ;
        RECT 136.200 115.800 137.000 120.400 ;
        RECT 140.400 111.800 141.200 120.400 ;
        RECT 142.600 115.800 143.400 120.400 ;
        RECT 146.800 111.800 147.600 120.400 ;
        RECT 153.800 115.800 154.600 120.400 ;
        RECT 158.000 111.800 158.800 120.400 ;
        RECT 159.600 111.800 160.400 120.400 ;
        RECT 162.800 111.800 163.600 120.400 ;
        RECT 166.000 111.800 166.800 120.400 ;
        RECT 169.200 111.800 170.000 120.400 ;
        RECT 172.400 111.800 173.200 120.400 ;
        RECT 175.600 112.200 176.400 120.400 ;
        RECT 180.800 111.800 181.600 120.400 ;
        RECT 185.200 112.200 186.000 120.400 ;
        RECT 190.400 111.800 191.200 120.400 ;
        RECT 195.000 119.800 195.800 120.400 ;
        RECT 194.800 113.200 195.800 119.800 ;
        RECT 201.000 113.200 202.000 120.400 ;
        RECT 206.600 111.800 207.400 120.400 ;
        RECT 214.000 113.000 214.800 120.400 ;
        RECT 217.200 115.800 218.000 120.400 ;
        RECT 220.400 116.200 221.200 120.400 ;
        RECT 225.200 115.800 226.000 120.400 ;
        RECT 229.400 111.800 230.200 120.400 ;
        RECT 233.200 111.800 234.000 120.400 ;
        RECT 238.600 115.800 239.400 120.400 ;
        RECT 242.800 111.800 243.600 120.400 ;
        RECT 244.400 115.800 245.200 120.400 ;
        RECT 247.600 115.800 248.400 120.400 ;
        RECT 250.800 115.800 251.600 120.400 ;
        RECT 257.200 115.800 258.000 120.400 ;
        RECT 260.400 115.800 261.200 120.400 ;
        RECT 268.400 115.800 269.200 120.400 ;
        RECT 271.600 115.800 272.400 120.400 ;
        RECT 274.800 115.800 275.600 120.400 ;
        RECT 278.000 115.800 278.800 120.400 ;
        RECT 280.200 115.800 281.000 120.400 ;
        RECT 284.400 111.800 285.200 120.400 ;
        RECT 286.000 111.800 286.800 120.400 ;
        RECT 289.200 113.000 290.000 120.400 ;
        RECT 294.200 119.800 295.000 120.400 ;
        RECT 294.000 113.200 295.000 119.800 ;
        RECT 300.200 113.200 301.200 120.400 ;
        RECT 308.400 115.800 309.200 120.400 ;
        RECT 311.600 115.800 312.400 120.400 ;
        RECT 313.200 115.800 314.000 120.400 ;
        RECT 316.400 115.800 317.200 120.400 ;
        RECT 319.600 115.800 320.400 120.400 ;
        RECT 322.800 115.800 323.600 120.400 ;
        RECT 330.800 115.800 331.600 120.400 ;
        RECT 334.000 115.800 334.800 120.400 ;
        RECT 340.400 115.800 341.200 120.400 ;
        RECT 343.600 115.800 344.400 120.400 ;
        RECT 346.800 115.800 347.600 120.400 ;
        RECT 340.200 111.800 341.200 112.000 ;
        RECT 343.600 111.800 344.400 112.400 ;
        RECT 348.400 111.800 349.200 120.400 ;
        RECT 351.600 113.000 352.400 120.400 ;
        RECT 356.400 113.000 357.200 120.400 ;
        RECT 359.600 111.800 360.400 120.400 ;
        RECT 362.800 115.800 363.600 120.400 ;
        RECT 364.400 111.800 365.200 120.400 ;
        RECT 368.600 115.800 369.400 120.400 ;
        RECT 370.800 115.800 371.600 120.400 ;
        RECT 374.000 115.800 374.800 120.400 ;
        RECT 377.200 115.800 378.000 120.400 ;
        RECT 383.600 115.800 384.400 120.400 ;
        RECT 386.800 115.800 387.600 120.400 ;
        RECT 394.800 115.800 395.600 120.400 ;
        RECT 398.000 115.800 398.800 120.400 ;
        RECT 401.200 115.800 402.000 120.400 ;
        RECT 404.400 115.800 405.200 120.400 ;
        RECT 374.000 111.800 374.800 112.400 ;
        RECT 377.400 111.800 378.200 112.000 ;
        RECT 407.600 111.800 408.400 120.400 ;
        RECT 413.200 115.800 414.000 120.400 ;
        RECT 416.400 115.800 417.200 120.400 ;
        RECT 422.000 112.000 422.800 120.400 ;
        RECT 425.200 115.800 426.000 120.400 ;
        RECT 429.000 115.800 429.800 120.400 ;
        RECT 433.200 111.800 434.000 120.400 ;
        RECT 436.000 111.800 436.800 120.400 ;
        RECT 441.200 112.200 442.000 120.400 ;
        RECT 445.000 115.800 445.800 120.400 ;
        RECT 449.200 111.800 450.000 120.400 ;
        RECT 451.400 115.800 452.200 120.400 ;
        RECT 455.600 111.800 456.400 120.400 ;
        RECT 462.000 115.800 462.800 120.400 ;
        RECT 465.200 115.800 466.000 120.400 ;
        RECT 468.400 115.800 469.200 120.400 ;
        RECT 471.600 115.800 472.400 120.400 ;
        RECT 473.200 115.800 474.000 120.400 ;
        RECT 476.400 115.800 477.200 120.400 ;
        RECT 478.000 111.800 478.800 120.400 ;
        RECT 483.400 115.800 484.200 120.400 ;
        RECT 487.600 111.800 488.400 120.400 ;
        RECT 489.200 115.800 490.000 120.400 ;
        RECT 492.400 115.800 493.200 120.400 ;
        RECT 494.000 111.800 494.800 120.400 ;
        RECT 498.200 115.800 499.000 120.400 ;
        RECT 500.400 115.800 501.200 120.400 ;
        RECT 503.600 115.800 504.400 120.400 ;
        RECT 506.800 115.800 507.600 120.400 ;
        RECT 508.400 111.800 509.200 120.400 ;
        RECT 512.600 115.800 513.400 120.400 ;
        RECT 516.000 111.800 516.800 120.400 ;
        RECT 521.200 112.200 522.000 120.400 ;
        RECT 524.400 111.800 525.200 120.400 ;
        RECT 528.600 115.800 529.400 120.400 ;
        RECT 531.400 115.800 532.200 120.400 ;
        RECT 535.600 111.800 536.400 120.400 ;
        RECT 538.800 111.800 539.600 120.400 ;
        RECT 544.400 115.800 545.200 120.400 ;
        RECT 547.600 115.800 548.400 120.400 ;
        RECT 553.200 112.000 554.000 120.400 ;
        RECT 558.000 113.000 558.800 120.400 ;
        RECT 561.200 111.800 562.000 120.400 ;
        RECT 562.800 111.800 563.600 120.400 ;
        RECT 567.000 115.800 567.800 120.400 ;
        RECT 569.200 115.800 570.000 120.400 ;
        RECT 572.400 115.800 573.200 120.400 ;
        RECT 575.600 115.800 576.400 120.400 ;
        RECT 578.800 115.800 579.600 120.400 ;
        RECT 586.800 115.800 587.600 120.400 ;
        RECT 590.000 115.800 590.800 120.400 ;
        RECT 596.400 115.800 597.200 120.400 ;
        RECT 599.600 115.800 600.400 120.400 ;
        RECT 602.800 115.800 603.600 120.400 ;
        RECT 605.000 115.800 605.800 120.400 ;
        RECT 596.200 111.800 597.200 112.000 ;
        RECT 599.600 111.800 600.400 112.400 ;
        RECT 609.200 111.800 610.000 120.400 ;
        RECT 317.400 111.200 344.400 111.800 ;
        RECT 374.000 111.200 401.000 111.800 ;
        RECT 317.400 111.000 318.200 111.200 ;
        RECT 400.200 111.000 401.000 111.200 ;
        RECT 573.400 111.200 600.400 111.800 ;
        RECT 573.400 111.000 574.200 111.200 ;
        RECT 245.800 110.000 269.200 110.600 ;
        RECT 245.800 109.800 246.600 110.000 ;
        RECT 250.800 109.600 251.600 110.000 ;
        RECT 268.400 109.400 269.200 110.000 ;
        RECT 340.400 92.000 341.200 92.600 ;
        RECT 358.000 92.000 358.800 92.400 ;
        RECT 363.000 92.000 363.800 92.200 ;
        RECT 340.400 91.400 363.800 92.000 ;
        RECT 206.600 90.800 207.400 91.000 ;
        RECT 180.400 90.200 207.400 90.800 ;
        RECT 253.400 90.800 254.200 91.000 ;
        RECT 313.800 90.800 314.600 91.000 ;
        RECT 395.400 90.800 396.200 91.000 ;
        RECT 605.000 90.800 605.800 91.000 ;
        RECT 253.400 90.200 280.400 90.800 ;
        RECT 2.800 81.600 3.600 90.200 ;
        RECT 8.400 81.600 9.200 86.200 ;
        RECT 11.600 81.600 12.400 86.200 ;
        RECT 17.200 81.600 18.000 90.000 ;
        RECT 21.000 81.600 21.800 86.200 ;
        RECT 25.200 81.600 26.000 90.200 ;
        RECT 26.800 81.600 27.600 90.200 ;
        RECT 31.000 81.600 31.800 86.200 ;
        RECT 34.400 81.600 35.200 90.200 ;
        RECT 39.600 81.600 40.400 89.800 ;
        RECT 43.400 81.600 44.200 86.200 ;
        RECT 47.600 81.600 48.400 90.200 ;
        RECT 50.800 81.600 51.600 90.000 ;
        RECT 56.400 81.600 57.200 86.200 ;
        RECT 59.600 81.600 60.400 86.200 ;
        RECT 65.200 81.600 66.000 90.200 ;
        RECT 69.000 81.600 69.800 86.200 ;
        RECT 73.200 81.600 74.000 90.200 ;
        RECT 76.400 81.600 77.200 89.800 ;
        RECT 81.600 81.600 82.400 90.200 ;
        RECT 85.000 81.600 85.800 86.200 ;
        RECT 89.200 81.600 90.000 90.200 ;
        RECT 90.800 81.600 91.600 86.200 ;
        RECT 94.000 81.600 94.800 85.800 ;
        RECT 97.800 81.600 98.600 86.200 ;
        RECT 102.000 81.600 102.800 90.200 ;
        RECT 103.600 81.600 104.400 86.200 ;
        RECT 106.800 81.600 107.600 85.800 ;
        RECT 113.200 81.600 114.000 90.200 ;
        RECT 115.400 81.600 116.200 86.200 ;
        RECT 119.600 81.600 120.400 90.200 ;
        RECT 121.200 81.600 122.000 86.200 ;
        RECT 124.400 81.600 125.200 86.200 ;
        RECT 127.200 81.600 128.000 90.200 ;
        RECT 132.400 81.600 133.200 89.800 ;
        RECT 135.600 81.600 136.400 90.200 ;
        RECT 139.800 81.600 140.600 86.200 ;
        RECT 142.000 81.600 142.800 86.200 ;
        RECT 145.200 81.600 146.000 86.200 ;
        RECT 148.400 81.600 149.200 85.800 ;
        RECT 151.600 81.600 152.400 86.200 ;
        RECT 159.600 81.600 160.400 90.200 ;
        RECT 165.200 81.600 166.000 86.200 ;
        RECT 168.400 81.600 169.200 86.200 ;
        RECT 174.000 81.600 174.800 90.000 ;
        RECT 180.400 89.600 181.200 90.200 ;
        RECT 183.600 90.000 184.600 90.200 ;
        RECT 177.200 81.600 178.000 86.200 ;
        RECT 180.400 81.600 181.200 86.200 ;
        RECT 183.600 81.600 184.400 86.200 ;
        RECT 190.000 81.600 190.800 86.200 ;
        RECT 193.200 81.600 194.000 86.200 ;
        RECT 201.200 81.600 202.000 86.200 ;
        RECT 204.400 81.600 205.200 86.200 ;
        RECT 207.600 81.600 208.400 86.200 ;
        RECT 210.800 81.600 211.600 86.200 ;
        RECT 213.000 81.600 213.800 86.200 ;
        RECT 217.200 81.600 218.000 90.200 ;
        RECT 218.800 81.600 219.600 86.200 ;
        RECT 222.000 81.600 222.800 86.200 ;
        RECT 223.600 81.600 224.400 86.200 ;
        RECT 226.800 81.600 227.600 86.200 ;
        RECT 230.000 81.600 230.800 89.800 ;
        RECT 233.200 81.600 234.000 86.200 ;
        RECT 234.800 81.600 235.600 86.200 ;
        RECT 238.000 81.600 238.800 86.200 ;
        RECT 239.600 81.600 240.400 90.200 ;
        RECT 276.200 90.000 277.200 90.200 ;
        RECT 279.600 89.600 280.400 90.200 ;
        RECT 287.600 90.200 314.600 90.800 ;
        RECT 369.200 90.200 396.200 90.800 ;
        RECT 578.800 90.200 605.800 90.800 ;
        RECT 287.600 89.600 288.400 90.200 ;
        RECT 291.000 90.000 291.800 90.200 ;
        RECT 243.800 81.600 244.600 86.200 ;
        RECT 246.000 81.600 246.800 86.200 ;
        RECT 249.200 81.600 250.000 86.200 ;
        RECT 252.400 81.600 253.200 86.200 ;
        RECT 255.600 81.600 256.400 86.200 ;
        RECT 258.800 81.600 259.600 86.200 ;
        RECT 266.800 81.600 267.600 86.200 ;
        RECT 270.000 81.600 270.800 86.200 ;
        RECT 276.400 81.600 277.200 86.200 ;
        RECT 279.600 81.600 280.400 86.200 ;
        RECT 282.800 81.600 283.600 86.200 ;
        RECT 284.400 81.600 285.200 86.200 ;
        RECT 287.600 81.600 288.400 86.200 ;
        RECT 290.800 81.600 291.600 86.200 ;
        RECT 297.200 81.600 298.000 86.200 ;
        RECT 300.400 81.600 301.200 86.200 ;
        RECT 308.400 81.600 309.200 86.200 ;
        RECT 311.600 81.600 312.400 86.200 ;
        RECT 314.800 81.600 315.600 86.200 ;
        RECT 318.000 81.600 318.800 86.200 ;
        RECT 324.400 81.600 325.200 90.200 ;
        RECT 369.200 89.600 370.000 90.200 ;
        RECT 372.400 90.000 373.400 90.200 ;
        RECT 327.600 81.600 328.400 89.000 ;
        RECT 330.800 81.600 331.600 86.200 ;
        RECT 334.000 81.600 334.800 86.200 ;
        RECT 337.200 81.600 338.000 86.200 ;
        RECT 340.400 81.600 341.200 86.200 ;
        RECT 348.400 81.600 349.200 86.200 ;
        RECT 351.600 81.600 352.400 86.200 ;
        RECT 358.000 81.600 358.800 86.200 ;
        RECT 361.200 81.600 362.000 86.200 ;
        RECT 364.400 81.600 365.200 86.200 ;
        RECT 366.000 81.600 366.800 86.200 ;
        RECT 369.200 81.600 370.000 86.200 ;
        RECT 372.400 81.600 373.200 86.200 ;
        RECT 378.800 81.600 379.600 86.200 ;
        RECT 382.000 81.600 382.800 86.200 ;
        RECT 390.000 81.600 390.800 86.200 ;
        RECT 393.200 81.600 394.000 86.200 ;
        RECT 396.400 81.600 397.200 86.200 ;
        RECT 399.600 81.600 400.400 86.200 ;
        RECT 401.800 81.600 402.600 86.200 ;
        RECT 406.000 81.600 406.800 90.200 ;
        RECT 407.600 81.600 408.400 86.200 ;
        RECT 410.800 81.600 411.600 90.200 ;
        RECT 415.000 81.600 415.800 86.200 ;
        RECT 418.400 81.600 419.200 90.200 ;
        RECT 423.600 81.600 424.400 89.800 ;
        RECT 430.000 81.600 430.800 90.200 ;
        RECT 431.600 81.600 432.400 90.200 ;
        RECT 434.800 81.600 435.600 89.000 ;
        RECT 438.000 81.600 438.800 90.200 ;
        RECT 442.200 81.600 443.000 86.200 ;
        RECT 447.600 81.600 448.400 90.200 ;
        RECT 449.800 81.600 450.600 86.200 ;
        RECT 454.000 81.600 454.800 90.200 ;
        RECT 455.600 81.600 456.400 86.200 ;
        RECT 458.800 81.600 459.600 86.200 ;
        RECT 466.800 81.600 467.600 89.800 ;
        RECT 472.000 81.600 472.800 90.200 ;
        RECT 476.400 81.600 477.200 86.200 ;
        RECT 478.000 81.600 478.800 90.200 ;
        RECT 481.200 81.600 482.000 89.000 ;
        RECT 486.000 81.600 486.800 89.000 ;
        RECT 489.200 81.600 490.000 90.200 ;
        RECT 490.800 81.600 491.600 90.200 ;
        RECT 495.000 81.600 495.800 86.200 ;
        RECT 498.800 81.600 499.600 89.800 ;
        RECT 504.000 81.600 504.800 90.200 ;
        RECT 508.400 81.600 509.200 89.000 ;
        RECT 511.600 81.600 512.400 90.200 ;
        RECT 513.200 81.600 514.000 86.200 ;
        RECT 516.400 81.600 517.200 86.200 ;
        RECT 519.600 81.600 520.400 89.800 ;
        RECT 524.800 81.600 525.600 90.200 ;
        RECT 527.600 81.600 528.400 90.200 ;
        RECT 531.800 81.600 532.600 86.200 ;
        RECT 534.600 81.600 535.400 86.200 ;
        RECT 538.800 81.600 539.600 90.200 ;
        RECT 540.400 81.600 541.200 86.200 ;
        RECT 543.600 81.600 544.400 86.200 ;
        RECT 546.800 81.600 547.600 90.200 ;
        RECT 552.400 81.600 553.200 86.200 ;
        RECT 555.600 81.600 556.400 86.200 ;
        RECT 561.200 81.600 562.000 90.000 ;
        RECT 564.400 81.600 565.200 86.200 ;
        RECT 567.600 81.600 568.400 86.200 ;
        RECT 569.200 81.600 570.000 90.200 ;
        RECT 578.800 89.600 579.600 90.200 ;
        RECT 582.000 90.000 583.000 90.200 ;
        RECT 573.400 81.600 574.200 86.200 ;
        RECT 575.600 81.600 576.400 86.200 ;
        RECT 578.800 81.600 579.600 86.200 ;
        RECT 582.000 81.600 582.800 86.200 ;
        RECT 588.400 81.600 589.200 86.200 ;
        RECT 591.600 81.600 592.400 86.200 ;
        RECT 599.600 81.600 600.400 86.200 ;
        RECT 602.800 81.600 603.600 86.200 ;
        RECT 606.000 81.600 606.800 86.200 ;
        RECT 609.200 81.600 610.000 86.200 ;
        RECT 0.400 80.400 614.000 81.600 ;
        RECT 1.200 75.800 2.000 80.400 ;
        RECT 4.400 71.800 5.200 80.400 ;
        RECT 8.600 75.800 9.400 80.400 ;
        RECT 11.400 75.800 12.200 80.400 ;
        RECT 15.600 71.800 16.400 80.400 ;
        RECT 17.200 75.800 18.000 80.400 ;
        RECT 20.400 75.800 21.200 80.400 ;
        RECT 23.200 71.800 24.000 80.400 ;
        RECT 28.400 72.200 29.200 80.400 ;
        RECT 31.600 71.800 32.400 80.400 ;
        RECT 35.800 75.800 36.600 80.400 ;
        RECT 38.600 75.800 39.400 80.400 ;
        RECT 42.800 71.800 43.600 80.400 ;
        RECT 46.000 72.000 46.800 80.400 ;
        RECT 51.600 75.800 52.400 80.400 ;
        RECT 54.800 75.800 55.600 80.400 ;
        RECT 60.400 71.800 61.200 80.400 ;
        RECT 63.600 71.800 64.400 80.400 ;
        RECT 67.800 75.800 68.600 80.400 ;
        RECT 70.000 71.800 70.800 80.400 ;
        RECT 74.200 75.800 75.000 80.400 ;
        RECT 77.000 75.800 77.800 80.400 ;
        RECT 81.200 71.800 82.000 80.400 ;
        RECT 84.400 72.200 85.200 80.400 ;
        RECT 89.600 71.800 90.400 80.400 ;
        RECT 92.400 71.800 93.200 80.400 ;
        RECT 95.600 73.000 96.400 80.400 ;
        RECT 98.800 75.800 99.600 80.400 ;
        RECT 102.000 75.800 102.800 80.400 ;
        RECT 105.200 75.800 106.000 80.400 ;
        RECT 110.000 71.800 110.800 80.400 ;
        RECT 115.600 75.800 116.400 80.400 ;
        RECT 118.800 75.800 119.600 80.400 ;
        RECT 124.400 72.000 125.200 80.400 ;
        RECT 129.200 75.800 130.000 80.400 ;
        RECT 130.800 75.800 131.600 80.400 ;
        RECT 135.600 73.000 136.400 80.400 ;
        RECT 138.800 71.800 139.600 80.400 ;
        RECT 140.400 71.800 141.200 80.400 ;
        RECT 144.600 75.800 145.400 80.400 ;
        RECT 147.400 75.800 148.200 80.400 ;
        RECT 151.600 71.800 152.400 80.400 ;
        RECT 159.600 72.000 160.400 80.400 ;
        RECT 165.200 75.800 166.000 80.400 ;
        RECT 168.400 75.800 169.200 80.400 ;
        RECT 174.000 71.800 174.800 80.400 ;
        RECT 177.200 71.800 178.000 80.400 ;
        RECT 181.400 75.800 182.200 80.400 ;
        RECT 184.200 75.800 185.000 80.400 ;
        RECT 188.400 71.800 189.200 80.400 ;
        RECT 191.600 72.200 192.400 80.400 ;
        RECT 196.800 71.800 197.600 80.400 ;
        RECT 199.600 75.800 200.400 80.400 ;
        RECT 202.800 75.800 203.600 80.400 ;
        RECT 204.400 75.800 205.200 80.400 ;
        RECT 207.600 75.800 208.400 80.400 ;
        RECT 210.800 75.800 211.600 80.400 ;
        RECT 217.200 75.800 218.000 80.400 ;
        RECT 220.400 75.800 221.200 80.400 ;
        RECT 228.400 75.800 229.200 80.400 ;
        RECT 231.600 75.800 232.400 80.400 ;
        RECT 234.800 75.800 235.600 80.400 ;
        RECT 238.000 75.800 238.800 80.400 ;
        RECT 240.200 75.800 241.000 80.400 ;
        RECT 207.600 71.800 208.400 72.400 ;
        RECT 211.000 71.800 211.800 72.000 ;
        RECT 244.400 71.800 245.200 80.400 ;
        RECT 246.000 71.800 246.800 80.400 ;
        RECT 250.200 75.800 251.000 80.400 ;
        RECT 252.400 75.800 253.200 80.400 ;
        RECT 255.600 75.800 256.400 80.400 ;
        RECT 257.200 75.800 258.000 80.400 ;
        RECT 260.400 75.800 261.200 80.400 ;
        RECT 263.600 75.800 264.400 80.400 ;
        RECT 266.800 75.800 267.600 80.400 ;
        RECT 274.800 75.800 275.600 80.400 ;
        RECT 278.000 75.800 278.800 80.400 ;
        RECT 284.400 75.800 285.200 80.400 ;
        RECT 287.600 75.800 288.400 80.400 ;
        RECT 290.800 75.800 291.600 80.400 ;
        RECT 292.400 75.800 293.200 80.400 ;
        RECT 295.600 75.800 296.400 80.400 ;
        RECT 302.000 75.800 302.800 80.400 ;
        RECT 305.200 75.800 306.000 80.400 ;
        RECT 308.400 75.800 309.200 80.400 ;
        RECT 311.600 75.800 312.400 80.400 ;
        RECT 319.600 75.800 320.400 80.400 ;
        RECT 322.800 75.800 323.600 80.400 ;
        RECT 329.200 75.800 330.000 80.400 ;
        RECT 332.400 75.800 333.200 80.400 ;
        RECT 335.600 75.800 336.400 80.400 ;
        RECT 284.200 71.800 285.200 72.000 ;
        RECT 287.600 71.800 288.400 72.400 ;
        RECT 329.000 71.800 329.800 72.000 ;
        RECT 332.400 71.800 333.200 72.400 ;
        RECT 337.200 71.800 338.000 80.400 ;
        RECT 341.400 75.800 342.200 80.400 ;
        RECT 345.400 79.800 346.200 80.400 ;
        RECT 345.200 73.200 346.200 79.800 ;
        RECT 351.400 73.200 352.400 80.400 ;
        RECT 355.400 75.800 356.200 80.400 ;
        RECT 359.600 71.800 360.400 80.400 ;
        RECT 361.200 75.800 362.000 80.400 ;
        RECT 364.400 75.800 365.200 80.400 ;
        RECT 368.600 71.800 369.400 80.400 ;
        RECT 372.400 71.800 373.200 80.400 ;
        RECT 377.200 71.800 378.000 80.400 ;
        RECT 381.400 75.800 382.200 80.400 ;
        RECT 383.600 75.800 384.400 80.400 ;
        RECT 386.800 75.800 387.600 80.400 ;
        RECT 388.400 71.800 389.200 80.400 ;
        RECT 392.600 75.800 393.400 80.400 ;
        RECT 396.600 79.800 397.400 80.400 ;
        RECT 396.400 73.200 397.400 79.800 ;
        RECT 402.600 73.200 403.600 80.400 ;
        RECT 406.000 71.800 406.800 80.400 ;
        RECT 409.200 71.800 410.000 80.400 ;
        RECT 413.400 75.800 414.200 80.400 ;
        RECT 415.600 71.800 416.400 80.400 ;
        RECT 419.800 75.800 420.600 80.400 ;
        RECT 422.000 75.800 422.800 80.400 ;
        RECT 425.200 75.800 426.000 80.400 ;
        RECT 426.800 75.800 427.600 80.400 ;
        RECT 430.000 76.200 430.800 80.400 ;
        RECT 433.200 71.800 434.000 80.400 ;
        RECT 436.400 73.000 437.200 80.400 ;
        RECT 439.600 71.800 440.400 80.400 ;
        RECT 443.800 75.800 444.600 80.400 ;
        RECT 446.600 75.800 447.400 80.400 ;
        RECT 450.800 71.800 451.600 80.400 ;
        RECT 453.000 75.800 453.800 80.400 ;
        RECT 457.200 71.800 458.000 80.400 ;
        RECT 465.200 71.800 466.000 80.400 ;
        RECT 470.800 75.800 471.600 80.400 ;
        RECT 474.000 75.800 474.800 80.400 ;
        RECT 479.600 72.000 480.400 80.400 ;
        RECT 482.800 71.800 483.600 80.400 ;
        RECT 487.000 75.800 487.800 80.400 ;
        RECT 489.800 75.800 490.600 80.400 ;
        RECT 494.000 71.800 494.800 80.400 ;
        RECT 495.600 71.800 496.400 80.400 ;
        RECT 499.800 75.800 500.600 80.400 ;
        RECT 502.600 75.800 503.400 80.400 ;
        RECT 506.800 71.800 507.600 80.400 ;
        RECT 508.400 71.800 509.200 80.400 ;
        RECT 512.600 75.800 513.400 80.400 ;
        RECT 516.400 71.800 517.200 80.400 ;
        RECT 522.000 75.800 522.800 80.400 ;
        RECT 525.200 75.800 526.000 80.400 ;
        RECT 530.800 72.000 531.600 80.400 ;
        RECT 534.000 71.800 534.800 80.400 ;
        RECT 538.200 75.800 539.000 80.400 ;
        RECT 540.400 75.800 541.200 80.400 ;
        RECT 543.600 75.800 544.400 80.400 ;
        RECT 545.200 75.800 546.000 80.400 ;
        RECT 548.400 75.800 549.200 80.400 ;
        RECT 551.600 73.000 552.400 80.400 ;
        RECT 554.800 71.800 555.600 80.400 ;
        RECT 556.400 71.800 557.200 80.400 ;
        RECT 560.600 75.800 561.400 80.400 ;
        RECT 564.400 72.200 565.200 80.400 ;
        RECT 569.600 71.800 570.400 80.400 ;
        RECT 573.000 75.800 573.800 80.400 ;
        RECT 577.200 71.800 578.000 80.400 ;
        RECT 580.400 72.000 581.200 80.400 ;
        RECT 586.000 75.800 586.800 80.400 ;
        RECT 589.200 75.800 590.000 80.400 ;
        RECT 594.800 71.800 595.600 80.400 ;
        RECT 598.000 75.800 598.800 80.400 ;
        RECT 601.200 75.800 602.000 80.400 ;
        RECT 603.400 75.800 604.200 80.400 ;
        RECT 607.600 71.800 608.400 80.400 ;
        RECT 207.600 71.200 234.600 71.800 ;
        RECT 233.800 71.000 234.600 71.200 ;
        RECT 261.400 71.200 288.400 71.800 ;
        RECT 306.200 71.200 333.200 71.800 ;
        RECT 261.400 71.000 262.200 71.200 ;
        RECT 306.200 71.000 307.000 71.200 ;
        RECT 30.600 50.800 31.400 51.000 ;
        RECT 209.800 50.800 210.600 51.000 ;
        RECT 272.200 50.800 273.000 51.000 ;
        RECT 325.000 50.800 325.800 51.000 ;
        RECT 401.800 50.800 402.600 51.000 ;
        RECT 4.400 50.200 31.400 50.800 ;
        RECT 183.600 50.200 210.600 50.800 ;
        RECT 246.000 50.200 273.000 50.800 ;
        RECT 298.800 50.200 325.800 50.800 ;
        RECT 375.600 50.200 402.600 50.800 ;
        RECT 581.400 50.800 582.200 51.000 ;
        RECT 581.400 50.200 608.400 50.800 ;
        RECT 4.400 49.600 5.200 50.200 ;
        RECT 7.800 50.000 8.600 50.200 ;
        RECT 1.200 41.600 2.000 46.200 ;
        RECT 4.400 41.600 5.200 46.200 ;
        RECT 7.600 41.600 8.400 46.200 ;
        RECT 14.000 41.600 14.800 46.200 ;
        RECT 17.200 41.600 18.000 46.200 ;
        RECT 25.200 41.600 26.000 46.200 ;
        RECT 28.400 41.600 29.200 46.200 ;
        RECT 31.600 41.600 32.400 46.200 ;
        RECT 34.800 41.600 35.600 46.200 ;
        RECT 36.400 41.600 37.200 50.200 ;
        RECT 40.600 41.600 41.400 46.200 ;
        RECT 42.800 41.600 43.600 46.200 ;
        RECT 46.000 41.600 46.800 46.200 ;
        RECT 47.600 41.600 48.400 50.200 ;
        RECT 50.800 41.600 51.600 50.200 ;
        RECT 54.000 41.600 54.800 50.200 ;
        RECT 57.200 41.600 58.000 50.200 ;
        RECT 60.400 41.600 61.200 50.200 ;
        RECT 63.200 41.600 64.000 50.200 ;
        RECT 68.400 41.600 69.200 49.800 ;
        RECT 71.600 41.600 72.400 46.200 ;
        RECT 74.800 41.600 75.600 46.200 ;
        RECT 78.000 41.600 78.800 49.800 ;
        RECT 83.200 41.600 84.000 50.200 ;
        RECT 87.200 41.600 88.000 50.200 ;
        RECT 92.400 41.600 93.200 49.800 ;
        RECT 95.600 41.600 96.400 46.200 ;
        RECT 98.800 41.600 99.600 50.200 ;
        RECT 102.000 41.600 102.800 50.200 ;
        RECT 105.200 41.600 106.000 50.200 ;
        RECT 108.400 41.600 109.200 50.200 ;
        RECT 111.600 41.600 112.400 50.200 ;
        RECT 114.400 41.600 115.200 50.200 ;
        RECT 119.600 41.600 120.400 49.800 ;
        RECT 124.400 41.600 125.200 49.800 ;
        RECT 129.600 41.600 130.400 50.200 ;
        RECT 132.400 41.600 133.200 50.200 ;
        RECT 135.600 41.600 136.400 49.000 ;
        RECT 140.000 41.600 140.800 50.200 ;
        RECT 145.200 41.600 146.000 49.800 ;
        RECT 153.200 41.600 154.000 50.200 ;
        RECT 157.400 41.600 158.200 46.200 ;
        RECT 160.200 41.600 161.000 46.200 ;
        RECT 164.400 41.600 165.200 50.200 ;
        RECT 166.000 41.600 166.800 50.200 ;
        RECT 169.200 41.600 170.000 50.200 ;
        RECT 172.400 41.600 173.200 50.200 ;
        RECT 175.600 41.600 176.400 50.200 ;
        RECT 178.800 41.600 179.600 50.200 ;
        RECT 183.600 49.600 184.400 50.200 ;
        RECT 187.000 50.000 187.800 50.200 ;
        RECT 180.400 41.600 181.200 46.200 ;
        RECT 183.600 41.600 184.400 46.200 ;
        RECT 186.800 41.600 187.600 46.200 ;
        RECT 193.200 41.600 194.000 46.200 ;
        RECT 196.400 41.600 197.200 46.200 ;
        RECT 204.400 41.600 205.200 46.200 ;
        RECT 207.600 41.600 208.400 46.200 ;
        RECT 210.800 41.600 211.600 46.200 ;
        RECT 214.000 41.600 214.800 46.200 ;
        RECT 215.600 41.600 216.400 46.200 ;
        RECT 218.800 41.600 219.600 46.200 ;
        RECT 222.000 41.600 222.800 46.200 ;
        RECT 223.600 41.600 224.400 46.200 ;
        RECT 226.800 41.600 227.600 46.200 ;
        RECT 228.400 41.600 229.200 46.200 ;
        RECT 231.600 41.600 232.400 46.200 ;
        RECT 233.800 41.600 234.600 46.200 ;
        RECT 238.000 41.600 238.800 50.200 ;
        RECT 246.000 49.600 246.800 50.200 ;
        RECT 249.400 50.000 250.200 50.200 ;
        RECT 241.200 41.600 242.000 46.200 ;
        RECT 242.800 41.600 243.600 46.200 ;
        RECT 246.000 41.600 246.800 46.200 ;
        RECT 249.200 41.600 250.000 46.200 ;
        RECT 255.600 41.600 256.400 46.200 ;
        RECT 258.800 41.600 259.600 46.200 ;
        RECT 266.800 41.600 267.600 46.200 ;
        RECT 270.000 41.600 270.800 46.200 ;
        RECT 273.200 41.600 274.000 46.200 ;
        RECT 276.400 41.600 277.200 46.200 ;
        RECT 278.000 41.600 278.800 50.200 ;
        RECT 282.200 41.600 283.000 46.200 ;
        RECT 285.000 41.600 285.800 46.200 ;
        RECT 289.200 41.600 290.000 50.200 ;
        RECT 298.800 49.600 299.600 50.200 ;
        RECT 302.000 50.000 303.000 50.200 ;
        RECT 295.600 41.600 296.400 46.200 ;
        RECT 298.800 41.600 299.600 46.200 ;
        RECT 302.000 41.600 302.800 46.200 ;
        RECT 308.400 41.600 309.200 46.200 ;
        RECT 311.600 41.600 312.400 46.200 ;
        RECT 319.600 41.600 320.400 46.200 ;
        RECT 322.800 41.600 323.600 46.200 ;
        RECT 326.000 41.600 326.800 46.200 ;
        RECT 329.200 41.600 330.000 46.200 ;
        RECT 332.000 41.600 332.800 50.200 ;
        RECT 337.200 41.600 338.000 49.800 ;
        RECT 340.400 41.600 341.200 46.200 ;
        RECT 343.600 41.600 344.400 46.200 ;
        RECT 345.200 41.600 346.000 46.200 ;
        RECT 348.400 41.600 349.200 46.200 ;
        RECT 351.600 41.600 352.400 49.000 ;
        RECT 356.400 41.600 357.200 50.200 ;
        RECT 360.600 41.600 361.400 46.200 ;
        RECT 362.800 41.600 363.600 46.200 ;
        RECT 366.000 41.600 366.800 49.800 ;
        RECT 375.600 49.600 376.400 50.200 ;
        RECT 378.800 50.000 379.800 50.200 ;
        RECT 369.200 41.600 370.000 46.200 ;
        RECT 372.400 41.600 373.200 46.200 ;
        RECT 375.600 41.600 376.400 46.200 ;
        RECT 378.800 41.600 379.600 46.200 ;
        RECT 385.200 41.600 386.000 46.200 ;
        RECT 388.400 41.600 389.200 46.200 ;
        RECT 396.400 41.600 397.200 46.200 ;
        RECT 399.600 41.600 400.400 46.200 ;
        RECT 402.800 41.600 403.600 46.200 ;
        RECT 406.000 41.600 406.800 46.200 ;
        RECT 409.200 41.600 410.000 50.000 ;
        RECT 414.800 41.600 415.600 46.200 ;
        RECT 418.000 41.600 418.800 46.200 ;
        RECT 423.600 41.600 424.400 50.200 ;
        RECT 426.800 41.600 427.600 46.200 ;
        RECT 430.000 41.600 430.800 50.200 ;
        RECT 434.200 41.600 435.000 46.200 ;
        RECT 437.000 41.600 437.800 46.200 ;
        RECT 441.200 41.600 442.000 50.200 ;
        RECT 443.400 41.600 444.200 46.200 ;
        RECT 447.600 41.600 448.400 50.200 ;
        RECT 450.400 41.600 451.200 50.200 ;
        RECT 455.600 41.600 456.400 49.800 ;
        RECT 464.200 41.600 465.000 46.200 ;
        RECT 468.400 41.600 469.200 50.200 ;
        RECT 471.600 41.600 472.400 46.200 ;
        RECT 474.800 41.600 475.600 49.800 ;
        RECT 480.000 41.600 480.800 50.200 ;
        RECT 484.400 41.600 485.200 50.000 ;
        RECT 490.000 41.600 490.800 46.200 ;
        RECT 493.200 41.600 494.000 46.200 ;
        RECT 498.800 41.600 499.600 50.200 ;
        RECT 502.000 41.600 502.800 46.200 ;
        RECT 506.800 41.600 507.600 49.800 ;
        RECT 512.000 41.600 512.800 50.200 ;
        RECT 514.800 41.600 515.600 50.200 ;
        RECT 518.000 41.600 518.800 49.000 ;
        RECT 522.400 41.600 523.200 50.200 ;
        RECT 527.600 41.600 528.400 49.800 ;
        RECT 530.800 41.600 531.600 50.200 ;
        RECT 535.000 41.600 535.800 46.200 ;
        RECT 537.800 41.600 538.600 46.200 ;
        RECT 542.000 41.600 542.800 50.200 ;
        RECT 545.200 41.600 546.000 50.200 ;
        RECT 550.800 41.600 551.600 46.200 ;
        RECT 554.000 41.600 554.800 46.200 ;
        RECT 559.600 41.600 560.400 50.000 ;
        RECT 562.800 41.600 563.600 50.200 ;
        RECT 566.000 41.600 566.800 50.200 ;
        RECT 569.200 41.600 570.000 50.200 ;
        RECT 572.400 41.600 573.200 50.200 ;
        RECT 575.600 41.600 576.400 50.200 ;
        RECT 604.200 50.000 605.200 50.200 ;
        RECT 607.600 49.600 608.400 50.200 ;
        RECT 577.200 41.600 578.000 46.200 ;
        RECT 580.400 41.600 581.200 46.200 ;
        RECT 583.600 41.600 584.400 46.200 ;
        RECT 586.800 41.600 587.600 46.200 ;
        RECT 594.800 41.600 595.600 46.200 ;
        RECT 598.000 41.600 598.800 46.200 ;
        RECT 604.400 41.600 605.200 46.200 ;
        RECT 607.600 41.600 608.400 46.200 ;
        RECT 610.800 41.600 611.600 46.200 ;
        RECT 0.400 40.400 614.000 41.600 ;
        RECT 2.800 33.000 3.600 40.400 ;
        RECT 6.000 35.800 6.800 40.400 ;
        RECT 9.200 35.800 10.000 40.400 ;
        RECT 12.400 35.800 13.200 40.400 ;
        RECT 18.800 35.800 19.600 40.400 ;
        RECT 22.000 35.800 22.800 40.400 ;
        RECT 30.000 35.800 30.800 40.400 ;
        RECT 33.200 35.800 34.000 40.400 ;
        RECT 36.400 35.800 37.200 40.400 ;
        RECT 39.600 35.800 40.400 40.400 ;
        RECT 41.800 35.800 42.600 40.400 ;
        RECT 9.200 31.800 10.000 32.400 ;
        RECT 12.600 31.800 13.400 32.000 ;
        RECT 46.000 31.800 46.800 40.400 ;
        RECT 49.200 35.800 50.000 40.400 ;
        RECT 50.800 31.800 51.600 40.400 ;
        RECT 55.000 35.800 55.800 40.400 ;
        RECT 57.800 35.800 58.600 40.400 ;
        RECT 62.000 31.800 62.800 40.400 ;
        RECT 65.200 31.800 66.000 40.400 ;
        RECT 70.800 35.800 71.600 40.400 ;
        RECT 74.000 35.800 74.800 40.400 ;
        RECT 79.600 32.000 80.400 40.400 ;
        RECT 82.800 31.800 83.600 40.400 ;
        RECT 87.000 35.800 87.800 40.400 ;
        RECT 89.800 35.800 90.600 40.400 ;
        RECT 94.000 31.800 94.800 40.400 ;
        RECT 97.200 32.000 98.000 40.400 ;
        RECT 102.800 35.800 103.600 40.400 ;
        RECT 106.000 35.800 106.800 40.400 ;
        RECT 111.600 31.800 112.400 40.400 ;
        RECT 114.800 31.800 115.600 40.400 ;
        RECT 119.000 35.800 119.800 40.400 ;
        RECT 121.800 35.800 122.600 40.400 ;
        RECT 126.000 31.800 126.800 40.400 ;
        RECT 127.600 31.800 128.400 40.400 ;
        RECT 131.800 35.800 132.600 40.400 ;
        RECT 134.600 35.800 135.400 40.400 ;
        RECT 138.800 31.800 139.600 40.400 ;
        RECT 142.000 31.800 142.800 40.400 ;
        RECT 147.600 35.800 148.400 40.400 ;
        RECT 150.800 35.800 151.600 40.400 ;
        RECT 156.400 32.000 157.200 40.400 ;
        RECT 164.400 35.800 165.200 40.400 ;
        RECT 167.600 31.800 168.400 40.400 ;
        RECT 171.800 35.800 172.600 40.400 ;
        RECT 174.000 35.800 174.800 40.400 ;
        RECT 177.200 35.800 178.000 40.400 ;
        RECT 178.800 35.800 179.600 40.400 ;
        RECT 182.000 35.800 182.800 40.400 ;
        RECT 185.200 35.800 186.000 40.400 ;
        RECT 188.400 35.800 189.200 40.400 ;
        RECT 196.400 35.800 197.200 40.400 ;
        RECT 199.600 35.800 200.400 40.400 ;
        RECT 206.000 35.800 206.800 40.400 ;
        RECT 209.200 35.800 210.000 40.400 ;
        RECT 212.400 35.800 213.200 40.400 ;
        RECT 215.600 35.800 216.400 40.400 ;
        RECT 217.800 35.800 218.600 40.400 ;
        RECT 205.800 31.800 206.800 32.000 ;
        RECT 209.200 31.800 210.000 32.400 ;
        RECT 222.000 31.800 222.800 40.400 ;
        RECT 224.200 35.800 225.000 40.400 ;
        RECT 228.400 31.800 229.200 40.400 ;
        RECT 231.600 35.800 232.400 40.400 ;
        RECT 233.200 35.800 234.000 40.400 ;
        RECT 236.400 35.800 237.200 40.400 ;
        RECT 239.600 35.800 240.400 40.400 ;
        RECT 246.000 35.800 246.800 40.400 ;
        RECT 249.200 35.800 250.000 40.400 ;
        RECT 257.200 35.800 258.000 40.400 ;
        RECT 260.400 35.800 261.200 40.400 ;
        RECT 263.600 35.800 264.400 40.400 ;
        RECT 266.800 35.800 267.600 40.400 ;
        RECT 268.400 35.800 269.200 40.400 ;
        RECT 271.600 35.800 272.400 40.400 ;
        RECT 274.800 35.800 275.600 40.400 ;
        RECT 278.000 35.800 278.800 40.400 ;
        RECT 284.400 35.800 285.200 40.400 ;
        RECT 287.600 35.800 288.400 40.400 ;
        RECT 295.600 35.800 296.400 40.400 ;
        RECT 298.800 35.800 299.600 40.400 ;
        RECT 302.000 35.800 302.800 40.400 ;
        RECT 305.200 35.800 306.000 40.400 ;
        RECT 311.600 35.800 312.400 40.400 ;
        RECT 316.400 33.200 317.400 40.400 ;
        RECT 322.600 39.800 323.400 40.400 ;
        RECT 322.600 33.200 323.600 39.800 ;
        RECT 236.400 31.800 237.200 32.400 ;
        RECT 239.600 31.800 240.600 32.000 ;
        RECT 274.800 31.800 275.600 32.400 ;
        RECT 327.600 32.200 328.400 40.400 ;
        RECT 278.000 31.800 279.000 32.000 ;
        RECT 332.800 31.800 333.600 40.400 ;
        RECT 337.400 39.800 338.200 40.400 ;
        RECT 337.200 33.200 338.200 39.800 ;
        RECT 343.400 33.200 344.400 40.400 ;
        RECT 346.800 35.800 347.600 40.400 ;
        RECT 350.000 36.200 350.800 40.400 ;
        RECT 353.200 31.800 354.000 40.400 ;
        RECT 358.000 35.800 358.800 40.400 ;
        RECT 361.200 35.800 362.000 40.400 ;
        RECT 364.400 35.800 365.200 40.400 ;
        RECT 367.600 35.800 368.400 40.400 ;
        RECT 375.600 35.800 376.400 40.400 ;
        RECT 378.800 35.800 379.600 40.400 ;
        RECT 385.200 35.800 386.000 40.400 ;
        RECT 388.400 35.800 389.200 40.400 ;
        RECT 391.600 35.800 392.400 40.400 ;
        RECT 385.000 31.800 385.800 32.000 ;
        RECT 388.400 31.800 389.200 32.400 ;
        RECT 393.200 31.800 394.000 40.400 ;
        RECT 396.400 31.800 397.200 40.400 ;
        RECT 399.600 31.800 400.400 40.400 ;
        RECT 402.800 31.800 403.600 40.400 ;
        RECT 406.000 31.800 406.800 40.400 ;
        RECT 407.600 31.800 408.400 40.400 ;
        RECT 410.800 31.800 411.600 40.400 ;
        RECT 414.000 31.800 414.800 40.400 ;
        RECT 417.200 31.800 418.000 40.400 ;
        RECT 420.400 31.800 421.200 40.400 ;
        RECT 422.000 31.800 422.800 40.400 ;
        RECT 426.200 35.800 427.000 40.400 ;
        RECT 430.000 36.200 430.800 40.400 ;
        RECT 433.200 35.800 434.000 40.400 ;
        RECT 435.400 35.800 436.200 40.400 ;
        RECT 439.600 31.800 440.400 40.400 ;
        RECT 442.800 36.200 443.600 40.400 ;
        RECT 446.000 35.800 446.800 40.400 ;
        RECT 448.200 35.800 449.000 40.400 ;
        RECT 452.400 31.800 453.200 40.400 ;
        RECT 460.400 32.000 461.200 40.400 ;
        RECT 466.000 35.800 466.800 40.400 ;
        RECT 469.200 35.800 470.000 40.400 ;
        RECT 474.800 31.800 475.600 40.400 ;
        RECT 478.000 31.800 478.800 40.400 ;
        RECT 482.200 35.800 483.000 40.400 ;
        RECT 485.000 35.800 485.800 40.400 ;
        RECT 489.200 31.800 490.000 40.400 ;
        RECT 492.400 32.000 493.200 40.400 ;
        RECT 498.000 35.800 498.800 40.400 ;
        RECT 501.200 35.800 502.000 40.400 ;
        RECT 506.800 31.800 507.600 40.400 ;
        RECT 510.000 31.800 510.800 40.400 ;
        RECT 514.200 35.800 515.000 40.400 ;
        RECT 517.000 35.800 517.800 40.400 ;
        RECT 521.200 31.800 522.000 40.400 ;
        RECT 522.800 31.800 523.600 40.400 ;
        RECT 526.000 31.800 526.800 40.400 ;
        RECT 529.200 31.800 530.000 40.400 ;
        RECT 532.400 31.800 533.200 40.400 ;
        RECT 535.600 31.800 536.400 40.400 ;
        RECT 538.800 35.800 539.600 40.400 ;
        RECT 541.000 35.800 541.800 40.400 ;
        RECT 545.200 31.800 546.000 40.400 ;
        RECT 546.800 31.800 547.600 40.400 ;
        RECT 551.000 35.800 551.800 40.400 ;
        RECT 553.800 35.800 554.600 40.400 ;
        RECT 558.000 31.800 558.800 40.400 ;
        RECT 560.200 35.800 561.000 40.400 ;
        RECT 564.400 31.800 565.200 40.400 ;
        RECT 567.600 35.800 568.400 40.400 ;
        RECT 569.200 35.800 570.000 40.400 ;
        RECT 572.400 35.800 573.200 40.400 ;
        RECT 575.600 35.800 576.400 40.400 ;
        RECT 578.800 35.800 579.600 40.400 ;
        RECT 586.800 35.800 587.600 40.400 ;
        RECT 590.000 35.800 590.800 40.400 ;
        RECT 596.400 35.800 597.200 40.400 ;
        RECT 599.600 35.800 600.400 40.400 ;
        RECT 602.800 35.800 603.600 40.400 ;
        RECT 606.000 35.800 606.800 40.400 ;
        RECT 609.200 33.000 610.000 40.400 ;
        RECT 596.200 31.800 597.200 32.000 ;
        RECT 599.600 31.800 600.400 32.400 ;
        RECT 9.200 31.200 36.200 31.800 ;
        RECT 35.400 31.000 36.200 31.200 ;
        RECT 183.000 31.200 210.000 31.800 ;
        RECT 236.400 31.200 263.400 31.800 ;
        RECT 274.800 31.200 301.800 31.800 ;
        RECT 183.000 31.000 183.800 31.200 ;
        RECT 262.600 31.000 263.400 31.200 ;
        RECT 301.000 31.000 301.800 31.200 ;
        RECT 362.200 31.200 389.200 31.800 ;
        RECT 573.400 31.200 600.400 31.800 ;
        RECT 362.200 31.000 363.000 31.200 ;
        RECT 573.400 31.000 574.200 31.200 ;
        RECT 30.600 10.800 31.400 11.000 ;
        RECT 4.400 10.200 31.400 10.800 ;
        RECT 149.400 10.800 150.200 11.000 ;
        RECT 209.800 10.800 210.600 11.000 ;
        RECT 249.800 10.800 250.600 11.000 ;
        RECT 299.400 10.800 300.200 11.000 ;
        RECT 344.200 10.800 345.000 11.000 ;
        RECT 393.800 10.800 394.600 11.000 ;
        RECT 149.400 10.200 176.400 10.800 ;
        RECT 4.400 9.600 5.200 10.200 ;
        RECT 7.800 10.000 8.600 10.200 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 4.400 1.600 5.200 6.200 ;
        RECT 7.600 1.600 8.400 6.200 ;
        RECT 14.000 1.600 14.800 6.200 ;
        RECT 17.200 1.600 18.000 6.200 ;
        RECT 25.200 1.600 26.000 6.200 ;
        RECT 28.400 1.600 29.200 6.200 ;
        RECT 31.600 1.600 32.400 6.200 ;
        RECT 34.800 1.600 35.600 6.200 ;
        RECT 36.400 1.600 37.200 10.200 ;
        RECT 40.600 1.600 41.400 6.200 ;
        RECT 43.400 1.600 44.200 6.200 ;
        RECT 47.600 1.600 48.400 10.200 ;
        RECT 50.800 1.600 51.600 6.200 ;
        RECT 54.000 1.600 54.800 10.000 ;
        RECT 59.600 1.600 60.400 6.200 ;
        RECT 62.800 1.600 63.600 6.200 ;
        RECT 68.400 1.600 69.200 10.200 ;
        RECT 71.600 1.600 72.400 10.200 ;
        RECT 74.800 1.600 75.600 9.000 ;
        RECT 78.000 1.600 78.800 10.200 ;
        RECT 82.200 1.600 83.000 6.200 ;
        RECT 85.000 1.600 85.800 6.200 ;
        RECT 89.200 1.600 90.000 10.200 ;
        RECT 92.400 1.600 93.200 10.200 ;
        RECT 98.000 1.600 98.800 6.200 ;
        RECT 101.200 1.600 102.000 6.200 ;
        RECT 106.800 1.600 107.600 10.000 ;
        RECT 111.600 1.600 112.400 10.200 ;
        RECT 117.200 1.600 118.000 6.200 ;
        RECT 120.400 1.600 121.200 6.200 ;
        RECT 126.000 1.600 126.800 10.000 ;
        RECT 129.200 1.600 130.000 10.200 ;
        RECT 172.200 10.000 173.000 10.200 ;
        RECT 175.600 9.600 176.400 10.200 ;
        RECT 183.600 10.200 210.600 10.800 ;
        RECT 223.600 10.200 250.600 10.800 ;
        RECT 273.200 10.200 300.200 10.800 ;
        RECT 318.000 10.200 345.000 10.800 ;
        RECT 367.600 10.200 394.600 10.800 ;
        RECT 576.600 10.800 577.400 11.000 ;
        RECT 576.600 10.200 603.600 10.800 ;
        RECT 183.600 9.600 184.400 10.200 ;
        RECT 186.800 10.000 187.800 10.200 ;
        RECT 223.600 9.600 224.400 10.200 ;
        RECT 227.000 10.000 227.800 10.200 ;
        RECT 273.200 9.600 274.000 10.200 ;
        RECT 276.400 10.000 277.400 10.200 ;
        RECT 318.000 9.600 318.800 10.200 ;
        RECT 321.200 10.000 322.200 10.200 ;
        RECT 132.400 1.600 133.200 9.000 ;
        RECT 137.200 1.600 138.000 9.000 ;
        RECT 145.200 1.600 146.000 6.200 ;
        RECT 148.400 1.600 149.200 6.200 ;
        RECT 151.600 1.600 152.400 6.200 ;
        RECT 154.800 1.600 155.600 6.200 ;
        RECT 162.800 1.600 163.600 6.200 ;
        RECT 166.000 1.600 166.800 6.200 ;
        RECT 172.400 1.600 173.200 6.200 ;
        RECT 175.600 1.600 176.400 6.200 ;
        RECT 178.800 1.600 179.600 6.200 ;
        RECT 180.400 1.600 181.200 6.200 ;
        RECT 183.600 1.600 184.400 6.200 ;
        RECT 186.800 1.600 187.600 6.200 ;
        RECT 193.200 1.600 194.000 6.200 ;
        RECT 196.400 1.600 197.200 6.200 ;
        RECT 204.400 1.600 205.200 6.200 ;
        RECT 207.600 1.600 208.400 6.200 ;
        RECT 210.800 1.600 211.600 6.200 ;
        RECT 214.000 1.600 214.800 6.200 ;
        RECT 217.200 1.600 218.000 9.000 ;
        RECT 220.400 1.600 221.200 6.200 ;
        RECT 223.600 1.600 224.400 6.200 ;
        RECT 226.800 1.600 227.600 6.200 ;
        RECT 233.200 1.600 234.000 6.200 ;
        RECT 236.400 1.600 237.200 6.200 ;
        RECT 244.400 1.600 245.200 6.200 ;
        RECT 247.600 1.600 248.400 6.200 ;
        RECT 250.800 1.600 251.600 6.200 ;
        RECT 254.000 1.600 254.800 6.200 ;
        RECT 257.200 1.600 258.000 9.000 ;
        RECT 262.000 1.600 262.800 9.000 ;
        RECT 266.800 1.600 267.600 9.000 ;
        RECT 270.000 1.600 270.800 6.200 ;
        RECT 273.200 1.600 274.000 6.200 ;
        RECT 276.400 1.600 277.200 6.200 ;
        RECT 282.800 1.600 283.600 6.200 ;
        RECT 286.000 1.600 286.800 6.200 ;
        RECT 294.000 1.600 294.800 6.200 ;
        RECT 297.200 1.600 298.000 6.200 ;
        RECT 300.400 1.600 301.200 6.200 ;
        RECT 303.600 1.600 304.400 6.200 ;
        RECT 311.600 1.600 312.400 9.000 ;
        RECT 314.800 1.600 315.600 6.200 ;
        RECT 318.000 1.600 318.800 6.200 ;
        RECT 321.200 1.600 322.000 6.200 ;
        RECT 327.600 1.600 328.400 6.200 ;
        RECT 330.800 1.600 331.600 6.200 ;
        RECT 338.800 1.600 339.600 6.200 ;
        RECT 342.000 1.600 342.800 6.200 ;
        RECT 345.200 1.600 346.000 6.200 ;
        RECT 348.400 1.600 349.200 6.200 ;
        RECT 352.600 1.600 353.400 10.200 ;
        RECT 359.600 1.600 360.400 10.200 ;
        RECT 367.600 9.600 368.400 10.200 ;
        RECT 371.000 10.000 371.800 10.200 ;
        RECT 362.800 1.600 363.600 6.200 ;
        RECT 364.400 1.600 365.200 6.200 ;
        RECT 367.600 1.600 368.400 6.200 ;
        RECT 370.800 1.600 371.600 6.200 ;
        RECT 377.200 1.600 378.000 6.200 ;
        RECT 380.400 1.600 381.200 6.200 ;
        RECT 388.400 1.600 389.200 6.200 ;
        RECT 391.600 1.600 392.400 6.200 ;
        RECT 394.800 1.600 395.600 6.200 ;
        RECT 398.000 1.600 398.800 6.200 ;
        RECT 401.200 1.600 402.000 9.000 ;
        RECT 406.000 1.600 406.800 10.000 ;
        RECT 411.600 1.600 412.400 6.200 ;
        RECT 414.800 1.600 415.600 6.200 ;
        RECT 420.400 1.600 421.200 10.200 ;
        RECT 425.200 1.600 426.000 9.800 ;
        RECT 430.400 1.600 431.200 10.200 ;
        RECT 434.800 1.600 435.600 10.200 ;
        RECT 440.400 1.600 441.200 6.200 ;
        RECT 443.600 1.600 444.400 6.200 ;
        RECT 449.200 1.600 450.000 10.000 ;
        RECT 453.000 1.600 453.800 6.200 ;
        RECT 457.200 1.600 458.000 10.200 ;
        RECT 465.200 1.600 466.000 9.800 ;
        RECT 470.400 1.600 471.200 10.200 ;
        RECT 474.400 1.600 475.200 10.200 ;
        RECT 479.600 1.600 480.400 9.800 ;
        RECT 482.800 1.600 483.600 10.200 ;
        RECT 487.000 1.600 487.800 6.200 ;
        RECT 489.800 1.600 490.600 6.200 ;
        RECT 494.000 1.600 494.800 10.200 ;
        RECT 497.200 1.600 498.000 10.000 ;
        RECT 502.800 1.600 503.600 6.200 ;
        RECT 506.000 1.600 506.800 6.200 ;
        RECT 511.600 1.600 512.400 10.200 ;
        RECT 516.000 1.600 516.800 10.200 ;
        RECT 521.200 1.600 522.000 9.800 ;
        RECT 524.400 1.600 525.200 10.200 ;
        RECT 528.600 1.600 529.400 6.200 ;
        RECT 531.400 1.600 532.200 6.200 ;
        RECT 535.600 1.600 536.400 10.200 ;
        RECT 537.200 1.600 538.000 10.200 ;
        RECT 540.400 1.600 541.200 9.000 ;
        RECT 545.200 1.600 546.000 10.200 ;
        RECT 550.800 1.600 551.600 6.200 ;
        RECT 554.000 1.600 554.800 6.200 ;
        RECT 559.600 1.600 560.400 10.000 ;
        RECT 564.400 1.600 565.200 6.200 ;
        RECT 566.000 1.600 566.800 10.200 ;
        RECT 599.400 10.000 600.400 10.200 ;
        RECT 602.800 9.600 603.600 10.200 ;
        RECT 570.200 1.600 571.000 6.200 ;
        RECT 572.400 1.600 573.200 6.200 ;
        RECT 575.600 1.600 576.400 6.200 ;
        RECT 578.800 1.600 579.600 6.200 ;
        RECT 582.000 1.600 582.800 6.200 ;
        RECT 590.000 1.600 590.800 6.200 ;
        RECT 593.200 1.600 594.000 6.200 ;
        RECT 599.600 1.600 600.400 6.200 ;
        RECT 602.800 1.600 603.600 6.200 ;
        RECT 606.000 1.600 606.800 6.200 ;
        RECT 609.200 1.600 610.000 6.200 ;
        RECT 0.400 0.400 614.000 1.600 ;
      LAYER via1 ;
        RECT 150.200 560.600 151.000 561.400 ;
        RECT 151.600 560.600 152.400 561.400 ;
        RECT 153.000 560.600 153.800 561.400 ;
        RECT 457.400 560.600 458.200 561.400 ;
        RECT 458.800 560.600 459.600 561.400 ;
        RECT 460.200 560.600 461.000 561.400 ;
        RECT 7.600 557.600 8.400 558.400 ;
        RECT 7.600 551.600 8.400 552.400 ;
        RECT 95.600 557.600 96.400 558.400 ;
        RECT 95.600 551.600 96.400 552.400 ;
        RECT 146.800 557.600 147.600 558.400 ;
        RECT 146.800 551.600 147.600 552.400 ;
        RECT 206.000 557.600 206.800 558.400 ;
        RECT 206.000 551.600 206.800 552.400 ;
        RECT 260.400 557.600 261.200 558.400 ;
        RECT 332.400 557.600 333.200 558.400 ;
        RECT 260.400 551.600 261.200 552.400 ;
        RECT 332.400 551.600 333.200 552.400 ;
        RECT 396.400 551.200 397.200 552.000 ;
        RECT 585.200 551.200 586.000 552.000 ;
        RECT 7.600 523.600 8.400 524.400 ;
        RECT 94.000 523.600 94.800 524.400 ;
        RECT 170.800 523.600 171.600 524.400 ;
        RECT 182.000 523.600 182.800 524.400 ;
        RECT 255.600 523.600 256.400 524.400 ;
        RECT 263.600 523.600 264.400 524.400 ;
        RECT 342.000 530.000 342.800 530.800 ;
        RECT 342.000 525.400 342.800 526.200 ;
        RECT 409.200 530.000 410.000 530.800 ;
        RECT 409.200 523.600 410.000 524.400 ;
        RECT 574.000 523.600 574.800 524.400 ;
        RECT 150.200 520.600 151.000 521.400 ;
        RECT 151.600 520.600 152.400 521.400 ;
        RECT 153.000 520.600 153.800 521.400 ;
        RECT 457.400 520.600 458.200 521.400 ;
        RECT 458.800 520.600 459.600 521.400 ;
        RECT 460.200 520.600 461.000 521.400 ;
        RECT 202.800 517.600 203.600 518.400 ;
        RECT 202.800 511.600 203.600 512.400 ;
        RECT 287.600 517.600 288.400 518.400 ;
        RECT 255.600 511.200 256.400 512.000 ;
        RECT 287.600 511.600 288.400 512.400 ;
        RECT 601.200 511.200 602.000 512.000 ;
        RECT 159.600 483.600 160.400 484.400 ;
        RECT 204.400 483.600 205.200 484.400 ;
        RECT 239.600 483.600 240.400 484.400 ;
        RECT 604.400 490.000 605.200 490.800 ;
        RECT 604.400 485.400 605.200 486.200 ;
        RECT 150.200 480.600 151.000 481.400 ;
        RECT 151.600 480.600 152.400 481.400 ;
        RECT 153.000 480.600 153.800 481.400 ;
        RECT 457.400 480.600 458.200 481.400 ;
        RECT 458.800 480.600 459.600 481.400 ;
        RECT 460.200 480.600 461.000 481.400 ;
        RECT 609.200 477.600 610.000 478.400 ;
        RECT 609.200 471.600 610.000 472.400 ;
        RECT 266.800 443.600 267.600 444.400 ;
        RECT 326.000 443.600 326.800 444.400 ;
        RECT 601.200 450.000 602.000 450.800 ;
        RECT 569.200 443.600 570.000 444.400 ;
        RECT 601.200 445.400 602.000 446.200 ;
        RECT 150.200 440.600 151.000 441.400 ;
        RECT 151.600 440.600 152.400 441.400 ;
        RECT 153.000 440.600 153.800 441.400 ;
        RECT 457.400 440.600 458.200 441.400 ;
        RECT 458.800 440.600 459.600 441.400 ;
        RECT 460.200 440.600 461.000 441.400 ;
        RECT 316.400 437.600 317.200 438.400 ;
        RECT 316.400 431.600 317.200 432.400 ;
        RECT 540.400 437.600 541.200 438.400 ;
        RECT 502.000 431.200 502.800 432.000 ;
        RECT 540.400 431.600 541.200 432.400 ;
        RECT 594.800 437.600 595.600 438.400 ;
        RECT 594.800 431.600 595.600 432.400 ;
        RECT 4.400 403.600 5.200 404.400 ;
        RECT 188.400 405.400 189.200 406.200 ;
        RECT 306.800 403.600 307.600 404.400 ;
        RECT 582.000 405.400 582.800 406.200 ;
        RECT 150.200 400.600 151.000 401.400 ;
        RECT 151.600 400.600 152.400 401.400 ;
        RECT 153.000 400.600 153.800 401.400 ;
        RECT 457.400 400.600 458.200 401.400 ;
        RECT 458.800 400.600 459.600 401.400 ;
        RECT 460.200 400.600 461.000 401.400 ;
        RECT 4.400 397.600 5.200 398.400 ;
        RECT 4.400 391.600 5.200 392.400 ;
        RECT 196.400 397.600 197.200 398.400 ;
        RECT 196.400 391.600 197.200 392.400 ;
        RECT 220.400 391.200 221.200 392.000 ;
        RECT 268.400 397.600 269.200 398.400 ;
        RECT 308.400 397.600 309.200 398.400 ;
        RECT 370.800 397.600 371.600 398.400 ;
        RECT 268.400 391.600 269.200 392.400 ;
        RECT 308.400 391.600 309.200 392.400 ;
        RECT 370.800 391.600 371.600 392.400 ;
        RECT 438.000 397.600 438.800 398.400 ;
        RECT 438.000 391.600 438.800 392.400 ;
        RECT 462.000 397.600 462.800 398.400 ;
        RECT 462.000 391.600 462.800 392.400 ;
        RECT 521.200 397.600 522.000 398.400 ;
        RECT 521.200 391.600 522.000 392.400 ;
        RECT 577.200 397.600 578.000 398.400 ;
        RECT 577.200 391.600 578.000 392.400 ;
        RECT 529.200 371.600 530.000 372.400 ;
        RECT 180.400 365.400 181.200 366.200 ;
        RECT 263.600 363.600 264.400 364.400 ;
        RECT 406.000 370.000 406.800 370.800 ;
        RECT 350.000 365.400 350.800 366.200 ;
        RECT 406.000 365.400 406.800 366.200 ;
        RECT 474.800 370.000 475.600 370.800 ;
        RECT 474.800 363.600 475.600 364.400 ;
        RECT 529.200 365.400 530.000 366.200 ;
        RECT 602.800 363.600 603.600 364.400 ;
        RECT 150.200 360.600 151.000 361.400 ;
        RECT 151.600 360.600 152.400 361.400 ;
        RECT 153.000 360.600 153.800 361.400 ;
        RECT 457.400 360.600 458.200 361.400 ;
        RECT 458.800 360.600 459.600 361.400 ;
        RECT 460.200 360.600 461.000 361.400 ;
        RECT 14.000 357.600 14.800 358.400 ;
        RECT 14.000 351.600 14.800 352.400 ;
        RECT 182.000 357.600 182.800 358.400 ;
        RECT 182.000 351.600 182.800 352.400 ;
        RECT 238.000 357.600 238.800 358.400 ;
        RECT 238.000 351.600 238.800 352.400 ;
        RECT 292.400 351.200 293.200 352.000 ;
        RECT 342.000 357.600 342.800 358.400 ;
        RECT 342.000 351.600 342.800 352.400 ;
        RECT 444.400 357.600 445.200 358.400 ;
        RECT 444.400 351.600 445.200 352.400 ;
        RECT 486.000 351.200 486.800 352.000 ;
        RECT 500.400 351.200 501.200 352.000 ;
        RECT 569.200 357.600 570.000 358.400 ;
        RECT 569.200 351.600 570.000 352.400 ;
        RECT 4.400 323.600 5.200 324.400 ;
        RECT 89.200 323.600 90.000 324.400 ;
        RECT 183.600 323.600 184.400 324.400 ;
        RECT 201.200 323.600 202.000 324.400 ;
        RECT 247.600 325.400 248.400 326.200 ;
        RECT 366.000 323.600 366.800 324.400 ;
        RECT 426.800 323.600 427.600 324.400 ;
        RECT 532.400 330.000 533.200 330.800 ;
        RECT 532.400 325.400 533.200 326.200 ;
        RECT 543.600 323.600 544.400 324.400 ;
        RECT 150.200 320.600 151.000 321.400 ;
        RECT 151.600 320.600 152.400 321.400 ;
        RECT 153.000 320.600 153.800 321.400 ;
        RECT 457.400 320.600 458.200 321.400 ;
        RECT 458.800 320.600 459.600 321.400 ;
        RECT 460.200 320.600 461.000 321.400 ;
        RECT 18.800 317.600 19.600 318.400 ;
        RECT 81.200 317.600 82.000 318.400 ;
        RECT 18.800 311.600 19.600 312.400 ;
        RECT 81.200 311.600 82.000 312.400 ;
        RECT 138.800 317.600 139.600 318.400 ;
        RECT 138.800 311.600 139.600 312.400 ;
        RECT 186.800 311.200 187.600 312.000 ;
        RECT 207.600 311.200 208.400 312.000 ;
        RECT 324.400 311.200 325.200 312.000 ;
        RECT 428.400 317.600 429.200 318.400 ;
        RECT 428.400 311.600 429.200 312.400 ;
        RECT 553.200 317.600 554.000 318.400 ;
        RECT 553.200 311.600 554.000 312.400 ;
        RECT 18.800 283.600 19.600 284.400 ;
        RECT 65.200 283.600 66.000 284.400 ;
        RECT 148.400 290.000 149.200 290.800 ;
        RECT 148.400 283.600 149.200 284.400 ;
        RECT 177.200 283.600 178.000 284.400 ;
        RECT 222.000 283.600 222.800 284.400 ;
        RECT 270.000 283.600 270.800 284.400 ;
        RECT 428.400 283.600 429.200 284.400 ;
        RECT 564.400 290.000 565.200 290.800 ;
        RECT 564.400 285.400 565.200 286.200 ;
        RECT 580.400 283.600 581.200 284.400 ;
        RECT 150.200 280.600 151.000 281.400 ;
        RECT 151.600 280.600 152.400 281.400 ;
        RECT 153.000 280.600 153.800 281.400 ;
        RECT 457.400 280.600 458.200 281.400 ;
        RECT 458.800 280.600 459.600 281.400 ;
        RECT 460.200 280.600 461.000 281.400 ;
        RECT 4.400 277.600 5.200 278.400 ;
        RECT 66.800 277.600 67.600 278.400 ;
        RECT 4.400 271.600 5.200 272.400 ;
        RECT 66.800 271.600 67.600 272.400 ;
        RECT 113.200 277.600 114.000 278.400 ;
        RECT 113.200 271.600 114.000 272.400 ;
        RECT 178.800 277.600 179.600 278.400 ;
        RECT 178.800 271.600 179.600 272.400 ;
        RECT 234.800 277.600 235.600 278.400 ;
        RECT 234.800 271.600 235.600 272.400 ;
        RECT 316.400 271.200 317.200 272.000 ;
        RECT 604.400 271.200 605.200 272.000 ;
        RECT 4.400 243.600 5.200 244.400 ;
        RECT 46.000 245.400 46.800 246.200 ;
        RECT 121.200 250.000 122.000 250.800 ;
        RECT 121.200 245.400 122.000 246.200 ;
        RECT 170.800 250.000 171.600 250.800 ;
        RECT 170.800 245.400 171.600 246.200 ;
        RECT 201.200 243.600 202.000 244.400 ;
        RECT 279.600 243.600 280.400 244.400 ;
        RECT 358.000 245.400 358.800 246.200 ;
        RECT 596.400 250.000 597.200 250.800 ;
        RECT 596.400 245.400 597.200 246.200 ;
        RECT 150.200 240.600 151.000 241.400 ;
        RECT 151.600 240.600 152.400 241.400 ;
        RECT 153.000 240.600 153.800 241.400 ;
        RECT 457.400 240.600 458.200 241.400 ;
        RECT 458.800 240.600 459.600 241.400 ;
        RECT 460.200 240.600 461.000 241.400 ;
        RECT 47.600 237.600 48.400 238.400 ;
        RECT 47.600 231.600 48.400 232.400 ;
        RECT 191.600 237.600 192.400 238.400 ;
        RECT 156.400 231.200 157.200 232.000 ;
        RECT 191.600 231.600 192.400 232.400 ;
        RECT 234.800 237.600 235.600 238.400 ;
        RECT 234.800 231.600 235.600 232.400 ;
        RECT 374.000 231.200 374.800 232.000 ;
        RECT 598.000 237.600 598.800 238.400 ;
        RECT 598.000 231.600 598.800 232.400 ;
        RECT 207.600 203.600 208.400 204.400 ;
        RECT 215.600 203.600 216.400 204.400 ;
        RECT 257.200 203.600 258.000 204.400 ;
        RECT 338.800 203.600 339.600 204.400 ;
        RECT 377.200 210.000 378.000 210.800 ;
        RECT 377.200 203.600 378.000 204.400 ;
        RECT 452.400 210.000 453.200 210.800 ;
        RECT 452.400 205.400 453.200 206.200 ;
        RECT 494.000 205.400 494.800 206.200 ;
        RECT 564.400 210.000 565.200 210.800 ;
        RECT 564.400 205.400 565.200 206.200 ;
        RECT 150.200 200.600 151.000 201.400 ;
        RECT 151.600 200.600 152.400 201.400 ;
        RECT 153.000 200.600 153.800 201.400 ;
        RECT 457.400 200.600 458.200 201.400 ;
        RECT 458.800 200.600 459.600 201.400 ;
        RECT 460.200 200.600 461.000 201.400 ;
        RECT 4.400 197.600 5.200 198.400 ;
        RECT 4.400 191.600 5.200 192.400 ;
        RECT 202.800 197.600 203.600 198.400 ;
        RECT 202.800 191.600 203.600 192.400 ;
        RECT 258.800 197.600 259.600 198.400 ;
        RECT 258.800 191.600 259.600 192.400 ;
        RECT 350.000 191.200 350.800 192.000 ;
        RECT 394.800 197.600 395.600 198.400 ;
        RECT 438.000 197.600 438.800 198.400 ;
        RECT 394.800 191.600 395.600 192.400 ;
        RECT 406.000 191.200 406.800 192.000 ;
        RECT 438.000 191.600 438.800 192.400 ;
        RECT 558.000 197.600 558.800 198.400 ;
        RECT 558.000 191.600 558.800 192.400 ;
        RECT 569.200 191.200 570.000 192.000 ;
        RECT 180.400 163.600 181.200 164.400 ;
        RECT 234.800 170.000 235.600 170.800 ;
        RECT 234.800 165.400 235.600 166.200 ;
        RECT 246.000 163.600 246.800 164.400 ;
        RECT 308.400 165.400 309.200 166.200 ;
        RECT 591.600 170.000 592.400 170.800 ;
        RECT 591.600 163.600 592.400 164.400 ;
        RECT 150.200 160.600 151.000 161.400 ;
        RECT 151.600 160.600 152.400 161.400 ;
        RECT 153.000 160.600 153.800 161.400 ;
        RECT 457.400 160.600 458.200 161.400 ;
        RECT 458.800 160.600 459.600 161.400 ;
        RECT 460.200 160.600 461.000 161.400 ;
        RECT 167.600 151.200 168.400 152.000 ;
        RECT 268.400 157.600 269.200 158.400 ;
        RECT 231.600 151.200 232.400 152.000 ;
        RECT 268.400 151.600 269.200 152.400 ;
        RECT 326.000 151.200 326.800 152.000 ;
        RECT 598.000 157.600 598.800 158.400 ;
        RECT 598.000 151.600 598.800 152.400 ;
        RECT 31.600 123.600 32.400 124.400 ;
        RECT 190.000 130.000 190.800 130.800 ;
        RECT 190.000 125.400 190.800 126.200 ;
        RECT 239.600 123.600 240.400 124.400 ;
        RECT 294.000 130.000 294.800 130.800 ;
        RECT 294.000 125.400 294.800 126.200 ;
        RECT 324.400 123.600 325.200 124.400 ;
        RECT 385.200 123.600 386.000 124.400 ;
        RECT 150.200 120.600 151.000 121.400 ;
        RECT 151.600 120.600 152.400 121.400 ;
        RECT 153.000 120.600 153.800 121.400 ;
        RECT 457.400 120.600 458.200 121.400 ;
        RECT 458.800 120.600 459.600 121.400 ;
        RECT 460.200 120.600 461.000 121.400 ;
        RECT 340.400 111.200 341.200 112.000 ;
        RECT 374.000 117.600 374.800 118.400 ;
        RECT 374.000 111.600 374.800 112.400 ;
        RECT 596.400 111.200 597.200 112.000 ;
        RECT 268.400 109.600 269.200 110.400 ;
        RECT 340.400 91.600 341.200 92.400 ;
        RECT 183.600 85.400 184.400 86.200 ;
        RECT 276.400 90.000 277.200 90.800 ;
        RECT 276.400 83.600 277.200 84.400 ;
        RECT 287.600 83.600 288.400 84.400 ;
        RECT 340.400 85.400 341.200 86.200 ;
        RECT 372.400 85.400 373.200 86.200 ;
        RECT 582.000 85.400 582.800 86.200 ;
        RECT 150.200 80.600 151.000 81.400 ;
        RECT 151.600 80.600 152.400 81.400 ;
        RECT 153.000 80.600 153.800 81.400 ;
        RECT 457.400 80.600 458.200 81.400 ;
        RECT 458.800 80.600 459.600 81.400 ;
        RECT 460.200 80.600 461.000 81.400 ;
        RECT 207.600 77.600 208.400 78.400 ;
        RECT 207.600 71.600 208.400 72.400 ;
        RECT 332.400 77.600 333.200 78.400 ;
        RECT 284.400 71.200 285.200 72.000 ;
        RECT 332.400 71.600 333.200 72.400 ;
        RECT 4.400 43.600 5.200 44.400 ;
        RECT 183.600 43.600 184.400 44.400 ;
        RECT 246.000 43.600 246.800 44.400 ;
        RECT 302.000 45.400 302.800 46.200 ;
        RECT 378.800 43.600 379.600 44.400 ;
        RECT 604.400 50.000 605.200 50.800 ;
        RECT 604.400 45.400 605.200 46.200 ;
        RECT 150.200 40.600 151.000 41.400 ;
        RECT 151.600 40.600 152.400 41.400 ;
        RECT 153.000 40.600 153.800 41.400 ;
        RECT 457.400 40.600 458.200 41.400 ;
        RECT 458.800 40.600 459.600 41.400 ;
        RECT 460.200 40.600 461.000 41.400 ;
        RECT 9.200 37.600 10.000 38.400 ;
        RECT 9.200 31.600 10.000 32.400 ;
        RECT 206.000 31.200 206.800 32.000 ;
        RECT 239.600 31.200 240.400 32.000 ;
        RECT 278.000 31.200 278.800 32.000 ;
        RECT 388.400 37.600 389.200 38.400 ;
        RECT 388.400 31.600 389.200 32.400 ;
        RECT 596.400 31.200 597.200 32.000 ;
        RECT 4.400 3.600 5.200 4.400 ;
        RECT 175.600 3.600 176.400 4.400 ;
        RECT 186.800 3.600 187.600 4.400 ;
        RECT 223.600 3.600 224.400 4.400 ;
        RECT 276.400 5.400 277.200 6.200 ;
        RECT 321.200 3.600 322.000 4.400 ;
        RECT 367.600 3.600 368.400 4.400 ;
        RECT 599.600 10.000 600.400 10.800 ;
        RECT 599.600 3.600 600.400 4.400 ;
        RECT 150.200 0.600 151.000 1.400 ;
        RECT 151.600 0.600 152.400 1.400 ;
        RECT 153.000 0.600 153.800 1.400 ;
        RECT 457.400 0.600 458.200 1.400 ;
        RECT 458.800 0.600 459.600 1.400 ;
        RECT 460.200 0.600 461.000 1.400 ;
      LAYER metal2 ;
        RECT 149.600 560.600 154.400 561.400 ;
        RECT 456.800 560.600 461.600 561.400 ;
        RECT 7.600 557.600 8.400 558.400 ;
        RECT 95.600 557.600 96.400 558.400 ;
        RECT 146.800 557.600 147.600 558.400 ;
        RECT 206.000 557.600 206.800 558.400 ;
        RECT 260.400 557.600 261.200 558.400 ;
        RECT 332.400 557.600 333.200 558.400 ;
        RECT 7.700 552.400 8.300 557.600 ;
        RECT 95.700 552.400 96.300 557.600 ;
        RECT 146.900 552.400 147.500 557.600 ;
        RECT 206.100 552.400 206.700 557.600 ;
        RECT 260.500 552.400 261.100 557.600 ;
        RECT 332.500 552.400 333.100 557.600 ;
        RECT 396.400 555.800 397.200 556.600 ;
        RECT 585.200 555.800 586.000 556.600 ;
        RECT 7.600 551.600 8.400 552.400 ;
        RECT 95.600 551.600 96.400 552.400 ;
        RECT 146.800 551.600 147.600 552.400 ;
        RECT 206.000 551.600 206.800 552.400 ;
        RECT 260.400 551.600 261.200 552.400 ;
        RECT 332.400 551.600 333.200 552.400 ;
        RECT 396.500 552.000 397.100 555.800 ;
        RECT 585.300 552.000 585.900 555.800 ;
        RECT 396.400 551.200 397.200 552.000 ;
        RECT 585.200 551.200 586.000 552.000 ;
        RECT 7.600 530.000 8.400 530.800 ;
        RECT 7.700 524.400 8.300 530.000 ;
        RECT 94.000 529.600 94.800 530.400 ;
        RECT 170.800 529.600 171.600 530.400 ;
        RECT 182.000 530.000 182.800 530.800 ;
        RECT 94.100 524.400 94.700 529.600 ;
        RECT 170.900 524.400 171.500 529.600 ;
        RECT 182.100 524.400 182.700 530.000 ;
        RECT 255.600 529.600 256.400 530.400 ;
        RECT 263.600 529.600 264.400 530.400 ;
        RECT 342.000 530.000 342.800 530.800 ;
        RECT 409.200 530.000 410.000 530.800 ;
        RECT 255.700 524.400 256.300 529.600 ;
        RECT 263.700 524.400 264.300 529.600 ;
        RECT 342.100 526.200 342.700 530.000 ;
        RECT 342.000 525.400 342.800 526.200 ;
        RECT 409.300 524.400 409.900 530.000 ;
        RECT 574.000 529.600 574.800 530.400 ;
        RECT 574.100 524.400 574.700 529.600 ;
        RECT 7.600 523.600 8.400 524.400 ;
        RECT 94.000 523.600 94.800 524.400 ;
        RECT 170.800 523.600 171.600 524.400 ;
        RECT 182.000 523.600 182.800 524.400 ;
        RECT 255.600 523.600 256.400 524.400 ;
        RECT 263.600 523.600 264.400 524.400 ;
        RECT 409.200 523.600 410.000 524.400 ;
        RECT 574.000 523.600 574.800 524.400 ;
        RECT 149.600 520.600 154.400 521.400 ;
        RECT 456.800 520.600 461.600 521.400 ;
        RECT 202.800 517.600 203.600 518.400 ;
        RECT 287.600 517.600 288.400 518.400 ;
        RECT 202.900 512.400 203.500 517.600 ;
        RECT 255.600 515.800 256.400 516.600 ;
        RECT 202.800 511.600 203.600 512.400 ;
        RECT 255.700 512.000 256.300 515.800 ;
        RECT 287.700 512.400 288.300 517.600 ;
        RECT 601.200 515.800 602.000 516.600 ;
        RECT 255.600 511.200 256.400 512.000 ;
        RECT 287.600 511.600 288.400 512.400 ;
        RECT 601.300 512.000 601.900 515.800 ;
        RECT 601.200 511.200 602.000 512.000 ;
        RECT 159.600 489.600 160.400 490.400 ;
        RECT 204.400 489.600 205.200 490.400 ;
        RECT 239.600 489.600 240.400 490.400 ;
        RECT 604.400 490.000 605.200 490.800 ;
        RECT 159.700 484.400 160.300 489.600 ;
        RECT 204.500 484.400 205.100 489.600 ;
        RECT 239.700 484.400 240.300 489.600 ;
        RECT 604.500 486.200 605.100 490.000 ;
        RECT 604.400 485.400 605.200 486.200 ;
        RECT 159.600 483.600 160.400 484.400 ;
        RECT 204.400 483.600 205.200 484.400 ;
        RECT 239.600 483.600 240.400 484.400 ;
        RECT 149.600 480.600 154.400 481.400 ;
        RECT 456.800 480.600 461.600 481.400 ;
        RECT 609.200 477.600 610.000 478.400 ;
        RECT 266.800 475.600 267.600 476.400 ;
        RECT 266.900 470.400 267.500 475.600 ;
        RECT 609.300 472.400 609.900 477.600 ;
        RECT 609.200 471.600 610.000 472.400 ;
        RECT 266.800 469.600 267.600 470.400 ;
        RECT 266.800 449.600 267.600 450.400 ;
        RECT 326.000 449.600 326.800 450.400 ;
        RECT 569.200 449.600 570.000 450.400 ;
        RECT 601.200 450.000 602.000 450.800 ;
        RECT 266.900 444.400 267.500 449.600 ;
        RECT 326.100 444.400 326.700 449.600 ;
        RECT 569.300 444.400 569.900 449.600 ;
        RECT 601.300 446.200 601.900 450.000 ;
        RECT 601.200 445.400 602.000 446.200 ;
        RECT 266.800 443.600 267.600 444.400 ;
        RECT 326.000 443.600 326.800 444.400 ;
        RECT 569.200 443.600 570.000 444.400 ;
        RECT 149.600 440.600 154.400 441.400 ;
        RECT 456.800 440.600 461.600 441.400 ;
        RECT 316.400 437.600 317.200 438.400 ;
        RECT 540.400 437.600 541.200 438.400 ;
        RECT 594.800 437.600 595.600 438.400 ;
        RECT 316.500 432.400 317.100 437.600 ;
        RECT 502.000 435.800 502.800 436.600 ;
        RECT 316.400 431.600 317.200 432.400 ;
        RECT 502.100 432.000 502.700 435.800 ;
        RECT 540.500 432.400 541.100 437.600 ;
        RECT 594.900 432.400 595.500 437.600 ;
        RECT 502.000 431.200 502.800 432.000 ;
        RECT 540.400 431.600 541.200 432.400 ;
        RECT 594.800 431.600 595.600 432.400 ;
        RECT 4.400 409.600 5.200 410.400 ;
        RECT 188.400 410.000 189.200 410.800 ;
        RECT 306.800 410.000 307.600 410.800 ;
        RECT 582.000 410.000 582.800 410.800 ;
        RECT 4.500 404.400 5.100 409.600 ;
        RECT 188.500 406.200 189.100 410.000 ;
        RECT 188.400 405.400 189.200 406.200 ;
        RECT 306.900 404.400 307.500 410.000 ;
        RECT 582.100 406.200 582.700 410.000 ;
        RECT 582.000 405.400 582.800 406.200 ;
        RECT 4.400 403.600 5.200 404.400 ;
        RECT 306.800 403.600 307.600 404.400 ;
        RECT 149.600 400.600 154.400 401.400 ;
        RECT 456.800 400.600 461.600 401.400 ;
        RECT 4.400 397.600 5.200 398.400 ;
        RECT 196.400 397.600 197.200 398.400 ;
        RECT 268.400 397.600 269.200 398.400 ;
        RECT 308.400 397.600 309.200 398.400 ;
        RECT 370.800 397.600 371.600 398.400 ;
        RECT 438.000 397.600 438.800 398.400 ;
        RECT 462.000 397.600 462.800 398.400 ;
        RECT 521.200 397.600 522.000 398.400 ;
        RECT 577.200 397.600 578.000 398.400 ;
        RECT 4.500 392.400 5.100 397.600 ;
        RECT 196.500 392.400 197.100 397.600 ;
        RECT 220.400 395.800 221.200 396.600 ;
        RECT 4.400 391.600 5.200 392.400 ;
        RECT 196.400 391.600 197.200 392.400 ;
        RECT 220.500 392.000 221.100 395.800 ;
        RECT 268.500 392.400 269.100 397.600 ;
        RECT 308.500 392.400 309.100 397.600 ;
        RECT 370.900 392.400 371.500 397.600 ;
        RECT 438.100 392.400 438.700 397.600 ;
        RECT 462.100 392.400 462.700 397.600 ;
        RECT 521.300 392.400 521.900 397.600 ;
        RECT 577.300 392.400 577.900 397.600 ;
        RECT 220.400 391.200 221.200 392.000 ;
        RECT 268.400 391.600 269.200 392.400 ;
        RECT 308.400 391.600 309.200 392.400 ;
        RECT 370.800 391.600 371.600 392.400 ;
        RECT 438.000 391.600 438.800 392.400 ;
        RECT 462.000 391.600 462.800 392.400 ;
        RECT 521.200 391.600 522.000 392.400 ;
        RECT 577.200 391.600 578.000 392.400 ;
        RECT 529.200 371.600 530.000 372.400 ;
        RECT 180.400 370.000 181.200 370.800 ;
        RECT 180.500 366.200 181.100 370.000 ;
        RECT 263.600 369.600 264.400 370.400 ;
        RECT 350.000 370.000 350.800 370.800 ;
        RECT 406.000 370.000 406.800 370.800 ;
        RECT 474.800 370.000 475.600 370.800 ;
        RECT 180.400 365.400 181.200 366.200 ;
        RECT 263.700 364.400 264.300 369.600 ;
        RECT 350.100 366.200 350.700 370.000 ;
        RECT 406.100 366.200 406.700 370.000 ;
        RECT 350.000 365.400 350.800 366.200 ;
        RECT 406.000 365.400 406.800 366.200 ;
        RECT 474.900 364.400 475.500 370.000 ;
        RECT 529.300 366.200 529.900 371.600 ;
        RECT 602.800 369.600 603.600 370.400 ;
        RECT 529.200 365.400 530.000 366.200 ;
        RECT 602.900 364.400 603.500 369.600 ;
        RECT 263.600 363.600 264.400 364.400 ;
        RECT 474.800 363.600 475.600 364.400 ;
        RECT 602.800 363.600 603.600 364.400 ;
        RECT 149.600 360.600 154.400 361.400 ;
        RECT 456.800 360.600 461.600 361.400 ;
        RECT 14.000 357.600 14.800 358.400 ;
        RECT 182.000 357.600 182.800 358.400 ;
        RECT 238.000 357.600 238.800 358.400 ;
        RECT 342.000 357.600 342.800 358.400 ;
        RECT 444.400 357.600 445.200 358.400 ;
        RECT 569.200 357.600 570.000 358.400 ;
        RECT 14.100 352.400 14.700 357.600 ;
        RECT 182.100 352.400 182.700 357.600 ;
        RECT 238.100 352.400 238.700 357.600 ;
        RECT 292.400 355.800 293.200 356.600 ;
        RECT 14.000 351.600 14.800 352.400 ;
        RECT 182.000 351.600 182.800 352.400 ;
        RECT 238.000 351.600 238.800 352.400 ;
        RECT 292.500 352.000 293.100 355.800 ;
        RECT 342.100 352.400 342.700 357.600 ;
        RECT 444.500 352.400 445.100 357.600 ;
        RECT 486.000 355.800 486.800 356.600 ;
        RECT 500.400 355.800 501.200 356.600 ;
        RECT 292.400 351.200 293.200 352.000 ;
        RECT 342.000 351.600 342.800 352.400 ;
        RECT 444.400 351.600 445.200 352.400 ;
        RECT 486.100 352.000 486.700 355.800 ;
        RECT 500.500 352.000 501.100 355.800 ;
        RECT 569.300 352.400 569.900 357.600 ;
        RECT 486.000 351.200 486.800 352.000 ;
        RECT 500.400 351.200 501.200 352.000 ;
        RECT 569.200 351.600 570.000 352.400 ;
        RECT 4.400 329.600 5.200 330.400 ;
        RECT 89.200 329.600 90.000 330.400 ;
        RECT 183.600 329.600 184.400 330.400 ;
        RECT 201.200 330.000 202.000 330.800 ;
        RECT 247.600 330.000 248.400 330.800 ;
        RECT 4.500 324.400 5.100 329.600 ;
        RECT 89.300 324.400 89.900 329.600 ;
        RECT 183.700 324.400 184.300 329.600 ;
        RECT 201.300 324.400 201.900 330.000 ;
        RECT 247.700 326.200 248.300 330.000 ;
        RECT 366.000 329.600 366.800 330.400 ;
        RECT 426.800 329.600 427.600 330.400 ;
        RECT 532.400 330.000 533.200 330.800 ;
        RECT 247.600 325.400 248.400 326.200 ;
        RECT 366.100 324.400 366.700 329.600 ;
        RECT 426.900 324.400 427.500 329.600 ;
        RECT 532.500 326.200 533.100 330.000 ;
        RECT 543.600 329.600 544.400 330.400 ;
        RECT 532.400 325.400 533.200 326.200 ;
        RECT 543.700 324.400 544.300 329.600 ;
        RECT 4.400 323.600 5.200 324.400 ;
        RECT 89.200 323.600 90.000 324.400 ;
        RECT 183.600 323.600 184.400 324.400 ;
        RECT 201.200 323.600 202.000 324.400 ;
        RECT 366.000 323.600 366.800 324.400 ;
        RECT 426.800 323.600 427.600 324.400 ;
        RECT 543.600 323.600 544.400 324.400 ;
        RECT 149.600 320.600 154.400 321.400 ;
        RECT 456.800 320.600 461.600 321.400 ;
        RECT 18.800 317.600 19.600 318.400 ;
        RECT 81.200 317.600 82.000 318.400 ;
        RECT 138.800 317.600 139.600 318.400 ;
        RECT 428.400 317.600 429.200 318.400 ;
        RECT 553.200 317.600 554.000 318.400 ;
        RECT 18.900 312.400 19.500 317.600 ;
        RECT 81.300 312.400 81.900 317.600 ;
        RECT 138.900 312.400 139.500 317.600 ;
        RECT 186.800 315.800 187.600 316.600 ;
        RECT 207.600 315.800 208.400 316.600 ;
        RECT 324.400 315.800 325.200 316.600 ;
        RECT 18.800 311.600 19.600 312.400 ;
        RECT 81.200 311.600 82.000 312.400 ;
        RECT 138.800 311.600 139.600 312.400 ;
        RECT 186.900 312.000 187.500 315.800 ;
        RECT 207.700 312.000 208.300 315.800 ;
        RECT 324.500 312.000 325.100 315.800 ;
        RECT 428.500 312.400 429.100 317.600 ;
        RECT 553.300 312.400 553.900 317.600 ;
        RECT 186.800 311.200 187.600 312.000 ;
        RECT 207.600 311.200 208.400 312.000 ;
        RECT 324.400 311.200 325.200 312.000 ;
        RECT 428.400 311.600 429.200 312.400 ;
        RECT 553.200 311.600 554.000 312.400 ;
        RECT 18.800 289.600 19.600 290.400 ;
        RECT 65.200 289.600 66.000 290.400 ;
        RECT 148.400 290.000 149.200 290.800 ;
        RECT 177.200 290.000 178.000 290.800 ;
        RECT 18.900 284.400 19.500 289.600 ;
        RECT 65.300 284.400 65.900 289.600 ;
        RECT 148.500 284.400 149.100 290.000 ;
        RECT 177.300 284.400 177.900 290.000 ;
        RECT 222.000 289.600 222.800 290.400 ;
        RECT 270.000 289.600 270.800 290.400 ;
        RECT 428.400 289.600 429.200 290.400 ;
        RECT 564.400 290.000 565.200 290.800 ;
        RECT 222.100 284.400 222.700 289.600 ;
        RECT 270.100 284.400 270.700 289.600 ;
        RECT 428.500 284.400 429.100 289.600 ;
        RECT 564.500 286.200 565.100 290.000 ;
        RECT 580.400 289.600 581.200 290.400 ;
        RECT 564.400 285.400 565.200 286.200 ;
        RECT 580.500 284.400 581.100 289.600 ;
        RECT 18.800 283.600 19.600 284.400 ;
        RECT 65.200 283.600 66.000 284.400 ;
        RECT 148.400 283.600 149.200 284.400 ;
        RECT 177.200 283.600 178.000 284.400 ;
        RECT 222.000 283.600 222.800 284.400 ;
        RECT 270.000 283.600 270.800 284.400 ;
        RECT 428.400 283.600 429.200 284.400 ;
        RECT 580.400 283.600 581.200 284.400 ;
        RECT 149.600 280.600 154.400 281.400 ;
        RECT 456.800 280.600 461.600 281.400 ;
        RECT 4.400 277.600 5.200 278.400 ;
        RECT 66.800 277.600 67.600 278.400 ;
        RECT 113.200 277.600 114.000 278.400 ;
        RECT 178.800 277.600 179.600 278.400 ;
        RECT 234.800 277.600 235.600 278.400 ;
        RECT 4.500 272.400 5.100 277.600 ;
        RECT 66.900 272.400 67.500 277.600 ;
        RECT 113.300 272.400 113.900 277.600 ;
        RECT 178.900 272.400 179.500 277.600 ;
        RECT 234.900 272.400 235.500 277.600 ;
        RECT 316.400 275.800 317.200 276.600 ;
        RECT 604.400 275.800 605.200 276.600 ;
        RECT 4.400 271.600 5.200 272.400 ;
        RECT 66.800 271.600 67.600 272.400 ;
        RECT 113.200 271.600 114.000 272.400 ;
        RECT 178.800 271.600 179.600 272.400 ;
        RECT 234.800 271.600 235.600 272.400 ;
        RECT 316.500 272.000 317.100 275.800 ;
        RECT 604.500 272.000 605.100 275.800 ;
        RECT 316.400 271.200 317.200 272.000 ;
        RECT 604.400 271.200 605.200 272.000 ;
        RECT 4.400 249.600 5.200 250.400 ;
        RECT 46.000 250.000 46.800 250.800 ;
        RECT 121.200 250.000 122.000 250.800 ;
        RECT 170.800 250.000 171.600 250.800 ;
        RECT 201.200 250.000 202.000 250.800 ;
        RECT 4.500 244.400 5.100 249.600 ;
        RECT 46.100 246.200 46.700 250.000 ;
        RECT 121.300 246.200 121.900 250.000 ;
        RECT 170.900 246.200 171.500 250.000 ;
        RECT 46.000 245.400 46.800 246.200 ;
        RECT 121.200 245.400 122.000 246.200 ;
        RECT 170.800 245.400 171.600 246.200 ;
        RECT 201.300 244.400 201.900 250.000 ;
        RECT 279.600 249.600 280.400 250.400 ;
        RECT 358.000 250.000 358.800 250.800 ;
        RECT 596.400 250.000 597.200 250.800 ;
        RECT 279.700 244.400 280.300 249.600 ;
        RECT 358.100 246.200 358.700 250.000 ;
        RECT 596.500 246.200 597.100 250.000 ;
        RECT 358.000 245.400 358.800 246.200 ;
        RECT 596.400 245.400 597.200 246.200 ;
        RECT 4.400 243.600 5.200 244.400 ;
        RECT 201.200 243.600 202.000 244.400 ;
        RECT 279.600 243.600 280.400 244.400 ;
        RECT 149.600 240.600 154.400 241.400 ;
        RECT 456.800 240.600 461.600 241.400 ;
        RECT 47.600 237.600 48.400 238.400 ;
        RECT 191.600 237.600 192.400 238.400 ;
        RECT 234.800 237.600 235.600 238.400 ;
        RECT 598.000 237.600 598.800 238.400 ;
        RECT 47.700 232.400 48.300 237.600 ;
        RECT 156.400 235.800 157.200 236.600 ;
        RECT 47.600 231.600 48.400 232.400 ;
        RECT 156.500 232.000 157.100 235.800 ;
        RECT 191.700 232.400 192.300 237.600 ;
        RECT 234.900 232.400 235.500 237.600 ;
        RECT 374.000 235.800 374.800 236.600 ;
        RECT 156.400 231.200 157.200 232.000 ;
        RECT 191.600 231.600 192.400 232.400 ;
        RECT 234.800 231.600 235.600 232.400 ;
        RECT 374.100 232.000 374.700 235.800 ;
        RECT 598.100 232.400 598.700 237.600 ;
        RECT 374.000 231.200 374.800 232.000 ;
        RECT 598.000 231.600 598.800 232.400 ;
        RECT 207.600 209.600 208.400 210.400 ;
        RECT 215.600 209.600 216.400 210.400 ;
        RECT 257.200 210.000 258.000 210.800 ;
        RECT 207.700 204.400 208.300 209.600 ;
        RECT 215.700 204.400 216.300 209.600 ;
        RECT 257.300 204.400 257.900 210.000 ;
        RECT 338.800 209.600 339.600 210.400 ;
        RECT 377.200 210.000 378.000 210.800 ;
        RECT 452.400 210.000 453.200 210.800 ;
        RECT 494.000 210.000 494.800 210.800 ;
        RECT 564.400 210.000 565.200 210.800 ;
        RECT 338.900 204.400 339.500 209.600 ;
        RECT 377.300 204.400 377.900 210.000 ;
        RECT 452.500 206.200 453.100 210.000 ;
        RECT 494.100 206.200 494.700 210.000 ;
        RECT 564.500 206.200 565.100 210.000 ;
        RECT 452.400 205.400 453.200 206.200 ;
        RECT 494.000 205.400 494.800 206.200 ;
        RECT 564.400 205.400 565.200 206.200 ;
        RECT 207.600 203.600 208.400 204.400 ;
        RECT 215.600 203.600 216.400 204.400 ;
        RECT 257.200 203.600 258.000 204.400 ;
        RECT 338.800 203.600 339.600 204.400 ;
        RECT 377.200 203.600 378.000 204.400 ;
        RECT 149.600 200.600 154.400 201.400 ;
        RECT 456.800 200.600 461.600 201.400 ;
        RECT 4.400 197.600 5.200 198.400 ;
        RECT 202.800 197.600 203.600 198.400 ;
        RECT 258.800 197.600 259.600 198.400 ;
        RECT 394.800 197.600 395.600 198.400 ;
        RECT 438.000 197.600 438.800 198.400 ;
        RECT 558.000 197.600 558.800 198.400 ;
        RECT 4.500 192.400 5.100 197.600 ;
        RECT 202.900 192.400 203.500 197.600 ;
        RECT 258.900 192.400 259.500 197.600 ;
        RECT 350.000 195.800 350.800 196.600 ;
        RECT 4.400 191.600 5.200 192.400 ;
        RECT 202.800 191.600 203.600 192.400 ;
        RECT 258.800 191.600 259.600 192.400 ;
        RECT 350.100 192.000 350.700 195.800 ;
        RECT 394.900 192.400 395.500 197.600 ;
        RECT 406.000 195.800 406.800 196.600 ;
        RECT 350.000 191.200 350.800 192.000 ;
        RECT 394.800 191.600 395.600 192.400 ;
        RECT 406.100 192.000 406.700 195.800 ;
        RECT 438.100 192.400 438.700 197.600 ;
        RECT 558.100 192.400 558.700 197.600 ;
        RECT 569.200 195.800 570.000 196.600 ;
        RECT 406.000 191.200 406.800 192.000 ;
        RECT 438.000 191.600 438.800 192.400 ;
        RECT 558.000 191.600 558.800 192.400 ;
        RECT 569.300 192.000 569.900 195.800 ;
        RECT 569.200 191.200 570.000 192.000 ;
        RECT 180.400 169.600 181.200 170.400 ;
        RECT 234.800 170.000 235.600 170.800 ;
        RECT 180.500 164.400 181.100 169.600 ;
        RECT 234.900 166.200 235.500 170.000 ;
        RECT 246.000 169.600 246.800 170.400 ;
        RECT 308.400 170.000 309.200 170.800 ;
        RECT 591.600 170.000 592.400 170.800 ;
        RECT 234.800 165.400 235.600 166.200 ;
        RECT 246.100 164.400 246.700 169.600 ;
        RECT 308.500 166.200 309.100 170.000 ;
        RECT 308.400 165.400 309.200 166.200 ;
        RECT 591.700 164.400 592.300 170.000 ;
        RECT 180.400 163.600 181.200 164.400 ;
        RECT 246.000 163.600 246.800 164.400 ;
        RECT 591.600 163.600 592.400 164.400 ;
        RECT 149.600 160.600 154.400 161.400 ;
        RECT 456.800 160.600 461.600 161.400 ;
        RECT 268.400 157.600 269.200 158.400 ;
        RECT 598.000 157.600 598.800 158.400 ;
        RECT 167.600 155.800 168.400 156.600 ;
        RECT 231.600 155.800 232.400 156.600 ;
        RECT 167.700 152.000 168.300 155.800 ;
        RECT 231.700 152.000 232.300 155.800 ;
        RECT 268.500 152.400 269.100 157.600 ;
        RECT 326.000 155.800 326.800 156.600 ;
        RECT 167.600 151.200 168.400 152.000 ;
        RECT 231.600 151.200 232.400 152.000 ;
        RECT 268.400 151.600 269.200 152.400 ;
        RECT 326.100 152.000 326.700 155.800 ;
        RECT 598.100 152.400 598.700 157.600 ;
        RECT 326.000 151.200 326.800 152.000 ;
        RECT 598.000 151.600 598.800 152.400 ;
        RECT 31.600 129.600 32.400 130.400 ;
        RECT 190.000 130.000 190.800 130.800 ;
        RECT 31.700 124.400 32.300 129.600 ;
        RECT 190.100 126.200 190.700 130.000 ;
        RECT 239.600 129.600 240.400 130.400 ;
        RECT 294.000 130.000 294.800 130.800 ;
        RECT 190.000 125.400 190.800 126.200 ;
        RECT 239.700 124.400 240.300 129.600 ;
        RECT 294.100 126.200 294.700 130.000 ;
        RECT 324.400 129.600 325.200 130.400 ;
        RECT 385.200 130.000 386.000 130.800 ;
        RECT 294.000 125.400 294.800 126.200 ;
        RECT 324.500 124.400 325.100 129.600 ;
        RECT 385.300 124.400 385.900 130.000 ;
        RECT 31.600 123.600 32.400 124.400 ;
        RECT 239.600 123.600 240.400 124.400 ;
        RECT 324.400 123.600 325.200 124.400 ;
        RECT 385.200 123.600 386.000 124.400 ;
        RECT 149.600 120.600 154.400 121.400 ;
        RECT 456.800 120.600 461.600 121.400 ;
        RECT 374.000 117.600 374.800 118.400 ;
        RECT 268.400 115.800 269.200 116.600 ;
        RECT 340.400 115.800 341.200 116.600 ;
        RECT 268.500 110.400 269.100 115.800 ;
        RECT 340.500 112.000 341.100 115.800 ;
        RECT 374.100 112.400 374.700 117.600 ;
        RECT 596.400 115.800 597.200 116.600 ;
        RECT 340.400 111.200 341.200 112.000 ;
        RECT 374.000 111.600 374.800 112.400 ;
        RECT 596.500 112.000 597.100 115.800 ;
        RECT 596.400 111.200 597.200 112.000 ;
        RECT 268.400 109.600 269.200 110.400 ;
        RECT 340.400 91.600 341.200 92.400 ;
        RECT 183.600 90.000 184.400 90.800 ;
        RECT 276.400 90.000 277.200 90.800 ;
        RECT 183.700 86.200 184.300 90.000 ;
        RECT 183.600 85.400 184.400 86.200 ;
        RECT 276.500 84.400 277.100 90.000 ;
        RECT 287.600 89.600 288.400 90.400 ;
        RECT 287.700 84.400 288.300 89.600 ;
        RECT 340.500 86.200 341.100 91.600 ;
        RECT 372.400 90.000 373.200 90.800 ;
        RECT 582.000 90.000 582.800 90.800 ;
        RECT 372.500 86.200 373.100 90.000 ;
        RECT 582.100 86.200 582.700 90.000 ;
        RECT 340.400 85.400 341.200 86.200 ;
        RECT 372.400 85.400 373.200 86.200 ;
        RECT 582.000 85.400 582.800 86.200 ;
        RECT 276.400 83.600 277.200 84.400 ;
        RECT 287.600 83.600 288.400 84.400 ;
        RECT 149.600 80.600 154.400 81.400 ;
        RECT 456.800 80.600 461.600 81.400 ;
        RECT 207.600 77.600 208.400 78.400 ;
        RECT 332.400 77.600 333.200 78.400 ;
        RECT 207.700 72.400 208.300 77.600 ;
        RECT 284.400 75.800 285.200 76.600 ;
        RECT 207.600 71.600 208.400 72.400 ;
        RECT 284.500 72.000 285.100 75.800 ;
        RECT 332.500 72.400 333.100 77.600 ;
        RECT 284.400 71.200 285.200 72.000 ;
        RECT 332.400 71.600 333.200 72.400 ;
        RECT 4.400 49.600 5.200 50.400 ;
        RECT 183.600 49.600 184.400 50.400 ;
        RECT 246.000 49.600 246.800 50.400 ;
        RECT 302.000 50.000 302.800 50.800 ;
        RECT 378.800 50.000 379.600 50.800 ;
        RECT 604.400 50.000 605.200 50.800 ;
        RECT 4.500 44.400 5.100 49.600 ;
        RECT 183.700 44.400 184.300 49.600 ;
        RECT 246.100 44.400 246.700 49.600 ;
        RECT 302.100 46.200 302.700 50.000 ;
        RECT 302.000 45.400 302.800 46.200 ;
        RECT 378.900 44.400 379.500 50.000 ;
        RECT 604.500 46.200 605.100 50.000 ;
        RECT 604.400 45.400 605.200 46.200 ;
        RECT 4.400 43.600 5.200 44.400 ;
        RECT 183.600 43.600 184.400 44.400 ;
        RECT 246.000 43.600 246.800 44.400 ;
        RECT 378.800 43.600 379.600 44.400 ;
        RECT 149.600 40.600 154.400 41.400 ;
        RECT 456.800 40.600 461.600 41.400 ;
        RECT 9.200 37.600 10.000 38.400 ;
        RECT 388.400 37.600 389.200 38.400 ;
        RECT 9.300 32.400 9.900 37.600 ;
        RECT 206.000 35.800 206.800 36.600 ;
        RECT 239.600 35.800 240.400 36.600 ;
        RECT 278.000 35.800 278.800 36.600 ;
        RECT 9.200 31.600 10.000 32.400 ;
        RECT 206.100 32.000 206.700 35.800 ;
        RECT 239.700 32.000 240.300 35.800 ;
        RECT 278.100 32.000 278.700 35.800 ;
        RECT 388.500 32.400 389.100 37.600 ;
        RECT 596.400 35.800 597.200 36.600 ;
        RECT 206.000 31.200 206.800 32.000 ;
        RECT 239.600 31.200 240.400 32.000 ;
        RECT 278.000 31.200 278.800 32.000 ;
        RECT 388.400 31.600 389.200 32.400 ;
        RECT 596.500 32.000 597.100 35.800 ;
        RECT 596.400 31.200 597.200 32.000 ;
        RECT 4.400 9.600 5.200 10.400 ;
        RECT 175.600 9.600 176.400 10.400 ;
        RECT 186.800 10.000 187.600 10.800 ;
        RECT 4.500 4.400 5.100 9.600 ;
        RECT 175.700 4.400 176.300 9.600 ;
        RECT 186.900 4.400 187.500 10.000 ;
        RECT 223.600 9.600 224.400 10.400 ;
        RECT 276.400 10.000 277.200 10.800 ;
        RECT 321.200 10.000 322.000 10.800 ;
        RECT 223.700 4.400 224.300 9.600 ;
        RECT 276.500 6.200 277.100 10.000 ;
        RECT 276.400 5.400 277.200 6.200 ;
        RECT 321.300 4.400 321.900 10.000 ;
        RECT 367.600 9.600 368.400 10.400 ;
        RECT 599.600 10.000 600.400 10.800 ;
        RECT 367.700 4.400 368.300 9.600 ;
        RECT 599.700 4.400 600.300 10.000 ;
        RECT 4.400 3.600 5.200 4.400 ;
        RECT 175.600 3.600 176.400 4.400 ;
        RECT 186.800 3.600 187.600 4.400 ;
        RECT 223.600 3.600 224.400 4.400 ;
        RECT 321.200 3.600 322.000 4.400 ;
        RECT 367.600 3.600 368.400 4.400 ;
        RECT 599.600 3.600 600.400 4.400 ;
        RECT 149.600 0.600 154.400 1.400 ;
        RECT 456.800 0.600 461.600 1.400 ;
      LAYER via2 ;
        RECT 150.200 560.600 151.000 561.400 ;
        RECT 151.600 560.600 152.400 561.400 ;
        RECT 153.000 560.600 153.800 561.400 ;
        RECT 457.400 560.600 458.200 561.400 ;
        RECT 458.800 560.600 459.600 561.400 ;
        RECT 460.200 560.600 461.000 561.400 ;
        RECT 150.200 520.600 151.000 521.400 ;
        RECT 151.600 520.600 152.400 521.400 ;
        RECT 153.000 520.600 153.800 521.400 ;
        RECT 457.400 520.600 458.200 521.400 ;
        RECT 458.800 520.600 459.600 521.400 ;
        RECT 460.200 520.600 461.000 521.400 ;
        RECT 150.200 480.600 151.000 481.400 ;
        RECT 151.600 480.600 152.400 481.400 ;
        RECT 153.000 480.600 153.800 481.400 ;
        RECT 457.400 480.600 458.200 481.400 ;
        RECT 458.800 480.600 459.600 481.400 ;
        RECT 460.200 480.600 461.000 481.400 ;
        RECT 150.200 440.600 151.000 441.400 ;
        RECT 151.600 440.600 152.400 441.400 ;
        RECT 153.000 440.600 153.800 441.400 ;
        RECT 457.400 440.600 458.200 441.400 ;
        RECT 458.800 440.600 459.600 441.400 ;
        RECT 460.200 440.600 461.000 441.400 ;
        RECT 150.200 400.600 151.000 401.400 ;
        RECT 151.600 400.600 152.400 401.400 ;
        RECT 153.000 400.600 153.800 401.400 ;
        RECT 457.400 400.600 458.200 401.400 ;
        RECT 458.800 400.600 459.600 401.400 ;
        RECT 460.200 400.600 461.000 401.400 ;
        RECT 150.200 360.600 151.000 361.400 ;
        RECT 151.600 360.600 152.400 361.400 ;
        RECT 153.000 360.600 153.800 361.400 ;
        RECT 457.400 360.600 458.200 361.400 ;
        RECT 458.800 360.600 459.600 361.400 ;
        RECT 460.200 360.600 461.000 361.400 ;
        RECT 150.200 320.600 151.000 321.400 ;
        RECT 151.600 320.600 152.400 321.400 ;
        RECT 153.000 320.600 153.800 321.400 ;
        RECT 457.400 320.600 458.200 321.400 ;
        RECT 458.800 320.600 459.600 321.400 ;
        RECT 460.200 320.600 461.000 321.400 ;
        RECT 150.200 280.600 151.000 281.400 ;
        RECT 151.600 280.600 152.400 281.400 ;
        RECT 153.000 280.600 153.800 281.400 ;
        RECT 457.400 280.600 458.200 281.400 ;
        RECT 458.800 280.600 459.600 281.400 ;
        RECT 460.200 280.600 461.000 281.400 ;
        RECT 150.200 240.600 151.000 241.400 ;
        RECT 151.600 240.600 152.400 241.400 ;
        RECT 153.000 240.600 153.800 241.400 ;
        RECT 457.400 240.600 458.200 241.400 ;
        RECT 458.800 240.600 459.600 241.400 ;
        RECT 460.200 240.600 461.000 241.400 ;
        RECT 150.200 200.600 151.000 201.400 ;
        RECT 151.600 200.600 152.400 201.400 ;
        RECT 153.000 200.600 153.800 201.400 ;
        RECT 457.400 200.600 458.200 201.400 ;
        RECT 458.800 200.600 459.600 201.400 ;
        RECT 460.200 200.600 461.000 201.400 ;
        RECT 150.200 160.600 151.000 161.400 ;
        RECT 151.600 160.600 152.400 161.400 ;
        RECT 153.000 160.600 153.800 161.400 ;
        RECT 457.400 160.600 458.200 161.400 ;
        RECT 458.800 160.600 459.600 161.400 ;
        RECT 460.200 160.600 461.000 161.400 ;
        RECT 150.200 120.600 151.000 121.400 ;
        RECT 151.600 120.600 152.400 121.400 ;
        RECT 153.000 120.600 153.800 121.400 ;
        RECT 457.400 120.600 458.200 121.400 ;
        RECT 458.800 120.600 459.600 121.400 ;
        RECT 460.200 120.600 461.000 121.400 ;
        RECT 150.200 80.600 151.000 81.400 ;
        RECT 151.600 80.600 152.400 81.400 ;
        RECT 153.000 80.600 153.800 81.400 ;
        RECT 457.400 80.600 458.200 81.400 ;
        RECT 458.800 80.600 459.600 81.400 ;
        RECT 460.200 80.600 461.000 81.400 ;
        RECT 150.200 40.600 151.000 41.400 ;
        RECT 151.600 40.600 152.400 41.400 ;
        RECT 153.000 40.600 153.800 41.400 ;
        RECT 457.400 40.600 458.200 41.400 ;
        RECT 458.800 40.600 459.600 41.400 ;
        RECT 460.200 40.600 461.000 41.400 ;
        RECT 150.200 0.600 151.000 1.400 ;
        RECT 151.600 0.600 152.400 1.400 ;
        RECT 153.000 0.600 153.800 1.400 ;
        RECT 457.400 0.600 458.200 1.400 ;
        RECT 458.800 0.600 459.600 1.400 ;
        RECT 460.200 0.600 461.000 1.400 ;
      LAYER metal3 ;
        RECT 149.600 560.400 154.400 561.600 ;
        RECT 456.800 560.400 461.600 561.600 ;
        RECT 149.600 520.400 154.400 521.600 ;
        RECT 456.800 520.400 461.600 521.600 ;
        RECT 149.600 480.400 154.400 481.600 ;
        RECT 456.800 480.400 461.600 481.600 ;
        RECT 149.600 440.400 154.400 441.600 ;
        RECT 456.800 440.400 461.600 441.600 ;
        RECT 149.600 400.400 154.400 401.600 ;
        RECT 456.800 400.400 461.600 401.600 ;
        RECT 149.600 360.400 154.400 361.600 ;
        RECT 456.800 360.400 461.600 361.600 ;
        RECT 149.600 320.400 154.400 321.600 ;
        RECT 456.800 320.400 461.600 321.600 ;
        RECT 149.600 280.400 154.400 281.600 ;
        RECT 456.800 280.400 461.600 281.600 ;
        RECT 149.600 240.400 154.400 241.600 ;
        RECT 456.800 240.400 461.600 241.600 ;
        RECT 149.600 200.400 154.400 201.600 ;
        RECT 456.800 200.400 461.600 201.600 ;
        RECT 149.600 160.400 154.400 161.600 ;
        RECT 456.800 160.400 461.600 161.600 ;
        RECT 149.600 120.400 154.400 121.600 ;
        RECT 456.800 120.400 461.600 121.600 ;
        RECT 149.600 80.400 154.400 81.600 ;
        RECT 456.800 80.400 461.600 81.600 ;
        RECT 149.600 40.400 154.400 41.600 ;
        RECT 456.800 40.400 461.600 41.600 ;
        RECT 149.600 0.400 154.400 1.600 ;
        RECT 456.800 0.400 461.600 1.600 ;
      LAYER via3 ;
        RECT 150.000 560.600 150.800 561.400 ;
        RECT 151.600 560.600 152.400 561.400 ;
        RECT 153.200 560.600 154.000 561.400 ;
        RECT 457.200 560.600 458.000 561.400 ;
        RECT 458.800 560.600 459.600 561.400 ;
        RECT 460.400 560.600 461.200 561.400 ;
        RECT 150.000 520.600 150.800 521.400 ;
        RECT 151.600 520.600 152.400 521.400 ;
        RECT 153.200 520.600 154.000 521.400 ;
        RECT 457.200 520.600 458.000 521.400 ;
        RECT 458.800 520.600 459.600 521.400 ;
        RECT 460.400 520.600 461.200 521.400 ;
        RECT 150.000 480.600 150.800 481.400 ;
        RECT 151.600 480.600 152.400 481.400 ;
        RECT 153.200 480.600 154.000 481.400 ;
        RECT 457.200 480.600 458.000 481.400 ;
        RECT 458.800 480.600 459.600 481.400 ;
        RECT 460.400 480.600 461.200 481.400 ;
        RECT 150.000 440.600 150.800 441.400 ;
        RECT 151.600 440.600 152.400 441.400 ;
        RECT 153.200 440.600 154.000 441.400 ;
        RECT 457.200 440.600 458.000 441.400 ;
        RECT 458.800 440.600 459.600 441.400 ;
        RECT 460.400 440.600 461.200 441.400 ;
        RECT 150.000 400.600 150.800 401.400 ;
        RECT 151.600 400.600 152.400 401.400 ;
        RECT 153.200 400.600 154.000 401.400 ;
        RECT 457.200 400.600 458.000 401.400 ;
        RECT 458.800 400.600 459.600 401.400 ;
        RECT 460.400 400.600 461.200 401.400 ;
        RECT 150.000 360.600 150.800 361.400 ;
        RECT 151.600 360.600 152.400 361.400 ;
        RECT 153.200 360.600 154.000 361.400 ;
        RECT 457.200 360.600 458.000 361.400 ;
        RECT 458.800 360.600 459.600 361.400 ;
        RECT 460.400 360.600 461.200 361.400 ;
        RECT 150.000 320.600 150.800 321.400 ;
        RECT 151.600 320.600 152.400 321.400 ;
        RECT 153.200 320.600 154.000 321.400 ;
        RECT 457.200 320.600 458.000 321.400 ;
        RECT 458.800 320.600 459.600 321.400 ;
        RECT 460.400 320.600 461.200 321.400 ;
        RECT 150.000 280.600 150.800 281.400 ;
        RECT 151.600 280.600 152.400 281.400 ;
        RECT 153.200 280.600 154.000 281.400 ;
        RECT 457.200 280.600 458.000 281.400 ;
        RECT 458.800 280.600 459.600 281.400 ;
        RECT 460.400 280.600 461.200 281.400 ;
        RECT 150.000 240.600 150.800 241.400 ;
        RECT 151.600 240.600 152.400 241.400 ;
        RECT 153.200 240.600 154.000 241.400 ;
        RECT 457.200 240.600 458.000 241.400 ;
        RECT 458.800 240.600 459.600 241.400 ;
        RECT 460.400 240.600 461.200 241.400 ;
        RECT 150.000 200.600 150.800 201.400 ;
        RECT 151.600 200.600 152.400 201.400 ;
        RECT 153.200 200.600 154.000 201.400 ;
        RECT 457.200 200.600 458.000 201.400 ;
        RECT 458.800 200.600 459.600 201.400 ;
        RECT 460.400 200.600 461.200 201.400 ;
        RECT 150.000 160.600 150.800 161.400 ;
        RECT 151.600 160.600 152.400 161.400 ;
        RECT 153.200 160.600 154.000 161.400 ;
        RECT 457.200 160.600 458.000 161.400 ;
        RECT 458.800 160.600 459.600 161.400 ;
        RECT 460.400 160.600 461.200 161.400 ;
        RECT 150.000 120.600 150.800 121.400 ;
        RECT 151.600 120.600 152.400 121.400 ;
        RECT 153.200 120.600 154.000 121.400 ;
        RECT 457.200 120.600 458.000 121.400 ;
        RECT 458.800 120.600 459.600 121.400 ;
        RECT 460.400 120.600 461.200 121.400 ;
        RECT 150.000 80.600 150.800 81.400 ;
        RECT 151.600 80.600 152.400 81.400 ;
        RECT 153.200 80.600 154.000 81.400 ;
        RECT 457.200 80.600 458.000 81.400 ;
        RECT 458.800 80.600 459.600 81.400 ;
        RECT 460.400 80.600 461.200 81.400 ;
        RECT 150.000 40.600 150.800 41.400 ;
        RECT 151.600 40.600 152.400 41.400 ;
        RECT 153.200 40.600 154.000 41.400 ;
        RECT 457.200 40.600 458.000 41.400 ;
        RECT 458.800 40.600 459.600 41.400 ;
        RECT 460.400 40.600 461.200 41.400 ;
        RECT 150.000 0.600 150.800 1.400 ;
        RECT 151.600 0.600 152.400 1.400 ;
        RECT 153.200 0.600 154.000 1.400 ;
        RECT 457.200 0.600 458.000 1.400 ;
        RECT 458.800 0.600 459.600 1.400 ;
        RECT 460.400 0.600 461.200 1.400 ;
      LAYER metal4 ;
        RECT 149.600 -4.000 154.400 564.000 ;
        RECT 456.800 -4.000 461.600 564.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 2.800 541.600 3.600 544.200 ;
        RECT 7.600 541.600 8.400 546.200 ;
        RECT 17.200 541.600 18.000 544.200 ;
        RECT 20.400 541.600 21.200 544.200 ;
        RECT 31.600 541.600 32.400 546.200 ;
        RECT 38.000 541.600 38.800 544.200 ;
        RECT 41.200 541.600 42.000 546.200 ;
        RECT 44.400 541.600 45.200 546.200 ;
        RECT 50.800 541.600 51.600 544.200 ;
        RECT 54.000 541.600 54.800 545.400 ;
        RECT 60.400 541.600 61.200 545.400 ;
        RECT 65.200 541.600 66.000 544.200 ;
        RECT 71.600 541.600 72.400 546.200 ;
        RECT 82.800 541.600 83.600 544.200 ;
        RECT 86.000 541.600 86.800 544.200 ;
        RECT 95.600 541.600 96.400 546.200 ;
        RECT 102.000 541.600 102.800 546.200 ;
        RECT 107.400 541.600 108.400 544.200 ;
        RECT 110.800 541.600 111.600 544.200 ;
        RECT 116.400 541.600 117.200 546.000 ;
        RECT 121.200 541.600 122.000 546.200 ;
        RECT 126.600 541.600 127.600 544.200 ;
        RECT 130.000 541.600 130.800 544.200 ;
        RECT 135.600 541.600 136.400 546.000 ;
        RECT 146.800 541.600 147.600 546.200 ;
        RECT 156.400 541.600 157.200 544.200 ;
        RECT 159.600 541.600 160.400 544.200 ;
        RECT 170.800 541.600 171.600 546.200 ;
        RECT 177.200 541.600 178.000 544.200 ;
        RECT 180.400 541.600 181.200 546.200 ;
        RECT 183.600 541.600 184.400 544.200 ;
        RECT 190.000 541.600 190.800 545.400 ;
        RECT 193.200 541.600 194.000 546.200 ;
        RECT 199.600 541.600 200.400 546.200 ;
        RECT 206.000 541.600 206.800 546.200 ;
        RECT 215.600 541.600 216.400 544.200 ;
        RECT 218.800 541.600 219.600 544.200 ;
        RECT 230.000 541.600 230.800 546.200 ;
        RECT 236.400 541.600 237.200 544.200 ;
        RECT 238.000 541.600 238.800 544.200 ;
        RECT 242.800 541.600 243.600 545.400 ;
        RECT 247.600 541.600 248.400 546.200 ;
        RECT 254.000 541.600 254.800 546.200 ;
        RECT 260.400 541.600 261.200 546.200 ;
        RECT 270.000 541.600 270.800 544.200 ;
        RECT 273.200 541.600 274.000 544.200 ;
        RECT 284.400 541.600 285.200 546.200 ;
        RECT 290.800 541.600 291.600 544.200 ;
        RECT 294.000 541.600 294.800 546.200 ;
        RECT 302.000 541.600 302.800 544.200 ;
        RECT 308.400 541.600 309.200 546.200 ;
        RECT 319.600 541.600 320.400 544.200 ;
        RECT 322.800 541.600 323.600 544.200 ;
        RECT 332.400 541.600 333.200 546.200 ;
        RECT 337.200 541.600 338.000 544.200 ;
        RECT 342.000 541.600 342.800 545.400 ;
        RECT 350.000 541.600 350.800 545.400 ;
        RECT 353.200 541.600 354.000 544.200 ;
        RECT 358.000 541.600 358.800 545.400 ;
        RECT 364.400 541.600 365.200 545.400 ;
        RECT 369.200 541.600 370.000 544.200 ;
        RECT 375.600 541.600 376.400 546.200 ;
        RECT 386.800 541.600 387.600 544.200 ;
        RECT 390.000 541.600 390.800 544.200 ;
        RECT 399.600 541.600 400.400 546.200 ;
        RECT 404.400 541.600 405.200 546.200 ;
        RECT 407.600 541.600 408.400 546.200 ;
        RECT 410.800 541.600 411.600 546.200 ;
        RECT 414.000 541.600 414.800 546.200 ;
        RECT 417.200 541.600 418.000 546.200 ;
        RECT 420.400 541.600 421.200 546.000 ;
        RECT 426.000 541.600 426.800 544.200 ;
        RECT 429.200 541.600 430.200 544.200 ;
        RECT 434.800 541.600 435.600 546.200 ;
        RECT 439.600 541.600 440.400 545.400 ;
        RECT 447.600 541.600 448.400 545.400 ;
        RECT 452.400 541.600 453.200 545.800 ;
        RECT 455.600 541.600 456.400 544.200 ;
        RECT 463.600 541.600 464.400 546.000 ;
        RECT 469.200 541.600 470.000 544.200 ;
        RECT 472.400 541.600 473.400 544.200 ;
        RECT 478.000 541.600 478.800 546.200 ;
        RECT 482.800 541.600 483.600 545.400 ;
        RECT 490.800 541.600 491.600 545.400 ;
        RECT 495.600 541.600 496.400 546.000 ;
        RECT 501.200 541.600 502.000 544.200 ;
        RECT 504.400 541.600 505.400 544.200 ;
        RECT 510.000 541.600 510.800 546.200 ;
        RECT 514.800 541.600 515.600 545.400 ;
        RECT 521.200 541.600 522.000 546.600 ;
        RECT 526.400 541.600 527.200 547.000 ;
        RECT 532.400 541.600 533.200 545.400 ;
        RECT 535.600 541.600 536.400 544.200 ;
        RECT 540.400 541.600 541.200 546.000 ;
        RECT 546.000 541.600 546.800 544.200 ;
        RECT 549.200 541.600 550.200 544.200 ;
        RECT 554.800 541.600 555.600 546.200 ;
        RECT 558.000 541.600 558.800 544.200 ;
        RECT 564.400 541.600 565.200 546.200 ;
        RECT 575.600 541.600 576.400 544.200 ;
        RECT 578.800 541.600 579.600 544.200 ;
        RECT 588.400 541.600 589.200 546.200 ;
        RECT 594.800 541.600 595.600 544.200 ;
        RECT 596.400 541.600 597.200 546.200 ;
        RECT 599.600 541.600 600.400 546.200 ;
        RECT 602.800 541.600 603.600 546.200 ;
        RECT 606.000 541.600 606.800 546.200 ;
        RECT 609.200 541.600 610.000 546.200 ;
        RECT 0.400 540.400 614.000 541.600 ;
        RECT 4.400 535.800 5.200 540.400 ;
        RECT 14.000 537.800 14.800 540.400 ;
        RECT 17.200 537.800 18.000 540.400 ;
        RECT 28.400 535.800 29.200 540.400 ;
        RECT 34.800 537.800 35.600 540.400 ;
        RECT 39.600 536.600 40.400 540.400 ;
        RECT 46.000 535.800 46.800 540.400 ;
        RECT 47.600 537.800 48.400 540.400 ;
        RECT 52.400 536.600 53.200 540.400 ;
        RECT 58.800 536.600 59.600 540.400 ;
        RECT 63.600 537.800 64.400 540.400 ;
        RECT 70.000 535.800 70.800 540.400 ;
        RECT 81.200 537.800 82.000 540.400 ;
        RECT 84.400 537.800 85.200 540.400 ;
        RECT 94.000 535.800 94.800 540.400 ;
        RECT 100.400 536.600 101.200 540.400 ;
        RECT 106.800 536.600 107.600 540.400 ;
        RECT 113.200 536.600 114.000 540.400 ;
        RECT 121.200 536.600 122.000 540.400 ;
        RECT 126.200 539.800 127.000 540.400 ;
        RECT 126.000 536.400 127.000 539.800 ;
        RECT 132.200 536.400 133.200 540.400 ;
        RECT 140.400 537.800 141.200 540.400 ;
        RECT 146.800 535.800 147.600 540.400 ;
        RECT 158.000 537.800 158.800 540.400 ;
        RECT 161.200 537.800 162.000 540.400 ;
        RECT 170.800 535.800 171.600 540.400 ;
        RECT 178.800 535.800 179.600 540.400 ;
        RECT 188.400 537.800 189.200 540.400 ;
        RECT 191.600 537.800 192.400 540.400 ;
        RECT 202.800 535.800 203.600 540.400 ;
        RECT 209.200 537.800 210.000 540.400 ;
        RECT 210.800 537.800 211.600 540.400 ;
        RECT 215.600 536.600 216.400 540.400 ;
        RECT 223.600 535.800 224.400 540.400 ;
        RECT 225.200 537.800 226.000 540.400 ;
        RECT 231.600 535.800 232.400 540.400 ;
        RECT 242.800 537.800 243.600 540.400 ;
        RECT 246.000 537.800 246.800 540.400 ;
        RECT 255.600 535.800 256.400 540.400 ;
        RECT 263.600 535.800 264.400 540.400 ;
        RECT 273.200 537.800 274.000 540.400 ;
        RECT 276.400 537.800 277.200 540.400 ;
        RECT 287.600 535.800 288.400 540.400 ;
        RECT 294.000 537.800 294.800 540.400 ;
        RECT 295.600 537.800 296.400 540.400 ;
        RECT 300.400 536.600 301.200 540.400 ;
        RECT 310.000 535.800 310.800 540.400 ;
        RECT 314.800 537.800 315.600 540.400 ;
        RECT 321.200 535.800 322.000 540.400 ;
        RECT 332.400 537.800 333.200 540.400 ;
        RECT 335.600 537.800 336.400 540.400 ;
        RECT 345.200 535.800 346.000 540.400 ;
        RECT 353.200 536.600 354.000 540.400 ;
        RECT 358.000 537.800 358.800 540.400 ;
        RECT 362.800 536.600 363.600 540.400 ;
        RECT 367.600 536.600 368.400 540.400 ;
        RECT 372.400 537.800 373.200 540.400 ;
        RECT 377.200 536.600 378.000 540.400 ;
        RECT 382.000 537.800 382.800 540.400 ;
        RECT 388.400 535.800 389.200 540.400 ;
        RECT 399.600 537.800 400.400 540.400 ;
        RECT 402.800 537.800 403.600 540.400 ;
        RECT 412.400 535.800 413.200 540.400 ;
        RECT 417.200 535.800 418.000 540.400 ;
        RECT 420.400 535.800 421.200 540.400 ;
        RECT 423.600 535.800 424.400 540.400 ;
        RECT 426.800 535.800 427.600 540.400 ;
        RECT 430.000 535.800 430.800 540.400 ;
        RECT 433.200 536.000 434.000 540.400 ;
        RECT 438.800 537.800 439.600 540.400 ;
        RECT 442.000 537.800 443.000 540.400 ;
        RECT 447.600 535.800 448.400 540.400 ;
        RECT 452.400 536.600 453.200 540.400 ;
        RECT 465.200 536.600 466.000 540.400 ;
        RECT 470.000 535.800 470.800 540.400 ;
        RECT 473.200 535.800 474.000 540.400 ;
        RECT 476.400 536.600 477.200 540.400 ;
        RECT 484.400 536.600 485.200 540.400 ;
        RECT 489.200 536.600 490.000 540.400 ;
        RECT 497.200 536.600 498.000 540.400 ;
        RECT 502.000 535.800 502.800 540.400 ;
        RECT 507.400 537.800 508.400 540.400 ;
        RECT 510.800 537.800 511.600 540.400 ;
        RECT 516.400 536.000 517.200 540.400 ;
        RECT 522.800 535.800 523.600 540.400 ;
        RECT 526.000 535.800 526.800 540.400 ;
        RECT 529.200 535.800 530.000 540.400 ;
        RECT 532.400 535.800 533.200 540.400 ;
        RECT 535.600 535.800 536.400 540.400 ;
        RECT 538.800 536.600 539.600 540.400 ;
        RECT 543.600 537.800 544.400 540.400 ;
        RECT 550.000 535.800 550.800 540.400 ;
        RECT 561.200 537.800 562.000 540.400 ;
        RECT 564.400 537.800 565.200 540.400 ;
        RECT 574.000 535.800 574.800 540.400 ;
        RECT 580.400 536.600 581.200 540.400 ;
        RECT 585.200 535.800 586.000 540.400 ;
        RECT 588.400 535.800 589.200 540.400 ;
        RECT 591.600 535.800 592.400 540.400 ;
        RECT 594.800 535.800 595.600 540.400 ;
        RECT 598.000 535.800 598.800 540.400 ;
        RECT 602.800 536.600 603.600 540.400 ;
        RECT 607.600 537.800 608.400 540.400 ;
        RECT 2.800 501.600 3.600 506.200 ;
        RECT 8.200 501.600 9.200 504.200 ;
        RECT 11.600 501.600 12.400 504.200 ;
        RECT 17.200 501.600 18.000 506.000 ;
        RECT 22.000 501.600 22.800 506.200 ;
        RECT 27.400 501.600 28.400 504.200 ;
        RECT 30.800 501.600 31.600 504.200 ;
        RECT 36.400 501.600 37.200 506.000 ;
        RECT 41.200 501.600 42.000 505.400 ;
        RECT 47.600 501.600 48.400 506.600 ;
        RECT 52.800 501.600 53.600 507.000 ;
        RECT 58.800 501.600 59.600 505.400 ;
        RECT 63.600 501.600 64.400 505.400 ;
        RECT 71.600 501.600 72.400 505.400 ;
        RECT 76.400 501.600 77.200 506.200 ;
        RECT 81.800 501.600 82.800 504.200 ;
        RECT 85.200 501.600 86.000 504.200 ;
        RECT 90.800 501.600 91.600 506.000 ;
        RECT 95.600 501.600 96.400 506.200 ;
        RECT 101.000 501.600 102.000 504.200 ;
        RECT 104.400 501.600 105.200 504.200 ;
        RECT 110.000 501.600 110.800 506.000 ;
        RECT 114.800 501.600 115.600 504.200 ;
        RECT 116.400 501.600 117.200 504.200 ;
        RECT 120.800 501.600 121.600 507.000 ;
        RECT 126.000 501.600 126.800 506.600 ;
        RECT 130.800 501.600 131.600 506.600 ;
        RECT 136.000 501.600 136.800 507.000 ;
        RECT 138.800 501.600 139.600 504.200 ;
        RECT 142.000 501.600 142.800 504.200 ;
        RECT 143.600 501.600 144.400 504.200 ;
        RECT 151.600 501.600 152.400 506.200 ;
        RECT 154.800 501.600 155.600 506.200 ;
        RECT 158.000 501.600 158.800 506.200 ;
        RECT 161.200 501.600 162.000 506.200 ;
        RECT 164.400 501.600 165.200 506.200 ;
        RECT 166.000 501.600 166.800 504.200 ;
        RECT 169.200 501.600 170.000 504.200 ;
        RECT 172.400 501.600 173.200 504.200 ;
        RECT 175.600 501.600 176.600 505.600 ;
        RECT 181.800 502.200 182.800 505.600 ;
        RECT 181.800 501.600 182.600 502.200 ;
        RECT 185.200 501.600 186.000 506.200 ;
        RECT 188.400 501.600 189.200 506.200 ;
        RECT 191.600 501.600 192.400 506.200 ;
        RECT 194.800 501.600 195.600 506.200 ;
        RECT 198.000 501.600 198.800 506.200 ;
        RECT 202.800 501.600 203.600 506.200 ;
        RECT 212.400 501.600 213.200 504.200 ;
        RECT 215.600 501.600 216.400 504.200 ;
        RECT 226.800 501.600 227.600 506.200 ;
        RECT 233.200 501.600 234.000 504.200 ;
        RECT 238.000 501.600 238.800 505.400 ;
        RECT 241.200 501.600 242.000 506.200 ;
        RECT 246.000 501.600 246.800 504.200 ;
        RECT 252.400 501.600 253.200 506.200 ;
        RECT 262.000 501.600 262.800 504.200 ;
        RECT 265.200 501.600 266.000 504.200 ;
        RECT 276.400 501.600 277.200 506.200 ;
        RECT 282.800 501.600 283.600 504.200 ;
        RECT 287.600 501.600 288.400 506.200 ;
        RECT 297.200 501.600 298.000 504.200 ;
        RECT 300.400 501.600 301.200 504.200 ;
        RECT 311.600 501.600 312.400 506.200 ;
        RECT 318.000 501.600 318.800 504.200 ;
        RECT 327.600 501.600 328.400 506.200 ;
        RECT 332.400 501.600 333.200 506.200 ;
        RECT 335.600 501.600 336.400 506.200 ;
        RECT 341.000 501.600 342.000 504.200 ;
        RECT 344.400 501.600 345.200 504.200 ;
        RECT 350.000 501.600 350.800 506.000 ;
        RECT 353.200 501.600 354.000 506.200 ;
        RECT 359.600 501.600 360.400 506.200 ;
        RECT 365.000 501.600 366.000 504.200 ;
        RECT 368.400 501.600 369.200 504.200 ;
        RECT 374.000 501.600 374.800 506.000 ;
        RECT 378.800 501.600 379.600 506.600 ;
        RECT 384.000 501.600 384.800 507.000 ;
        RECT 388.400 501.600 389.200 505.400 ;
        RECT 396.400 501.600 397.200 506.200 ;
        RECT 401.200 501.600 402.000 505.400 ;
        RECT 404.400 501.600 405.200 506.200 ;
        RECT 407.600 501.600 408.400 506.200 ;
        RECT 410.800 501.600 411.600 504.200 ;
        RECT 415.200 501.600 416.000 507.000 ;
        RECT 420.400 501.600 421.200 506.600 ;
        RECT 425.200 501.600 426.000 505.400 ;
        RECT 430.000 501.600 430.800 506.200 ;
        RECT 433.200 501.600 434.000 506.200 ;
        RECT 439.600 501.600 440.400 506.200 ;
        RECT 442.800 501.600 443.600 506.200 ;
        RECT 446.000 501.600 446.800 506.200 ;
        RECT 448.800 501.600 449.600 507.000 ;
        RECT 454.000 501.600 454.800 506.600 ;
        RECT 463.600 501.600 464.400 504.200 ;
        RECT 468.400 501.600 469.200 506.200 ;
        RECT 471.600 501.600 472.400 506.600 ;
        RECT 476.800 501.600 477.600 507.000 ;
        RECT 479.600 501.600 480.400 506.200 ;
        RECT 485.600 501.600 486.400 507.000 ;
        RECT 490.800 501.600 491.600 506.600 ;
        RECT 494.000 501.600 494.800 506.200 ;
        RECT 497.200 501.600 498.000 506.200 ;
        RECT 500.400 501.600 501.200 506.200 ;
        RECT 506.800 501.600 507.600 506.200 ;
        RECT 510.000 501.600 510.800 506.200 ;
        RECT 513.200 501.600 514.000 505.400 ;
        RECT 519.600 501.600 520.400 504.200 ;
        RECT 522.800 501.600 523.600 506.600 ;
        RECT 528.000 501.600 528.800 507.000 ;
        RECT 532.400 501.600 533.200 505.400 ;
        RECT 538.800 501.600 539.600 505.400 ;
        RECT 545.200 501.600 546.000 505.400 ;
        RECT 551.600 501.600 552.400 506.000 ;
        RECT 557.200 501.600 558.000 504.200 ;
        RECT 560.400 501.600 561.400 504.200 ;
        RECT 566.000 501.600 566.800 506.200 ;
        RECT 572.400 501.600 573.200 506.200 ;
        RECT 574.000 501.600 574.800 504.200 ;
        RECT 580.400 501.600 581.200 506.200 ;
        RECT 591.600 501.600 592.400 504.200 ;
        RECT 594.800 501.600 595.600 504.200 ;
        RECT 604.400 501.600 605.200 506.200 ;
        RECT 0.400 500.400 614.000 501.600 ;
        RECT 4.400 496.600 5.200 500.400 ;
        RECT 8.800 495.000 9.600 500.400 ;
        RECT 14.000 495.400 14.800 500.400 ;
        RECT 20.400 496.600 21.200 500.400 ;
        RECT 25.200 495.800 26.000 500.400 ;
        RECT 30.600 497.800 31.600 500.400 ;
        RECT 34.000 497.800 34.800 500.400 ;
        RECT 39.600 496.000 40.400 500.400 ;
        RECT 44.400 496.600 45.200 500.400 ;
        RECT 50.400 495.000 51.200 500.400 ;
        RECT 55.600 495.400 56.400 500.400 ;
        RECT 62.000 496.600 62.800 500.400 ;
        RECT 66.800 495.400 67.600 500.400 ;
        RECT 72.000 495.000 72.800 500.400 ;
        RECT 74.800 495.800 75.600 500.400 ;
        RECT 79.600 495.800 80.400 500.400 ;
        RECT 84.400 497.800 85.200 500.400 ;
        RECT 89.200 496.600 90.000 500.400 ;
        RECT 97.200 496.600 98.000 500.400 ;
        RECT 103.600 496.600 104.400 500.400 ;
        RECT 106.800 493.800 107.600 500.400 ;
        RECT 116.400 496.600 117.200 500.400 ;
        RECT 119.600 495.800 120.400 500.400 ;
        RECT 124.400 497.800 125.200 500.400 ;
        RECT 127.600 497.800 128.400 500.400 ;
        RECT 129.200 497.800 130.000 500.400 ;
        RECT 135.600 495.800 136.400 500.400 ;
        RECT 146.800 497.800 147.600 500.400 ;
        RECT 150.000 497.800 150.800 500.400 ;
        RECT 159.600 495.800 160.400 500.400 ;
        RECT 169.200 497.800 170.000 500.400 ;
        RECT 172.400 497.800 173.200 500.400 ;
        RECT 174.000 497.800 174.800 500.400 ;
        RECT 180.400 495.800 181.200 500.400 ;
        RECT 191.600 497.800 192.400 500.400 ;
        RECT 194.800 497.800 195.600 500.400 ;
        RECT 204.400 495.800 205.200 500.400 ;
        RECT 209.200 497.800 210.000 500.400 ;
        RECT 215.600 495.800 216.400 500.400 ;
        RECT 226.800 497.800 227.600 500.400 ;
        RECT 230.000 497.800 230.800 500.400 ;
        RECT 239.600 495.800 240.400 500.400 ;
        RECT 246.000 495.800 246.800 500.400 ;
        RECT 249.200 495.800 250.000 500.400 ;
        RECT 250.800 495.800 251.600 500.400 ;
        RECT 254.000 495.800 254.800 500.400 ;
        RECT 257.200 495.800 258.000 500.400 ;
        RECT 260.400 495.800 261.200 500.400 ;
        RECT 263.600 495.800 264.400 500.400 ;
        RECT 265.200 495.800 266.000 500.400 ;
        RECT 268.400 495.800 269.200 500.400 ;
        RECT 271.600 495.800 272.400 500.400 ;
        RECT 274.800 495.800 275.600 500.400 ;
        RECT 278.000 495.800 278.800 500.400 ;
        RECT 282.800 496.600 283.600 500.400 ;
        RECT 286.000 495.800 286.800 500.400 ;
        RECT 292.400 496.600 293.200 500.400 ;
        RECT 298.800 496.600 299.600 500.400 ;
        RECT 309.600 495.000 310.400 500.400 ;
        RECT 314.800 495.400 315.600 500.400 ;
        RECT 318.000 495.800 318.800 500.400 ;
        RECT 321.200 495.800 322.000 500.400 ;
        RECT 326.000 496.600 326.800 500.400 ;
        RECT 330.800 497.800 331.600 500.400 ;
        RECT 334.000 497.800 334.800 500.400 ;
        RECT 337.200 495.800 338.000 500.400 ;
        RECT 340.400 495.800 341.200 500.400 ;
        RECT 345.200 496.600 346.000 500.400 ;
        RECT 349.600 495.000 350.400 500.400 ;
        RECT 354.800 495.400 355.600 500.400 ;
        RECT 359.600 496.600 360.400 500.400 ;
        RECT 367.600 496.600 368.400 500.400 ;
        RECT 372.000 495.000 372.800 500.400 ;
        RECT 377.200 495.400 378.000 500.400 ;
        RECT 382.000 496.000 382.800 500.400 ;
        RECT 387.600 497.800 388.400 500.400 ;
        RECT 390.800 497.800 391.800 500.400 ;
        RECT 396.400 495.800 397.200 500.400 ;
        RECT 401.200 496.600 402.000 500.400 ;
        RECT 409.200 496.600 410.000 500.400 ;
        RECT 414.000 495.800 414.800 500.400 ;
        RECT 419.400 497.800 420.400 500.400 ;
        RECT 422.800 497.800 423.600 500.400 ;
        RECT 428.400 496.000 429.200 500.400 ;
        RECT 432.800 495.000 433.600 500.400 ;
        RECT 438.000 495.400 438.800 500.400 ;
        RECT 442.800 496.600 443.600 500.400 ;
        RECT 450.800 496.600 451.600 500.400 ;
        RECT 455.600 496.600 456.400 500.400 ;
        RECT 466.800 496.600 467.600 500.400 ;
        RECT 474.800 496.600 475.600 500.400 ;
        RECT 479.600 496.000 480.400 500.400 ;
        RECT 485.200 497.800 486.000 500.400 ;
        RECT 488.400 497.800 489.400 500.400 ;
        RECT 494.000 495.800 494.800 500.400 ;
        RECT 498.800 495.400 499.600 500.400 ;
        RECT 504.000 495.000 504.800 500.400 ;
        RECT 508.400 496.600 509.200 500.400 ;
        RECT 516.400 496.600 517.200 500.400 ;
        RECT 521.200 496.000 522.000 500.400 ;
        RECT 526.800 497.800 527.600 500.400 ;
        RECT 530.000 497.800 531.000 500.400 ;
        RECT 535.600 495.800 536.400 500.400 ;
        RECT 540.400 496.600 541.200 500.400 ;
        RECT 546.800 496.600 547.600 500.400 ;
        RECT 553.200 496.000 554.000 500.400 ;
        RECT 558.800 497.800 559.600 500.400 ;
        RECT 562.000 497.800 563.000 500.400 ;
        RECT 567.600 495.800 568.400 500.400 ;
        RECT 574.000 496.600 574.800 500.400 ;
        RECT 577.200 497.800 578.000 500.400 ;
        RECT 583.600 495.800 584.400 500.400 ;
        RECT 594.800 497.800 595.600 500.400 ;
        RECT 598.000 497.800 598.800 500.400 ;
        RECT 607.600 495.800 608.400 500.400 ;
        RECT 2.800 461.600 3.600 466.200 ;
        RECT 8.200 461.600 9.200 464.200 ;
        RECT 11.600 461.600 12.400 464.200 ;
        RECT 17.200 461.600 18.000 466.000 ;
        RECT 22.000 461.600 22.800 465.400 ;
        RECT 30.000 461.600 30.800 465.400 ;
        RECT 34.800 461.600 35.600 466.200 ;
        RECT 40.200 461.600 41.200 464.200 ;
        RECT 43.600 461.600 44.400 464.200 ;
        RECT 49.200 461.600 50.000 466.000 ;
        RECT 54.000 461.600 54.800 465.400 ;
        RECT 62.000 461.600 62.800 465.400 ;
        RECT 66.400 461.600 67.200 467.000 ;
        RECT 71.600 461.600 72.400 466.600 ;
        RECT 78.000 461.600 78.800 466.200 ;
        RECT 80.800 461.600 81.600 467.000 ;
        RECT 86.000 461.600 86.800 466.600 ;
        RECT 89.200 461.600 90.000 466.200 ;
        RECT 92.400 461.600 93.200 466.200 ;
        RECT 96.800 461.600 97.600 467.000 ;
        RECT 102.000 461.600 102.800 466.600 ;
        RECT 105.200 461.600 106.000 466.200 ;
        RECT 108.400 461.600 109.200 466.200 ;
        RECT 111.600 461.600 112.400 464.200 ;
        RECT 114.800 461.600 115.600 468.200 ;
        RECT 124.400 461.600 125.200 465.400 ;
        RECT 130.800 461.600 131.600 465.400 ;
        RECT 135.600 461.600 136.400 465.400 ;
        RECT 140.400 461.600 141.200 464.200 ;
        RECT 143.600 461.600 144.400 464.200 ;
        RECT 146.800 461.600 147.600 465.400 ;
        RECT 158.000 461.600 158.800 466.200 ;
        RECT 161.200 461.600 162.000 466.200 ;
        RECT 164.000 461.600 164.800 467.000 ;
        RECT 169.200 461.600 170.000 466.600 ;
        RECT 174.000 461.600 174.800 465.400 ;
        RECT 180.400 461.600 181.200 465.400 ;
        RECT 186.800 461.600 187.600 466.000 ;
        RECT 192.400 461.600 193.200 464.200 ;
        RECT 195.600 461.600 196.600 464.200 ;
        RECT 201.200 461.600 202.000 466.200 ;
        RECT 204.400 461.600 205.200 466.200 ;
        RECT 209.200 461.600 210.000 466.200 ;
        RECT 214.000 461.600 214.800 465.400 ;
        RECT 222.000 461.600 222.800 465.400 ;
        RECT 226.800 461.600 227.800 465.600 ;
        RECT 233.000 462.200 234.000 465.600 ;
        RECT 233.000 461.600 233.800 462.200 ;
        RECT 239.600 461.600 240.400 465.400 ;
        RECT 242.800 461.600 243.600 464.200 ;
        RECT 246.000 461.600 246.800 464.200 ;
        RECT 249.200 461.600 250.000 466.200 ;
        RECT 252.400 461.600 253.200 466.200 ;
        RECT 257.200 461.600 258.000 466.200 ;
        RECT 266.800 461.600 267.600 464.200 ;
        RECT 270.000 461.600 270.800 464.200 ;
        RECT 281.200 461.600 282.000 466.200 ;
        RECT 287.600 461.600 288.400 464.200 ;
        RECT 289.200 461.600 290.000 466.200 ;
        RECT 294.000 461.600 294.800 464.200 ;
        RECT 297.200 461.600 298.000 464.200 ;
        RECT 298.800 461.600 299.600 466.200 ;
        RECT 302.000 461.600 302.800 466.200 ;
        RECT 311.600 461.600 312.400 466.200 ;
        RECT 317.000 461.600 318.000 464.200 ;
        RECT 320.400 461.600 321.200 464.200 ;
        RECT 326.000 461.600 326.800 466.000 ;
        RECT 332.400 461.600 333.200 465.400 ;
        RECT 337.200 461.600 338.000 465.400 ;
        RECT 343.600 461.600 344.400 464.200 ;
        RECT 346.800 461.600 347.600 465.400 ;
        RECT 354.800 461.600 355.600 465.400 ;
        RECT 359.200 461.600 360.000 467.000 ;
        RECT 364.400 461.600 365.200 466.600 ;
        RECT 369.200 461.600 370.000 466.200 ;
        RECT 374.600 461.600 375.600 464.200 ;
        RECT 378.000 461.600 378.800 464.200 ;
        RECT 383.600 461.600 384.400 466.000 ;
        RECT 386.800 461.600 387.600 466.200 ;
        RECT 390.000 461.600 390.800 466.200 ;
        RECT 396.400 461.600 397.200 465.400 ;
        RECT 399.600 461.600 400.400 464.200 ;
        RECT 404.400 461.600 405.200 466.200 ;
        RECT 409.800 461.600 410.800 464.200 ;
        RECT 413.200 461.600 414.000 464.200 ;
        RECT 418.800 461.600 419.600 466.000 ;
        RECT 422.000 461.600 422.800 466.200 ;
        RECT 426.800 461.600 427.600 466.200 ;
        RECT 433.200 461.600 434.000 465.400 ;
        RECT 441.200 461.600 442.000 465.400 ;
        RECT 446.000 461.600 446.800 466.600 ;
        RECT 451.200 461.600 452.000 467.000 ;
        RECT 460.000 461.600 460.800 467.000 ;
        RECT 465.200 461.600 466.000 466.600 ;
        RECT 468.400 461.600 469.200 466.200 ;
        RECT 474.800 461.600 475.600 465.400 ;
        RECT 479.600 461.600 480.400 466.200 ;
        RECT 482.800 461.600 483.600 466.200 ;
        RECT 487.600 461.600 488.400 466.600 ;
        RECT 492.800 461.600 493.600 467.000 ;
        RECT 495.600 461.600 496.400 464.200 ;
        RECT 500.400 461.600 501.200 465.400 ;
        RECT 505.200 461.600 506.000 466.200 ;
        RECT 510.000 461.600 510.800 464.200 ;
        RECT 513.200 461.600 514.000 464.200 ;
        RECT 514.800 461.600 515.600 464.200 ;
        RECT 518.000 461.600 518.800 464.200 ;
        RECT 521.200 461.600 522.000 466.600 ;
        RECT 526.400 461.600 527.200 467.000 ;
        RECT 529.200 461.600 530.000 464.200 ;
        RECT 532.400 461.600 533.200 464.200 ;
        RECT 535.600 461.600 536.400 464.200 ;
        RECT 538.800 461.600 539.800 465.600 ;
        RECT 545.000 462.200 546.000 465.600 ;
        RECT 545.000 461.600 545.800 462.200 ;
        RECT 548.400 461.600 549.200 464.200 ;
        RECT 551.600 461.600 552.400 464.200 ;
        RECT 554.800 461.600 555.600 464.200 ;
        RECT 558.000 462.200 559.000 465.600 ;
        RECT 558.200 461.600 559.000 462.200 ;
        RECT 564.200 461.600 565.200 465.600 ;
        RECT 569.200 462.200 570.200 465.600 ;
        RECT 569.400 461.600 570.200 462.200 ;
        RECT 575.400 461.600 576.400 465.600 ;
        RECT 578.800 461.600 579.600 464.200 ;
        RECT 585.200 461.600 586.000 466.200 ;
        RECT 596.400 461.600 597.200 464.200 ;
        RECT 599.600 461.600 600.400 464.200 ;
        RECT 609.200 461.600 610.000 466.200 ;
        RECT 0.400 460.400 614.000 461.600 ;
        RECT 2.800 456.000 3.600 460.400 ;
        RECT 8.400 457.800 9.200 460.400 ;
        RECT 11.600 457.800 12.600 460.400 ;
        RECT 17.200 455.800 18.000 460.400 ;
        RECT 22.000 456.600 22.800 460.400 ;
        RECT 28.000 455.000 28.800 460.400 ;
        RECT 33.200 455.400 34.000 460.400 ;
        RECT 36.400 457.800 37.200 460.400 ;
        RECT 39.600 455.800 40.400 460.400 ;
        RECT 42.800 455.800 43.600 460.400 ;
        RECT 49.200 456.600 50.000 460.400 ;
        RECT 54.000 455.800 54.800 460.400 ;
        RECT 59.400 457.800 60.400 460.400 ;
        RECT 62.800 457.800 63.600 460.400 ;
        RECT 68.400 456.000 69.200 460.400 ;
        RECT 73.200 455.400 74.000 460.400 ;
        RECT 78.400 455.000 79.200 460.400 ;
        RECT 82.800 456.600 83.600 460.400 ;
        RECT 90.800 456.600 91.600 460.400 ;
        RECT 94.000 455.800 94.800 460.400 ;
        RECT 97.200 455.800 98.000 460.400 ;
        RECT 102.000 456.600 102.800 460.400 ;
        RECT 106.800 453.800 107.600 460.400 ;
        RECT 113.200 453.800 114.000 460.400 ;
        RECT 120.800 455.000 121.600 460.400 ;
        RECT 126.000 455.400 126.800 460.400 ;
        RECT 129.200 457.800 130.000 460.400 ;
        RECT 134.000 456.600 134.800 460.400 ;
        RECT 140.400 456.600 141.200 460.400 ;
        RECT 145.200 455.800 146.000 460.400 ;
        RECT 156.000 455.000 156.800 460.400 ;
        RECT 161.200 455.400 162.000 460.400 ;
        RECT 169.200 453.800 170.000 460.400 ;
        RECT 172.400 456.600 173.200 460.400 ;
        RECT 178.800 456.000 179.600 460.400 ;
        RECT 184.400 457.800 185.200 460.400 ;
        RECT 187.600 457.800 188.600 460.400 ;
        RECT 193.200 455.800 194.000 460.400 ;
        RECT 196.400 453.800 197.200 460.400 ;
        RECT 202.800 457.800 203.600 460.400 ;
        RECT 209.200 455.800 210.000 460.400 ;
        RECT 210.800 455.800 211.600 460.400 ;
        RECT 214.000 455.800 214.800 460.400 ;
        RECT 217.200 455.800 218.000 460.400 ;
        RECT 220.400 455.800 221.200 460.400 ;
        RECT 223.600 455.800 224.400 460.400 ;
        RECT 228.400 455.800 229.200 460.400 ;
        RECT 231.600 455.800 232.400 460.400 ;
        RECT 234.800 455.800 235.600 460.400 ;
        RECT 236.400 457.800 237.200 460.400 ;
        RECT 242.800 455.800 243.600 460.400 ;
        RECT 254.000 457.800 254.800 460.400 ;
        RECT 257.200 457.800 258.000 460.400 ;
        RECT 266.800 455.800 267.600 460.400 ;
        RECT 273.200 456.200 274.000 460.400 ;
        RECT 276.400 457.800 277.200 460.400 ;
        RECT 279.600 455.800 280.400 460.400 ;
        RECT 282.800 455.800 283.600 460.400 ;
        RECT 286.000 456.600 286.800 460.400 ;
        RECT 295.600 457.800 296.400 460.400 ;
        RECT 302.000 455.800 302.800 460.400 ;
        RECT 313.200 457.800 314.000 460.400 ;
        RECT 316.400 457.800 317.200 460.400 ;
        RECT 326.000 455.800 326.800 460.400 ;
        RECT 332.400 456.000 333.200 460.400 ;
        RECT 338.000 457.800 338.800 460.400 ;
        RECT 341.200 457.800 342.200 460.400 ;
        RECT 346.800 455.800 347.600 460.400 ;
        RECT 350.000 457.800 350.800 460.400 ;
        RECT 354.800 455.800 355.600 460.400 ;
        RECT 358.000 455.800 358.800 460.400 ;
        RECT 361.200 456.600 362.000 460.400 ;
        RECT 367.600 455.400 368.400 460.400 ;
        RECT 372.800 455.000 373.600 460.400 ;
        RECT 377.200 455.400 378.000 460.400 ;
        RECT 382.400 455.000 383.200 460.400 ;
        RECT 386.800 456.600 387.600 460.400 ;
        RECT 393.200 455.800 394.000 460.400 ;
        RECT 398.600 457.800 399.600 460.400 ;
        RECT 402.000 457.800 402.800 460.400 ;
        RECT 407.600 456.000 408.400 460.400 ;
        RECT 414.000 456.600 414.800 460.400 ;
        RECT 420.400 456.600 421.200 460.400 ;
        RECT 426.800 456.600 427.600 460.400 ;
        RECT 431.600 456.600 432.400 460.400 ;
        RECT 438.000 456.600 438.800 460.400 ;
        RECT 442.800 453.800 443.600 460.400 ;
        RECT 449.200 453.800 450.000 460.400 ;
        RECT 455.600 457.800 456.400 460.400 ;
        RECT 465.200 456.600 466.000 460.400 ;
        RECT 471.600 456.600 472.400 460.400 ;
        RECT 479.600 456.600 480.400 460.400 ;
        RECT 484.400 455.400 485.200 460.400 ;
        RECT 489.600 455.000 490.400 460.400 ;
        RECT 495.600 456.600 496.400 460.400 ;
        RECT 500.400 456.600 501.200 460.400 ;
        RECT 505.200 457.800 506.000 460.400 ;
        RECT 508.400 457.800 509.200 460.400 ;
        RECT 514.800 453.800 515.600 460.400 ;
        RECT 519.600 456.600 520.400 460.400 ;
        RECT 522.800 457.800 523.600 460.400 ;
        RECT 529.200 456.600 530.000 460.400 ;
        RECT 534.000 455.800 534.800 460.400 ;
        RECT 537.200 455.800 538.000 460.400 ;
        RECT 538.800 457.800 539.600 460.400 ;
        RECT 545.200 455.800 546.000 460.400 ;
        RECT 556.400 457.800 557.200 460.400 ;
        RECT 559.600 457.800 560.400 460.400 ;
        RECT 569.200 455.800 570.000 460.400 ;
        RECT 574.000 457.800 574.800 460.400 ;
        RECT 580.400 455.800 581.200 460.400 ;
        RECT 591.600 457.800 592.400 460.400 ;
        RECT 594.800 457.800 595.600 460.400 ;
        RECT 604.400 455.800 605.200 460.400 ;
        RECT 1.200 421.600 2.000 424.200 ;
        RECT 6.000 421.600 6.800 425.400 ;
        RECT 10.800 421.600 11.600 426.200 ;
        RECT 14.000 421.600 14.800 426.200 ;
        RECT 17.200 421.600 18.000 426.200 ;
        RECT 20.400 421.600 21.200 426.200 ;
        RECT 23.600 421.600 24.400 426.200 ;
        RECT 28.400 421.600 29.200 425.400 ;
        RECT 31.600 421.600 32.400 424.200 ;
        RECT 34.800 421.600 35.600 425.800 ;
        RECT 38.000 421.600 38.800 426.200 ;
        RECT 41.200 421.600 42.000 426.200 ;
        RECT 44.400 421.600 45.200 426.200 ;
        RECT 47.600 421.600 48.400 426.200 ;
        RECT 50.800 421.600 51.600 426.200 ;
        RECT 54.000 421.600 54.800 426.200 ;
        RECT 59.400 421.600 60.400 424.200 ;
        RECT 62.800 421.600 63.600 424.200 ;
        RECT 68.400 421.600 69.200 426.000 ;
        RECT 73.200 421.600 74.000 426.600 ;
        RECT 78.400 421.600 79.200 427.000 ;
        RECT 82.800 421.600 83.600 425.400 ;
        RECT 90.800 421.600 91.600 425.400 ;
        RECT 94.000 421.600 94.800 426.200 ;
        RECT 100.400 421.600 101.200 426.600 ;
        RECT 105.600 421.600 106.400 427.000 ;
        RECT 110.000 421.600 110.800 425.400 ;
        RECT 118.000 421.600 118.800 425.400 ;
        RECT 121.200 421.600 122.000 424.200 ;
        RECT 126.000 421.600 126.800 425.400 ;
        RECT 130.800 421.600 131.600 424.200 ;
        RECT 135.600 421.600 136.400 426.000 ;
        RECT 141.200 421.600 142.000 424.200 ;
        RECT 144.400 421.600 145.400 424.200 ;
        RECT 150.000 421.600 150.800 426.200 ;
        RECT 159.600 421.600 160.400 425.400 ;
        RECT 167.600 421.600 168.400 425.400 ;
        RECT 172.400 421.600 173.200 425.400 ;
        RECT 180.400 421.600 181.200 425.400 ;
        RECT 185.200 421.600 186.000 426.000 ;
        RECT 190.800 421.600 191.600 424.200 ;
        RECT 194.000 421.600 195.000 424.200 ;
        RECT 199.600 421.600 200.400 426.200 ;
        RECT 204.400 421.600 205.200 425.400 ;
        RECT 210.800 421.600 211.600 425.400 ;
        RECT 218.800 421.600 219.600 426.200 ;
        RECT 223.600 421.600 224.400 425.400 ;
        RECT 229.000 421.600 229.800 426.000 ;
        RECT 233.200 421.600 234.000 426.200 ;
        RECT 238.000 421.600 238.800 426.200 ;
        RECT 246.000 421.600 246.800 425.400 ;
        RECT 250.800 421.600 251.600 424.200 ;
        RECT 255.600 421.600 256.400 425.400 ;
        RECT 260.400 421.600 261.200 426.600 ;
        RECT 265.600 421.600 266.400 427.000 ;
        RECT 270.000 421.600 270.800 426.600 ;
        RECT 275.200 421.600 276.000 427.000 ;
        RECT 281.200 421.600 282.000 426.200 ;
        RECT 282.800 421.600 283.600 424.200 ;
        RECT 286.000 421.600 286.800 424.200 ;
        RECT 292.400 421.600 293.200 426.200 ;
        RECT 303.600 421.600 304.400 424.200 ;
        RECT 306.800 421.600 307.600 424.200 ;
        RECT 316.400 421.600 317.200 426.200 ;
        RECT 326.000 421.600 326.800 424.200 ;
        RECT 330.800 421.600 331.600 426.200 ;
        RECT 336.200 421.600 337.200 424.200 ;
        RECT 339.600 421.600 340.400 424.200 ;
        RECT 345.200 421.600 346.000 426.000 ;
        RECT 350.000 421.600 350.800 426.600 ;
        RECT 355.200 421.600 356.000 427.000 ;
        RECT 359.600 421.600 360.400 425.400 ;
        RECT 367.600 421.600 368.400 425.400 ;
        RECT 372.000 421.600 372.800 427.000 ;
        RECT 377.200 421.600 378.000 426.600 ;
        RECT 382.000 421.600 382.800 425.400 ;
        RECT 388.000 421.600 388.800 427.000 ;
        RECT 393.200 421.600 394.000 426.600 ;
        RECT 396.400 421.600 397.200 424.200 ;
        RECT 400.800 421.600 401.600 427.000 ;
        RECT 406.000 421.600 406.800 426.600 ;
        RECT 410.800 421.600 411.600 425.400 ;
        RECT 417.200 421.600 418.000 426.000 ;
        RECT 422.800 421.600 423.600 424.200 ;
        RECT 426.000 421.600 427.000 424.200 ;
        RECT 431.600 421.600 432.400 426.200 ;
        RECT 434.800 421.600 435.600 424.200 ;
        RECT 439.600 421.600 440.400 425.400 ;
        RECT 446.000 421.600 446.800 426.200 ;
        RECT 451.400 421.600 452.400 424.200 ;
        RECT 454.800 421.600 455.600 424.200 ;
        RECT 460.400 421.600 461.200 426.000 ;
        RECT 473.200 421.600 474.000 428.200 ;
        RECT 474.800 421.600 475.600 424.200 ;
        RECT 481.200 421.600 482.000 426.200 ;
        RECT 492.400 421.600 493.200 424.200 ;
        RECT 495.600 421.600 496.400 424.200 ;
        RECT 505.200 421.600 506.000 426.200 ;
        RECT 510.000 421.600 510.800 424.200 ;
        RECT 516.400 421.600 517.200 426.200 ;
        RECT 527.600 421.600 528.400 424.200 ;
        RECT 530.800 421.600 531.600 424.200 ;
        RECT 540.400 421.600 541.200 426.200 ;
        RECT 546.800 421.600 547.600 426.600 ;
        RECT 552.000 421.600 552.800 427.000 ;
        RECT 556.400 421.600 557.200 426.600 ;
        RECT 561.600 421.600 562.400 427.000 ;
        RECT 564.400 421.600 565.200 424.200 ;
        RECT 570.800 421.600 571.600 426.200 ;
        RECT 582.000 421.600 582.800 424.200 ;
        RECT 585.200 421.600 586.000 424.200 ;
        RECT 594.800 421.600 595.600 426.200 ;
        RECT 599.600 421.600 600.400 426.200 ;
        RECT 602.800 421.600 603.600 426.200 ;
        RECT 606.000 421.600 606.800 426.200 ;
        RECT 609.200 421.600 610.000 426.200 ;
        RECT 612.400 421.600 613.200 426.200 ;
        RECT 0.400 420.400 614.000 421.600 ;
        RECT 4.400 415.800 5.200 420.400 ;
        RECT 14.000 417.800 14.800 420.400 ;
        RECT 17.200 417.800 18.000 420.400 ;
        RECT 28.400 415.800 29.200 420.400 ;
        RECT 34.800 417.800 35.600 420.400 ;
        RECT 39.600 416.600 40.400 420.400 ;
        RECT 44.400 416.600 45.200 420.400 ;
        RECT 50.800 415.400 51.600 420.400 ;
        RECT 56.000 415.000 56.800 420.400 ;
        RECT 62.000 416.600 62.800 420.400 ;
        RECT 66.800 415.800 67.600 420.400 ;
        RECT 72.200 417.800 73.200 420.400 ;
        RECT 75.600 417.800 76.400 420.400 ;
        RECT 81.200 416.000 82.000 420.400 ;
        RECT 86.000 416.600 86.800 420.400 ;
        RECT 94.000 416.600 94.800 420.400 ;
        RECT 97.200 415.800 98.000 420.400 ;
        RECT 103.600 416.600 104.400 420.400 ;
        RECT 108.400 415.800 109.200 420.400 ;
        RECT 111.600 415.800 112.400 420.400 ;
        RECT 114.800 415.800 115.600 420.400 ;
        RECT 118.000 415.800 118.800 420.400 ;
        RECT 122.800 415.800 123.600 420.400 ;
        RECT 126.000 415.800 126.800 420.400 ;
        RECT 127.600 417.800 128.400 420.400 ;
        RECT 132.400 416.600 133.200 420.400 ;
        RECT 138.800 415.400 139.600 420.400 ;
        RECT 144.000 415.000 144.800 420.400 ;
        RECT 146.800 415.800 147.600 420.400 ;
        RECT 158.000 416.600 158.800 420.400 ;
        RECT 164.400 416.600 165.200 420.400 ;
        RECT 170.800 415.800 171.600 420.400 ;
        RECT 174.000 415.800 174.800 420.400 ;
        RECT 177.200 416.600 178.000 420.400 ;
        RECT 185.200 415.800 186.000 420.400 ;
        RECT 194.800 417.800 195.600 420.400 ;
        RECT 198.000 417.800 198.800 420.400 ;
        RECT 209.200 415.800 210.000 420.400 ;
        RECT 215.600 417.800 216.400 420.400 ;
        RECT 217.200 417.800 218.000 420.400 ;
        RECT 220.400 417.800 221.200 420.400 ;
        RECT 223.600 417.800 224.400 420.400 ;
        RECT 225.200 417.800 226.000 420.400 ;
        RECT 229.400 415.800 230.200 420.400 ;
        RECT 236.400 413.800 237.200 420.400 ;
        RECT 238.000 417.800 238.800 420.400 ;
        RECT 241.200 416.200 242.000 420.400 ;
        RECT 244.400 417.800 245.200 420.400 ;
        RECT 247.600 417.800 248.400 420.400 ;
        RECT 251.000 419.800 251.800 420.400 ;
        RECT 250.800 416.400 251.800 419.800 ;
        RECT 257.000 416.400 258.000 420.400 ;
        RECT 263.600 416.600 264.400 420.400 ;
        RECT 268.600 419.800 269.400 420.400 ;
        RECT 268.400 416.400 269.400 419.800 ;
        RECT 274.600 416.400 275.600 420.400 ;
        RECT 279.600 416.600 280.400 420.400 ;
        RECT 286.000 416.600 286.800 420.400 ;
        RECT 290.800 415.800 291.600 420.400 ;
        RECT 303.600 415.800 304.400 420.400 ;
        RECT 313.200 417.800 314.000 420.400 ;
        RECT 316.400 417.800 317.200 420.400 ;
        RECT 327.600 415.800 328.400 420.400 ;
        RECT 334.000 417.800 334.800 420.400 ;
        RECT 337.200 415.800 338.000 420.400 ;
        RECT 342.600 417.800 343.600 420.400 ;
        RECT 346.000 417.800 346.800 420.400 ;
        RECT 351.600 416.000 352.400 420.400 ;
        RECT 356.400 416.600 357.200 420.400 ;
        RECT 364.400 416.600 365.200 420.400 ;
        RECT 367.600 417.800 368.400 420.400 ;
        RECT 372.400 416.600 373.200 420.400 ;
        RECT 380.400 416.600 381.200 420.400 ;
        RECT 383.600 417.800 384.400 420.400 ;
        RECT 388.400 416.600 389.200 420.400 ;
        RECT 393.200 413.800 394.000 420.400 ;
        RECT 399.600 413.800 400.400 420.400 ;
        RECT 407.600 416.600 408.400 420.400 ;
        RECT 412.400 417.800 413.200 420.400 ;
        RECT 417.200 416.600 418.000 420.400 ;
        RECT 423.600 416.600 424.400 420.400 ;
        RECT 430.000 416.600 430.800 420.400 ;
        RECT 434.800 415.800 435.600 420.400 ;
        RECT 441.200 417.800 442.000 420.400 ;
        RECT 444.400 416.600 445.200 420.400 ;
        RECT 449.200 415.800 450.000 420.400 ;
        RECT 454.000 415.800 454.800 420.400 ;
        RECT 465.200 416.600 466.000 420.400 ;
        RECT 471.600 416.600 472.400 420.400 ;
        RECT 476.400 416.400 477.400 420.400 ;
        RECT 482.600 419.800 483.400 420.400 ;
        RECT 482.600 416.400 483.600 419.800 ;
        RECT 489.200 416.600 490.000 420.400 ;
        RECT 494.600 416.000 495.400 420.400 ;
        RECT 498.800 417.800 499.600 420.400 ;
        RECT 503.000 415.800 503.800 420.400 ;
        RECT 505.200 415.800 506.000 420.400 ;
        RECT 510.000 415.800 510.800 420.400 ;
        RECT 514.800 413.800 515.600 420.400 ;
        RECT 521.200 417.800 522.000 420.400 ;
        RECT 524.400 417.800 525.200 420.400 ;
        RECT 527.600 417.800 528.400 420.400 ;
        RECT 530.800 416.200 531.600 420.400 ;
        RECT 534.000 417.800 534.800 420.400 ;
        RECT 537.400 419.800 538.200 420.400 ;
        RECT 537.200 416.400 538.200 419.800 ;
        RECT 543.400 416.400 544.400 420.400 ;
        RECT 548.400 416.600 549.200 420.400 ;
        RECT 554.800 416.600 555.600 420.400 ;
        RECT 561.400 419.800 562.200 420.400 ;
        RECT 561.200 416.400 562.200 419.800 ;
        RECT 567.400 416.400 568.400 420.400 ;
        RECT 570.800 415.800 571.600 420.400 ;
        RECT 578.800 415.800 579.600 420.400 ;
        RECT 588.400 417.800 589.200 420.400 ;
        RECT 591.600 417.800 592.400 420.400 ;
        RECT 602.800 415.800 603.600 420.400 ;
        RECT 609.200 417.800 610.000 420.400 ;
        RECT 4.400 381.600 5.200 386.200 ;
        RECT 14.000 381.600 14.800 384.200 ;
        RECT 17.200 381.600 18.000 384.200 ;
        RECT 28.400 381.600 29.200 386.200 ;
        RECT 34.800 381.600 35.600 384.200 ;
        RECT 39.600 381.600 40.400 386.200 ;
        RECT 41.200 381.600 42.000 386.200 ;
        RECT 44.400 381.600 45.200 386.200 ;
        RECT 49.200 381.600 50.000 386.200 ;
        RECT 54.600 381.600 55.600 384.200 ;
        RECT 58.000 381.600 58.800 384.200 ;
        RECT 63.600 381.600 64.400 386.000 ;
        RECT 68.400 381.600 69.200 386.200 ;
        RECT 71.600 381.600 72.400 386.200 ;
        RECT 76.400 381.600 77.200 385.400 ;
        RECT 80.800 381.600 81.600 387.000 ;
        RECT 86.000 381.600 86.800 386.600 ;
        RECT 90.400 381.600 91.200 387.000 ;
        RECT 95.600 381.600 96.400 386.600 ;
        RECT 100.400 381.600 101.200 384.200 ;
        RECT 102.000 381.600 102.800 386.200 ;
        RECT 105.200 381.600 106.000 386.200 ;
        RECT 108.400 381.600 109.200 384.200 ;
        RECT 111.600 381.600 112.400 384.200 ;
        RECT 114.800 381.600 115.600 386.200 ;
        RECT 120.200 381.600 121.200 384.200 ;
        RECT 123.600 381.600 124.400 384.200 ;
        RECT 129.200 381.600 130.000 386.000 ;
        RECT 134.000 381.600 134.800 385.400 ;
        RECT 142.000 381.600 142.800 385.400 ;
        RECT 145.200 381.600 146.000 386.200 ;
        RECT 148.400 381.600 149.200 386.200 ;
        RECT 156.400 381.600 157.200 384.200 ;
        RECT 159.600 381.600 160.400 386.200 ;
        RECT 162.800 381.600 163.600 386.200 ;
        RECT 166.000 381.600 166.800 384.200 ;
        RECT 172.400 381.600 173.200 386.200 ;
        RECT 183.600 381.600 184.400 384.200 ;
        RECT 186.800 381.600 187.600 384.200 ;
        RECT 196.400 381.600 197.200 386.200 ;
        RECT 201.200 381.600 202.000 384.200 ;
        RECT 207.600 381.600 208.400 386.200 ;
        RECT 212.400 381.600 213.200 386.200 ;
        RECT 217.200 381.600 218.000 386.200 ;
        RECT 226.800 381.600 227.600 384.200 ;
        RECT 230.000 381.600 230.800 384.200 ;
        RECT 241.200 381.600 242.000 386.200 ;
        RECT 247.600 381.600 248.400 384.200 ;
        RECT 249.200 381.600 250.000 386.200 ;
        RECT 257.200 381.600 258.000 385.400 ;
        RECT 262.000 381.600 262.800 386.200 ;
        RECT 268.400 381.600 269.200 386.200 ;
        RECT 278.000 381.600 278.800 384.200 ;
        RECT 281.200 381.600 282.000 384.200 ;
        RECT 292.400 381.600 293.200 386.200 ;
        RECT 298.800 381.600 299.600 384.200 ;
        RECT 308.400 381.600 309.200 386.200 ;
        RECT 318.000 381.600 318.800 384.200 ;
        RECT 321.200 381.600 322.000 384.200 ;
        RECT 332.400 381.600 333.200 386.200 ;
        RECT 338.800 381.600 339.600 384.200 ;
        RECT 340.400 381.600 341.200 384.200 ;
        RECT 346.800 381.600 347.600 386.200 ;
        RECT 358.000 381.600 358.800 384.200 ;
        RECT 361.200 381.600 362.000 384.200 ;
        RECT 370.800 381.600 371.600 386.200 ;
        RECT 377.200 381.600 378.000 386.200 ;
        RECT 382.600 381.600 383.600 384.200 ;
        RECT 386.000 381.600 386.800 384.200 ;
        RECT 391.600 381.600 392.400 386.000 ;
        RECT 394.800 381.600 395.600 384.200 ;
        RECT 398.000 381.600 398.800 384.200 ;
        RECT 402.800 381.600 403.600 386.200 ;
        RECT 406.000 381.600 406.800 386.200 ;
        RECT 407.600 381.600 408.400 384.200 ;
        RECT 414.000 381.600 414.800 386.200 ;
        RECT 425.200 381.600 426.000 384.200 ;
        RECT 428.400 381.600 429.200 384.200 ;
        RECT 438.000 381.600 438.800 386.200 ;
        RECT 446.000 381.600 446.800 386.200 ;
        RECT 450.800 381.600 451.600 385.400 ;
        RECT 462.000 381.600 462.800 386.200 ;
        RECT 471.600 381.600 472.400 384.200 ;
        RECT 474.800 381.600 475.600 384.200 ;
        RECT 486.000 381.600 486.800 386.200 ;
        RECT 492.400 381.600 493.200 384.200 ;
        RECT 494.000 381.600 494.800 386.200 ;
        RECT 497.200 381.600 498.000 386.200 ;
        RECT 500.400 381.600 501.200 386.200 ;
        RECT 503.600 381.600 504.400 386.200 ;
        RECT 506.800 381.600 507.600 386.200 ;
        RECT 508.400 381.600 509.200 384.200 ;
        RECT 511.600 381.600 512.400 384.200 ;
        RECT 516.400 381.600 517.200 386.200 ;
        RECT 521.200 381.600 522.000 386.200 ;
        RECT 530.800 381.600 531.600 384.200 ;
        RECT 534.000 381.600 534.800 384.200 ;
        RECT 545.200 381.600 546.000 386.200 ;
        RECT 551.600 381.600 552.400 384.200 ;
        RECT 553.200 381.600 554.000 384.200 ;
        RECT 556.400 381.600 557.200 384.200 ;
        RECT 561.200 381.600 562.000 385.400 ;
        RECT 566.000 381.600 566.800 384.200 ;
        RECT 569.200 381.600 570.000 385.800 ;
        RECT 572.400 381.600 573.200 384.200 ;
        RECT 577.200 381.600 578.000 386.200 ;
        RECT 586.800 381.600 587.600 384.200 ;
        RECT 590.000 381.600 590.800 384.200 ;
        RECT 601.200 381.600 602.000 386.200 ;
        RECT 607.600 381.600 608.400 384.200 ;
        RECT 0.400 380.400 614.000 381.600 ;
        RECT 1.200 377.800 2.000 380.400 ;
        RECT 4.400 377.800 5.200 380.400 ;
        RECT 9.200 376.600 10.000 380.400 ;
        RECT 15.600 376.600 16.400 380.400 ;
        RECT 23.600 376.600 24.400 380.400 ;
        RECT 28.400 376.600 29.200 380.400 ;
        RECT 36.400 376.600 37.200 380.400 ;
        RECT 42.800 376.600 43.600 380.400 ;
        RECT 49.200 375.800 50.000 380.400 ;
        RECT 54.000 376.600 54.800 380.400 ;
        RECT 58.800 375.400 59.600 380.400 ;
        RECT 64.000 375.000 64.800 380.400 ;
        RECT 68.400 376.600 69.200 380.400 ;
        RECT 76.400 376.600 77.200 380.400 ;
        RECT 81.200 376.600 82.000 380.400 ;
        RECT 89.200 376.600 90.000 380.400 ;
        RECT 94.000 376.000 94.800 380.400 ;
        RECT 99.600 377.800 100.400 380.400 ;
        RECT 102.800 377.800 103.800 380.400 ;
        RECT 108.400 375.800 109.200 380.400 ;
        RECT 111.600 377.800 112.400 380.400 ;
        RECT 118.000 376.600 118.800 380.400 ;
        RECT 122.800 376.600 123.600 380.400 ;
        RECT 129.200 375.400 130.000 380.400 ;
        RECT 134.400 375.000 135.200 380.400 ;
        RECT 138.800 376.600 139.600 380.400 ;
        RECT 145.200 376.600 146.000 380.400 ;
        RECT 156.400 375.800 157.200 380.400 ;
        RECT 161.800 377.800 162.800 380.400 ;
        RECT 165.200 377.800 166.000 380.400 ;
        RECT 170.800 376.000 171.600 380.400 ;
        RECT 177.200 375.800 178.000 380.400 ;
        RECT 186.800 377.800 187.600 380.400 ;
        RECT 190.000 377.800 190.800 380.400 ;
        RECT 201.200 375.800 202.000 380.400 ;
        RECT 207.600 377.800 208.400 380.400 ;
        RECT 212.400 375.800 213.200 380.400 ;
        RECT 217.200 376.600 218.000 380.400 ;
        RECT 223.600 376.600 224.400 380.400 ;
        RECT 228.400 376.600 229.200 380.400 ;
        RECT 233.200 377.800 234.000 380.400 ;
        RECT 239.600 375.800 240.400 380.400 ;
        RECT 250.800 377.800 251.600 380.400 ;
        RECT 254.000 377.800 254.800 380.400 ;
        RECT 263.600 375.800 264.400 380.400 ;
        RECT 268.400 375.800 269.200 380.400 ;
        RECT 271.600 375.800 272.400 380.400 ;
        RECT 274.800 375.800 275.600 380.400 ;
        RECT 278.000 375.800 278.800 380.400 ;
        RECT 281.200 375.800 282.000 380.400 ;
        RECT 284.400 375.800 285.200 380.400 ;
        RECT 287.600 375.800 288.400 380.400 ;
        RECT 289.200 375.800 290.000 380.400 ;
        RECT 292.400 375.800 293.200 380.400 ;
        RECT 295.600 375.800 296.400 380.400 ;
        RECT 298.800 375.800 299.600 380.400 ;
        RECT 302.000 375.800 302.800 380.400 ;
        RECT 310.000 375.400 310.800 380.400 ;
        RECT 315.200 375.000 316.000 380.400 ;
        RECT 319.600 377.800 320.400 380.400 ;
        RECT 324.400 376.600 325.200 380.400 ;
        RECT 329.200 377.800 330.000 380.400 ;
        RECT 332.400 375.400 333.200 380.400 ;
        RECT 337.600 375.000 338.400 380.400 ;
        RECT 342.000 377.800 342.800 380.400 ;
        RECT 346.800 375.800 347.600 380.400 ;
        RECT 356.400 377.800 357.200 380.400 ;
        RECT 359.600 377.800 360.400 380.400 ;
        RECT 370.800 375.800 371.600 380.400 ;
        RECT 377.200 377.800 378.000 380.400 ;
        RECT 378.800 377.800 379.600 380.400 ;
        RECT 385.200 375.800 386.000 380.400 ;
        RECT 396.400 377.800 397.200 380.400 ;
        RECT 399.600 377.800 400.400 380.400 ;
        RECT 409.200 375.800 410.000 380.400 ;
        RECT 415.600 375.800 416.400 380.400 ;
        RECT 418.800 375.800 419.600 380.400 ;
        RECT 423.600 375.800 424.400 380.400 ;
        RECT 428.400 376.600 429.200 380.400 ;
        RECT 433.200 376.600 434.000 380.400 ;
        RECT 438.000 375.800 438.800 380.400 ;
        RECT 447.600 377.800 448.400 380.400 ;
        RECT 454.000 375.800 454.800 380.400 ;
        RECT 465.200 377.800 466.000 380.400 ;
        RECT 468.400 377.800 469.200 380.400 ;
        RECT 478.000 375.800 478.800 380.400 ;
        RECT 484.400 377.800 485.200 380.400 ;
        RECT 486.000 375.800 486.800 380.400 ;
        RECT 489.200 375.800 490.000 380.400 ;
        RECT 492.400 375.800 493.200 380.400 ;
        RECT 495.600 375.800 496.400 380.400 ;
        RECT 498.800 375.800 499.600 380.400 ;
        RECT 500.400 375.800 501.200 380.400 ;
        RECT 503.600 375.800 504.400 380.400 ;
        RECT 506.800 375.800 507.600 380.400 ;
        RECT 510.000 375.800 510.800 380.400 ;
        RECT 513.200 375.800 514.000 380.400 ;
        RECT 516.400 375.800 517.200 380.400 ;
        RECT 519.600 377.800 520.400 380.400 ;
        RECT 526.000 375.800 526.800 380.400 ;
        RECT 537.200 377.800 538.000 380.400 ;
        RECT 540.400 377.800 541.200 380.400 ;
        RECT 550.000 375.800 550.800 380.400 ;
        RECT 556.400 375.800 557.200 380.400 ;
        RECT 559.600 375.800 560.400 380.400 ;
        RECT 564.400 375.800 565.200 380.400 ;
        RECT 567.600 376.600 568.400 380.400 ;
        RECT 572.400 377.800 573.200 380.400 ;
        RECT 578.800 375.800 579.600 380.400 ;
        RECT 590.000 377.800 590.800 380.400 ;
        RECT 593.200 377.800 594.000 380.400 ;
        RECT 602.800 375.800 603.600 380.400 ;
        RECT 609.200 375.800 610.000 380.400 ;
        RECT 1.200 341.600 2.000 344.200 ;
        RECT 6.000 341.600 6.800 345.400 ;
        RECT 14.000 341.600 14.800 346.200 ;
        RECT 23.600 341.600 24.400 344.200 ;
        RECT 26.800 341.600 27.600 344.200 ;
        RECT 38.000 341.600 38.800 346.200 ;
        RECT 44.400 341.600 45.200 344.200 ;
        RECT 46.000 341.600 46.800 344.200 ;
        RECT 50.800 341.600 51.600 344.200 ;
        RECT 55.600 341.600 56.400 346.200 ;
        RECT 58.800 341.600 59.600 344.200 ;
        RECT 62.000 341.600 62.800 346.200 ;
        RECT 67.400 341.600 68.400 344.200 ;
        RECT 70.800 341.600 71.600 344.200 ;
        RECT 76.400 341.600 77.200 346.000 ;
        RECT 81.200 341.600 82.000 344.200 ;
        RECT 86.000 341.600 86.800 346.200 ;
        RECT 90.800 341.600 91.600 345.400 ;
        RECT 97.200 341.600 98.000 345.400 ;
        RECT 102.000 341.600 102.800 344.200 ;
        RECT 105.200 341.600 106.000 346.600 ;
        RECT 110.400 341.600 111.200 347.000 ;
        RECT 114.800 341.600 115.600 345.400 ;
        RECT 122.800 341.600 123.600 345.400 ;
        RECT 129.200 341.600 130.000 345.400 ;
        RECT 134.000 341.600 134.800 346.600 ;
        RECT 139.200 341.600 140.000 347.000 ;
        RECT 142.000 341.600 142.800 346.200 ;
        RECT 145.200 341.600 146.000 346.200 ;
        RECT 148.400 341.600 149.200 346.200 ;
        RECT 151.600 341.600 152.400 346.200 ;
        RECT 154.800 341.600 155.600 346.200 ;
        RECT 161.200 341.600 162.000 344.200 ;
        RECT 165.600 341.600 166.400 347.000 ;
        RECT 170.800 341.600 171.600 346.600 ;
        RECT 175.600 341.600 176.400 346.200 ;
        RECT 182.000 341.600 182.800 346.200 ;
        RECT 191.600 341.600 192.400 344.200 ;
        RECT 194.800 341.600 195.600 344.200 ;
        RECT 206.000 341.600 206.800 346.200 ;
        RECT 212.400 341.600 213.200 344.200 ;
        RECT 214.000 341.600 214.800 346.200 ;
        RECT 217.200 341.600 218.000 346.200 ;
        RECT 220.400 341.600 221.200 346.200 ;
        RECT 223.600 341.600 224.400 346.200 ;
        RECT 226.800 341.600 227.600 346.200 ;
        RECT 230.000 341.600 230.800 346.200 ;
        RECT 233.200 341.600 234.000 346.200 ;
        RECT 238.000 341.600 238.800 346.200 ;
        RECT 247.600 341.600 248.400 344.200 ;
        RECT 250.800 341.600 251.600 344.200 ;
        RECT 262.000 341.600 262.800 346.200 ;
        RECT 268.400 341.600 269.200 344.200 ;
        RECT 271.600 341.600 272.400 346.600 ;
        RECT 276.800 341.600 277.600 347.000 ;
        RECT 281.200 341.600 282.000 344.200 ;
        RECT 282.800 341.600 283.600 344.200 ;
        RECT 289.200 341.600 290.000 346.200 ;
        RECT 298.800 341.600 299.600 344.200 ;
        RECT 302.000 341.600 302.800 344.200 ;
        RECT 313.200 341.600 314.000 346.200 ;
        RECT 319.600 341.600 320.400 344.200 ;
        RECT 327.600 341.600 328.400 346.600 ;
        RECT 332.800 341.600 333.600 347.000 ;
        RECT 337.200 341.600 338.000 344.200 ;
        RECT 342.000 341.600 342.800 346.200 ;
        RECT 351.600 341.600 352.400 344.200 ;
        RECT 354.800 341.600 355.600 344.200 ;
        RECT 366.000 341.600 366.800 346.200 ;
        RECT 372.400 341.600 373.200 344.200 ;
        RECT 374.000 341.600 374.800 344.200 ;
        RECT 377.200 341.600 378.000 346.200 ;
        RECT 383.200 341.600 384.000 347.000 ;
        RECT 388.400 341.600 389.200 346.600 ;
        RECT 392.800 341.600 393.600 347.000 ;
        RECT 398.000 341.600 398.800 346.600 ;
        RECT 404.400 341.600 405.200 346.200 ;
        RECT 407.600 341.600 408.400 344.200 ;
        RECT 409.200 341.600 410.000 346.200 ;
        RECT 414.000 341.600 414.800 344.200 ;
        RECT 420.400 341.600 421.200 346.200 ;
        RECT 431.600 341.600 432.400 344.200 ;
        RECT 434.800 341.600 435.600 344.200 ;
        RECT 444.400 341.600 445.200 346.200 ;
        RECT 449.200 341.600 450.000 344.200 ;
        RECT 452.400 341.600 453.200 344.200 ;
        RECT 458.800 341.600 459.600 344.200 ;
        RECT 465.200 341.600 466.000 346.200 ;
        RECT 476.400 341.600 477.200 344.200 ;
        RECT 479.600 341.600 480.400 344.200 ;
        RECT 489.200 341.600 490.000 346.200 ;
        RECT 497.200 341.600 498.000 346.200 ;
        RECT 506.800 341.600 507.600 344.200 ;
        RECT 510.000 341.600 510.800 344.200 ;
        RECT 521.200 341.600 522.000 346.200 ;
        RECT 527.600 341.600 528.400 344.200 ;
        RECT 529.200 341.600 530.000 346.200 ;
        RECT 534.000 341.600 534.800 346.200 ;
        RECT 537.200 341.600 538.000 346.200 ;
        RECT 542.000 341.600 542.800 346.200 ;
        RECT 545.200 341.600 546.000 346.200 ;
        RECT 546.800 341.600 547.600 346.200 ;
        RECT 550.000 341.600 550.800 346.200 ;
        RECT 553.200 341.600 554.000 346.200 ;
        RECT 558.000 341.600 558.800 346.200 ;
        RECT 561.200 341.600 562.000 345.400 ;
        RECT 569.200 341.600 570.000 346.200 ;
        RECT 578.800 341.600 579.600 344.200 ;
        RECT 582.000 341.600 582.800 344.200 ;
        RECT 593.200 341.600 594.000 346.200 ;
        RECT 599.600 341.600 600.400 344.200 ;
        RECT 601.200 341.600 602.000 346.200 ;
        RECT 607.600 341.600 608.400 346.200 ;
        RECT 0.400 340.400 614.000 341.600 ;
        RECT 4.400 335.800 5.200 340.400 ;
        RECT 14.000 337.800 14.800 340.400 ;
        RECT 17.200 337.800 18.000 340.400 ;
        RECT 28.400 335.800 29.200 340.400 ;
        RECT 34.800 337.800 35.600 340.400 ;
        RECT 36.400 335.800 37.200 340.400 ;
        RECT 39.600 335.800 40.400 340.400 ;
        RECT 44.400 337.800 45.200 340.400 ;
        RECT 47.200 335.000 48.000 340.400 ;
        RECT 52.400 335.400 53.200 340.400 ;
        RECT 55.600 337.800 56.400 340.400 ;
        RECT 58.800 337.800 59.600 340.400 ;
        RECT 65.200 335.800 66.000 340.400 ;
        RECT 76.400 337.800 77.200 340.400 ;
        RECT 79.600 337.800 80.400 340.400 ;
        RECT 89.200 335.800 90.000 340.400 ;
        RECT 94.000 337.800 94.800 340.400 ;
        RECT 98.400 335.000 99.200 340.400 ;
        RECT 103.600 335.400 104.400 340.400 ;
        RECT 108.400 335.800 109.200 340.400 ;
        RECT 113.800 337.800 114.800 340.400 ;
        RECT 117.200 337.800 118.000 340.400 ;
        RECT 122.800 336.000 123.600 340.400 ;
        RECT 127.600 335.800 128.400 340.400 ;
        RECT 133.000 337.800 134.000 340.400 ;
        RECT 136.400 337.800 137.200 340.400 ;
        RECT 142.000 336.000 142.800 340.400 ;
        RECT 146.800 337.800 147.600 340.400 ;
        RECT 153.200 337.800 154.000 340.400 ;
        RECT 159.600 335.800 160.400 340.400 ;
        RECT 170.800 337.800 171.600 340.400 ;
        RECT 174.000 337.800 174.800 340.400 ;
        RECT 183.600 335.800 184.400 340.400 ;
        RECT 190.000 335.800 190.800 340.400 ;
        RECT 193.200 335.800 194.000 340.400 ;
        RECT 198.000 335.800 198.800 340.400 ;
        RECT 207.600 337.800 208.400 340.400 ;
        RECT 210.800 337.800 211.600 340.400 ;
        RECT 222.000 335.800 222.800 340.400 ;
        RECT 228.400 337.800 229.200 340.400 ;
        RECT 230.000 335.800 230.800 340.400 ;
        RECT 233.200 335.800 234.000 340.400 ;
        RECT 236.400 335.800 237.200 340.400 ;
        RECT 238.000 337.800 238.800 340.400 ;
        RECT 244.400 335.800 245.200 340.400 ;
        RECT 254.000 337.800 254.800 340.400 ;
        RECT 257.200 337.800 258.000 340.400 ;
        RECT 268.400 335.800 269.200 340.400 ;
        RECT 274.800 337.800 275.600 340.400 ;
        RECT 278.000 337.800 278.800 340.400 ;
        RECT 284.400 334.300 285.200 340.400 ;
        RECT 290.800 334.300 291.600 340.400 ;
        RECT 297.200 334.300 298.000 340.400 ;
        RECT 303.600 334.300 304.400 340.400 ;
        RECT 310.000 335.800 310.800 340.400 ;
        RECT 313.200 335.800 314.000 340.400 ;
        RECT 316.400 335.800 317.200 340.400 ;
        RECT 322.800 336.600 323.600 340.400 ;
        RECT 332.400 336.600 333.200 340.400 ;
        RECT 335.600 337.800 336.400 340.400 ;
        RECT 342.000 335.800 342.800 340.400 ;
        RECT 353.200 337.800 354.000 340.400 ;
        RECT 356.400 337.800 357.200 340.400 ;
        RECT 366.000 335.800 366.800 340.400 ;
        RECT 374.000 336.600 374.800 340.400 ;
        RECT 382.000 336.600 382.800 340.400 ;
        RECT 388.400 335.800 389.200 340.400 ;
        RECT 390.000 335.800 390.800 340.400 ;
        RECT 393.200 335.800 394.000 340.400 ;
        RECT 396.400 337.800 397.200 340.400 ;
        RECT 402.800 335.800 403.600 340.400 ;
        RECT 414.000 337.800 414.800 340.400 ;
        RECT 417.200 337.800 418.000 340.400 ;
        RECT 426.800 335.800 427.600 340.400 ;
        RECT 434.800 335.800 435.600 340.400 ;
        RECT 436.400 337.800 437.200 340.400 ;
        RECT 441.200 336.600 442.000 340.400 ;
        RECT 447.600 336.600 448.400 340.400 ;
        RECT 452.400 335.800 453.200 340.400 ;
        RECT 462.600 335.800 463.400 340.400 ;
        RECT 466.800 337.800 467.600 340.400 ;
        RECT 468.400 337.800 469.200 340.400 ;
        RECT 471.600 337.800 472.400 340.400 ;
        RECT 473.200 337.800 474.000 340.400 ;
        RECT 476.400 337.800 477.200 340.400 ;
        RECT 481.200 336.600 482.000 340.400 ;
        RECT 484.400 335.800 485.200 340.400 ;
        RECT 489.200 335.800 490.000 340.400 ;
        RECT 492.400 335.800 493.200 340.400 ;
        RECT 282.900 333.800 285.200 334.300 ;
        RECT 289.300 333.800 291.600 334.300 ;
        RECT 295.700 333.800 298.000 334.300 ;
        RECT 302.100 333.800 304.400 334.300 ;
        RECT 388.400 334.300 389.200 335.200 ;
        RECT 390.100 334.300 390.700 335.800 ;
        RECT 282.900 333.700 285.100 333.800 ;
        RECT 289.300 333.700 291.500 333.800 ;
        RECT 295.700 333.700 297.900 333.800 ;
        RECT 302.100 333.700 304.300 333.800 ;
        RECT 388.400 333.700 390.700 334.300 ;
        RECT 494.000 333.800 494.800 340.400 ;
        RECT 500.400 337.800 501.200 340.400 ;
        RECT 503.600 337.800 504.400 340.400 ;
        RECT 505.200 337.800 506.000 340.400 ;
        RECT 511.600 335.800 512.400 340.400 ;
        RECT 522.800 337.800 523.600 340.400 ;
        RECT 526.000 337.800 526.800 340.400 ;
        RECT 535.600 335.800 536.400 340.400 ;
        RECT 543.600 335.800 544.400 340.400 ;
        RECT 553.200 337.800 554.000 340.400 ;
        RECT 556.400 337.800 557.200 340.400 ;
        RECT 567.600 335.800 568.400 340.400 ;
        RECT 574.000 337.800 574.800 340.400 ;
        RECT 578.800 335.800 579.600 340.400 ;
        RECT 583.600 336.600 584.400 340.400 ;
        RECT 588.400 337.800 589.200 340.400 ;
        RECT 590.000 335.800 590.800 340.400 ;
        RECT 598.000 336.600 598.800 340.400 ;
        RECT 602.800 337.800 603.600 340.400 ;
        RECT 604.400 335.800 605.200 340.400 ;
        RECT 607.600 335.800 608.400 340.400 ;
        RECT 610.800 335.800 611.600 340.400 ;
        RECT 282.900 332.400 283.500 333.700 ;
        RECT 289.300 332.400 289.900 333.700 ;
        RECT 295.700 332.400 296.300 333.700 ;
        RECT 302.100 332.400 302.700 333.700 ;
        RECT 388.400 333.600 389.200 333.700 ;
        RECT 282.000 331.600 283.600 332.400 ;
        RECT 288.400 331.600 290.000 332.400 ;
        RECT 294.800 331.600 296.400 332.400 ;
        RECT 301.200 331.600 302.800 332.400 ;
        RECT 319.600 328.800 320.400 330.400 ;
        RECT 198.000 311.600 198.800 314.400 ;
        RECT 358.000 310.800 358.800 312.400 ;
        RECT 369.200 310.800 370.000 312.400 ;
        RECT 358.100 308.200 358.700 310.800 ;
        RECT 367.600 308.300 368.400 308.400 ;
        RECT 369.300 308.300 369.900 310.800 ;
        RECT 367.600 308.200 369.900 308.300 ;
        RECT 1.200 301.600 2.000 306.200 ;
        RECT 4.400 301.600 5.200 306.200 ;
        RECT 7.600 301.600 8.400 306.200 ;
        RECT 10.800 301.600 11.600 306.200 ;
        RECT 14.000 301.600 14.800 306.200 ;
        RECT 18.800 301.600 19.600 306.200 ;
        RECT 28.400 301.600 29.200 304.200 ;
        RECT 31.600 301.600 32.400 304.200 ;
        RECT 42.800 301.600 43.600 306.200 ;
        RECT 49.200 301.600 50.000 304.200 ;
        RECT 50.800 301.600 51.600 304.200 ;
        RECT 57.200 301.600 58.000 306.200 ;
        RECT 68.400 301.600 69.200 304.200 ;
        RECT 71.600 301.600 72.400 304.200 ;
        RECT 81.200 301.600 82.000 306.200 ;
        RECT 87.200 301.600 88.000 307.000 ;
        RECT 92.400 301.600 93.200 306.600 ;
        RECT 97.200 301.600 98.000 306.600 ;
        RECT 102.400 301.600 103.200 307.000 ;
        RECT 106.800 301.600 107.600 304.200 ;
        RECT 108.400 301.600 109.200 304.200 ;
        RECT 114.800 301.600 115.600 306.200 ;
        RECT 126.000 301.600 126.800 304.200 ;
        RECT 129.200 301.600 130.000 304.200 ;
        RECT 138.800 301.600 139.600 306.200 ;
        RECT 143.600 301.600 144.400 304.200 ;
        RECT 146.800 301.600 147.600 304.200 ;
        RECT 153.200 301.600 154.000 304.200 ;
        RECT 157.400 301.600 158.200 306.200 ;
        RECT 159.600 301.600 160.400 304.200 ;
        RECT 166.000 301.600 166.800 306.200 ;
        RECT 177.200 301.600 178.000 304.200 ;
        RECT 180.400 301.600 181.200 304.200 ;
        RECT 190.000 301.600 190.800 306.200 ;
        RECT 194.800 301.600 195.600 308.200 ;
        RECT 204.400 301.600 205.200 306.200 ;
        RECT 214.000 301.600 214.800 304.200 ;
        RECT 217.200 301.600 218.000 304.200 ;
        RECT 228.400 301.600 229.200 306.200 ;
        RECT 234.800 301.600 235.600 304.200 ;
        RECT 238.000 301.600 238.800 306.200 ;
        RECT 239.600 301.600 240.400 306.200 ;
        RECT 244.400 301.600 245.200 306.200 ;
        RECT 250.800 301.600 251.600 306.200 ;
        RECT 254.000 301.600 254.800 306.200 ;
        RECT 256.800 301.600 257.600 307.000 ;
        RECT 262.000 301.600 262.800 306.600 ;
        RECT 266.800 301.600 267.600 306.600 ;
        RECT 272.000 301.600 272.800 307.000 ;
        RECT 278.000 301.600 278.800 305.400 ;
        RECT 281.200 301.600 282.000 306.200 ;
        RECT 287.600 301.600 288.400 306.200 ;
        RECT 290.800 301.600 291.600 306.200 ;
        RECT 297.200 301.600 298.000 304.200 ;
        RECT 303.600 301.600 304.400 306.200 ;
        RECT 314.800 301.600 315.600 304.200 ;
        RECT 318.000 301.600 318.800 304.200 ;
        RECT 327.600 301.600 328.400 306.200 ;
        RECT 332.400 301.600 333.200 306.200 ;
        RECT 337.200 301.600 338.000 306.200 ;
        RECT 345.200 301.600 346.000 305.400 ;
        RECT 351.600 301.600 352.400 305.400 ;
        RECT 356.400 301.600 357.200 304.200 ;
        RECT 358.000 301.600 358.800 308.200 ;
        RECT 367.600 307.700 370.000 308.200 ;
        RECT 367.600 306.800 368.400 307.700 ;
        RECT 364.400 301.600 365.200 306.200 ;
        RECT 367.600 301.600 368.400 306.200 ;
        RECT 369.200 301.600 370.000 307.700 ;
        RECT 375.600 301.600 376.400 306.200 ;
        RECT 381.600 301.600 382.400 306.200 ;
        RECT 383.600 301.600 384.400 306.200 ;
        RECT 388.800 301.600 389.600 306.200 ;
        RECT 394.800 301.600 395.600 306.200 ;
        RECT 398.000 301.600 398.800 305.400 ;
        RECT 404.400 301.600 405.200 305.400 ;
        RECT 410.800 301.600 411.600 304.200 ;
        RECT 415.600 301.600 416.400 305.400 ;
        RECT 420.400 301.600 421.200 305.400 ;
        RECT 428.400 301.600 429.200 306.200 ;
        RECT 438.000 301.600 438.800 304.200 ;
        RECT 441.200 301.600 442.000 304.200 ;
        RECT 452.400 301.600 453.200 306.200 ;
        RECT 458.800 301.600 459.600 304.200 ;
        RECT 466.800 301.600 467.600 305.400 ;
        RECT 471.600 301.600 472.400 304.200 ;
        RECT 476.400 301.600 477.200 305.400 ;
        RECT 484.400 301.600 485.200 305.400 ;
        RECT 490.800 301.600 491.600 305.400 ;
        RECT 494.000 301.600 494.800 304.200 ;
        RECT 498.200 301.600 499.000 306.200 ;
        RECT 502.000 301.600 502.800 305.400 ;
        RECT 508.400 301.600 509.200 305.400 ;
        RECT 516.400 301.600 517.200 306.200 ;
        RECT 521.200 301.600 522.000 306.200 ;
        RECT 526.000 301.600 526.800 305.400 ;
        RECT 530.800 301.600 531.600 306.200 ;
        RECT 534.000 301.600 534.800 306.200 ;
        RECT 540.400 301.600 541.200 306.200 ;
        RECT 543.600 301.600 544.400 306.200 ;
        RECT 545.200 301.600 546.000 306.200 ;
        RECT 548.400 301.600 549.200 306.200 ;
        RECT 553.200 301.600 554.000 306.200 ;
        RECT 562.800 301.600 563.600 304.200 ;
        RECT 566.000 301.600 566.800 304.200 ;
        RECT 577.200 301.600 578.000 306.200 ;
        RECT 583.600 301.600 584.400 304.200 ;
        RECT 588.400 301.600 589.200 305.400 ;
        RECT 593.200 301.600 594.000 304.200 ;
        RECT 598.000 301.600 598.800 305.400 ;
        RECT 602.800 301.600 603.600 304.200 ;
        RECT 606.000 301.600 606.800 306.200 ;
        RECT 0.400 300.400 614.000 301.600 ;
        RECT 1.200 295.800 2.000 300.400 ;
        RECT 4.400 295.800 5.200 300.400 ;
        RECT 7.600 295.800 8.400 300.400 ;
        RECT 10.800 295.800 11.600 300.400 ;
        RECT 14.000 295.800 14.800 300.400 ;
        RECT 18.800 295.800 19.600 300.400 ;
        RECT 28.400 297.800 29.200 300.400 ;
        RECT 31.600 297.800 32.400 300.400 ;
        RECT 42.800 295.800 43.600 300.400 ;
        RECT 49.200 297.800 50.000 300.400 ;
        RECT 50.800 297.800 51.600 300.400 ;
        RECT 54.000 297.800 54.800 300.400 ;
        RECT 55.600 297.800 56.400 300.400 ;
        RECT 59.800 295.800 60.600 300.400 ;
        RECT 65.200 295.800 66.000 300.400 ;
        RECT 74.800 297.800 75.600 300.400 ;
        RECT 78.000 297.800 78.800 300.400 ;
        RECT 89.200 295.800 90.000 300.400 ;
        RECT 95.600 297.800 96.400 300.400 ;
        RECT 97.200 297.800 98.000 300.400 ;
        RECT 100.400 297.800 101.200 300.400 ;
        RECT 102.000 297.800 102.800 300.400 ;
        RECT 106.200 295.800 107.000 300.400 ;
        RECT 108.400 297.800 109.200 300.400 ;
        RECT 113.200 295.400 114.000 300.400 ;
        RECT 118.400 295.000 119.200 300.400 ;
        RECT 121.200 297.800 122.000 300.400 ;
        RECT 127.600 295.800 128.400 300.400 ;
        RECT 138.800 297.800 139.600 300.400 ;
        RECT 142.000 297.800 142.800 300.400 ;
        RECT 151.600 295.800 152.400 300.400 ;
        RECT 161.200 297.800 162.000 300.400 ;
        RECT 166.000 296.600 166.800 300.400 ;
        RECT 174.000 295.800 174.800 300.400 ;
        RECT 183.600 297.800 184.400 300.400 ;
        RECT 186.800 297.800 187.600 300.400 ;
        RECT 198.000 295.800 198.800 300.400 ;
        RECT 204.400 297.800 205.200 300.400 ;
        RECT 206.000 295.800 206.800 300.400 ;
        RECT 209.200 295.800 210.000 300.400 ;
        RECT 214.000 295.800 214.800 300.400 ;
        RECT 222.000 295.800 222.800 300.400 ;
        RECT 231.600 297.800 232.400 300.400 ;
        RECT 234.800 297.800 235.600 300.400 ;
        RECT 246.000 295.800 246.800 300.400 ;
        RECT 252.400 297.800 253.200 300.400 ;
        RECT 254.000 297.800 254.800 300.400 ;
        RECT 258.400 295.000 259.200 300.400 ;
        RECT 263.600 295.400 264.400 300.400 ;
        RECT 270.000 295.800 270.800 300.400 ;
        RECT 279.600 297.800 280.400 300.400 ;
        RECT 282.800 297.800 283.600 300.400 ;
        RECT 294.000 295.800 294.800 300.400 ;
        RECT 300.400 297.800 301.200 300.400 ;
        RECT 302.000 295.800 302.800 300.400 ;
        RECT 311.600 295.800 312.400 300.400 ;
        RECT 316.400 295.800 317.200 300.400 ;
        RECT 322.800 296.600 323.600 300.400 ;
        RECT 329.200 296.600 330.000 300.400 ;
        RECT 334.000 295.800 334.800 300.400 ;
        RECT 338.800 297.800 339.600 300.400 ;
        RECT 342.000 297.800 342.800 300.400 ;
        RECT 345.200 297.800 346.000 300.400 ;
        RECT 345.200 296.300 346.000 297.200 ;
        RECT 346.800 296.300 347.600 300.400 ;
        RECT 345.200 295.700 347.600 296.300 ;
        RECT 345.200 295.600 346.000 295.700 ;
        RECT 346.800 293.800 347.600 295.700 ;
        RECT 353.200 293.800 354.000 300.400 ;
        RECT 361.200 295.400 362.000 300.400 ;
        RECT 366.400 295.000 367.200 300.400 ;
        RECT 372.400 295.800 373.200 300.400 ;
        RECT 374.000 294.300 374.800 300.400 ;
        RECT 380.400 295.800 381.200 300.400 ;
        RECT 383.600 295.800 384.400 300.400 ;
        RECT 385.200 295.800 386.000 300.400 ;
        RECT 391.200 295.800 392.000 300.400 ;
        RECT 393.200 295.800 394.000 300.400 ;
        RECT 398.000 297.800 398.800 300.400 ;
        RECT 404.400 295.800 405.200 300.400 ;
        RECT 415.600 297.800 416.400 300.400 ;
        RECT 418.800 297.800 419.600 300.400 ;
        RECT 428.400 295.800 429.200 300.400 ;
        RECT 433.200 295.800 434.000 300.400 ;
        RECT 439.200 295.800 440.000 300.400 ;
        RECT 441.200 295.800 442.000 300.400 ;
        RECT 447.200 295.800 448.000 300.400 ;
        RECT 450.800 297.800 451.600 300.400 ;
        RECT 454.000 297.800 454.800 300.400 ;
        RECT 374.000 293.800 376.300 294.300 ;
        RECT 460.400 293.800 461.200 300.400 ;
        RECT 466.800 293.800 467.600 300.400 ;
        RECT 473.800 295.800 474.600 300.400 ;
        RECT 478.000 297.800 478.800 300.400 ;
        RECT 482.800 295.800 483.600 300.400 ;
        RECT 485.000 295.800 485.800 300.400 ;
        RECT 489.200 297.800 490.000 300.400 ;
        RECT 490.800 297.800 491.600 300.400 ;
        RECT 494.000 297.800 494.800 300.400 ;
        RECT 495.600 295.800 496.400 300.400 ;
        RECT 503.600 296.600 504.400 300.400 ;
        RECT 508.400 296.600 509.200 300.400 ;
        RECT 513.200 295.800 514.000 300.400 ;
        RECT 518.000 297.800 518.800 300.400 ;
        RECT 521.200 297.800 522.000 300.400 ;
        RECT 522.800 297.800 523.600 300.400 ;
        RECT 526.000 297.800 526.800 300.400 ;
        RECT 527.600 295.800 528.400 300.400 ;
        RECT 534.000 296.600 534.800 300.400 ;
        RECT 537.200 297.800 538.000 300.400 ;
        RECT 543.600 295.800 544.400 300.400 ;
        RECT 554.800 297.800 555.600 300.400 ;
        RECT 558.000 297.800 558.800 300.400 ;
        RECT 567.600 295.800 568.400 300.400 ;
        RECT 572.400 295.800 573.200 300.400 ;
        RECT 580.400 295.800 581.200 300.400 ;
        RECT 590.000 297.800 590.800 300.400 ;
        RECT 593.200 297.800 594.000 300.400 ;
        RECT 604.400 295.800 605.200 300.400 ;
        RECT 610.800 297.800 611.600 300.400 ;
        RECT 353.300 291.200 353.900 293.800 ;
        RECT 374.100 293.700 376.300 293.800 ;
        RECT 375.700 292.400 376.300 293.700 ;
        RECT 375.600 291.600 377.200 292.400 ;
        RECT 353.200 289.600 354.000 291.200 ;
        RECT 388.400 270.800 389.200 272.400 ;
        RECT 370.800 269.600 372.400 270.400 ;
        RECT 172.000 268.400 172.800 269.200 ;
        RECT 172.200 267.600 173.200 268.400 ;
        RECT 370.900 268.300 371.500 269.600 ;
        RECT 369.300 268.200 371.500 268.300 ;
        RECT 388.500 268.200 389.100 270.800 ;
        RECT 369.200 267.700 371.500 268.200 ;
        RECT 4.400 261.600 5.200 266.200 ;
        RECT 14.000 261.600 14.800 264.200 ;
        RECT 17.200 261.600 18.000 264.200 ;
        RECT 28.400 261.600 29.200 266.200 ;
        RECT 34.800 261.600 35.600 264.200 ;
        RECT 36.400 261.600 37.200 264.200 ;
        RECT 42.800 261.600 43.600 266.200 ;
        RECT 54.000 261.600 54.800 264.200 ;
        RECT 57.200 261.600 58.000 264.200 ;
        RECT 66.800 261.600 67.600 266.200 ;
        RECT 71.600 261.600 72.400 264.200 ;
        RECT 74.800 261.600 75.600 264.200 ;
        RECT 76.400 261.600 77.200 264.200 ;
        RECT 80.600 261.600 81.400 266.200 ;
        RECT 82.800 261.600 83.600 264.200 ;
        RECT 89.200 261.600 90.000 266.200 ;
        RECT 100.400 261.600 101.200 264.200 ;
        RECT 103.600 261.600 104.400 264.200 ;
        RECT 113.200 261.600 114.000 266.200 ;
        RECT 118.000 261.600 118.800 264.200 ;
        RECT 122.200 261.600 123.000 266.200 ;
        RECT 124.400 261.600 125.200 266.200 ;
        RECT 127.600 261.600 128.400 266.200 ;
        RECT 130.800 261.600 131.600 266.200 ;
        RECT 134.000 261.600 134.800 266.200 ;
        RECT 137.200 261.600 138.000 266.200 ;
        RECT 138.800 261.600 139.600 266.200 ;
        RECT 142.000 261.600 142.800 266.200 ;
        RECT 145.200 261.600 146.000 266.200 ;
        RECT 148.400 261.600 149.200 266.200 ;
        RECT 151.600 261.600 152.400 266.200 ;
        RECT 159.600 261.600 160.400 266.200 ;
        RECT 162.800 261.600 163.600 266.200 ;
        RECT 164.400 261.600 165.200 264.200 ;
        RECT 167.600 261.600 168.400 264.200 ;
        RECT 170.800 261.600 171.600 265.800 ;
        RECT 174.000 261.600 174.800 264.200 ;
        RECT 178.800 261.600 179.600 266.200 ;
        RECT 188.400 261.600 189.200 264.200 ;
        RECT 191.600 261.600 192.400 264.200 ;
        RECT 202.800 261.600 203.600 266.200 ;
        RECT 209.200 261.600 210.000 264.200 ;
        RECT 212.400 261.600 213.200 266.200 ;
        RECT 214.000 261.600 214.800 266.200 ;
        RECT 218.800 261.600 219.600 266.200 ;
        RECT 223.600 261.600 224.400 266.200 ;
        RECT 226.800 261.600 227.600 266.200 ;
        RECT 230.000 261.600 230.800 266.200 ;
        RECT 234.800 261.600 235.600 266.200 ;
        RECT 244.400 261.600 245.200 264.200 ;
        RECT 247.600 261.600 248.400 264.200 ;
        RECT 258.800 261.600 259.600 266.200 ;
        RECT 265.200 261.600 266.000 264.200 ;
        RECT 268.400 261.600 269.200 266.600 ;
        RECT 273.600 261.600 274.400 267.000 ;
        RECT 278.000 261.600 278.800 264.200 ;
        RECT 282.800 261.600 283.600 265.400 ;
        RECT 287.600 261.600 288.400 265.400 ;
        RECT 292.400 261.600 293.200 264.200 ;
        RECT 297.200 261.600 298.000 266.600 ;
        RECT 302.400 261.600 303.200 267.000 ;
        RECT 313.200 261.600 314.000 266.200 ;
        RECT 322.800 261.600 323.600 264.200 ;
        RECT 326.000 261.600 326.800 264.200 ;
        RECT 337.200 261.600 338.000 266.200 ;
        RECT 343.600 261.600 344.400 264.200 ;
        RECT 346.800 261.600 347.600 264.200 ;
        RECT 351.600 261.600 352.400 265.400 ;
        RECT 356.400 261.600 357.200 265.400 ;
        RECT 362.800 261.600 363.600 264.200 ;
        RECT 367.600 261.600 368.400 266.200 ;
        RECT 369.200 261.600 370.000 267.700 ;
        RECT 375.600 261.600 376.400 268.200 ;
        RECT 382.000 261.600 382.800 268.200 ;
        RECT 388.400 261.600 389.200 268.200 ;
        RECT 395.200 261.600 396.000 266.200 ;
        RECT 401.200 261.600 402.000 266.200 ;
        RECT 403.200 261.600 404.000 266.200 ;
        RECT 409.200 261.600 410.000 266.200 ;
        RECT 410.800 261.600 411.600 266.200 ;
        RECT 415.600 261.600 416.400 266.200 ;
        RECT 421.600 261.600 422.400 266.200 ;
        RECT 423.600 261.600 424.400 266.200 ;
        RECT 429.600 261.600 430.400 266.200 ;
        RECT 431.600 261.600 432.400 268.200 ;
        RECT 442.800 261.600 443.600 268.200 ;
        RECT 444.400 261.600 445.200 266.200 ;
        RECT 450.400 261.600 451.200 266.200 ;
        RECT 457.200 261.600 458.000 268.200 ;
        RECT 463.600 261.600 464.400 268.200 ;
        RECT 470.000 261.600 470.800 268.200 ;
        RECT 476.400 261.600 477.200 268.200 ;
        RECT 482.800 261.600 483.600 264.200 ;
        RECT 486.000 261.600 486.800 264.200 ;
        RECT 492.400 261.600 493.200 265.400 ;
        RECT 496.200 261.600 497.000 266.200 ;
        RECT 500.400 261.600 501.200 264.200 ;
        RECT 502.000 261.600 502.800 264.200 ;
        RECT 505.200 261.600 506.000 264.200 ;
        RECT 510.000 261.600 510.800 265.400 ;
        RECT 513.200 261.600 514.000 264.200 ;
        RECT 516.400 261.600 517.200 264.200 ;
        RECT 518.000 261.600 518.800 264.200 ;
        RECT 521.200 261.600 522.000 264.200 ;
        RECT 524.400 261.600 525.200 265.400 ;
        RECT 530.800 261.600 531.600 265.400 ;
        RECT 540.400 261.600 541.200 266.200 ;
        RECT 543.600 261.600 544.400 264.200 ;
        RECT 548.400 261.600 549.200 266.200 ;
        RECT 553.200 261.600 554.000 266.200 ;
        RECT 556.400 261.600 557.200 265.400 ;
        RECT 561.200 261.600 562.000 266.200 ;
        RECT 567.600 261.600 568.400 265.400 ;
        RECT 572.400 261.600 573.200 266.200 ;
        RECT 577.200 261.600 578.000 264.200 ;
        RECT 583.600 261.600 584.400 266.200 ;
        RECT 594.800 261.600 595.600 264.200 ;
        RECT 598.000 261.600 598.800 264.200 ;
        RECT 607.600 261.600 608.400 266.200 ;
        RECT 0.400 260.400 614.000 261.600 ;
        RECT 4.400 255.800 5.200 260.400 ;
        RECT 14.000 257.800 14.800 260.400 ;
        RECT 17.200 257.800 18.000 260.400 ;
        RECT 28.400 255.800 29.200 260.400 ;
        RECT 34.800 257.800 35.600 260.400 ;
        RECT 38.000 257.800 38.800 260.400 ;
        RECT 42.800 255.800 43.600 260.400 ;
        RECT 52.400 257.800 53.200 260.400 ;
        RECT 55.600 257.800 56.400 260.400 ;
        RECT 66.800 255.800 67.600 260.400 ;
        RECT 73.200 257.800 74.000 260.400 ;
        RECT 74.800 257.800 75.600 260.400 ;
        RECT 78.000 257.800 78.800 260.400 ;
        RECT 79.600 257.800 80.400 260.400 ;
        RECT 83.800 255.800 84.600 260.400 ;
        RECT 87.600 257.800 88.400 260.400 ;
        RECT 89.200 257.800 90.000 260.400 ;
        RECT 92.400 257.800 93.200 260.400 ;
        RECT 94.000 257.800 94.800 260.400 ;
        RECT 100.400 255.800 101.200 260.400 ;
        RECT 111.600 257.800 112.400 260.400 ;
        RECT 114.800 257.800 115.600 260.400 ;
        RECT 124.400 255.800 125.200 260.400 ;
        RECT 130.800 257.800 131.600 260.400 ;
        RECT 132.400 255.800 133.200 260.400 ;
        RECT 135.600 255.800 136.400 260.400 ;
        RECT 143.600 257.800 144.400 260.400 ;
        RECT 150.000 255.800 150.800 260.400 ;
        RECT 161.200 257.800 162.000 260.400 ;
        RECT 164.400 257.800 165.200 260.400 ;
        RECT 172.400 258.300 173.200 258.400 ;
        RECT 174.000 258.300 174.800 260.400 ;
        RECT 172.400 257.700 174.800 258.300 ;
        RECT 172.400 257.600 173.200 257.700 ;
        RECT 174.000 255.800 174.800 257.700 ;
        RECT 178.800 255.800 179.600 260.400 ;
        RECT 186.800 256.600 187.600 260.400 ;
        RECT 190.000 255.800 190.800 260.400 ;
        RECT 193.200 255.800 194.000 260.400 ;
        RECT 198.000 255.800 198.800 260.400 ;
        RECT 207.600 257.800 208.400 260.400 ;
        RECT 210.800 257.800 211.600 260.400 ;
        RECT 222.000 255.800 222.800 260.400 ;
        RECT 228.400 257.800 229.200 260.400 ;
        RECT 230.000 257.800 230.800 260.400 ;
        RECT 234.400 255.000 235.200 260.400 ;
        RECT 239.600 255.400 240.400 260.400 ;
        RECT 242.800 255.800 243.600 260.400 ;
        RECT 246.000 255.800 246.800 260.400 ;
        RECT 249.200 257.800 250.000 260.400 ;
        RECT 255.600 255.800 256.400 260.400 ;
        RECT 266.800 257.800 267.600 260.400 ;
        RECT 270.000 257.800 270.800 260.400 ;
        RECT 279.600 255.800 280.400 260.400 ;
        RECT 289.200 256.600 290.000 260.400 ;
        RECT 295.600 256.600 296.400 260.400 ;
        RECT 298.800 255.800 299.600 260.400 ;
        RECT 308.400 257.800 309.200 260.400 ;
        RECT 311.600 256.200 312.400 260.400 ;
        RECT 314.800 255.800 315.600 260.400 ;
        RECT 318.000 255.800 318.800 260.400 ;
        RECT 324.400 256.600 325.200 260.400 ;
        RECT 332.400 256.600 333.200 260.400 ;
        RECT 338.800 255.800 339.600 260.400 ;
        RECT 325.200 254.400 326.000 254.800 ;
        RECT 310.000 253.600 311.000 254.400 ;
        RECT 325.200 253.800 326.800 254.400 ;
        RECT 340.400 253.800 341.200 260.400 ;
        RECT 348.400 255.800 349.200 260.400 ;
        RECT 354.800 255.800 355.600 260.400 ;
        RECT 364.400 257.800 365.200 260.400 ;
        RECT 367.600 257.800 368.400 260.400 ;
        RECT 378.800 255.800 379.600 260.400 ;
        RECT 385.200 257.800 386.000 260.400 ;
        RECT 388.400 257.800 389.200 260.400 ;
        RECT 390.000 253.800 390.800 260.400 ;
        RECT 396.400 255.800 397.200 260.400 ;
        RECT 402.400 255.800 403.200 260.400 ;
        RECT 404.400 255.800 405.200 260.400 ;
        RECT 410.400 255.800 411.200 260.400 ;
        RECT 412.400 255.800 413.200 260.400 ;
        RECT 417.200 253.800 418.000 260.400 ;
        RECT 426.800 255.800 427.600 260.400 ;
        RECT 428.800 255.800 429.600 260.400 ;
        RECT 434.800 255.800 435.600 260.400 ;
        RECT 436.400 255.800 437.200 260.400 ;
        RECT 444.400 255.800 445.200 260.400 ;
        RECT 446.000 253.800 446.800 260.400 ;
        RECT 452.400 255.800 453.200 260.400 ;
        RECT 458.400 255.800 459.200 260.400 ;
        RECT 465.200 255.800 466.000 260.400 ;
        RECT 471.200 255.800 472.000 260.400 ;
        RECT 473.200 253.800 474.000 260.400 ;
        RECT 479.600 257.800 480.400 260.400 ;
        RECT 482.800 257.800 483.600 260.400 ;
        RECT 484.400 257.800 485.200 260.400 ;
        RECT 487.600 257.800 488.400 260.400 ;
        RECT 490.800 257.800 491.600 260.400 ;
        RECT 494.000 257.800 494.800 260.400 ;
        RECT 496.200 255.800 497.000 260.400 ;
        RECT 500.400 257.800 501.200 260.400 ;
        RECT 505.200 255.800 506.000 260.400 ;
        RECT 511.600 253.800 512.400 260.400 ;
        RECT 513.200 257.800 514.000 260.400 ;
        RECT 516.400 257.800 517.200 260.400 ;
        RECT 522.800 256.600 523.600 260.400 ;
        RECT 530.800 256.600 531.600 260.400 ;
        RECT 534.000 257.800 534.800 260.400 ;
        RECT 542.000 256.600 542.800 260.400 ;
        RECT 545.200 255.800 546.000 260.400 ;
        RECT 550.000 256.600 550.800 260.400 ;
        RECT 554.800 255.800 555.600 260.400 ;
        RECT 558.000 255.800 558.800 260.400 ;
        RECT 561.200 255.800 562.000 260.400 ;
        RECT 564.400 255.800 565.200 260.400 ;
        RECT 567.600 255.800 568.400 260.400 ;
        RECT 569.200 257.800 570.000 260.400 ;
        RECT 575.600 255.800 576.400 260.400 ;
        RECT 586.800 257.800 587.600 260.400 ;
        RECT 590.000 257.800 590.800 260.400 ;
        RECT 599.600 255.800 600.400 260.400 ;
        RECT 606.000 255.800 606.800 260.400 ;
        RECT 326.000 253.600 326.800 253.800 ;
        RECT 295.600 251.600 296.400 253.200 ;
        RECT 310.400 252.800 311.200 253.600 ;
        RECT 340.500 251.200 341.100 253.800 ;
        RECT 390.100 251.200 390.700 253.800 ;
        RECT 340.400 249.600 341.200 251.200 ;
        RECT 390.000 249.600 390.800 251.200 ;
        RECT 1.200 221.600 2.000 224.200 ;
        RECT 4.400 221.600 5.200 224.200 ;
        RECT 9.200 221.600 10.000 225.400 ;
        RECT 15.600 221.600 16.400 225.400 ;
        RECT 22.000 221.600 22.800 225.400 ;
        RECT 26.800 221.600 27.600 226.200 ;
        RECT 33.200 221.600 34.000 225.400 ;
        RECT 39.600 221.600 40.400 224.200 ;
        RECT 41.200 221.600 42.000 224.200 ;
        RECT 47.600 221.600 48.400 226.200 ;
        RECT 57.200 221.600 58.000 224.200 ;
        RECT 60.400 221.600 61.200 224.200 ;
        RECT 71.600 221.600 72.400 226.200 ;
        RECT 78.000 221.600 78.800 224.200 ;
        RECT 82.800 221.600 83.600 226.200 ;
        RECT 84.400 221.600 85.200 226.200 ;
        RECT 87.600 221.600 88.400 226.200 ;
        RECT 90.800 221.600 91.600 226.200 ;
        RECT 94.000 221.600 94.800 226.200 ;
        RECT 97.200 221.600 98.000 226.200 ;
        RECT 100.400 221.600 101.200 226.200 ;
        RECT 103.600 221.600 104.400 226.200 ;
        RECT 106.800 221.600 107.600 226.200 ;
        RECT 112.200 221.600 113.200 224.200 ;
        RECT 115.600 221.600 116.400 224.200 ;
        RECT 121.200 221.600 122.000 226.000 ;
        RECT 127.600 221.600 128.400 225.400 ;
        RECT 130.800 221.600 131.600 224.200 ;
        RECT 134.000 221.600 134.800 224.200 ;
        RECT 137.200 221.600 138.000 225.400 ;
        RECT 143.600 221.600 144.400 224.200 ;
        RECT 153.200 221.600 154.000 226.200 ;
        RECT 162.800 221.600 163.600 224.200 ;
        RECT 166.000 221.600 166.800 224.200 ;
        RECT 177.200 221.600 178.000 226.200 ;
        RECT 183.600 221.600 184.400 224.200 ;
        RECT 185.200 221.600 186.000 224.200 ;
        RECT 191.600 221.600 192.400 226.200 ;
        RECT 201.200 221.600 202.000 224.200 ;
        RECT 204.400 221.600 205.200 224.200 ;
        RECT 215.600 221.600 216.400 226.200 ;
        RECT 222.000 221.600 222.800 224.200 ;
        RECT 223.600 221.600 224.400 226.200 ;
        RECT 226.800 221.600 227.600 226.200 ;
        RECT 230.000 221.600 230.800 226.200 ;
        RECT 234.800 221.600 235.600 226.200 ;
        RECT 244.400 221.600 245.200 224.200 ;
        RECT 247.600 221.600 248.400 224.200 ;
        RECT 258.800 221.600 259.600 226.200 ;
        RECT 265.200 221.600 266.000 224.200 ;
        RECT 270.000 221.600 270.800 226.200 ;
        RECT 274.800 221.600 275.600 226.200 ;
        RECT 276.400 221.600 277.200 226.200 ;
        RECT 282.800 221.600 283.600 225.400 ;
        RECT 287.600 221.600 288.400 224.200 ;
        RECT 292.400 221.600 293.200 225.400 ;
        RECT 297.200 221.600 298.000 225.400 ;
        RECT 302.000 221.600 302.800 226.200 ;
        RECT 313.200 221.600 314.000 225.400 ;
        RECT 318.000 221.600 318.800 228.200 ;
        RECT 324.400 221.600 325.200 226.200 ;
        RECT 327.600 221.600 328.400 226.200 ;
        RECT 330.800 221.600 331.600 226.200 ;
        RECT 334.000 221.600 334.800 226.200 ;
        RECT 337.200 221.600 338.000 226.200 ;
        RECT 338.800 221.600 339.600 228.200 ;
        RECT 345.200 221.600 346.000 228.200 ;
        RECT 351.600 221.600 352.400 228.200 ;
        RECT 359.600 221.600 360.400 226.600 ;
        RECT 364.800 221.600 365.600 227.000 ;
        RECT 370.800 221.600 371.600 226.200 ;
        RECT 380.400 221.600 381.200 224.200 ;
        RECT 383.600 221.600 384.400 224.200 ;
        RECT 394.800 221.600 395.600 226.200 ;
        RECT 401.200 221.600 402.000 224.200 ;
        RECT 404.400 221.600 405.200 224.200 ;
        RECT 409.200 221.600 410.000 226.200 ;
        RECT 412.400 221.600 413.200 226.200 ;
        RECT 415.600 221.600 416.400 226.200 ;
        RECT 417.200 221.600 418.000 226.200 ;
        RECT 420.400 221.600 421.200 226.200 ;
        RECT 423.600 221.600 424.400 226.200 ;
        RECT 426.800 221.600 427.600 226.200 ;
        RECT 430.000 221.600 430.800 226.200 ;
        RECT 431.600 221.600 432.400 226.200 ;
        RECT 434.800 221.600 435.600 226.200 ;
        RECT 438.000 221.600 438.800 226.200 ;
        RECT 441.200 221.600 442.000 226.200 ;
        RECT 444.400 221.600 445.200 226.200 ;
        RECT 446.400 221.600 447.200 226.200 ;
        RECT 452.400 221.600 453.200 226.200 ;
        RECT 454.000 221.600 454.800 226.200 ;
        RECT 460.000 221.600 460.800 226.200 ;
        RECT 466.800 221.600 467.600 226.200 ;
        RECT 471.600 221.600 472.400 228.200 ;
        RECT 478.000 221.600 478.800 226.200 ;
        RECT 483.200 221.600 484.000 226.200 ;
        RECT 489.200 221.600 490.000 226.200 ;
        RECT 495.600 221.600 496.400 228.200 ;
        RECT 497.200 221.600 498.000 224.200 ;
        RECT 501.400 221.600 502.200 226.200 ;
        RECT 508.400 221.600 509.200 228.200 ;
        RECT 514.800 221.600 515.600 228.200 ;
        RECT 516.400 221.600 517.200 228.200 ;
        RECT 522.800 221.600 523.600 228.200 ;
        RECT 529.200 221.600 530.000 228.200 ;
        RECT 540.400 221.600 541.200 228.200 ;
        RECT 546.800 221.600 547.600 228.200 ;
        RECT 551.600 221.600 552.400 226.200 ;
        RECT 553.200 221.600 554.000 226.200 ;
        RECT 556.400 221.600 557.200 228.200 ;
        RECT 566.000 221.600 566.800 226.200 ;
        RECT 567.600 221.600 568.400 224.200 ;
        RECT 574.000 221.600 574.800 226.200 ;
        RECT 585.200 221.600 586.000 224.200 ;
        RECT 588.400 221.600 589.200 224.200 ;
        RECT 598.000 221.600 598.800 226.200 ;
        RECT 604.400 221.600 605.200 225.400 ;
        RECT 0.400 220.400 614.000 221.600 ;
        RECT 1.200 217.800 2.000 220.400 ;
        RECT 6.000 216.600 6.800 220.400 ;
        RECT 12.400 216.200 13.200 220.400 ;
        RECT 15.600 217.800 16.400 220.400 ;
        RECT 18.800 216.600 19.600 220.400 ;
        RECT 23.600 215.800 24.400 220.400 ;
        RECT 31.600 216.600 32.400 220.400 ;
        RECT 38.000 216.600 38.800 220.400 ;
        RECT 41.200 215.800 42.000 220.400 ;
        RECT 44.400 215.800 45.200 220.400 ;
        RECT 47.600 215.800 48.400 220.400 ;
        RECT 50.800 215.800 51.600 220.400 ;
        RECT 54.000 215.800 54.800 220.400 ;
        RECT 55.600 215.800 56.400 220.400 ;
        RECT 58.800 215.800 59.600 220.400 ;
        RECT 62.000 215.800 62.800 220.400 ;
        RECT 65.200 215.800 66.000 220.400 ;
        RECT 68.400 215.800 69.200 220.400 ;
        RECT 71.200 215.000 72.000 220.400 ;
        RECT 76.400 215.400 77.200 220.400 ;
        RECT 81.200 216.000 82.000 220.400 ;
        RECT 86.800 217.800 87.600 220.400 ;
        RECT 90.000 217.800 91.000 220.400 ;
        RECT 95.600 215.800 96.400 220.400 ;
        RECT 100.400 216.600 101.200 220.400 ;
        RECT 108.400 216.600 109.200 220.400 ;
        RECT 113.200 216.600 114.000 220.400 ;
        RECT 121.200 216.600 122.000 220.400 ;
        RECT 126.000 216.600 126.800 220.400 ;
        RECT 134.000 216.600 134.800 220.400 ;
        RECT 138.800 216.000 139.600 220.400 ;
        RECT 144.400 217.800 145.200 220.400 ;
        RECT 147.600 217.800 148.600 220.400 ;
        RECT 153.200 215.800 154.000 220.400 ;
        RECT 161.200 217.800 162.000 220.400 ;
        RECT 164.400 217.800 165.200 220.400 ;
        RECT 167.600 216.400 168.600 220.400 ;
        RECT 173.800 219.800 174.600 220.400 ;
        RECT 173.800 216.400 174.800 219.800 ;
        RECT 177.200 217.800 178.000 220.400 ;
        RECT 183.600 215.800 184.400 220.400 ;
        RECT 194.800 217.800 195.600 220.400 ;
        RECT 198.000 217.800 198.800 220.400 ;
        RECT 207.600 215.800 208.400 220.400 ;
        RECT 215.600 215.800 216.400 220.400 ;
        RECT 225.200 217.800 226.000 220.400 ;
        RECT 228.400 217.800 229.200 220.400 ;
        RECT 239.600 215.800 240.400 220.400 ;
        RECT 246.000 217.800 246.800 220.400 ;
        RECT 247.600 217.800 248.400 220.400 ;
        RECT 254.000 215.800 254.800 220.400 ;
        RECT 263.600 217.800 264.400 220.400 ;
        RECT 266.800 217.800 267.600 220.400 ;
        RECT 278.000 215.800 278.800 220.400 ;
        RECT 284.400 217.800 285.200 220.400 ;
        RECT 287.600 217.800 288.400 220.400 ;
        RECT 289.200 215.800 290.000 220.400 ;
        RECT 292.400 215.800 293.200 220.400 ;
        RECT 295.600 215.800 296.400 220.400 ;
        RECT 298.800 215.800 299.600 220.400 ;
        RECT 302.000 215.800 302.800 220.400 ;
        RECT 308.400 217.800 309.200 220.400 ;
        RECT 314.800 215.800 315.600 220.400 ;
        RECT 326.000 217.800 326.800 220.400 ;
        RECT 329.200 217.800 330.000 220.400 ;
        RECT 338.800 215.800 339.600 220.400 ;
        RECT 345.200 216.600 346.000 220.400 ;
        RECT 350.000 217.800 350.800 220.400 ;
        RECT 356.400 215.800 357.200 220.400 ;
        RECT 367.600 217.800 368.400 220.400 ;
        RECT 370.800 217.800 371.600 220.400 ;
        RECT 380.400 215.800 381.200 220.400 ;
        RECT 385.200 215.800 386.000 220.400 ;
        RECT 390.000 215.800 390.800 220.400 ;
        RECT 393.200 215.800 394.000 220.400 ;
        RECT 396.400 215.800 397.200 220.400 ;
        RECT 399.600 215.800 400.400 220.400 ;
        RECT 402.800 215.800 403.600 220.400 ;
        RECT 406.000 216.600 406.800 220.400 ;
        RECT 410.800 217.800 411.600 220.400 ;
        RECT 415.600 215.800 416.400 220.400 ;
        RECT 418.800 215.800 419.600 220.400 ;
        RECT 420.400 215.800 421.200 220.400 ;
        RECT 425.200 217.800 426.000 220.400 ;
        RECT 431.600 215.800 432.400 220.400 ;
        RECT 442.800 217.800 443.600 220.400 ;
        RECT 446.000 217.800 446.800 220.400 ;
        RECT 455.600 215.800 456.400 220.400 ;
        RECT 465.200 217.800 466.000 220.400 ;
        RECT 468.400 217.800 469.200 220.400 ;
        RECT 471.600 217.800 472.400 220.400 ;
        RECT 474.800 217.800 475.600 220.400 ;
        RECT 478.000 217.800 478.800 220.400 ;
        RECT 483.400 216.000 484.200 220.400 ;
        RECT 490.800 215.800 491.600 220.400 ;
        RECT 500.400 217.800 501.200 220.400 ;
        RECT 503.600 217.800 504.400 220.400 ;
        RECT 514.800 215.800 515.600 220.400 ;
        RECT 521.200 217.800 522.000 220.400 ;
        RECT 522.800 217.800 523.600 220.400 ;
        RECT 527.600 216.600 528.400 220.400 ;
        RECT 535.600 215.800 536.400 220.400 ;
        RECT 537.200 217.800 538.000 220.400 ;
        RECT 543.600 215.800 544.400 220.400 ;
        RECT 554.800 217.800 555.600 220.400 ;
        RECT 558.000 217.800 558.800 220.400 ;
        RECT 567.600 215.800 568.400 220.400 ;
        RECT 574.000 216.600 574.800 220.400 ;
        RECT 578.800 215.800 579.600 220.400 ;
        RECT 582.000 215.800 582.800 220.400 ;
        RECT 585.200 215.800 586.000 220.400 ;
        RECT 588.400 215.800 589.200 220.400 ;
        RECT 591.600 215.800 592.400 220.400 ;
        RECT 593.200 215.800 594.000 220.400 ;
        RECT 596.400 215.800 597.200 220.400 ;
        RECT 599.600 215.800 600.400 220.400 ;
        RECT 602.800 215.800 603.600 220.400 ;
        RECT 606.000 215.800 606.800 220.400 ;
        RECT 4.400 181.600 5.200 186.200 ;
        RECT 14.000 181.600 14.800 184.200 ;
        RECT 17.200 181.600 18.000 184.200 ;
        RECT 28.400 181.600 29.200 186.200 ;
        RECT 34.800 181.600 35.600 184.200 ;
        RECT 38.000 181.600 38.800 184.200 ;
        RECT 41.200 181.600 42.000 186.200 ;
        RECT 46.600 181.600 47.600 184.200 ;
        RECT 50.000 181.600 50.800 184.200 ;
        RECT 55.600 181.600 56.400 186.000 ;
        RECT 62.000 181.600 62.800 185.400 ;
        RECT 66.800 181.600 67.600 185.400 ;
        RECT 72.800 181.600 73.600 187.000 ;
        RECT 78.000 181.600 78.800 186.600 ;
        RECT 81.200 181.600 82.000 186.200 ;
        RECT 84.400 181.600 85.200 186.200 ;
        RECT 89.200 181.600 90.000 186.200 ;
        RECT 94.600 181.600 95.600 184.200 ;
        RECT 98.000 181.600 98.800 184.200 ;
        RECT 103.600 181.600 104.400 186.000 ;
        RECT 108.400 181.600 109.200 185.400 ;
        RECT 114.800 181.600 115.600 186.600 ;
        RECT 120.000 181.600 120.800 187.000 ;
        RECT 126.000 181.600 126.800 185.400 ;
        RECT 130.800 181.600 131.600 186.600 ;
        RECT 136.000 181.600 136.800 187.000 ;
        RECT 140.400 181.600 141.200 186.200 ;
        RECT 143.600 181.600 144.400 186.200 ;
        RECT 146.800 181.600 147.600 184.200 ;
        RECT 148.400 181.600 149.200 184.200 ;
        RECT 151.600 181.600 152.400 184.200 ;
        RECT 159.600 181.600 160.400 184.200 ;
        RECT 162.800 182.200 163.800 185.600 ;
        RECT 163.000 181.600 163.800 182.200 ;
        RECT 169.000 181.600 170.000 185.600 ;
        RECT 172.400 181.600 173.200 184.200 ;
        RECT 178.800 181.600 179.600 186.200 ;
        RECT 190.000 181.600 190.800 184.200 ;
        RECT 193.200 181.600 194.000 184.200 ;
        RECT 202.800 181.600 203.600 186.200 ;
        RECT 210.800 181.600 211.600 186.200 ;
        RECT 214.000 181.600 214.800 185.400 ;
        RECT 220.400 181.600 221.200 186.200 ;
        RECT 223.600 181.600 224.400 186.200 ;
        RECT 226.800 181.600 227.600 186.200 ;
        RECT 230.000 181.600 230.800 186.200 ;
        RECT 233.200 181.600 234.000 185.400 ;
        RECT 239.600 181.600 240.400 185.400 ;
        RECT 244.400 181.600 245.200 186.200 ;
        RECT 249.200 181.600 250.000 186.200 ;
        RECT 252.400 181.600 253.200 186.200 ;
        RECT 258.800 181.600 259.600 186.200 ;
        RECT 268.400 181.600 269.200 184.200 ;
        RECT 271.600 181.600 272.400 184.200 ;
        RECT 282.800 181.600 283.600 186.200 ;
        RECT 289.200 181.600 290.000 184.200 ;
        RECT 294.000 181.600 294.800 185.400 ;
        RECT 298.800 181.600 299.600 186.200 ;
        RECT 302.000 181.600 302.800 186.200 ;
        RECT 308.400 181.600 309.200 184.200 ;
        RECT 311.600 181.600 312.400 184.200 ;
        RECT 314.800 181.600 315.600 184.200 ;
        RECT 318.000 181.600 318.800 185.400 ;
        RECT 322.800 181.600 323.600 184.200 ;
        RECT 329.200 181.600 330.000 186.200 ;
        RECT 340.400 181.600 341.200 184.200 ;
        RECT 343.600 181.600 344.400 184.200 ;
        RECT 353.200 181.600 354.000 186.200 ;
        RECT 361.200 181.600 362.000 185.400 ;
        RECT 364.400 181.600 365.200 184.200 ;
        RECT 370.800 181.600 371.600 186.200 ;
        RECT 382.000 181.600 382.800 184.200 ;
        RECT 385.200 181.600 386.000 184.200 ;
        RECT 394.800 181.600 395.600 186.200 ;
        RECT 402.800 181.600 403.600 186.200 ;
        RECT 412.400 181.600 413.200 184.200 ;
        RECT 415.600 181.600 416.400 184.200 ;
        RECT 426.800 181.600 427.600 186.200 ;
        RECT 433.200 181.600 434.000 184.200 ;
        RECT 438.000 181.600 438.800 186.200 ;
        RECT 447.600 181.600 448.400 184.200 ;
        RECT 450.800 181.600 451.600 184.200 ;
        RECT 462.000 181.600 462.800 186.200 ;
        RECT 468.400 181.600 469.200 184.200 ;
        RECT 476.400 181.600 477.200 186.200 ;
        RECT 481.800 181.600 482.800 184.200 ;
        RECT 485.200 181.600 486.000 184.200 ;
        RECT 490.800 181.600 491.600 186.000 ;
        RECT 495.600 181.600 496.400 185.400 ;
        RECT 503.600 181.600 504.400 186.200 ;
        RECT 505.200 181.600 506.000 186.200 ;
        RECT 508.400 181.600 509.200 186.200 ;
        RECT 511.600 181.600 512.400 186.200 ;
        RECT 513.200 181.600 514.000 184.200 ;
        RECT 516.400 181.600 517.200 184.200 ;
        RECT 521.200 181.600 522.000 185.400 ;
        RECT 526.000 181.600 526.800 184.200 ;
        RECT 527.600 181.600 528.400 184.200 ;
        RECT 534.000 181.600 534.800 186.200 ;
        RECT 545.200 181.600 546.000 184.200 ;
        RECT 548.400 181.600 549.200 184.200 ;
        RECT 558.000 181.600 558.800 186.200 ;
        RECT 566.000 181.600 566.800 186.200 ;
        RECT 575.600 181.600 576.400 184.200 ;
        RECT 578.800 181.600 579.600 184.200 ;
        RECT 590.000 181.600 590.800 186.200 ;
        RECT 596.400 181.600 597.200 184.200 ;
        RECT 601.200 181.600 602.000 185.400 ;
        RECT 606.000 181.600 606.800 186.200 ;
        RECT 0.400 180.400 614.000 181.600 ;
        RECT 2.800 175.800 3.600 180.400 ;
        RECT 8.200 177.800 9.200 180.400 ;
        RECT 11.600 177.800 12.400 180.400 ;
        RECT 17.200 176.000 18.000 180.400 ;
        RECT 23.600 176.600 24.400 180.400 ;
        RECT 28.400 175.400 29.200 180.400 ;
        RECT 33.600 175.000 34.400 180.400 ;
        RECT 36.400 175.800 37.200 180.400 ;
        RECT 39.600 175.800 40.400 180.400 ;
        RECT 46.000 176.600 46.800 180.400 ;
        RECT 50.800 177.800 51.600 180.400 ;
        RECT 54.000 176.000 54.800 180.400 ;
        RECT 59.600 177.800 60.400 180.400 ;
        RECT 62.800 177.800 63.800 180.400 ;
        RECT 68.400 175.800 69.200 180.400 ;
        RECT 72.800 175.000 73.600 180.400 ;
        RECT 78.000 175.400 78.800 180.400 ;
        RECT 82.800 176.600 83.600 180.400 ;
        RECT 90.800 176.600 91.600 180.400 ;
        RECT 94.000 177.800 94.800 180.400 ;
        RECT 98.400 175.000 99.200 180.400 ;
        RECT 103.600 175.400 104.400 180.400 ;
        RECT 106.800 177.800 107.600 180.400 ;
        RECT 110.000 175.800 110.800 180.400 ;
        RECT 114.800 177.800 115.600 180.400 ;
        RECT 118.000 177.800 118.800 180.400 ;
        RECT 124.400 175.800 125.200 180.400 ;
        RECT 126.000 177.800 126.800 180.400 ;
        RECT 129.200 177.800 130.000 180.400 ;
        RECT 130.800 175.800 131.600 180.400 ;
        RECT 134.000 175.800 134.800 180.400 ;
        RECT 137.200 177.800 138.000 180.400 ;
        RECT 140.400 177.800 141.200 180.400 ;
        RECT 143.600 177.800 144.400 180.400 ;
        RECT 150.000 177.800 150.800 180.400 ;
        RECT 156.400 175.800 157.200 180.400 ;
        RECT 167.600 177.800 168.400 180.400 ;
        RECT 170.800 177.800 171.600 180.400 ;
        RECT 180.400 175.800 181.200 180.400 ;
        RECT 185.200 175.800 186.000 180.400 ;
        RECT 188.400 175.800 189.200 180.400 ;
        RECT 194.800 175.800 195.600 180.400 ;
        RECT 199.600 175.800 200.400 180.400 ;
        RECT 204.400 176.600 205.200 180.400 ;
        RECT 207.600 177.800 208.400 180.400 ;
        RECT 214.000 175.800 214.800 180.400 ;
        RECT 225.200 177.800 226.000 180.400 ;
        RECT 228.400 177.800 229.200 180.400 ;
        RECT 238.000 175.800 238.800 180.400 ;
        RECT 246.000 175.800 246.800 180.400 ;
        RECT 255.600 177.800 256.400 180.400 ;
        RECT 258.800 177.800 259.600 180.400 ;
        RECT 270.000 175.800 270.800 180.400 ;
        RECT 276.400 177.800 277.200 180.400 ;
        RECT 281.200 175.800 282.000 180.400 ;
        RECT 282.800 175.800 283.600 180.400 ;
        RECT 286.000 175.800 286.800 180.400 ;
        RECT 289.200 175.800 290.000 180.400 ;
        RECT 292.400 175.800 293.200 180.400 ;
        RECT 295.600 175.800 296.400 180.400 ;
        RECT 305.200 175.800 306.000 180.400 ;
        RECT 314.800 177.800 315.600 180.400 ;
        RECT 318.000 177.800 318.800 180.400 ;
        RECT 329.200 175.800 330.000 180.400 ;
        RECT 335.600 177.800 336.400 180.400 ;
        RECT 337.200 175.800 338.000 180.400 ;
        RECT 345.200 176.600 346.000 180.400 ;
        RECT 348.400 175.800 349.200 180.400 ;
        RECT 354.800 175.800 355.600 180.400 ;
        RECT 358.000 175.800 358.800 180.400 ;
        RECT 359.600 175.800 360.400 180.400 ;
        RECT 366.000 176.600 366.800 180.400 ;
        RECT 372.400 175.800 373.200 180.400 ;
        RECT 375.600 175.800 376.400 180.400 ;
        RECT 377.200 175.800 378.000 180.400 ;
        RECT 383.600 177.800 384.400 180.400 ;
        RECT 386.800 176.000 387.600 180.400 ;
        RECT 392.400 177.800 393.200 180.400 ;
        RECT 395.600 177.800 396.600 180.400 ;
        RECT 401.200 175.800 402.000 180.400 ;
        RECT 406.000 176.600 406.800 180.400 ;
        RECT 414.000 176.600 414.800 180.400 ;
        RECT 418.400 175.000 419.200 180.400 ;
        RECT 423.600 175.400 424.400 180.400 ;
        RECT 428.400 175.800 429.200 180.400 ;
        RECT 433.800 177.800 434.800 180.400 ;
        RECT 437.200 177.800 438.000 180.400 ;
        RECT 442.800 176.000 443.600 180.400 ;
        RECT 447.600 176.600 448.400 180.400 ;
        RECT 455.600 176.600 456.400 180.400 ;
        RECT 465.200 176.600 466.000 180.400 ;
        RECT 471.600 176.600 472.400 180.400 ;
        RECT 477.600 175.000 478.400 180.400 ;
        RECT 482.800 175.400 483.600 180.400 ;
        RECT 487.600 176.000 488.400 180.400 ;
        RECT 493.200 177.800 494.000 180.400 ;
        RECT 496.400 177.800 497.400 180.400 ;
        RECT 502.000 175.800 502.800 180.400 ;
        RECT 506.800 176.600 507.600 180.400 ;
        RECT 514.800 176.600 515.600 180.400 ;
        RECT 519.600 175.400 520.400 180.400 ;
        RECT 524.800 175.000 525.600 180.400 ;
        RECT 529.200 175.400 530.000 180.400 ;
        RECT 534.400 175.000 535.200 180.400 ;
        RECT 538.800 176.600 539.600 180.400 ;
        RECT 545.200 176.600 546.000 180.400 ;
        RECT 551.600 177.800 552.400 180.400 ;
        RECT 553.200 175.800 554.000 180.400 ;
        RECT 559.600 176.600 560.400 180.400 ;
        RECT 564.400 177.800 565.200 180.400 ;
        RECT 570.800 175.800 571.600 180.400 ;
        RECT 582.000 177.800 582.800 180.400 ;
        RECT 585.200 177.800 586.000 180.400 ;
        RECT 594.800 175.800 595.600 180.400 ;
        RECT 602.800 176.600 603.600 180.400 ;
        RECT 607.600 177.800 608.400 180.400 ;
        RECT 2.800 141.600 3.600 146.200 ;
        RECT 8.200 141.600 9.200 144.200 ;
        RECT 11.600 141.600 12.400 144.200 ;
        RECT 17.200 141.600 18.000 146.000 ;
        RECT 23.600 141.600 24.400 145.400 ;
        RECT 28.400 141.600 29.200 145.400 ;
        RECT 36.400 141.600 37.200 145.400 ;
        RECT 40.800 141.600 41.600 147.000 ;
        RECT 46.000 141.600 46.800 146.600 ;
        RECT 50.400 141.600 51.200 147.000 ;
        RECT 55.600 141.600 56.400 146.600 ;
        RECT 60.400 141.600 61.200 145.400 ;
        RECT 68.400 141.600 69.200 145.400 ;
        RECT 73.200 141.600 74.000 146.200 ;
        RECT 78.600 141.600 79.600 144.200 ;
        RECT 82.000 141.600 82.800 144.200 ;
        RECT 87.600 141.600 88.400 146.000 ;
        RECT 90.800 141.600 91.600 148.200 ;
        RECT 98.800 141.600 99.600 145.400 ;
        RECT 103.600 141.600 104.400 148.200 ;
        RECT 111.600 141.600 112.400 145.400 ;
        RECT 119.600 141.600 120.400 145.400 ;
        RECT 124.400 141.600 125.200 145.400 ;
        RECT 130.800 141.600 131.600 145.400 ;
        RECT 137.200 141.600 138.000 145.400 ;
        RECT 142.000 141.600 142.800 146.200 ;
        RECT 146.800 141.600 147.800 145.600 ;
        RECT 153.000 142.200 154.000 145.600 ;
        RECT 153.000 141.600 153.800 142.200 ;
        RECT 164.400 141.600 165.200 146.200 ;
        RECT 174.000 141.600 174.800 144.200 ;
        RECT 177.200 141.600 178.000 144.200 ;
        RECT 188.400 141.600 189.200 146.200 ;
        RECT 194.800 141.600 195.600 144.200 ;
        RECT 199.600 141.600 200.400 145.400 ;
        RECT 202.800 141.600 203.600 146.200 ;
        RECT 206.000 141.600 206.800 146.200 ;
        RECT 209.200 141.600 210.000 144.200 ;
        RECT 212.400 141.600 213.200 144.200 ;
        RECT 217.200 141.600 218.000 146.200 ;
        RECT 220.400 141.600 221.200 145.400 ;
        RECT 228.400 141.600 229.200 146.200 ;
        RECT 238.000 141.600 238.800 144.200 ;
        RECT 241.200 141.600 242.000 144.200 ;
        RECT 252.400 141.600 253.200 146.200 ;
        RECT 258.800 141.600 259.600 144.200 ;
        RECT 263.600 141.600 264.400 146.200 ;
        RECT 268.400 141.600 269.200 146.200 ;
        RECT 278.000 141.600 278.800 144.200 ;
        RECT 281.200 141.600 282.000 144.200 ;
        RECT 292.400 141.600 293.200 146.200 ;
        RECT 298.800 141.600 299.600 144.200 ;
        RECT 302.000 141.600 302.800 144.200 ;
        RECT 310.000 141.600 310.800 145.400 ;
        RECT 314.800 141.600 315.600 146.200 ;
        RECT 322.800 141.600 323.600 146.200 ;
        RECT 332.400 141.600 333.200 144.200 ;
        RECT 335.600 141.600 336.400 144.200 ;
        RECT 346.800 141.600 347.600 146.200 ;
        RECT 353.200 141.600 354.000 144.200 ;
        RECT 358.000 141.600 358.800 146.200 ;
        RECT 362.800 141.600 363.600 145.400 ;
        RECT 366.000 141.600 366.800 146.200 ;
        RECT 374.000 141.600 374.800 145.400 ;
        RECT 380.400 141.600 381.200 145.400 ;
        RECT 385.200 141.600 386.000 145.400 ;
        RECT 393.200 141.600 394.000 145.400 ;
        RECT 401.200 141.600 402.000 148.200 ;
        RECT 407.600 141.600 408.400 148.200 ;
        RECT 410.800 141.600 411.600 145.400 ;
        RECT 418.800 141.600 419.600 145.400 ;
        RECT 423.200 141.600 424.000 147.000 ;
        RECT 428.400 141.600 429.200 146.600 ;
        RECT 434.800 141.600 435.600 145.400 ;
        RECT 439.600 141.600 440.400 144.200 ;
        RECT 442.800 141.600 443.600 146.600 ;
        RECT 448.000 141.600 448.800 147.000 ;
        RECT 454.000 141.600 454.800 146.200 ;
        RECT 462.000 141.600 462.800 146.000 ;
        RECT 467.600 141.600 468.400 144.200 ;
        RECT 470.800 141.600 471.800 144.200 ;
        RECT 476.400 141.600 477.200 146.200 ;
        RECT 481.200 141.600 482.000 144.200 ;
        RECT 484.400 141.600 485.200 146.600 ;
        RECT 489.600 141.600 490.400 147.000 ;
        RECT 492.400 141.600 493.200 146.200 ;
        RECT 500.400 141.600 501.200 145.400 ;
        RECT 505.200 141.600 506.000 145.400 ;
        RECT 513.200 141.600 514.000 145.400 ;
        RECT 518.000 141.600 518.800 146.000 ;
        RECT 523.600 141.600 524.400 144.200 ;
        RECT 526.800 141.600 527.800 144.200 ;
        RECT 532.400 141.600 533.200 146.200 ;
        RECT 537.200 141.600 538.000 145.400 ;
        RECT 543.600 141.600 544.400 146.000 ;
        RECT 549.200 141.600 550.000 144.200 ;
        RECT 552.400 141.600 553.400 144.200 ;
        RECT 558.000 141.600 558.800 146.200 ;
        RECT 561.200 141.600 562.000 144.200 ;
        RECT 564.400 141.600 565.200 145.800 ;
        RECT 567.600 141.600 568.400 144.200 ;
        RECT 574.000 141.600 574.800 146.200 ;
        RECT 585.200 141.600 586.000 144.200 ;
        RECT 588.400 141.600 589.200 144.200 ;
        RECT 598.000 141.600 598.800 146.200 ;
        RECT 604.400 141.600 605.200 144.200 ;
        RECT 607.600 141.600 608.400 146.200 ;
        RECT 0.400 140.400 614.000 141.600 ;
        RECT 1.200 137.800 2.000 140.400 ;
        RECT 7.600 135.800 8.400 140.400 ;
        RECT 18.800 137.800 19.600 140.400 ;
        RECT 22.000 137.800 22.800 140.400 ;
        RECT 31.600 135.800 32.400 140.400 ;
        RECT 36.400 135.800 37.200 140.400 ;
        RECT 44.400 136.600 45.200 140.400 ;
        RECT 48.800 135.000 49.600 140.400 ;
        RECT 54.000 135.400 54.800 140.400 ;
        RECT 58.800 136.600 59.600 140.400 ;
        RECT 66.800 136.600 67.600 140.400 ;
        RECT 71.600 135.800 72.400 140.400 ;
        RECT 77.000 137.800 78.000 140.400 ;
        RECT 80.400 137.800 81.200 140.400 ;
        RECT 86.000 136.000 86.800 140.400 ;
        RECT 89.200 135.800 90.000 140.400 ;
        RECT 92.400 135.800 93.200 140.400 ;
        RECT 98.800 136.600 99.600 140.400 ;
        RECT 103.600 135.800 104.400 140.400 ;
        RECT 109.000 137.800 110.000 140.400 ;
        RECT 112.400 137.800 113.200 140.400 ;
        RECT 118.000 136.000 118.800 140.400 ;
        RECT 121.200 135.800 122.000 140.400 ;
        RECT 126.000 137.800 126.800 140.400 ;
        RECT 129.200 135.800 130.000 140.400 ;
        RECT 135.600 136.600 136.400 140.400 ;
        RECT 142.000 136.600 142.800 140.400 ;
        RECT 150.000 135.800 150.800 140.400 ;
        RECT 158.000 136.600 158.800 140.400 ;
        RECT 162.800 137.800 163.600 140.400 ;
        RECT 169.200 135.800 170.000 140.400 ;
        RECT 180.400 137.800 181.200 140.400 ;
        RECT 183.600 137.800 184.400 140.400 ;
        RECT 193.200 135.800 194.000 140.400 ;
        RECT 201.200 135.800 202.000 140.400 ;
        RECT 202.800 135.800 203.600 140.400 ;
        RECT 206.000 135.800 206.800 140.400 ;
        RECT 209.200 137.800 210.000 140.400 ;
        RECT 215.600 135.800 216.400 140.400 ;
        RECT 226.800 137.800 227.600 140.400 ;
        RECT 230.000 137.800 230.800 140.400 ;
        RECT 239.600 135.800 240.400 140.400 ;
        RECT 244.400 137.800 245.200 140.400 ;
        RECT 247.600 137.800 248.400 140.400 ;
        RECT 249.200 137.800 250.000 140.400 ;
        RECT 252.400 137.800 253.200 140.400 ;
        RECT 255.600 135.800 256.400 140.400 ;
        RECT 258.800 135.800 259.600 140.400 ;
        RECT 262.000 136.600 262.800 140.400 ;
        RECT 266.800 137.800 267.600 140.400 ;
        RECT 273.200 135.800 274.000 140.400 ;
        RECT 284.400 137.800 285.200 140.400 ;
        RECT 287.600 137.800 288.400 140.400 ;
        RECT 297.200 135.800 298.000 140.400 ;
        RECT 306.800 135.800 307.600 140.400 ;
        RECT 310.000 135.800 310.800 140.400 ;
        RECT 313.200 135.800 314.000 140.400 ;
        RECT 316.400 135.800 317.200 140.400 ;
        RECT 319.600 135.800 320.400 140.400 ;
        RECT 324.400 135.800 325.200 140.400 ;
        RECT 334.000 137.800 334.800 140.400 ;
        RECT 337.200 137.800 338.000 140.400 ;
        RECT 348.400 135.800 349.200 140.400 ;
        RECT 354.800 137.800 355.600 140.400 ;
        RECT 358.000 135.800 358.800 140.400 ;
        RECT 361.200 135.800 362.000 140.400 ;
        RECT 364.400 135.800 365.200 140.400 ;
        RECT 369.200 136.600 370.000 140.400 ;
        RECT 374.000 135.800 374.800 140.400 ;
        RECT 382.000 135.800 382.800 140.400 ;
        RECT 391.600 137.800 392.400 140.400 ;
        RECT 394.800 137.800 395.600 140.400 ;
        RECT 406.000 135.800 406.800 140.400 ;
        RECT 412.400 137.800 413.200 140.400 ;
        RECT 414.000 135.800 414.800 140.400 ;
        RECT 417.200 135.800 418.000 140.400 ;
        RECT 420.400 135.800 421.200 140.400 ;
        RECT 423.600 135.800 424.400 140.400 ;
        RECT 426.800 135.800 427.600 140.400 ;
        RECT 431.600 136.600 432.400 140.400 ;
        RECT 436.400 135.800 437.200 140.400 ;
        RECT 439.600 135.800 440.400 140.400 ;
        RECT 446.000 133.800 446.800 140.400 ;
        RECT 447.600 137.800 448.400 140.400 ;
        RECT 450.800 137.800 451.600 140.400 ;
        RECT 454.200 139.800 455.000 140.400 ;
        RECT 454.000 136.400 455.000 139.800 ;
        RECT 460.200 136.400 461.200 140.400 ;
        RECT 470.000 137.800 470.800 140.400 ;
        RECT 471.600 137.800 472.400 140.400 ;
        RECT 474.800 137.800 475.600 140.400 ;
        RECT 478.000 136.600 478.800 140.400 ;
        RECT 482.800 135.800 483.600 140.400 ;
        RECT 486.000 135.800 486.800 140.400 ;
        RECT 492.400 136.600 493.200 140.400 ;
        RECT 496.800 135.000 497.600 140.400 ;
        RECT 502.000 135.400 502.800 140.400 ;
        RECT 505.200 135.800 506.000 140.400 ;
        RECT 508.400 135.800 509.200 140.400 ;
        RECT 513.200 136.600 514.000 140.400 ;
        RECT 519.600 136.000 520.400 140.400 ;
        RECT 525.200 137.800 526.000 140.400 ;
        RECT 528.400 137.800 529.400 140.400 ;
        RECT 534.000 135.800 534.800 140.400 ;
        RECT 538.800 136.600 539.600 140.400 ;
        RECT 545.200 137.800 546.000 140.400 ;
        RECT 548.400 135.800 549.200 140.400 ;
        RECT 551.600 135.800 552.400 140.400 ;
        RECT 554.800 135.800 555.600 140.400 ;
        RECT 558.000 135.800 558.800 140.400 ;
        RECT 561.200 137.800 562.000 140.400 ;
        RECT 564.400 136.600 565.200 140.400 ;
        RECT 570.800 135.400 571.600 140.400 ;
        RECT 576.000 135.000 576.800 140.400 ;
        RECT 580.400 136.600 581.200 140.400 ;
        RECT 588.400 135.800 589.200 140.400 ;
        RECT 591.600 135.800 592.400 140.400 ;
        RECT 597.000 137.800 598.000 140.400 ;
        RECT 600.400 137.800 601.200 140.400 ;
        RECT 606.000 136.000 606.800 140.400 ;
        RECT 2.800 101.600 3.600 106.200 ;
        RECT 8.200 101.600 9.200 104.200 ;
        RECT 11.600 101.600 12.400 104.200 ;
        RECT 17.200 101.600 18.000 106.000 ;
        RECT 23.600 101.600 24.400 105.400 ;
        RECT 30.000 101.600 30.800 105.400 ;
        RECT 33.200 101.600 34.000 106.200 ;
        RECT 36.400 101.600 37.200 106.200 ;
        RECT 40.800 101.600 41.600 107.000 ;
        RECT 46.000 101.600 46.800 106.600 ;
        RECT 50.800 101.600 51.600 105.400 ;
        RECT 58.800 101.600 59.600 105.400 ;
        RECT 63.200 101.600 64.000 107.000 ;
        RECT 68.400 101.600 69.200 106.600 ;
        RECT 71.600 101.600 72.400 106.200 ;
        RECT 74.800 101.600 75.600 106.200 ;
        RECT 78.000 101.600 78.800 106.200 ;
        RECT 81.200 101.600 82.000 106.200 ;
        RECT 84.400 101.600 85.200 106.200 ;
        RECT 89.200 101.600 90.000 108.200 ;
        RECT 98.800 101.600 99.600 105.400 ;
        RECT 103.600 101.600 104.400 105.400 ;
        RECT 110.000 101.600 110.800 105.400 ;
        RECT 116.400 101.600 117.200 105.400 ;
        RECT 122.800 101.600 123.600 106.200 ;
        RECT 126.000 101.600 126.800 106.200 ;
        RECT 130.800 101.600 131.600 106.200 ;
        RECT 132.400 101.600 133.200 104.200 ;
        RECT 138.800 101.600 139.600 105.400 ;
        RECT 145.200 101.600 146.000 105.400 ;
        RECT 156.400 101.600 157.200 105.400 ;
        RECT 159.600 101.600 160.400 106.200 ;
        RECT 162.800 101.600 163.600 106.200 ;
        RECT 166.000 101.600 166.800 106.200 ;
        RECT 169.200 101.600 170.000 106.200 ;
        RECT 172.400 101.600 173.200 106.200 ;
        RECT 175.600 101.600 176.400 106.600 ;
        RECT 180.800 101.600 181.600 107.000 ;
        RECT 185.200 101.600 186.000 106.600 ;
        RECT 190.400 101.600 191.200 107.000 ;
        RECT 194.800 102.200 195.800 105.600 ;
        RECT 195.000 101.600 195.800 102.200 ;
        RECT 201.000 101.600 202.000 105.600 ;
        RECT 206.000 101.600 206.800 105.800 ;
        RECT 209.200 101.600 210.000 104.200 ;
        RECT 210.800 101.600 211.600 104.200 ;
        RECT 215.000 101.600 215.800 106.200 ;
        RECT 217.200 101.600 218.000 108.200 ;
        RECT 225.200 101.600 226.000 104.200 ;
        RECT 226.800 101.600 227.600 104.200 ;
        RECT 230.000 101.600 230.800 105.800 ;
        RECT 233.200 101.600 234.000 104.200 ;
        RECT 236.400 101.600 237.200 104.200 ;
        RECT 241.200 101.600 242.000 105.400 ;
        RECT 247.600 101.600 248.400 106.200 ;
        RECT 257.200 101.600 258.000 104.200 ;
        RECT 260.400 101.600 261.200 104.200 ;
        RECT 271.600 101.600 272.400 106.200 ;
        RECT 278.000 101.600 278.800 104.200 ;
        RECT 282.800 101.600 283.600 105.400 ;
        RECT 286.000 101.600 286.800 106.200 ;
        RECT 289.200 101.600 290.000 106.200 ;
        RECT 294.000 102.200 295.000 105.600 ;
        RECT 294.200 101.600 295.000 102.200 ;
        RECT 300.200 101.600 301.200 105.600 ;
        RECT 308.400 101.600 309.200 106.200 ;
        RECT 313.200 101.600 314.000 104.200 ;
        RECT 319.600 101.600 320.400 106.200 ;
        RECT 330.800 101.600 331.600 104.200 ;
        RECT 334.000 101.600 334.800 104.200 ;
        RECT 343.600 101.600 344.400 106.200 ;
        RECT 348.400 101.600 349.200 106.200 ;
        RECT 351.600 101.600 352.400 106.200 ;
        RECT 356.400 101.600 357.200 106.200 ;
        RECT 359.600 101.600 360.400 106.200 ;
        RECT 362.800 101.600 363.600 104.200 ;
        RECT 366.000 101.600 366.800 105.400 ;
        RECT 374.000 101.600 374.800 106.200 ;
        RECT 383.600 101.600 384.400 104.200 ;
        RECT 386.800 101.600 387.600 104.200 ;
        RECT 398.000 101.600 398.800 106.200 ;
        RECT 404.400 101.600 405.200 104.200 ;
        RECT 407.600 101.600 408.400 106.000 ;
        RECT 413.200 101.600 414.000 104.200 ;
        RECT 416.400 101.600 417.400 104.200 ;
        RECT 422.000 101.600 422.800 106.200 ;
        RECT 425.200 101.600 426.000 104.200 ;
        RECT 431.600 101.600 432.400 105.400 ;
        RECT 436.000 101.600 436.800 107.000 ;
        RECT 441.200 101.600 442.000 106.600 ;
        RECT 447.600 101.600 448.400 105.400 ;
        RECT 454.000 101.600 454.800 105.400 ;
        RECT 462.000 101.600 462.800 106.200 ;
        RECT 468.400 101.600 469.200 104.200 ;
        RECT 471.600 101.600 472.400 104.200 ;
        RECT 473.200 101.600 474.000 106.200 ;
        RECT 478.000 101.600 478.800 104.200 ;
        RECT 481.200 101.600 482.000 104.200 ;
        RECT 486.000 101.600 486.800 105.400 ;
        RECT 492.400 101.600 493.200 106.200 ;
        RECT 495.600 101.600 496.400 105.400 ;
        RECT 500.400 101.600 501.200 106.200 ;
        RECT 506.800 101.600 507.600 104.200 ;
        RECT 510.000 101.600 510.800 105.400 ;
        RECT 516.000 101.600 516.800 107.000 ;
        RECT 521.200 101.600 522.000 106.600 ;
        RECT 526.000 101.600 526.800 105.400 ;
        RECT 534.000 101.600 534.800 105.400 ;
        RECT 538.800 101.600 539.600 106.000 ;
        RECT 544.400 101.600 545.200 104.200 ;
        RECT 547.600 101.600 548.600 104.200 ;
        RECT 553.200 101.600 554.000 106.200 ;
        RECT 558.000 101.600 558.800 106.200 ;
        RECT 561.200 101.600 562.000 106.200 ;
        RECT 564.400 101.600 565.200 105.400 ;
        RECT 569.200 101.600 570.000 104.200 ;
        RECT 575.600 101.600 576.400 106.200 ;
        RECT 586.800 101.600 587.600 104.200 ;
        RECT 590.000 101.600 590.800 104.200 ;
        RECT 599.600 101.600 600.400 106.200 ;
        RECT 607.600 101.600 608.400 105.400 ;
        RECT 0.400 100.400 614.000 101.600 ;
        RECT 2.800 96.000 3.600 100.400 ;
        RECT 8.400 97.800 9.200 100.400 ;
        RECT 11.600 97.800 12.600 100.400 ;
        RECT 17.200 95.800 18.000 100.400 ;
        RECT 23.600 96.600 24.400 100.400 ;
        RECT 28.400 96.600 29.200 100.400 ;
        RECT 34.400 95.000 35.200 100.400 ;
        RECT 39.600 95.400 40.400 100.400 ;
        RECT 46.000 96.600 46.800 100.400 ;
        RECT 50.800 95.800 51.600 100.400 ;
        RECT 56.200 97.800 57.200 100.400 ;
        RECT 59.600 97.800 60.400 100.400 ;
        RECT 65.200 96.000 66.000 100.400 ;
        RECT 71.600 96.600 72.400 100.400 ;
        RECT 76.400 95.400 77.200 100.400 ;
        RECT 81.600 95.000 82.400 100.400 ;
        RECT 87.600 96.600 88.400 100.400 ;
        RECT 90.800 93.800 91.600 100.400 ;
        RECT 100.400 96.600 101.200 100.400 ;
        RECT 103.600 93.800 104.400 100.400 ;
        RECT 110.000 97.800 110.800 100.400 ;
        RECT 113.200 97.800 114.000 100.400 ;
        RECT 118.000 96.600 118.800 100.400 ;
        RECT 124.400 95.800 125.200 100.400 ;
        RECT 127.200 95.000 128.000 100.400 ;
        RECT 132.400 95.400 133.200 100.400 ;
        RECT 137.200 96.600 138.000 100.400 ;
        RECT 145.200 95.800 146.000 100.400 ;
        RECT 151.600 93.800 152.400 100.400 ;
        RECT 159.600 96.000 160.400 100.400 ;
        RECT 165.200 97.800 166.000 100.400 ;
        RECT 168.400 97.800 169.400 100.400 ;
        RECT 174.000 95.800 174.800 100.400 ;
        RECT 180.400 95.800 181.200 100.400 ;
        RECT 190.000 97.800 190.800 100.400 ;
        RECT 193.200 97.800 194.000 100.400 ;
        RECT 204.400 95.800 205.200 100.400 ;
        RECT 210.800 97.800 211.600 100.400 ;
        RECT 215.600 96.600 216.400 100.400 ;
        RECT 218.800 95.800 219.600 100.400 ;
        RECT 226.800 95.800 227.600 100.400 ;
        RECT 230.600 96.000 231.400 100.400 ;
        RECT 238.000 95.800 238.800 100.400 ;
        RECT 241.200 96.600 242.000 100.400 ;
        RECT 246.000 97.800 246.800 100.400 ;
        RECT 249.200 97.800 250.000 100.400 ;
        RECT 255.600 95.800 256.400 100.400 ;
        RECT 266.800 97.800 267.600 100.400 ;
        RECT 270.000 97.800 270.800 100.400 ;
        RECT 279.600 95.800 280.400 100.400 ;
        RECT 287.600 95.800 288.400 100.400 ;
        RECT 297.200 97.800 298.000 100.400 ;
        RECT 300.400 97.800 301.200 100.400 ;
        RECT 311.600 95.800 312.400 100.400 ;
        RECT 318.000 97.800 318.800 100.400 ;
        RECT 324.400 95.800 325.200 100.400 ;
        RECT 327.600 95.800 328.400 100.400 ;
        RECT 330.800 97.800 331.600 100.400 ;
        RECT 337.200 95.800 338.000 100.400 ;
        RECT 348.400 97.800 349.200 100.400 ;
        RECT 351.600 97.800 352.400 100.400 ;
        RECT 361.200 95.800 362.000 100.400 ;
        RECT 369.200 95.800 370.000 100.400 ;
        RECT 378.800 97.800 379.600 100.400 ;
        RECT 382.000 97.800 382.800 100.400 ;
        RECT 393.200 95.800 394.000 100.400 ;
        RECT 399.600 97.800 400.400 100.400 ;
        RECT 404.400 96.600 405.200 100.400 ;
        RECT 407.600 97.800 408.400 100.400 ;
        RECT 412.400 96.600 413.200 100.400 ;
        RECT 418.400 95.000 419.200 100.400 ;
        RECT 423.600 95.400 424.400 100.400 ;
        RECT 426.800 97.800 427.600 100.400 ;
        RECT 430.000 97.800 430.800 100.400 ;
        RECT 431.600 95.800 432.400 100.400 ;
        RECT 434.800 95.800 435.600 100.400 ;
        RECT 439.600 96.600 440.400 100.400 ;
        RECT 444.400 97.800 445.200 100.400 ;
        RECT 447.600 97.800 448.400 100.400 ;
        RECT 452.400 96.600 453.200 100.400 ;
        RECT 458.800 95.800 459.600 100.400 ;
        RECT 466.800 95.400 467.600 100.400 ;
        RECT 472.000 95.000 472.800 100.400 ;
        RECT 476.400 97.800 477.200 100.400 ;
        RECT 478.000 95.800 478.800 100.400 ;
        RECT 481.200 95.800 482.000 100.400 ;
        RECT 486.000 95.800 486.800 100.400 ;
        RECT 489.200 95.800 490.000 100.400 ;
        RECT 492.400 96.600 493.200 100.400 ;
        RECT 498.800 95.400 499.600 100.400 ;
        RECT 504.000 95.000 504.800 100.400 ;
        RECT 508.400 95.800 509.200 100.400 ;
        RECT 511.600 95.800 512.400 100.400 ;
        RECT 513.200 95.800 514.000 100.400 ;
        RECT 519.600 95.400 520.400 100.400 ;
        RECT 524.800 95.000 525.600 100.400 ;
        RECT 529.200 96.600 530.000 100.400 ;
        RECT 537.200 96.600 538.000 100.400 ;
        RECT 540.400 95.800 541.200 100.400 ;
        RECT 546.800 96.000 547.600 100.400 ;
        RECT 552.400 97.800 553.200 100.400 ;
        RECT 555.600 97.800 556.600 100.400 ;
        RECT 561.200 95.800 562.000 100.400 ;
        RECT 564.400 95.800 565.200 100.400 ;
        RECT 570.800 96.600 571.600 100.400 ;
        RECT 578.800 95.800 579.600 100.400 ;
        RECT 588.400 97.800 589.200 100.400 ;
        RECT 591.600 97.800 592.400 100.400 ;
        RECT 602.800 95.800 603.600 100.400 ;
        RECT 609.200 97.800 610.000 100.400 ;
        RECT 1.200 61.600 2.000 64.200 ;
        RECT 6.000 61.600 6.800 65.400 ;
        RECT 14.000 61.600 14.800 65.400 ;
        RECT 20.400 61.600 21.200 66.200 ;
        RECT 23.200 61.600 24.000 67.000 ;
        RECT 28.400 61.600 29.200 66.600 ;
        RECT 33.200 61.600 34.000 65.400 ;
        RECT 41.200 61.600 42.000 65.400 ;
        RECT 46.000 61.600 46.800 66.200 ;
        RECT 51.400 61.600 52.400 64.200 ;
        RECT 54.800 61.600 55.600 64.200 ;
        RECT 60.400 61.600 61.200 66.000 ;
        RECT 65.200 61.600 66.000 65.400 ;
        RECT 71.600 61.600 72.400 65.400 ;
        RECT 79.600 61.600 80.400 65.400 ;
        RECT 84.400 61.600 85.200 66.600 ;
        RECT 89.600 61.600 90.400 67.000 ;
        RECT 92.400 61.600 93.200 66.200 ;
        RECT 95.600 61.600 96.400 66.200 ;
        RECT 98.800 61.600 99.600 64.200 ;
        RECT 102.000 61.600 102.800 64.200 ;
        RECT 105.200 61.600 106.000 64.200 ;
        RECT 110.000 61.600 110.800 66.000 ;
        RECT 115.600 61.600 116.400 64.200 ;
        RECT 118.800 61.600 119.800 64.200 ;
        RECT 124.400 61.600 125.200 66.200 ;
        RECT 129.200 61.600 130.000 64.200 ;
        RECT 130.800 61.600 131.600 64.200 ;
        RECT 135.600 61.600 136.400 66.200 ;
        RECT 138.800 61.600 139.600 66.200 ;
        RECT 142.000 61.600 142.800 65.400 ;
        RECT 150.000 61.600 150.800 65.400 ;
        RECT 159.600 61.600 160.400 66.200 ;
        RECT 165.000 61.600 166.000 64.200 ;
        RECT 168.400 61.600 169.200 64.200 ;
        RECT 174.000 61.600 174.800 66.000 ;
        RECT 178.800 61.600 179.600 65.400 ;
        RECT 186.800 61.600 187.600 65.400 ;
        RECT 191.600 61.600 192.400 66.600 ;
        RECT 196.800 61.600 197.600 67.000 ;
        RECT 202.800 61.600 203.600 66.200 ;
        RECT 207.600 61.600 208.400 66.200 ;
        RECT 217.200 61.600 218.000 64.200 ;
        RECT 220.400 61.600 221.200 64.200 ;
        RECT 231.600 61.600 232.400 66.200 ;
        RECT 238.000 61.600 238.800 64.200 ;
        RECT 242.800 61.600 243.600 65.400 ;
        RECT 247.600 61.600 248.400 65.400 ;
        RECT 252.400 61.600 253.200 66.200 ;
        RECT 257.200 61.600 258.000 64.200 ;
        RECT 263.600 61.600 264.400 66.200 ;
        RECT 274.800 61.600 275.600 64.200 ;
        RECT 278.000 61.600 278.800 64.200 ;
        RECT 287.600 61.600 288.400 66.200 ;
        RECT 292.400 61.600 293.200 66.200 ;
        RECT 302.000 61.600 302.800 64.200 ;
        RECT 308.400 61.600 309.200 66.200 ;
        RECT 319.600 61.600 320.400 64.200 ;
        RECT 322.800 61.600 323.600 64.200 ;
        RECT 332.400 61.600 333.200 66.200 ;
        RECT 338.800 61.600 339.600 65.400 ;
        RECT 345.200 62.200 346.200 65.600 ;
        RECT 345.400 61.600 346.200 62.200 ;
        RECT 351.400 61.600 352.400 65.600 ;
        RECT 358.000 61.600 358.800 65.400 ;
        RECT 361.200 61.600 362.000 66.200 ;
        RECT 366.000 61.600 366.800 64.200 ;
        RECT 369.200 61.600 370.000 65.800 ;
        RECT 372.400 61.600 373.200 64.200 ;
        RECT 375.600 61.600 376.400 64.200 ;
        RECT 378.800 61.600 379.600 65.400 ;
        RECT 383.600 61.600 384.400 66.200 ;
        RECT 390.000 61.600 390.800 65.400 ;
        RECT 396.400 62.200 397.400 65.600 ;
        RECT 396.600 61.600 397.400 62.200 ;
        RECT 402.600 61.600 403.600 65.600 ;
        RECT 406.000 61.600 406.800 66.200 ;
        RECT 410.800 61.600 411.600 65.400 ;
        RECT 417.200 61.600 418.000 65.400 ;
        RECT 425.200 61.600 426.000 66.200 ;
        RECT 426.800 61.600 427.600 68.200 ;
        RECT 433.200 61.600 434.000 66.200 ;
        RECT 436.400 61.600 437.200 66.200 ;
        RECT 441.200 61.600 442.000 65.400 ;
        RECT 449.200 61.600 450.000 65.400 ;
        RECT 455.600 61.600 456.400 65.400 ;
        RECT 465.200 61.600 466.000 66.000 ;
        RECT 470.800 61.600 471.600 64.200 ;
        RECT 474.000 61.600 475.000 64.200 ;
        RECT 479.600 61.600 480.400 66.200 ;
        RECT 484.400 61.600 485.200 65.400 ;
        RECT 492.400 61.600 493.200 65.400 ;
        RECT 497.200 61.600 498.000 65.400 ;
        RECT 505.200 61.600 506.000 65.400 ;
        RECT 510.000 61.600 510.800 65.400 ;
        RECT 516.400 61.600 517.200 66.000 ;
        RECT 522.000 61.600 522.800 64.200 ;
        RECT 525.200 61.600 526.200 64.200 ;
        RECT 530.800 61.600 531.600 66.200 ;
        RECT 535.600 61.600 536.400 65.400 ;
        RECT 540.400 61.600 541.200 66.200 ;
        RECT 548.400 61.600 549.200 66.200 ;
        RECT 551.600 61.600 552.400 66.200 ;
        RECT 554.800 61.600 555.600 66.200 ;
        RECT 558.000 61.600 558.800 65.400 ;
        RECT 564.400 61.600 565.200 66.600 ;
        RECT 569.600 61.600 570.400 67.000 ;
        RECT 575.600 61.600 576.400 65.400 ;
        RECT 580.400 61.600 581.200 66.200 ;
        RECT 585.800 61.600 586.800 64.200 ;
        RECT 589.200 61.600 590.000 64.200 ;
        RECT 594.800 61.600 595.600 66.000 ;
        RECT 598.000 61.600 598.800 66.200 ;
        RECT 606.000 61.600 606.800 65.400 ;
        RECT 0.400 60.400 614.000 61.600 ;
        RECT 4.400 55.800 5.200 60.400 ;
        RECT 14.000 57.800 14.800 60.400 ;
        RECT 17.200 57.800 18.000 60.400 ;
        RECT 28.400 55.800 29.200 60.400 ;
        RECT 34.800 57.800 35.600 60.400 ;
        RECT 38.000 56.600 38.800 60.400 ;
        RECT 46.000 55.800 46.800 60.400 ;
        RECT 47.600 55.800 48.400 60.400 ;
        RECT 50.800 55.800 51.600 60.400 ;
        RECT 54.000 55.800 54.800 60.400 ;
        RECT 57.200 55.800 58.000 60.400 ;
        RECT 60.400 55.800 61.200 60.400 ;
        RECT 63.200 55.000 64.000 60.400 ;
        RECT 68.400 55.400 69.200 60.400 ;
        RECT 74.800 55.800 75.600 60.400 ;
        RECT 78.000 55.400 78.800 60.400 ;
        RECT 83.200 55.000 84.000 60.400 ;
        RECT 87.200 55.000 88.000 60.400 ;
        RECT 92.400 55.400 93.200 60.400 ;
        RECT 95.600 57.800 96.400 60.400 ;
        RECT 98.800 55.800 99.600 60.400 ;
        RECT 102.000 55.800 102.800 60.400 ;
        RECT 105.200 55.800 106.000 60.400 ;
        RECT 108.400 55.800 109.200 60.400 ;
        RECT 111.600 55.800 112.400 60.400 ;
        RECT 114.400 55.000 115.200 60.400 ;
        RECT 119.600 55.400 120.400 60.400 ;
        RECT 124.400 55.400 125.200 60.400 ;
        RECT 129.600 55.000 130.400 60.400 ;
        RECT 132.400 55.800 133.200 60.400 ;
        RECT 135.600 55.800 136.400 60.400 ;
        RECT 140.000 55.000 140.800 60.400 ;
        RECT 145.200 55.400 146.000 60.400 ;
        RECT 154.800 56.600 155.600 60.400 ;
        RECT 162.800 56.600 163.600 60.400 ;
        RECT 166.000 55.800 166.800 60.400 ;
        RECT 169.200 55.800 170.000 60.400 ;
        RECT 172.400 55.800 173.200 60.400 ;
        RECT 175.600 55.800 176.400 60.400 ;
        RECT 178.800 55.800 179.600 60.400 ;
        RECT 183.600 55.800 184.400 60.400 ;
        RECT 193.200 57.800 194.000 60.400 ;
        RECT 196.400 57.800 197.200 60.400 ;
        RECT 207.600 55.800 208.400 60.400 ;
        RECT 214.000 57.800 214.800 60.400 ;
        RECT 215.600 55.800 216.400 60.400 ;
        RECT 222.000 57.800 222.800 60.400 ;
        RECT 223.600 55.800 224.400 60.400 ;
        RECT 228.400 55.800 229.200 60.400 ;
        RECT 236.400 56.600 237.200 60.400 ;
        RECT 241.200 57.800 242.000 60.400 ;
        RECT 246.000 55.800 246.800 60.400 ;
        RECT 255.600 57.800 256.400 60.400 ;
        RECT 258.800 57.800 259.600 60.400 ;
        RECT 270.000 55.800 270.800 60.400 ;
        RECT 276.400 57.800 277.200 60.400 ;
        RECT 279.600 56.600 280.400 60.400 ;
        RECT 287.600 56.600 288.400 60.400 ;
        RECT 298.800 55.800 299.600 60.400 ;
        RECT 308.400 57.800 309.200 60.400 ;
        RECT 311.600 57.800 312.400 60.400 ;
        RECT 322.800 55.800 323.600 60.400 ;
        RECT 329.200 57.800 330.000 60.400 ;
        RECT 332.000 55.000 332.800 60.400 ;
        RECT 337.200 55.400 338.000 60.400 ;
        RECT 340.400 55.800 341.200 60.400 ;
        RECT 348.400 55.800 349.200 60.400 ;
        RECT 350.600 55.800 351.400 60.400 ;
        RECT 354.800 57.800 355.600 60.400 ;
        RECT 358.000 56.600 358.800 60.400 ;
        RECT 365.400 56.000 366.200 60.400 ;
        RECT 369.200 57.800 370.000 60.400 ;
        RECT 375.600 55.800 376.400 60.400 ;
        RECT 385.200 57.800 386.000 60.400 ;
        RECT 388.400 57.800 389.200 60.400 ;
        RECT 399.600 55.800 400.400 60.400 ;
        RECT 406.000 57.800 406.800 60.400 ;
        RECT 409.200 55.800 410.000 60.400 ;
        RECT 414.600 57.800 415.600 60.400 ;
        RECT 418.000 57.800 418.800 60.400 ;
        RECT 423.600 56.000 424.400 60.400 ;
        RECT 426.800 57.800 427.600 60.400 ;
        RECT 431.600 56.600 432.400 60.400 ;
        RECT 439.600 56.600 440.400 60.400 ;
        RECT 446.000 56.600 446.800 60.400 ;
        RECT 450.400 55.000 451.200 60.400 ;
        RECT 455.600 55.400 456.400 60.400 ;
        RECT 466.800 56.600 467.600 60.400 ;
        RECT 471.600 57.800 472.400 60.400 ;
        RECT 474.800 55.400 475.600 60.400 ;
        RECT 480.000 55.000 480.800 60.400 ;
        RECT 484.400 55.800 485.200 60.400 ;
        RECT 489.800 57.800 490.800 60.400 ;
        RECT 493.200 57.800 494.000 60.400 ;
        RECT 498.800 56.000 499.600 60.400 ;
        RECT 502.000 57.800 502.800 60.400 ;
        RECT 506.800 55.400 507.600 60.400 ;
        RECT 512.000 55.000 512.800 60.400 ;
        RECT 514.800 55.800 515.600 60.400 ;
        RECT 518.000 55.800 518.800 60.400 ;
        RECT 522.400 55.000 523.200 60.400 ;
        RECT 527.600 55.400 528.400 60.400 ;
        RECT 532.400 56.600 533.200 60.400 ;
        RECT 540.400 56.600 541.200 60.400 ;
        RECT 545.200 56.000 546.000 60.400 ;
        RECT 550.800 57.800 551.600 60.400 ;
        RECT 554.000 57.800 555.000 60.400 ;
        RECT 559.600 55.800 560.400 60.400 ;
        RECT 562.800 55.800 563.600 60.400 ;
        RECT 566.000 55.800 566.800 60.400 ;
        RECT 569.200 55.800 570.000 60.400 ;
        RECT 572.400 55.800 573.200 60.400 ;
        RECT 575.600 55.800 576.400 60.400 ;
        RECT 577.200 57.800 578.000 60.400 ;
        RECT 583.600 55.800 584.400 60.400 ;
        RECT 594.800 57.800 595.600 60.400 ;
        RECT 598.000 57.800 598.800 60.400 ;
        RECT 607.600 55.800 608.400 60.400 ;
        RECT 2.800 21.600 3.600 26.200 ;
        RECT 9.200 21.600 10.000 26.200 ;
        RECT 18.800 21.600 19.600 24.200 ;
        RECT 22.000 21.600 22.800 24.200 ;
        RECT 33.200 21.600 34.000 26.200 ;
        RECT 39.600 21.600 40.400 24.200 ;
        RECT 44.400 21.600 45.200 25.400 ;
        RECT 49.200 21.600 50.000 24.200 ;
        RECT 52.400 21.600 53.200 25.400 ;
        RECT 60.400 21.600 61.200 25.400 ;
        RECT 65.200 21.600 66.000 26.000 ;
        RECT 70.800 21.600 71.600 24.200 ;
        RECT 74.000 21.600 75.000 24.200 ;
        RECT 79.600 21.600 80.400 26.200 ;
        RECT 84.400 21.600 85.200 25.400 ;
        RECT 92.400 21.600 93.200 25.400 ;
        RECT 97.200 21.600 98.000 26.200 ;
        RECT 102.600 21.600 103.600 24.200 ;
        RECT 106.000 21.600 106.800 24.200 ;
        RECT 111.600 21.600 112.400 26.000 ;
        RECT 116.400 21.600 117.200 25.400 ;
        RECT 124.400 21.600 125.200 25.400 ;
        RECT 129.200 21.600 130.000 25.400 ;
        RECT 137.200 21.600 138.000 25.400 ;
        RECT 142.000 21.600 142.800 26.000 ;
        RECT 147.600 21.600 148.400 24.200 ;
        RECT 150.800 21.600 151.800 24.200 ;
        RECT 156.400 21.600 157.200 26.200 ;
        RECT 164.400 21.600 165.200 24.200 ;
        RECT 169.200 21.600 170.000 25.400 ;
        RECT 177.200 21.600 178.000 26.200 ;
        RECT 178.800 21.600 179.600 24.200 ;
        RECT 185.200 21.600 186.000 26.200 ;
        RECT 196.400 21.600 197.200 24.200 ;
        RECT 199.600 21.600 200.400 24.200 ;
        RECT 209.200 21.600 210.000 26.200 ;
        RECT 215.600 21.600 216.400 24.200 ;
        RECT 220.400 21.600 221.200 25.400 ;
        RECT 226.800 21.600 227.600 25.400 ;
        RECT 231.600 21.600 232.400 24.200 ;
        RECT 236.400 21.600 237.200 26.200 ;
        RECT 246.000 21.600 246.800 24.200 ;
        RECT 249.200 21.600 250.000 24.200 ;
        RECT 260.400 21.600 261.200 26.200 ;
        RECT 266.800 21.600 267.600 24.200 ;
        RECT 268.400 21.600 269.200 24.200 ;
        RECT 274.800 21.600 275.600 26.200 ;
        RECT 284.400 21.600 285.200 24.200 ;
        RECT 287.600 21.600 288.400 24.200 ;
        RECT 298.800 21.600 299.600 26.200 ;
        RECT 305.200 21.600 306.000 24.200 ;
        RECT 311.600 21.600 312.400 24.200 ;
        RECT 316.400 21.600 317.400 25.600 ;
        RECT 322.600 22.200 323.600 25.600 ;
        RECT 322.600 21.600 323.400 22.200 ;
        RECT 327.600 21.600 328.400 26.600 ;
        RECT 332.800 21.600 333.600 27.000 ;
        RECT 337.200 22.200 338.200 25.600 ;
        RECT 337.400 21.600 338.200 22.200 ;
        RECT 343.400 21.600 344.400 25.600 ;
        RECT 346.800 21.600 347.600 28.200 ;
        RECT 353.200 21.600 354.000 24.200 ;
        RECT 356.400 21.600 357.200 24.200 ;
        RECT 358.000 21.600 358.800 24.200 ;
        RECT 364.400 21.600 365.200 26.200 ;
        RECT 375.600 21.600 376.400 24.200 ;
        RECT 378.800 21.600 379.600 24.200 ;
        RECT 388.400 21.600 389.200 26.200 ;
        RECT 393.200 21.600 394.000 26.200 ;
        RECT 396.400 21.600 397.200 26.200 ;
        RECT 399.600 21.600 400.400 26.200 ;
        RECT 402.800 21.600 403.600 26.200 ;
        RECT 406.000 21.600 406.800 26.200 ;
        RECT 407.600 21.600 408.400 26.200 ;
        RECT 410.800 21.600 411.600 26.200 ;
        RECT 414.000 21.600 414.800 26.200 ;
        RECT 417.200 21.600 418.000 26.200 ;
        RECT 420.400 21.600 421.200 26.200 ;
        RECT 423.600 21.600 424.400 25.400 ;
        RECT 433.200 21.600 434.000 28.200 ;
        RECT 438.000 21.600 438.800 25.400 ;
        RECT 446.000 21.600 446.800 28.200 ;
        RECT 450.800 21.600 451.600 25.400 ;
        RECT 460.400 21.600 461.200 26.200 ;
        RECT 465.800 21.600 466.800 24.200 ;
        RECT 469.200 21.600 470.000 24.200 ;
        RECT 474.800 21.600 475.600 26.000 ;
        RECT 479.600 21.600 480.400 25.400 ;
        RECT 487.600 21.600 488.400 25.400 ;
        RECT 492.400 21.600 493.200 26.200 ;
        RECT 497.800 21.600 498.800 24.200 ;
        RECT 501.200 21.600 502.000 24.200 ;
        RECT 506.800 21.600 507.600 26.000 ;
        RECT 511.600 21.600 512.400 25.400 ;
        RECT 519.600 21.600 520.400 25.400 ;
        RECT 522.800 21.600 523.600 26.200 ;
        RECT 526.000 21.600 526.800 26.200 ;
        RECT 529.200 21.600 530.000 26.200 ;
        RECT 532.400 21.600 533.200 26.200 ;
        RECT 535.600 21.600 536.400 26.200 ;
        RECT 538.800 21.600 539.600 24.200 ;
        RECT 543.600 21.600 544.400 25.400 ;
        RECT 548.400 21.600 549.200 25.400 ;
        RECT 556.400 21.600 557.200 25.400 ;
        RECT 562.800 21.600 563.600 25.400 ;
        RECT 567.600 21.600 568.400 24.200 ;
        RECT 569.200 21.600 570.000 24.200 ;
        RECT 575.600 21.600 576.400 26.200 ;
        RECT 586.800 21.600 587.600 24.200 ;
        RECT 590.000 21.600 590.800 24.200 ;
        RECT 599.600 21.600 600.400 26.200 ;
        RECT 606.000 21.600 606.800 24.200 ;
        RECT 609.200 21.600 610.000 26.200 ;
        RECT 0.400 20.400 614.000 21.600 ;
        RECT 4.400 15.800 5.200 20.400 ;
        RECT 14.000 17.800 14.800 20.400 ;
        RECT 17.200 17.800 18.000 20.400 ;
        RECT 28.400 15.800 29.200 20.400 ;
        RECT 34.800 17.800 35.600 20.400 ;
        RECT 38.000 16.600 38.800 20.400 ;
        RECT 46.000 16.600 46.800 20.400 ;
        RECT 50.800 17.800 51.600 20.400 ;
        RECT 54.000 15.800 54.800 20.400 ;
        RECT 59.400 17.800 60.400 20.400 ;
        RECT 62.800 17.800 63.600 20.400 ;
        RECT 68.400 16.000 69.200 20.400 ;
        RECT 71.600 15.800 72.400 20.400 ;
        RECT 74.800 15.800 75.600 20.400 ;
        RECT 79.600 16.600 80.400 20.400 ;
        RECT 87.600 16.600 88.400 20.400 ;
        RECT 92.400 16.000 93.200 20.400 ;
        RECT 98.000 17.800 98.800 20.400 ;
        RECT 101.200 17.800 102.200 20.400 ;
        RECT 106.800 15.800 107.600 20.400 ;
        RECT 111.600 16.000 112.400 20.400 ;
        RECT 117.200 17.800 118.000 20.400 ;
        RECT 120.400 17.800 121.400 20.400 ;
        RECT 126.000 15.800 126.800 20.400 ;
        RECT 129.200 15.800 130.000 20.400 ;
        RECT 132.400 15.800 133.200 20.400 ;
        RECT 137.200 15.800 138.000 20.400 ;
        RECT 145.200 17.800 146.000 20.400 ;
        RECT 151.600 15.800 152.400 20.400 ;
        RECT 162.800 17.800 163.600 20.400 ;
        RECT 166.000 17.800 166.800 20.400 ;
        RECT 175.600 15.800 176.400 20.400 ;
        RECT 183.600 15.800 184.400 20.400 ;
        RECT 193.200 17.800 194.000 20.400 ;
        RECT 196.400 17.800 197.200 20.400 ;
        RECT 207.600 15.800 208.400 20.400 ;
        RECT 214.000 17.800 214.800 20.400 ;
        RECT 217.200 15.800 218.000 20.400 ;
        RECT 223.600 15.800 224.400 20.400 ;
        RECT 233.200 17.800 234.000 20.400 ;
        RECT 236.400 17.800 237.200 20.400 ;
        RECT 247.600 15.800 248.400 20.400 ;
        RECT 254.000 17.800 254.800 20.400 ;
        RECT 257.200 15.800 258.000 20.400 ;
        RECT 262.000 15.800 262.800 20.400 ;
        RECT 266.800 15.800 267.600 20.400 ;
        RECT 273.200 15.800 274.000 20.400 ;
        RECT 282.800 17.800 283.600 20.400 ;
        RECT 286.000 17.800 286.800 20.400 ;
        RECT 297.200 15.800 298.000 20.400 ;
        RECT 303.600 17.800 304.400 20.400 ;
        RECT 311.600 15.800 312.400 20.400 ;
        RECT 318.000 15.800 318.800 20.400 ;
        RECT 327.600 17.800 328.400 20.400 ;
        RECT 330.800 17.800 331.600 20.400 ;
        RECT 342.000 15.800 342.800 20.400 ;
        RECT 348.400 17.800 349.200 20.400 ;
        RECT 350.000 17.800 350.800 20.400 ;
        RECT 353.200 16.200 354.000 20.400 ;
        RECT 356.400 17.800 357.200 20.400 ;
        RECT 359.600 17.800 360.400 20.400 ;
        RECT 362.800 17.800 363.600 20.400 ;
        RECT 367.600 15.800 368.400 20.400 ;
        RECT 377.200 17.800 378.000 20.400 ;
        RECT 380.400 17.800 381.200 20.400 ;
        RECT 391.600 15.800 392.400 20.400 ;
        RECT 398.000 17.800 398.800 20.400 ;
        RECT 401.200 15.800 402.000 20.400 ;
        RECT 406.000 15.800 406.800 20.400 ;
        RECT 411.400 17.800 412.400 20.400 ;
        RECT 414.800 17.800 415.600 20.400 ;
        RECT 420.400 16.000 421.200 20.400 ;
        RECT 425.200 15.400 426.000 20.400 ;
        RECT 430.400 15.000 431.200 20.400 ;
        RECT 434.800 16.000 435.600 20.400 ;
        RECT 440.400 17.800 441.200 20.400 ;
        RECT 443.600 17.800 444.600 20.400 ;
        RECT 449.200 15.800 450.000 20.400 ;
        RECT 455.600 16.600 456.400 20.400 ;
        RECT 465.200 15.400 466.000 20.400 ;
        RECT 470.400 15.000 471.200 20.400 ;
        RECT 474.400 15.000 475.200 20.400 ;
        RECT 479.600 15.400 480.400 20.400 ;
        RECT 484.400 16.600 485.200 20.400 ;
        RECT 492.400 16.600 493.200 20.400 ;
        RECT 497.200 15.800 498.000 20.400 ;
        RECT 502.600 17.800 503.600 20.400 ;
        RECT 506.000 17.800 506.800 20.400 ;
        RECT 511.600 16.000 512.400 20.400 ;
        RECT 516.000 15.000 516.800 20.400 ;
        RECT 521.200 15.400 522.000 20.400 ;
        RECT 526.000 16.600 526.800 20.400 ;
        RECT 534.000 16.600 534.800 20.400 ;
        RECT 537.200 15.800 538.000 20.400 ;
        RECT 540.400 15.800 541.200 20.400 ;
        RECT 545.200 16.000 546.000 20.400 ;
        RECT 550.800 17.800 551.600 20.400 ;
        RECT 554.000 17.800 555.000 20.400 ;
        RECT 559.600 15.800 560.400 20.400 ;
        RECT 564.400 17.800 565.200 20.400 ;
        RECT 567.600 16.600 568.400 20.400 ;
        RECT 572.400 17.800 573.200 20.400 ;
        RECT 578.800 15.800 579.600 20.400 ;
        RECT 590.000 17.800 590.800 20.400 ;
        RECT 593.200 17.800 594.000 20.400 ;
        RECT 602.800 15.800 603.600 20.400 ;
        RECT 609.200 17.800 610.000 20.400 ;
      LAYER via1 ;
        RECT 303.800 540.600 304.600 541.400 ;
        RECT 305.200 540.600 306.000 541.400 ;
        RECT 306.600 540.600 307.400 541.400 ;
        RECT 303.800 500.600 304.600 501.400 ;
        RECT 305.200 500.600 306.000 501.400 ;
        RECT 306.600 500.600 307.400 501.400 ;
        RECT 303.800 460.600 304.600 461.400 ;
        RECT 305.200 460.600 306.000 461.400 ;
        RECT 306.600 460.600 307.400 461.400 ;
        RECT 303.800 420.600 304.600 421.400 ;
        RECT 305.200 420.600 306.000 421.400 ;
        RECT 306.600 420.600 307.400 421.400 ;
        RECT 303.800 380.600 304.600 381.400 ;
        RECT 305.200 380.600 306.000 381.400 ;
        RECT 306.600 380.600 307.400 381.400 ;
        RECT 303.800 340.600 304.600 341.400 ;
        RECT 305.200 340.600 306.000 341.400 ;
        RECT 306.600 340.600 307.400 341.400 ;
        RECT 319.600 329.600 320.400 330.400 ;
        RECT 303.800 300.600 304.600 301.400 ;
        RECT 305.200 300.600 306.000 301.400 ;
        RECT 306.600 300.600 307.400 301.400 ;
        RECT 198.000 299.600 198.800 300.400 ;
        RECT 172.400 267.600 173.200 268.400 ;
        RECT 303.800 260.600 304.600 261.400 ;
        RECT 305.200 260.600 306.000 261.400 ;
        RECT 306.600 260.600 307.400 261.400 ;
        RECT 295.600 257.600 296.400 258.400 ;
        RECT 311.600 257.600 312.400 258.400 ;
        RECT 303.800 220.600 304.600 221.400 ;
        RECT 305.200 220.600 306.000 221.400 ;
        RECT 306.600 220.600 307.400 221.400 ;
        RECT 303.800 180.600 304.600 181.400 ;
        RECT 305.200 180.600 306.000 181.400 ;
        RECT 306.600 180.600 307.400 181.400 ;
        RECT 303.800 140.600 304.600 141.400 ;
        RECT 305.200 140.600 306.000 141.400 ;
        RECT 306.600 140.600 307.400 141.400 ;
        RECT 303.800 100.600 304.600 101.400 ;
        RECT 305.200 100.600 306.000 101.400 ;
        RECT 306.600 100.600 307.400 101.400 ;
        RECT 303.800 60.600 304.600 61.400 ;
        RECT 305.200 60.600 306.000 61.400 ;
        RECT 306.600 60.600 307.400 61.400 ;
        RECT 303.800 20.600 304.600 21.400 ;
        RECT 305.200 20.600 306.000 21.400 ;
        RECT 306.600 20.600 307.400 21.400 ;
      LAYER metal2 ;
        RECT 303.200 540.600 308.000 541.400 ;
        RECT 303.200 500.600 308.000 501.400 ;
        RECT 303.200 460.600 308.000 461.400 ;
        RECT 303.200 420.600 308.000 421.400 ;
        RECT 303.200 380.600 308.000 381.400 ;
        RECT 319.600 341.600 320.400 342.400 ;
        RECT 303.200 340.600 308.000 341.400 ;
        RECT 319.700 330.400 320.300 341.600 ;
        RECT 319.600 329.600 320.400 330.400 ;
        RECT 198.000 311.600 198.800 312.400 ;
        RECT 198.100 300.400 198.700 311.600 ;
        RECT 303.200 300.600 308.000 301.400 ;
        RECT 198.000 299.600 198.800 300.400 ;
        RECT 172.400 267.600 173.200 268.400 ;
        RECT 172.500 258.400 173.100 267.600 ;
        RECT 326.000 261.600 326.800 262.400 ;
        RECT 303.200 260.600 308.000 261.400 ;
        RECT 172.400 257.600 173.200 258.400 ;
        RECT 295.600 257.600 296.400 258.400 ;
        RECT 311.600 258.300 312.400 258.400 ;
        RECT 310.100 257.700 312.400 258.300 ;
        RECT 295.700 252.400 296.300 257.600 ;
        RECT 310.100 254.400 310.700 257.700 ;
        RECT 311.600 257.600 312.400 257.700 ;
        RECT 326.100 254.400 326.700 261.600 ;
        RECT 310.000 253.600 310.800 254.400 ;
        RECT 326.000 253.600 326.800 254.400 ;
        RECT 295.600 251.600 296.400 252.400 ;
        RECT 303.200 220.600 308.000 221.400 ;
        RECT 303.200 180.600 308.000 181.400 ;
        RECT 303.200 140.600 308.000 141.400 ;
        RECT 303.200 100.600 308.000 101.400 ;
        RECT 303.200 60.600 308.000 61.400 ;
        RECT 303.200 20.600 308.000 21.400 ;
      LAYER via2 ;
        RECT 303.800 540.600 304.600 541.400 ;
        RECT 305.200 540.600 306.000 541.400 ;
        RECT 306.600 540.600 307.400 541.400 ;
        RECT 303.800 500.600 304.600 501.400 ;
        RECT 305.200 500.600 306.000 501.400 ;
        RECT 306.600 500.600 307.400 501.400 ;
        RECT 303.800 460.600 304.600 461.400 ;
        RECT 305.200 460.600 306.000 461.400 ;
        RECT 306.600 460.600 307.400 461.400 ;
        RECT 303.800 420.600 304.600 421.400 ;
        RECT 305.200 420.600 306.000 421.400 ;
        RECT 306.600 420.600 307.400 421.400 ;
        RECT 303.800 380.600 304.600 381.400 ;
        RECT 305.200 380.600 306.000 381.400 ;
        RECT 306.600 380.600 307.400 381.400 ;
        RECT 303.800 340.600 304.600 341.400 ;
        RECT 305.200 340.600 306.000 341.400 ;
        RECT 306.600 340.600 307.400 341.400 ;
        RECT 303.800 300.600 304.600 301.400 ;
        RECT 305.200 300.600 306.000 301.400 ;
        RECT 306.600 300.600 307.400 301.400 ;
        RECT 303.800 260.600 304.600 261.400 ;
        RECT 305.200 260.600 306.000 261.400 ;
        RECT 306.600 260.600 307.400 261.400 ;
        RECT 303.800 220.600 304.600 221.400 ;
        RECT 305.200 220.600 306.000 221.400 ;
        RECT 306.600 220.600 307.400 221.400 ;
        RECT 303.800 180.600 304.600 181.400 ;
        RECT 305.200 180.600 306.000 181.400 ;
        RECT 306.600 180.600 307.400 181.400 ;
        RECT 303.800 140.600 304.600 141.400 ;
        RECT 305.200 140.600 306.000 141.400 ;
        RECT 306.600 140.600 307.400 141.400 ;
        RECT 303.800 100.600 304.600 101.400 ;
        RECT 305.200 100.600 306.000 101.400 ;
        RECT 306.600 100.600 307.400 101.400 ;
        RECT 303.800 60.600 304.600 61.400 ;
        RECT 305.200 60.600 306.000 61.400 ;
        RECT 306.600 60.600 307.400 61.400 ;
        RECT 303.800 20.600 304.600 21.400 ;
        RECT 305.200 20.600 306.000 21.400 ;
        RECT 306.600 20.600 307.400 21.400 ;
      LAYER metal3 ;
        RECT 303.200 540.400 308.000 541.600 ;
        RECT 303.200 500.400 308.000 501.600 ;
        RECT 303.200 460.400 308.000 461.600 ;
        RECT 303.200 420.400 308.000 421.600 ;
        RECT 303.200 380.400 308.000 381.600 ;
        RECT 303.200 340.400 308.000 341.600 ;
        RECT 303.200 300.400 308.000 301.600 ;
        RECT 303.200 260.400 308.000 261.600 ;
        RECT 303.200 220.400 308.000 221.600 ;
        RECT 303.200 180.400 308.000 181.600 ;
        RECT 303.200 140.400 308.000 141.600 ;
        RECT 303.200 100.400 308.000 101.600 ;
        RECT 303.200 60.400 308.000 61.600 ;
        RECT 303.200 20.400 308.000 21.600 ;
      LAYER via3 ;
        RECT 303.600 540.600 304.400 541.400 ;
        RECT 305.200 540.600 306.000 541.400 ;
        RECT 306.800 540.600 307.600 541.400 ;
        RECT 303.600 500.600 304.400 501.400 ;
        RECT 305.200 500.600 306.000 501.400 ;
        RECT 306.800 500.600 307.600 501.400 ;
        RECT 303.600 460.600 304.400 461.400 ;
        RECT 305.200 460.600 306.000 461.400 ;
        RECT 306.800 460.600 307.600 461.400 ;
        RECT 303.600 420.600 304.400 421.400 ;
        RECT 305.200 420.600 306.000 421.400 ;
        RECT 306.800 420.600 307.600 421.400 ;
        RECT 303.600 380.600 304.400 381.400 ;
        RECT 305.200 380.600 306.000 381.400 ;
        RECT 306.800 380.600 307.600 381.400 ;
        RECT 303.600 340.600 304.400 341.400 ;
        RECT 305.200 340.600 306.000 341.400 ;
        RECT 306.800 340.600 307.600 341.400 ;
        RECT 303.600 300.600 304.400 301.400 ;
        RECT 305.200 300.600 306.000 301.400 ;
        RECT 306.800 300.600 307.600 301.400 ;
        RECT 303.600 260.600 304.400 261.400 ;
        RECT 305.200 260.600 306.000 261.400 ;
        RECT 306.800 260.600 307.600 261.400 ;
        RECT 303.600 220.600 304.400 221.400 ;
        RECT 305.200 220.600 306.000 221.400 ;
        RECT 306.800 220.600 307.600 221.400 ;
        RECT 303.600 180.600 304.400 181.400 ;
        RECT 305.200 180.600 306.000 181.400 ;
        RECT 306.800 180.600 307.600 181.400 ;
        RECT 303.600 140.600 304.400 141.400 ;
        RECT 305.200 140.600 306.000 141.400 ;
        RECT 306.800 140.600 307.600 141.400 ;
        RECT 303.600 100.600 304.400 101.400 ;
        RECT 305.200 100.600 306.000 101.400 ;
        RECT 306.800 100.600 307.600 101.400 ;
        RECT 303.600 60.600 304.400 61.400 ;
        RECT 305.200 60.600 306.000 61.400 ;
        RECT 306.800 60.600 307.600 61.400 ;
        RECT 303.600 20.600 304.400 21.400 ;
        RECT 305.200 20.600 306.000 21.400 ;
        RECT 306.800 20.600 307.600 21.400 ;
      LAYER metal4 ;
        RECT 303.200 -4.000 308.000 564.000 ;
    END
  END gnd
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 273.000 372.400 273.800 373.200 ;
        RECT 414.200 372.400 415.000 373.200 ;
        RECT 273.000 371.600 274.000 372.400 ;
        RECT 414.000 371.600 415.000 372.400 ;
        RECT 41.000 332.400 41.800 333.200 ;
        RECT 41.000 331.600 42.000 332.400 ;
        RECT 98.800 229.600 99.800 230.400 ;
        RECT 410.800 229.600 411.800 230.400 ;
        RECT 99.000 228.800 99.800 229.600 ;
        RECT 411.000 228.800 411.800 229.600 ;
        RECT 414.200 212.400 415.000 213.200 ;
        RECT 414.000 211.600 415.000 212.400 ;
      LAYER via1 ;
        RECT 273.200 371.600 274.000 372.400 ;
        RECT 41.200 331.600 42.000 332.400 ;
      LAYER metal2 ;
        RECT 273.200 371.600 274.000 372.400 ;
        RECT 414.000 371.600 414.800 372.400 ;
        RECT 273.300 368.400 273.900 371.600 ;
        RECT 414.100 368.400 414.700 371.600 ;
        RECT 273.200 367.600 274.000 368.400 ;
        RECT 414.000 367.600 414.800 368.400 ;
        RECT 273.300 356.400 273.900 367.600 ;
        RECT 41.200 355.600 42.000 356.400 ;
        RECT 273.200 355.600 274.000 356.400 ;
        RECT 41.300 332.400 41.900 355.600 ;
        RECT 414.100 354.400 414.700 367.600 ;
        RECT 414.000 353.600 414.800 354.400 ;
        RECT 41.200 331.600 42.000 332.400 ;
        RECT 98.800 231.600 99.600 232.400 ;
        RECT 98.900 230.400 99.500 231.600 ;
        RECT 98.800 229.600 99.600 230.400 ;
        RECT 410.800 229.600 411.600 230.400 ;
        RECT 414.000 229.600 414.800 230.400 ;
        RECT 414.100 212.400 414.700 229.600 ;
        RECT 414.000 211.600 414.800 212.400 ;
      LAYER metal3 ;
        RECT 273.200 368.300 274.000 368.400 ;
        RECT 414.000 368.300 414.800 368.400 ;
        RECT 273.200 367.700 414.800 368.300 ;
        RECT 273.200 367.600 274.000 367.700 ;
        RECT 414.000 367.600 414.800 367.700 ;
        RECT 41.200 356.300 42.000 356.400 ;
        RECT 94.000 356.300 94.800 356.400 ;
        RECT 273.200 356.300 274.000 356.400 ;
        RECT 41.200 355.700 274.000 356.300 ;
        RECT 41.200 355.600 42.000 355.700 ;
        RECT 94.000 355.600 94.800 355.700 ;
        RECT 273.200 355.600 274.000 355.700 ;
        RECT 414.000 353.600 414.800 354.400 ;
        RECT 41.200 332.300 42.000 332.400 ;
        RECT -1.900 331.700 42.000 332.300 ;
        RECT 41.200 331.600 42.000 331.700 ;
        RECT 94.000 232.300 94.800 232.400 ;
        RECT 98.800 232.300 99.600 232.400 ;
        RECT 94.000 231.700 99.600 232.300 ;
        RECT 94.000 231.600 94.800 231.700 ;
        RECT 98.800 231.600 99.600 231.700 ;
        RECT 410.800 230.300 411.600 230.400 ;
        RECT 414.000 230.300 414.800 230.400 ;
        RECT 410.800 229.700 414.800 230.300 ;
        RECT 410.800 229.600 411.600 229.700 ;
        RECT 414.000 229.600 414.800 229.700 ;
      LAYER metal4 ;
        RECT 93.800 231.400 95.000 356.600 ;
        RECT 413.800 229.400 415.000 354.600 ;
    END
  END clk
  PIN rst
    PORT
      LAYER metal1 ;
        RECT 226.800 346.800 227.600 348.400 ;
        RECT 545.200 348.300 546.000 348.400 ;
        RECT 546.800 348.300 547.600 348.400 ;
        RECT 545.200 347.700 547.600 348.300 ;
        RECT 545.200 347.600 546.000 347.700 ;
        RECT 546.800 346.800 547.600 347.700 ;
        RECT 230.000 333.600 230.800 335.200 ;
        RECT 610.800 333.600 611.600 335.200 ;
        RECT 545.200 306.800 546.000 308.400 ;
        RECT 230.000 266.800 230.800 268.400 ;
        RECT 230.000 226.800 230.800 228.400 ;
        RECT 390.000 213.600 390.800 215.200 ;
        RECT 230.000 186.800 230.800 188.400 ;
        RECT 511.600 186.800 512.400 188.400 ;
      LAYER via1 ;
        RECT 226.800 347.600 227.600 348.400 ;
        RECT 545.200 307.600 546.000 308.400 ;
        RECT 230.000 267.600 230.800 268.400 ;
        RECT 230.000 227.600 230.800 228.400 ;
        RECT 230.000 187.600 230.800 188.400 ;
        RECT 511.600 187.600 512.400 188.400 ;
      LAYER metal2 ;
        RECT 226.800 347.600 227.600 348.400 ;
        RECT 230.000 347.600 230.800 348.400 ;
        RECT 545.200 347.600 546.000 348.400 ;
        RECT 230.100 334.400 230.700 347.600 ;
        RECT 545.300 340.400 545.900 347.600 ;
        RECT 545.200 339.600 546.000 340.400 ;
        RECT 610.800 339.600 611.600 340.400 ;
        RECT 230.000 333.600 230.800 334.400 ;
        RECT 230.100 328.400 230.700 333.600 ;
        RECT 230.000 327.600 230.800 328.400 ;
        RECT 545.300 308.400 545.900 339.600 ;
        RECT 610.900 334.400 611.500 339.600 ;
        RECT 610.800 333.600 611.600 334.400 ;
        RECT 545.200 307.600 546.000 308.400 ;
        RECT 545.300 284.400 545.900 307.600 ;
        RECT 545.200 283.600 546.000 284.400 ;
        RECT 230.000 277.600 230.800 278.400 ;
        RECT 230.100 268.400 230.700 277.600 ;
        RECT 230.000 267.600 230.800 268.400 ;
        RECT 230.100 228.400 230.700 267.600 ;
        RECT 230.000 227.600 230.800 228.400 ;
        RECT 390.000 213.600 390.800 214.400 ;
        RECT 390.100 212.400 390.700 213.600 ;
        RECT 390.000 211.600 390.800 212.400 ;
        RECT 390.100 204.400 390.700 211.600 ;
        RECT 511.600 209.600 512.400 210.400 ;
        RECT 511.700 204.400 512.300 209.600 ;
        RECT 230.000 203.600 230.800 204.400 ;
        RECT 390.000 203.600 390.800 204.400 ;
        RECT 511.600 203.600 512.400 204.400 ;
        RECT 230.100 188.400 230.700 203.600 ;
        RECT 511.700 188.400 512.300 203.600 ;
        RECT 230.000 187.600 230.800 188.400 ;
        RECT 511.600 187.600 512.400 188.400 ;
      LAYER metal3 ;
        RECT 226.800 348.300 227.600 348.400 ;
        RECT 230.000 348.300 230.800 348.400 ;
        RECT 226.800 347.700 230.800 348.300 ;
        RECT 226.800 347.600 227.600 347.700 ;
        RECT 230.000 347.600 230.800 347.700 ;
        RECT 545.200 340.300 546.000 340.400 ;
        RECT 610.800 340.300 611.600 340.400 ;
        RECT 545.200 339.700 611.600 340.300 ;
        RECT 545.200 339.600 546.000 339.700 ;
        RECT 610.800 339.600 611.600 339.700 ;
        RECT 610.800 334.300 611.600 334.400 ;
        RECT 610.800 333.700 616.300 334.300 ;
        RECT 610.800 333.600 611.600 333.700 ;
        RECT 230.000 328.300 230.800 328.400 ;
        RECT 231.600 328.300 232.400 328.400 ;
        RECT 230.000 327.700 232.400 328.300 ;
        RECT 230.000 327.600 230.800 327.700 ;
        RECT 231.600 327.600 232.400 327.700 ;
        RECT 513.200 284.300 514.000 284.400 ;
        RECT 545.200 284.300 546.000 284.400 ;
        RECT 513.200 283.700 546.000 284.300 ;
        RECT 513.200 283.600 514.000 283.700 ;
        RECT 545.200 283.600 546.000 283.700 ;
        RECT 230.000 278.300 230.800 278.400 ;
        RECT 231.600 278.300 232.400 278.400 ;
        RECT 230.000 277.700 232.400 278.300 ;
        RECT 230.000 277.600 230.800 277.700 ;
        RECT 231.600 277.600 232.400 277.700 ;
        RECT 230.000 228.300 230.800 228.400 ;
        RECT 231.600 228.300 232.400 228.400 ;
        RECT 230.000 227.700 232.400 228.300 ;
        RECT 230.000 227.600 230.800 227.700 ;
        RECT 231.600 227.600 232.400 227.700 ;
        RECT 231.600 212.300 232.400 212.400 ;
        RECT 390.000 212.300 390.800 212.400 ;
        RECT 231.600 211.700 390.800 212.300 ;
        RECT 231.600 211.600 232.400 211.700 ;
        RECT 390.000 211.600 390.800 211.700 ;
        RECT 511.600 210.300 512.400 210.400 ;
        RECT 513.200 210.300 514.000 210.400 ;
        RECT 511.600 209.700 514.000 210.300 ;
        RECT 511.600 209.600 512.400 209.700 ;
        RECT 513.200 209.600 514.000 209.700 ;
        RECT 230.000 204.300 230.800 204.400 ;
        RECT 231.600 204.300 232.400 204.400 ;
        RECT 230.000 203.700 232.400 204.300 ;
        RECT 230.000 203.600 230.800 203.700 ;
        RECT 231.600 203.600 232.400 203.700 ;
        RECT 390.000 204.300 390.800 204.400 ;
        RECT 511.600 204.300 512.400 204.400 ;
        RECT 390.000 203.700 512.400 204.300 ;
        RECT 390.000 203.600 390.800 203.700 ;
        RECT 511.600 203.600 512.400 203.700 ;
      LAYER metal4 ;
        RECT 231.400 277.400 232.600 328.600 ;
        RECT 231.400 203.400 232.600 228.600 ;
        RECT 513.000 209.400 514.200 284.600 ;
    END
  END rst
  PIN dest[0]
    PORT
      LAYER metal1 ;
        RECT 1.200 64.800 2.000 66.400 ;
      LAYER via1 ;
        RECT 1.200 65.600 2.000 66.400 ;
      LAYER metal2 ;
        RECT 1.200 69.600 2.000 70.400 ;
        RECT 1.300 66.400 1.900 69.600 ;
        RECT 1.200 65.600 2.000 66.400 ;
      LAYER metal3 ;
        RECT 1.200 70.300 2.000 70.400 ;
        RECT -1.900 69.700 2.000 70.300 ;
        RECT 1.200 69.600 2.000 69.700 ;
    END
  END dest[0]
  PIN dest[1]
    PORT
      LAYER metal1 ;
        RECT 1.200 224.800 2.000 226.400 ;
      LAYER via1 ;
        RECT 1.200 225.600 2.000 226.400 ;
      LAYER metal2 ;
        RECT 1.200 233.600 2.000 234.400 ;
        RECT 1.300 226.400 1.900 233.600 ;
        RECT 1.200 225.600 2.000 226.400 ;
      LAYER metal3 ;
        RECT 1.200 234.300 2.000 234.400 ;
        RECT -1.900 233.700 2.000 234.300 ;
        RECT 1.200 233.600 2.000 233.700 ;
    END
  END dest[1]
  PIN dest[2]
    PORT
      LAYER metal1 ;
        RECT 604.400 144.800 605.200 146.400 ;
      LAYER via1 ;
        RECT 604.400 145.600 605.200 146.400 ;
      LAYER metal2 ;
        RECT 604.400 147.600 605.200 148.400 ;
        RECT 604.500 146.400 605.100 147.600 ;
        RECT 604.400 145.600 605.200 146.400 ;
      LAYER metal3 ;
        RECT 604.400 148.300 605.200 148.400 ;
        RECT 604.400 147.700 616.300 148.300 ;
        RECT 604.400 147.600 605.200 147.700 ;
    END
  END dest[2]
  PIN dest[3]
    PORT
      LAYER metal1 ;
        RECT 609.200 16.300 610.000 17.200 ;
        RECT 610.800 16.300 611.600 16.400 ;
        RECT 609.200 15.700 611.600 16.300 ;
        RECT 609.200 15.600 610.000 15.700 ;
        RECT 610.800 15.600 611.600 15.700 ;
      LAYER metal2 ;
        RECT 610.800 15.600 611.600 16.400 ;
        RECT 610.900 10.400 611.500 15.600 ;
        RECT 610.800 9.600 611.600 10.400 ;
      LAYER metal3 ;
        RECT 610.800 10.300 611.600 10.400 ;
        RECT 610.800 9.700 616.300 10.300 ;
        RECT 610.800 9.600 611.600 9.700 ;
    END
  END dest[3]
  PIN dest[4]
    PORT
      LAYER metal1 ;
        RECT 372.400 535.600 373.200 537.200 ;
      LAYER metal2 ;
        RECT 372.500 536.400 373.100 564.300 ;
        RECT 372.400 535.600 373.200 536.400 ;
    END
  END dest[4]
  PIN dest[5]
    PORT
      LAYER metal1 ;
        RECT 337.200 544.800 338.000 546.400 ;
      LAYER via1 ;
        RECT 337.200 545.600 338.000 546.400 ;
      LAYER metal2 ;
        RECT 337.300 546.400 337.900 564.300 ;
        RECT 337.200 545.600 338.000 546.400 ;
    END
  END dest[5]
  PIN dest[6]
    PORT
      LAYER metal1 ;
        RECT 1.200 344.800 2.000 346.400 ;
      LAYER via1 ;
        RECT 1.200 345.600 2.000 346.400 ;
      LAYER metal2 ;
        RECT 1.200 349.600 2.000 350.400 ;
        RECT 1.300 346.400 1.900 349.600 ;
        RECT 1.200 345.600 2.000 346.400 ;
      LAYER metal3 ;
        RECT 1.200 350.300 2.000 350.400 ;
        RECT -1.900 349.700 2.000 350.300 ;
        RECT 1.200 349.600 2.000 349.700 ;
    END
  END dest[6]
  PIN dest[7]
    PORT
      LAYER metal1 ;
        RECT 1.200 424.800 2.000 426.400 ;
      LAYER via1 ;
        RECT 1.200 425.600 2.000 426.400 ;
      LAYER metal2 ;
        RECT 1.200 429.600 2.000 430.400 ;
        RECT 1.300 426.400 1.900 429.600 ;
        RECT 1.200 425.600 2.000 426.400 ;
      LAYER metal3 ;
        RECT 1.200 430.300 2.000 430.400 ;
        RECT -1.900 429.700 2.000 430.300 ;
        RECT 1.200 429.600 2.000 429.700 ;
    END
  END dest[7]
  PIN ext_data_in[0]
    PORT
      LAYER metal1 ;
        RECT 50.800 15.600 51.600 17.200 ;
      LAYER metal2 ;
        RECT 50.800 15.600 51.600 16.400 ;
        RECT 50.900 -2.300 51.500 15.600 ;
    END
  END ext_data_in[0]
  PIN ext_data_in[1]
    PORT
      LAYER metal1 ;
        RECT 4.400 224.800 5.200 226.400 ;
      LAYER via1 ;
        RECT 4.400 225.600 5.200 226.400 ;
      LAYER metal2 ;
        RECT 4.400 229.600 5.200 230.400 ;
        RECT 4.500 226.400 5.100 229.600 ;
        RECT 4.400 225.600 5.200 226.400 ;
      LAYER metal3 ;
        RECT 4.400 230.300 5.200 230.400 ;
        RECT -1.900 229.700 5.200 230.300 ;
        RECT 4.400 229.600 5.200 229.700 ;
    END
  END ext_data_in[1]
  PIN ext_data_in[2]
    PORT
      LAYER metal1 ;
        RECT 49.200 24.800 50.000 26.400 ;
      LAYER via1 ;
        RECT 49.200 25.600 50.000 26.400 ;
      LAYER metal2 ;
        RECT 49.200 25.600 50.000 26.400 ;
        RECT 49.300 -1.700 49.900 25.600 ;
        RECT 47.700 -2.300 49.900 -1.700 ;
    END
  END ext_data_in[2]
  PIN ext_data_in[3]
    PORT
      LAYER metal1 ;
        RECT 1.200 215.600 2.000 217.200 ;
      LAYER metal2 ;
        RECT 1.200 215.600 2.000 216.400 ;
        RECT 1.300 210.400 1.900 215.600 ;
        RECT 1.200 209.600 2.000 210.400 ;
      LAYER metal3 ;
        RECT 1.200 210.300 2.000 210.400 ;
        RECT -1.900 209.700 2.000 210.300 ;
        RECT 1.200 209.600 2.000 209.700 ;
    END
  END ext_data_in[3]
  PIN ext_data_in[4]
    PORT
      LAYER metal1 ;
        RECT 607.600 176.300 608.400 177.200 ;
        RECT 612.400 176.300 613.200 176.400 ;
        RECT 607.600 175.700 613.200 176.300 ;
        RECT 607.600 175.600 608.400 175.700 ;
        RECT 612.400 175.600 613.200 175.700 ;
      LAYER metal2 ;
        RECT 612.400 175.600 613.200 176.400 ;
        RECT 612.500 170.400 613.100 175.600 ;
        RECT 612.400 169.600 613.200 170.400 ;
      LAYER metal3 ;
        RECT 612.400 170.300 613.200 170.400 ;
        RECT 612.400 169.700 616.300 170.300 ;
        RECT 612.400 169.600 613.200 169.700 ;
    END
  END ext_data_in[4]
  PIN ext_data_in[5]
    PORT
      LAYER metal1 ;
        RECT 567.600 24.800 568.400 26.400 ;
      LAYER via1 ;
        RECT 567.600 25.600 568.400 26.400 ;
      LAYER metal2 ;
        RECT 567.600 25.600 568.400 26.400 ;
        RECT 567.700 14.400 568.300 25.600 ;
        RECT 567.600 13.600 568.400 14.400 ;
        RECT 566.000 1.600 566.800 2.400 ;
        RECT 566.100 -2.300 566.700 1.600 ;
      LAYER metal3 ;
        RECT 567.600 13.600 568.400 14.400 ;
        RECT 566.000 2.300 566.800 2.400 ;
        RECT 567.600 2.300 568.400 2.400 ;
        RECT 566.000 1.700 568.400 2.300 ;
        RECT 566.000 1.600 566.800 1.700 ;
        RECT 567.600 1.600 568.400 1.700 ;
      LAYER metal4 ;
        RECT 567.400 1.400 568.600 14.600 ;
    END
  END ext_data_in[5]
  PIN ext_data_in[6]
    PORT
      LAYER metal1 ;
        RECT 564.400 15.600 565.200 17.200 ;
      LAYER metal2 ;
        RECT 564.400 15.600 565.200 16.400 ;
        RECT 564.500 -1.700 565.100 15.600 ;
        RECT 562.900 -2.300 565.100 -1.700 ;
    END
  END ext_data_in[6]
  PIN ext_data_in[7]
    PORT
      LAYER metal1 ;
        RECT 606.000 24.800 606.800 26.400 ;
      LAYER via1 ;
        RECT 606.000 25.600 606.800 26.400 ;
      LAYER metal2 ;
        RECT 606.000 27.600 606.800 28.400 ;
        RECT 606.100 26.400 606.700 27.600 ;
        RECT 606.000 25.600 606.800 26.400 ;
      LAYER metal3 ;
        RECT 606.000 28.300 606.800 28.400 ;
        RECT 606.000 27.700 616.300 28.300 ;
        RECT 606.000 27.600 606.800 27.700 ;
    END
  END ext_data_in[7]
  PIN ext_data_in[8]
    PORT
      LAYER metal1 ;
        RECT 535.600 544.800 536.400 546.400 ;
      LAYER via1 ;
        RECT 535.600 545.600 536.400 546.400 ;
      LAYER metal2 ;
        RECT 535.700 546.400 536.300 564.300 ;
        RECT 535.600 545.600 536.400 546.400 ;
    END
  END ext_data_in[8]
  PIN ext_data_in[9]
    PORT
      LAYER metal1 ;
        RECT 353.200 544.800 354.000 546.400 ;
      LAYER via1 ;
        RECT 353.200 545.600 354.000 546.400 ;
      LAYER metal2 ;
        RECT 353.300 546.400 353.900 564.300 ;
        RECT 353.200 545.600 354.000 546.400 ;
    END
  END ext_data_in[9]
  PIN ext_data_in[10]
    PORT
      LAYER metal1 ;
        RECT 358.000 535.600 358.800 537.200 ;
      LAYER metal2 ;
        RECT 356.500 538.300 357.100 564.300 ;
        RECT 356.500 537.700 358.700 538.300 ;
        RECT 358.100 536.400 358.700 537.700 ;
        RECT 358.000 535.600 358.800 536.400 ;
    END
  END ext_data_in[10]
  PIN ext_data_in[11]
    PORT
      LAYER metal1 ;
        RECT 607.600 535.600 608.400 537.200 ;
      LAYER metal2 ;
        RECT 606.100 554.300 606.700 564.300 ;
        RECT 606.100 553.700 608.300 554.300 ;
        RECT 607.700 536.400 608.300 553.700 ;
        RECT 607.600 535.600 608.400 536.400 ;
    END
  END ext_data_in[11]
  PIN ext_data_in[12]
    PORT
      LAYER metal1 ;
        RECT 47.600 535.600 48.400 537.200 ;
      LAYER metal2 ;
        RECT 46.100 563.700 48.300 564.300 ;
        RECT 46.100 552.300 46.700 563.700 ;
        RECT 46.100 551.700 48.300 552.300 ;
        RECT 47.700 536.400 48.300 551.700 ;
        RECT 47.600 535.600 48.400 536.400 ;
    END
  END ext_data_in[12]
  PIN ext_data_in[13]
    PORT
      LAYER metal1 ;
        RECT 4.400 375.600 5.200 377.200 ;
      LAYER metal2 ;
        RECT 4.400 375.600 5.200 376.400 ;
        RECT 4.500 374.300 5.100 375.600 ;
        RECT 2.900 373.700 5.100 374.300 ;
        RECT 2.900 370.400 3.500 373.700 ;
        RECT 2.800 369.600 3.600 370.400 ;
      LAYER metal3 ;
        RECT 2.800 370.300 3.600 370.400 ;
        RECT -1.900 369.700 3.600 370.300 ;
        RECT 2.800 369.600 3.600 369.700 ;
    END
  END ext_data_in[13]
  PIN ext_data_in[14]
    PORT
      LAYER metal1 ;
        RECT 1.200 375.600 2.000 377.200 ;
      LAYER metal2 ;
        RECT 1.200 375.600 2.000 376.400 ;
        RECT 1.300 374.400 1.900 375.600 ;
        RECT 1.200 373.600 2.000 374.400 ;
      LAYER metal3 ;
        RECT 1.200 374.300 2.000 374.400 ;
        RECT -1.900 373.700 2.000 374.300 ;
        RECT 1.200 373.600 2.000 373.700 ;
    END
  END ext_data_in[14]
  PIN ext_data_in[15]
    PORT
      LAYER metal1 ;
        RECT 50.800 544.800 51.600 546.400 ;
      LAYER via1 ;
        RECT 50.800 545.600 51.600 546.400 ;
      LAYER metal2 ;
        RECT 50.900 546.400 51.500 564.300 ;
        RECT 50.800 545.600 51.600 546.400 ;
    END
  END ext_data_in[15]
  PIN ext_data_out[0]
    PORT
      LAYER metal1 ;
        RECT 218.800 12.400 219.600 19.800 ;
        RECT 219.000 10.200 219.600 12.400 ;
        RECT 218.800 2.200 219.600 10.200 ;
      LAYER via1 ;
        RECT 218.800 3.600 219.600 4.400 ;
      LAYER metal2 ;
        RECT 218.800 3.600 219.600 4.400 ;
        RECT 218.900 -1.700 219.500 3.600 ;
        RECT 217.300 -2.300 219.500 -1.700 ;
    END
  END ext_data_out[0]
  PIN ext_data_out[1]
    PORT
      LAYER metal1 ;
        RECT 135.600 12.400 136.400 19.800 ;
        RECT 135.600 10.200 136.200 12.400 ;
        RECT 135.600 2.200 136.400 10.200 ;
      LAYER via1 ;
        RECT 135.600 3.600 136.400 4.400 ;
      LAYER metal2 ;
        RECT 135.600 3.600 136.400 4.400 ;
        RECT 135.700 -1.700 136.300 3.600 ;
        RECT 135.700 -2.300 137.900 -1.700 ;
    END
  END ext_data_out[1]
  PIN ext_data_out[2]
    PORT
      LAYER metal1 ;
        RECT 263.600 12.400 264.400 19.800 ;
        RECT 263.800 10.200 264.400 12.400 ;
        RECT 263.600 2.200 264.400 10.200 ;
      LAYER via1 ;
        RECT 263.600 3.600 264.400 4.400 ;
      LAYER metal2 ;
        RECT 263.600 3.600 264.400 4.400 ;
        RECT 263.700 -1.700 264.300 3.600 ;
        RECT 262.100 -2.300 264.300 -1.700 ;
    END
  END ext_data_out[2]
  PIN ext_data_out[3]
    PORT
      LAYER metal1 ;
        RECT 258.800 12.400 259.600 19.800 ;
        RECT 259.000 10.200 259.600 12.400 ;
        RECT 258.800 2.200 259.600 10.200 ;
      LAYER via1 ;
        RECT 258.800 3.600 259.600 4.400 ;
      LAYER metal2 ;
        RECT 258.800 3.600 259.600 4.400 ;
        RECT 258.900 -1.700 259.500 3.600 ;
        RECT 257.300 -2.300 259.500 -1.700 ;
    END
  END ext_data_out[3]
  PIN ext_data_out[4]
    PORT
      LAYER metal1 ;
        RECT 402.800 12.400 403.600 19.800 ;
        RECT 403.000 10.200 403.600 12.400 ;
        RECT 402.800 2.200 403.600 10.200 ;
      LAYER via1 ;
        RECT 402.800 3.600 403.600 4.400 ;
      LAYER metal2 ;
        RECT 402.800 3.600 403.600 4.400 ;
        RECT 402.900 -1.700 403.500 3.600 ;
        RECT 401.300 -2.300 403.500 -1.700 ;
    END
  END ext_data_out[4]
  PIN ext_data_out[5]
    PORT
      LAYER metal1 ;
        RECT 268.400 12.400 269.200 19.800 ;
        RECT 268.600 10.200 269.200 12.400 ;
        RECT 268.400 2.200 269.200 10.200 ;
      LAYER via1 ;
        RECT 268.400 3.600 269.200 4.400 ;
      LAYER metal2 ;
        RECT 268.400 3.600 269.200 4.400 ;
        RECT 268.500 -1.700 269.100 3.600 ;
        RECT 266.900 -2.300 269.100 -1.700 ;
    END
  END ext_data_out[5]
  PIN ext_data_out[6]
    PORT
      LAYER metal1 ;
        RECT 607.600 191.800 608.400 199.800 ;
        RECT 607.800 189.600 608.400 191.800 ;
        RECT 607.600 188.300 608.400 189.600 ;
        RECT 612.400 188.300 613.200 188.400 ;
        RECT 607.600 187.700 613.200 188.300 ;
        RECT 607.600 182.200 608.400 187.700 ;
        RECT 612.400 187.600 613.200 187.700 ;
      LAYER metal2 ;
        RECT 612.400 189.600 613.200 190.400 ;
        RECT 612.500 188.400 613.100 189.600 ;
        RECT 612.400 187.600 613.200 188.400 ;
      LAYER metal3 ;
        RECT 612.400 190.300 613.200 190.400 ;
        RECT 612.400 189.700 616.300 190.300 ;
        RECT 612.400 189.600 613.200 189.700 ;
    END
  END ext_data_out[6]
  PIN ext_data_out[7]
    PORT
      LAYER metal1 ;
        RECT 313.200 12.400 314.000 19.800 ;
        RECT 313.400 10.200 314.000 12.400 ;
        RECT 313.200 2.200 314.000 10.200 ;
      LAYER via1 ;
        RECT 313.200 3.600 314.000 4.400 ;
      LAYER metal2 ;
        RECT 313.200 3.600 314.000 4.400 ;
        RECT 313.300 -1.700 313.900 3.600 ;
        RECT 311.700 -2.300 313.900 -1.700 ;
    END
  END ext_data_out[7]
  PIN ext_data_out[8]
    PORT
      LAYER metal1 ;
        RECT 609.200 154.300 610.000 159.800 ;
        RECT 612.400 154.300 613.200 154.400 ;
        RECT 609.200 153.700 613.200 154.300 ;
        RECT 609.200 151.800 610.000 153.700 ;
        RECT 612.400 153.600 613.200 153.700 ;
        RECT 609.400 149.600 610.000 151.800 ;
        RECT 609.200 142.200 610.000 149.600 ;
      LAYER metal2 ;
        RECT 612.400 153.600 613.200 154.400 ;
        RECT 612.500 152.400 613.100 153.600 ;
        RECT 612.400 151.600 613.200 152.400 ;
      LAYER metal3 ;
        RECT 612.400 152.300 613.200 152.400 ;
        RECT 612.400 151.700 616.300 152.300 ;
        RECT 612.400 151.600 613.200 151.700 ;
    END
  END ext_data_out[8]
  PIN ext_data_out[9]
    PORT
      LAYER metal1 ;
        RECT 609.200 351.800 610.000 359.800 ;
        RECT 609.400 349.600 610.000 351.800 ;
        RECT 609.200 348.300 610.000 349.600 ;
        RECT 612.400 348.300 613.200 348.400 ;
        RECT 609.200 347.700 613.200 348.300 ;
        RECT 609.200 342.200 610.000 347.700 ;
        RECT 612.400 347.600 613.200 347.700 ;
      LAYER metal2 ;
        RECT 612.400 349.600 613.200 350.400 ;
        RECT 612.500 348.400 613.100 349.600 ;
        RECT 612.400 347.600 613.200 348.400 ;
      LAYER metal3 ;
        RECT 612.400 350.300 613.200 350.400 ;
        RECT 612.400 349.700 616.300 350.300 ;
        RECT 612.400 349.600 613.200 349.700 ;
    END
  END ext_data_out[9]
  PIN ext_data_out[10]
    PORT
      LAYER metal1 ;
        RECT 610.800 372.400 611.600 379.800 ;
        RECT 611.000 370.200 611.600 372.400 ;
        RECT 610.800 368.300 611.600 370.200 ;
        RECT 612.400 368.300 613.200 368.400 ;
        RECT 610.800 367.700 613.200 368.300 ;
        RECT 610.800 362.200 611.600 367.700 ;
        RECT 612.400 367.600 613.200 367.700 ;
      LAYER metal2 ;
        RECT 612.400 369.600 613.200 370.400 ;
        RECT 612.500 368.400 613.100 369.600 ;
        RECT 612.400 367.600 613.200 368.400 ;
      LAYER metal3 ;
        RECT 612.400 370.300 613.200 370.400 ;
        RECT 612.400 369.700 616.300 370.300 ;
        RECT 612.400 369.600 613.200 369.700 ;
    END
  END ext_data_out[10]
  PIN ext_data_out[11]
    PORT
      LAYER metal1 ;
        RECT 607.600 311.800 608.400 319.800 ;
        RECT 607.800 309.600 608.400 311.800 ;
        RECT 607.600 308.300 608.400 309.600 ;
        RECT 612.400 308.300 613.200 308.400 ;
        RECT 607.600 307.700 613.200 308.300 ;
        RECT 607.600 302.200 608.400 307.700 ;
        RECT 612.400 307.600 613.200 307.700 ;
      LAYER metal2 ;
        RECT 612.400 309.600 613.200 310.400 ;
        RECT 612.500 308.400 613.100 309.600 ;
        RECT 612.400 307.600 613.200 308.400 ;
      LAYER metal3 ;
        RECT 612.400 310.300 613.200 310.400 ;
        RECT 612.400 309.700 616.300 310.300 ;
        RECT 612.400 309.600 613.200 309.700 ;
    END
  END ext_data_out[11]
  PIN ext_data_out[12]
    PORT
      LAYER metal1 ;
        RECT 198.000 551.800 198.800 559.800 ;
        RECT 198.000 549.600 198.600 551.800 ;
        RECT 198.000 542.200 198.800 549.600 ;
      LAYER via1 ;
        RECT 198.000 557.600 198.800 558.400 ;
      LAYER metal2 ;
        RECT 198.100 563.700 200.300 564.300 ;
        RECT 198.100 558.400 198.700 563.700 ;
        RECT 198.000 557.600 198.800 558.400 ;
    END
  END ext_data_out[12]
  PIN ext_data_out[13]
    PORT
      LAYER metal1 ;
        RECT 252.400 551.800 253.200 559.800 ;
        RECT 252.400 549.600 253.000 551.800 ;
        RECT 252.400 542.200 253.200 549.600 ;
      LAYER via1 ;
        RECT 252.400 557.600 253.200 558.400 ;
      LAYER metal2 ;
        RECT 252.500 563.700 254.700 564.300 ;
        RECT 252.500 558.400 253.100 563.700 ;
        RECT 252.400 557.600 253.200 558.400 ;
    END
  END ext_data_out[13]
  PIN ext_data_out[14]
    PORT
      LAYER metal1 ;
        RECT 295.600 551.800 296.400 559.800 ;
        RECT 295.800 549.600 296.400 551.800 ;
        RECT 295.600 542.200 296.400 549.600 ;
      LAYER via1 ;
        RECT 295.600 557.600 296.400 558.400 ;
      LAYER metal2 ;
        RECT 294.100 563.700 296.300 564.300 ;
        RECT 295.700 558.400 296.300 563.700 ;
        RECT 295.600 557.600 296.400 558.400 ;
    END
  END ext_data_out[14]
  PIN ext_data_out[15]
    PORT
      LAYER metal1 ;
        RECT 178.800 551.800 179.600 559.800 ;
        RECT 178.800 549.600 179.400 551.800 ;
        RECT 178.800 542.200 179.600 549.600 ;
      LAYER via1 ;
        RECT 178.800 557.600 179.600 558.400 ;
      LAYER metal2 ;
        RECT 178.900 563.700 181.100 564.300 ;
        RECT 178.900 558.400 179.500 563.700 ;
        RECT 178.800 557.600 179.600 558.400 ;
    END
  END ext_data_out[15]
  PIN pe_busy[0]
    PORT
      LAYER metal1 ;
        RECT 1.200 31.800 2.000 39.800 ;
        RECT 1.200 29.600 1.800 31.800 ;
        RECT 1.200 22.200 2.000 29.600 ;
      LAYER via1 ;
        RECT 1.200 27.600 2.000 28.400 ;
      LAYER metal2 ;
        RECT 1.200 29.600 2.000 30.400 ;
        RECT 1.300 28.400 1.900 29.600 ;
        RECT 1.200 27.600 2.000 28.400 ;
      LAYER metal3 ;
        RECT 1.200 30.300 2.000 30.400 ;
        RECT -1.900 29.700 2.000 30.300 ;
        RECT 1.200 29.600 2.000 29.700 ;
    END
  END pe_busy[0]
  PIN pe_busy[1]
    PORT
      LAYER metal1 ;
        RECT 610.800 34.300 611.600 39.800 ;
        RECT 612.400 34.300 613.200 34.400 ;
        RECT 610.800 33.700 613.200 34.300 ;
        RECT 610.800 31.800 611.600 33.700 ;
        RECT 612.400 33.600 613.200 33.700 ;
        RECT 611.000 29.600 611.600 31.800 ;
        RECT 610.800 22.200 611.600 29.600 ;
      LAYER metal2 ;
        RECT 612.400 33.600 613.200 34.400 ;
        RECT 612.500 32.400 613.100 33.600 ;
        RECT 612.400 31.600 613.200 32.400 ;
      LAYER metal3 ;
        RECT 612.400 32.300 613.200 32.400 ;
        RECT 612.400 31.700 616.300 32.300 ;
        RECT 612.400 31.600 613.200 31.700 ;
    END
  END pe_busy[1]
  PIN pe_busy[2]
    PORT
      LAYER metal1 ;
        RECT 607.600 252.400 608.400 259.800 ;
        RECT 607.800 250.200 608.400 252.400 ;
        RECT 607.600 242.200 608.400 250.200 ;
      LAYER via1 ;
        RECT 607.600 257.600 608.400 258.400 ;
      LAYER metal2 ;
        RECT 609.300 560.400 609.900 564.300 ;
        RECT 609.200 559.600 610.000 560.400 ;
        RECT 607.600 333.600 608.400 334.400 ;
        RECT 607.700 258.400 608.300 333.600 ;
        RECT 607.600 257.600 608.400 258.400 ;
      LAYER metal3 ;
        RECT 609.200 559.600 610.000 560.400 ;
        RECT 607.600 334.300 608.400 334.400 ;
        RECT 609.200 334.300 610.000 334.400 ;
        RECT 607.600 333.700 610.000 334.300 ;
        RECT 607.600 333.600 608.400 333.700 ;
        RECT 609.200 333.600 610.000 333.700 ;
      LAYER metal4 ;
        RECT 609.000 333.400 610.200 560.600 ;
    END
  END pe_busy[2]
  PIN pe_busy[3]
    PORT
      LAYER metal1 ;
        RECT 39.600 551.800 40.400 559.800 ;
        RECT 39.600 549.600 40.200 551.800 ;
        RECT 39.600 542.200 40.400 549.600 ;
      LAYER via1 ;
        RECT 39.600 557.600 40.400 558.400 ;
      LAYER metal2 ;
        RECT 39.700 563.700 41.900 564.300 ;
        RECT 39.700 558.400 40.300 563.700 ;
        RECT 39.600 557.600 40.400 558.400 ;
    END
  END pe_busy[3]
  OBS
      LAYER metal1 ;
        RECT 1.200 548.300 2.000 559.800 ;
        RECT 6.000 556.400 6.800 559.800 ;
        RECT 5.800 555.800 6.800 556.400 ;
        RECT 5.800 555.200 6.400 555.800 ;
        RECT 9.200 555.200 10.000 559.800 ;
        RECT 12.400 557.000 13.200 559.800 ;
        RECT 14.000 557.000 14.800 559.800 ;
        RECT 4.400 554.600 6.400 555.200 ;
        RECT 4.400 549.000 5.200 554.600 ;
        RECT 7.000 554.400 11.200 555.200 ;
        RECT 15.600 555.000 16.400 559.800 ;
        RECT 18.800 555.000 19.600 559.800 ;
        RECT 7.000 554.000 7.600 554.400 ;
        RECT 6.000 553.200 7.600 554.000 ;
        RECT 10.600 553.800 16.400 554.400 ;
        RECT 8.600 553.200 10.000 553.800 ;
        RECT 8.600 553.000 14.800 553.200 ;
        RECT 9.400 552.600 14.800 553.000 ;
        RECT 14.000 552.400 14.800 552.600 ;
        RECT 15.800 553.000 16.400 553.800 ;
        RECT 17.000 553.600 19.600 554.400 ;
        RECT 22.000 553.600 22.800 559.800 ;
        RECT 23.600 557.000 24.400 559.800 ;
        RECT 25.200 557.000 26.000 559.800 ;
        RECT 26.800 557.000 27.600 559.800 ;
        RECT 25.200 554.400 29.400 555.200 ;
        RECT 30.000 554.400 30.800 559.800 ;
        RECT 33.200 555.200 34.000 559.800 ;
        RECT 33.200 554.600 35.800 555.200 ;
        RECT 30.000 553.600 32.600 554.400 ;
        RECT 23.600 553.000 24.400 553.200 ;
        RECT 15.800 552.400 24.400 553.000 ;
        RECT 26.800 553.000 27.600 553.200 ;
        RECT 35.200 553.000 35.800 554.600 ;
        RECT 26.800 552.400 35.800 553.000 ;
        RECT 35.200 550.600 35.800 552.400 ;
        RECT 36.400 552.000 37.200 559.800 ;
        RECT 42.800 552.400 43.600 559.800 ;
        RECT 36.400 551.200 37.400 552.000 ;
        RECT 41.400 551.800 43.600 552.400 ;
        RECT 41.400 551.200 42.000 551.800 ;
        RECT 5.800 550.000 29.200 550.600 ;
        RECT 35.200 550.000 36.000 550.600 ;
        RECT 5.800 549.800 6.800 550.000 ;
        RECT 6.000 549.600 6.800 549.800 ;
        RECT 10.800 549.600 11.600 550.000 ;
        RECT 28.400 549.400 29.200 550.000 ;
        RECT 2.800 548.300 3.600 548.400 ;
        RECT 1.200 547.700 3.600 548.300 ;
        RECT 1.200 542.200 2.000 547.700 ;
        RECT 2.800 547.600 3.600 547.700 ;
        RECT 4.400 548.200 13.200 549.000 ;
        RECT 13.800 548.600 15.800 549.400 ;
        RECT 19.600 548.600 22.800 549.400 ;
        RECT 2.800 544.800 3.600 546.400 ;
        RECT 4.400 542.200 5.200 548.200 ;
        RECT 6.800 546.800 9.800 547.600 ;
        RECT 9.000 546.200 9.800 546.800 ;
        RECT 15.000 546.200 15.800 548.600 ;
        RECT 17.200 546.800 18.000 548.400 ;
        RECT 22.400 547.800 23.200 548.000 ;
        RECT 18.800 547.200 23.200 547.800 ;
        RECT 18.800 547.000 19.600 547.200 ;
        RECT 25.200 546.400 26.000 549.200 ;
        RECT 31.000 548.600 34.800 549.400 ;
        RECT 31.000 547.400 31.800 548.600 ;
        RECT 35.400 548.000 36.000 550.000 ;
        RECT 18.800 546.200 19.600 546.400 ;
        RECT 9.000 545.400 11.600 546.200 ;
        RECT 15.000 545.600 19.600 546.200 ;
        RECT 20.400 545.600 22.000 546.400 ;
        RECT 25.000 545.600 26.000 546.400 ;
        RECT 30.000 546.800 31.800 547.400 ;
        RECT 34.800 547.400 36.000 548.000 ;
        RECT 30.000 546.200 30.800 546.800 ;
        RECT 10.800 542.200 11.600 545.400 ;
        RECT 28.400 545.400 30.800 546.200 ;
        RECT 12.400 542.200 13.200 545.000 ;
        RECT 14.000 542.200 14.800 545.000 ;
        RECT 15.600 542.200 16.400 545.000 ;
        RECT 18.800 542.200 19.600 545.000 ;
        RECT 22.000 542.200 22.800 545.000 ;
        RECT 23.600 542.200 24.400 545.000 ;
        RECT 25.200 542.200 26.000 545.000 ;
        RECT 26.800 542.200 27.600 545.000 ;
        RECT 28.400 542.200 29.200 545.400 ;
        RECT 34.800 542.200 35.600 547.400 ;
        RECT 36.600 546.800 37.400 551.200 ;
        RECT 40.800 550.400 42.000 551.200 ;
        RECT 41.400 547.400 42.000 550.400 ;
        RECT 42.800 550.300 43.600 550.400 ;
        RECT 44.400 550.300 45.200 550.400 ;
        RECT 42.800 549.700 45.200 550.300 ;
        RECT 42.800 548.800 43.600 549.700 ;
        RECT 44.400 549.600 45.200 549.700 ;
        RECT 41.400 546.800 43.600 547.400 ;
        RECT 44.400 546.800 45.200 548.400 ;
        RECT 36.400 546.300 37.400 546.800 ;
        RECT 38.000 546.300 38.800 546.400 ;
        RECT 36.400 545.700 38.800 546.300 ;
        RECT 36.400 542.200 37.200 545.700 ;
        RECT 38.000 545.600 38.800 545.700 ;
        RECT 42.800 542.200 43.600 546.800 ;
        RECT 46.000 546.200 46.800 559.800 ;
        RECT 47.600 551.600 48.400 554.400 ;
        RECT 49.200 548.300 50.000 559.800 ;
        RECT 55.000 552.400 55.800 559.800 ;
        RECT 56.400 553.600 57.200 554.400 ;
        RECT 56.600 552.400 57.200 553.600 ;
        RECT 61.400 552.400 62.200 559.800 ;
        RECT 62.800 554.300 63.600 554.400 ;
        RECT 66.800 554.300 67.600 559.800 ;
        RECT 70.000 555.200 70.800 559.800 ;
        RECT 62.800 553.700 67.600 554.300 ;
        RECT 62.800 553.600 63.600 553.700 ;
        RECT 63.000 552.400 63.600 553.600 ;
        RECT 55.000 551.800 56.000 552.400 ;
        RECT 56.600 551.800 58.000 552.400 ;
        RECT 52.400 550.300 53.200 550.400 ;
        RECT 54.000 550.300 54.800 550.400 ;
        RECT 52.400 549.700 54.800 550.300 ;
        RECT 52.400 549.600 53.200 549.700 ;
        RECT 54.000 548.800 54.800 549.700 ;
        RECT 55.400 548.400 56.000 551.800 ;
        RECT 57.200 551.600 58.000 551.800 ;
        RECT 60.400 551.600 62.400 552.400 ;
        RECT 63.000 551.800 64.400 552.400 ;
        RECT 66.800 552.000 67.600 553.700 ;
        RECT 63.600 551.600 64.400 551.800 ;
        RECT 60.400 548.800 61.200 550.400 ;
        RECT 61.800 548.400 62.400 551.600 ;
        RECT 66.600 551.200 67.600 552.000 ;
        RECT 68.200 554.600 70.800 555.200 ;
        RECT 68.200 553.000 68.800 554.600 ;
        RECT 73.200 554.400 74.000 559.800 ;
        RECT 76.400 557.000 77.200 559.800 ;
        RECT 78.000 557.000 78.800 559.800 ;
        RECT 79.600 557.000 80.400 559.800 ;
        RECT 74.600 554.400 78.800 555.200 ;
        RECT 71.400 553.600 74.000 554.400 ;
        RECT 81.200 553.600 82.000 559.800 ;
        RECT 84.400 555.000 85.200 559.800 ;
        RECT 87.600 555.000 88.400 559.800 ;
        RECT 89.200 557.000 90.000 559.800 ;
        RECT 90.800 557.000 91.600 559.800 ;
        RECT 94.000 555.200 94.800 559.800 ;
        RECT 97.200 556.400 98.000 559.800 ;
        RECT 97.200 555.800 98.200 556.400 ;
        RECT 97.600 555.200 98.200 555.800 ;
        RECT 92.800 554.400 97.000 555.200 ;
        RECT 97.600 554.600 99.600 555.200 ;
        RECT 84.400 553.600 87.000 554.400 ;
        RECT 87.600 553.800 93.400 554.400 ;
        RECT 96.400 554.000 97.000 554.400 ;
        RECT 76.400 553.000 77.200 553.200 ;
        RECT 68.200 552.400 77.200 553.000 ;
        RECT 79.600 553.000 80.400 553.200 ;
        RECT 87.600 553.000 88.200 553.800 ;
        RECT 94.000 553.200 95.400 553.800 ;
        RECT 96.400 553.200 98.000 554.000 ;
        RECT 79.600 552.400 88.200 553.000 ;
        RECT 89.200 553.000 95.400 553.200 ;
        RECT 89.200 552.600 94.600 553.000 ;
        RECT 89.200 552.400 90.000 552.600 ;
        RECT 52.400 548.300 53.200 548.400 ;
        RECT 49.200 548.200 53.200 548.300 ;
        RECT 49.200 547.700 54.000 548.200 ;
        RECT 46.000 545.600 47.800 546.200 ;
        RECT 47.000 544.400 47.800 545.600 ;
        RECT 46.000 543.600 47.800 544.400 ;
        RECT 47.000 542.200 47.800 543.600 ;
        RECT 49.200 542.200 50.000 547.700 ;
        RECT 52.400 547.600 54.000 547.700 ;
        RECT 55.400 547.600 58.000 548.400 ;
        RECT 58.800 548.200 59.600 548.400 ;
        RECT 58.800 547.600 60.400 548.200 ;
        RECT 61.800 547.600 64.400 548.400 ;
        RECT 53.200 547.200 54.000 547.600 ;
        RECT 52.600 546.200 56.200 546.600 ;
        RECT 57.200 546.200 57.800 547.600 ;
        RECT 59.600 547.200 60.400 547.600 ;
        RECT 59.000 546.200 62.600 546.600 ;
        RECT 63.600 546.200 64.200 547.600 ;
        RECT 66.600 546.800 67.400 551.200 ;
        RECT 68.200 550.600 68.800 552.400 ;
        RECT 68.000 550.000 68.800 550.600 ;
        RECT 74.800 550.000 98.200 550.600 ;
        RECT 68.000 548.000 68.600 550.000 ;
        RECT 74.800 549.400 75.600 550.000 ;
        RECT 92.400 549.600 93.200 550.000 ;
        RECT 95.600 549.600 96.400 550.000 ;
        RECT 97.400 549.800 98.200 550.000 ;
        RECT 69.200 548.600 73.000 549.400 ;
        RECT 68.000 547.400 69.200 548.000 ;
        RECT 52.400 546.000 56.400 546.200 ;
        RECT 52.400 542.200 53.200 546.000 ;
        RECT 55.600 542.200 56.400 546.000 ;
        RECT 57.200 542.200 58.000 546.200 ;
        RECT 58.800 546.000 62.800 546.200 ;
        RECT 58.800 542.200 59.600 546.000 ;
        RECT 62.000 542.200 62.800 546.000 ;
        RECT 63.600 542.200 64.400 546.200 ;
        RECT 66.600 546.000 67.600 546.800 ;
        RECT 66.800 542.200 67.600 546.000 ;
        RECT 68.400 542.200 69.200 547.400 ;
        RECT 72.200 547.400 73.000 548.600 ;
        RECT 72.200 546.800 74.000 547.400 ;
        RECT 73.200 546.200 74.000 546.800 ;
        RECT 78.000 546.400 78.800 549.200 ;
        RECT 81.200 548.600 84.400 549.400 ;
        RECT 88.200 548.600 90.200 549.400 ;
        RECT 98.800 549.000 99.600 554.600 ;
        RECT 100.400 551.400 101.200 559.800 ;
        RECT 104.800 556.400 105.600 559.800 ;
        RECT 103.600 555.800 105.600 556.400 ;
        RECT 109.200 555.800 110.000 559.800 ;
        RECT 113.400 555.800 114.600 559.800 ;
        RECT 103.600 555.000 104.400 555.800 ;
        RECT 109.200 555.200 109.800 555.800 ;
        RECT 107.000 554.600 110.600 555.200 ;
        RECT 113.200 555.000 114.000 555.800 ;
        RECT 107.000 554.400 107.800 554.600 ;
        RECT 109.800 554.400 110.600 554.600 ;
        RECT 103.600 553.000 104.400 553.200 ;
        RECT 108.200 553.000 109.000 553.200 ;
        RECT 103.600 552.400 109.000 553.000 ;
        RECT 109.600 553.000 111.800 553.600 ;
        RECT 109.600 551.800 110.200 553.000 ;
        RECT 111.000 552.800 111.800 553.000 ;
        RECT 113.400 553.200 114.800 554.000 ;
        RECT 113.400 552.200 114.000 553.200 ;
        RECT 105.400 551.400 110.200 551.800 ;
        RECT 100.400 551.200 110.200 551.400 ;
        RECT 111.600 551.600 114.000 552.200 ;
        RECT 100.400 551.000 106.200 551.200 ;
        RECT 100.400 550.800 106.000 551.000 ;
        RECT 106.800 550.200 107.600 550.400 ;
        RECT 102.600 549.600 107.600 550.200 ;
        RECT 102.600 549.400 103.400 549.600 ;
        RECT 105.200 549.400 106.000 549.600 ;
        RECT 80.800 547.800 81.600 548.000 ;
        RECT 80.800 547.200 85.200 547.800 ;
        RECT 84.400 547.000 85.200 547.200 ;
        RECT 86.000 546.800 86.800 548.400 ;
        RECT 73.200 545.400 75.600 546.200 ;
        RECT 78.000 545.600 79.000 546.400 ;
        RECT 82.000 545.600 83.600 546.400 ;
        RECT 84.400 546.200 85.200 546.400 ;
        RECT 88.200 546.200 89.000 548.600 ;
        RECT 90.800 548.200 99.600 549.000 ;
        RECT 104.200 548.400 105.000 548.600 ;
        RECT 111.600 548.400 112.200 551.600 ;
        RECT 118.000 551.200 118.800 559.800 ;
        RECT 114.600 550.600 118.800 551.200 ;
        RECT 119.600 551.400 120.400 559.800 ;
        RECT 124.000 556.400 124.800 559.800 ;
        RECT 122.800 555.800 124.800 556.400 ;
        RECT 128.400 555.800 129.200 559.800 ;
        RECT 132.600 555.800 133.800 559.800 ;
        RECT 122.800 555.000 123.600 555.800 ;
        RECT 128.400 555.200 129.000 555.800 ;
        RECT 126.200 554.600 129.800 555.200 ;
        RECT 132.400 555.000 133.200 555.800 ;
        RECT 126.200 554.400 127.000 554.600 ;
        RECT 129.000 554.400 129.800 554.600 ;
        RECT 122.800 553.000 123.600 553.200 ;
        RECT 127.400 553.000 128.200 553.200 ;
        RECT 122.800 552.400 128.200 553.000 ;
        RECT 128.800 553.000 131.000 553.600 ;
        RECT 128.800 551.800 129.400 553.000 ;
        RECT 130.200 552.800 131.000 553.000 ;
        RECT 132.600 553.200 134.000 554.000 ;
        RECT 132.600 552.200 133.200 553.200 ;
        RECT 124.600 551.400 129.400 551.800 ;
        RECT 119.600 551.200 129.400 551.400 ;
        RECT 130.800 551.600 133.200 552.200 ;
        RECT 119.600 551.000 125.400 551.200 ;
        RECT 119.600 550.800 125.200 551.000 ;
        RECT 114.600 550.400 115.400 550.600 ;
        RECT 116.200 549.800 117.000 550.000 ;
        RECT 113.200 549.200 117.000 549.800 ;
        RECT 113.200 549.000 114.000 549.200 ;
        RECT 94.200 546.800 97.200 547.600 ;
        RECT 94.200 546.200 95.000 546.800 ;
        RECT 84.400 545.600 89.000 546.200 ;
        RECT 74.800 542.200 75.600 545.400 ;
        RECT 92.400 545.400 95.000 546.200 ;
        RECT 76.400 542.200 77.200 545.000 ;
        RECT 78.000 542.200 78.800 545.000 ;
        RECT 79.600 542.200 80.400 545.000 ;
        RECT 81.200 542.200 82.000 545.000 ;
        RECT 84.400 542.200 85.200 545.000 ;
        RECT 87.600 542.200 88.400 545.000 ;
        RECT 89.200 542.200 90.000 545.000 ;
        RECT 90.800 542.200 91.600 545.000 ;
        RECT 92.400 542.200 93.200 545.400 ;
        RECT 98.800 542.200 99.600 548.200 ;
        RECT 101.200 547.800 112.400 548.400 ;
        RECT 101.200 547.600 102.800 547.800 ;
        RECT 100.400 542.200 101.200 547.000 ;
        RECT 105.400 545.600 106.000 547.800 ;
        RECT 111.000 547.600 112.400 547.800 ;
        RECT 118.000 547.200 118.800 550.600 ;
        RECT 126.000 550.200 126.800 550.400 ;
        RECT 121.800 549.600 126.800 550.200 ;
        RECT 121.800 549.400 122.600 549.600 ;
        RECT 124.400 549.400 125.200 549.600 ;
        RECT 123.400 548.400 124.200 548.600 ;
        RECT 130.800 548.400 131.400 551.600 ;
        RECT 137.200 551.200 138.000 559.800 ;
        RECT 145.200 556.400 146.000 559.800 ;
        RECT 145.000 555.800 146.000 556.400 ;
        RECT 145.000 555.200 145.600 555.800 ;
        RECT 148.400 555.200 149.200 559.800 ;
        RECT 151.600 557.000 152.400 559.800 ;
        RECT 153.200 557.000 154.000 559.800 ;
        RECT 133.800 550.600 138.000 551.200 ;
        RECT 133.800 550.400 134.600 550.600 ;
        RECT 135.400 549.800 136.200 550.000 ;
        RECT 132.400 549.200 136.200 549.800 ;
        RECT 132.400 549.000 133.200 549.200 ;
        RECT 120.400 547.800 131.400 548.400 ;
        RECT 120.400 547.600 122.000 547.800 ;
        RECT 115.000 546.600 118.800 547.200 ;
        RECT 115.000 546.400 115.800 546.600 ;
        RECT 103.600 544.200 104.400 545.000 ;
        RECT 105.200 544.800 106.000 545.600 ;
        RECT 107.000 545.400 107.800 545.600 ;
        RECT 107.000 544.800 109.800 545.400 ;
        RECT 109.200 544.200 109.800 544.800 ;
        RECT 113.200 544.200 114.000 545.000 ;
        RECT 103.600 543.600 105.600 544.200 ;
        RECT 104.800 542.200 105.600 543.600 ;
        RECT 109.200 542.200 110.000 544.200 ;
        RECT 113.200 543.600 114.600 544.200 ;
        RECT 113.400 542.200 114.600 543.600 ;
        RECT 118.000 542.200 118.800 546.600 ;
        RECT 119.600 542.200 120.400 547.000 ;
        RECT 124.600 545.600 125.200 547.800 ;
        RECT 130.200 547.600 131.000 547.800 ;
        RECT 137.200 547.200 138.000 550.600 ;
        RECT 134.200 546.600 138.000 547.200 ;
        RECT 134.200 546.400 135.000 546.600 ;
        RECT 122.800 544.200 123.600 545.000 ;
        RECT 124.400 544.800 125.200 545.600 ;
        RECT 126.200 545.400 127.000 545.600 ;
        RECT 126.200 544.800 129.000 545.400 ;
        RECT 128.400 544.200 129.000 544.800 ;
        RECT 132.400 544.200 133.200 545.000 ;
        RECT 122.800 543.600 124.800 544.200 ;
        RECT 124.000 542.200 124.800 543.600 ;
        RECT 128.400 542.200 129.200 544.200 ;
        RECT 132.400 543.600 133.800 544.200 ;
        RECT 132.600 542.200 133.800 543.600 ;
        RECT 137.200 542.200 138.000 546.600 ;
        RECT 143.600 554.600 145.600 555.200 ;
        RECT 143.600 549.000 144.400 554.600 ;
        RECT 146.200 554.400 150.400 555.200 ;
        RECT 154.800 555.000 155.600 559.800 ;
        RECT 158.000 555.000 158.800 559.800 ;
        RECT 146.200 554.000 146.800 554.400 ;
        RECT 145.200 553.200 146.800 554.000 ;
        RECT 149.800 553.800 155.600 554.400 ;
        RECT 147.800 553.200 149.200 553.800 ;
        RECT 147.800 553.000 154.000 553.200 ;
        RECT 148.600 552.600 154.000 553.000 ;
        RECT 153.200 552.400 154.000 552.600 ;
        RECT 155.000 553.000 155.600 553.800 ;
        RECT 156.200 553.600 158.800 554.400 ;
        RECT 161.200 553.600 162.000 559.800 ;
        RECT 162.800 557.000 163.600 559.800 ;
        RECT 164.400 557.000 165.200 559.800 ;
        RECT 166.000 557.000 166.800 559.800 ;
        RECT 164.400 554.400 168.600 555.200 ;
        RECT 169.200 554.400 170.000 559.800 ;
        RECT 172.400 555.200 173.200 559.800 ;
        RECT 172.400 554.600 175.000 555.200 ;
        RECT 169.200 553.600 171.800 554.400 ;
        RECT 162.800 553.000 163.600 553.200 ;
        RECT 155.000 552.400 163.600 553.000 ;
        RECT 166.000 553.000 166.800 553.200 ;
        RECT 174.400 553.000 175.000 554.600 ;
        RECT 166.000 552.400 175.000 553.000 ;
        RECT 174.400 550.600 175.000 552.400 ;
        RECT 175.600 552.000 176.400 559.800 ;
        RECT 182.000 552.400 182.800 559.800 ;
        RECT 175.600 551.200 176.600 552.000 ;
        RECT 180.600 551.800 182.800 552.400 ;
        RECT 180.600 551.200 181.200 551.800 ;
        RECT 145.000 550.000 168.400 550.600 ;
        RECT 174.400 550.000 175.200 550.600 ;
        RECT 145.000 549.800 146.000 550.000 ;
        RECT 145.200 549.600 146.000 549.800 ;
        RECT 150.000 549.600 150.800 550.000 ;
        RECT 167.600 549.400 168.400 550.000 ;
        RECT 143.600 548.200 152.400 549.000 ;
        RECT 153.000 548.600 155.000 549.400 ;
        RECT 158.800 548.600 162.000 549.400 ;
        RECT 143.600 542.200 144.400 548.200 ;
        RECT 146.000 546.800 149.000 547.600 ;
        RECT 148.200 546.200 149.000 546.800 ;
        RECT 154.200 546.200 155.000 548.600 ;
        RECT 156.400 546.800 157.200 548.400 ;
        RECT 161.600 547.800 162.400 548.000 ;
        RECT 158.000 547.200 162.400 547.800 ;
        RECT 158.000 547.000 158.800 547.200 ;
        RECT 164.400 546.400 165.200 549.200 ;
        RECT 170.200 548.600 174.000 549.400 ;
        RECT 170.200 547.400 171.000 548.600 ;
        RECT 174.600 548.000 175.200 550.000 ;
        RECT 158.000 546.200 158.800 546.400 ;
        RECT 148.200 545.400 150.800 546.200 ;
        RECT 154.200 545.600 158.800 546.200 ;
        RECT 159.600 545.600 161.200 546.400 ;
        RECT 164.200 545.600 165.200 546.400 ;
        RECT 169.200 546.800 171.000 547.400 ;
        RECT 174.000 547.400 175.200 548.000 ;
        RECT 169.200 546.200 170.000 546.800 ;
        RECT 150.000 542.200 150.800 545.400 ;
        RECT 167.600 545.400 170.000 546.200 ;
        RECT 151.600 542.200 152.400 545.000 ;
        RECT 153.200 542.200 154.000 545.000 ;
        RECT 154.800 542.200 155.600 545.000 ;
        RECT 158.000 542.200 158.800 545.000 ;
        RECT 161.200 542.200 162.000 545.000 ;
        RECT 162.800 542.200 163.600 545.000 ;
        RECT 164.400 542.200 165.200 545.000 ;
        RECT 166.000 542.200 166.800 545.000 ;
        RECT 167.600 542.200 168.400 545.400 ;
        RECT 174.000 542.200 174.800 547.400 ;
        RECT 175.800 546.800 176.600 551.200 ;
        RECT 180.000 550.400 181.200 551.200 ;
        RECT 180.600 547.400 181.200 550.400 ;
        RECT 182.000 550.300 182.800 550.400 ;
        RECT 183.600 550.300 184.400 550.400 ;
        RECT 182.000 549.700 184.400 550.300 ;
        RECT 182.000 548.800 182.800 549.700 ;
        RECT 183.600 549.600 184.400 549.700 ;
        RECT 185.200 550.300 186.000 559.800 ;
        RECT 189.000 554.400 189.800 559.800 ;
        RECT 187.600 553.600 188.400 554.400 ;
        RECT 189.000 553.600 190.800 554.400 ;
        RECT 187.600 552.400 188.200 553.600 ;
        RECT 189.000 552.400 189.800 553.600 ;
        RECT 186.800 551.800 188.200 552.400 ;
        RECT 188.800 551.800 189.800 552.400 ;
        RECT 193.200 552.300 194.000 552.400 ;
        RECT 194.800 552.300 195.600 559.800 ;
        RECT 186.800 551.600 187.600 551.800 ;
        RECT 186.800 550.300 187.600 550.400 ;
        RECT 185.200 549.700 187.600 550.300 ;
        RECT 180.600 546.800 182.800 547.400 ;
        RECT 175.600 546.000 176.600 546.800 ;
        RECT 175.600 542.200 176.400 546.000 ;
        RECT 182.000 542.200 182.800 546.800 ;
        RECT 183.600 544.800 184.400 546.400 ;
        RECT 185.200 542.200 186.000 549.700 ;
        RECT 186.800 549.600 187.600 549.700 ;
        RECT 188.800 548.400 189.400 551.800 ;
        RECT 193.200 551.700 195.600 552.300 ;
        RECT 193.200 551.600 194.000 551.700 ;
        RECT 190.000 548.800 190.800 550.400 ;
        RECT 186.800 547.600 189.400 548.400 ;
        RECT 191.600 548.300 192.400 548.400 ;
        RECT 193.200 548.300 194.000 548.400 ;
        RECT 191.600 548.200 194.000 548.300 ;
        RECT 190.800 547.700 194.000 548.200 ;
        RECT 190.800 547.600 192.400 547.700 ;
        RECT 187.000 546.200 187.600 547.600 ;
        RECT 190.800 547.200 191.600 547.600 ;
        RECT 193.200 546.800 194.000 547.700 ;
        RECT 188.600 546.200 192.200 546.600 ;
        RECT 194.800 546.200 195.600 551.700 ;
        RECT 196.400 551.600 197.200 553.200 ;
        RECT 201.200 552.400 202.000 559.800 ;
        RECT 204.400 556.400 205.200 559.800 ;
        RECT 204.200 555.800 205.200 556.400 ;
        RECT 204.200 555.200 204.800 555.800 ;
        RECT 207.600 555.200 208.400 559.800 ;
        RECT 210.800 557.000 211.600 559.800 ;
        RECT 212.400 557.000 213.200 559.800 ;
        RECT 199.800 551.800 202.000 552.400 ;
        RECT 202.800 554.600 204.800 555.200 ;
        RECT 199.800 551.200 200.400 551.800 ;
        RECT 199.200 550.400 200.400 551.200 ;
        RECT 199.800 547.400 200.400 550.400 ;
        RECT 201.200 548.800 202.000 550.400 ;
        RECT 202.800 549.000 203.600 554.600 ;
        RECT 205.400 554.400 209.600 555.200 ;
        RECT 214.000 555.000 214.800 559.800 ;
        RECT 217.200 555.000 218.000 559.800 ;
        RECT 205.400 554.000 206.000 554.400 ;
        RECT 204.400 553.200 206.000 554.000 ;
        RECT 209.000 553.800 214.800 554.400 ;
        RECT 207.000 553.200 208.400 553.800 ;
        RECT 207.000 553.000 213.200 553.200 ;
        RECT 207.800 552.600 213.200 553.000 ;
        RECT 212.400 552.400 213.200 552.600 ;
        RECT 214.200 553.000 214.800 553.800 ;
        RECT 215.400 553.600 218.000 554.400 ;
        RECT 220.400 553.600 221.200 559.800 ;
        RECT 222.000 557.000 222.800 559.800 ;
        RECT 223.600 557.000 224.400 559.800 ;
        RECT 225.200 557.000 226.000 559.800 ;
        RECT 223.600 554.400 227.800 555.200 ;
        RECT 228.400 554.400 229.200 559.800 ;
        RECT 231.600 555.200 232.400 559.800 ;
        RECT 231.600 554.600 234.200 555.200 ;
        RECT 228.400 553.600 231.000 554.400 ;
        RECT 222.000 553.000 222.800 553.200 ;
        RECT 214.200 552.400 222.800 553.000 ;
        RECT 225.200 553.000 226.000 553.200 ;
        RECT 233.600 553.000 234.200 554.600 ;
        RECT 225.200 552.400 234.200 553.000 ;
        RECT 233.600 550.600 234.200 552.400 ;
        RECT 234.800 552.000 235.600 559.800 ;
        RECT 234.800 551.200 235.800 552.000 ;
        RECT 204.200 550.000 227.600 550.600 ;
        RECT 233.600 550.000 234.400 550.600 ;
        RECT 204.200 549.800 205.200 550.000 ;
        RECT 204.400 549.600 205.200 549.800 ;
        RECT 209.200 549.600 210.000 550.000 ;
        RECT 226.800 549.400 227.600 550.000 ;
        RECT 202.800 548.200 211.600 549.000 ;
        RECT 212.200 548.600 214.200 549.400 ;
        RECT 218.000 548.600 221.200 549.400 ;
        RECT 199.800 546.800 202.000 547.400 ;
        RECT 186.800 542.200 187.600 546.200 ;
        RECT 188.400 546.000 192.400 546.200 ;
        RECT 188.400 542.200 189.200 546.000 ;
        RECT 191.600 542.200 192.400 546.000 ;
        RECT 194.800 545.600 196.600 546.200 ;
        RECT 195.800 542.200 196.600 545.600 ;
        RECT 201.200 542.200 202.000 546.800 ;
        RECT 202.800 542.200 203.600 548.200 ;
        RECT 205.200 546.800 208.200 547.600 ;
        RECT 207.400 546.200 208.200 546.800 ;
        RECT 213.400 546.200 214.200 548.600 ;
        RECT 215.600 546.800 216.400 548.400 ;
        RECT 220.800 547.800 221.600 548.000 ;
        RECT 217.200 547.200 221.600 547.800 ;
        RECT 217.200 547.000 218.000 547.200 ;
        RECT 223.600 546.400 224.400 549.200 ;
        RECT 229.400 548.600 233.200 549.400 ;
        RECT 229.400 547.400 230.200 548.600 ;
        RECT 233.800 548.000 234.400 550.000 ;
        RECT 217.200 546.200 218.000 546.400 ;
        RECT 207.400 545.400 210.000 546.200 ;
        RECT 213.400 545.600 218.000 546.200 ;
        RECT 218.800 545.600 220.400 546.400 ;
        RECT 223.400 545.600 224.400 546.400 ;
        RECT 228.400 546.800 230.200 547.400 ;
        RECT 233.200 547.400 234.400 548.000 ;
        RECT 228.400 546.200 229.200 546.800 ;
        RECT 209.200 542.200 210.000 545.400 ;
        RECT 226.800 545.400 229.200 546.200 ;
        RECT 210.800 542.200 211.600 545.000 ;
        RECT 212.400 542.200 213.200 545.000 ;
        RECT 214.000 542.200 214.800 545.000 ;
        RECT 217.200 542.200 218.000 545.000 ;
        RECT 220.400 542.200 221.200 545.000 ;
        RECT 222.000 542.200 222.800 545.000 ;
        RECT 223.600 542.200 224.400 545.000 ;
        RECT 225.200 542.200 226.000 545.000 ;
        RECT 226.800 542.200 227.600 545.400 ;
        RECT 233.200 542.200 234.000 547.400 ;
        RECT 235.000 546.800 235.800 551.200 ;
        RECT 234.800 546.300 235.800 546.800 ;
        RECT 239.600 550.300 240.400 559.800 ;
        RECT 243.800 552.400 244.600 559.800 ;
        RECT 245.200 553.600 246.000 554.400 ;
        RECT 245.400 552.400 246.000 553.600 ;
        RECT 243.800 551.800 244.800 552.400 ;
        RECT 245.400 552.300 246.800 552.400 ;
        RECT 249.200 552.300 250.000 559.800 ;
        RECT 245.400 551.800 250.000 552.300 ;
        RECT 244.200 550.400 244.800 551.800 ;
        RECT 246.000 551.700 250.000 551.800 ;
        RECT 246.000 551.600 246.800 551.700 ;
        RECT 242.800 550.300 243.600 550.400 ;
        RECT 239.600 549.700 243.600 550.300 ;
        RECT 238.000 546.300 238.800 546.400 ;
        RECT 234.800 545.700 238.800 546.300 ;
        RECT 234.800 542.200 235.600 545.700 ;
        RECT 238.000 544.800 238.800 545.700 ;
        RECT 239.600 542.200 240.400 549.700 ;
        RECT 242.800 548.800 243.600 549.700 ;
        RECT 244.200 549.600 245.200 550.400 ;
        RECT 244.200 548.400 244.800 549.600 ;
        RECT 241.200 548.200 242.000 548.400 ;
        RECT 241.200 547.600 242.800 548.200 ;
        RECT 244.200 547.600 246.800 548.400 ;
        RECT 242.000 547.200 242.800 547.600 ;
        RECT 241.400 546.200 245.000 546.600 ;
        RECT 246.000 546.200 246.600 547.600 ;
        RECT 247.600 546.800 248.400 548.400 ;
        RECT 249.200 546.200 250.000 551.700 ;
        RECT 250.800 551.600 251.600 553.200 ;
        RECT 255.600 552.400 256.400 559.800 ;
        RECT 258.800 556.400 259.600 559.800 ;
        RECT 258.600 555.800 259.600 556.400 ;
        RECT 258.600 555.200 259.200 555.800 ;
        RECT 262.000 555.200 262.800 559.800 ;
        RECT 265.200 557.000 266.000 559.800 ;
        RECT 266.800 557.000 267.600 559.800 ;
        RECT 254.200 551.800 256.400 552.400 ;
        RECT 257.200 554.600 259.200 555.200 ;
        RECT 254.200 551.200 254.800 551.800 ;
        RECT 253.600 550.400 254.800 551.200 ;
        RECT 254.200 547.400 254.800 550.400 ;
        RECT 255.600 548.800 256.400 550.400 ;
        RECT 257.200 549.000 258.000 554.600 ;
        RECT 259.800 554.400 264.000 555.200 ;
        RECT 268.400 555.000 269.200 559.800 ;
        RECT 271.600 555.000 272.400 559.800 ;
        RECT 259.800 554.000 260.400 554.400 ;
        RECT 258.800 553.200 260.400 554.000 ;
        RECT 263.400 553.800 269.200 554.400 ;
        RECT 261.400 553.200 262.800 553.800 ;
        RECT 261.400 553.000 267.600 553.200 ;
        RECT 262.200 552.600 267.600 553.000 ;
        RECT 266.800 552.400 267.600 552.600 ;
        RECT 268.600 553.000 269.200 553.800 ;
        RECT 269.800 553.600 272.400 554.400 ;
        RECT 274.800 553.600 275.600 559.800 ;
        RECT 276.400 557.000 277.200 559.800 ;
        RECT 278.000 557.000 278.800 559.800 ;
        RECT 279.600 557.000 280.400 559.800 ;
        RECT 278.000 554.400 282.200 555.200 ;
        RECT 282.800 554.400 283.600 559.800 ;
        RECT 286.000 555.200 286.800 559.800 ;
        RECT 286.000 554.600 288.600 555.200 ;
        RECT 282.800 553.600 285.400 554.400 ;
        RECT 276.400 553.000 277.200 553.200 ;
        RECT 268.600 552.400 277.200 553.000 ;
        RECT 279.600 553.000 280.400 553.200 ;
        RECT 288.000 553.000 288.600 554.600 ;
        RECT 279.600 552.400 288.600 553.000 ;
        RECT 288.000 550.600 288.600 552.400 ;
        RECT 289.200 552.000 290.000 559.800 ;
        RECT 292.400 552.400 293.200 559.800 ;
        RECT 289.200 551.200 290.200 552.000 ;
        RECT 292.400 551.800 294.600 552.400 ;
        RECT 303.600 552.000 304.400 559.800 ;
        RECT 306.800 555.200 307.600 559.800 ;
        RECT 258.600 550.000 282.000 550.600 ;
        RECT 288.000 550.000 288.800 550.600 ;
        RECT 258.600 549.800 259.400 550.000 ;
        RECT 262.000 549.600 262.800 550.000 ;
        RECT 263.600 549.600 264.400 550.000 ;
        RECT 281.200 549.400 282.000 550.000 ;
        RECT 257.200 548.200 266.000 549.000 ;
        RECT 266.600 548.600 268.600 549.400 ;
        RECT 272.400 548.600 275.600 549.400 ;
        RECT 254.200 546.800 256.400 547.400 ;
        RECT 241.200 546.000 245.200 546.200 ;
        RECT 241.200 542.200 242.000 546.000 ;
        RECT 244.400 542.200 245.200 546.000 ;
        RECT 246.000 542.200 246.800 546.200 ;
        RECT 249.200 545.600 251.000 546.200 ;
        RECT 250.200 542.200 251.000 545.600 ;
        RECT 255.600 542.200 256.400 546.800 ;
        RECT 257.200 542.200 258.000 548.200 ;
        RECT 259.600 546.800 262.600 547.600 ;
        RECT 261.800 546.200 262.600 546.800 ;
        RECT 267.800 546.200 268.600 548.600 ;
        RECT 270.000 546.800 270.800 548.400 ;
        RECT 275.200 547.800 276.000 548.000 ;
        RECT 271.600 547.200 276.000 547.800 ;
        RECT 271.600 547.000 272.400 547.200 ;
        RECT 278.000 546.400 278.800 549.200 ;
        RECT 283.800 548.600 287.600 549.400 ;
        RECT 283.800 547.400 284.600 548.600 ;
        RECT 288.200 548.000 288.800 550.000 ;
        RECT 271.600 546.200 272.400 546.400 ;
        RECT 261.800 545.400 264.400 546.200 ;
        RECT 267.800 545.600 272.400 546.200 ;
        RECT 273.200 545.600 274.800 546.400 ;
        RECT 277.800 545.600 278.800 546.400 ;
        RECT 282.800 546.800 284.600 547.400 ;
        RECT 287.600 547.400 288.800 548.000 ;
        RECT 289.400 550.300 290.200 551.200 ;
        RECT 294.000 551.200 294.600 551.800 ;
        RECT 303.400 551.200 304.400 552.000 ;
        RECT 305.000 554.600 307.600 555.200 ;
        RECT 305.000 553.000 305.600 554.600 ;
        RECT 310.000 554.400 310.800 559.800 ;
        RECT 313.200 557.000 314.000 559.800 ;
        RECT 314.800 557.000 315.600 559.800 ;
        RECT 316.400 557.000 317.200 559.800 ;
        RECT 311.400 554.400 315.600 555.200 ;
        RECT 308.200 553.600 310.800 554.400 ;
        RECT 318.000 553.600 318.800 559.800 ;
        RECT 321.200 555.000 322.000 559.800 ;
        RECT 324.400 555.000 325.200 559.800 ;
        RECT 326.000 557.000 326.800 559.800 ;
        RECT 327.600 557.000 328.400 559.800 ;
        RECT 330.800 555.200 331.600 559.800 ;
        RECT 334.000 556.400 334.800 559.800 ;
        RECT 334.000 555.800 335.000 556.400 ;
        RECT 334.400 555.200 335.000 555.800 ;
        RECT 329.600 554.400 333.800 555.200 ;
        RECT 334.400 554.600 336.400 555.200 ;
        RECT 321.200 553.600 323.800 554.400 ;
        RECT 324.400 553.800 330.200 554.400 ;
        RECT 333.200 554.000 333.800 554.400 ;
        RECT 313.200 553.000 314.000 553.200 ;
        RECT 305.000 552.400 314.000 553.000 ;
        RECT 316.400 553.000 317.200 553.200 ;
        RECT 324.400 553.000 325.000 553.800 ;
        RECT 330.800 553.200 332.200 553.800 ;
        RECT 333.200 553.200 334.800 554.000 ;
        RECT 316.400 552.400 325.000 553.000 ;
        RECT 326.000 553.000 332.200 553.200 ;
        RECT 326.000 552.600 331.400 553.000 ;
        RECT 326.000 552.400 326.800 552.600 ;
        RECT 294.000 550.400 295.200 551.200 ;
        RECT 292.400 550.300 293.200 550.400 ;
        RECT 289.400 549.700 293.200 550.300 ;
        RECT 282.800 546.200 283.600 546.800 ;
        RECT 263.600 542.200 264.400 545.400 ;
        RECT 281.200 545.400 283.600 546.200 ;
        RECT 265.200 542.200 266.000 545.000 ;
        RECT 266.800 542.200 267.600 545.000 ;
        RECT 268.400 542.200 269.200 545.000 ;
        RECT 271.600 542.200 272.400 545.000 ;
        RECT 274.800 542.200 275.600 545.000 ;
        RECT 276.400 542.200 277.200 545.000 ;
        RECT 278.000 542.200 278.800 545.000 ;
        RECT 279.600 542.200 280.400 545.000 ;
        RECT 281.200 542.200 282.000 545.400 ;
        RECT 287.600 542.200 288.400 547.400 ;
        RECT 289.400 546.800 290.200 549.700 ;
        RECT 292.400 548.800 293.200 549.700 ;
        RECT 294.000 547.400 294.600 550.400 ;
        RECT 289.200 546.000 290.200 546.800 ;
        RECT 292.400 546.800 294.600 547.400 ;
        RECT 303.400 546.800 304.200 551.200 ;
        RECT 305.000 550.600 305.600 552.400 ;
        RECT 304.800 550.000 305.600 550.600 ;
        RECT 311.600 550.000 335.000 550.600 ;
        RECT 304.800 548.000 305.400 550.000 ;
        RECT 311.600 549.400 312.400 550.000 ;
        RECT 329.200 549.600 330.000 550.000 ;
        RECT 332.400 549.600 333.200 550.000 ;
        RECT 334.200 549.800 335.000 550.000 ;
        RECT 306.000 548.600 309.800 549.400 ;
        RECT 304.800 547.400 306.000 548.000 ;
        RECT 289.200 542.200 290.000 546.000 ;
        RECT 292.400 542.200 293.200 546.800 ;
        RECT 300.400 546.300 301.200 546.400 ;
        RECT 303.400 546.300 304.400 546.800 ;
        RECT 300.400 545.700 304.400 546.300 ;
        RECT 300.400 545.600 301.200 545.700 ;
        RECT 303.600 542.200 304.400 545.700 ;
        RECT 305.200 542.200 306.000 547.400 ;
        RECT 309.000 547.400 309.800 548.600 ;
        RECT 309.000 546.800 310.800 547.400 ;
        RECT 310.000 546.200 310.800 546.800 ;
        RECT 314.800 546.400 315.600 549.200 ;
        RECT 318.000 548.600 321.200 549.400 ;
        RECT 325.000 548.600 327.000 549.400 ;
        RECT 335.600 549.000 336.400 554.600 ;
        RECT 317.600 547.800 318.400 548.000 ;
        RECT 317.600 547.200 322.000 547.800 ;
        RECT 321.200 547.000 322.000 547.200 ;
        RECT 322.800 546.800 323.600 548.400 ;
        RECT 310.000 545.400 312.400 546.200 ;
        RECT 314.800 545.600 315.800 546.400 ;
        RECT 318.800 545.600 320.400 546.400 ;
        RECT 321.200 546.200 322.000 546.400 ;
        RECT 325.000 546.200 325.800 548.600 ;
        RECT 327.600 548.200 336.400 549.000 ;
        RECT 331.000 546.800 334.000 547.600 ;
        RECT 331.000 546.200 331.800 546.800 ;
        RECT 321.200 545.600 325.800 546.200 ;
        RECT 311.600 542.200 312.400 545.400 ;
        RECT 329.200 545.400 331.800 546.200 ;
        RECT 313.200 542.200 314.000 545.000 ;
        RECT 314.800 542.200 315.600 545.000 ;
        RECT 316.400 542.200 317.200 545.000 ;
        RECT 318.000 542.200 318.800 545.000 ;
        RECT 321.200 542.200 322.000 545.000 ;
        RECT 324.400 542.200 325.200 545.000 ;
        RECT 326.000 542.200 326.800 545.000 ;
        RECT 327.600 542.200 328.400 545.000 ;
        RECT 329.200 542.200 330.000 545.400 ;
        RECT 335.600 542.200 336.400 548.200 ;
        RECT 338.800 548.300 339.600 559.800 ;
        RECT 343.000 552.400 343.800 559.800 ;
        RECT 344.400 553.600 345.200 554.400 ;
        RECT 344.600 552.400 345.200 553.600 ;
        RECT 347.600 553.600 348.400 554.400 ;
        RECT 347.600 552.400 348.200 553.600 ;
        RECT 349.000 552.400 349.800 559.800 ;
        RECT 343.000 551.800 344.000 552.400 ;
        RECT 344.600 551.800 346.000 552.400 ;
        RECT 342.000 548.800 342.800 550.400 ;
        RECT 343.400 548.400 344.000 551.800 ;
        RECT 345.200 551.600 346.000 551.800 ;
        RECT 346.800 551.800 348.200 552.400 ;
        RECT 348.800 551.800 349.800 552.400 ;
        RECT 346.800 551.600 347.600 551.800 ;
        RECT 345.300 550.300 345.900 551.600 ;
        RECT 348.800 550.300 349.400 551.800 ;
        RECT 345.300 549.700 349.400 550.300 ;
        RECT 348.800 548.400 349.400 549.700 ;
        RECT 350.000 548.800 350.800 550.400 ;
        RECT 340.400 548.300 341.200 548.400 ;
        RECT 338.800 548.200 341.200 548.300 ;
        RECT 338.800 547.700 342.000 548.200 ;
        RECT 338.800 542.200 339.600 547.700 ;
        RECT 340.400 547.600 342.000 547.700 ;
        RECT 343.400 547.600 346.000 548.400 ;
        RECT 346.800 547.600 349.400 548.400 ;
        RECT 351.600 548.200 352.400 548.400 ;
        RECT 350.800 547.600 352.400 548.200 ;
        RECT 354.800 548.300 355.600 559.800 ;
        RECT 359.000 552.400 359.800 559.800 ;
        RECT 360.400 553.600 361.200 554.400 ;
        RECT 360.600 552.400 361.200 553.600 ;
        RECT 365.400 552.400 366.200 559.800 ;
        RECT 366.800 553.600 367.600 554.400 ;
        RECT 367.000 552.400 367.600 553.600 ;
        RECT 359.000 551.800 360.000 552.400 ;
        RECT 360.600 551.800 362.000 552.400 ;
        RECT 358.000 548.800 358.800 550.400 ;
        RECT 359.400 550.300 360.000 551.800 ;
        RECT 361.200 551.600 362.000 551.800 ;
        RECT 364.400 551.600 366.400 552.400 ;
        RECT 367.000 552.300 368.400 552.400 ;
        RECT 370.800 552.300 371.600 559.800 ;
        RECT 374.000 555.200 374.800 559.800 ;
        RECT 367.000 551.800 371.600 552.300 ;
        RECT 367.600 551.700 371.600 551.800 ;
        RECT 367.600 551.600 368.400 551.700 ;
        RECT 362.800 550.300 363.600 550.400 ;
        RECT 359.400 549.700 363.600 550.300 ;
        RECT 359.400 548.400 360.000 549.700 ;
        RECT 362.800 549.600 363.600 549.700 ;
        RECT 364.400 548.800 365.200 550.400 ;
        RECT 365.800 548.400 366.400 551.600 ;
        RECT 370.600 551.200 371.600 551.700 ;
        RECT 372.200 554.600 374.800 555.200 ;
        RECT 372.200 553.000 372.800 554.600 ;
        RECT 377.200 554.400 378.000 559.800 ;
        RECT 380.400 557.000 381.200 559.800 ;
        RECT 382.000 557.000 382.800 559.800 ;
        RECT 383.600 557.000 384.400 559.800 ;
        RECT 378.600 554.400 382.800 555.200 ;
        RECT 375.400 553.600 378.000 554.400 ;
        RECT 385.200 553.600 386.000 559.800 ;
        RECT 388.400 555.000 389.200 559.800 ;
        RECT 391.600 555.000 392.400 559.800 ;
        RECT 393.200 557.000 394.000 559.800 ;
        RECT 394.800 557.000 395.600 559.800 ;
        RECT 398.000 555.200 398.800 559.800 ;
        RECT 401.200 556.400 402.000 559.800 ;
        RECT 401.200 555.800 402.200 556.400 ;
        RECT 401.600 555.200 402.200 555.800 ;
        RECT 396.800 554.400 401.000 555.200 ;
        RECT 401.600 554.600 403.600 555.200 ;
        RECT 388.400 553.600 391.000 554.400 ;
        RECT 391.600 553.800 397.400 554.400 ;
        RECT 400.400 554.000 401.000 554.400 ;
        RECT 380.400 553.000 381.200 553.200 ;
        RECT 372.200 552.400 381.200 553.000 ;
        RECT 383.600 553.000 384.400 553.200 ;
        RECT 391.600 553.000 392.200 553.800 ;
        RECT 398.000 553.200 399.400 553.800 ;
        RECT 400.400 553.200 402.000 554.000 ;
        RECT 383.600 552.400 392.200 553.000 ;
        RECT 393.200 553.000 399.400 553.200 ;
        RECT 393.200 552.600 398.600 553.000 ;
        RECT 393.200 552.400 394.000 552.600 ;
        RECT 356.400 548.300 357.200 548.400 ;
        RECT 354.800 548.200 357.200 548.300 ;
        RECT 354.800 547.700 358.000 548.200 ;
        RECT 341.200 547.200 342.000 547.600 ;
        RECT 340.600 546.200 344.200 546.600 ;
        RECT 345.200 546.200 345.800 547.600 ;
        RECT 347.000 546.200 347.600 547.600 ;
        RECT 350.800 547.200 351.600 547.600 ;
        RECT 348.600 546.200 352.200 546.600 ;
        RECT 340.400 546.000 344.400 546.200 ;
        RECT 340.400 542.200 341.200 546.000 ;
        RECT 343.600 542.200 344.400 546.000 ;
        RECT 345.200 542.200 346.000 546.200 ;
        RECT 346.800 542.200 347.600 546.200 ;
        RECT 348.400 546.000 352.400 546.200 ;
        RECT 348.400 542.200 349.200 546.000 ;
        RECT 351.600 542.200 352.400 546.000 ;
        RECT 354.800 542.200 355.600 547.700 ;
        RECT 356.400 547.600 358.000 547.700 ;
        RECT 359.400 547.600 362.000 548.400 ;
        RECT 362.800 548.200 363.600 548.400 ;
        RECT 362.800 547.600 364.400 548.200 ;
        RECT 365.800 547.600 368.400 548.400 ;
        RECT 357.200 547.200 358.000 547.600 ;
        RECT 356.600 546.200 360.200 546.600 ;
        RECT 361.200 546.200 361.800 547.600 ;
        RECT 363.600 547.200 364.400 547.600 ;
        RECT 363.000 546.200 366.600 546.600 ;
        RECT 367.600 546.200 368.200 547.600 ;
        RECT 370.600 546.800 371.400 551.200 ;
        RECT 372.200 550.600 372.800 552.400 ;
        RECT 372.000 550.000 372.800 550.600 ;
        RECT 378.800 550.000 402.200 550.600 ;
        RECT 372.000 548.000 372.600 550.000 ;
        RECT 378.800 549.400 379.600 550.000 ;
        RECT 396.400 549.600 397.200 550.000 ;
        RECT 399.600 549.600 400.400 550.000 ;
        RECT 401.400 549.800 402.200 550.000 ;
        RECT 373.200 548.600 377.000 549.400 ;
        RECT 372.000 547.400 373.200 548.000 ;
        RECT 356.400 546.000 360.400 546.200 ;
        RECT 356.400 542.200 357.200 546.000 ;
        RECT 359.600 542.200 360.400 546.000 ;
        RECT 361.200 542.200 362.000 546.200 ;
        RECT 362.800 546.000 366.800 546.200 ;
        RECT 362.800 542.200 363.600 546.000 ;
        RECT 366.000 542.200 366.800 546.000 ;
        RECT 367.600 542.200 368.400 546.200 ;
        RECT 370.600 546.000 371.600 546.800 ;
        RECT 370.800 542.200 371.600 546.000 ;
        RECT 372.400 542.200 373.200 547.400 ;
        RECT 376.200 547.400 377.000 548.600 ;
        RECT 376.200 546.800 378.000 547.400 ;
        RECT 377.200 546.200 378.000 546.800 ;
        RECT 382.000 546.400 382.800 549.200 ;
        RECT 385.200 548.600 388.400 549.400 ;
        RECT 392.200 548.600 394.200 549.400 ;
        RECT 402.800 549.000 403.600 554.600 ;
        RECT 406.000 551.200 406.800 559.800 ;
        RECT 409.200 551.200 410.000 559.800 ;
        RECT 412.400 551.200 413.200 559.800 ;
        RECT 415.600 551.200 416.400 559.800 ;
        RECT 384.800 547.800 385.600 548.000 ;
        RECT 384.800 547.200 389.200 547.800 ;
        RECT 388.400 547.000 389.200 547.200 ;
        RECT 390.000 546.800 390.800 548.400 ;
        RECT 377.200 545.400 379.600 546.200 ;
        RECT 382.000 545.600 383.000 546.400 ;
        RECT 386.000 545.600 387.600 546.400 ;
        RECT 388.400 546.200 389.200 546.400 ;
        RECT 392.200 546.200 393.000 548.600 ;
        RECT 394.800 548.200 403.600 549.000 ;
        RECT 398.200 546.800 401.200 547.600 ;
        RECT 398.200 546.200 399.000 546.800 ;
        RECT 388.400 545.600 393.000 546.200 ;
        RECT 378.800 542.200 379.600 545.400 ;
        RECT 396.400 545.400 399.000 546.200 ;
        RECT 380.400 542.200 381.200 545.000 ;
        RECT 382.000 542.200 382.800 545.000 ;
        RECT 383.600 542.200 384.400 545.000 ;
        RECT 385.200 542.200 386.000 545.000 ;
        RECT 388.400 542.200 389.200 545.000 ;
        RECT 391.600 542.200 392.400 545.000 ;
        RECT 393.200 542.200 394.000 545.000 ;
        RECT 394.800 542.200 395.600 545.000 ;
        RECT 396.400 542.200 397.200 545.400 ;
        RECT 402.800 542.200 403.600 548.200 ;
        RECT 404.400 550.400 406.800 551.200 ;
        RECT 407.800 550.400 410.000 551.200 ;
        RECT 411.000 550.400 413.200 551.200 ;
        RECT 414.600 550.400 416.400 551.200 ;
        RECT 418.800 551.200 419.600 559.800 ;
        RECT 423.000 555.800 424.200 559.800 ;
        RECT 427.600 555.800 428.400 559.800 ;
        RECT 432.000 556.400 432.800 559.800 ;
        RECT 432.000 555.800 434.000 556.400 ;
        RECT 423.600 555.000 424.400 555.800 ;
        RECT 427.800 555.200 428.400 555.800 ;
        RECT 427.000 554.600 430.600 555.200 ;
        RECT 433.200 555.000 434.000 555.800 ;
        RECT 427.000 554.400 427.800 554.600 ;
        RECT 429.800 554.400 430.600 554.600 ;
        RECT 422.800 553.200 424.200 554.000 ;
        RECT 423.600 552.200 424.200 553.200 ;
        RECT 425.800 553.000 428.000 553.600 ;
        RECT 425.800 552.800 426.600 553.000 ;
        RECT 423.600 551.600 426.000 552.200 ;
        RECT 418.800 550.600 423.000 551.200 ;
        RECT 404.400 547.600 405.200 550.400 ;
        RECT 407.800 549.000 408.600 550.400 ;
        RECT 411.000 549.000 411.800 550.400 ;
        RECT 414.600 549.000 415.400 550.400 ;
        RECT 406.000 548.200 408.600 549.000 ;
        RECT 409.400 548.200 411.800 549.000 ;
        RECT 412.800 548.200 415.400 549.000 ;
        RECT 416.200 548.200 418.000 549.000 ;
        RECT 407.800 547.600 408.600 548.200 ;
        RECT 411.000 547.600 411.800 548.200 ;
        RECT 414.600 547.600 415.400 548.200 ;
        RECT 417.200 547.600 418.000 548.200 ;
        RECT 404.400 546.800 406.800 547.600 ;
        RECT 407.800 546.800 410.000 547.600 ;
        RECT 411.000 546.800 413.200 547.600 ;
        RECT 414.600 546.800 416.400 547.600 ;
        RECT 406.000 542.200 406.800 546.800 ;
        RECT 409.200 542.200 410.000 546.800 ;
        RECT 412.400 542.200 413.200 546.800 ;
        RECT 415.600 542.200 416.400 546.800 ;
        RECT 418.800 547.200 419.600 550.600 ;
        RECT 422.200 550.400 423.000 550.600 ;
        RECT 425.400 550.400 426.000 551.600 ;
        RECT 427.400 551.800 428.000 553.000 ;
        RECT 428.600 553.000 429.400 553.200 ;
        RECT 433.200 553.000 434.000 553.200 ;
        RECT 428.600 552.400 434.000 553.000 ;
        RECT 427.400 551.400 432.200 551.800 ;
        RECT 436.400 551.400 437.200 559.800 ;
        RECT 440.600 552.400 441.400 559.800 ;
        RECT 442.000 553.600 442.800 554.400 ;
        RECT 442.200 552.400 442.800 553.600 ;
        RECT 445.200 553.600 446.000 554.400 ;
        RECT 445.200 552.400 445.800 553.600 ;
        RECT 446.600 552.400 447.400 559.800 ;
        RECT 451.400 552.400 452.200 559.800 ;
        RECT 440.600 551.800 441.600 552.400 ;
        RECT 442.200 551.800 443.600 552.400 ;
        RECT 427.400 551.200 437.200 551.400 ;
        RECT 431.400 551.000 437.200 551.200 ;
        RECT 431.600 550.800 437.200 551.000 ;
        RECT 441.000 550.400 441.600 551.800 ;
        RECT 442.800 551.600 443.600 551.800 ;
        RECT 444.400 551.800 445.800 552.400 ;
        RECT 446.400 551.800 447.400 552.400 ;
        RECT 450.800 551.800 452.200 552.400 ;
        RECT 444.400 551.600 445.200 551.800 ;
        RECT 420.600 549.800 421.400 550.000 ;
        RECT 420.600 549.200 424.400 549.800 ;
        RECT 425.200 549.600 426.000 550.400 ;
        RECT 430.000 550.200 430.800 550.400 ;
        RECT 430.000 549.600 435.000 550.200 ;
        RECT 423.600 549.000 424.400 549.200 ;
        RECT 425.400 548.400 426.000 549.600 ;
        RECT 431.600 549.400 432.400 549.600 ;
        RECT 434.200 549.400 435.000 549.600 ;
        RECT 439.600 548.800 440.400 550.400 ;
        RECT 441.000 549.600 442.000 550.400 ;
        RECT 442.900 550.300 443.500 551.600 ;
        RECT 446.400 550.300 447.000 551.800 ;
        RECT 450.800 550.400 451.400 551.800 ;
        RECT 455.600 551.200 456.400 559.800 ;
        RECT 452.400 550.800 456.400 551.200 ;
        RECT 452.200 550.600 456.400 550.800 ;
        RECT 462.000 551.200 462.800 559.800 ;
        RECT 466.200 555.800 467.400 559.800 ;
        RECT 470.800 555.800 471.600 559.800 ;
        RECT 475.200 556.400 476.000 559.800 ;
        RECT 475.200 555.800 477.200 556.400 ;
        RECT 466.800 555.000 467.600 555.800 ;
        RECT 471.000 555.200 471.600 555.800 ;
        RECT 470.200 554.600 473.800 555.200 ;
        RECT 476.400 555.000 477.200 555.800 ;
        RECT 470.200 554.400 471.000 554.600 ;
        RECT 473.000 554.400 473.800 554.600 ;
        RECT 466.000 553.200 467.400 554.000 ;
        RECT 466.800 552.200 467.400 553.200 ;
        RECT 469.000 553.000 471.200 553.600 ;
        RECT 469.000 552.800 469.800 553.000 ;
        RECT 466.800 551.600 469.200 552.200 ;
        RECT 462.000 550.600 466.200 551.200 ;
        RECT 442.900 549.700 447.000 550.300 ;
        RECT 432.600 548.400 433.400 548.600 ;
        RECT 441.000 548.400 441.600 549.600 ;
        RECT 446.400 548.400 447.000 549.700 ;
        RECT 447.600 548.800 448.400 550.400 ;
        RECT 450.800 549.600 451.600 550.400 ;
        RECT 452.200 550.000 453.000 550.600 ;
        RECT 425.400 547.800 436.400 548.400 ;
        RECT 425.800 547.600 426.600 547.800 ;
        RECT 418.800 546.600 422.600 547.200 ;
        RECT 418.800 542.200 419.600 546.600 ;
        RECT 421.800 546.400 422.600 546.600 ;
        RECT 431.600 545.600 432.200 547.800 ;
        RECT 434.800 547.600 436.400 547.800 ;
        RECT 438.000 548.200 438.800 548.400 ;
        RECT 438.000 547.600 439.600 548.200 ;
        RECT 441.000 547.600 443.600 548.400 ;
        RECT 444.400 547.600 447.000 548.400 ;
        RECT 449.200 548.200 450.000 548.400 ;
        RECT 448.400 547.600 450.000 548.200 ;
        RECT 438.800 547.200 439.600 547.600 ;
        RECT 429.800 545.400 430.600 545.600 ;
        RECT 423.600 544.200 424.400 545.000 ;
        RECT 427.800 544.800 430.600 545.400 ;
        RECT 431.600 544.800 432.400 545.600 ;
        RECT 427.800 544.200 428.400 544.800 ;
        RECT 433.200 544.200 434.000 545.000 ;
        RECT 423.000 543.600 424.400 544.200 ;
        RECT 423.000 542.200 424.200 543.600 ;
        RECT 427.600 542.200 428.400 544.200 ;
        RECT 432.000 543.600 434.000 544.200 ;
        RECT 432.000 542.200 432.800 543.600 ;
        RECT 436.400 542.200 437.200 547.000 ;
        RECT 438.200 546.200 441.800 546.600 ;
        RECT 442.800 546.200 443.400 547.600 ;
        RECT 444.600 546.200 445.200 547.600 ;
        RECT 448.400 547.200 449.200 547.600 ;
        RECT 446.200 546.200 449.800 546.600 ;
        RECT 450.800 546.200 451.400 549.600 ;
        RECT 452.200 547.000 452.800 550.000 ;
        RECT 453.600 548.400 454.400 549.200 ;
        RECT 453.800 548.300 454.800 548.400 ;
        RECT 457.200 548.300 458.000 548.400 ;
        RECT 453.800 547.700 458.000 548.300 ;
        RECT 453.800 547.600 454.800 547.700 ;
        RECT 457.200 547.600 458.000 547.700 ;
        RECT 462.000 547.200 462.800 550.600 ;
        RECT 465.400 550.400 466.200 550.600 ;
        RECT 468.600 550.400 469.200 551.600 ;
        RECT 470.600 551.800 471.200 553.000 ;
        RECT 471.800 553.000 472.600 553.200 ;
        RECT 476.400 553.000 477.200 553.200 ;
        RECT 471.800 552.400 477.200 553.000 ;
        RECT 470.600 551.400 475.400 551.800 ;
        RECT 479.600 551.400 480.400 559.800 ;
        RECT 483.800 552.400 484.600 559.800 ;
        RECT 485.200 553.600 486.000 554.400 ;
        RECT 485.400 552.400 486.000 553.600 ;
        RECT 488.400 553.600 489.200 554.400 ;
        RECT 488.400 552.400 489.000 553.600 ;
        RECT 489.800 552.400 490.600 559.800 ;
        RECT 483.800 551.800 484.800 552.400 ;
        RECT 485.400 551.800 486.800 552.400 ;
        RECT 470.600 551.200 480.400 551.400 ;
        RECT 474.600 551.000 480.400 551.200 ;
        RECT 474.800 550.800 480.400 551.000 ;
        RECT 463.800 549.800 464.600 550.000 ;
        RECT 463.800 549.200 467.600 549.800 ;
        RECT 468.400 549.600 469.200 550.400 ;
        RECT 473.200 550.200 474.000 550.400 ;
        RECT 473.200 549.600 478.200 550.200 ;
        RECT 466.800 549.000 467.600 549.200 ;
        RECT 468.600 548.400 469.200 549.600 ;
        RECT 474.800 549.400 475.600 549.600 ;
        RECT 477.400 549.400 478.200 549.600 ;
        RECT 482.800 548.800 483.600 550.400 ;
        RECT 475.800 548.400 476.600 548.600 ;
        RECT 484.200 548.400 484.800 551.800 ;
        RECT 486.000 551.600 486.800 551.800 ;
        RECT 487.600 551.800 489.000 552.400 ;
        RECT 489.600 551.800 490.600 552.400 ;
        RECT 487.600 551.600 488.400 551.800 ;
        RECT 486.100 550.300 486.700 551.600 ;
        RECT 489.600 550.300 490.200 551.800 ;
        RECT 494.000 551.200 494.800 559.800 ;
        RECT 498.200 555.800 499.400 559.800 ;
        RECT 502.800 555.800 503.600 559.800 ;
        RECT 507.200 556.400 508.000 559.800 ;
        RECT 507.200 555.800 509.200 556.400 ;
        RECT 498.800 555.000 499.600 555.800 ;
        RECT 503.000 555.200 503.600 555.800 ;
        RECT 502.200 554.600 505.800 555.200 ;
        RECT 508.400 555.000 509.200 555.800 ;
        RECT 502.200 554.400 503.000 554.600 ;
        RECT 505.000 554.400 505.800 554.600 ;
        RECT 498.000 553.200 499.400 554.000 ;
        RECT 498.800 552.200 499.400 553.200 ;
        RECT 501.000 553.000 503.200 553.600 ;
        RECT 501.000 552.800 501.800 553.000 ;
        RECT 498.800 551.600 501.200 552.200 ;
        RECT 494.000 550.600 498.200 551.200 ;
        RECT 486.100 549.700 490.200 550.300 ;
        RECT 489.600 548.400 490.200 549.700 ;
        RECT 490.800 548.800 491.600 550.400 ;
        RECT 468.600 547.800 479.600 548.400 ;
        RECT 469.000 547.600 469.800 547.800 ;
        RECT 452.200 546.400 454.600 547.000 ;
        RECT 462.000 546.600 465.800 547.200 ;
        RECT 438.000 546.000 442.000 546.200 ;
        RECT 438.000 542.200 438.800 546.000 ;
        RECT 441.200 542.200 442.000 546.000 ;
        RECT 442.800 542.200 443.600 546.200 ;
        RECT 444.400 542.200 445.200 546.200 ;
        RECT 446.000 546.000 450.000 546.200 ;
        RECT 446.000 542.200 446.800 546.000 ;
        RECT 449.200 542.200 450.000 546.000 ;
        RECT 450.800 542.200 451.600 546.200 ;
        RECT 454.000 544.200 454.600 546.400 ;
        RECT 455.600 544.800 456.400 546.400 ;
        RECT 458.800 544.300 459.600 544.400 ;
        RECT 462.000 544.300 462.800 546.600 ;
        RECT 465.000 546.400 465.800 546.600 ;
        RECT 474.800 545.600 475.400 547.800 ;
        RECT 478.000 547.600 479.600 547.800 ;
        RECT 481.200 548.200 482.000 548.400 ;
        RECT 481.200 547.600 482.800 548.200 ;
        RECT 484.200 547.600 486.800 548.400 ;
        RECT 487.600 547.600 490.200 548.400 ;
        RECT 492.400 548.200 493.200 548.400 ;
        RECT 491.600 547.600 493.200 548.200 ;
        RECT 482.000 547.200 482.800 547.600 ;
        RECT 473.000 545.400 473.800 545.600 ;
        RECT 454.000 542.200 454.800 544.200 ;
        RECT 458.800 543.700 462.800 544.300 ;
        RECT 466.800 544.200 467.600 545.000 ;
        RECT 471.000 544.800 473.800 545.400 ;
        RECT 474.800 544.800 475.600 545.600 ;
        RECT 471.000 544.200 471.600 544.800 ;
        RECT 476.400 544.200 477.200 545.000 ;
        RECT 458.800 543.600 459.600 543.700 ;
        RECT 462.000 542.200 462.800 543.700 ;
        RECT 466.200 543.600 467.600 544.200 ;
        RECT 466.200 542.200 467.400 543.600 ;
        RECT 470.800 542.200 471.600 544.200 ;
        RECT 475.200 543.600 477.200 544.200 ;
        RECT 475.200 542.200 476.000 543.600 ;
        RECT 479.600 542.200 480.400 547.000 ;
        RECT 481.400 546.200 485.000 546.600 ;
        RECT 486.000 546.200 486.600 547.600 ;
        RECT 487.800 546.200 488.400 547.600 ;
        RECT 491.600 547.200 492.400 547.600 ;
        RECT 494.000 547.200 494.800 550.600 ;
        RECT 497.400 550.400 498.200 550.600 ;
        RECT 495.800 549.800 496.600 550.000 ;
        RECT 495.800 549.200 499.600 549.800 ;
        RECT 498.800 549.000 499.600 549.200 ;
        RECT 500.600 548.400 501.200 551.600 ;
        RECT 502.600 551.800 503.200 553.000 ;
        RECT 503.800 553.000 504.600 553.200 ;
        RECT 508.400 553.000 509.200 553.200 ;
        RECT 503.800 552.400 509.200 553.000 ;
        RECT 502.600 551.400 507.400 551.800 ;
        RECT 511.600 551.400 512.400 559.800 ;
        RECT 515.800 552.400 516.600 559.800 ;
        RECT 519.600 555.000 520.400 559.000 ;
        RECT 517.200 553.600 518.000 554.400 ;
        RECT 517.400 552.400 518.000 553.600 ;
        RECT 515.800 551.800 516.800 552.400 ;
        RECT 517.400 551.800 518.800 552.400 ;
        RECT 502.600 551.200 512.400 551.400 ;
        RECT 506.600 551.000 512.400 551.200 ;
        RECT 506.800 550.800 512.400 551.000 ;
        RECT 505.200 550.200 506.000 550.400 ;
        RECT 505.200 549.600 510.200 550.200 ;
        RECT 509.400 549.400 510.200 549.600 ;
        RECT 514.800 548.800 515.600 550.400 ;
        RECT 507.800 548.400 508.600 548.600 ;
        RECT 516.200 548.400 516.800 551.800 ;
        RECT 518.000 551.600 518.800 551.800 ;
        RECT 519.600 551.600 520.200 555.000 ;
        RECT 523.800 552.800 524.600 559.800 ;
        RECT 530.000 553.600 530.800 554.400 ;
        RECT 523.800 552.200 525.400 552.800 ;
        RECT 530.000 552.400 530.600 553.600 ;
        RECT 531.400 552.400 532.200 559.800 ;
        RECT 519.600 551.000 523.400 551.600 ;
        RECT 519.600 548.800 520.400 550.400 ;
        RECT 521.200 548.800 522.000 550.400 ;
        RECT 522.800 549.000 523.400 551.000 ;
        RECT 500.600 547.800 511.600 548.400 ;
        RECT 501.000 547.600 501.800 547.800 ;
        RECT 494.000 546.600 497.800 547.200 ;
        RECT 489.400 546.200 493.000 546.600 ;
        RECT 481.200 546.000 485.200 546.200 ;
        RECT 481.200 542.200 482.000 546.000 ;
        RECT 484.400 542.200 485.200 546.000 ;
        RECT 486.000 542.200 486.800 546.200 ;
        RECT 487.600 542.200 488.400 546.200 ;
        RECT 489.200 546.000 493.200 546.200 ;
        RECT 489.200 542.200 490.000 546.000 ;
        RECT 492.400 542.200 493.200 546.000 ;
        RECT 494.000 542.200 494.800 546.600 ;
        RECT 497.000 546.400 497.800 546.600 ;
        RECT 506.800 545.600 507.400 547.800 ;
        RECT 510.000 547.600 511.600 547.800 ;
        RECT 513.200 548.200 514.000 548.400 ;
        RECT 513.200 547.600 514.800 548.200 ;
        RECT 516.200 547.600 518.800 548.400 ;
        RECT 522.800 548.200 524.200 549.000 ;
        RECT 524.800 548.400 525.400 552.200 ;
        RECT 529.200 551.800 530.600 552.400 ;
        RECT 529.200 551.600 530.000 551.800 ;
        RECT 531.200 551.600 533.200 552.400 ;
        RECT 526.000 549.600 526.800 551.200 ;
        RECT 531.200 548.400 531.800 551.600 ;
        RECT 532.400 548.800 533.200 550.400 ;
        RECT 524.800 548.300 526.800 548.400 ;
        RECT 527.600 548.300 528.400 548.400 ;
        RECT 522.800 547.800 523.800 548.200 ;
        RECT 514.000 547.200 514.800 547.600 ;
        RECT 505.000 545.400 505.800 545.600 ;
        RECT 498.800 544.200 499.600 545.000 ;
        RECT 503.000 544.800 505.800 545.400 ;
        RECT 506.800 544.800 507.600 545.600 ;
        RECT 503.000 544.200 503.600 544.800 ;
        RECT 508.400 544.200 509.200 545.000 ;
        RECT 498.200 543.600 499.600 544.200 ;
        RECT 498.200 542.200 499.400 543.600 ;
        RECT 502.800 542.200 503.600 544.200 ;
        RECT 507.200 543.600 509.200 544.200 ;
        RECT 507.200 542.200 508.000 543.600 ;
        RECT 511.600 542.200 512.400 547.000 ;
        RECT 513.400 546.200 517.000 546.600 ;
        RECT 518.000 546.200 518.600 547.600 ;
        RECT 519.600 547.200 523.800 547.800 ;
        RECT 524.800 547.700 528.400 548.300 ;
        RECT 524.800 547.600 526.800 547.700 ;
        RECT 527.600 547.600 528.400 547.700 ;
        RECT 529.200 547.600 531.800 548.400 ;
        RECT 534.000 548.200 534.800 548.400 ;
        RECT 533.200 547.600 534.800 548.200 ;
        RECT 513.200 546.000 517.200 546.200 ;
        RECT 513.200 542.200 514.000 546.000 ;
        RECT 516.400 542.200 517.200 546.000 ;
        RECT 518.000 542.200 518.800 546.200 ;
        RECT 519.600 545.000 520.200 547.200 ;
        RECT 524.800 547.000 525.400 547.600 ;
        RECT 524.600 546.600 525.400 547.000 ;
        RECT 523.800 546.000 525.400 546.600 ;
        RECT 529.400 546.200 530.000 547.600 ;
        RECT 533.200 547.200 534.000 547.600 ;
        RECT 531.000 546.200 534.600 546.600 ;
        RECT 519.600 543.000 520.400 545.000 ;
        RECT 523.800 543.000 524.600 546.000 ;
        RECT 529.200 542.200 530.000 546.200 ;
        RECT 530.800 546.000 534.800 546.200 ;
        RECT 530.800 542.200 531.600 546.000 ;
        RECT 534.000 542.200 534.800 546.000 ;
        RECT 537.200 542.200 538.000 559.800 ;
        RECT 538.800 551.200 539.600 559.800 ;
        RECT 543.000 555.800 544.200 559.800 ;
        RECT 547.600 555.800 548.400 559.800 ;
        RECT 552.000 556.400 552.800 559.800 ;
        RECT 552.000 555.800 554.000 556.400 ;
        RECT 543.600 555.000 544.400 555.800 ;
        RECT 547.800 555.200 548.400 555.800 ;
        RECT 547.000 554.600 550.600 555.200 ;
        RECT 553.200 555.000 554.000 555.800 ;
        RECT 547.000 554.400 547.800 554.600 ;
        RECT 549.800 554.400 550.600 554.600 ;
        RECT 542.800 553.200 544.200 554.000 ;
        RECT 543.600 552.200 544.200 553.200 ;
        RECT 545.800 553.000 548.000 553.600 ;
        RECT 545.800 552.800 546.600 553.000 ;
        RECT 543.600 551.600 546.000 552.200 ;
        RECT 538.800 550.600 543.000 551.200 ;
        RECT 538.800 547.200 539.600 550.600 ;
        RECT 542.200 550.400 543.000 550.600 ;
        RECT 540.600 549.800 541.400 550.000 ;
        RECT 540.600 549.200 544.400 549.800 ;
        RECT 543.600 549.000 544.400 549.200 ;
        RECT 545.400 548.400 546.000 551.600 ;
        RECT 547.400 551.800 548.000 553.000 ;
        RECT 548.600 553.000 549.400 553.200 ;
        RECT 553.200 553.000 554.000 553.200 ;
        RECT 548.600 552.400 554.000 553.000 ;
        RECT 547.400 551.400 552.200 551.800 ;
        RECT 556.400 551.400 557.200 559.800 ;
        RECT 559.600 552.000 560.400 559.800 ;
        RECT 562.800 555.200 563.600 559.800 ;
        RECT 547.400 551.200 557.200 551.400 ;
        RECT 551.400 551.000 557.200 551.200 ;
        RECT 551.600 550.800 557.200 551.000 ;
        RECT 559.400 551.200 560.400 552.000 ;
        RECT 561.000 554.600 563.600 555.200 ;
        RECT 561.000 553.000 561.600 554.600 ;
        RECT 566.000 554.400 566.800 559.800 ;
        RECT 569.200 557.000 570.000 559.800 ;
        RECT 570.800 557.000 571.600 559.800 ;
        RECT 572.400 557.000 573.200 559.800 ;
        RECT 567.400 554.400 571.600 555.200 ;
        RECT 564.200 553.600 566.800 554.400 ;
        RECT 574.000 553.600 574.800 559.800 ;
        RECT 577.200 555.000 578.000 559.800 ;
        RECT 580.400 555.000 581.200 559.800 ;
        RECT 582.000 557.000 582.800 559.800 ;
        RECT 583.600 557.000 584.400 559.800 ;
        RECT 586.800 555.200 587.600 559.800 ;
        RECT 590.000 556.400 590.800 559.800 ;
        RECT 590.000 555.800 591.000 556.400 ;
        RECT 590.400 555.200 591.000 555.800 ;
        RECT 585.600 554.400 589.800 555.200 ;
        RECT 590.400 554.600 592.400 555.200 ;
        RECT 577.200 553.600 579.800 554.400 ;
        RECT 580.400 553.800 586.200 554.400 ;
        RECT 589.200 554.000 589.800 554.400 ;
        RECT 569.200 553.000 570.000 553.200 ;
        RECT 561.000 552.400 570.000 553.000 ;
        RECT 572.400 553.000 573.200 553.200 ;
        RECT 580.400 553.000 581.000 553.800 ;
        RECT 586.800 553.200 588.200 553.800 ;
        RECT 589.200 553.200 590.800 554.000 ;
        RECT 572.400 552.400 581.000 553.000 ;
        RECT 582.000 553.000 588.200 553.200 ;
        RECT 582.000 552.600 587.400 553.000 ;
        RECT 582.000 552.400 582.800 552.600 ;
        RECT 550.000 550.200 550.800 550.400 ;
        RECT 550.000 549.600 555.000 550.200 ;
        RECT 554.200 549.400 555.000 549.600 ;
        RECT 552.600 548.400 553.400 548.600 ;
        RECT 545.200 547.800 556.400 548.400 ;
        RECT 545.200 547.600 546.600 547.800 ;
        RECT 538.800 546.600 542.600 547.200 ;
        RECT 538.800 542.200 539.600 546.600 ;
        RECT 541.800 546.400 542.600 546.600 ;
        RECT 551.600 545.600 552.200 547.800 ;
        RECT 554.800 547.600 556.400 547.800 ;
        RECT 549.800 545.400 550.600 545.600 ;
        RECT 543.600 544.200 544.400 545.000 ;
        RECT 547.800 544.800 550.600 545.400 ;
        RECT 551.600 544.800 552.400 545.600 ;
        RECT 547.800 544.200 548.400 544.800 ;
        RECT 553.200 544.200 554.000 545.000 ;
        RECT 543.000 543.600 544.400 544.200 ;
        RECT 543.000 542.200 544.200 543.600 ;
        RECT 547.600 542.200 548.400 544.200 ;
        RECT 552.000 543.600 554.000 544.200 ;
        RECT 552.000 542.200 552.800 543.600 ;
        RECT 556.400 542.200 557.200 547.000 ;
        RECT 559.400 546.800 560.200 551.200 ;
        RECT 561.000 550.600 561.600 552.400 ;
        RECT 560.800 550.000 561.600 550.600 ;
        RECT 567.600 550.000 591.000 550.600 ;
        RECT 560.800 548.000 561.400 550.000 ;
        RECT 567.600 549.400 568.400 550.000 ;
        RECT 585.200 549.600 586.000 550.000 ;
        RECT 588.400 549.600 589.200 550.000 ;
        RECT 590.200 549.800 591.000 550.000 ;
        RECT 562.000 548.600 565.800 549.400 ;
        RECT 560.800 547.400 562.000 548.000 ;
        RECT 559.400 546.000 560.400 546.800 ;
        RECT 559.600 542.200 560.400 546.000 ;
        RECT 561.200 542.200 562.000 547.400 ;
        RECT 565.000 547.400 565.800 548.600 ;
        RECT 565.000 546.800 566.800 547.400 ;
        RECT 566.000 546.200 566.800 546.800 ;
        RECT 570.800 546.400 571.600 549.200 ;
        RECT 574.000 548.600 577.200 549.400 ;
        RECT 581.000 548.600 583.000 549.400 ;
        RECT 591.600 549.000 592.400 554.600 ;
        RECT 573.600 547.800 574.400 548.000 ;
        RECT 573.600 547.200 578.000 547.800 ;
        RECT 577.200 547.000 578.000 547.200 ;
        RECT 578.800 546.800 579.600 548.400 ;
        RECT 566.000 545.400 568.400 546.200 ;
        RECT 570.800 545.600 571.800 546.400 ;
        RECT 574.800 545.600 576.400 546.400 ;
        RECT 577.200 546.200 578.000 546.400 ;
        RECT 581.000 546.200 581.800 548.600 ;
        RECT 583.600 548.200 592.400 549.000 ;
        RECT 587.000 546.800 590.000 547.600 ;
        RECT 587.000 546.200 587.800 546.800 ;
        RECT 577.200 545.600 581.800 546.200 ;
        RECT 567.600 542.200 568.400 545.400 ;
        RECT 585.200 545.400 587.800 546.200 ;
        RECT 569.200 542.200 570.000 545.000 ;
        RECT 570.800 542.200 571.600 545.000 ;
        RECT 572.400 542.200 573.200 545.000 ;
        RECT 574.000 542.200 574.800 545.000 ;
        RECT 577.200 542.200 578.000 545.000 ;
        RECT 580.400 542.200 581.200 545.000 ;
        RECT 582.000 542.200 582.800 545.000 ;
        RECT 583.600 542.200 584.400 545.000 ;
        RECT 585.200 542.200 586.000 545.400 ;
        RECT 591.600 542.200 592.400 548.200 ;
        RECT 593.200 542.200 594.000 559.800 ;
        RECT 598.000 551.200 598.800 559.800 ;
        RECT 601.200 551.200 602.000 559.800 ;
        RECT 604.400 551.200 605.200 559.800 ;
        RECT 607.600 551.200 608.400 559.800 ;
        RECT 598.000 550.400 599.800 551.200 ;
        RECT 601.200 550.400 603.400 551.200 ;
        RECT 604.400 550.400 606.600 551.200 ;
        RECT 607.600 550.400 610.000 551.200 ;
        RECT 599.000 549.000 599.800 550.400 ;
        RECT 602.600 549.000 603.400 550.400 ;
        RECT 605.800 549.000 606.600 550.400 ;
        RECT 596.400 548.200 598.200 549.000 ;
        RECT 599.000 548.200 601.600 549.000 ;
        RECT 602.600 548.200 605.000 549.000 ;
        RECT 605.800 548.200 608.400 549.000 ;
        RECT 596.400 547.600 597.200 548.200 ;
        RECT 599.000 547.600 599.800 548.200 ;
        RECT 602.600 547.600 603.400 548.200 ;
        RECT 605.800 547.600 606.600 548.200 ;
        RECT 609.200 547.600 610.000 550.400 ;
        RECT 598.000 546.800 599.800 547.600 ;
        RECT 601.200 546.800 603.400 547.600 ;
        RECT 604.400 546.800 606.600 547.600 ;
        RECT 607.600 546.800 610.000 547.600 ;
        RECT 594.800 544.800 595.600 546.400 ;
        RECT 598.000 542.200 598.800 546.800 ;
        RECT 601.200 542.200 602.000 546.800 ;
        RECT 604.400 542.200 605.200 546.800 ;
        RECT 607.600 542.200 608.400 546.800 ;
        RECT 1.200 533.800 2.000 539.800 ;
        RECT 7.600 536.600 8.400 539.800 ;
        RECT 9.200 537.000 10.000 539.800 ;
        RECT 10.800 537.000 11.600 539.800 ;
        RECT 12.400 537.000 13.200 539.800 ;
        RECT 15.600 537.000 16.400 539.800 ;
        RECT 18.800 537.000 19.600 539.800 ;
        RECT 20.400 537.000 21.200 539.800 ;
        RECT 22.000 537.000 22.800 539.800 ;
        RECT 23.600 537.000 24.400 539.800 ;
        RECT 5.800 535.800 8.400 536.600 ;
        RECT 25.200 536.600 26.000 539.800 ;
        RECT 11.800 535.800 16.400 536.400 ;
        RECT 5.800 535.200 6.600 535.800 ;
        RECT 3.600 534.400 6.600 535.200 ;
        RECT 1.200 533.000 10.000 533.800 ;
        RECT 11.800 533.400 12.600 535.800 ;
        RECT 15.600 535.600 16.400 535.800 ;
        RECT 17.200 535.600 18.800 536.400 ;
        RECT 21.800 535.600 22.800 536.400 ;
        RECT 25.200 535.800 27.600 536.600 ;
        RECT 14.000 533.600 14.800 535.200 ;
        RECT 15.600 534.800 16.400 535.000 ;
        RECT 15.600 534.200 20.000 534.800 ;
        RECT 19.200 534.000 20.000 534.200 ;
        RECT 1.200 527.400 2.000 533.000 ;
        RECT 10.600 532.600 12.600 533.400 ;
        RECT 16.400 532.600 19.600 533.400 ;
        RECT 22.000 532.800 22.800 535.600 ;
        RECT 26.800 535.200 27.600 535.800 ;
        RECT 26.800 534.600 28.600 535.200 ;
        RECT 27.800 533.400 28.600 534.600 ;
        RECT 31.600 534.600 32.400 539.800 ;
        RECT 33.200 536.000 34.000 539.800 ;
        RECT 33.200 535.200 34.200 536.000 ;
        RECT 36.400 535.800 37.200 539.800 ;
        RECT 38.000 536.000 38.800 539.800 ;
        RECT 41.200 536.000 42.000 539.800 ;
        RECT 43.400 536.400 44.200 539.800 ;
        RECT 38.000 535.800 42.000 536.000 ;
        RECT 31.600 534.000 32.800 534.600 ;
        RECT 27.800 532.600 31.600 533.400 ;
        RECT 2.600 532.000 3.400 532.200 ;
        RECT 6.000 532.000 6.800 532.400 ;
        RECT 7.600 532.000 8.400 532.400 ;
        RECT 25.200 532.000 26.000 532.600 ;
        RECT 32.200 532.000 32.800 534.000 ;
        RECT 2.600 531.400 26.000 532.000 ;
        RECT 32.000 531.400 32.800 532.000 ;
        RECT 32.000 529.600 32.600 531.400 ;
        RECT 33.400 530.800 34.200 535.200 ;
        RECT 36.600 534.400 37.200 535.800 ;
        RECT 38.200 535.400 41.800 535.800 ;
        RECT 42.800 535.600 45.200 536.400 ;
        RECT 40.400 534.400 41.200 534.800 ;
        RECT 36.400 533.600 39.000 534.400 ;
        RECT 40.400 533.800 42.000 534.400 ;
        RECT 41.200 533.600 42.000 533.800 ;
        RECT 10.800 529.400 11.600 529.600 ;
        RECT 6.200 529.000 11.600 529.400 ;
        RECT 5.400 528.800 11.600 529.000 ;
        RECT 12.600 529.000 21.200 529.600 ;
        RECT 2.800 528.000 4.400 528.800 ;
        RECT 5.400 528.200 6.800 528.800 ;
        RECT 12.600 528.200 13.200 529.000 ;
        RECT 20.400 528.800 21.200 529.000 ;
        RECT 23.600 529.000 32.600 529.600 ;
        RECT 23.600 528.800 24.400 529.000 ;
        RECT 3.800 527.600 4.400 528.000 ;
        RECT 7.400 527.600 13.200 528.200 ;
        RECT 13.800 527.600 16.400 528.400 ;
        RECT 1.200 526.800 3.200 527.400 ;
        RECT 3.800 526.800 8.000 527.600 ;
        RECT 2.600 526.200 3.200 526.800 ;
        RECT 2.600 525.600 3.600 526.200 ;
        RECT 2.800 522.200 3.600 525.600 ;
        RECT 6.000 522.200 6.800 526.800 ;
        RECT 9.200 522.200 10.000 525.000 ;
        RECT 10.800 522.200 11.600 525.000 ;
        RECT 12.400 522.200 13.200 527.000 ;
        RECT 15.600 522.200 16.400 527.000 ;
        RECT 18.800 522.200 19.600 528.400 ;
        RECT 26.800 527.600 29.400 528.400 ;
        RECT 22.000 526.800 26.200 527.600 ;
        RECT 20.400 522.200 21.200 525.000 ;
        RECT 22.000 522.200 22.800 525.000 ;
        RECT 23.600 522.200 24.400 525.000 ;
        RECT 26.800 522.200 27.600 527.600 ;
        RECT 32.000 527.400 32.600 529.000 ;
        RECT 30.000 526.800 32.600 527.400 ;
        RECT 33.200 530.000 34.200 530.800 ;
        RECT 34.800 530.300 35.600 530.400 ;
        RECT 36.400 530.300 37.200 530.400 ;
        RECT 34.800 530.200 37.200 530.300 ;
        RECT 38.400 530.200 39.000 533.600 ;
        RECT 39.600 531.600 40.400 533.200 ;
        RECT 30.000 522.200 30.800 526.800 ;
        RECT 33.200 522.200 34.000 530.000 ;
        RECT 34.800 529.700 37.800 530.200 ;
        RECT 34.800 529.600 35.600 529.700 ;
        RECT 36.400 529.600 37.800 529.700 ;
        RECT 38.400 529.600 39.400 530.200 ;
        RECT 37.200 528.400 37.800 529.600 ;
        RECT 37.200 527.600 38.000 528.400 ;
        RECT 38.600 522.200 39.400 529.600 ;
        RECT 42.800 528.800 43.600 530.400 ;
        RECT 44.400 522.200 45.200 535.600 ;
        RECT 46.000 533.600 46.800 535.200 ;
        RECT 49.200 534.300 50.000 539.800 ;
        RECT 50.800 536.000 51.600 539.800 ;
        RECT 54.000 536.000 54.800 539.800 ;
        RECT 50.800 535.800 54.800 536.000 ;
        RECT 55.600 535.800 56.400 539.800 ;
        RECT 57.200 536.000 58.000 539.800 ;
        RECT 60.400 536.000 61.200 539.800 ;
        RECT 57.200 535.800 61.200 536.000 ;
        RECT 62.000 535.800 62.800 539.800 ;
        RECT 65.200 536.000 66.000 539.800 ;
        RECT 51.000 535.400 54.600 535.800 ;
        RECT 51.600 534.400 52.400 534.800 ;
        RECT 55.600 534.400 56.200 535.800 ;
        RECT 57.400 535.400 61.000 535.800 ;
        RECT 58.000 534.400 58.800 534.800 ;
        RECT 62.000 534.400 62.600 535.800 ;
        RECT 65.000 535.200 66.000 536.000 ;
        RECT 50.800 534.300 52.400 534.400 ;
        RECT 49.200 533.800 52.400 534.300 ;
        RECT 49.200 533.700 51.600 533.800 ;
        RECT 49.200 522.200 50.000 533.700 ;
        RECT 50.800 533.600 51.600 533.700 ;
        RECT 53.800 533.600 56.400 534.400 ;
        RECT 57.200 533.800 58.800 534.400 ;
        RECT 57.200 533.600 58.000 533.800 ;
        RECT 60.200 533.600 62.800 534.400 ;
        RECT 52.400 531.600 53.200 533.200 ;
        RECT 53.800 530.200 54.400 533.600 ;
        RECT 58.800 531.600 59.600 533.200 ;
        RECT 60.200 530.400 60.800 533.600 ;
        RECT 65.000 530.800 65.800 535.200 ;
        RECT 66.800 534.600 67.600 539.800 ;
        RECT 73.200 536.600 74.000 539.800 ;
        RECT 74.800 537.000 75.600 539.800 ;
        RECT 76.400 537.000 77.200 539.800 ;
        RECT 78.000 537.000 78.800 539.800 ;
        RECT 79.600 537.000 80.400 539.800 ;
        RECT 82.800 537.000 83.600 539.800 ;
        RECT 86.000 537.000 86.800 539.800 ;
        RECT 87.600 537.000 88.400 539.800 ;
        RECT 89.200 537.000 90.000 539.800 ;
        RECT 71.600 535.800 74.000 536.600 ;
        RECT 90.800 536.600 91.600 539.800 ;
        RECT 71.600 535.200 72.400 535.800 ;
        RECT 66.400 534.000 67.600 534.600 ;
        RECT 70.600 534.600 72.400 535.200 ;
        RECT 76.400 535.600 77.400 536.400 ;
        RECT 80.400 535.600 82.000 536.400 ;
        RECT 82.800 535.800 87.400 536.400 ;
        RECT 90.800 535.800 93.400 536.600 ;
        RECT 82.800 535.600 83.600 535.800 ;
        RECT 66.400 532.000 67.000 534.000 ;
        RECT 70.600 533.400 71.400 534.600 ;
        RECT 67.600 532.600 71.400 533.400 ;
        RECT 76.400 532.800 77.200 535.600 ;
        RECT 82.800 534.800 83.600 535.000 ;
        RECT 79.200 534.200 83.600 534.800 ;
        RECT 79.200 534.000 80.000 534.200 ;
        RECT 84.400 533.600 85.200 535.200 ;
        RECT 86.600 533.400 87.400 535.800 ;
        RECT 92.600 535.200 93.400 535.800 ;
        RECT 92.600 534.400 95.600 535.200 ;
        RECT 97.200 533.800 98.000 539.800 ;
        RECT 98.800 536.000 99.600 539.800 ;
        RECT 102.000 536.000 102.800 539.800 ;
        RECT 98.800 535.800 102.800 536.000 ;
        RECT 103.600 535.800 104.400 539.800 ;
        RECT 105.200 536.000 106.000 539.800 ;
        RECT 108.400 536.000 109.200 539.800 ;
        RECT 105.200 535.800 109.200 536.000 ;
        RECT 110.000 535.800 110.800 539.800 ;
        RECT 111.600 536.000 112.400 539.800 ;
        RECT 114.800 536.000 115.600 539.800 ;
        RECT 111.600 535.800 115.600 536.000 ;
        RECT 116.400 535.800 117.200 539.800 ;
        RECT 118.000 535.800 118.800 539.800 ;
        RECT 119.600 536.000 120.400 539.800 ;
        RECT 122.800 536.000 123.600 539.800 ;
        RECT 119.600 535.800 123.600 536.000 ;
        RECT 124.400 535.800 125.200 539.800 ;
        RECT 128.800 536.200 130.400 539.800 ;
        RECT 99.000 535.400 102.600 535.800 ;
        RECT 99.600 534.400 100.400 534.800 ;
        RECT 103.600 534.400 104.200 535.800 ;
        RECT 105.400 535.400 109.000 535.800 ;
        RECT 106.000 534.400 106.800 534.800 ;
        RECT 110.000 534.400 110.600 535.800 ;
        RECT 111.800 535.400 115.400 535.800 ;
        RECT 112.400 534.400 113.200 534.800 ;
        RECT 116.400 534.400 117.000 535.800 ;
        RECT 118.200 534.400 118.800 535.800 ;
        RECT 119.800 535.400 123.400 535.800 ;
        RECT 124.400 535.200 126.600 535.800 ;
        RECT 127.600 535.400 129.200 535.600 ;
        RECT 125.800 535.000 126.600 535.200 ;
        RECT 127.200 534.800 129.200 535.400 ;
        RECT 122.000 534.400 122.800 534.800 ;
        RECT 127.200 534.400 127.800 534.800 ;
        RECT 79.600 532.600 82.800 533.400 ;
        RECT 86.600 532.600 88.600 533.400 ;
        RECT 89.200 533.000 98.000 533.800 ;
        RECT 98.800 533.800 100.400 534.400 ;
        RECT 98.800 533.600 99.600 533.800 ;
        RECT 101.800 533.600 104.400 534.400 ;
        RECT 105.200 533.800 106.800 534.400 ;
        RECT 105.200 533.600 106.000 533.800 ;
        RECT 108.200 533.600 110.800 534.400 ;
        RECT 111.600 533.800 113.200 534.400 ;
        RECT 111.600 533.600 112.400 533.800 ;
        RECT 114.600 533.600 117.200 534.400 ;
        RECT 118.000 533.600 120.600 534.400 ;
        RECT 122.000 534.300 123.600 534.400 ;
        RECT 124.400 534.300 127.800 534.400 ;
        RECT 122.000 533.800 127.800 534.300 ;
        RECT 122.800 533.700 126.000 533.800 ;
        RECT 122.800 533.600 123.600 533.700 ;
        RECT 124.400 533.600 126.000 533.700 ;
        RECT 73.200 532.000 74.000 532.600 ;
        RECT 90.800 532.000 91.600 532.400 ;
        RECT 94.000 532.000 94.800 532.400 ;
        RECT 95.800 532.000 96.600 532.200 ;
        RECT 66.400 531.400 67.200 532.000 ;
        RECT 73.200 531.400 96.600 532.000 ;
        RECT 55.600 530.200 56.400 530.400 ;
        RECT 53.400 529.600 54.400 530.200 ;
        RECT 55.000 529.600 56.400 530.200 ;
        RECT 58.800 529.600 60.800 530.400 ;
        RECT 62.000 530.300 62.800 530.400 ;
        RECT 65.000 530.300 66.000 530.800 ;
        RECT 62.000 530.200 66.000 530.300 ;
        RECT 61.400 529.700 66.000 530.200 ;
        RECT 61.400 529.600 62.800 529.700 ;
        RECT 53.400 522.200 54.200 529.600 ;
        RECT 55.000 528.400 55.600 529.600 ;
        RECT 54.800 527.600 55.600 528.400 ;
        RECT 59.800 522.200 60.600 529.600 ;
        RECT 61.400 528.400 62.000 529.600 ;
        RECT 61.200 527.600 62.000 528.400 ;
        RECT 65.200 522.200 66.000 529.700 ;
        RECT 66.600 529.600 67.200 531.400 ;
        RECT 66.600 529.000 75.600 529.600 ;
        RECT 66.600 527.400 67.200 529.000 ;
        RECT 74.800 528.800 75.600 529.000 ;
        RECT 78.000 529.000 86.600 529.600 ;
        RECT 78.000 528.800 78.800 529.000 ;
        RECT 69.800 527.600 72.400 528.400 ;
        RECT 66.600 526.800 69.200 527.400 ;
        RECT 68.400 522.200 69.200 526.800 ;
        RECT 71.600 522.200 72.400 527.600 ;
        RECT 73.000 526.800 77.200 527.600 ;
        RECT 74.800 522.200 75.600 525.000 ;
        RECT 76.400 522.200 77.200 525.000 ;
        RECT 78.000 522.200 78.800 525.000 ;
        RECT 79.600 522.200 80.400 528.400 ;
        RECT 82.800 527.600 85.400 528.400 ;
        RECT 86.000 528.200 86.600 529.000 ;
        RECT 87.600 529.400 88.400 529.600 ;
        RECT 87.600 529.000 93.000 529.400 ;
        RECT 87.600 528.800 93.800 529.000 ;
        RECT 92.400 528.200 93.800 528.800 ;
        RECT 86.000 527.600 91.800 528.200 ;
        RECT 94.800 528.000 96.400 528.800 ;
        RECT 94.800 527.600 95.400 528.000 ;
        RECT 82.800 522.200 83.600 527.000 ;
        RECT 86.000 522.200 86.800 527.000 ;
        RECT 91.200 526.800 95.400 527.600 ;
        RECT 97.200 527.400 98.000 533.000 ;
        RECT 100.400 531.600 101.200 533.200 ;
        RECT 101.800 530.200 102.400 533.600 ;
        RECT 105.200 532.300 106.000 532.400 ;
        RECT 106.800 532.300 107.600 533.200 ;
        RECT 105.200 531.700 107.600 532.300 ;
        RECT 105.200 531.600 106.000 531.700 ;
        RECT 106.800 531.600 107.600 531.700 ;
        RECT 103.600 530.200 104.400 530.400 ;
        RECT 108.200 530.200 108.800 533.600 ;
        RECT 113.200 531.600 114.000 533.200 ;
        RECT 114.600 532.300 115.200 533.600 ;
        RECT 114.600 531.700 118.700 532.300 ;
        RECT 110.000 530.200 110.800 530.400 ;
        RECT 114.600 530.200 115.200 531.700 ;
        RECT 118.100 530.400 118.700 531.700 ;
        RECT 116.400 530.200 117.200 530.400 ;
        RECT 96.000 526.800 98.000 527.400 ;
        RECT 101.400 529.600 102.400 530.200 ;
        RECT 103.000 529.600 104.400 530.200 ;
        RECT 107.800 529.600 108.800 530.200 ;
        RECT 109.400 529.600 110.800 530.200 ;
        RECT 114.200 529.600 115.200 530.200 ;
        RECT 115.800 529.600 117.200 530.200 ;
        RECT 118.000 530.200 118.800 530.400 ;
        RECT 120.000 530.200 120.600 533.600 ;
        RECT 128.400 533.400 129.200 534.200 ;
        RECT 121.200 532.300 122.000 533.200 ;
        RECT 128.400 532.800 129.000 533.400 ;
        RECT 122.800 532.300 123.600 532.400 ;
        RECT 121.200 531.700 123.600 532.300 ;
        RECT 126.400 532.200 129.000 532.800 ;
        RECT 129.800 532.800 130.400 536.200 ;
        RECT 134.000 535.800 134.800 539.800 ;
        RECT 142.000 536.000 142.800 539.800 ;
        RECT 131.000 534.800 131.800 535.600 ;
        RECT 132.400 535.200 134.800 535.800 ;
        RECT 141.800 535.200 142.800 536.000 ;
        RECT 132.400 535.000 133.200 535.200 ;
        RECT 131.200 534.400 131.800 534.800 ;
        RECT 131.200 533.600 132.000 534.400 ;
        RECT 133.200 534.300 134.800 534.400 ;
        RECT 141.800 534.300 142.600 535.200 ;
        RECT 143.600 534.600 144.400 539.800 ;
        RECT 150.000 536.600 150.800 539.800 ;
        RECT 151.600 537.000 152.400 539.800 ;
        RECT 153.200 537.000 154.000 539.800 ;
        RECT 154.800 537.000 155.600 539.800 ;
        RECT 156.400 537.000 157.200 539.800 ;
        RECT 159.600 537.000 160.400 539.800 ;
        RECT 162.800 537.000 163.600 539.800 ;
        RECT 164.400 537.000 165.200 539.800 ;
        RECT 166.000 537.000 166.800 539.800 ;
        RECT 148.400 535.800 150.800 536.600 ;
        RECT 167.600 536.600 168.400 539.800 ;
        RECT 148.400 535.200 149.200 535.800 ;
        RECT 133.200 533.700 142.600 534.300 ;
        RECT 133.200 533.600 134.800 533.700 ;
        RECT 129.800 532.400 130.800 532.800 ;
        RECT 129.800 532.300 131.600 532.400 ;
        RECT 140.400 532.300 141.200 532.400 ;
        RECT 129.800 532.200 141.200 532.300 ;
        RECT 126.400 532.000 127.200 532.200 ;
        RECT 121.200 531.600 122.000 531.700 ;
        RECT 122.800 531.600 123.600 531.700 ;
        RECT 130.200 531.700 141.200 532.200 ;
        RECT 130.200 531.600 131.600 531.700 ;
        RECT 140.400 531.600 141.200 531.700 ;
        RECT 128.600 531.400 129.400 531.600 ;
        RECT 126.000 530.800 129.400 531.400 ;
        RECT 126.000 530.200 126.600 530.800 ;
        RECT 130.200 530.200 130.800 531.600 ;
        RECT 141.800 530.800 142.600 533.700 ;
        RECT 143.200 534.000 144.400 534.600 ;
        RECT 147.400 534.600 149.200 535.200 ;
        RECT 153.200 535.600 154.200 536.400 ;
        RECT 157.200 535.600 158.800 536.400 ;
        RECT 159.600 535.800 164.200 536.400 ;
        RECT 167.600 535.800 170.200 536.600 ;
        RECT 159.600 535.600 160.400 535.800 ;
        RECT 143.200 532.000 143.800 534.000 ;
        RECT 147.400 533.400 148.200 534.600 ;
        RECT 144.400 532.600 148.200 533.400 ;
        RECT 153.200 532.800 154.000 535.600 ;
        RECT 159.600 534.800 160.400 535.000 ;
        RECT 156.000 534.200 160.400 534.800 ;
        RECT 156.000 534.000 156.800 534.200 ;
        RECT 161.200 533.600 162.000 535.200 ;
        RECT 163.400 533.400 164.200 535.800 ;
        RECT 169.400 535.200 170.200 535.800 ;
        RECT 169.400 534.400 172.400 535.200 ;
        RECT 174.000 533.800 174.800 539.800 ;
        RECT 156.400 532.600 159.600 533.400 ;
        RECT 163.400 532.600 165.400 533.400 ;
        RECT 166.000 533.000 174.800 533.800 ;
        RECT 150.000 532.000 150.800 532.600 ;
        RECT 167.600 532.000 168.400 532.400 ;
        RECT 172.600 532.000 173.400 532.200 ;
        RECT 143.200 531.400 144.000 532.000 ;
        RECT 150.000 531.400 173.400 532.000 ;
        RECT 118.000 529.600 119.400 530.200 ;
        RECT 120.000 529.600 121.000 530.200 ;
        RECT 87.600 522.200 88.400 525.000 ;
        RECT 89.200 522.200 90.000 525.000 ;
        RECT 92.400 522.200 93.200 526.800 ;
        RECT 96.000 526.200 96.600 526.800 ;
        RECT 95.600 525.600 96.600 526.200 ;
        RECT 95.600 522.200 96.400 525.600 ;
        RECT 101.400 522.200 102.200 529.600 ;
        RECT 103.000 528.400 103.600 529.600 ;
        RECT 102.800 527.600 103.600 528.400 ;
        RECT 107.800 522.200 108.600 529.600 ;
        RECT 109.400 528.400 110.000 529.600 ;
        RECT 109.200 527.600 110.000 528.400 ;
        RECT 114.200 522.200 115.000 529.600 ;
        RECT 115.800 528.400 116.400 529.600 ;
        RECT 115.600 527.600 116.400 528.400 ;
        RECT 118.800 528.400 119.400 529.600 ;
        RECT 118.800 527.600 119.600 528.400 ;
        RECT 120.200 522.200 121.000 529.600 ;
        RECT 124.400 529.600 126.600 530.200 ;
        RECT 124.400 522.200 125.200 529.600 ;
        RECT 125.800 529.400 126.600 529.600 ;
        RECT 128.800 529.600 130.800 530.200 ;
        RECT 132.400 529.600 134.800 530.200 ;
        RECT 141.800 530.000 142.800 530.800 ;
        RECT 128.800 522.200 130.400 529.600 ;
        RECT 132.400 529.400 133.200 529.600 ;
        RECT 134.000 522.200 134.800 529.600 ;
        RECT 142.000 522.200 142.800 530.000 ;
        RECT 143.400 529.600 144.000 531.400 ;
        RECT 143.400 529.000 152.400 529.600 ;
        RECT 143.400 527.400 144.000 529.000 ;
        RECT 151.600 528.800 152.400 529.000 ;
        RECT 154.800 529.000 163.400 529.600 ;
        RECT 154.800 528.800 155.600 529.000 ;
        RECT 146.600 527.600 149.200 528.400 ;
        RECT 143.400 526.800 146.000 527.400 ;
        RECT 145.200 522.200 146.000 526.800 ;
        RECT 148.400 522.200 149.200 527.600 ;
        RECT 149.800 526.800 154.000 527.600 ;
        RECT 151.600 522.200 152.400 525.000 ;
        RECT 153.200 522.200 154.000 525.000 ;
        RECT 154.800 522.200 155.600 525.000 ;
        RECT 156.400 522.200 157.200 528.400 ;
        RECT 159.600 527.600 162.200 528.400 ;
        RECT 162.800 528.200 163.400 529.000 ;
        RECT 164.400 529.400 165.200 529.600 ;
        RECT 164.400 529.000 169.800 529.400 ;
        RECT 164.400 528.800 170.600 529.000 ;
        RECT 169.200 528.200 170.600 528.800 ;
        RECT 162.800 527.600 168.600 528.200 ;
        RECT 171.600 528.000 173.200 528.800 ;
        RECT 171.600 527.600 172.200 528.000 ;
        RECT 159.600 522.200 160.400 527.000 ;
        RECT 162.800 522.200 163.600 527.000 ;
        RECT 168.000 526.800 172.200 527.600 ;
        RECT 174.000 527.400 174.800 533.000 ;
        RECT 172.800 526.800 174.800 527.400 ;
        RECT 175.600 533.800 176.400 539.800 ;
        RECT 182.000 536.600 182.800 539.800 ;
        RECT 183.600 537.000 184.400 539.800 ;
        RECT 185.200 537.000 186.000 539.800 ;
        RECT 186.800 537.000 187.600 539.800 ;
        RECT 190.000 537.000 190.800 539.800 ;
        RECT 193.200 537.000 194.000 539.800 ;
        RECT 194.800 537.000 195.600 539.800 ;
        RECT 196.400 537.000 197.200 539.800 ;
        RECT 198.000 537.000 198.800 539.800 ;
        RECT 180.200 535.800 182.800 536.600 ;
        RECT 199.600 536.600 200.400 539.800 ;
        RECT 186.200 535.800 190.800 536.400 ;
        RECT 180.200 535.200 181.000 535.800 ;
        RECT 178.000 534.400 181.000 535.200 ;
        RECT 175.600 533.000 184.400 533.800 ;
        RECT 186.200 533.400 187.000 535.800 ;
        RECT 190.000 535.600 190.800 535.800 ;
        RECT 191.600 535.600 193.200 536.400 ;
        RECT 196.200 535.600 197.200 536.400 ;
        RECT 199.600 535.800 202.000 536.600 ;
        RECT 188.400 533.600 189.200 535.200 ;
        RECT 190.000 534.800 190.800 535.000 ;
        RECT 190.000 534.200 194.400 534.800 ;
        RECT 193.600 534.000 194.400 534.200 ;
        RECT 175.600 527.400 176.400 533.000 ;
        RECT 185.000 532.600 187.000 533.400 ;
        RECT 190.800 532.600 194.000 533.400 ;
        RECT 196.400 532.800 197.200 535.600 ;
        RECT 201.200 535.200 202.000 535.800 ;
        RECT 201.200 534.600 203.000 535.200 ;
        RECT 202.200 533.400 203.000 534.600 ;
        RECT 206.000 534.600 206.800 539.800 ;
        RECT 207.600 536.300 208.400 539.800 ;
        RECT 210.800 536.300 211.600 537.200 ;
        RECT 207.600 535.700 211.600 536.300 ;
        RECT 207.600 535.200 208.600 535.700 ;
        RECT 210.800 535.600 211.600 535.700 ;
        RECT 206.000 534.000 207.200 534.600 ;
        RECT 202.200 532.600 206.000 533.400 ;
        RECT 177.200 532.200 178.000 532.400 ;
        RECT 177.000 532.000 178.000 532.200 ;
        RECT 182.000 532.000 182.800 532.400 ;
        RECT 199.600 532.000 200.400 532.600 ;
        RECT 206.600 532.000 207.200 534.000 ;
        RECT 177.000 531.400 200.400 532.000 ;
        RECT 206.400 531.400 207.200 532.000 ;
        RECT 206.400 529.600 207.000 531.400 ;
        RECT 207.800 530.800 208.600 535.200 ;
        RECT 185.200 529.400 186.000 529.600 ;
        RECT 180.600 529.000 186.000 529.400 ;
        RECT 179.800 528.800 186.000 529.000 ;
        RECT 187.000 529.000 195.600 529.600 ;
        RECT 177.200 528.000 178.800 528.800 ;
        RECT 179.800 528.200 181.200 528.800 ;
        RECT 187.000 528.200 187.600 529.000 ;
        RECT 194.800 528.800 195.600 529.000 ;
        RECT 198.000 529.000 207.000 529.600 ;
        RECT 198.000 528.800 198.800 529.000 ;
        RECT 178.200 527.600 178.800 528.000 ;
        RECT 181.800 527.600 187.600 528.200 ;
        RECT 188.200 527.600 190.800 528.400 ;
        RECT 175.600 526.800 177.600 527.400 ;
        RECT 178.200 526.800 182.400 527.600 ;
        RECT 164.400 522.200 165.200 525.000 ;
        RECT 166.000 522.200 166.800 525.000 ;
        RECT 169.200 522.200 170.000 526.800 ;
        RECT 172.800 526.200 173.400 526.800 ;
        RECT 172.400 525.600 173.400 526.200 ;
        RECT 177.000 526.200 177.600 526.800 ;
        RECT 177.000 525.600 178.000 526.200 ;
        RECT 172.400 522.200 173.200 525.600 ;
        RECT 177.200 522.200 178.000 525.600 ;
        RECT 180.400 522.200 181.200 526.800 ;
        RECT 183.600 522.200 184.400 525.000 ;
        RECT 185.200 522.200 186.000 525.000 ;
        RECT 186.800 522.200 187.600 527.000 ;
        RECT 190.000 522.200 190.800 527.000 ;
        RECT 193.200 522.200 194.000 528.400 ;
        RECT 201.200 527.600 203.800 528.400 ;
        RECT 196.400 526.800 200.600 527.600 ;
        RECT 194.800 522.200 195.600 525.000 ;
        RECT 196.400 522.200 197.200 525.000 ;
        RECT 198.000 522.200 198.800 525.000 ;
        RECT 201.200 522.200 202.000 527.600 ;
        RECT 206.400 527.400 207.000 529.000 ;
        RECT 204.400 526.800 207.000 527.400 ;
        RECT 207.600 530.000 208.600 530.800 ;
        RECT 212.400 532.300 213.200 539.800 ;
        RECT 214.000 536.000 214.800 539.800 ;
        RECT 217.200 536.000 218.000 539.800 ;
        RECT 214.000 535.800 218.000 536.000 ;
        RECT 218.800 535.800 219.600 539.800 ;
        RECT 221.000 536.400 221.800 539.800 ;
        RECT 221.000 535.800 222.800 536.400 ;
        RECT 226.800 536.000 227.600 539.800 ;
        RECT 214.200 535.400 217.800 535.800 ;
        RECT 214.800 534.400 215.600 534.800 ;
        RECT 218.800 534.400 219.400 535.800 ;
        RECT 214.000 533.800 215.600 534.400 ;
        RECT 214.000 533.600 214.800 533.800 ;
        RECT 217.000 533.600 219.600 534.400 ;
        RECT 215.600 532.300 216.400 533.200 ;
        RECT 212.400 531.700 216.400 532.300 ;
        RECT 204.400 522.200 205.200 526.800 ;
        RECT 207.600 522.200 208.400 530.000 ;
        RECT 212.400 522.200 213.200 531.700 ;
        RECT 215.600 531.600 216.400 531.700 ;
        RECT 217.000 530.200 217.600 533.600 ;
        RECT 222.000 532.300 222.800 535.800 ;
        RECT 226.600 535.200 227.600 536.000 ;
        RECT 223.600 534.300 224.400 535.200 ;
        RECT 225.200 534.300 226.000 534.400 ;
        RECT 223.600 533.700 226.000 534.300 ;
        RECT 223.600 533.600 224.400 533.700 ;
        RECT 225.200 533.600 226.000 533.700 ;
        RECT 218.900 531.700 222.800 532.300 ;
        RECT 218.900 530.400 219.500 531.700 ;
        RECT 218.800 530.200 219.600 530.400 ;
        RECT 216.600 529.600 217.600 530.200 ;
        RECT 218.200 529.600 219.600 530.200 ;
        RECT 216.600 522.200 217.400 529.600 ;
        RECT 218.200 528.400 218.800 529.600 ;
        RECT 220.400 528.800 221.200 530.400 ;
        RECT 218.000 527.600 218.800 528.400 ;
        RECT 222.000 522.200 222.800 531.700 ;
        RECT 226.600 530.800 227.400 535.200 ;
        RECT 228.400 534.600 229.200 539.800 ;
        RECT 234.800 536.600 235.600 539.800 ;
        RECT 236.400 537.000 237.200 539.800 ;
        RECT 238.000 537.000 238.800 539.800 ;
        RECT 239.600 537.000 240.400 539.800 ;
        RECT 241.200 537.000 242.000 539.800 ;
        RECT 244.400 537.000 245.200 539.800 ;
        RECT 247.600 537.000 248.400 539.800 ;
        RECT 249.200 537.000 250.000 539.800 ;
        RECT 250.800 537.000 251.600 539.800 ;
        RECT 233.200 535.800 235.600 536.600 ;
        RECT 252.400 536.600 253.200 539.800 ;
        RECT 233.200 535.200 234.000 535.800 ;
        RECT 228.000 534.000 229.200 534.600 ;
        RECT 232.200 534.600 234.000 535.200 ;
        RECT 238.000 535.600 239.000 536.400 ;
        RECT 242.000 535.600 243.600 536.400 ;
        RECT 244.400 535.800 249.000 536.400 ;
        RECT 252.400 535.800 255.000 536.600 ;
        RECT 244.400 535.600 245.200 535.800 ;
        RECT 228.000 532.000 228.600 534.000 ;
        RECT 232.200 533.400 233.000 534.600 ;
        RECT 229.200 532.600 233.000 533.400 ;
        RECT 238.000 532.800 238.800 535.600 ;
        RECT 244.400 534.800 245.200 535.000 ;
        RECT 240.800 534.200 245.200 534.800 ;
        RECT 240.800 534.000 241.600 534.200 ;
        RECT 246.000 533.600 246.800 535.200 ;
        RECT 248.200 533.400 249.000 535.800 ;
        RECT 254.200 535.200 255.000 535.800 ;
        RECT 254.200 534.400 257.200 535.200 ;
        RECT 258.800 533.800 259.600 539.800 ;
        RECT 241.200 532.600 244.400 533.400 ;
        RECT 248.200 532.600 250.200 533.400 ;
        RECT 250.800 533.000 259.600 533.800 ;
        RECT 234.800 532.000 235.600 532.600 ;
        RECT 252.400 532.000 253.200 532.400 ;
        RECT 257.400 532.000 258.200 532.200 ;
        RECT 228.000 531.400 228.800 532.000 ;
        RECT 234.800 531.400 258.200 532.000 ;
        RECT 226.600 530.000 227.600 530.800 ;
        RECT 226.800 522.200 227.600 530.000 ;
        RECT 228.200 529.600 228.800 531.400 ;
        RECT 228.200 529.000 237.200 529.600 ;
        RECT 228.200 527.400 228.800 529.000 ;
        RECT 236.400 528.800 237.200 529.000 ;
        RECT 239.600 529.000 248.200 529.600 ;
        RECT 239.600 528.800 240.400 529.000 ;
        RECT 231.400 527.600 234.000 528.400 ;
        RECT 228.200 526.800 230.800 527.400 ;
        RECT 230.000 522.200 230.800 526.800 ;
        RECT 233.200 522.200 234.000 527.600 ;
        RECT 234.600 526.800 238.800 527.600 ;
        RECT 236.400 522.200 237.200 525.000 ;
        RECT 238.000 522.200 238.800 525.000 ;
        RECT 239.600 522.200 240.400 525.000 ;
        RECT 241.200 522.200 242.000 528.400 ;
        RECT 244.400 527.600 247.000 528.400 ;
        RECT 247.600 528.200 248.200 529.000 ;
        RECT 249.200 529.400 250.000 529.600 ;
        RECT 249.200 529.000 254.600 529.400 ;
        RECT 249.200 528.800 255.400 529.000 ;
        RECT 254.000 528.200 255.400 528.800 ;
        RECT 247.600 527.600 253.400 528.200 ;
        RECT 256.400 528.000 258.000 528.800 ;
        RECT 256.400 527.600 257.000 528.000 ;
        RECT 244.400 522.200 245.200 527.000 ;
        RECT 247.600 522.200 248.400 527.000 ;
        RECT 252.800 526.800 257.000 527.600 ;
        RECT 258.800 527.400 259.600 533.000 ;
        RECT 257.600 526.800 259.600 527.400 ;
        RECT 260.400 533.800 261.200 539.800 ;
        RECT 266.800 536.600 267.600 539.800 ;
        RECT 268.400 537.000 269.200 539.800 ;
        RECT 270.000 537.000 270.800 539.800 ;
        RECT 271.600 537.000 272.400 539.800 ;
        RECT 274.800 537.000 275.600 539.800 ;
        RECT 278.000 537.000 278.800 539.800 ;
        RECT 279.600 537.000 280.400 539.800 ;
        RECT 281.200 537.000 282.000 539.800 ;
        RECT 282.800 537.000 283.600 539.800 ;
        RECT 265.000 535.800 267.600 536.600 ;
        RECT 284.400 536.600 285.200 539.800 ;
        RECT 271.000 535.800 275.600 536.400 ;
        RECT 265.000 535.200 265.800 535.800 ;
        RECT 262.800 534.400 265.800 535.200 ;
        RECT 260.400 533.000 269.200 533.800 ;
        RECT 271.000 533.400 271.800 535.800 ;
        RECT 274.800 535.600 275.600 535.800 ;
        RECT 276.400 535.600 278.000 536.400 ;
        RECT 281.000 535.600 282.000 536.400 ;
        RECT 284.400 535.800 286.800 536.600 ;
        RECT 273.200 533.600 274.000 535.200 ;
        RECT 274.800 534.800 275.600 535.000 ;
        RECT 274.800 534.200 279.200 534.800 ;
        RECT 278.400 534.000 279.200 534.200 ;
        RECT 260.400 527.400 261.200 533.000 ;
        RECT 269.800 532.600 271.800 533.400 ;
        RECT 275.600 532.600 278.800 533.400 ;
        RECT 281.200 532.800 282.000 535.600 ;
        RECT 286.000 535.200 286.800 535.800 ;
        RECT 286.000 534.600 287.800 535.200 ;
        RECT 287.000 533.400 287.800 534.600 ;
        RECT 290.800 534.600 291.600 539.800 ;
        RECT 292.400 536.000 293.200 539.800 ;
        RECT 292.400 535.200 293.400 536.000 ;
        RECT 295.600 535.600 296.400 537.200 ;
        RECT 290.800 534.000 292.000 534.600 ;
        RECT 287.000 532.600 290.800 533.400 ;
        RECT 261.800 532.000 262.600 532.200 ;
        RECT 263.600 532.000 264.400 532.400 ;
        RECT 266.800 532.000 267.600 532.400 ;
        RECT 284.400 532.000 285.200 532.600 ;
        RECT 291.400 532.000 292.000 534.000 ;
        RECT 261.800 531.400 285.200 532.000 ;
        RECT 291.200 531.400 292.000 532.000 ;
        RECT 291.200 529.600 291.800 531.400 ;
        RECT 292.600 530.800 293.400 535.200 ;
        RECT 270.000 529.400 270.800 529.600 ;
        RECT 265.400 529.000 270.800 529.400 ;
        RECT 264.600 528.800 270.800 529.000 ;
        RECT 271.800 529.000 280.400 529.600 ;
        RECT 262.000 528.000 263.600 528.800 ;
        RECT 264.600 528.200 266.000 528.800 ;
        RECT 271.800 528.200 272.400 529.000 ;
        RECT 279.600 528.800 280.400 529.000 ;
        RECT 282.800 529.000 291.800 529.600 ;
        RECT 282.800 528.800 283.600 529.000 ;
        RECT 263.000 527.600 263.600 528.000 ;
        RECT 266.600 527.600 272.400 528.200 ;
        RECT 273.000 527.600 275.600 528.400 ;
        RECT 260.400 526.800 262.400 527.400 ;
        RECT 263.000 526.800 267.200 527.600 ;
        RECT 249.200 522.200 250.000 525.000 ;
        RECT 250.800 522.200 251.600 525.000 ;
        RECT 254.000 522.200 254.800 526.800 ;
        RECT 257.600 526.200 258.200 526.800 ;
        RECT 257.200 525.600 258.200 526.200 ;
        RECT 261.800 526.200 262.400 526.800 ;
        RECT 261.800 525.600 262.800 526.200 ;
        RECT 257.200 522.200 258.000 525.600 ;
        RECT 262.000 522.200 262.800 525.600 ;
        RECT 265.200 522.200 266.000 526.800 ;
        RECT 268.400 522.200 269.200 525.000 ;
        RECT 270.000 522.200 270.800 525.000 ;
        RECT 271.600 522.200 272.400 527.000 ;
        RECT 274.800 522.200 275.600 527.000 ;
        RECT 278.000 522.200 278.800 528.400 ;
        RECT 286.000 527.600 288.600 528.400 ;
        RECT 281.200 526.800 285.400 527.600 ;
        RECT 279.600 522.200 280.400 525.000 ;
        RECT 281.200 522.200 282.000 525.000 ;
        RECT 282.800 522.200 283.600 525.000 ;
        RECT 286.000 522.200 286.800 527.600 ;
        RECT 291.200 527.400 291.800 529.000 ;
        RECT 289.200 526.800 291.800 527.400 ;
        RECT 292.400 530.000 293.400 530.800 ;
        RECT 297.200 532.300 298.000 539.800 ;
        RECT 298.800 536.000 299.600 539.800 ;
        RECT 302.000 536.000 302.800 539.800 ;
        RECT 298.800 535.800 302.800 536.000 ;
        RECT 303.600 535.800 304.400 539.800 ;
        RECT 312.600 536.400 313.400 539.800 ;
        RECT 311.600 535.800 313.400 536.400 ;
        RECT 316.400 536.000 317.200 539.800 ;
        RECT 299.000 535.400 302.600 535.800 ;
        RECT 299.600 534.400 300.400 534.800 ;
        RECT 303.600 534.400 304.200 535.800 ;
        RECT 298.800 533.800 300.400 534.400 ;
        RECT 298.800 533.600 299.600 533.800 ;
        RECT 301.800 533.600 304.400 534.400 ;
        RECT 310.000 533.600 310.800 535.200 ;
        RECT 300.400 532.300 301.200 533.200 ;
        RECT 297.200 531.700 301.200 532.300 ;
        RECT 289.200 522.200 290.000 526.800 ;
        RECT 292.400 522.200 293.200 530.000 ;
        RECT 297.200 522.200 298.000 531.700 ;
        RECT 300.400 531.600 301.200 531.700 ;
        RECT 301.800 530.200 302.400 533.600 ;
        RECT 303.600 530.300 304.400 530.400 ;
        RECT 311.600 530.300 312.400 535.800 ;
        RECT 316.200 535.200 317.200 536.000 ;
        RECT 316.200 530.800 317.000 535.200 ;
        RECT 318.000 534.600 318.800 539.800 ;
        RECT 324.400 536.600 325.200 539.800 ;
        RECT 326.000 537.000 326.800 539.800 ;
        RECT 327.600 537.000 328.400 539.800 ;
        RECT 329.200 537.000 330.000 539.800 ;
        RECT 330.800 537.000 331.600 539.800 ;
        RECT 334.000 537.000 334.800 539.800 ;
        RECT 337.200 537.000 338.000 539.800 ;
        RECT 338.800 537.000 339.600 539.800 ;
        RECT 340.400 537.000 341.200 539.800 ;
        RECT 322.800 535.800 325.200 536.600 ;
        RECT 342.000 536.600 342.800 539.800 ;
        RECT 322.800 535.200 323.600 535.800 ;
        RECT 317.600 534.000 318.800 534.600 ;
        RECT 321.800 534.600 323.600 535.200 ;
        RECT 327.600 535.600 328.600 536.400 ;
        RECT 331.600 535.600 333.200 536.400 ;
        RECT 334.000 535.800 338.600 536.400 ;
        RECT 342.000 535.800 344.600 536.600 ;
        RECT 334.000 535.600 334.800 535.800 ;
        RECT 317.600 532.000 318.200 534.000 ;
        RECT 321.800 533.400 322.600 534.600 ;
        RECT 318.800 532.600 322.600 533.400 ;
        RECT 327.600 532.800 328.400 535.600 ;
        RECT 334.000 534.800 334.800 535.000 ;
        RECT 330.400 534.200 334.800 534.800 ;
        RECT 330.400 534.000 331.200 534.200 ;
        RECT 335.600 533.600 336.400 535.200 ;
        RECT 337.800 533.400 338.600 535.800 ;
        RECT 343.800 535.200 344.600 535.800 ;
        RECT 343.800 534.400 346.800 535.200 ;
        RECT 348.400 533.800 349.200 539.800 ;
        RECT 350.000 535.600 350.800 539.800 ;
        RECT 351.600 536.000 352.400 539.800 ;
        RECT 354.800 536.000 355.600 539.800 ;
        RECT 351.600 535.800 355.600 536.000 ;
        RECT 350.200 534.400 350.800 535.600 ;
        RECT 351.800 535.400 355.400 535.800 ;
        RECT 354.000 534.400 354.800 534.800 ;
        RECT 330.800 532.600 334.000 533.400 ;
        RECT 337.800 532.600 339.800 533.400 ;
        RECT 340.400 533.000 349.200 533.800 ;
        RECT 350.000 533.600 352.600 534.400 ;
        RECT 354.000 534.300 355.600 534.400 ;
        RECT 356.400 534.300 357.200 539.800 ;
        RECT 359.600 535.800 360.400 539.800 ;
        RECT 361.200 536.000 362.000 539.800 ;
        RECT 364.400 536.000 365.200 539.800 ;
        RECT 361.200 535.800 365.200 536.000 ;
        RECT 366.000 536.000 366.800 539.800 ;
        RECT 369.200 536.000 370.000 539.800 ;
        RECT 366.000 535.800 370.000 536.000 ;
        RECT 370.800 535.800 371.600 539.800 ;
        RECT 359.800 534.400 360.400 535.800 ;
        RECT 361.400 535.400 365.000 535.800 ;
        RECT 366.200 535.400 369.800 535.800 ;
        RECT 363.600 534.400 364.400 534.800 ;
        RECT 366.800 534.400 367.600 534.800 ;
        RECT 370.800 534.400 371.400 535.800 ;
        RECT 354.000 533.800 357.200 534.300 ;
        RECT 354.800 533.700 357.200 533.800 ;
        RECT 354.800 533.600 355.600 533.700 ;
        RECT 324.400 532.000 325.200 532.600 ;
        RECT 342.000 532.000 342.800 532.400 ;
        RECT 345.200 532.000 346.000 532.400 ;
        RECT 347.000 532.000 347.800 532.200 ;
        RECT 317.600 531.400 318.400 532.000 ;
        RECT 324.400 531.400 347.800 532.000 ;
        RECT 303.600 530.200 312.400 530.300 ;
        RECT 301.400 529.600 302.400 530.200 ;
        RECT 303.000 529.700 312.400 530.200 ;
        RECT 303.000 529.600 304.400 529.700 ;
        RECT 301.400 522.200 302.200 529.600 ;
        RECT 303.000 528.400 303.600 529.600 ;
        RECT 302.800 527.600 303.600 528.400 ;
        RECT 311.600 522.200 312.400 529.700 ;
        RECT 313.200 528.800 314.000 530.400 ;
        RECT 316.200 530.000 317.200 530.800 ;
        RECT 316.400 522.200 317.200 530.000 ;
        RECT 317.800 529.600 318.400 531.400 ;
        RECT 317.800 529.000 326.800 529.600 ;
        RECT 317.800 527.400 318.400 529.000 ;
        RECT 326.000 528.800 326.800 529.000 ;
        RECT 329.200 529.000 337.800 529.600 ;
        RECT 329.200 528.800 330.000 529.000 ;
        RECT 321.000 527.600 323.600 528.400 ;
        RECT 317.800 526.800 320.400 527.400 ;
        RECT 319.600 522.200 320.400 526.800 ;
        RECT 322.800 522.200 323.600 527.600 ;
        RECT 324.200 526.800 328.400 527.600 ;
        RECT 326.000 522.200 326.800 525.000 ;
        RECT 327.600 522.200 328.400 525.000 ;
        RECT 329.200 522.200 330.000 525.000 ;
        RECT 330.800 522.200 331.600 528.400 ;
        RECT 334.000 527.600 336.600 528.400 ;
        RECT 337.200 528.200 337.800 529.000 ;
        RECT 338.800 529.400 339.600 529.600 ;
        RECT 338.800 529.000 344.200 529.400 ;
        RECT 338.800 528.800 345.000 529.000 ;
        RECT 343.600 528.200 345.000 528.800 ;
        RECT 337.200 527.600 343.000 528.200 ;
        RECT 346.000 528.000 347.600 528.800 ;
        RECT 346.000 527.600 346.600 528.000 ;
        RECT 334.000 522.200 334.800 527.000 ;
        RECT 337.200 522.200 338.000 527.000 ;
        RECT 342.400 526.800 346.600 527.600 ;
        RECT 348.400 527.400 349.200 533.000 ;
        RECT 350.000 530.200 350.800 530.400 ;
        RECT 352.000 530.200 352.600 533.600 ;
        RECT 353.200 531.600 354.000 533.200 ;
        RECT 350.000 529.600 351.400 530.200 ;
        RECT 352.000 529.600 353.000 530.200 ;
        RECT 350.800 528.400 351.400 529.600 ;
        RECT 350.800 527.600 351.600 528.400 ;
        RECT 347.200 526.800 349.200 527.400 ;
        RECT 338.800 522.200 339.600 525.000 ;
        RECT 340.400 522.200 341.200 525.000 ;
        RECT 343.600 522.200 344.400 526.800 ;
        RECT 347.200 526.200 347.800 526.800 ;
        RECT 346.800 525.600 347.800 526.200 ;
        RECT 346.800 522.200 347.600 525.600 ;
        RECT 352.200 522.200 353.000 529.600 ;
        RECT 356.400 522.200 357.200 533.700 ;
        RECT 358.000 534.300 358.800 534.400 ;
        RECT 359.600 534.300 362.200 534.400 ;
        RECT 358.000 533.700 362.200 534.300 ;
        RECT 363.600 534.300 365.200 534.400 ;
        RECT 366.000 534.300 367.600 534.400 ;
        RECT 363.600 533.800 367.600 534.300 ;
        RECT 358.000 533.600 358.800 533.700 ;
        RECT 359.600 533.600 362.200 533.700 ;
        RECT 364.400 533.700 366.800 533.800 ;
        RECT 364.400 533.600 365.200 533.700 ;
        RECT 366.000 533.600 366.800 533.700 ;
        RECT 369.000 533.600 371.600 534.400 ;
        RECT 374.000 534.300 374.800 539.800 ;
        RECT 375.600 536.000 376.400 539.800 ;
        RECT 378.800 536.000 379.600 539.800 ;
        RECT 375.600 535.800 379.600 536.000 ;
        RECT 380.400 535.800 381.200 539.800 ;
        RECT 383.600 536.000 384.400 539.800 ;
        RECT 375.800 535.400 379.400 535.800 ;
        RECT 376.400 534.400 377.200 534.800 ;
        RECT 380.400 534.400 381.000 535.800 ;
        RECT 383.400 535.200 384.400 536.000 ;
        RECT 375.600 534.300 377.200 534.400 ;
        RECT 374.000 533.800 377.200 534.300 ;
        RECT 378.600 534.300 381.200 534.400 ;
        RECT 382.000 534.300 382.800 534.400 ;
        RECT 374.000 533.700 376.400 533.800 ;
        RECT 359.600 530.200 360.400 530.400 ;
        RECT 361.600 530.200 362.200 533.600 ;
        RECT 362.800 532.300 363.600 533.200 ;
        RECT 364.400 532.300 365.200 532.400 ;
        RECT 367.600 532.300 368.400 533.200 ;
        RECT 362.800 531.700 368.400 532.300 ;
        RECT 362.800 531.600 363.600 531.700 ;
        RECT 364.400 531.600 365.200 531.700 ;
        RECT 367.600 531.600 368.400 531.700 ;
        RECT 369.000 532.300 369.600 533.600 ;
        RECT 372.400 532.300 373.200 532.400 ;
        RECT 369.000 531.700 373.200 532.300 ;
        RECT 369.000 530.200 369.600 531.700 ;
        RECT 372.400 531.600 373.200 531.700 ;
        RECT 370.800 530.200 371.600 530.400 ;
        RECT 359.600 529.600 361.000 530.200 ;
        RECT 361.600 529.600 362.600 530.200 ;
        RECT 360.400 528.400 361.000 529.600 ;
        RECT 360.400 527.600 361.200 528.400 ;
        RECT 361.800 522.200 362.600 529.600 ;
        RECT 368.600 529.600 369.600 530.200 ;
        RECT 370.200 529.600 371.600 530.200 ;
        RECT 368.600 522.200 369.400 529.600 ;
        RECT 370.200 528.400 370.800 529.600 ;
        RECT 370.000 527.600 370.800 528.400 ;
        RECT 374.000 522.200 374.800 533.700 ;
        RECT 375.600 533.600 376.400 533.700 ;
        RECT 378.600 533.700 382.800 534.300 ;
        RECT 378.600 533.600 381.200 533.700 ;
        RECT 382.000 533.600 382.800 533.700 ;
        RECT 377.200 531.600 378.000 533.200 ;
        RECT 378.600 530.200 379.200 533.600 ;
        RECT 383.400 530.800 384.200 535.200 ;
        RECT 385.200 534.600 386.000 539.800 ;
        RECT 391.600 536.600 392.400 539.800 ;
        RECT 393.200 537.000 394.000 539.800 ;
        RECT 394.800 537.000 395.600 539.800 ;
        RECT 396.400 537.000 397.200 539.800 ;
        RECT 398.000 537.000 398.800 539.800 ;
        RECT 401.200 537.000 402.000 539.800 ;
        RECT 404.400 537.000 405.200 539.800 ;
        RECT 406.000 537.000 406.800 539.800 ;
        RECT 407.600 537.000 408.400 539.800 ;
        RECT 390.000 535.800 392.400 536.600 ;
        RECT 409.200 536.600 410.000 539.800 ;
        RECT 390.000 535.200 390.800 535.800 ;
        RECT 384.800 534.000 386.000 534.600 ;
        RECT 389.000 534.600 390.800 535.200 ;
        RECT 394.800 535.600 395.800 536.400 ;
        RECT 398.800 535.600 400.400 536.400 ;
        RECT 401.200 535.800 405.800 536.400 ;
        RECT 409.200 535.800 411.800 536.600 ;
        RECT 401.200 535.600 402.000 535.800 ;
        RECT 384.800 532.000 385.400 534.000 ;
        RECT 389.000 533.400 389.800 534.600 ;
        RECT 386.000 532.600 389.800 533.400 ;
        RECT 394.800 532.800 395.600 535.600 ;
        RECT 401.200 534.800 402.000 535.000 ;
        RECT 397.600 534.200 402.000 534.800 ;
        RECT 397.600 534.000 398.400 534.200 ;
        RECT 402.800 533.600 403.600 535.200 ;
        RECT 405.000 533.400 405.800 535.800 ;
        RECT 411.000 535.200 411.800 535.800 ;
        RECT 411.000 534.400 414.000 535.200 ;
        RECT 415.600 533.800 416.400 539.800 ;
        RECT 418.800 535.200 419.600 539.800 ;
        RECT 422.000 535.200 422.800 539.800 ;
        RECT 425.200 535.200 426.000 539.800 ;
        RECT 428.400 535.200 429.200 539.800 ;
        RECT 398.000 532.600 401.200 533.400 ;
        RECT 405.000 532.600 407.000 533.400 ;
        RECT 407.600 533.000 416.400 533.800 ;
        RECT 391.600 532.000 392.400 532.600 ;
        RECT 409.200 532.000 410.000 532.400 ;
        RECT 412.400 532.000 413.200 532.400 ;
        RECT 414.200 532.000 415.000 532.200 ;
        RECT 384.800 531.400 385.600 532.000 ;
        RECT 391.600 531.400 415.000 532.000 ;
        RECT 380.400 530.200 381.200 530.400 ;
        RECT 378.200 529.600 379.200 530.200 ;
        RECT 379.800 529.600 381.200 530.200 ;
        RECT 383.400 530.000 384.400 530.800 ;
        RECT 378.200 522.200 379.000 529.600 ;
        RECT 379.800 528.400 380.400 529.600 ;
        RECT 379.600 527.600 380.400 528.400 ;
        RECT 383.600 522.200 384.400 530.000 ;
        RECT 385.000 529.600 385.600 531.400 ;
        RECT 385.000 529.000 394.000 529.600 ;
        RECT 385.000 527.400 385.600 529.000 ;
        RECT 393.200 528.800 394.000 529.000 ;
        RECT 396.400 529.000 405.000 529.600 ;
        RECT 396.400 528.800 397.200 529.000 ;
        RECT 388.200 527.600 390.800 528.400 ;
        RECT 385.000 526.800 387.600 527.400 ;
        RECT 386.800 522.200 387.600 526.800 ;
        RECT 390.000 522.200 390.800 527.600 ;
        RECT 391.400 526.800 395.600 527.600 ;
        RECT 393.200 522.200 394.000 525.000 ;
        RECT 394.800 522.200 395.600 525.000 ;
        RECT 396.400 522.200 397.200 525.000 ;
        RECT 398.000 522.200 398.800 528.400 ;
        RECT 401.200 527.600 403.800 528.400 ;
        RECT 404.400 528.200 405.000 529.000 ;
        RECT 406.000 529.400 406.800 529.600 ;
        RECT 406.000 529.000 411.400 529.400 ;
        RECT 406.000 528.800 412.200 529.000 ;
        RECT 410.800 528.200 412.200 528.800 ;
        RECT 404.400 527.600 410.200 528.200 ;
        RECT 413.200 528.000 414.800 528.800 ;
        RECT 413.200 527.600 413.800 528.000 ;
        RECT 401.200 522.200 402.000 527.000 ;
        RECT 404.400 522.200 405.200 527.000 ;
        RECT 409.600 526.800 413.800 527.600 ;
        RECT 415.600 527.400 416.400 533.000 ;
        RECT 417.200 534.400 419.600 535.200 ;
        RECT 420.600 534.400 422.800 535.200 ;
        RECT 423.800 534.400 426.000 535.200 ;
        RECT 427.400 534.400 429.200 535.200 ;
        RECT 431.600 535.400 432.400 539.800 ;
        RECT 435.800 538.400 437.000 539.800 ;
        RECT 435.800 537.800 437.200 538.400 ;
        RECT 440.400 537.800 441.200 539.800 ;
        RECT 444.800 538.400 445.600 539.800 ;
        RECT 444.800 537.800 446.800 538.400 ;
        RECT 436.400 537.000 437.200 537.800 ;
        RECT 440.600 537.200 441.200 537.800 ;
        RECT 440.600 536.600 443.400 537.200 ;
        RECT 442.600 536.400 443.400 536.600 ;
        RECT 444.400 536.400 445.200 537.200 ;
        RECT 446.000 537.000 446.800 537.800 ;
        RECT 434.600 535.400 435.400 535.600 ;
        RECT 431.600 534.800 435.400 535.400 ;
        RECT 417.200 531.600 418.000 534.400 ;
        RECT 420.600 533.800 421.400 534.400 ;
        RECT 423.800 533.800 424.600 534.400 ;
        RECT 427.400 533.800 428.200 534.400 ;
        RECT 430.000 533.800 430.800 534.400 ;
        RECT 418.800 533.000 421.400 533.800 ;
        RECT 422.200 533.000 424.600 533.800 ;
        RECT 425.600 533.000 428.200 533.800 ;
        RECT 429.000 533.000 430.800 533.800 ;
        RECT 420.600 531.600 421.400 533.000 ;
        RECT 423.800 531.600 424.600 533.000 ;
        RECT 427.400 531.600 428.200 533.000 ;
        RECT 417.200 530.800 419.600 531.600 ;
        RECT 420.600 530.800 422.800 531.600 ;
        RECT 423.800 530.800 426.000 531.600 ;
        RECT 427.400 530.800 429.200 531.600 ;
        RECT 414.400 526.800 416.400 527.400 ;
        RECT 406.000 522.200 406.800 525.000 ;
        RECT 407.600 522.200 408.400 525.000 ;
        RECT 410.800 522.200 411.600 526.800 ;
        RECT 414.400 526.200 415.000 526.800 ;
        RECT 414.000 525.600 415.000 526.200 ;
        RECT 414.000 522.200 414.800 525.600 ;
        RECT 418.800 522.200 419.600 530.800 ;
        RECT 422.000 522.200 422.800 530.800 ;
        RECT 425.200 522.200 426.000 530.800 ;
        RECT 428.400 522.200 429.200 530.800 ;
        RECT 431.600 531.400 432.400 534.800 ;
        RECT 438.600 534.200 439.400 534.400 ;
        RECT 444.400 534.200 445.000 536.400 ;
        RECT 449.200 535.000 450.000 539.800 ;
        RECT 450.800 536.000 451.600 539.800 ;
        RECT 454.000 536.000 454.800 539.800 ;
        RECT 450.800 535.800 454.800 536.000 ;
        RECT 455.600 535.800 456.400 539.800 ;
        RECT 462.000 535.800 462.800 539.800 ;
        RECT 463.600 536.000 464.400 539.800 ;
        RECT 466.800 536.000 467.600 539.800 ;
        RECT 463.600 535.800 467.600 536.000 ;
        RECT 451.000 535.400 454.600 535.800 ;
        RECT 451.600 534.400 452.400 534.800 ;
        RECT 455.600 534.400 456.200 535.800 ;
        RECT 462.200 534.400 462.800 535.800 ;
        RECT 463.800 535.400 467.400 535.800 ;
        RECT 468.400 535.200 469.200 539.800 ;
        RECT 471.600 536.400 472.400 539.800 ;
        RECT 471.600 535.800 472.600 536.400 ;
        RECT 474.800 536.000 475.600 539.800 ;
        RECT 478.000 536.000 478.800 539.800 ;
        RECT 474.800 535.800 478.800 536.000 ;
        RECT 479.600 535.800 480.400 539.800 ;
        RECT 481.200 535.800 482.000 539.800 ;
        RECT 482.800 536.000 483.600 539.800 ;
        RECT 486.000 536.000 486.800 539.800 ;
        RECT 482.800 535.800 486.800 536.000 ;
        RECT 487.600 536.000 488.400 539.800 ;
        RECT 490.800 536.000 491.600 539.800 ;
        RECT 487.600 535.800 491.600 536.000 ;
        RECT 492.400 535.800 493.200 539.800 ;
        RECT 494.000 535.800 494.800 539.800 ;
        RECT 495.600 536.000 496.400 539.800 ;
        RECT 498.800 536.000 499.600 539.800 ;
        RECT 495.600 535.800 499.600 536.000 ;
        RECT 466.000 534.400 466.800 534.800 ;
        RECT 468.400 534.600 471.000 535.200 ;
        RECT 447.600 534.200 449.200 534.400 ;
        RECT 438.200 533.600 449.200 534.200 ;
        RECT 450.800 533.800 452.400 534.400 ;
        RECT 450.800 533.600 451.600 533.800 ;
        RECT 453.800 533.600 456.400 534.400 ;
        RECT 462.000 533.600 464.600 534.400 ;
        RECT 466.000 533.800 467.600 534.400 ;
        RECT 466.800 533.600 467.600 533.800 ;
        RECT 436.400 532.800 437.200 533.000 ;
        RECT 433.400 532.200 437.200 532.800 ;
        RECT 438.200 532.400 438.800 533.600 ;
        RECT 445.400 533.400 446.200 533.600 ;
        RECT 444.400 532.400 445.200 532.600 ;
        RECT 447.000 532.400 447.800 532.600 ;
        RECT 433.400 532.000 434.200 532.200 ;
        RECT 438.000 531.600 438.800 532.400 ;
        RECT 442.800 531.800 447.800 532.400 ;
        RECT 442.800 531.600 443.600 531.800 ;
        RECT 452.400 531.600 453.200 533.200 ;
        RECT 435.000 531.400 435.800 531.600 ;
        RECT 431.600 530.800 435.800 531.400 ;
        RECT 431.600 522.200 432.400 530.800 ;
        RECT 438.200 530.400 438.800 531.600 ;
        RECT 444.400 531.000 450.000 531.200 ;
        RECT 444.200 530.800 450.000 531.000 ;
        RECT 436.400 529.800 438.800 530.400 ;
        RECT 440.200 530.600 450.000 530.800 ;
        RECT 440.200 530.200 445.000 530.600 ;
        RECT 436.400 528.800 437.000 529.800 ;
        RECT 435.600 528.000 437.000 528.800 ;
        RECT 438.600 529.000 439.400 529.200 ;
        RECT 440.200 529.000 440.800 530.200 ;
        RECT 438.600 528.400 440.800 529.000 ;
        RECT 441.400 529.000 446.800 529.600 ;
        RECT 441.400 528.800 442.200 529.000 ;
        RECT 446.000 528.800 446.800 529.000 ;
        RECT 439.800 527.400 440.600 527.600 ;
        RECT 442.600 527.400 443.400 527.600 ;
        RECT 436.400 526.200 437.200 527.000 ;
        RECT 439.800 526.800 443.400 527.400 ;
        RECT 440.600 526.200 441.200 526.800 ;
        RECT 446.000 526.200 446.800 527.000 ;
        RECT 435.800 522.200 437.000 526.200 ;
        RECT 440.400 522.200 441.200 526.200 ;
        RECT 444.800 525.600 446.800 526.200 ;
        RECT 444.800 522.200 445.600 525.600 ;
        RECT 449.200 522.200 450.000 530.600 ;
        RECT 453.800 530.200 454.400 533.600 ;
        RECT 464.000 532.300 464.600 533.600 ;
        RECT 455.700 531.700 464.600 532.300 ;
        RECT 455.700 530.400 456.300 531.700 ;
        RECT 455.600 530.200 456.400 530.400 ;
        RECT 453.400 529.600 454.400 530.200 ;
        RECT 455.000 529.600 456.400 530.200 ;
        RECT 462.000 530.200 462.800 530.400 ;
        RECT 464.000 530.200 464.600 531.700 ;
        RECT 465.200 531.600 466.000 533.200 ;
        RECT 468.600 532.400 469.400 533.200 ;
        RECT 466.800 532.300 467.600 532.400 ;
        RECT 468.400 532.300 469.400 532.400 ;
        RECT 466.800 531.700 469.400 532.300 ;
        RECT 466.800 531.600 467.600 531.700 ;
        RECT 468.400 531.600 469.400 531.700 ;
        RECT 470.400 533.000 471.000 534.600 ;
        RECT 472.000 534.400 472.600 535.800 ;
        RECT 475.000 535.400 478.600 535.800 ;
        RECT 475.600 534.400 476.400 534.800 ;
        RECT 479.600 534.400 480.200 535.800 ;
        RECT 481.400 534.400 482.000 535.800 ;
        RECT 483.000 535.400 486.600 535.800 ;
        RECT 487.800 535.400 491.400 535.800 ;
        RECT 485.200 534.400 486.000 534.800 ;
        RECT 488.400 534.400 489.200 534.800 ;
        RECT 492.400 534.400 493.000 535.800 ;
        RECT 494.200 534.400 494.800 535.800 ;
        RECT 495.800 535.400 499.400 535.800 ;
        RECT 500.400 535.000 501.200 539.800 ;
        RECT 504.800 538.400 505.600 539.800 ;
        RECT 503.600 537.800 505.600 538.400 ;
        RECT 509.200 537.800 510.000 539.800 ;
        RECT 513.400 538.400 514.600 539.800 ;
        RECT 513.200 537.800 514.600 538.400 ;
        RECT 503.600 537.000 504.400 537.800 ;
        RECT 509.200 537.200 509.800 537.800 ;
        RECT 505.200 536.400 506.000 537.200 ;
        RECT 507.000 536.600 509.800 537.200 ;
        RECT 513.200 537.000 514.000 537.800 ;
        RECT 507.000 536.400 507.800 536.600 ;
        RECT 498.000 534.400 498.800 534.800 ;
        RECT 471.600 533.600 472.600 534.400 ;
        RECT 474.800 533.800 476.400 534.400 ;
        RECT 474.800 533.600 475.600 533.800 ;
        RECT 477.800 533.600 480.400 534.400 ;
        RECT 481.200 533.600 483.800 534.400 ;
        RECT 485.200 533.800 486.800 534.400 ;
        RECT 486.000 533.600 486.800 533.800 ;
        RECT 487.600 533.800 489.200 534.400 ;
        RECT 487.600 533.600 488.400 533.800 ;
        RECT 490.600 533.600 493.200 534.400 ;
        RECT 494.000 533.600 496.600 534.400 ;
        RECT 498.000 533.800 499.600 534.400 ;
        RECT 498.800 533.600 499.600 533.800 ;
        RECT 501.200 534.200 502.800 534.400 ;
        RECT 505.400 534.200 506.000 536.400 ;
        RECT 515.000 535.400 515.800 535.600 ;
        RECT 518.000 535.400 518.800 539.800 ;
        RECT 520.200 536.400 521.000 539.800 ;
        RECT 520.200 535.800 522.000 536.400 ;
        RECT 515.000 534.800 518.800 535.400 ;
        RECT 511.000 534.200 511.800 534.400 ;
        RECT 501.200 533.600 512.200 534.200 ;
        RECT 470.400 532.200 471.400 533.000 ;
        RECT 470.400 530.200 471.000 532.200 ;
        RECT 472.000 530.200 472.600 533.600 ;
        RECT 473.200 532.300 474.000 532.400 ;
        RECT 476.400 532.300 477.200 533.200 ;
        RECT 473.200 531.700 477.200 532.300 ;
        RECT 473.200 531.600 474.000 531.700 ;
        RECT 476.400 531.600 477.200 531.700 ;
        RECT 477.800 530.200 478.400 533.600 ;
        RECT 483.200 532.300 483.800 533.600 ;
        RECT 479.700 531.700 483.800 532.300 ;
        RECT 479.700 530.400 480.300 531.700 ;
        RECT 479.600 530.200 480.400 530.400 ;
        RECT 462.000 529.600 463.400 530.200 ;
        RECT 464.000 529.600 465.000 530.200 ;
        RECT 453.400 528.400 454.200 529.600 ;
        RECT 455.000 528.400 455.600 529.600 ;
        RECT 452.400 527.600 454.200 528.400 ;
        RECT 454.800 527.600 455.600 528.400 ;
        RECT 462.800 528.400 463.400 529.600 ;
        RECT 462.800 527.600 463.600 528.400 ;
        RECT 453.400 522.200 454.200 527.600 ;
        RECT 464.200 522.200 465.000 529.600 ;
        RECT 468.400 529.600 471.000 530.200 ;
        RECT 468.400 522.200 469.200 529.600 ;
        RECT 471.600 529.200 472.600 530.200 ;
        RECT 477.400 529.600 478.400 530.200 ;
        RECT 479.000 529.600 480.400 530.200 ;
        RECT 481.200 530.200 482.000 530.400 ;
        RECT 483.200 530.200 483.800 531.700 ;
        RECT 484.400 531.600 485.200 533.200 ;
        RECT 489.200 531.600 490.000 533.200 ;
        RECT 490.600 530.200 491.200 533.600 ;
        RECT 496.000 532.300 496.600 533.600 ;
        RECT 504.200 533.400 505.000 533.600 ;
        RECT 492.500 531.700 496.600 532.300 ;
        RECT 492.500 530.400 493.100 531.700 ;
        RECT 492.400 530.200 493.200 530.400 ;
        RECT 481.200 529.600 482.600 530.200 ;
        RECT 483.200 529.600 484.200 530.200 ;
        RECT 471.600 522.200 472.400 529.200 ;
        RECT 477.400 522.200 478.200 529.600 ;
        RECT 479.000 528.400 479.600 529.600 ;
        RECT 478.800 527.600 479.600 528.400 ;
        RECT 482.000 528.400 482.600 529.600 ;
        RECT 482.000 527.600 482.800 528.400 ;
        RECT 483.400 522.200 484.200 529.600 ;
        RECT 490.200 529.600 491.200 530.200 ;
        RECT 491.800 529.600 493.200 530.200 ;
        RECT 494.000 530.200 494.800 530.400 ;
        RECT 496.000 530.200 496.600 531.700 ;
        RECT 497.200 531.600 498.000 533.200 ;
        RECT 502.600 532.400 503.400 532.600 ;
        RECT 505.200 532.400 506.000 532.600 ;
        RECT 502.600 531.800 507.600 532.400 ;
        RECT 506.800 531.600 507.600 531.800 ;
        RECT 500.400 531.000 506.000 531.200 ;
        RECT 500.400 530.800 506.200 531.000 ;
        RECT 500.400 530.600 510.200 530.800 ;
        RECT 494.000 529.600 495.400 530.200 ;
        RECT 496.000 529.600 497.000 530.200 ;
        RECT 490.200 522.200 491.000 529.600 ;
        RECT 491.800 528.400 492.400 529.600 ;
        RECT 491.600 527.600 492.400 528.400 ;
        RECT 494.800 528.400 495.400 529.600 ;
        RECT 494.800 527.600 495.600 528.400 ;
        RECT 496.200 522.200 497.000 529.600 ;
        RECT 500.400 522.200 501.200 530.600 ;
        RECT 505.400 530.200 510.200 530.600 ;
        RECT 503.600 529.000 509.000 529.600 ;
        RECT 503.600 528.800 504.400 529.000 ;
        RECT 508.200 528.800 509.000 529.000 ;
        RECT 509.600 529.000 510.200 530.200 ;
        RECT 511.600 530.400 512.200 533.600 ;
        RECT 513.200 532.800 514.000 533.000 ;
        RECT 513.200 532.200 517.000 532.800 ;
        RECT 516.200 532.000 517.000 532.200 ;
        RECT 514.600 531.400 515.400 531.600 ;
        RECT 518.000 531.400 518.800 534.800 ;
        RECT 514.600 530.800 518.800 531.400 ;
        RECT 511.600 529.800 514.000 530.400 ;
        RECT 511.000 529.000 511.800 529.200 ;
        RECT 509.600 528.400 511.800 529.000 ;
        RECT 513.400 528.800 514.000 529.800 ;
        RECT 513.400 528.000 514.800 528.800 ;
        RECT 507.000 527.400 507.800 527.600 ;
        RECT 509.800 527.400 510.600 527.600 ;
        RECT 503.600 526.200 504.400 527.000 ;
        RECT 507.000 526.800 510.600 527.400 ;
        RECT 509.200 526.200 509.800 526.800 ;
        RECT 513.200 526.200 514.000 527.000 ;
        RECT 503.600 525.600 505.600 526.200 ;
        RECT 504.800 522.200 505.600 525.600 ;
        RECT 509.200 522.200 510.000 526.200 ;
        RECT 513.400 522.200 514.600 526.200 ;
        RECT 518.000 522.200 518.800 530.800 ;
        RECT 519.600 528.800 520.400 530.400 ;
        RECT 521.200 522.200 522.000 535.800 ;
        RECT 524.400 535.200 525.200 539.800 ;
        RECT 527.600 536.400 528.400 539.800 ;
        RECT 527.600 535.800 528.600 536.400 ;
        RECT 522.800 533.600 523.600 535.200 ;
        RECT 524.400 534.600 527.000 535.200 ;
        RECT 524.600 532.400 525.400 533.200 ;
        RECT 522.800 532.300 523.600 532.400 ;
        RECT 524.400 532.300 525.400 532.400 ;
        RECT 522.800 531.700 525.400 532.300 ;
        RECT 522.800 531.600 523.600 531.700 ;
        RECT 524.400 531.600 525.400 531.700 ;
        RECT 526.400 533.000 527.000 534.600 ;
        RECT 528.000 534.400 528.600 535.800 ;
        RECT 530.800 535.200 531.600 539.800 ;
        RECT 534.000 536.400 534.800 539.800 ;
        RECT 534.000 535.800 535.000 536.400 ;
        RECT 537.200 536.000 538.000 539.800 ;
        RECT 540.400 536.000 541.200 539.800 ;
        RECT 537.200 535.800 541.200 536.000 ;
        RECT 542.000 536.300 542.800 539.800 ;
        RECT 543.600 536.300 544.400 536.400 ;
        RECT 530.800 534.600 533.400 535.200 ;
        RECT 527.600 533.600 528.600 534.400 ;
        RECT 526.400 532.200 527.400 533.000 ;
        RECT 526.400 530.200 527.000 532.200 ;
        RECT 528.000 530.200 528.600 533.600 ;
        RECT 531.000 532.400 531.800 533.200 ;
        RECT 530.800 531.600 531.800 532.400 ;
        RECT 532.800 533.000 533.400 534.600 ;
        RECT 534.400 534.400 535.000 535.800 ;
        RECT 537.400 535.400 541.000 535.800 ;
        RECT 542.000 535.700 544.400 536.300 ;
        RECT 545.200 536.000 546.000 539.800 ;
        RECT 538.000 534.400 538.800 534.800 ;
        RECT 542.000 534.400 542.600 535.700 ;
        RECT 543.600 535.600 544.400 535.700 ;
        RECT 545.000 535.200 546.000 536.000 ;
        RECT 534.000 533.600 535.000 534.400 ;
        RECT 537.200 533.800 538.800 534.400 ;
        RECT 537.200 533.600 538.000 533.800 ;
        RECT 540.200 533.600 542.800 534.400 ;
        RECT 532.800 532.200 533.800 533.000 ;
        RECT 532.800 530.200 533.400 532.200 ;
        RECT 534.400 530.200 535.000 533.600 ;
        RECT 538.800 531.600 539.600 533.200 ;
        RECT 540.200 530.200 540.800 533.600 ;
        RECT 545.000 530.800 545.800 535.200 ;
        RECT 546.800 534.600 547.600 539.800 ;
        RECT 553.200 536.600 554.000 539.800 ;
        RECT 554.800 537.000 555.600 539.800 ;
        RECT 556.400 537.000 557.200 539.800 ;
        RECT 558.000 537.000 558.800 539.800 ;
        RECT 559.600 537.000 560.400 539.800 ;
        RECT 562.800 537.000 563.600 539.800 ;
        RECT 566.000 537.000 566.800 539.800 ;
        RECT 567.600 537.000 568.400 539.800 ;
        RECT 569.200 537.000 570.000 539.800 ;
        RECT 551.600 535.800 554.000 536.600 ;
        RECT 570.800 536.600 571.600 539.800 ;
        RECT 551.600 535.200 552.400 535.800 ;
        RECT 546.400 534.000 547.600 534.600 ;
        RECT 550.600 534.600 552.400 535.200 ;
        RECT 556.400 535.600 557.400 536.400 ;
        RECT 560.400 535.600 562.000 536.400 ;
        RECT 562.800 535.800 567.400 536.400 ;
        RECT 570.800 535.800 573.400 536.600 ;
        RECT 562.800 535.600 563.600 535.800 ;
        RECT 546.400 532.000 547.000 534.000 ;
        RECT 550.600 533.400 551.400 534.600 ;
        RECT 547.600 532.600 551.400 533.400 ;
        RECT 556.400 532.800 557.200 535.600 ;
        RECT 562.800 534.800 563.600 535.000 ;
        RECT 559.200 534.200 563.600 534.800 ;
        RECT 559.200 534.000 560.000 534.200 ;
        RECT 564.400 533.600 565.200 535.200 ;
        RECT 566.600 533.400 567.400 535.800 ;
        RECT 572.600 535.200 573.400 535.800 ;
        RECT 572.600 534.400 575.600 535.200 ;
        RECT 577.200 533.800 578.000 539.800 ;
        RECT 578.800 536.000 579.600 539.800 ;
        RECT 582.000 536.000 582.800 539.800 ;
        RECT 578.800 535.800 582.800 536.000 ;
        RECT 583.600 535.800 584.400 539.800 ;
        RECT 579.000 535.400 582.600 535.800 ;
        RECT 579.600 534.400 580.400 534.800 ;
        RECT 583.600 534.400 584.200 535.800 ;
        RECT 586.800 535.200 587.600 539.800 ;
        RECT 590.000 535.200 590.800 539.800 ;
        RECT 593.200 535.200 594.000 539.800 ;
        RECT 596.400 535.200 597.200 539.800 ;
        RECT 599.600 535.800 600.400 539.800 ;
        RECT 601.200 536.000 602.000 539.800 ;
        RECT 604.400 536.000 605.200 539.800 ;
        RECT 601.200 535.800 605.200 536.000 ;
        RECT 585.200 534.400 587.600 535.200 ;
        RECT 588.600 534.400 590.800 535.200 ;
        RECT 591.800 534.400 594.000 535.200 ;
        RECT 595.400 534.400 597.200 535.200 ;
        RECT 599.800 534.400 600.400 535.800 ;
        RECT 601.400 535.400 605.000 535.800 ;
        RECT 603.600 534.400 604.400 534.800 ;
        RECT 559.600 532.600 562.800 533.400 ;
        RECT 566.600 532.600 568.600 533.400 ;
        RECT 569.200 533.000 578.000 533.800 ;
        RECT 578.800 533.800 580.400 534.400 ;
        RECT 578.800 533.600 579.600 533.800 ;
        RECT 581.800 533.600 584.400 534.400 ;
        RECT 553.200 532.000 554.000 532.600 ;
        RECT 570.800 532.000 571.600 532.400 ;
        RECT 572.400 532.000 573.200 532.400 ;
        RECT 575.800 532.000 576.600 532.200 ;
        RECT 546.400 531.400 547.200 532.000 ;
        RECT 553.200 531.400 576.600 532.000 ;
        RECT 542.000 530.300 542.800 530.400 ;
        RECT 543.600 530.300 544.400 530.400 ;
        RECT 542.000 530.200 544.400 530.300 ;
        RECT 524.400 529.600 527.000 530.200 ;
        RECT 524.400 522.200 525.200 529.600 ;
        RECT 527.600 529.200 528.600 530.200 ;
        RECT 530.800 529.600 533.400 530.200 ;
        RECT 527.600 522.200 528.400 529.200 ;
        RECT 530.800 522.200 531.600 529.600 ;
        RECT 534.000 529.200 535.000 530.200 ;
        RECT 539.800 529.600 540.800 530.200 ;
        RECT 541.400 529.700 544.400 530.200 ;
        RECT 545.000 530.000 546.000 530.800 ;
        RECT 541.400 529.600 542.800 529.700 ;
        RECT 543.600 529.600 544.400 529.700 ;
        RECT 534.000 522.200 534.800 529.200 ;
        RECT 539.800 522.200 540.600 529.600 ;
        RECT 541.400 528.400 542.000 529.600 ;
        RECT 541.200 527.600 542.000 528.400 ;
        RECT 545.200 522.200 546.000 530.000 ;
        RECT 546.600 529.600 547.200 531.400 ;
        RECT 546.600 529.000 555.600 529.600 ;
        RECT 546.600 527.400 547.200 529.000 ;
        RECT 554.800 528.800 555.600 529.000 ;
        RECT 558.000 529.000 566.600 529.600 ;
        RECT 558.000 528.800 558.800 529.000 ;
        RECT 549.800 527.600 552.400 528.400 ;
        RECT 546.600 526.800 549.200 527.400 ;
        RECT 548.400 522.200 549.200 526.800 ;
        RECT 551.600 522.200 552.400 527.600 ;
        RECT 553.000 526.800 557.200 527.600 ;
        RECT 554.800 522.200 555.600 525.000 ;
        RECT 556.400 522.200 557.200 525.000 ;
        RECT 558.000 522.200 558.800 525.000 ;
        RECT 559.600 522.200 560.400 528.400 ;
        RECT 562.800 527.600 565.400 528.400 ;
        RECT 566.000 528.200 566.600 529.000 ;
        RECT 567.600 529.400 568.400 529.600 ;
        RECT 567.600 529.000 573.000 529.400 ;
        RECT 567.600 528.800 573.800 529.000 ;
        RECT 572.400 528.200 573.800 528.800 ;
        RECT 566.000 527.600 571.800 528.200 ;
        RECT 574.800 528.000 576.400 528.800 ;
        RECT 574.800 527.600 575.400 528.000 ;
        RECT 562.800 522.200 563.600 527.000 ;
        RECT 566.000 522.200 566.800 527.000 ;
        RECT 571.200 526.800 575.400 527.600 ;
        RECT 577.200 527.400 578.000 533.000 ;
        RECT 580.400 531.600 581.200 533.200 ;
        RECT 581.800 532.400 582.400 533.600 ;
        RECT 581.800 531.600 582.800 532.400 ;
        RECT 585.200 531.600 586.000 534.400 ;
        RECT 588.600 533.800 589.400 534.400 ;
        RECT 591.800 533.800 592.600 534.400 ;
        RECT 595.400 533.800 596.200 534.400 ;
        RECT 598.000 533.800 598.800 534.400 ;
        RECT 586.800 533.000 589.400 533.800 ;
        RECT 590.200 533.000 592.600 533.800 ;
        RECT 593.600 533.000 596.200 533.800 ;
        RECT 597.000 533.000 598.800 533.800 ;
        RECT 599.600 533.600 602.200 534.400 ;
        RECT 603.600 534.300 605.200 534.400 ;
        RECT 606.000 534.300 606.800 539.800 ;
        RECT 603.600 533.800 606.800 534.300 ;
        RECT 604.400 533.700 606.800 533.800 ;
        RECT 604.400 533.600 605.200 533.700 ;
        RECT 588.600 531.600 589.400 533.000 ;
        RECT 591.800 531.600 592.600 533.000 ;
        RECT 595.400 531.600 596.200 533.000 ;
        RECT 598.000 532.300 598.800 532.400 ;
        RECT 601.600 532.300 602.200 533.600 ;
        RECT 598.000 531.700 602.200 532.300 ;
        RECT 598.000 531.600 598.800 531.700 ;
        RECT 581.800 530.200 582.400 531.600 ;
        RECT 585.200 530.800 587.600 531.600 ;
        RECT 588.600 530.800 590.800 531.600 ;
        RECT 591.800 530.800 594.000 531.600 ;
        RECT 595.400 530.800 597.200 531.600 ;
        RECT 583.600 530.200 584.400 530.400 ;
        RECT 576.000 526.800 578.000 527.400 ;
        RECT 581.400 529.600 582.400 530.200 ;
        RECT 583.000 529.600 584.400 530.200 ;
        RECT 567.600 522.200 568.400 525.000 ;
        RECT 569.200 522.200 570.000 525.000 ;
        RECT 572.400 522.200 573.200 526.800 ;
        RECT 576.000 526.200 576.600 526.800 ;
        RECT 575.600 525.600 576.600 526.200 ;
        RECT 575.600 522.200 576.400 525.600 ;
        RECT 581.400 522.200 582.200 529.600 ;
        RECT 583.000 528.400 583.600 529.600 ;
        RECT 582.800 527.600 584.400 528.400 ;
        RECT 586.800 522.200 587.600 530.800 ;
        RECT 590.000 522.200 590.800 530.800 ;
        RECT 593.200 522.200 594.000 530.800 ;
        RECT 596.400 522.200 597.200 530.800 ;
        RECT 599.600 530.200 600.400 530.400 ;
        RECT 601.600 530.200 602.200 531.700 ;
        RECT 602.800 531.600 603.600 533.200 ;
        RECT 599.600 529.600 601.000 530.200 ;
        RECT 601.600 529.600 602.600 530.200 ;
        RECT 600.400 528.400 601.000 529.600 ;
        RECT 600.400 527.600 601.200 528.400 ;
        RECT 601.800 522.200 602.600 529.600 ;
        RECT 606.000 522.200 606.800 533.700 ;
        RECT 1.200 511.400 2.000 519.800 ;
        RECT 5.600 516.400 6.400 519.800 ;
        RECT 4.400 515.800 6.400 516.400 ;
        RECT 10.000 515.800 10.800 519.800 ;
        RECT 14.200 515.800 15.400 519.800 ;
        RECT 4.400 515.000 5.200 515.800 ;
        RECT 10.000 515.200 10.600 515.800 ;
        RECT 7.800 514.600 11.400 515.200 ;
        RECT 14.000 515.000 14.800 515.800 ;
        RECT 7.800 514.400 8.600 514.600 ;
        RECT 10.600 514.400 11.400 514.600 ;
        RECT 4.400 513.000 5.200 513.200 ;
        RECT 9.000 513.000 9.800 513.200 ;
        RECT 4.400 512.400 9.800 513.000 ;
        RECT 10.400 513.000 12.600 513.600 ;
        RECT 10.400 511.800 11.000 513.000 ;
        RECT 11.800 512.800 12.600 513.000 ;
        RECT 14.200 513.200 15.600 514.000 ;
        RECT 14.200 512.200 14.800 513.200 ;
        RECT 6.200 511.400 11.000 511.800 ;
        RECT 1.200 511.200 11.000 511.400 ;
        RECT 12.400 511.600 14.800 512.200 ;
        RECT 1.200 511.000 7.000 511.200 ;
        RECT 1.200 510.800 6.800 511.000 ;
        RECT 12.400 510.400 13.000 511.600 ;
        RECT 18.800 511.200 19.600 519.800 ;
        RECT 15.400 510.600 19.600 511.200 ;
        RECT 20.400 511.400 21.200 519.800 ;
        RECT 24.800 516.400 25.600 519.800 ;
        RECT 23.600 515.800 25.600 516.400 ;
        RECT 29.200 515.800 30.000 519.800 ;
        RECT 33.400 515.800 34.600 519.800 ;
        RECT 23.600 515.000 24.400 515.800 ;
        RECT 29.200 515.200 29.800 515.800 ;
        RECT 27.000 514.600 30.600 515.200 ;
        RECT 33.200 515.000 34.000 515.800 ;
        RECT 27.000 514.400 27.800 514.600 ;
        RECT 29.800 514.400 30.600 514.600 ;
        RECT 23.600 513.000 24.400 513.200 ;
        RECT 28.200 513.000 29.000 513.200 ;
        RECT 23.600 512.400 29.000 513.000 ;
        RECT 29.600 513.000 31.800 513.600 ;
        RECT 29.600 511.800 30.200 513.000 ;
        RECT 31.000 512.800 31.800 513.000 ;
        RECT 33.400 513.200 34.800 514.000 ;
        RECT 33.400 512.200 34.000 513.200 ;
        RECT 25.400 511.400 30.200 511.800 ;
        RECT 20.400 511.200 30.200 511.400 ;
        RECT 31.600 511.600 34.000 512.200 ;
        RECT 20.400 511.000 26.200 511.200 ;
        RECT 20.400 510.800 26.000 511.000 ;
        RECT 15.400 510.400 16.200 510.600 ;
        RECT 7.600 510.200 8.400 510.400 ;
        RECT 3.400 509.600 8.400 510.200 ;
        RECT 12.400 509.600 13.200 510.400 ;
        RECT 17.000 509.800 17.800 510.000 ;
        RECT 3.400 509.400 4.200 509.600 ;
        RECT 6.000 509.400 6.800 509.600 ;
        RECT 5.000 508.400 5.800 508.600 ;
        RECT 12.400 508.400 13.000 509.600 ;
        RECT 14.000 509.200 17.800 509.800 ;
        RECT 14.000 509.000 14.800 509.200 ;
        RECT 2.000 507.800 13.000 508.400 ;
        RECT 2.000 507.600 3.600 507.800 ;
        RECT 1.200 502.200 2.000 507.000 ;
        RECT 6.200 505.600 6.800 507.800 ;
        RECT 11.800 507.600 12.600 507.800 ;
        RECT 18.800 507.200 19.600 510.600 ;
        RECT 26.800 510.200 27.600 510.400 ;
        RECT 22.600 509.600 27.600 510.200 ;
        RECT 22.600 509.400 23.400 509.600 ;
        RECT 24.200 508.400 25.000 508.600 ;
        RECT 31.600 508.400 32.200 511.600 ;
        RECT 38.000 511.200 38.800 519.800 ;
        RECT 42.200 512.400 43.000 519.800 ;
        RECT 46.000 515.000 46.800 519.000 ;
        RECT 43.600 513.600 44.400 514.400 ;
        RECT 43.800 512.400 44.400 513.600 ;
        RECT 42.200 511.800 43.200 512.400 ;
        RECT 43.800 511.800 45.200 512.400 ;
        RECT 34.600 510.600 38.800 511.200 ;
        RECT 34.600 510.400 35.400 510.600 ;
        RECT 36.200 509.800 37.000 510.000 ;
        RECT 33.200 509.200 37.000 509.800 ;
        RECT 33.200 509.000 34.000 509.200 ;
        RECT 21.200 507.800 32.200 508.400 ;
        RECT 21.200 507.600 22.800 507.800 ;
        RECT 15.800 506.600 19.600 507.200 ;
        RECT 15.800 506.400 16.600 506.600 ;
        RECT 4.400 504.200 5.200 505.000 ;
        RECT 6.000 504.800 6.800 505.600 ;
        RECT 7.800 505.400 8.600 505.600 ;
        RECT 7.800 504.800 10.600 505.400 ;
        RECT 10.000 504.200 10.600 504.800 ;
        RECT 14.000 504.200 14.800 505.000 ;
        RECT 4.400 503.600 6.400 504.200 ;
        RECT 5.600 502.200 6.400 503.600 ;
        RECT 10.000 502.200 10.800 504.200 ;
        RECT 14.000 503.600 15.400 504.200 ;
        RECT 14.200 502.200 15.400 503.600 ;
        RECT 18.800 502.200 19.600 506.600 ;
        RECT 20.400 502.200 21.200 507.000 ;
        RECT 25.400 506.400 26.000 507.800 ;
        RECT 31.000 507.600 31.800 507.800 ;
        RECT 38.000 507.200 38.800 510.600 ;
        RECT 42.600 510.400 43.200 511.800 ;
        RECT 44.400 511.600 45.200 511.800 ;
        RECT 46.000 511.600 46.600 515.000 ;
        RECT 50.200 512.800 51.000 519.800 ;
        RECT 56.400 513.600 57.200 514.400 ;
        RECT 50.200 512.200 51.800 512.800 ;
        RECT 56.400 512.400 57.000 513.600 ;
        RECT 57.800 512.400 58.600 519.800 ;
        RECT 46.000 511.000 49.800 511.600 ;
        RECT 41.200 508.800 42.000 510.400 ;
        RECT 42.600 509.600 43.600 510.400 ;
        RECT 42.600 508.400 43.200 509.600 ;
        RECT 46.000 508.800 46.800 510.400 ;
        RECT 47.600 508.800 48.400 510.400 ;
        RECT 49.200 509.000 49.800 511.000 ;
        RECT 39.600 508.200 40.400 508.400 ;
        RECT 39.600 507.600 41.200 508.200 ;
        RECT 42.600 507.600 45.200 508.400 ;
        RECT 49.200 508.200 50.600 509.000 ;
        RECT 51.200 508.400 51.800 512.200 ;
        RECT 55.600 511.800 57.000 512.400 ;
        RECT 57.600 511.800 58.600 512.400 ;
        RECT 64.600 512.400 65.400 519.800 ;
        RECT 66.000 513.600 66.800 514.400 ;
        RECT 66.200 512.400 66.800 513.600 ;
        RECT 69.200 513.600 70.000 514.400 ;
        RECT 69.200 512.400 69.800 513.600 ;
        RECT 70.600 512.400 71.400 519.800 ;
        RECT 64.600 511.800 65.600 512.400 ;
        RECT 66.200 511.800 67.600 512.400 ;
        RECT 55.600 511.600 56.400 511.800 ;
        RECT 52.400 509.600 53.200 511.200 ;
        RECT 54.000 510.300 54.800 510.400 ;
        RECT 57.600 510.300 58.200 511.800 ;
        RECT 54.000 509.700 58.200 510.300 ;
        RECT 54.000 509.600 54.800 509.700 ;
        RECT 57.600 508.400 58.200 509.700 ;
        RECT 58.800 510.300 59.600 510.400 ;
        RECT 60.400 510.300 61.200 510.400 ;
        RECT 63.600 510.300 64.400 510.400 ;
        RECT 58.800 509.700 64.400 510.300 ;
        RECT 58.800 508.800 59.600 509.700 ;
        RECT 60.400 509.600 61.200 509.700 ;
        RECT 63.600 508.800 64.400 509.700 ;
        RECT 65.000 510.300 65.600 511.800 ;
        RECT 66.800 511.600 67.600 511.800 ;
        RECT 68.400 511.800 69.800 512.400 ;
        RECT 68.400 511.600 69.200 511.800 ;
        RECT 70.400 511.600 72.400 512.400 ;
        RECT 68.500 510.300 69.100 511.600 ;
        RECT 65.000 509.700 69.100 510.300 ;
        RECT 65.000 508.400 65.600 509.700 ;
        RECT 70.400 508.400 71.000 511.600 ;
        RECT 74.800 511.400 75.600 519.800 ;
        RECT 79.200 516.400 80.000 519.800 ;
        RECT 78.000 515.800 80.000 516.400 ;
        RECT 83.600 515.800 84.400 519.800 ;
        RECT 87.800 515.800 89.000 519.800 ;
        RECT 78.000 515.000 78.800 515.800 ;
        RECT 83.600 515.200 84.200 515.800 ;
        RECT 81.400 514.600 85.000 515.200 ;
        RECT 87.600 515.000 88.400 515.800 ;
        RECT 81.400 514.400 82.200 514.600 ;
        RECT 84.200 514.400 85.000 514.600 ;
        RECT 78.000 513.000 78.800 513.200 ;
        RECT 82.600 513.000 83.400 513.200 ;
        RECT 78.000 512.400 83.400 513.000 ;
        RECT 84.000 513.000 86.200 513.600 ;
        RECT 84.000 511.800 84.600 513.000 ;
        RECT 85.400 512.800 86.200 513.000 ;
        RECT 87.800 513.200 89.200 514.000 ;
        RECT 87.800 512.200 88.400 513.200 ;
        RECT 79.800 511.400 84.600 511.800 ;
        RECT 74.800 511.200 84.600 511.400 ;
        RECT 86.000 511.600 88.400 512.200 ;
        RECT 74.800 511.000 80.600 511.200 ;
        RECT 74.800 510.800 80.400 511.000 ;
        RECT 86.000 510.400 86.600 511.600 ;
        RECT 92.400 511.200 93.200 519.800 ;
        RECT 89.000 510.600 93.200 511.200 ;
        RECT 94.000 511.400 94.800 519.800 ;
        RECT 98.400 516.400 99.200 519.800 ;
        RECT 97.200 515.800 99.200 516.400 ;
        RECT 102.800 515.800 103.600 519.800 ;
        RECT 107.000 515.800 108.200 519.800 ;
        RECT 97.200 515.000 98.000 515.800 ;
        RECT 102.800 515.200 103.400 515.800 ;
        RECT 100.600 514.600 104.200 515.200 ;
        RECT 106.800 515.000 107.600 515.800 ;
        RECT 100.600 514.400 101.400 514.600 ;
        RECT 103.400 514.400 104.200 514.600 ;
        RECT 97.200 513.000 98.000 513.200 ;
        RECT 101.800 513.000 102.600 513.200 ;
        RECT 97.200 512.400 102.600 513.000 ;
        RECT 103.200 513.000 105.400 513.600 ;
        RECT 103.200 511.800 103.800 513.000 ;
        RECT 104.600 512.800 105.400 513.000 ;
        RECT 107.000 513.200 108.400 514.000 ;
        RECT 107.000 512.200 107.600 513.200 ;
        RECT 99.000 511.400 103.800 511.800 ;
        RECT 94.000 511.200 103.800 511.400 ;
        RECT 105.200 511.600 107.600 512.200 ;
        RECT 94.000 511.000 99.800 511.200 ;
        RECT 94.000 510.800 99.600 511.000 ;
        RECT 89.000 510.400 89.800 510.600 ;
        RECT 71.600 508.800 72.400 510.400 ;
        RECT 81.200 510.200 82.000 510.400 ;
        RECT 77.000 509.600 82.000 510.200 ;
        RECT 86.000 509.600 86.800 510.400 ;
        RECT 90.600 509.800 91.400 510.000 ;
        RECT 77.000 509.400 77.800 509.600 ;
        RECT 79.600 509.400 80.400 509.600 ;
        RECT 78.600 508.400 79.400 508.600 ;
        RECT 86.000 508.400 86.600 509.600 ;
        RECT 87.600 509.200 91.400 509.800 ;
        RECT 87.600 509.000 88.400 509.200 ;
        RECT 49.200 507.800 50.200 508.200 ;
        RECT 40.400 507.200 41.200 507.600 ;
        RECT 35.000 506.600 38.800 507.200 ;
        RECT 35.000 506.400 35.800 506.600 ;
        RECT 23.600 504.200 24.400 505.000 ;
        RECT 25.200 504.800 26.000 506.400 ;
        RECT 27.000 505.400 27.800 505.600 ;
        RECT 27.000 504.800 29.800 505.400 ;
        RECT 29.200 504.200 29.800 504.800 ;
        RECT 33.200 504.200 34.000 505.000 ;
        RECT 23.600 503.600 25.600 504.200 ;
        RECT 24.800 502.200 25.600 503.600 ;
        RECT 29.200 502.200 30.000 504.200 ;
        RECT 33.200 503.600 34.600 504.200 ;
        RECT 33.400 502.200 34.600 503.600 ;
        RECT 38.000 502.200 38.800 506.600 ;
        RECT 39.800 506.200 43.400 506.600 ;
        RECT 44.400 506.200 45.000 507.600 ;
        RECT 46.000 507.200 50.200 507.800 ;
        RECT 51.200 507.600 53.200 508.400 ;
        RECT 55.600 507.600 58.200 508.400 ;
        RECT 60.400 508.300 61.200 508.400 ;
        RECT 62.000 508.300 62.800 508.400 ;
        RECT 60.400 508.200 62.800 508.300 ;
        RECT 59.600 507.700 63.600 508.200 ;
        RECT 59.600 507.600 61.200 507.700 ;
        RECT 62.000 507.600 63.600 507.700 ;
        RECT 65.000 507.600 67.600 508.400 ;
        RECT 68.400 507.600 71.000 508.400 ;
        RECT 73.200 508.200 74.000 508.400 ;
        RECT 72.400 507.600 74.000 508.200 ;
        RECT 75.600 507.800 86.600 508.400 ;
        RECT 75.600 507.600 77.200 507.800 ;
        RECT 39.600 506.000 43.600 506.200 ;
        RECT 39.600 502.200 40.400 506.000 ;
        RECT 42.800 502.200 43.600 506.000 ;
        RECT 44.400 502.200 45.200 506.200 ;
        RECT 46.000 505.000 46.600 507.200 ;
        RECT 51.200 507.000 51.800 507.600 ;
        RECT 51.000 506.600 51.800 507.000 ;
        RECT 50.200 506.400 51.800 506.600 ;
        RECT 49.200 506.000 51.800 506.400 ;
        RECT 55.800 506.200 56.400 507.600 ;
        RECT 59.600 507.200 60.400 507.600 ;
        RECT 62.800 507.200 63.600 507.600 ;
        RECT 57.400 506.200 61.000 506.600 ;
        RECT 62.200 506.200 65.800 506.600 ;
        RECT 66.800 506.200 67.400 507.600 ;
        RECT 68.600 506.200 69.200 507.600 ;
        RECT 72.400 507.200 73.200 507.600 ;
        RECT 70.200 506.200 73.800 506.600 ;
        RECT 49.200 505.600 51.000 506.000 ;
        RECT 46.000 503.000 46.800 505.000 ;
        RECT 50.200 503.000 51.000 505.600 ;
        RECT 55.600 502.200 56.400 506.200 ;
        RECT 57.200 506.000 61.200 506.200 ;
        RECT 57.200 502.200 58.000 506.000 ;
        RECT 60.400 502.200 61.200 506.000 ;
        RECT 62.000 506.000 66.000 506.200 ;
        RECT 62.000 502.200 62.800 506.000 ;
        RECT 65.200 502.200 66.000 506.000 ;
        RECT 66.800 502.200 67.600 506.200 ;
        RECT 68.400 502.200 69.200 506.200 ;
        RECT 70.000 506.000 74.000 506.200 ;
        RECT 70.000 502.200 70.800 506.000 ;
        RECT 73.200 502.200 74.000 506.000 ;
        RECT 74.800 502.200 75.600 507.000 ;
        RECT 79.800 505.600 80.400 507.800 ;
        RECT 85.400 507.600 86.200 507.800 ;
        RECT 92.400 507.200 93.200 510.600 ;
        RECT 105.200 510.400 105.800 511.600 ;
        RECT 111.600 511.200 112.400 519.800 ;
        RECT 108.200 510.600 112.400 511.200 ;
        RECT 108.200 510.400 109.000 510.600 ;
        RECT 100.400 510.200 101.200 510.400 ;
        RECT 96.200 509.600 101.200 510.200 ;
        RECT 105.200 509.600 106.000 510.400 ;
        RECT 109.800 509.800 110.600 510.000 ;
        RECT 96.200 509.400 97.000 509.600 ;
        RECT 97.800 508.400 98.600 508.600 ;
        RECT 105.200 508.400 105.800 509.600 ;
        RECT 106.800 509.200 110.600 509.800 ;
        RECT 106.800 509.000 107.600 509.200 ;
        RECT 94.800 507.800 105.800 508.400 ;
        RECT 94.800 507.600 96.400 507.800 ;
        RECT 89.400 506.600 93.200 507.200 ;
        RECT 89.400 506.400 90.200 506.600 ;
        RECT 78.000 504.200 78.800 505.000 ;
        RECT 79.600 504.800 80.400 505.600 ;
        RECT 81.400 505.400 82.200 505.600 ;
        RECT 81.400 504.800 84.200 505.400 ;
        RECT 83.600 504.200 84.200 504.800 ;
        RECT 87.600 504.200 88.400 505.000 ;
        RECT 78.000 503.600 80.000 504.200 ;
        RECT 79.200 502.200 80.000 503.600 ;
        RECT 83.600 502.200 84.400 504.200 ;
        RECT 87.600 503.600 89.000 504.200 ;
        RECT 87.800 502.200 89.000 503.600 ;
        RECT 92.400 502.200 93.200 506.600 ;
        RECT 94.000 502.200 94.800 507.000 ;
        RECT 99.000 505.600 99.600 507.800 ;
        RECT 104.600 507.600 105.400 507.800 ;
        RECT 111.600 507.200 112.400 510.600 ;
        RECT 108.600 506.600 112.400 507.200 ;
        RECT 108.600 506.400 109.400 506.600 ;
        RECT 97.200 504.200 98.000 505.000 ;
        RECT 98.800 504.800 99.600 505.600 ;
        RECT 100.600 505.400 101.400 505.600 ;
        RECT 100.600 504.800 103.400 505.400 ;
        RECT 102.800 504.200 103.400 504.800 ;
        RECT 106.800 504.200 107.600 505.000 ;
        RECT 97.200 503.600 99.200 504.200 ;
        RECT 98.400 502.200 99.200 503.600 ;
        RECT 102.800 502.200 103.600 504.200 ;
        RECT 106.800 503.600 108.200 504.200 ;
        RECT 107.000 502.200 108.200 503.600 ;
        RECT 111.600 502.200 112.400 506.600 ;
        RECT 113.200 502.200 114.000 519.800 ;
        RECT 114.800 504.800 115.600 506.400 ;
        RECT 116.400 504.800 117.200 506.400 ;
        RECT 118.000 502.200 118.800 519.800 ;
        RECT 123.400 518.400 124.200 519.800 ;
        RECT 122.800 517.600 124.200 518.400 ;
        RECT 123.400 512.800 124.200 517.600 ;
        RECT 127.600 515.000 128.400 519.000 ;
        RECT 122.600 512.200 124.200 512.800 ;
        RECT 121.200 509.600 122.000 511.200 ;
        RECT 122.600 508.400 123.200 512.200 ;
        RECT 127.800 511.600 128.400 515.000 ;
        RECT 124.600 511.000 128.400 511.600 ;
        RECT 129.200 515.000 130.000 519.000 ;
        RECT 133.400 518.400 134.200 519.800 ;
        RECT 132.400 517.600 134.200 518.400 ;
        RECT 129.200 511.600 129.800 515.000 ;
        RECT 133.400 512.800 134.200 517.600 ;
        RECT 133.400 512.200 135.000 512.800 ;
        RECT 141.400 512.600 142.200 519.800 ;
        RECT 129.200 511.000 133.000 511.600 ;
        RECT 124.600 509.000 125.200 511.000 ;
        RECT 121.200 507.600 123.200 508.400 ;
        RECT 123.800 508.200 125.200 509.000 ;
        RECT 126.000 508.800 126.800 510.400 ;
        RECT 127.600 510.300 128.400 510.400 ;
        RECT 129.200 510.300 130.000 510.400 ;
        RECT 127.600 509.700 130.000 510.300 ;
        RECT 127.600 508.800 128.400 509.700 ;
        RECT 129.200 508.800 130.000 509.700 ;
        RECT 130.800 508.800 131.600 510.400 ;
        RECT 132.400 509.000 133.000 511.000 ;
        RECT 122.600 507.000 123.200 507.600 ;
        RECT 124.200 507.800 125.200 508.200 ;
        RECT 132.400 508.200 133.800 509.000 ;
        RECT 134.400 508.400 135.000 512.200 ;
        RECT 140.400 511.800 142.200 512.600 ;
        RECT 135.600 510.300 136.400 511.200 ;
        RECT 137.200 510.300 138.000 510.400 ;
        RECT 135.600 509.700 138.000 510.300 ;
        RECT 135.600 509.600 136.400 509.700 ;
        RECT 137.200 509.600 138.000 509.700 ;
        RECT 140.600 508.400 141.200 511.800 ;
        RECT 142.000 509.600 142.800 511.200 ;
        RECT 132.400 507.800 133.400 508.200 ;
        RECT 124.200 507.200 128.400 507.800 ;
        RECT 122.600 506.600 123.400 507.000 ;
        RECT 122.600 506.000 124.200 506.600 ;
        RECT 123.400 503.000 124.200 506.000 ;
        RECT 127.800 505.000 128.400 507.200 ;
        RECT 127.600 503.000 128.400 505.000 ;
        RECT 129.200 507.200 133.400 507.800 ;
        RECT 134.400 507.600 136.400 508.400 ;
        RECT 140.400 507.600 141.200 508.400 ;
        RECT 129.200 505.000 129.800 507.200 ;
        RECT 134.400 507.000 135.000 507.600 ;
        RECT 134.200 506.600 135.000 507.000 ;
        RECT 133.400 506.000 135.000 506.600 ;
        RECT 129.200 503.000 130.000 505.000 ;
        RECT 133.400 503.000 134.200 506.000 ;
        RECT 138.800 504.800 139.600 506.400 ;
        RECT 140.600 504.400 141.200 507.600 ;
        RECT 142.000 506.300 142.800 506.400 ;
        RECT 143.600 506.300 144.400 506.400 ;
        RECT 142.000 505.700 144.400 506.300 ;
        RECT 142.000 505.600 142.800 505.700 ;
        RECT 143.600 504.800 144.400 505.700 ;
        RECT 140.400 502.200 141.200 504.400 ;
        RECT 145.200 504.300 146.000 519.800 ;
        RECT 153.200 511.200 154.000 519.800 ;
        RECT 156.400 511.200 157.200 519.800 ;
        RECT 159.600 511.200 160.400 519.800 ;
        RECT 162.800 511.200 163.600 519.800 ;
        RECT 151.600 510.400 154.000 511.200 ;
        RECT 155.000 510.400 157.200 511.200 ;
        RECT 158.200 510.400 160.400 511.200 ;
        RECT 161.800 510.400 163.600 511.200 ;
        RECT 151.600 507.600 152.400 510.400 ;
        RECT 155.000 509.000 155.800 510.400 ;
        RECT 158.200 509.000 159.000 510.400 ;
        RECT 161.800 509.000 162.600 510.400 ;
        RECT 153.200 508.200 155.800 509.000 ;
        RECT 156.600 508.200 159.000 509.000 ;
        RECT 160.000 508.200 162.600 509.000 ;
        RECT 163.400 508.200 165.200 509.000 ;
        RECT 155.000 507.600 155.800 508.200 ;
        RECT 158.200 507.600 159.000 508.200 ;
        RECT 161.800 507.600 162.600 508.200 ;
        RECT 164.400 507.600 165.200 508.200 ;
        RECT 151.600 506.800 154.000 507.600 ;
        RECT 155.000 506.800 157.200 507.600 ;
        RECT 158.200 506.800 160.400 507.600 ;
        RECT 161.800 506.800 163.600 507.600 ;
        RECT 150.000 504.300 150.800 504.400 ;
        RECT 145.200 503.700 150.800 504.300 ;
        RECT 145.200 502.200 146.000 503.700 ;
        RECT 150.000 503.600 150.800 503.700 ;
        RECT 153.200 502.200 154.000 506.800 ;
        RECT 156.400 502.200 157.200 506.800 ;
        RECT 159.600 502.200 160.400 506.800 ;
        RECT 162.800 502.200 163.600 506.800 ;
        RECT 166.000 504.800 166.800 506.400 ;
        RECT 167.600 502.200 168.400 519.800 ;
        RECT 171.800 512.600 172.600 519.800 ;
        RECT 170.800 511.800 172.600 512.600 ;
        RECT 174.000 512.400 174.800 519.800 ;
        RECT 175.600 512.400 176.400 512.600 ;
        RECT 178.400 512.400 180.000 519.800 ;
        RECT 174.000 511.800 176.400 512.400 ;
        RECT 178.000 511.800 180.000 512.400 ;
        RECT 182.200 512.400 183.000 512.600 ;
        RECT 183.600 512.400 184.400 519.800 ;
        RECT 182.200 511.800 184.400 512.400 ;
        RECT 171.000 510.400 171.600 511.800 ;
        RECT 170.800 509.600 171.600 510.400 ;
        RECT 172.400 509.600 173.200 511.200 ;
        RECT 178.000 510.400 178.600 511.800 ;
        RECT 182.200 511.200 182.800 511.800 ;
        RECT 179.400 510.600 182.800 511.200 ;
        RECT 186.800 511.200 187.600 519.800 ;
        RECT 190.000 511.200 190.800 519.800 ;
        RECT 193.200 511.200 194.000 519.800 ;
        RECT 196.400 511.200 197.200 519.800 ;
        RECT 201.200 516.400 202.000 519.800 ;
        RECT 201.000 515.800 202.000 516.400 ;
        RECT 201.000 515.200 201.600 515.800 ;
        RECT 204.400 515.200 205.200 519.800 ;
        RECT 207.600 517.000 208.400 519.800 ;
        RECT 209.200 517.000 210.000 519.800 ;
        RECT 199.600 514.600 201.600 515.200 ;
        RECT 179.400 510.400 180.200 510.600 ;
        RECT 186.800 510.400 188.600 511.200 ;
        RECT 190.000 510.400 192.200 511.200 ;
        RECT 193.200 510.400 195.400 511.200 ;
        RECT 196.400 510.400 198.800 511.200 ;
        RECT 177.200 509.800 178.600 510.400 ;
        RECT 181.600 509.800 182.400 510.000 ;
        RECT 177.200 509.600 179.000 509.800 ;
        RECT 171.000 508.400 171.600 509.600 ;
        RECT 178.000 509.200 179.000 509.600 ;
        RECT 170.800 507.600 171.600 508.400 ;
        RECT 174.000 507.600 175.600 508.400 ;
        RECT 176.800 507.600 177.600 508.400 ;
        RECT 169.200 504.800 170.000 506.400 ;
        RECT 171.000 504.200 171.600 507.600 ;
        RECT 177.000 507.200 177.600 507.600 ;
        RECT 175.600 506.800 176.400 507.000 ;
        RECT 170.800 502.200 171.600 504.200 ;
        RECT 174.000 506.200 176.400 506.800 ;
        RECT 177.000 506.400 177.800 507.200 ;
        RECT 174.000 502.200 174.800 506.200 ;
        RECT 178.400 505.800 179.000 509.200 ;
        RECT 179.800 509.200 182.400 509.800 ;
        RECT 179.800 508.600 180.400 509.200 ;
        RECT 187.800 509.000 188.600 510.400 ;
        RECT 191.400 509.000 192.200 510.400 ;
        RECT 194.600 509.000 195.400 510.400 ;
        RECT 179.600 507.800 180.400 508.600 ;
        RECT 182.800 508.200 184.400 508.400 ;
        RECT 181.000 507.600 184.400 508.200 ;
        RECT 185.200 508.200 187.000 509.000 ;
        RECT 187.800 508.200 190.400 509.000 ;
        RECT 191.400 508.200 193.800 509.000 ;
        RECT 194.600 508.200 197.200 509.000 ;
        RECT 185.200 507.600 186.000 508.200 ;
        RECT 187.800 507.600 188.600 508.200 ;
        RECT 191.400 507.600 192.200 508.200 ;
        RECT 194.600 507.600 195.400 508.200 ;
        RECT 198.000 507.600 198.800 510.400 ;
        RECT 181.000 507.200 181.600 507.600 ;
        RECT 179.600 506.600 181.600 507.200 ;
        RECT 182.200 506.800 183.000 507.000 ;
        RECT 186.800 506.800 188.600 507.600 ;
        RECT 190.000 506.800 192.200 507.600 ;
        RECT 193.200 506.800 195.400 507.600 ;
        RECT 196.400 506.800 198.800 507.600 ;
        RECT 199.600 509.000 200.400 514.600 ;
        RECT 202.200 514.400 206.400 515.200 ;
        RECT 210.800 515.000 211.600 519.800 ;
        RECT 214.000 515.000 214.800 519.800 ;
        RECT 202.200 514.000 202.800 514.400 ;
        RECT 201.200 513.200 202.800 514.000 ;
        RECT 205.800 513.800 211.600 514.400 ;
        RECT 203.800 513.200 205.200 513.800 ;
        RECT 203.800 513.000 210.000 513.200 ;
        RECT 204.600 512.600 210.000 513.000 ;
        RECT 209.200 512.400 210.000 512.600 ;
        RECT 211.000 513.000 211.600 513.800 ;
        RECT 212.200 513.600 214.800 514.400 ;
        RECT 217.200 513.600 218.000 519.800 ;
        RECT 218.800 517.000 219.600 519.800 ;
        RECT 220.400 517.000 221.200 519.800 ;
        RECT 222.000 517.000 222.800 519.800 ;
        RECT 220.400 514.400 224.600 515.200 ;
        RECT 225.200 514.400 226.000 519.800 ;
        RECT 228.400 515.200 229.200 519.800 ;
        RECT 228.400 514.600 231.000 515.200 ;
        RECT 225.200 513.600 227.800 514.400 ;
        RECT 218.800 513.000 219.600 513.200 ;
        RECT 211.000 512.400 219.600 513.000 ;
        RECT 222.000 513.000 222.800 513.200 ;
        RECT 230.400 513.000 231.000 514.600 ;
        RECT 222.000 512.400 231.000 513.000 ;
        RECT 230.400 510.600 231.000 512.400 ;
        RECT 231.600 512.000 232.400 519.800 ;
        RECT 233.200 514.300 234.000 514.400 ;
        RECT 235.600 514.300 236.400 514.400 ;
        RECT 233.200 513.700 236.400 514.300 ;
        RECT 233.200 513.600 234.000 513.700 ;
        RECT 235.600 513.600 236.400 513.700 ;
        RECT 235.600 512.400 236.200 513.600 ;
        RECT 237.000 512.400 237.800 519.800 ;
        RECT 231.600 511.200 232.600 512.000 ;
        RECT 234.800 511.800 236.200 512.400 ;
        RECT 236.800 511.800 237.800 512.400 ;
        RECT 234.800 511.600 235.600 511.800 ;
        RECT 201.000 510.000 224.400 510.600 ;
        RECT 230.400 510.000 231.200 510.600 ;
        RECT 201.000 509.800 201.800 510.000 ;
        RECT 204.400 509.600 205.200 510.000 ;
        RECT 206.000 509.600 206.800 510.000 ;
        RECT 223.600 509.400 224.400 510.000 ;
        RECT 199.600 508.200 208.400 509.000 ;
        RECT 209.000 508.600 211.000 509.400 ;
        RECT 214.800 508.600 218.000 509.400 ;
        RECT 179.600 506.400 181.200 506.600 ;
        RECT 182.200 506.200 184.400 506.800 ;
        RECT 178.400 504.400 180.000 505.800 ;
        RECT 177.200 503.600 180.000 504.400 ;
        RECT 178.400 502.200 180.000 503.600 ;
        RECT 183.600 502.200 184.400 506.200 ;
        RECT 186.800 502.200 187.600 506.800 ;
        RECT 190.000 502.200 190.800 506.800 ;
        RECT 193.200 502.200 194.000 506.800 ;
        RECT 196.400 502.200 197.200 506.800 ;
        RECT 199.600 502.200 200.400 508.200 ;
        RECT 202.000 506.800 205.000 507.600 ;
        RECT 204.200 506.200 205.000 506.800 ;
        RECT 210.200 506.200 211.000 508.600 ;
        RECT 212.400 506.800 213.200 508.400 ;
        RECT 217.600 507.800 218.400 508.000 ;
        RECT 214.000 507.200 218.400 507.800 ;
        RECT 214.000 507.000 214.800 507.200 ;
        RECT 220.400 506.400 221.200 509.200 ;
        RECT 226.200 508.600 230.000 509.400 ;
        RECT 226.200 507.400 227.000 508.600 ;
        RECT 230.600 508.000 231.200 510.000 ;
        RECT 214.000 506.200 214.800 506.400 ;
        RECT 204.200 505.400 206.800 506.200 ;
        RECT 210.200 505.600 214.800 506.200 ;
        RECT 215.600 505.600 217.200 506.400 ;
        RECT 220.200 505.600 221.200 506.400 ;
        RECT 225.200 506.800 227.000 507.400 ;
        RECT 230.000 507.400 231.200 508.000 ;
        RECT 225.200 506.200 226.000 506.800 ;
        RECT 206.000 502.200 206.800 505.400 ;
        RECT 223.600 505.400 226.000 506.200 ;
        RECT 207.600 502.200 208.400 505.000 ;
        RECT 209.200 502.200 210.000 505.000 ;
        RECT 210.800 502.200 211.600 505.000 ;
        RECT 214.000 502.200 214.800 505.000 ;
        RECT 217.200 502.200 218.000 505.000 ;
        RECT 218.800 502.200 219.600 505.000 ;
        RECT 220.400 502.200 221.200 505.000 ;
        RECT 222.000 502.200 222.800 505.000 ;
        RECT 223.600 502.200 224.400 505.400 ;
        RECT 230.000 502.200 230.800 507.400 ;
        RECT 231.800 506.800 232.600 511.200 ;
        RECT 236.800 510.400 237.400 511.800 ;
        RECT 236.400 509.600 237.400 510.400 ;
        RECT 236.800 508.400 237.400 509.600 ;
        RECT 238.000 508.800 238.800 510.400 ;
        RECT 234.800 507.600 237.400 508.400 ;
        RECT 239.600 508.200 240.400 508.400 ;
        RECT 238.800 507.600 240.400 508.200 ;
        RECT 231.600 506.000 232.600 506.800 ;
        RECT 235.000 506.200 235.600 507.600 ;
        RECT 238.800 507.200 239.600 507.600 ;
        RECT 241.200 506.800 242.000 508.400 ;
        RECT 236.600 506.200 240.200 506.600 ;
        RECT 242.800 506.200 243.600 519.800 ;
        RECT 244.400 511.600 245.200 513.200 ;
        RECT 231.600 502.200 232.400 506.000 ;
        RECT 234.800 502.200 235.600 506.200 ;
        RECT 236.400 506.000 240.400 506.200 ;
        RECT 236.400 502.200 237.200 506.000 ;
        RECT 239.600 502.200 240.400 506.000 ;
        RECT 242.800 505.600 244.600 506.200 ;
        RECT 243.800 502.200 244.600 505.600 ;
        RECT 246.000 504.800 246.800 506.400 ;
        RECT 247.600 502.200 248.400 519.800 ;
        RECT 250.800 516.400 251.600 519.800 ;
        RECT 250.600 515.800 251.600 516.400 ;
        RECT 250.600 515.200 251.200 515.800 ;
        RECT 254.000 515.200 254.800 519.800 ;
        RECT 257.200 517.000 258.000 519.800 ;
        RECT 258.800 517.000 259.600 519.800 ;
        RECT 249.200 514.600 251.200 515.200 ;
        RECT 249.200 509.000 250.000 514.600 ;
        RECT 251.800 514.400 256.000 515.200 ;
        RECT 260.400 515.000 261.200 519.800 ;
        RECT 263.600 515.000 264.400 519.800 ;
        RECT 251.800 514.000 252.400 514.400 ;
        RECT 250.800 513.200 252.400 514.000 ;
        RECT 255.400 513.800 261.200 514.400 ;
        RECT 253.400 513.200 254.800 513.800 ;
        RECT 253.400 513.000 259.600 513.200 ;
        RECT 254.200 512.600 259.600 513.000 ;
        RECT 258.800 512.400 259.600 512.600 ;
        RECT 260.600 513.000 261.200 513.800 ;
        RECT 261.800 513.600 264.400 514.400 ;
        RECT 266.800 513.600 267.600 519.800 ;
        RECT 268.400 517.000 269.200 519.800 ;
        RECT 270.000 517.000 270.800 519.800 ;
        RECT 271.600 517.000 272.400 519.800 ;
        RECT 270.000 514.400 274.200 515.200 ;
        RECT 274.800 514.400 275.600 519.800 ;
        RECT 278.000 515.200 278.800 519.800 ;
        RECT 278.000 514.600 280.600 515.200 ;
        RECT 274.800 513.600 277.400 514.400 ;
        RECT 268.400 513.000 269.200 513.200 ;
        RECT 260.600 512.400 269.200 513.000 ;
        RECT 271.600 513.000 272.400 513.200 ;
        RECT 280.000 513.000 280.600 514.600 ;
        RECT 271.600 512.400 280.600 513.000 ;
        RECT 280.000 510.600 280.600 512.400 ;
        RECT 281.200 512.000 282.000 519.800 ;
        RECT 286.000 516.400 286.800 519.800 ;
        RECT 285.800 515.800 286.800 516.400 ;
        RECT 285.800 515.200 286.400 515.800 ;
        RECT 289.200 515.200 290.000 519.800 ;
        RECT 292.400 517.000 293.200 519.800 ;
        RECT 294.000 517.000 294.800 519.800 ;
        RECT 284.400 514.600 286.400 515.200 ;
        RECT 281.200 511.200 282.200 512.000 ;
        RECT 250.600 510.000 274.000 510.600 ;
        RECT 280.000 510.000 280.800 510.600 ;
        RECT 250.600 509.800 251.400 510.000 ;
        RECT 254.000 509.600 254.800 510.000 ;
        RECT 255.600 509.600 256.400 510.000 ;
        RECT 262.000 509.600 262.800 510.000 ;
        RECT 273.200 509.400 274.000 510.000 ;
        RECT 249.200 508.200 258.000 509.000 ;
        RECT 258.600 508.600 260.600 509.400 ;
        RECT 264.400 508.600 267.600 509.400 ;
        RECT 249.200 502.200 250.000 508.200 ;
        RECT 251.600 506.800 254.600 507.600 ;
        RECT 253.800 506.200 254.600 506.800 ;
        RECT 259.800 506.200 260.600 508.600 ;
        RECT 262.000 506.800 262.800 508.400 ;
        RECT 267.200 507.800 268.000 508.000 ;
        RECT 263.600 507.200 268.000 507.800 ;
        RECT 263.600 507.000 264.400 507.200 ;
        RECT 270.000 506.400 270.800 509.200 ;
        RECT 275.800 508.600 279.600 509.400 ;
        RECT 275.800 507.400 276.600 508.600 ;
        RECT 280.200 508.000 280.800 510.000 ;
        RECT 263.600 506.200 264.400 506.400 ;
        RECT 253.800 505.400 256.400 506.200 ;
        RECT 259.800 505.600 264.400 506.200 ;
        RECT 265.200 505.600 266.800 506.400 ;
        RECT 269.800 505.600 270.800 506.400 ;
        RECT 274.800 506.800 276.600 507.400 ;
        RECT 279.600 507.400 280.800 508.000 ;
        RECT 274.800 506.200 275.600 506.800 ;
        RECT 255.600 502.200 256.400 505.400 ;
        RECT 273.200 505.400 275.600 506.200 ;
        RECT 257.200 502.200 258.000 505.000 ;
        RECT 258.800 502.200 259.600 505.000 ;
        RECT 260.400 502.200 261.200 505.000 ;
        RECT 263.600 502.200 264.400 505.000 ;
        RECT 266.800 502.200 267.600 505.000 ;
        RECT 268.400 502.200 269.200 505.000 ;
        RECT 270.000 502.200 270.800 505.000 ;
        RECT 271.600 502.200 272.400 505.000 ;
        RECT 273.200 502.200 274.000 505.400 ;
        RECT 279.600 502.200 280.400 507.400 ;
        RECT 281.400 506.800 282.200 511.200 ;
        RECT 281.200 506.000 282.200 506.800 ;
        RECT 284.400 509.000 285.200 514.600 ;
        RECT 287.000 514.400 291.200 515.200 ;
        RECT 295.600 515.000 296.400 519.800 ;
        RECT 298.800 515.000 299.600 519.800 ;
        RECT 287.000 514.000 287.600 514.400 ;
        RECT 286.000 513.200 287.600 514.000 ;
        RECT 290.600 513.800 296.400 514.400 ;
        RECT 288.600 513.200 290.000 513.800 ;
        RECT 288.600 513.000 294.800 513.200 ;
        RECT 289.400 512.600 294.800 513.000 ;
        RECT 294.000 512.400 294.800 512.600 ;
        RECT 295.800 513.000 296.400 513.800 ;
        RECT 297.000 513.600 299.600 514.400 ;
        RECT 302.000 513.600 302.800 519.800 ;
        RECT 303.600 517.000 304.400 519.800 ;
        RECT 305.200 517.000 306.000 519.800 ;
        RECT 306.800 517.000 307.600 519.800 ;
        RECT 305.200 514.400 309.400 515.200 ;
        RECT 310.000 514.400 310.800 519.800 ;
        RECT 313.200 515.200 314.000 519.800 ;
        RECT 313.200 514.600 315.800 515.200 ;
        RECT 310.000 513.600 312.600 514.400 ;
        RECT 303.600 513.000 304.400 513.200 ;
        RECT 295.800 512.400 304.400 513.000 ;
        RECT 306.800 513.000 307.600 513.200 ;
        RECT 315.200 513.000 315.800 514.600 ;
        RECT 306.800 512.400 315.800 513.000 ;
        RECT 315.200 510.600 315.800 512.400 ;
        RECT 316.400 512.000 317.200 519.800 ;
        RECT 318.000 514.300 318.800 514.400 ;
        RECT 318.000 513.700 325.200 514.300 ;
        RECT 318.000 513.600 318.800 513.700 ;
        RECT 316.400 511.200 317.400 512.000 ;
        RECT 324.400 511.600 325.200 513.700 ;
        RECT 285.800 510.000 309.200 510.600 ;
        RECT 315.200 510.000 316.000 510.600 ;
        RECT 285.800 509.800 286.600 510.000 ;
        RECT 287.600 509.600 288.400 510.000 ;
        RECT 290.800 509.600 291.600 510.000 ;
        RECT 308.400 509.400 309.200 510.000 ;
        RECT 284.400 508.200 293.200 509.000 ;
        RECT 293.800 508.600 295.800 509.400 ;
        RECT 299.600 508.600 302.800 509.400 ;
        RECT 281.200 502.200 282.000 506.000 ;
        RECT 284.400 502.200 285.200 508.200 ;
        RECT 286.800 506.800 289.800 507.600 ;
        RECT 289.000 506.200 289.800 506.800 ;
        RECT 295.000 506.200 295.800 508.600 ;
        RECT 297.200 506.800 298.000 508.400 ;
        RECT 302.400 507.800 303.200 508.000 ;
        RECT 298.800 507.200 303.200 507.800 ;
        RECT 298.800 507.000 299.600 507.200 ;
        RECT 305.200 506.400 306.000 509.200 ;
        RECT 311.000 508.600 314.800 509.400 ;
        RECT 311.000 507.400 311.800 508.600 ;
        RECT 315.400 508.000 316.000 510.000 ;
        RECT 298.800 506.200 299.600 506.400 ;
        RECT 289.000 505.400 291.600 506.200 ;
        RECT 295.000 505.600 299.600 506.200 ;
        RECT 300.400 505.600 302.000 506.400 ;
        RECT 305.000 505.600 306.000 506.400 ;
        RECT 310.000 506.800 311.800 507.400 ;
        RECT 314.800 507.400 316.000 508.000 ;
        RECT 310.000 506.200 310.800 506.800 ;
        RECT 290.800 502.200 291.600 505.400 ;
        RECT 308.400 505.400 310.800 506.200 ;
        RECT 292.400 502.200 293.200 505.000 ;
        RECT 294.000 502.200 294.800 505.000 ;
        RECT 295.600 502.200 296.400 505.000 ;
        RECT 298.800 502.200 299.600 505.000 ;
        RECT 302.000 502.200 302.800 505.000 ;
        RECT 303.600 502.200 304.400 505.000 ;
        RECT 305.200 502.200 306.000 505.000 ;
        RECT 306.800 502.200 307.600 505.000 ;
        RECT 308.400 502.200 309.200 505.400 ;
        RECT 314.800 502.200 315.600 507.400 ;
        RECT 316.600 506.800 317.400 511.200 ;
        RECT 316.400 506.000 317.400 506.800 ;
        RECT 326.000 506.200 326.800 519.800 ;
        RECT 329.200 511.600 330.000 514.400 ;
        RECT 327.600 506.800 328.400 508.400 ;
        RECT 330.800 506.200 331.600 519.800 ;
        RECT 334.000 511.400 334.800 519.800 ;
        RECT 338.400 516.400 339.200 519.800 ;
        RECT 337.200 515.800 339.200 516.400 ;
        RECT 342.800 515.800 343.600 519.800 ;
        RECT 347.000 515.800 348.200 519.800 ;
        RECT 337.200 515.000 338.000 515.800 ;
        RECT 342.800 515.200 343.400 515.800 ;
        RECT 340.600 514.600 344.200 515.200 ;
        RECT 346.800 515.000 347.600 515.800 ;
        RECT 340.600 514.400 341.400 514.600 ;
        RECT 343.400 514.400 344.200 514.600 ;
        RECT 337.200 513.000 338.000 513.200 ;
        RECT 341.800 513.000 342.600 513.200 ;
        RECT 337.200 512.400 342.600 513.000 ;
        RECT 343.200 513.000 345.400 513.600 ;
        RECT 343.200 511.800 343.800 513.000 ;
        RECT 344.600 512.800 345.400 513.000 ;
        RECT 347.000 513.200 348.400 514.000 ;
        RECT 347.000 512.200 347.600 513.200 ;
        RECT 339.000 511.400 343.800 511.800 ;
        RECT 334.000 511.200 343.800 511.400 ;
        RECT 345.200 511.600 347.600 512.200 ;
        RECT 334.000 511.000 339.800 511.200 ;
        RECT 334.000 510.800 339.600 511.000 ;
        RECT 340.400 510.200 341.200 510.400 ;
        RECT 336.200 509.600 341.200 510.200 ;
        RECT 336.200 509.400 337.000 509.600 ;
        RECT 338.800 509.400 339.600 509.600 ;
        RECT 337.800 508.400 338.600 508.600 ;
        RECT 345.200 508.400 345.800 511.600 ;
        RECT 351.600 511.200 352.400 519.800 ;
        RECT 348.200 510.600 352.400 511.200 ;
        RECT 348.200 510.400 349.000 510.600 ;
        RECT 349.800 509.800 350.600 510.000 ;
        RECT 346.800 509.200 350.600 509.800 ;
        RECT 346.800 509.000 347.600 509.200 ;
        RECT 332.400 506.800 333.200 508.400 ;
        RECT 334.800 507.800 345.800 508.400 ;
        RECT 334.800 507.600 336.400 507.800 ;
        RECT 316.400 502.200 317.200 506.000 ;
        RECT 325.000 505.600 326.800 506.200 ;
        RECT 329.800 505.600 331.600 506.200 ;
        RECT 319.600 504.300 320.400 504.400 ;
        RECT 325.000 504.300 325.800 505.600 ;
        RECT 319.600 503.700 325.800 504.300 ;
        RECT 319.600 503.600 320.400 503.700 ;
        RECT 325.000 502.200 325.800 503.700 ;
        RECT 329.800 504.400 330.600 505.600 ;
        RECT 329.800 503.600 331.600 504.400 ;
        RECT 329.800 502.200 330.600 503.600 ;
        RECT 334.000 502.200 334.800 507.000 ;
        RECT 339.000 505.600 339.600 507.800 ;
        RECT 344.600 507.600 345.400 507.800 ;
        RECT 351.600 507.200 352.400 510.600 ;
        RECT 348.600 506.600 352.400 507.200 ;
        RECT 353.200 506.800 354.000 508.400 ;
        RECT 348.600 506.400 349.400 506.600 ;
        RECT 337.200 504.200 338.000 505.000 ;
        RECT 338.800 504.800 339.600 505.600 ;
        RECT 340.600 505.400 341.400 505.600 ;
        RECT 340.600 504.800 343.400 505.400 ;
        RECT 342.800 504.200 343.400 504.800 ;
        RECT 346.800 504.200 347.600 505.000 ;
        RECT 337.200 503.600 339.200 504.200 ;
        RECT 338.400 502.200 339.200 503.600 ;
        RECT 342.800 502.200 343.600 504.200 ;
        RECT 346.800 503.600 348.200 504.200 ;
        RECT 347.000 502.200 348.200 503.600 ;
        RECT 351.600 502.200 352.400 506.600 ;
        RECT 354.800 506.200 355.600 519.800 ;
        RECT 356.400 511.600 357.200 514.400 ;
        RECT 358.000 511.400 358.800 519.800 ;
        RECT 362.400 516.400 363.200 519.800 ;
        RECT 361.200 515.800 363.200 516.400 ;
        RECT 366.800 515.800 367.600 519.800 ;
        RECT 371.000 515.800 372.200 519.800 ;
        RECT 361.200 515.000 362.000 515.800 ;
        RECT 366.800 515.200 367.400 515.800 ;
        RECT 364.600 514.600 368.200 515.200 ;
        RECT 370.800 515.000 371.600 515.800 ;
        RECT 364.600 514.400 365.400 514.600 ;
        RECT 367.400 514.400 368.200 514.600 ;
        RECT 371.800 514.000 373.200 514.400 ;
        RECT 371.000 513.600 373.200 514.000 ;
        RECT 361.200 513.000 362.000 513.200 ;
        RECT 365.800 513.000 366.600 513.200 ;
        RECT 361.200 512.400 366.600 513.000 ;
        RECT 367.200 513.000 369.400 513.600 ;
        RECT 367.200 511.800 367.800 513.000 ;
        RECT 368.600 512.800 369.400 513.000 ;
        RECT 371.000 513.200 372.400 513.600 ;
        RECT 371.000 512.200 371.600 513.200 ;
        RECT 363.000 511.400 367.800 511.800 ;
        RECT 358.000 511.200 367.800 511.400 ;
        RECT 369.200 511.600 371.600 512.200 ;
        RECT 358.000 511.000 363.800 511.200 ;
        RECT 358.000 510.800 363.600 511.000 ;
        RECT 364.400 510.200 365.200 510.400 ;
        RECT 360.200 509.600 365.200 510.200 ;
        RECT 367.600 510.300 368.400 510.400 ;
        RECT 369.200 510.300 369.800 511.600 ;
        RECT 375.600 511.200 376.400 519.800 ;
        RECT 372.200 510.600 376.400 511.200 ;
        RECT 377.200 515.000 378.000 519.000 ;
        RECT 377.200 511.600 377.800 515.000 ;
        RECT 381.400 512.800 382.200 519.800 ;
        RECT 381.400 512.200 383.000 512.800 ;
        RECT 377.200 511.000 381.000 511.600 ;
        RECT 372.200 510.400 373.000 510.600 ;
        RECT 367.600 509.700 369.900 510.300 ;
        RECT 373.800 509.800 374.600 510.000 ;
        RECT 367.600 509.600 368.400 509.700 ;
        RECT 360.200 509.400 361.000 509.600 ;
        RECT 361.800 508.400 362.600 508.600 ;
        RECT 369.200 508.400 369.800 509.700 ;
        RECT 370.800 509.200 374.600 509.800 ;
        RECT 370.800 509.000 371.600 509.200 ;
        RECT 358.800 507.800 369.800 508.400 ;
        RECT 358.800 507.600 360.400 507.800 ;
        RECT 354.800 505.600 356.600 506.200 ;
        RECT 355.800 504.400 356.600 505.600 ;
        RECT 354.800 503.600 356.600 504.400 ;
        RECT 355.800 502.200 356.600 503.600 ;
        RECT 358.000 502.200 358.800 507.000 ;
        RECT 363.000 505.600 363.600 507.800 ;
        RECT 368.600 507.600 369.400 507.800 ;
        RECT 375.600 507.200 376.400 510.600 ;
        RECT 377.200 508.800 378.000 510.400 ;
        RECT 378.800 508.800 379.600 510.400 ;
        RECT 380.400 509.000 381.000 511.000 ;
        RECT 380.400 508.200 381.800 509.000 ;
        RECT 382.400 508.400 383.000 512.200 ;
        RECT 389.400 512.400 390.200 519.800 ;
        RECT 390.800 513.600 391.600 514.400 ;
        RECT 391.000 512.400 391.600 513.600 ;
        RECT 389.400 511.800 390.400 512.400 ;
        RECT 391.000 511.800 392.400 512.400 ;
        RECT 383.600 509.600 384.400 511.200 ;
        RECT 389.800 510.400 390.400 511.800 ;
        RECT 391.600 511.600 392.400 511.800 ;
        RECT 393.200 511.600 394.000 514.400 ;
        RECT 388.400 510.300 389.200 510.400 ;
        RECT 385.300 509.700 389.200 510.300 ;
        RECT 382.400 508.300 384.400 508.400 ;
        RECT 385.300 508.300 385.900 509.700 ;
        RECT 388.400 508.800 389.200 509.700 ;
        RECT 389.800 509.600 390.800 510.400 ;
        RECT 389.800 508.400 390.400 509.600 ;
        RECT 380.400 507.800 381.400 508.200 ;
        RECT 372.600 506.600 376.400 507.200 ;
        RECT 372.600 506.400 373.400 506.600 ;
        RECT 361.200 504.200 362.000 505.000 ;
        RECT 362.800 504.800 363.600 505.600 ;
        RECT 364.600 505.400 365.400 505.600 ;
        RECT 364.600 504.800 367.400 505.400 ;
        RECT 366.800 504.200 367.400 504.800 ;
        RECT 370.800 504.200 371.600 505.000 ;
        RECT 361.200 503.600 363.200 504.200 ;
        RECT 362.400 502.200 363.200 503.600 ;
        RECT 366.800 502.200 367.600 504.200 ;
        RECT 370.800 503.600 372.200 504.200 ;
        RECT 371.000 502.200 372.200 503.600 ;
        RECT 375.600 502.200 376.400 506.600 ;
        RECT 377.200 507.200 381.400 507.800 ;
        RECT 382.400 507.700 385.900 508.300 ;
        RECT 386.800 508.200 387.600 508.400 ;
        RECT 382.400 507.600 384.400 507.700 ;
        RECT 386.800 507.600 388.400 508.200 ;
        RECT 389.800 507.600 392.400 508.400 ;
        RECT 377.200 505.000 377.800 507.200 ;
        RECT 382.400 507.000 383.000 507.600 ;
        RECT 387.600 507.200 388.400 507.600 ;
        RECT 382.200 506.600 383.000 507.000 ;
        RECT 381.400 506.000 383.000 506.600 ;
        RECT 387.000 506.200 390.600 506.600 ;
        RECT 391.600 506.200 392.200 507.600 ;
        RECT 394.800 506.200 395.600 519.800 ;
        RECT 398.800 513.600 399.600 514.400 ;
        RECT 398.800 512.400 399.400 513.600 ;
        RECT 400.200 512.400 401.000 519.800 ;
        RECT 406.000 512.800 406.800 519.800 ;
        RECT 398.000 511.800 399.400 512.400 ;
        RECT 400.000 511.800 401.000 512.400 ;
        RECT 405.800 511.800 406.800 512.800 ;
        RECT 409.200 512.400 410.000 519.800 ;
        RECT 407.400 511.800 410.000 512.400 ;
        RECT 398.000 511.600 398.800 511.800 ;
        RECT 396.400 510.300 397.200 510.400 ;
        RECT 400.000 510.300 400.600 511.800 ;
        RECT 396.400 509.700 400.600 510.300 ;
        RECT 396.400 509.600 397.200 509.700 ;
        RECT 400.000 508.400 400.600 509.700 ;
        RECT 401.200 510.300 402.000 510.400 ;
        RECT 402.800 510.300 403.600 510.400 ;
        RECT 401.200 509.700 403.600 510.300 ;
        RECT 401.200 508.800 402.000 509.700 ;
        RECT 402.800 509.600 403.600 509.700 ;
        RECT 405.800 508.400 406.400 511.800 ;
        RECT 407.400 509.800 408.000 511.800 ;
        RECT 407.000 509.000 408.000 509.800 ;
        RECT 396.400 506.800 397.200 508.400 ;
        RECT 398.000 507.600 400.600 508.400 ;
        RECT 402.800 508.300 403.600 508.400 ;
        RECT 405.800 508.300 406.800 508.400 ;
        RECT 402.800 508.200 406.800 508.300 ;
        RECT 402.000 507.700 406.800 508.200 ;
        RECT 402.000 507.600 403.600 507.700 ;
        RECT 405.800 507.600 406.800 507.700 ;
        RECT 398.200 506.200 398.800 507.600 ;
        RECT 402.000 507.200 402.800 507.600 ;
        RECT 399.800 506.200 403.400 506.600 ;
        RECT 405.800 506.200 406.400 507.600 ;
        RECT 407.400 507.400 408.000 509.000 ;
        RECT 409.000 509.600 410.000 510.400 ;
        RECT 409.000 508.800 409.800 509.600 ;
        RECT 412.400 508.300 413.200 519.800 ;
        RECT 417.800 518.400 418.600 519.800 ;
        RECT 417.200 517.600 418.600 518.400 ;
        RECT 417.800 512.800 418.600 517.600 ;
        RECT 422.000 515.000 422.800 519.000 ;
        RECT 417.000 512.200 418.600 512.800 ;
        RECT 415.600 509.600 416.400 511.200 ;
        RECT 417.000 508.400 417.600 512.200 ;
        RECT 422.200 511.600 422.800 515.000 ;
        RECT 426.200 512.400 427.000 519.800 ;
        RECT 427.600 513.600 428.400 514.400 ;
        RECT 427.800 512.400 428.400 513.600 ;
        RECT 431.600 512.800 432.400 519.800 ;
        RECT 426.200 511.800 427.200 512.400 ;
        RECT 427.800 511.800 429.200 512.400 ;
        RECT 419.000 511.000 422.800 511.600 ;
        RECT 419.000 509.000 419.600 511.000 ;
        RECT 414.000 508.300 414.800 508.400 ;
        RECT 412.400 507.700 414.800 508.300 ;
        RECT 407.400 506.800 410.000 507.400 ;
        RECT 386.800 506.000 390.800 506.200 ;
        RECT 377.200 503.000 378.000 505.000 ;
        RECT 381.400 503.000 382.200 506.000 ;
        RECT 386.800 502.200 387.600 506.000 ;
        RECT 390.000 502.200 390.800 506.000 ;
        RECT 391.600 502.200 392.400 506.200 ;
        RECT 393.800 505.600 395.600 506.200 ;
        RECT 393.800 504.400 394.600 505.600 ;
        RECT 393.200 503.600 394.600 504.400 ;
        RECT 393.800 502.200 394.600 503.600 ;
        RECT 398.000 502.200 398.800 506.200 ;
        RECT 399.600 506.000 403.600 506.200 ;
        RECT 399.600 502.200 400.400 506.000 ;
        RECT 402.800 502.200 403.600 506.000 ;
        RECT 405.800 505.600 406.800 506.200 ;
        RECT 406.000 502.200 406.800 505.600 ;
        RECT 409.200 502.200 410.000 506.800 ;
        RECT 410.800 504.800 411.600 506.400 ;
        RECT 412.400 502.200 413.200 507.700 ;
        RECT 414.000 507.600 414.800 507.700 ;
        RECT 415.600 507.600 417.600 508.400 ;
        RECT 418.200 508.200 419.600 509.000 ;
        RECT 420.400 508.800 421.200 510.400 ;
        RECT 422.000 508.800 422.800 510.400 ;
        RECT 425.200 508.800 426.000 510.400 ;
        RECT 426.600 508.400 427.200 511.800 ;
        RECT 428.400 511.600 429.200 511.800 ;
        RECT 431.400 511.800 432.400 512.800 ;
        RECT 434.800 512.400 435.600 519.800 ;
        RECT 433.000 511.800 435.600 512.400 ;
        RECT 431.400 508.400 432.000 511.800 ;
        RECT 433.000 509.800 433.600 511.800 ;
        RECT 436.400 511.600 437.200 513.200 ;
        RECT 432.600 509.000 433.600 509.800 ;
        RECT 417.000 507.000 417.600 507.600 ;
        RECT 418.600 507.800 419.600 508.200 ;
        RECT 423.600 508.200 424.400 508.400 ;
        RECT 418.600 507.200 422.800 507.800 ;
        RECT 423.600 507.600 425.200 508.200 ;
        RECT 426.600 507.600 429.200 508.400 ;
        RECT 431.400 507.600 432.400 508.400 ;
        RECT 424.400 507.200 425.200 507.600 ;
        RECT 417.000 506.600 417.800 507.000 ;
        RECT 417.000 506.000 418.600 506.600 ;
        RECT 417.800 503.000 418.600 506.000 ;
        RECT 422.200 505.000 422.800 507.200 ;
        RECT 423.800 506.200 427.400 506.600 ;
        RECT 428.400 506.200 429.000 507.600 ;
        RECT 431.400 506.200 432.000 507.600 ;
        RECT 433.000 507.400 433.600 509.000 ;
        RECT 434.600 509.600 435.600 510.400 ;
        RECT 434.600 508.800 435.400 509.600 ;
        RECT 436.400 508.300 437.200 508.400 ;
        RECT 438.000 508.300 438.800 519.800 ;
        RECT 441.200 512.400 442.000 519.800 ;
        RECT 444.400 512.800 445.200 519.800 ;
        RECT 451.400 518.400 452.200 519.800 ;
        RECT 451.400 517.600 453.200 518.400 ;
        RECT 451.400 512.800 452.200 517.600 ;
        RECT 455.600 515.000 456.400 519.000 ;
        RECT 441.200 511.800 443.800 512.400 ;
        RECT 444.400 511.800 445.400 512.800 ;
        RECT 441.200 509.600 442.200 510.400 ;
        RECT 441.400 508.800 442.200 509.600 ;
        RECT 443.200 509.800 443.800 511.800 ;
        RECT 443.200 509.000 444.200 509.800 ;
        RECT 436.400 507.700 438.800 508.300 ;
        RECT 436.400 507.600 437.200 507.700 ;
        RECT 433.000 506.800 435.600 507.400 ;
        RECT 422.000 503.000 422.800 505.000 ;
        RECT 423.600 506.000 427.600 506.200 ;
        RECT 423.600 502.200 424.400 506.000 ;
        RECT 426.800 502.200 427.600 506.000 ;
        RECT 428.400 502.200 429.200 506.200 ;
        RECT 431.400 505.600 432.400 506.200 ;
        RECT 431.600 502.200 432.400 505.600 ;
        RECT 434.800 502.200 435.600 506.800 ;
        RECT 438.000 506.200 438.800 507.700 ;
        RECT 439.600 506.800 440.400 508.400 ;
        RECT 443.200 507.400 443.800 509.000 ;
        RECT 444.800 508.400 445.400 511.800 ;
        RECT 450.600 512.200 452.200 512.800 ;
        RECT 447.600 510.300 448.400 510.400 ;
        RECT 449.200 510.300 450.000 511.200 ;
        RECT 447.600 509.700 450.000 510.300 ;
        RECT 447.600 509.600 448.400 509.700 ;
        RECT 449.200 509.600 450.000 509.700 ;
        RECT 450.600 508.400 451.200 512.200 ;
        RECT 455.800 511.600 456.400 515.000 ;
        RECT 452.600 511.000 456.400 511.600 ;
        RECT 452.600 509.000 453.200 511.000 ;
        RECT 444.400 507.600 445.400 508.400 ;
        RECT 449.200 507.600 451.200 508.400 ;
        RECT 451.800 508.200 453.200 509.000 ;
        RECT 454.000 508.800 454.800 510.400 ;
        RECT 455.600 508.800 456.400 510.400 ;
        RECT 441.200 506.800 443.800 507.400 ;
        RECT 437.000 505.600 438.800 506.200 ;
        RECT 437.000 502.200 437.800 505.600 ;
        RECT 441.200 502.200 442.000 506.800 ;
        RECT 444.800 506.200 445.400 507.600 ;
        RECT 444.400 505.600 445.400 506.200 ;
        RECT 450.600 507.000 451.200 507.600 ;
        RECT 452.200 507.800 453.200 508.200 ;
        RECT 452.200 507.200 456.400 507.800 ;
        RECT 450.600 506.600 451.400 507.000 ;
        RECT 450.600 506.000 452.200 506.600 ;
        RECT 444.400 502.200 445.200 505.600 ;
        RECT 451.400 503.000 452.200 506.000 ;
        RECT 455.800 505.000 456.400 507.200 ;
        RECT 455.600 503.000 456.400 505.000 ;
        RECT 457.200 504.300 458.000 504.400 ;
        RECT 462.000 504.300 462.800 519.800 ;
        RECT 465.200 511.600 466.000 513.200 ;
        RECT 463.600 504.800 464.400 506.400 ;
        RECT 466.800 506.200 467.600 519.800 ;
        RECT 470.000 515.000 470.800 519.000 ;
        RECT 474.200 518.400 475.000 519.800 ;
        RECT 474.200 517.600 475.600 518.400 ;
        RECT 470.000 511.600 470.600 515.000 ;
        RECT 474.200 512.800 475.000 517.600 ;
        RECT 474.200 512.200 475.800 512.800 ;
        RECT 470.000 511.000 473.800 511.600 ;
        RECT 470.000 508.800 470.800 510.400 ;
        RECT 471.600 508.800 472.400 510.400 ;
        RECT 473.200 509.000 473.800 511.000 ;
        RECT 468.400 506.800 469.200 508.400 ;
        RECT 473.200 508.200 474.600 509.000 ;
        RECT 475.200 508.400 475.800 512.200 ;
        RECT 476.400 509.600 477.200 511.200 ;
        RECT 473.200 507.800 474.200 508.200 ;
        RECT 470.000 507.200 474.200 507.800 ;
        RECT 475.200 507.600 477.200 508.400 ;
        RECT 465.800 505.600 467.600 506.200 ;
        RECT 465.800 504.400 466.600 505.600 ;
        RECT 457.200 503.700 462.800 504.300 ;
        RECT 457.200 503.600 458.000 503.700 ;
        RECT 462.000 502.200 462.800 503.700 ;
        RECT 465.200 503.600 466.600 504.400 ;
        RECT 465.800 502.200 466.600 503.600 ;
        RECT 470.000 505.000 470.600 507.200 ;
        RECT 475.200 507.000 475.800 507.600 ;
        RECT 475.000 506.600 475.800 507.000 ;
        RECT 479.600 506.800 480.400 508.400 ;
        RECT 474.200 506.000 475.800 506.600 ;
        RECT 481.200 506.200 482.000 519.800 ;
        RECT 488.200 518.400 489.000 519.800 ;
        RECT 488.200 517.600 490.000 518.400 ;
        RECT 482.800 511.600 483.600 514.400 ;
        RECT 488.200 512.800 489.000 517.600 ;
        RECT 492.400 515.000 493.200 519.000 ;
        RECT 487.400 512.200 489.000 512.800 ;
        RECT 486.000 509.600 486.800 511.200 ;
        RECT 487.400 508.400 488.000 512.200 ;
        RECT 492.600 511.600 493.200 515.000 ;
        RECT 495.600 512.800 496.400 519.800 ;
        RECT 489.400 511.000 493.200 511.600 ;
        RECT 495.400 511.800 496.400 512.800 ;
        RECT 498.800 512.400 499.600 519.800 ;
        RECT 497.000 511.800 499.600 512.400 ;
        RECT 489.400 509.000 490.000 511.000 ;
        RECT 486.000 507.600 488.000 508.400 ;
        RECT 488.600 508.200 490.000 509.000 ;
        RECT 490.800 508.800 491.600 510.400 ;
        RECT 492.400 510.300 493.200 510.400 ;
        RECT 494.000 510.300 494.800 510.400 ;
        RECT 492.400 509.700 494.800 510.300 ;
        RECT 492.400 508.800 493.200 509.700 ;
        RECT 494.000 509.600 494.800 509.700 ;
        RECT 487.400 507.000 488.000 507.600 ;
        RECT 489.000 507.800 490.000 508.200 ;
        RECT 495.400 508.400 496.000 511.800 ;
        RECT 497.000 509.800 497.600 511.800 ;
        RECT 496.600 509.000 497.600 509.800 ;
        RECT 489.000 507.200 493.200 507.800 ;
        RECT 487.400 506.600 488.200 507.000 ;
        RECT 470.000 503.000 470.800 505.000 ;
        RECT 474.200 503.000 475.000 506.000 ;
        RECT 481.200 505.600 483.000 506.200 ;
        RECT 487.400 506.000 489.000 506.600 ;
        RECT 482.200 504.400 483.000 505.600 ;
        RECT 481.200 503.600 483.000 504.400 ;
        RECT 482.200 502.200 483.000 503.600 ;
        RECT 488.200 503.000 489.000 506.000 ;
        RECT 492.600 505.000 493.200 507.200 ;
        RECT 495.400 507.600 496.400 508.400 ;
        RECT 495.400 506.200 496.000 507.600 ;
        RECT 497.000 507.400 497.600 509.000 ;
        RECT 498.600 509.600 499.600 510.400 ;
        RECT 498.600 508.800 499.400 509.600 ;
        RECT 497.000 506.800 499.600 507.400 ;
        RECT 500.400 506.800 501.200 508.400 ;
        RECT 495.400 505.600 496.400 506.200 ;
        RECT 492.400 503.000 493.200 505.000 ;
        RECT 495.600 502.200 496.400 505.600 ;
        RECT 498.800 502.200 499.600 506.800 ;
        RECT 502.000 506.200 502.800 519.800 ;
        RECT 503.600 511.600 504.400 514.400 ;
        RECT 505.200 512.400 506.000 519.800 ;
        RECT 508.400 512.800 509.200 519.800 ;
        RECT 505.200 511.800 507.800 512.400 ;
        RECT 508.400 511.800 509.400 512.800 ;
        RECT 514.200 512.400 515.000 519.800 ;
        RECT 515.600 513.600 516.400 514.400 ;
        RECT 515.800 512.400 516.400 513.600 ;
        RECT 514.200 511.800 515.200 512.400 ;
        RECT 515.800 511.800 517.200 512.400 ;
        RECT 505.200 509.600 506.200 510.400 ;
        RECT 505.400 508.800 506.200 509.600 ;
        RECT 507.200 509.800 507.800 511.800 ;
        RECT 507.200 509.000 508.200 509.800 ;
        RECT 507.200 507.400 507.800 509.000 ;
        RECT 508.800 508.400 509.400 511.800 ;
        RECT 510.000 510.300 510.800 510.400 ;
        RECT 513.200 510.300 514.000 510.400 ;
        RECT 510.000 509.700 514.000 510.300 ;
        RECT 510.000 509.600 510.800 509.700 ;
        RECT 513.200 508.800 514.000 509.700 ;
        RECT 514.600 508.400 515.200 511.800 ;
        RECT 516.400 511.600 517.200 511.800 ;
        RECT 508.400 507.600 509.400 508.400 ;
        RECT 511.600 508.200 512.400 508.400 ;
        RECT 511.600 507.600 513.200 508.200 ;
        RECT 514.600 507.600 517.200 508.400 ;
        RECT 505.200 506.800 507.800 507.400 ;
        RECT 502.000 505.600 503.800 506.200 ;
        RECT 503.000 504.400 503.800 505.600 ;
        RECT 503.000 503.600 504.400 504.400 ;
        RECT 503.000 502.200 503.800 503.600 ;
        RECT 505.200 502.200 506.000 506.800 ;
        RECT 508.800 506.200 509.400 507.600 ;
        RECT 512.400 507.200 513.200 507.600 ;
        RECT 511.800 506.200 515.400 506.600 ;
        RECT 516.400 506.200 517.000 507.600 ;
        RECT 508.400 505.600 509.400 506.200 ;
        RECT 511.600 506.000 515.600 506.200 ;
        RECT 508.400 502.200 509.200 505.600 ;
        RECT 511.600 502.200 512.400 506.000 ;
        RECT 514.800 502.200 515.600 506.000 ;
        RECT 516.400 502.200 517.200 506.200 ;
        RECT 518.000 502.200 518.800 519.800 ;
        RECT 521.200 515.000 522.000 519.000 ;
        RECT 521.200 511.600 521.800 515.000 ;
        RECT 525.400 512.800 526.200 519.800 ;
        RECT 525.400 512.200 527.000 512.800 ;
        RECT 526.000 511.600 527.000 512.200 ;
        RECT 533.400 512.400 534.200 519.800 ;
        RECT 534.800 513.600 535.600 514.400 ;
        RECT 535.000 512.400 535.600 513.600 ;
        RECT 539.800 512.400 540.600 519.800 ;
        RECT 546.200 514.400 547.000 519.800 ;
        RECT 541.200 513.600 542.000 514.400 ;
        RECT 545.200 513.600 547.000 514.400 ;
        RECT 547.600 514.300 548.400 514.400 ;
        RECT 550.000 514.300 550.800 519.800 ;
        RECT 554.200 515.800 555.400 519.800 ;
        RECT 558.800 515.800 559.600 519.800 ;
        RECT 563.200 516.400 564.000 519.800 ;
        RECT 563.200 515.800 565.200 516.400 ;
        RECT 554.800 515.000 555.600 515.800 ;
        RECT 559.000 515.200 559.600 515.800 ;
        RECT 558.200 514.600 561.800 515.200 ;
        RECT 564.400 515.000 565.200 515.800 ;
        RECT 558.200 514.400 559.000 514.600 ;
        RECT 561.000 514.400 561.800 514.600 ;
        RECT 547.600 513.700 550.800 514.300 ;
        RECT 547.600 513.600 548.400 513.700 ;
        RECT 541.400 512.400 542.000 513.600 ;
        RECT 546.200 512.400 547.000 513.600 ;
        RECT 547.800 512.400 548.400 513.600 ;
        RECT 533.400 511.800 534.400 512.400 ;
        RECT 535.000 511.800 536.400 512.400 ;
        RECT 539.800 511.800 540.800 512.400 ;
        RECT 541.400 511.800 542.800 512.400 ;
        RECT 546.200 511.800 547.200 512.400 ;
        RECT 547.800 511.800 549.200 512.400 ;
        RECT 521.200 511.000 525.000 511.600 ;
        RECT 521.200 508.800 522.000 510.400 ;
        RECT 522.800 508.800 523.600 510.400 ;
        RECT 524.400 509.000 525.000 511.000 ;
        RECT 524.400 508.200 525.800 509.000 ;
        RECT 526.400 508.400 527.000 511.600 ;
        RECT 527.600 509.600 528.400 511.200 ;
        RECT 529.200 510.300 530.000 510.400 ;
        RECT 532.400 510.300 533.200 510.400 ;
        RECT 529.200 509.700 533.200 510.300 ;
        RECT 529.200 509.600 530.000 509.700 ;
        RECT 532.400 508.800 533.200 509.700 ;
        RECT 533.800 508.400 534.400 511.800 ;
        RECT 535.600 511.600 536.400 511.800 ;
        RECT 538.800 508.800 539.600 510.400 ;
        RECT 540.200 510.300 540.800 511.800 ;
        RECT 542.000 511.600 542.800 511.800 ;
        RECT 543.600 510.300 544.400 510.400 ;
        RECT 540.200 509.700 544.400 510.300 ;
        RECT 540.200 508.400 540.800 509.700 ;
        RECT 543.600 509.600 544.400 509.700 ;
        RECT 545.200 508.800 546.000 510.400 ;
        RECT 546.600 508.400 547.200 511.800 ;
        RECT 548.400 511.600 549.200 511.800 ;
        RECT 550.000 511.200 550.800 513.700 ;
        RECT 554.000 513.200 555.400 514.000 ;
        RECT 554.800 512.200 555.400 513.200 ;
        RECT 557.000 513.000 559.200 513.600 ;
        RECT 557.000 512.800 557.800 513.000 ;
        RECT 554.800 511.600 557.200 512.200 ;
        RECT 550.000 510.600 554.200 511.200 ;
        RECT 524.400 507.800 525.400 508.200 ;
        RECT 521.200 507.200 525.400 507.800 ;
        RECT 526.400 507.600 528.400 508.400 ;
        RECT 529.200 508.300 530.000 508.400 ;
        RECT 530.800 508.300 531.600 508.400 ;
        RECT 529.200 508.200 531.600 508.300 ;
        RECT 529.200 507.700 532.400 508.200 ;
        RECT 529.200 507.600 530.000 507.700 ;
        RECT 530.800 507.600 532.400 507.700 ;
        RECT 533.800 507.600 536.400 508.400 ;
        RECT 537.200 508.200 538.000 508.400 ;
        RECT 537.200 507.600 538.800 508.200 ;
        RECT 540.200 507.600 542.800 508.400 ;
        RECT 543.600 508.200 544.400 508.400 ;
        RECT 543.600 507.600 545.200 508.200 ;
        RECT 546.600 507.600 549.200 508.400 ;
        RECT 519.600 504.800 520.400 506.400 ;
        RECT 521.200 505.000 521.800 507.200 ;
        RECT 526.400 507.000 527.000 507.600 ;
        RECT 531.600 507.200 532.400 507.600 ;
        RECT 526.200 506.600 527.000 507.000 ;
        RECT 525.400 506.000 527.000 506.600 ;
        RECT 531.000 506.200 534.600 506.600 ;
        RECT 535.600 506.400 536.200 507.600 ;
        RECT 538.000 507.200 538.800 507.600 ;
        RECT 530.800 506.000 534.800 506.200 ;
        RECT 521.200 503.000 522.000 505.000 ;
        RECT 525.400 503.000 526.200 506.000 ;
        RECT 530.800 502.200 531.600 506.000 ;
        RECT 534.000 502.200 534.800 506.000 ;
        RECT 535.600 502.200 536.400 506.400 ;
        RECT 537.400 506.200 541.000 506.600 ;
        RECT 542.000 506.200 542.600 507.600 ;
        RECT 544.400 507.200 545.200 507.600 ;
        RECT 543.800 506.200 547.400 506.600 ;
        RECT 548.400 506.200 549.000 507.600 ;
        RECT 550.000 507.200 550.800 510.600 ;
        RECT 553.400 510.400 554.200 510.600 ;
        RECT 551.800 509.800 552.600 510.000 ;
        RECT 551.800 509.200 555.600 509.800 ;
        RECT 554.800 509.000 555.600 509.200 ;
        RECT 556.600 508.400 557.200 511.600 ;
        RECT 558.600 511.800 559.200 513.000 ;
        RECT 559.800 513.000 560.600 513.200 ;
        RECT 564.400 513.000 565.200 513.200 ;
        RECT 559.800 512.400 565.200 513.000 ;
        RECT 558.600 511.400 563.400 511.800 ;
        RECT 567.600 511.400 568.400 519.800 ;
        RECT 569.200 511.600 570.000 513.200 ;
        RECT 558.600 511.200 568.400 511.400 ;
        RECT 562.600 511.000 568.400 511.200 ;
        RECT 562.800 510.800 568.400 511.000 ;
        RECT 561.200 510.200 562.000 510.400 ;
        RECT 561.200 509.600 566.200 510.200 ;
        RECT 565.400 509.400 566.200 509.600 ;
        RECT 563.800 508.400 564.600 508.600 ;
        RECT 556.600 507.800 567.600 508.400 ;
        RECT 557.000 507.600 557.800 507.800 ;
        RECT 550.000 506.600 553.800 507.200 ;
        RECT 537.200 506.000 541.200 506.200 ;
        RECT 537.200 502.200 538.000 506.000 ;
        RECT 540.400 502.200 541.200 506.000 ;
        RECT 542.000 502.200 542.800 506.200 ;
        RECT 543.600 506.000 547.600 506.200 ;
        RECT 543.600 502.200 544.400 506.000 ;
        RECT 546.800 502.200 547.600 506.000 ;
        RECT 548.400 502.200 549.200 506.200 ;
        RECT 550.000 502.200 550.800 506.600 ;
        RECT 553.000 506.400 553.800 506.600 ;
        RECT 562.800 505.600 563.400 507.800 ;
        RECT 566.000 507.600 567.600 507.800 ;
        RECT 561.000 505.400 561.800 505.600 ;
        RECT 554.800 504.200 555.600 505.000 ;
        RECT 559.000 504.800 561.800 505.400 ;
        RECT 562.800 504.800 563.600 505.600 ;
        RECT 559.000 504.200 559.600 504.800 ;
        RECT 564.400 504.200 565.200 505.000 ;
        RECT 554.200 503.600 555.600 504.200 ;
        RECT 554.200 502.200 555.400 503.600 ;
        RECT 558.800 502.200 559.600 504.200 ;
        RECT 563.200 503.600 565.200 504.200 ;
        RECT 563.200 502.200 564.000 503.600 ;
        RECT 567.600 502.200 568.400 507.000 ;
        RECT 570.800 506.200 571.600 519.800 ;
        RECT 575.600 512.000 576.400 519.800 ;
        RECT 578.800 515.200 579.600 519.800 ;
        RECT 575.400 511.200 576.400 512.000 ;
        RECT 577.000 514.600 579.600 515.200 ;
        RECT 577.000 513.000 577.600 514.600 ;
        RECT 582.000 514.400 582.800 519.800 ;
        RECT 585.200 517.000 586.000 519.800 ;
        RECT 586.800 517.000 587.600 519.800 ;
        RECT 588.400 517.000 589.200 519.800 ;
        RECT 583.400 514.400 587.600 515.200 ;
        RECT 580.200 513.600 582.800 514.400 ;
        RECT 590.000 513.600 590.800 519.800 ;
        RECT 593.200 515.000 594.000 519.800 ;
        RECT 596.400 515.000 597.200 519.800 ;
        RECT 598.000 517.000 598.800 519.800 ;
        RECT 599.600 517.000 600.400 519.800 ;
        RECT 602.800 515.200 603.600 519.800 ;
        RECT 606.000 516.400 606.800 519.800 ;
        RECT 606.000 515.800 607.000 516.400 ;
        RECT 606.400 515.200 607.000 515.800 ;
        RECT 601.600 514.400 605.800 515.200 ;
        RECT 606.400 514.600 608.400 515.200 ;
        RECT 593.200 513.600 595.800 514.400 ;
        RECT 596.400 513.800 602.200 514.400 ;
        RECT 605.200 514.000 605.800 514.400 ;
        RECT 585.200 513.000 586.000 513.200 ;
        RECT 577.000 512.400 586.000 513.000 ;
        RECT 588.400 513.000 589.200 513.200 ;
        RECT 596.400 513.000 597.000 513.800 ;
        RECT 602.800 513.200 604.200 513.800 ;
        RECT 605.200 513.200 606.800 514.000 ;
        RECT 588.400 512.400 597.000 513.000 ;
        RECT 598.000 513.000 604.200 513.200 ;
        RECT 598.000 512.600 603.400 513.000 ;
        RECT 598.000 512.400 598.800 512.600 ;
        RECT 572.400 506.800 573.200 508.400 ;
        RECT 575.400 506.800 576.200 511.200 ;
        RECT 577.000 510.600 577.600 512.400 ;
        RECT 576.800 510.000 577.600 510.600 ;
        RECT 583.600 510.000 607.000 510.600 ;
        RECT 576.800 508.000 577.400 510.000 ;
        RECT 583.600 509.400 584.400 510.000 ;
        RECT 601.200 509.600 602.000 510.000 ;
        RECT 604.400 509.600 605.200 510.000 ;
        RECT 606.200 509.800 607.000 510.000 ;
        RECT 578.000 508.600 581.800 509.400 ;
        RECT 576.800 507.400 578.000 508.000 ;
        RECT 569.800 505.600 571.600 506.200 ;
        RECT 575.400 506.000 576.400 506.800 ;
        RECT 569.800 504.400 570.600 505.600 ;
        RECT 569.800 503.600 571.600 504.400 ;
        RECT 569.800 502.200 570.600 503.600 ;
        RECT 575.600 502.200 576.400 506.000 ;
        RECT 577.200 502.200 578.000 507.400 ;
        RECT 581.000 507.400 581.800 508.600 ;
        RECT 581.000 506.800 582.800 507.400 ;
        RECT 582.000 506.200 582.800 506.800 ;
        RECT 586.800 506.400 587.600 509.200 ;
        RECT 590.000 508.600 593.200 509.400 ;
        RECT 597.000 508.600 599.000 509.400 ;
        RECT 607.600 509.000 608.400 514.600 ;
        RECT 589.600 507.800 590.400 508.000 ;
        RECT 589.600 507.200 594.000 507.800 ;
        RECT 593.200 507.000 594.000 507.200 ;
        RECT 594.800 506.800 595.600 508.400 ;
        RECT 582.000 505.400 584.400 506.200 ;
        RECT 586.800 505.600 587.800 506.400 ;
        RECT 590.800 505.600 592.400 506.400 ;
        RECT 593.200 506.200 594.000 506.400 ;
        RECT 597.000 506.200 597.800 508.600 ;
        RECT 599.600 508.200 608.400 509.000 ;
        RECT 603.000 506.800 606.000 507.600 ;
        RECT 603.000 506.200 603.800 506.800 ;
        RECT 593.200 505.600 597.800 506.200 ;
        RECT 583.600 502.200 584.400 505.400 ;
        RECT 601.200 505.400 603.800 506.200 ;
        RECT 585.200 502.200 586.000 505.000 ;
        RECT 586.800 502.200 587.600 505.000 ;
        RECT 588.400 502.200 589.200 505.000 ;
        RECT 590.000 502.200 590.800 505.000 ;
        RECT 593.200 502.200 594.000 505.000 ;
        RECT 596.400 502.200 597.200 505.000 ;
        RECT 598.000 502.200 598.800 505.000 ;
        RECT 599.600 502.200 600.400 505.000 ;
        RECT 601.200 502.200 602.000 505.400 ;
        RECT 607.600 502.200 608.400 508.200 ;
        RECT 1.200 495.800 2.000 499.800 ;
        RECT 2.800 496.000 3.600 499.800 ;
        RECT 6.000 496.000 6.800 499.800 ;
        RECT 11.400 496.000 12.200 499.000 ;
        RECT 15.600 497.000 16.400 499.000 ;
        RECT 2.800 495.800 6.800 496.000 ;
        RECT 1.400 494.400 2.000 495.800 ;
        RECT 3.000 495.400 6.600 495.800 ;
        RECT 10.600 495.400 12.200 496.000 ;
        RECT 10.600 495.000 11.400 495.400 ;
        RECT 5.200 494.400 6.000 494.800 ;
        RECT 10.600 494.400 11.200 495.000 ;
        RECT 15.800 494.800 16.400 497.000 ;
        RECT 17.200 495.800 18.000 499.800 ;
        RECT 18.800 496.000 19.600 499.800 ;
        RECT 22.000 496.000 22.800 499.800 ;
        RECT 18.800 495.800 22.800 496.000 ;
        RECT 1.200 493.600 3.800 494.400 ;
        RECT 5.200 493.800 6.800 494.400 ;
        RECT 9.200 494.300 11.200 494.400 ;
        RECT 6.000 493.600 6.800 493.800 ;
        RECT 7.700 493.700 11.200 494.300 ;
        RECT 12.200 494.200 16.400 494.800 ;
        RECT 17.400 494.400 18.000 495.800 ;
        RECT 19.000 495.400 22.600 495.800 ;
        RECT 23.600 495.000 24.400 499.800 ;
        RECT 28.000 498.400 28.800 499.800 ;
        RECT 26.800 497.800 28.800 498.400 ;
        RECT 32.400 497.800 33.200 499.800 ;
        RECT 36.600 498.400 37.800 499.800 ;
        RECT 36.400 497.800 37.800 498.400 ;
        RECT 26.800 497.000 27.600 497.800 ;
        RECT 32.400 497.200 33.000 497.800 ;
        RECT 28.400 496.400 29.200 497.200 ;
        RECT 30.200 496.600 33.000 497.200 ;
        RECT 36.400 497.000 37.200 497.800 ;
        RECT 30.200 496.400 31.000 496.600 ;
        RECT 21.200 494.400 22.000 494.800 ;
        RECT 12.200 493.800 13.200 494.200 ;
        RECT 1.200 490.200 2.000 490.400 ;
        RECT 3.200 490.200 3.800 493.600 ;
        RECT 4.400 492.300 5.200 493.200 ;
        RECT 7.700 492.300 8.300 493.700 ;
        RECT 9.200 493.600 11.200 493.700 ;
        RECT 4.400 491.700 8.300 492.300 ;
        RECT 4.400 491.600 5.200 491.700 ;
        RECT 9.200 490.800 10.000 492.400 ;
        RECT 1.200 489.600 2.600 490.200 ;
        RECT 3.200 489.600 4.200 490.200 ;
        RECT 2.000 488.400 2.600 489.600 ;
        RECT 2.000 487.600 2.800 488.400 ;
        RECT 3.400 482.200 4.200 489.600 ;
        RECT 10.600 489.800 11.200 493.600 ;
        RECT 11.800 493.000 13.200 493.800 ;
        RECT 17.200 493.600 19.800 494.400 ;
        RECT 21.200 493.800 22.800 494.400 ;
        RECT 22.000 493.600 22.800 493.800 ;
        RECT 24.400 494.200 26.000 494.400 ;
        RECT 28.600 494.200 29.200 496.400 ;
        RECT 38.200 495.400 39.000 495.600 ;
        RECT 41.200 495.400 42.000 499.800 ;
        RECT 42.800 496.000 43.600 499.800 ;
        RECT 46.000 496.000 46.800 499.800 ;
        RECT 42.800 495.800 46.800 496.000 ;
        RECT 47.600 495.800 48.400 499.800 ;
        RECT 53.000 496.000 53.800 499.000 ;
        RECT 57.200 497.000 58.000 499.000 ;
        RECT 43.000 495.400 46.600 495.800 ;
        RECT 38.200 494.800 42.000 495.400 ;
        RECT 34.200 494.200 35.000 494.400 ;
        RECT 24.400 493.600 35.400 494.200 ;
        RECT 12.600 491.000 13.200 493.000 ;
        RECT 14.000 491.600 14.800 493.200 ;
        RECT 15.600 491.600 16.400 493.200 ;
        RECT 12.600 490.400 16.400 491.000 ;
        RECT 10.600 489.200 12.200 489.800 ;
        RECT 11.400 482.200 12.200 489.200 ;
        RECT 15.800 487.000 16.400 490.400 ;
        RECT 17.200 490.200 18.000 490.400 ;
        RECT 19.200 490.200 19.800 493.600 ;
        RECT 27.400 493.400 28.200 493.600 ;
        RECT 20.400 491.600 21.200 493.200 ;
        RECT 25.800 492.400 26.600 492.600 ;
        RECT 25.800 491.800 30.800 492.400 ;
        RECT 30.000 491.600 30.800 491.800 ;
        RECT 23.600 491.000 29.200 491.200 ;
        RECT 23.600 490.800 29.400 491.000 ;
        RECT 23.600 490.600 33.400 490.800 ;
        RECT 17.200 489.600 18.600 490.200 ;
        RECT 19.200 489.600 20.200 490.200 ;
        RECT 18.000 488.400 18.600 489.600 ;
        RECT 18.000 487.600 18.800 488.400 ;
        RECT 15.600 483.000 16.400 487.000 ;
        RECT 19.400 482.200 20.200 489.600 ;
        RECT 23.600 482.200 24.400 490.600 ;
        RECT 28.600 490.200 33.400 490.600 ;
        RECT 26.800 489.000 32.200 489.600 ;
        RECT 26.800 488.800 27.600 489.000 ;
        RECT 31.400 488.800 32.200 489.000 ;
        RECT 32.800 489.000 33.400 490.200 ;
        RECT 34.800 490.400 35.400 493.600 ;
        RECT 36.400 492.800 37.200 493.000 ;
        RECT 36.400 492.200 40.200 492.800 ;
        RECT 39.400 492.000 40.200 492.200 ;
        RECT 37.800 491.400 38.600 491.600 ;
        RECT 41.200 491.400 42.000 494.800 ;
        RECT 43.600 494.400 44.400 494.800 ;
        RECT 47.600 494.400 48.200 495.800 ;
        RECT 52.200 495.400 53.800 496.000 ;
        RECT 52.200 495.000 53.000 495.400 ;
        RECT 52.200 494.400 52.800 495.000 ;
        RECT 57.400 494.800 58.000 497.000 ;
        RECT 58.800 495.800 59.600 499.800 ;
        RECT 60.400 496.000 61.200 499.800 ;
        RECT 63.600 496.000 64.400 499.800 ;
        RECT 60.400 495.800 64.400 496.000 ;
        RECT 65.200 497.000 66.000 499.000 ;
        RECT 42.800 493.800 44.400 494.400 ;
        RECT 42.800 493.600 43.600 493.800 ;
        RECT 45.800 493.600 48.400 494.400 ;
        RECT 49.200 494.300 50.000 494.400 ;
        RECT 50.800 494.300 52.800 494.400 ;
        RECT 49.200 493.700 52.800 494.300 ;
        RECT 53.800 494.200 58.000 494.800 ;
        RECT 59.000 494.400 59.600 495.800 ;
        RECT 60.600 495.400 64.200 495.800 ;
        RECT 65.200 494.800 65.800 497.000 ;
        RECT 69.400 496.000 70.200 499.000 ;
        RECT 77.400 496.400 78.200 499.800 ;
        RECT 82.200 496.400 83.000 499.800 ;
        RECT 69.400 495.400 71.000 496.000 ;
        RECT 70.200 495.000 71.000 495.400 ;
        RECT 76.400 495.800 78.200 496.400 ;
        RECT 81.200 495.800 83.000 496.400 ;
        RECT 62.800 494.400 63.600 494.800 ;
        RECT 53.800 493.800 54.800 494.200 ;
        RECT 49.200 493.600 50.000 493.700 ;
        RECT 50.800 493.600 52.800 493.700 ;
        RECT 44.400 491.600 45.200 493.200 ;
        RECT 45.800 492.400 46.400 493.600 ;
        RECT 45.800 491.600 46.800 492.400 ;
        RECT 49.200 492.300 50.000 492.400 ;
        RECT 50.800 492.300 51.600 492.400 ;
        RECT 49.200 491.700 51.600 492.300 ;
        RECT 49.200 491.600 50.000 491.700 ;
        RECT 37.800 490.800 42.000 491.400 ;
        RECT 34.800 489.800 37.200 490.400 ;
        RECT 34.200 489.000 35.000 489.200 ;
        RECT 32.800 488.400 35.000 489.000 ;
        RECT 36.600 488.800 37.200 489.800 ;
        RECT 36.600 488.400 38.000 488.800 ;
        RECT 36.600 488.000 38.800 488.400 ;
        RECT 37.400 487.600 38.800 488.000 ;
        RECT 30.200 487.400 31.000 487.600 ;
        RECT 33.000 487.400 33.800 487.600 ;
        RECT 26.800 486.200 27.600 487.000 ;
        RECT 30.200 486.800 33.800 487.400 ;
        RECT 32.400 486.200 33.000 486.800 ;
        RECT 36.400 486.200 37.200 487.000 ;
        RECT 26.800 485.600 28.800 486.200 ;
        RECT 28.000 482.200 28.800 485.600 ;
        RECT 32.400 482.200 33.200 486.200 ;
        RECT 36.600 482.200 37.800 486.200 ;
        RECT 41.200 482.200 42.000 490.800 ;
        RECT 45.800 490.200 46.400 491.600 ;
        RECT 50.800 490.800 51.600 491.700 ;
        RECT 47.600 490.200 48.400 490.400 ;
        RECT 45.400 489.600 46.400 490.200 ;
        RECT 47.000 489.600 48.400 490.200 ;
        RECT 52.200 489.800 52.800 493.600 ;
        RECT 53.400 493.000 54.800 493.800 ;
        RECT 58.800 493.600 61.400 494.400 ;
        RECT 62.800 493.800 64.400 494.400 ;
        RECT 65.200 494.200 69.400 494.800 ;
        RECT 63.600 493.600 64.400 493.800 ;
        RECT 68.400 493.800 69.400 494.200 ;
        RECT 70.400 494.400 71.000 495.000 ;
        RECT 54.200 491.000 54.800 493.000 ;
        RECT 55.600 491.600 56.400 493.200 ;
        RECT 57.200 491.600 58.000 493.200 ;
        RECT 58.800 492.300 59.600 492.400 ;
        RECT 60.800 492.300 61.400 493.600 ;
        RECT 58.800 491.700 61.400 492.300 ;
        RECT 58.800 491.600 59.600 491.700 ;
        RECT 54.200 490.400 58.000 491.000 ;
        RECT 45.400 482.200 46.200 489.600 ;
        RECT 47.000 488.400 47.600 489.600 ;
        RECT 52.200 489.200 53.800 489.800 ;
        RECT 46.800 487.600 47.600 488.400 ;
        RECT 53.000 482.200 53.800 489.200 ;
        RECT 57.400 487.000 58.000 490.400 ;
        RECT 58.800 490.200 59.600 490.400 ;
        RECT 60.800 490.200 61.400 491.700 ;
        RECT 62.000 491.600 62.800 493.200 ;
        RECT 65.200 491.600 66.000 493.200 ;
        RECT 66.800 491.600 67.600 493.200 ;
        RECT 68.400 493.000 69.800 493.800 ;
        RECT 70.400 493.600 72.400 494.400 ;
        RECT 74.800 493.600 75.600 495.200 ;
        RECT 68.400 491.000 69.000 493.000 ;
        RECT 65.200 490.400 69.000 491.000 ;
        RECT 58.800 489.600 60.200 490.200 ;
        RECT 60.800 489.600 61.800 490.200 ;
        RECT 59.600 488.400 60.200 489.600 ;
        RECT 59.600 487.600 60.400 488.400 ;
        RECT 57.200 483.000 58.000 487.000 ;
        RECT 61.000 482.200 61.800 489.600 ;
        RECT 65.200 487.000 65.800 490.400 ;
        RECT 70.400 489.800 71.000 493.600 ;
        RECT 71.600 490.800 72.400 492.400 ;
        RECT 76.400 492.300 77.200 495.800 ;
        RECT 79.600 493.600 80.400 495.200 ;
        RECT 79.600 492.300 80.400 492.400 ;
        RECT 76.400 491.700 80.400 492.300 ;
        RECT 69.400 489.200 71.000 489.800 ;
        RECT 65.200 483.000 66.000 487.000 ;
        RECT 69.400 482.200 70.200 489.200 ;
        RECT 76.400 482.200 77.200 491.700 ;
        RECT 79.600 491.600 80.400 491.700 ;
        RECT 78.000 488.800 78.800 490.400 ;
        RECT 81.200 482.200 82.000 495.800 ;
        RECT 84.400 495.600 85.200 497.200 ;
        RECT 82.800 488.800 83.600 490.400 ;
        RECT 86.000 482.200 86.800 499.800 ;
        RECT 87.600 496.000 88.400 499.800 ;
        RECT 90.800 496.000 91.600 499.800 ;
        RECT 87.600 495.800 91.600 496.000 ;
        RECT 92.400 495.800 93.200 499.800 ;
        RECT 94.000 495.800 94.800 499.800 ;
        RECT 95.600 496.000 96.400 499.800 ;
        RECT 98.800 496.000 99.600 499.800 ;
        RECT 95.600 495.800 99.600 496.000 ;
        RECT 100.400 495.800 101.200 499.800 ;
        RECT 102.000 496.000 102.800 499.800 ;
        RECT 105.200 496.000 106.000 499.800 ;
        RECT 102.000 495.800 106.000 496.000 ;
        RECT 87.800 495.400 91.400 495.800 ;
        RECT 88.400 494.400 89.200 494.800 ;
        RECT 92.400 494.400 93.000 495.800 ;
        RECT 94.200 494.400 94.800 495.800 ;
        RECT 95.800 495.400 99.400 495.800 ;
        RECT 98.000 494.400 98.800 494.800 ;
        RECT 100.600 494.400 101.200 495.800 ;
        RECT 102.200 495.400 105.800 495.800 ;
        RECT 104.400 494.400 105.200 494.800 ;
        RECT 87.600 493.800 89.200 494.400 ;
        RECT 87.600 493.600 88.400 493.800 ;
        RECT 90.600 493.600 93.200 494.400 ;
        RECT 94.000 493.600 96.600 494.400 ;
        RECT 98.000 493.800 99.600 494.400 ;
        RECT 98.800 493.600 99.600 493.800 ;
        RECT 100.400 493.600 103.000 494.400 ;
        RECT 104.400 493.800 106.000 494.400 ;
        RECT 110.400 494.200 111.200 499.800 ;
        RECT 113.200 495.800 114.000 499.800 ;
        RECT 114.800 496.000 115.600 499.800 ;
        RECT 118.000 496.000 118.800 499.800 ;
        RECT 122.200 496.400 123.000 499.800 ;
        RECT 114.800 495.800 118.800 496.000 ;
        RECT 121.200 495.800 123.000 496.400 ;
        RECT 126.000 497.800 126.800 499.800 ;
        RECT 113.400 494.400 114.000 495.800 ;
        RECT 115.000 495.400 118.600 495.800 ;
        RECT 117.200 494.400 118.000 494.800 ;
        RECT 110.400 493.800 112.200 494.200 ;
        RECT 105.200 493.600 106.000 493.800 ;
        RECT 110.600 493.600 112.200 493.800 ;
        RECT 113.200 493.600 115.800 494.400 ;
        RECT 117.200 493.800 118.800 494.400 ;
        RECT 118.000 493.600 118.800 493.800 ;
        RECT 119.600 493.600 120.400 495.200 ;
        RECT 89.200 491.600 90.000 493.200 ;
        RECT 90.600 492.300 91.200 493.600 ;
        RECT 90.600 491.700 94.700 492.300 ;
        RECT 90.600 490.200 91.200 491.700 ;
        RECT 94.100 490.400 94.700 491.700 ;
        RECT 92.400 490.200 93.200 490.400 ;
        RECT 90.200 489.600 91.200 490.200 ;
        RECT 91.800 489.600 93.200 490.200 ;
        RECT 94.000 490.200 94.800 490.400 ;
        RECT 96.000 490.200 96.600 493.600 ;
        RECT 97.200 492.300 98.000 493.200 ;
        RECT 98.800 492.300 99.600 492.400 ;
        RECT 97.200 491.700 99.600 492.300 ;
        RECT 97.200 491.600 98.000 491.700 ;
        RECT 98.800 491.600 99.600 491.700 ;
        RECT 100.400 490.200 101.200 490.400 ;
        RECT 102.400 490.200 103.000 493.600 ;
        RECT 103.600 491.600 104.400 493.200 ;
        RECT 108.400 491.600 110.000 492.400 ;
        RECT 94.000 489.600 95.400 490.200 ;
        RECT 96.000 489.600 97.000 490.200 ;
        RECT 100.400 489.600 101.800 490.200 ;
        RECT 102.400 489.600 103.400 490.200 ;
        RECT 106.800 489.600 107.600 491.200 ;
        RECT 111.600 490.400 112.200 493.600 ;
        RECT 111.600 489.600 112.400 490.400 ;
        RECT 113.200 490.200 114.000 490.400 ;
        RECT 115.200 490.200 115.800 493.600 ;
        RECT 116.400 491.600 117.200 493.200 ;
        RECT 113.200 489.600 114.600 490.200 ;
        RECT 115.200 489.600 116.200 490.200 ;
        RECT 90.200 482.200 91.000 489.600 ;
        RECT 91.800 488.400 92.400 489.600 ;
        RECT 91.600 487.600 92.400 488.400 ;
        RECT 94.800 488.400 95.400 489.600 ;
        RECT 94.800 487.600 95.600 488.400 ;
        RECT 96.200 482.200 97.000 489.600 ;
        RECT 101.200 488.400 101.800 489.600 ;
        RECT 101.200 487.600 102.000 488.400 ;
        RECT 102.600 486.400 103.400 489.600 ;
        RECT 110.000 487.600 110.800 489.200 ;
        RECT 111.600 487.000 112.200 489.600 ;
        RECT 114.000 488.400 114.600 489.600 ;
        RECT 114.000 487.600 114.800 488.400 ;
        RECT 108.600 486.400 112.200 487.000 ;
        RECT 102.600 485.600 104.400 486.400 ;
        RECT 108.600 486.200 109.200 486.400 ;
        RECT 102.600 482.200 103.400 485.600 ;
        RECT 108.400 482.200 109.200 486.200 ;
        RECT 111.600 486.200 112.200 486.400 ;
        RECT 111.600 482.200 112.400 486.200 ;
        RECT 115.400 484.400 116.200 489.600 ;
        RECT 115.400 483.600 117.200 484.400 ;
        RECT 115.400 482.200 116.200 483.600 ;
        RECT 121.200 482.200 122.000 495.800 ;
        RECT 126.000 494.400 126.600 497.800 ;
        RECT 127.600 496.300 128.400 497.200 ;
        RECT 130.800 496.300 131.600 499.800 ;
        RECT 127.600 495.700 131.600 496.300 ;
        RECT 127.600 495.600 128.400 495.700 ;
        RECT 130.600 495.200 131.600 495.700 ;
        RECT 126.000 494.300 126.800 494.400 ;
        RECT 127.600 494.300 128.400 494.400 ;
        RECT 126.000 493.700 128.400 494.300 ;
        RECT 126.000 493.600 126.800 493.700 ;
        RECT 127.600 493.600 128.400 493.700 ;
        RECT 124.400 492.300 125.200 492.400 ;
        RECT 122.900 491.700 125.200 492.300 ;
        RECT 122.900 490.400 123.500 491.700 ;
        RECT 124.400 490.800 125.200 491.700 ;
        RECT 122.800 488.800 123.600 490.400 ;
        RECT 126.000 490.200 126.600 493.600 ;
        RECT 130.600 490.800 131.400 495.200 ;
        RECT 132.400 494.600 133.200 499.800 ;
        RECT 138.800 496.600 139.600 499.800 ;
        RECT 140.400 497.000 141.200 499.800 ;
        RECT 142.000 497.000 142.800 499.800 ;
        RECT 143.600 497.000 144.400 499.800 ;
        RECT 145.200 497.000 146.000 499.800 ;
        RECT 148.400 497.000 149.200 499.800 ;
        RECT 151.600 497.000 152.400 499.800 ;
        RECT 153.200 497.000 154.000 499.800 ;
        RECT 154.800 497.000 155.600 499.800 ;
        RECT 137.200 495.800 139.600 496.600 ;
        RECT 156.400 496.600 157.200 499.800 ;
        RECT 137.200 495.200 138.000 495.800 ;
        RECT 132.000 494.000 133.200 494.600 ;
        RECT 136.200 494.600 138.000 495.200 ;
        RECT 142.000 495.600 143.000 496.400 ;
        RECT 146.000 495.600 147.600 496.400 ;
        RECT 148.400 495.800 153.000 496.400 ;
        RECT 156.400 495.800 159.000 496.600 ;
        RECT 148.400 495.600 149.200 495.800 ;
        RECT 132.000 492.000 132.600 494.000 ;
        RECT 136.200 493.400 137.000 494.600 ;
        RECT 133.200 492.600 137.000 493.400 ;
        RECT 142.000 492.800 142.800 495.600 ;
        RECT 148.400 494.800 149.200 495.000 ;
        RECT 144.800 494.200 149.200 494.800 ;
        RECT 144.800 494.000 145.600 494.200 ;
        RECT 150.000 493.600 150.800 495.200 ;
        RECT 152.200 493.400 153.000 495.800 ;
        RECT 158.200 495.200 159.000 495.800 ;
        RECT 158.200 494.400 161.200 495.200 ;
        RECT 162.800 493.800 163.600 499.800 ;
        RECT 145.200 492.600 148.400 493.400 ;
        RECT 152.200 492.600 154.200 493.400 ;
        RECT 154.800 493.000 163.600 493.800 ;
        RECT 138.800 492.000 139.600 492.600 ;
        RECT 156.400 492.000 157.200 492.400 ;
        RECT 159.600 492.000 160.400 492.400 ;
        RECT 161.400 492.000 162.200 492.200 ;
        RECT 132.000 491.400 132.800 492.000 ;
        RECT 138.800 491.400 162.200 492.000 ;
        RECT 125.000 489.400 126.800 490.200 ;
        RECT 130.600 490.000 131.600 490.800 ;
        RECT 125.000 482.200 125.800 489.400 ;
        RECT 130.800 482.200 131.600 490.000 ;
        RECT 132.200 489.600 132.800 491.400 ;
        RECT 132.200 489.000 141.200 489.600 ;
        RECT 132.200 487.400 132.800 489.000 ;
        RECT 140.400 488.800 141.200 489.000 ;
        RECT 143.600 489.000 152.200 489.600 ;
        RECT 143.600 488.800 144.400 489.000 ;
        RECT 135.400 487.600 138.000 488.400 ;
        RECT 132.200 486.800 134.800 487.400 ;
        RECT 134.000 482.200 134.800 486.800 ;
        RECT 137.200 482.200 138.000 487.600 ;
        RECT 138.600 486.800 142.800 487.600 ;
        RECT 140.400 482.200 141.200 485.000 ;
        RECT 142.000 482.200 142.800 485.000 ;
        RECT 143.600 482.200 144.400 485.000 ;
        RECT 145.200 482.200 146.000 488.400 ;
        RECT 148.400 487.600 151.000 488.400 ;
        RECT 151.600 488.200 152.200 489.000 ;
        RECT 153.200 489.400 154.000 489.600 ;
        RECT 153.200 489.000 158.600 489.400 ;
        RECT 153.200 488.800 159.400 489.000 ;
        RECT 158.000 488.200 159.400 488.800 ;
        RECT 151.600 487.600 157.400 488.200 ;
        RECT 160.400 488.000 162.000 488.800 ;
        RECT 160.400 487.600 161.000 488.000 ;
        RECT 148.400 482.200 149.200 487.000 ;
        RECT 151.600 482.200 152.400 487.000 ;
        RECT 156.800 486.800 161.000 487.600 ;
        RECT 162.800 487.400 163.600 493.000 ;
        RECT 170.800 497.800 171.600 499.800 ;
        RECT 170.800 494.400 171.400 497.800 ;
        RECT 172.400 496.300 173.200 497.200 ;
        RECT 174.000 496.300 174.800 496.400 ;
        RECT 172.400 495.700 174.800 496.300 ;
        RECT 175.600 496.000 176.400 499.800 ;
        RECT 172.400 495.600 173.200 495.700 ;
        RECT 174.000 495.600 174.800 495.700 ;
        RECT 175.400 495.200 176.400 496.000 ;
        RECT 170.800 493.600 171.600 494.400 ;
        RECT 169.200 490.800 170.000 492.400 ;
        RECT 170.800 490.200 171.400 493.600 ;
        RECT 175.400 490.800 176.200 495.200 ;
        RECT 177.200 494.600 178.000 499.800 ;
        RECT 183.600 496.600 184.400 499.800 ;
        RECT 185.200 497.000 186.000 499.800 ;
        RECT 186.800 497.000 187.600 499.800 ;
        RECT 188.400 497.000 189.200 499.800 ;
        RECT 190.000 497.000 190.800 499.800 ;
        RECT 193.200 497.000 194.000 499.800 ;
        RECT 196.400 497.000 197.200 499.800 ;
        RECT 198.000 497.000 198.800 499.800 ;
        RECT 199.600 497.000 200.400 499.800 ;
        RECT 182.000 495.800 184.400 496.600 ;
        RECT 201.200 496.600 202.000 499.800 ;
        RECT 182.000 495.200 182.800 495.800 ;
        RECT 176.800 494.000 178.000 494.600 ;
        RECT 181.000 494.600 182.800 495.200 ;
        RECT 186.800 495.600 187.800 496.400 ;
        RECT 190.800 495.600 192.400 496.400 ;
        RECT 193.200 495.800 197.800 496.400 ;
        RECT 201.200 495.800 203.800 496.600 ;
        RECT 193.200 495.600 194.000 495.800 ;
        RECT 176.800 492.000 177.400 494.000 ;
        RECT 181.000 493.400 181.800 494.600 ;
        RECT 178.000 492.600 181.800 493.400 ;
        RECT 186.800 492.800 187.600 495.600 ;
        RECT 193.200 494.800 194.000 495.000 ;
        RECT 189.600 494.200 194.000 494.800 ;
        RECT 189.600 494.000 190.400 494.200 ;
        RECT 194.800 493.600 195.600 495.200 ;
        RECT 197.000 493.400 197.800 495.800 ;
        RECT 203.000 495.200 203.800 495.800 ;
        RECT 203.000 494.400 206.000 495.200 ;
        RECT 207.600 493.800 208.400 499.800 ;
        RECT 210.800 496.000 211.600 499.800 ;
        RECT 190.000 492.600 193.200 493.400 ;
        RECT 197.000 492.600 199.000 493.400 ;
        RECT 199.600 493.000 208.400 493.800 ;
        RECT 183.600 492.000 184.400 492.600 ;
        RECT 201.200 492.000 202.000 492.400 ;
        RECT 204.400 492.000 205.200 492.400 ;
        RECT 206.200 492.000 207.000 492.200 ;
        RECT 176.800 491.400 177.600 492.000 ;
        RECT 183.600 491.400 207.000 492.000 ;
        RECT 161.600 486.800 163.600 487.400 ;
        RECT 169.800 489.400 171.600 490.200 ;
        RECT 175.400 490.000 176.400 490.800 ;
        RECT 153.200 482.200 154.000 485.000 ;
        RECT 154.800 482.200 155.600 485.000 ;
        RECT 158.000 482.200 158.800 486.800 ;
        RECT 161.600 486.200 162.200 486.800 ;
        RECT 161.200 485.600 162.200 486.200 ;
        RECT 161.200 482.200 162.000 485.600 ;
        RECT 169.800 484.400 170.600 489.400 ;
        RECT 169.800 483.600 171.600 484.400 ;
        RECT 169.800 482.200 170.600 483.600 ;
        RECT 175.600 482.200 176.400 490.000 ;
        RECT 177.000 489.600 177.600 491.400 ;
        RECT 177.000 489.000 186.000 489.600 ;
        RECT 177.000 487.400 177.600 489.000 ;
        RECT 185.200 488.800 186.000 489.000 ;
        RECT 188.400 489.000 197.000 489.600 ;
        RECT 188.400 488.800 189.200 489.000 ;
        RECT 180.200 487.600 182.800 488.400 ;
        RECT 177.000 486.800 179.600 487.400 ;
        RECT 178.800 482.200 179.600 486.800 ;
        RECT 182.000 482.200 182.800 487.600 ;
        RECT 183.400 486.800 187.600 487.600 ;
        RECT 185.200 482.200 186.000 485.000 ;
        RECT 186.800 482.200 187.600 485.000 ;
        RECT 188.400 482.200 189.200 485.000 ;
        RECT 190.000 482.200 190.800 488.400 ;
        RECT 193.200 487.600 195.800 488.400 ;
        RECT 196.400 488.200 197.000 489.000 ;
        RECT 198.000 489.400 198.800 489.600 ;
        RECT 198.000 489.000 203.400 489.400 ;
        RECT 198.000 488.800 204.200 489.000 ;
        RECT 202.800 488.200 204.200 488.800 ;
        RECT 196.400 487.600 202.200 488.200 ;
        RECT 205.200 488.000 206.800 488.800 ;
        RECT 205.200 487.600 205.800 488.000 ;
        RECT 193.200 482.200 194.000 487.000 ;
        RECT 196.400 482.200 197.200 487.000 ;
        RECT 201.600 486.800 205.800 487.600 ;
        RECT 207.600 487.400 208.400 493.000 ;
        RECT 210.600 495.200 211.600 496.000 ;
        RECT 210.600 490.800 211.400 495.200 ;
        RECT 212.400 494.600 213.200 499.800 ;
        RECT 218.800 496.600 219.600 499.800 ;
        RECT 220.400 497.000 221.200 499.800 ;
        RECT 222.000 497.000 222.800 499.800 ;
        RECT 223.600 497.000 224.400 499.800 ;
        RECT 225.200 497.000 226.000 499.800 ;
        RECT 228.400 497.000 229.200 499.800 ;
        RECT 231.600 497.000 232.400 499.800 ;
        RECT 233.200 497.000 234.000 499.800 ;
        RECT 234.800 497.000 235.600 499.800 ;
        RECT 217.200 495.800 219.600 496.600 ;
        RECT 236.400 496.600 237.200 499.800 ;
        RECT 217.200 495.200 218.000 495.800 ;
        RECT 212.000 494.000 213.200 494.600 ;
        RECT 216.200 494.600 218.000 495.200 ;
        RECT 222.000 495.600 223.000 496.400 ;
        RECT 226.000 495.600 227.600 496.400 ;
        RECT 228.400 495.800 233.000 496.400 ;
        RECT 236.400 495.800 239.000 496.600 ;
        RECT 228.400 495.600 229.200 495.800 ;
        RECT 212.000 492.000 212.600 494.000 ;
        RECT 216.200 493.400 217.000 494.600 ;
        RECT 213.200 492.600 217.000 493.400 ;
        RECT 222.000 492.800 222.800 495.600 ;
        RECT 228.400 494.800 229.200 495.000 ;
        RECT 224.800 494.200 229.200 494.800 ;
        RECT 224.800 494.000 225.600 494.200 ;
        RECT 230.000 493.600 230.800 495.200 ;
        RECT 232.200 493.400 233.000 495.800 ;
        RECT 238.200 495.200 239.000 495.800 ;
        RECT 238.200 494.400 241.200 495.200 ;
        RECT 242.800 493.800 243.600 499.800 ;
        RECT 244.400 495.200 245.200 499.800 ;
        RECT 247.600 496.400 248.400 499.800 ;
        RECT 247.600 495.800 248.600 496.400 ;
        RECT 244.400 494.600 247.000 495.200 ;
        RECT 225.200 492.600 228.400 493.400 ;
        RECT 232.200 492.600 234.200 493.400 ;
        RECT 234.800 493.000 243.600 493.800 ;
        RECT 218.800 492.000 219.600 492.600 ;
        RECT 236.400 492.000 237.200 492.400 ;
        RECT 238.000 492.000 238.800 492.400 ;
        RECT 241.400 492.000 242.200 492.200 ;
        RECT 212.000 491.400 212.800 492.000 ;
        RECT 218.800 491.400 242.200 492.000 ;
        RECT 210.600 490.000 211.600 490.800 ;
        RECT 209.200 488.300 210.000 488.400 ;
        RECT 210.800 488.300 211.600 490.000 ;
        RECT 209.200 487.700 211.600 488.300 ;
        RECT 209.200 487.600 210.000 487.700 ;
        RECT 206.400 486.800 208.400 487.400 ;
        RECT 198.000 482.200 198.800 485.000 ;
        RECT 199.600 482.200 200.400 485.000 ;
        RECT 202.800 482.200 203.600 486.800 ;
        RECT 206.400 486.200 207.000 486.800 ;
        RECT 206.000 485.600 207.000 486.200 ;
        RECT 206.000 482.200 206.800 485.600 ;
        RECT 210.800 482.200 211.600 487.700 ;
        RECT 212.200 489.600 212.800 491.400 ;
        RECT 212.200 489.000 221.200 489.600 ;
        RECT 212.200 487.400 212.800 489.000 ;
        RECT 220.400 488.800 221.200 489.000 ;
        RECT 223.600 489.000 232.200 489.600 ;
        RECT 223.600 488.800 224.400 489.000 ;
        RECT 215.400 487.600 218.000 488.400 ;
        RECT 212.200 486.800 214.800 487.400 ;
        RECT 214.000 482.200 214.800 486.800 ;
        RECT 217.200 482.200 218.000 487.600 ;
        RECT 218.600 486.800 222.800 487.600 ;
        RECT 220.400 482.200 221.200 485.000 ;
        RECT 222.000 482.200 222.800 485.000 ;
        RECT 223.600 482.200 224.400 485.000 ;
        RECT 225.200 482.200 226.000 488.400 ;
        RECT 228.400 487.600 231.000 488.400 ;
        RECT 231.600 488.200 232.200 489.000 ;
        RECT 233.200 489.400 234.000 489.600 ;
        RECT 233.200 489.000 238.600 489.400 ;
        RECT 233.200 488.800 239.400 489.000 ;
        RECT 238.000 488.200 239.400 488.800 ;
        RECT 231.600 487.600 237.400 488.200 ;
        RECT 240.400 488.000 242.000 488.800 ;
        RECT 240.400 487.600 241.000 488.000 ;
        RECT 228.400 482.200 229.200 487.000 ;
        RECT 231.600 482.200 232.400 487.000 ;
        RECT 236.800 486.800 241.000 487.600 ;
        RECT 242.800 487.400 243.600 493.000 ;
        RECT 244.600 492.400 245.400 493.200 ;
        RECT 244.400 491.600 245.400 492.400 ;
        RECT 246.400 493.000 247.000 494.600 ;
        RECT 248.000 494.400 248.600 495.800 ;
        RECT 252.400 495.200 253.200 499.800 ;
        RECT 255.600 495.200 256.400 499.800 ;
        RECT 258.800 495.200 259.600 499.800 ;
        RECT 262.000 495.200 262.800 499.800 ;
        RECT 266.800 495.200 267.600 499.800 ;
        RECT 270.000 495.200 270.800 499.800 ;
        RECT 273.200 495.200 274.000 499.800 ;
        RECT 276.400 495.200 277.200 499.800 ;
        RECT 279.600 495.800 280.400 499.800 ;
        RECT 281.200 496.000 282.000 499.800 ;
        RECT 284.400 496.000 285.200 499.800 ;
        RECT 288.600 498.400 289.400 499.800 ;
        RECT 288.600 497.600 290.000 498.400 ;
        RECT 288.600 496.400 289.400 497.600 ;
        RECT 281.200 495.800 285.200 496.000 ;
        RECT 287.600 495.800 289.400 496.400 ;
        RECT 290.800 496.000 291.600 499.800 ;
        RECT 294.000 496.000 294.800 499.800 ;
        RECT 290.800 495.800 294.800 496.000 ;
        RECT 247.600 493.600 248.600 494.400 ;
        RECT 246.400 492.200 247.400 493.000 ;
        RECT 246.400 490.200 247.000 492.200 ;
        RECT 248.000 490.200 248.600 493.600 ;
        RECT 250.800 494.400 253.200 495.200 ;
        RECT 254.200 494.400 256.400 495.200 ;
        RECT 257.400 494.400 259.600 495.200 ;
        RECT 261.000 494.400 262.800 495.200 ;
        RECT 265.200 494.400 267.600 495.200 ;
        RECT 268.600 494.400 270.800 495.200 ;
        RECT 271.800 494.400 274.000 495.200 ;
        RECT 275.400 494.400 277.200 495.200 ;
        RECT 279.800 494.400 280.400 495.800 ;
        RECT 281.400 495.400 285.000 495.800 ;
        RECT 283.600 494.400 284.400 494.800 ;
        RECT 250.800 491.600 251.600 494.400 ;
        RECT 254.200 493.800 255.000 494.400 ;
        RECT 257.400 493.800 258.200 494.400 ;
        RECT 261.000 493.800 261.800 494.400 ;
        RECT 263.600 493.800 264.400 494.400 ;
        RECT 252.400 493.000 255.000 493.800 ;
        RECT 255.800 493.000 258.200 493.800 ;
        RECT 259.200 493.000 261.800 493.800 ;
        RECT 262.600 493.000 264.400 493.800 ;
        RECT 254.200 491.600 255.000 493.000 ;
        RECT 257.400 491.600 258.200 493.000 ;
        RECT 261.000 491.600 261.800 493.000 ;
        RECT 265.200 491.600 266.000 494.400 ;
        RECT 268.600 493.800 269.400 494.400 ;
        RECT 271.800 493.800 272.600 494.400 ;
        RECT 275.400 493.800 276.200 494.400 ;
        RECT 278.000 493.800 278.800 494.400 ;
        RECT 266.800 493.000 269.400 493.800 ;
        RECT 270.200 493.000 272.600 493.800 ;
        RECT 273.600 493.000 276.200 493.800 ;
        RECT 277.000 493.000 278.800 493.800 ;
        RECT 279.600 493.600 282.200 494.400 ;
        RECT 283.600 493.800 285.200 494.400 ;
        RECT 284.400 493.600 285.200 493.800 ;
        RECT 286.000 493.600 286.800 495.200 ;
        RECT 268.600 491.600 269.400 493.000 ;
        RECT 271.800 491.600 272.600 493.000 ;
        RECT 275.400 491.600 276.200 493.000 ;
        RECT 250.800 490.800 253.200 491.600 ;
        RECT 254.200 490.800 256.400 491.600 ;
        RECT 257.400 490.800 259.600 491.600 ;
        RECT 261.000 490.800 262.800 491.600 ;
        RECT 265.200 490.800 267.600 491.600 ;
        RECT 268.600 490.800 270.800 491.600 ;
        RECT 271.800 490.800 274.000 491.600 ;
        RECT 275.400 490.800 277.200 491.600 ;
        RECT 241.600 486.800 243.600 487.400 ;
        RECT 244.400 489.600 247.000 490.200 ;
        RECT 233.200 482.200 234.000 485.000 ;
        RECT 234.800 482.200 235.600 485.000 ;
        RECT 238.000 482.200 238.800 486.800 ;
        RECT 241.600 486.200 242.200 486.800 ;
        RECT 241.200 485.600 242.200 486.200 ;
        RECT 241.200 482.200 242.000 485.600 ;
        RECT 244.400 482.200 245.200 489.600 ;
        RECT 247.600 489.200 248.600 490.200 ;
        RECT 247.600 482.200 248.400 489.200 ;
        RECT 252.400 482.200 253.200 490.800 ;
        RECT 255.600 482.200 256.400 490.800 ;
        RECT 258.800 482.200 259.600 490.800 ;
        RECT 262.000 482.200 262.800 490.800 ;
        RECT 266.800 482.200 267.600 490.800 ;
        RECT 270.000 482.200 270.800 490.800 ;
        RECT 273.200 482.200 274.000 490.800 ;
        RECT 276.400 482.200 277.200 490.800 ;
        RECT 279.600 490.200 280.400 490.400 ;
        RECT 281.600 490.200 282.200 493.600 ;
        RECT 282.800 491.600 283.600 493.200 ;
        RECT 279.600 489.600 281.000 490.200 ;
        RECT 281.600 489.600 282.600 490.200 ;
        RECT 280.400 488.400 281.000 489.600 ;
        RECT 280.400 487.600 281.200 488.400 ;
        RECT 281.800 482.200 282.600 489.600 ;
        RECT 287.600 482.200 288.400 495.800 ;
        RECT 291.000 495.400 294.600 495.800 ;
        RECT 295.600 495.600 296.400 499.800 ;
        RECT 297.200 496.000 298.000 499.800 ;
        RECT 300.400 496.000 301.200 499.800 ;
        RECT 297.200 495.800 301.200 496.000 ;
        RECT 302.000 495.800 302.800 499.800 ;
        RECT 312.200 496.000 313.000 499.000 ;
        RECT 316.400 497.000 317.200 499.000 ;
        RECT 291.600 494.400 292.400 494.800 ;
        RECT 295.600 494.400 296.200 495.600 ;
        RECT 297.400 495.400 301.000 495.800 ;
        RECT 298.000 494.400 298.800 494.800 ;
        RECT 302.000 494.400 302.600 495.800 ;
        RECT 311.400 495.400 313.000 496.000 ;
        RECT 311.400 495.000 312.200 495.400 ;
        RECT 311.400 494.400 312.000 495.000 ;
        RECT 316.600 494.800 317.200 497.000 ;
        RECT 319.600 496.400 320.400 499.800 ;
        RECT 290.800 493.800 292.400 494.400 ;
        RECT 290.800 493.600 291.600 493.800 ;
        RECT 293.800 493.600 296.400 494.400 ;
        RECT 297.200 493.800 298.800 494.400 ;
        RECT 297.200 493.600 298.000 493.800 ;
        RECT 300.200 493.600 302.800 494.400 ;
        RECT 310.000 493.600 312.000 494.400 ;
        RECT 313.000 494.200 317.200 494.800 ;
        RECT 319.400 495.600 320.400 496.400 ;
        RECT 319.400 494.400 320.000 495.600 ;
        RECT 322.800 495.200 323.600 499.800 ;
        RECT 324.400 496.000 325.200 499.800 ;
        RECT 327.600 496.000 328.400 499.800 ;
        RECT 324.400 495.800 328.400 496.000 ;
        RECT 329.200 495.800 330.000 499.800 ;
        RECT 332.400 497.800 333.200 499.800 ;
        RECT 324.600 495.400 328.200 495.800 ;
        RECT 321.000 494.600 323.600 495.200 ;
        RECT 313.000 493.800 314.000 494.200 ;
        RECT 292.400 491.600 293.200 493.200 ;
        RECT 289.200 488.800 290.000 490.400 ;
        RECT 293.800 490.200 294.400 493.600 ;
        RECT 298.800 491.600 299.600 493.200 ;
        RECT 295.600 490.200 296.400 490.400 ;
        RECT 300.200 490.200 300.800 493.600 ;
        RECT 311.400 492.400 312.000 493.600 ;
        RECT 312.600 493.000 314.000 493.800 ;
        RECT 319.400 493.600 320.400 494.400 ;
        RECT 310.000 490.800 310.800 492.400 ;
        RECT 311.400 491.600 312.400 492.400 ;
        RECT 302.000 490.200 302.800 490.400 ;
        RECT 293.400 489.600 294.400 490.200 ;
        RECT 295.000 489.600 296.400 490.200 ;
        RECT 299.800 489.600 300.800 490.200 ;
        RECT 301.400 489.600 302.800 490.200 ;
        RECT 311.400 489.800 312.000 491.600 ;
        RECT 313.400 491.000 314.000 493.000 ;
        RECT 314.800 491.600 315.600 493.200 ;
        RECT 316.400 492.300 317.200 493.200 ;
        RECT 318.000 492.300 318.800 492.400 ;
        RECT 316.400 491.700 318.800 492.300 ;
        RECT 316.400 491.600 317.200 491.700 ;
        RECT 318.000 491.600 318.800 491.700 ;
        RECT 313.400 490.400 317.200 491.000 ;
        RECT 293.400 482.200 294.200 489.600 ;
        RECT 295.000 488.400 295.600 489.600 ;
        RECT 294.800 487.600 295.600 488.400 ;
        RECT 299.800 484.400 300.600 489.600 ;
        RECT 301.400 488.400 302.000 489.600 ;
        RECT 311.400 489.200 313.000 489.800 ;
        RECT 301.200 487.600 302.000 488.400 ;
        RECT 298.800 483.600 300.600 484.400 ;
        RECT 299.800 482.200 300.600 483.600 ;
        RECT 312.200 482.200 313.000 489.200 ;
        RECT 316.600 487.000 317.200 490.400 ;
        RECT 319.400 490.200 320.000 493.600 ;
        RECT 321.000 493.000 321.600 494.600 ;
        RECT 325.200 494.400 326.000 494.800 ;
        RECT 329.200 494.400 329.800 495.800 ;
        RECT 330.800 495.600 331.600 497.200 ;
        RECT 332.600 494.400 333.200 497.800 ;
        RECT 335.600 495.200 336.400 499.800 ;
        RECT 338.800 496.400 339.600 499.800 ;
        RECT 338.800 495.800 339.800 496.400 ;
        RECT 342.000 495.800 342.800 499.800 ;
        RECT 343.600 496.000 344.400 499.800 ;
        RECT 346.800 496.000 347.600 499.800 ;
        RECT 352.200 496.000 353.000 499.000 ;
        RECT 356.400 497.000 357.200 499.000 ;
        RECT 343.600 495.800 347.600 496.000 ;
        RECT 335.600 494.600 338.200 495.200 ;
        RECT 324.400 493.800 326.000 494.400 ;
        RECT 324.400 493.600 325.200 493.800 ;
        RECT 327.400 493.600 330.000 494.400 ;
        RECT 332.400 493.600 333.200 494.400 ;
        RECT 320.600 492.200 321.600 493.000 ;
        RECT 321.000 490.200 321.600 492.200 ;
        RECT 322.600 492.400 323.400 493.200 ;
        RECT 322.600 491.600 323.600 492.400 ;
        RECT 326.000 491.600 326.800 493.200 ;
        RECT 327.400 490.200 328.000 493.600 ;
        RECT 332.600 492.400 333.200 493.600 ;
        RECT 335.800 492.400 336.600 493.200 ;
        RECT 332.400 491.600 333.200 492.400 ;
        RECT 329.200 490.200 330.000 490.400 ;
        RECT 332.600 490.200 333.200 491.600 ;
        RECT 334.000 490.800 334.800 492.400 ;
        RECT 335.600 491.600 336.600 492.400 ;
        RECT 337.600 493.000 338.200 494.600 ;
        RECT 339.200 494.400 339.800 495.800 ;
        RECT 342.200 494.400 342.800 495.800 ;
        RECT 343.800 495.400 347.400 495.800 ;
        RECT 351.400 495.400 353.000 496.000 ;
        RECT 351.400 495.000 352.200 495.400 ;
        RECT 346.000 494.400 346.800 494.800 ;
        RECT 351.400 494.400 352.000 495.000 ;
        RECT 356.600 494.800 357.200 497.000 ;
        RECT 358.000 496.000 358.800 499.800 ;
        RECT 361.200 496.000 362.000 499.800 ;
        RECT 358.000 495.800 362.000 496.000 ;
        RECT 362.800 495.800 363.600 499.800 ;
        RECT 364.400 495.800 365.200 499.800 ;
        RECT 366.000 496.000 366.800 499.800 ;
        RECT 369.200 496.000 370.000 499.800 ;
        RECT 374.600 496.000 375.400 499.000 ;
        RECT 378.800 497.000 379.600 499.000 ;
        RECT 366.000 495.800 370.000 496.000 ;
        RECT 358.200 495.400 361.800 495.800 ;
        RECT 338.800 494.300 339.800 494.400 ;
        RECT 340.400 494.300 341.200 494.400 ;
        RECT 338.800 493.700 341.200 494.300 ;
        RECT 338.800 493.600 339.800 493.700 ;
        RECT 340.400 493.600 341.200 493.700 ;
        RECT 342.000 493.600 344.600 494.400 ;
        RECT 346.000 493.800 347.600 494.400 ;
        RECT 346.800 493.600 347.600 493.800 ;
        RECT 350.000 493.600 352.000 494.400 ;
        RECT 353.000 494.200 357.200 494.800 ;
        RECT 358.800 494.400 359.600 494.800 ;
        RECT 362.800 494.400 363.400 495.800 ;
        RECT 364.600 494.400 365.200 495.800 ;
        RECT 366.200 495.400 369.800 495.800 ;
        RECT 373.800 495.400 375.400 496.000 ;
        RECT 373.800 495.000 374.600 495.400 ;
        RECT 368.400 494.400 369.200 494.800 ;
        RECT 373.800 494.400 374.400 495.000 ;
        RECT 379.000 494.800 379.600 497.000 ;
        RECT 353.000 493.800 354.000 494.200 ;
        RECT 337.600 492.200 338.600 493.000 ;
        RECT 337.600 490.200 338.200 492.200 ;
        RECT 339.200 490.200 339.800 493.600 ;
        RECT 319.400 489.200 320.400 490.200 ;
        RECT 321.000 489.600 323.600 490.200 ;
        RECT 316.400 483.000 317.200 487.000 ;
        RECT 319.600 482.200 320.400 489.200 ;
        RECT 322.800 482.200 323.600 489.600 ;
        RECT 327.000 489.600 328.000 490.200 ;
        RECT 328.600 489.600 330.000 490.200 ;
        RECT 327.000 482.200 327.800 489.600 ;
        RECT 328.600 488.400 329.200 489.600 ;
        RECT 332.400 489.400 334.200 490.200 ;
        RECT 328.400 487.600 329.200 488.400 ;
        RECT 333.400 482.200 334.200 489.400 ;
        RECT 335.600 489.600 338.200 490.200 ;
        RECT 335.600 482.200 336.400 489.600 ;
        RECT 338.800 489.200 339.800 490.200 ;
        RECT 342.000 490.200 342.800 490.400 ;
        RECT 344.000 490.200 344.600 493.600 ;
        RECT 345.200 491.600 346.000 493.200 ;
        RECT 351.400 492.400 352.000 493.600 ;
        RECT 352.600 493.000 354.000 493.800 ;
        RECT 358.000 493.800 359.600 494.400 ;
        RECT 358.000 493.600 358.800 493.800 ;
        RECT 361.000 493.600 363.600 494.400 ;
        RECT 364.400 493.600 367.000 494.400 ;
        RECT 368.400 493.800 370.000 494.400 ;
        RECT 369.200 493.600 370.000 493.800 ;
        RECT 372.400 493.600 374.400 494.400 ;
        RECT 375.400 494.200 379.600 494.800 ;
        RECT 380.400 495.400 381.200 499.800 ;
        RECT 384.600 498.400 385.800 499.800 ;
        RECT 384.600 497.800 386.000 498.400 ;
        RECT 389.200 497.800 390.000 499.800 ;
        RECT 393.600 498.400 394.400 499.800 ;
        RECT 393.600 497.800 395.600 498.400 ;
        RECT 385.200 497.000 386.000 497.800 ;
        RECT 389.400 497.200 390.000 497.800 ;
        RECT 389.400 496.600 392.200 497.200 ;
        RECT 391.400 496.400 392.200 496.600 ;
        RECT 393.200 495.600 394.000 497.200 ;
        RECT 394.800 497.000 395.600 497.800 ;
        RECT 383.400 495.400 384.200 495.600 ;
        RECT 380.400 494.800 384.200 495.400 ;
        RECT 375.400 493.800 376.400 494.200 ;
        RECT 348.400 492.300 349.200 492.400 ;
        RECT 350.000 492.300 350.800 492.400 ;
        RECT 348.400 491.700 350.800 492.300 ;
        RECT 348.400 491.600 349.200 491.700 ;
        RECT 350.000 490.800 350.800 491.700 ;
        RECT 351.400 491.600 352.400 492.400 ;
        RECT 342.000 489.600 343.400 490.200 ;
        RECT 344.000 489.600 345.000 490.200 ;
        RECT 338.800 482.200 339.600 489.200 ;
        RECT 342.800 488.400 343.400 489.600 ;
        RECT 344.200 488.400 345.000 489.600 ;
        RECT 351.400 489.800 352.000 491.600 ;
        RECT 353.400 491.000 354.000 493.000 ;
        RECT 354.800 491.600 355.600 493.200 ;
        RECT 356.400 491.600 357.200 493.200 ;
        RECT 359.600 491.600 360.400 493.200 ;
        RECT 353.400 490.400 357.200 491.000 ;
        RECT 351.400 489.200 353.000 489.800 ;
        RECT 342.800 487.600 343.600 488.400 ;
        RECT 344.200 487.600 346.000 488.400 ;
        RECT 344.200 482.200 345.000 487.600 ;
        RECT 352.200 482.200 353.000 489.200 ;
        RECT 356.600 487.000 357.200 490.400 ;
        RECT 361.000 490.200 361.600 493.600 ;
        RECT 366.400 492.300 367.000 493.600 ;
        RECT 362.900 491.700 367.000 492.300 ;
        RECT 362.900 490.400 363.500 491.700 ;
        RECT 362.800 490.200 363.600 490.400 ;
        RECT 356.400 483.000 357.200 487.000 ;
        RECT 360.600 489.600 361.600 490.200 ;
        RECT 362.200 489.600 363.600 490.200 ;
        RECT 364.400 490.200 365.200 490.400 ;
        RECT 366.400 490.200 367.000 491.700 ;
        RECT 367.600 491.600 368.400 493.200 ;
        RECT 373.800 492.400 374.400 493.600 ;
        RECT 375.000 493.000 376.400 493.800 ;
        RECT 370.800 492.300 371.600 492.400 ;
        RECT 372.400 492.300 373.200 492.400 ;
        RECT 370.800 491.700 373.200 492.300 ;
        RECT 370.800 491.600 371.600 491.700 ;
        RECT 372.400 490.800 373.200 491.700 ;
        RECT 373.800 491.600 374.800 492.400 ;
        RECT 364.400 489.600 365.800 490.200 ;
        RECT 366.400 489.600 367.400 490.200 ;
        RECT 360.600 484.400 361.400 489.600 ;
        RECT 362.200 488.400 362.800 489.600 ;
        RECT 362.000 487.600 362.800 488.400 ;
        RECT 365.200 488.400 365.800 489.600 ;
        RECT 365.200 487.600 366.000 488.400 ;
        RECT 359.600 483.600 361.400 484.400 ;
        RECT 360.600 482.200 361.400 483.600 ;
        RECT 366.600 482.200 367.400 489.600 ;
        RECT 373.800 489.800 374.400 491.600 ;
        RECT 375.800 491.000 376.400 493.000 ;
        RECT 377.200 491.600 378.000 493.200 ;
        RECT 378.800 491.600 379.600 493.200 ;
        RECT 380.400 491.400 381.200 494.800 ;
        RECT 387.400 494.200 388.200 494.400 ;
        RECT 393.200 494.200 393.800 495.600 ;
        RECT 398.000 495.000 398.800 499.800 ;
        RECT 399.600 496.000 400.400 499.800 ;
        RECT 402.800 496.000 403.600 499.800 ;
        RECT 399.600 495.800 403.600 496.000 ;
        RECT 404.400 495.800 405.200 499.800 ;
        RECT 406.000 495.800 406.800 499.800 ;
        RECT 407.600 496.000 408.400 499.800 ;
        RECT 410.800 496.000 411.600 499.800 ;
        RECT 407.600 495.800 411.600 496.000 ;
        RECT 399.800 495.400 403.400 495.800 ;
        RECT 400.400 494.400 401.200 494.800 ;
        RECT 404.400 494.400 405.000 495.800 ;
        RECT 406.200 494.400 406.800 495.800 ;
        RECT 407.800 495.400 411.400 495.800 ;
        RECT 412.400 495.000 413.200 499.800 ;
        RECT 416.800 498.400 417.600 499.800 ;
        RECT 415.600 497.800 417.600 498.400 ;
        RECT 421.200 497.800 422.000 499.800 ;
        RECT 425.400 498.400 426.600 499.800 ;
        RECT 425.200 497.800 426.600 498.400 ;
        RECT 415.600 497.000 416.400 497.800 ;
        RECT 421.200 497.200 421.800 497.800 ;
        RECT 417.200 496.400 418.000 497.200 ;
        RECT 419.000 496.600 421.800 497.200 ;
        RECT 425.200 497.000 426.000 497.800 ;
        RECT 419.000 496.400 419.800 496.600 ;
        RECT 410.000 494.400 410.800 494.800 ;
        RECT 396.400 494.200 398.000 494.400 ;
        RECT 387.000 493.600 398.000 494.200 ;
        RECT 399.600 493.800 401.200 494.400 ;
        RECT 399.600 493.600 400.400 493.800 ;
        RECT 402.600 493.600 405.200 494.400 ;
        RECT 406.000 493.600 408.600 494.400 ;
        RECT 410.000 493.800 411.600 494.400 ;
        RECT 410.800 493.600 411.600 493.800 ;
        RECT 413.200 494.200 414.800 494.400 ;
        RECT 417.400 494.200 418.000 496.400 ;
        RECT 427.000 495.400 427.800 495.600 ;
        RECT 430.000 495.400 430.800 499.800 ;
        RECT 435.400 498.400 436.200 499.000 ;
        RECT 434.800 497.600 436.200 498.400 ;
        RECT 435.400 496.000 436.200 497.600 ;
        RECT 439.600 497.000 440.400 499.000 ;
        RECT 427.000 494.800 430.800 495.400 ;
        RECT 418.800 494.200 419.600 494.400 ;
        RECT 423.000 494.200 423.800 494.400 ;
        RECT 413.200 493.600 424.200 494.200 ;
        RECT 385.200 492.800 386.000 493.000 ;
        RECT 382.200 492.200 386.000 492.800 ;
        RECT 382.200 492.000 383.000 492.200 ;
        RECT 383.800 491.400 384.600 491.600 ;
        RECT 375.800 490.400 379.600 491.000 ;
        RECT 373.800 489.200 375.400 489.800 ;
        RECT 374.600 482.200 375.400 489.200 ;
        RECT 379.000 487.000 379.600 490.400 ;
        RECT 378.800 483.000 379.600 487.000 ;
        RECT 380.400 490.800 384.600 491.400 ;
        RECT 380.400 482.200 381.200 490.800 ;
        RECT 387.000 490.400 387.600 493.600 ;
        RECT 394.200 493.400 395.000 493.600 ;
        RECT 395.800 492.400 396.600 492.600 ;
        RECT 391.600 491.800 396.600 492.400 ;
        RECT 391.600 491.600 392.400 491.800 ;
        RECT 401.200 491.600 402.000 493.200 ;
        RECT 393.200 491.000 398.800 491.200 ;
        RECT 393.000 490.800 398.800 491.000 ;
        RECT 385.200 489.800 387.600 490.400 ;
        RECT 389.000 490.600 398.800 490.800 ;
        RECT 389.000 490.200 393.800 490.600 ;
        RECT 385.200 488.800 385.800 489.800 ;
        RECT 384.400 488.000 385.800 488.800 ;
        RECT 387.400 489.000 388.200 489.200 ;
        RECT 389.000 489.000 389.600 490.200 ;
        RECT 387.400 488.400 389.600 489.000 ;
        RECT 390.200 489.000 395.600 489.600 ;
        RECT 390.200 488.800 391.000 489.000 ;
        RECT 394.800 488.800 395.600 489.000 ;
        RECT 388.600 487.400 389.400 487.600 ;
        RECT 391.400 487.400 392.200 487.600 ;
        RECT 385.200 486.200 386.000 487.000 ;
        RECT 388.600 486.800 392.200 487.400 ;
        RECT 389.400 486.200 390.000 486.800 ;
        RECT 394.800 486.200 395.600 487.000 ;
        RECT 384.600 482.200 385.800 486.200 ;
        RECT 389.200 482.200 390.000 486.200 ;
        RECT 393.600 485.600 395.600 486.200 ;
        RECT 393.600 482.200 394.400 485.600 ;
        RECT 398.000 482.200 398.800 490.600 ;
        RECT 402.600 490.200 403.200 493.600 ;
        RECT 408.000 492.300 408.600 493.600 ;
        RECT 416.200 493.400 417.000 493.600 ;
        RECT 404.500 491.700 408.600 492.300 ;
        RECT 404.500 490.400 405.100 491.700 ;
        RECT 404.400 490.200 405.200 490.400 ;
        RECT 402.200 489.600 403.200 490.200 ;
        RECT 403.800 489.600 405.200 490.200 ;
        RECT 406.000 490.200 406.800 490.400 ;
        RECT 408.000 490.200 408.600 491.700 ;
        RECT 409.200 491.600 410.000 493.200 ;
        RECT 414.600 492.400 415.400 492.600 ;
        RECT 414.600 492.300 419.600 492.400 ;
        RECT 420.400 492.300 421.200 492.400 ;
        RECT 414.600 491.800 421.200 492.300 ;
        RECT 418.800 491.700 421.200 491.800 ;
        RECT 418.800 491.600 419.600 491.700 ;
        RECT 420.400 491.600 421.200 491.700 ;
        RECT 412.400 491.000 418.000 491.200 ;
        RECT 412.400 490.800 418.200 491.000 ;
        RECT 412.400 490.600 422.200 490.800 ;
        RECT 406.000 489.600 407.400 490.200 ;
        RECT 408.000 489.600 409.000 490.200 ;
        RECT 402.200 482.200 403.000 489.600 ;
        RECT 403.800 488.400 404.400 489.600 ;
        RECT 403.600 487.600 404.400 488.400 ;
        RECT 406.800 488.400 407.400 489.600 ;
        RECT 406.800 487.600 407.600 488.400 ;
        RECT 408.200 482.200 409.000 489.600 ;
        RECT 412.400 482.200 413.200 490.600 ;
        RECT 417.400 490.200 422.200 490.600 ;
        RECT 415.600 489.000 421.000 489.600 ;
        RECT 415.600 488.800 416.400 489.000 ;
        RECT 420.200 488.800 421.000 489.000 ;
        RECT 421.600 489.000 422.200 490.200 ;
        RECT 423.600 490.400 424.200 493.600 ;
        RECT 425.200 492.800 426.000 493.000 ;
        RECT 425.200 492.200 429.000 492.800 ;
        RECT 428.200 492.000 429.000 492.200 ;
        RECT 426.600 491.400 427.400 491.600 ;
        RECT 430.000 491.400 430.800 494.800 ;
        RECT 434.600 495.400 436.200 496.000 ;
        RECT 434.600 495.000 435.400 495.400 ;
        RECT 434.600 494.400 435.200 495.000 ;
        RECT 439.800 494.800 440.400 497.000 ;
        RECT 441.200 496.000 442.000 499.800 ;
        RECT 444.400 496.000 445.200 499.800 ;
        RECT 441.200 495.800 445.200 496.000 ;
        RECT 446.000 495.800 446.800 499.800 ;
        RECT 441.400 495.400 445.000 495.800 ;
        RECT 433.200 493.600 435.200 494.400 ;
        RECT 436.200 494.200 440.400 494.800 ;
        RECT 442.000 494.400 442.800 494.800 ;
        RECT 446.000 494.400 446.600 495.800 ;
        RECT 447.600 495.600 448.400 499.800 ;
        RECT 449.200 496.000 450.000 499.800 ;
        RECT 452.400 496.000 453.200 499.800 ;
        RECT 449.200 495.800 453.200 496.000 ;
        RECT 454.000 496.000 454.800 499.800 ;
        RECT 457.200 496.000 458.000 499.800 ;
        RECT 454.000 495.800 458.000 496.000 ;
        RECT 458.800 495.800 459.600 499.800 ;
        RECT 465.200 496.000 466.000 499.800 ;
        RECT 468.400 496.000 469.200 499.800 ;
        RECT 465.200 495.800 469.200 496.000 ;
        RECT 470.000 495.800 470.800 499.800 ;
        RECT 447.800 494.400 448.400 495.600 ;
        RECT 449.400 495.400 453.000 495.800 ;
        RECT 454.200 495.400 457.800 495.800 ;
        RECT 451.600 494.400 452.400 494.800 ;
        RECT 454.800 494.400 455.600 494.800 ;
        RECT 458.800 494.400 459.400 495.800 ;
        RECT 465.400 495.400 469.000 495.800 ;
        RECT 466.000 494.400 466.800 494.800 ;
        RECT 470.000 494.400 470.600 495.800 ;
        RECT 471.600 495.600 472.400 499.800 ;
        RECT 473.200 496.000 474.000 499.800 ;
        RECT 476.400 496.000 477.200 499.800 ;
        RECT 473.200 495.800 477.200 496.000 ;
        RECT 471.800 494.400 472.400 495.600 ;
        RECT 473.400 495.400 477.000 495.800 ;
        RECT 478.000 495.400 478.800 499.800 ;
        RECT 482.200 498.400 483.400 499.800 ;
        RECT 482.200 497.800 483.600 498.400 ;
        RECT 486.800 497.800 487.600 499.800 ;
        RECT 491.200 498.400 492.000 499.800 ;
        RECT 491.200 497.800 493.200 498.400 ;
        RECT 482.800 497.000 483.600 497.800 ;
        RECT 487.000 497.200 487.600 497.800 ;
        RECT 487.000 496.600 489.800 497.200 ;
        RECT 489.000 496.400 489.800 496.600 ;
        RECT 490.800 495.600 491.600 497.200 ;
        RECT 492.400 497.000 493.200 497.800 ;
        RECT 481.000 495.400 481.800 495.600 ;
        RECT 478.000 494.800 481.800 495.400 ;
        RECT 475.600 494.400 476.400 494.800 ;
        RECT 436.200 493.800 437.200 494.200 ;
        RECT 426.600 490.800 430.800 491.400 ;
        RECT 433.200 490.800 434.000 492.400 ;
        RECT 423.600 489.800 426.000 490.400 ;
        RECT 423.000 489.000 423.800 489.200 ;
        RECT 421.600 488.400 423.800 489.000 ;
        RECT 425.400 488.800 426.000 489.800 ;
        RECT 425.400 488.000 426.800 488.800 ;
        RECT 419.000 487.400 419.800 487.600 ;
        RECT 421.800 487.400 422.600 487.600 ;
        RECT 415.600 486.200 416.400 487.000 ;
        RECT 419.000 486.800 422.600 487.400 ;
        RECT 421.200 486.200 421.800 486.800 ;
        RECT 425.200 486.200 426.000 487.000 ;
        RECT 415.600 485.600 417.600 486.200 ;
        RECT 416.800 482.200 417.600 485.600 ;
        RECT 421.200 482.200 422.000 486.200 ;
        RECT 425.400 482.200 426.600 486.200 ;
        RECT 430.000 482.200 430.800 490.800 ;
        RECT 434.600 489.800 435.200 493.600 ;
        RECT 435.800 493.000 437.200 493.800 ;
        RECT 441.200 493.800 442.800 494.400 ;
        RECT 441.200 493.600 442.000 493.800 ;
        RECT 444.200 493.600 446.800 494.400 ;
        RECT 447.600 493.600 450.200 494.400 ;
        RECT 451.600 493.800 453.200 494.400 ;
        RECT 452.400 493.600 453.200 493.800 ;
        RECT 454.000 493.800 455.600 494.400 ;
        RECT 454.000 493.600 454.800 493.800 ;
        RECT 457.000 493.600 459.600 494.400 ;
        RECT 465.200 493.800 466.800 494.400 ;
        RECT 465.200 493.600 466.000 493.800 ;
        RECT 468.200 493.600 470.800 494.400 ;
        RECT 471.600 493.600 474.200 494.400 ;
        RECT 475.600 493.800 477.200 494.400 ;
        RECT 476.400 493.600 477.200 493.800 ;
        RECT 436.600 491.000 437.200 493.000 ;
        RECT 438.000 491.600 438.800 493.200 ;
        RECT 439.600 491.600 440.400 493.200 ;
        RECT 442.800 491.600 443.600 493.200 ;
        RECT 444.200 492.300 444.800 493.600 ;
        RECT 444.200 491.700 448.300 492.300 ;
        RECT 436.600 490.400 440.400 491.000 ;
        RECT 434.600 489.200 436.200 489.800 ;
        RECT 435.400 482.200 436.200 489.200 ;
        RECT 439.800 487.000 440.400 490.400 ;
        RECT 444.200 490.200 444.800 491.700 ;
        RECT 447.700 490.400 448.300 491.700 ;
        RECT 446.000 490.200 446.800 490.400 ;
        RECT 439.600 483.000 440.400 487.000 ;
        RECT 443.800 489.600 444.800 490.200 ;
        RECT 445.400 489.600 446.800 490.200 ;
        RECT 447.600 490.200 448.400 490.400 ;
        RECT 449.600 490.200 450.200 493.600 ;
        RECT 450.800 492.300 451.600 493.200 ;
        RECT 452.400 492.300 453.200 492.400 ;
        RECT 450.800 491.700 453.200 492.300 ;
        RECT 450.800 491.600 451.600 491.700 ;
        RECT 452.400 491.600 453.200 491.700 ;
        RECT 454.000 492.300 454.800 492.400 ;
        RECT 455.600 492.300 456.400 493.200 ;
        RECT 454.000 491.700 456.400 492.300 ;
        RECT 454.000 491.600 454.800 491.700 ;
        RECT 455.600 491.600 456.400 491.700 ;
        RECT 457.000 490.200 457.600 493.600 ;
        RECT 466.800 491.600 467.600 493.200 ;
        RECT 468.200 492.300 468.800 493.600 ;
        RECT 468.200 491.700 472.300 492.300 ;
        RECT 458.800 490.300 459.600 490.400 ;
        RECT 463.600 490.300 464.400 490.400 ;
        RECT 458.800 490.200 464.400 490.300 ;
        RECT 468.200 490.200 468.800 491.700 ;
        RECT 471.700 490.400 472.300 491.700 ;
        RECT 470.000 490.200 470.800 490.400 ;
        RECT 447.600 489.600 449.000 490.200 ;
        RECT 449.600 489.600 450.600 490.200 ;
        RECT 443.800 482.200 444.600 489.600 ;
        RECT 445.400 488.400 446.000 489.600 ;
        RECT 445.200 487.600 446.000 488.400 ;
        RECT 448.400 488.400 449.000 489.600 ;
        RECT 448.400 487.600 449.200 488.400 ;
        RECT 449.800 482.200 450.600 489.600 ;
        RECT 456.600 489.600 457.600 490.200 ;
        RECT 458.200 489.700 464.400 490.200 ;
        RECT 458.200 489.600 459.600 489.700 ;
        RECT 463.600 489.600 464.400 489.700 ;
        RECT 467.800 489.600 468.800 490.200 ;
        RECT 469.400 489.600 470.800 490.200 ;
        RECT 471.600 490.200 472.400 490.400 ;
        RECT 473.600 490.200 474.200 493.600 ;
        RECT 474.800 491.600 475.600 493.200 ;
        RECT 478.000 491.400 478.800 494.800 ;
        RECT 485.000 494.200 485.800 494.400 ;
        RECT 490.800 494.200 491.400 495.600 ;
        RECT 495.600 495.000 496.400 499.800 ;
        RECT 497.200 497.000 498.000 499.000 ;
        RECT 497.200 494.800 497.800 497.000 ;
        RECT 501.400 496.000 502.200 499.000 ;
        RECT 506.800 496.000 507.600 499.800 ;
        RECT 510.000 496.000 510.800 499.800 ;
        RECT 501.400 495.400 503.000 496.000 ;
        RECT 506.800 495.800 510.800 496.000 ;
        RECT 507.000 495.400 510.600 495.800 ;
        RECT 511.600 495.600 512.400 499.800 ;
        RECT 513.200 495.800 514.000 499.800 ;
        RECT 514.800 496.000 515.600 499.800 ;
        RECT 518.000 496.000 518.800 499.800 ;
        RECT 514.800 495.800 518.800 496.000 ;
        RECT 502.200 495.000 503.000 495.400 ;
        RECT 494.000 494.200 495.600 494.400 ;
        RECT 497.200 494.200 501.400 494.800 ;
        RECT 484.600 493.600 495.600 494.200 ;
        RECT 500.400 493.800 501.400 494.200 ;
        RECT 502.400 494.400 503.000 495.000 ;
        RECT 507.600 494.400 508.400 494.800 ;
        RECT 511.600 494.400 512.200 495.600 ;
        RECT 513.400 494.400 514.000 495.800 ;
        RECT 515.000 495.400 518.600 495.800 ;
        RECT 519.600 495.400 520.400 499.800 ;
        RECT 523.800 498.400 525.000 499.800 ;
        RECT 523.800 497.800 525.200 498.400 ;
        RECT 528.400 497.800 529.200 499.800 ;
        RECT 532.800 498.400 533.600 499.800 ;
        RECT 532.800 497.800 534.800 498.400 ;
        RECT 524.400 497.000 525.200 497.800 ;
        RECT 528.600 497.200 529.200 497.800 ;
        RECT 528.600 496.600 531.400 497.200 ;
        RECT 530.600 496.400 531.400 496.600 ;
        RECT 532.400 495.600 533.200 497.200 ;
        RECT 534.000 497.000 534.800 497.800 ;
        RECT 522.600 495.400 523.400 495.600 ;
        RECT 519.600 494.800 523.400 495.400 ;
        RECT 517.200 494.400 518.000 494.800 ;
        RECT 502.400 494.300 504.400 494.400 ;
        RECT 482.800 492.800 483.600 493.000 ;
        RECT 479.800 492.200 483.600 492.800 ;
        RECT 479.800 492.000 480.600 492.200 ;
        RECT 481.400 491.400 482.200 491.600 ;
        RECT 478.000 490.800 482.200 491.400 ;
        RECT 471.600 489.600 473.000 490.200 ;
        RECT 473.600 489.600 474.600 490.200 ;
        RECT 456.600 484.400 457.400 489.600 ;
        RECT 458.200 488.400 458.800 489.600 ;
        RECT 458.000 487.600 458.800 488.400 ;
        RECT 455.600 483.600 457.400 484.400 ;
        RECT 456.600 482.200 457.400 483.600 ;
        RECT 467.800 482.200 468.600 489.600 ;
        RECT 469.400 488.400 470.000 489.600 ;
        RECT 469.200 487.600 470.000 488.400 ;
        RECT 472.400 488.400 473.000 489.600 ;
        RECT 472.400 487.600 473.200 488.400 ;
        RECT 473.800 482.200 474.600 489.600 ;
        RECT 478.000 482.200 478.800 490.800 ;
        RECT 484.600 490.400 485.200 493.600 ;
        RECT 491.800 493.400 492.600 493.600 ;
        RECT 493.400 492.400 494.200 492.600 ;
        RECT 489.200 491.800 494.200 492.400 ;
        RECT 489.200 491.600 490.000 491.800 ;
        RECT 497.200 491.600 498.000 493.200 ;
        RECT 498.800 491.600 499.600 493.200 ;
        RECT 500.400 493.000 501.800 493.800 ;
        RECT 502.400 493.700 505.900 494.300 ;
        RECT 502.400 493.600 504.400 493.700 ;
        RECT 490.800 491.000 496.400 491.200 ;
        RECT 500.400 491.000 501.000 493.000 ;
        RECT 490.600 490.800 496.400 491.000 ;
        RECT 482.800 489.800 485.200 490.400 ;
        RECT 486.600 490.600 496.400 490.800 ;
        RECT 486.600 490.200 491.400 490.600 ;
        RECT 482.800 488.800 483.400 489.800 ;
        RECT 482.000 488.000 483.400 488.800 ;
        RECT 485.000 489.000 485.800 489.200 ;
        RECT 486.600 489.000 487.200 490.200 ;
        RECT 485.000 488.400 487.200 489.000 ;
        RECT 487.800 489.000 493.200 489.600 ;
        RECT 487.800 488.800 488.600 489.000 ;
        RECT 492.400 488.800 493.200 489.000 ;
        RECT 486.200 487.400 487.000 487.600 ;
        RECT 489.000 487.400 489.800 487.600 ;
        RECT 482.800 486.200 483.600 487.000 ;
        RECT 486.200 486.800 489.800 487.400 ;
        RECT 487.000 486.200 487.600 486.800 ;
        RECT 492.400 486.200 493.200 487.000 ;
        RECT 482.200 482.200 483.400 486.200 ;
        RECT 486.800 482.200 487.600 486.200 ;
        RECT 491.200 485.600 493.200 486.200 ;
        RECT 491.200 482.200 492.000 485.600 ;
        RECT 495.600 482.200 496.400 490.600 ;
        RECT 497.200 490.400 501.000 491.000 ;
        RECT 497.200 487.000 497.800 490.400 ;
        RECT 502.400 489.800 503.000 493.600 ;
        RECT 503.600 490.800 504.400 492.400 ;
        RECT 505.300 492.300 505.900 493.700 ;
        RECT 506.800 493.800 508.400 494.400 ;
        RECT 506.800 493.600 507.600 493.800 ;
        RECT 509.800 493.600 512.400 494.400 ;
        RECT 513.200 493.600 515.800 494.400 ;
        RECT 517.200 493.800 518.800 494.400 ;
        RECT 518.000 493.600 518.800 493.800 ;
        RECT 508.400 492.300 509.200 493.200 ;
        RECT 505.300 491.700 509.200 492.300 ;
        RECT 508.400 491.600 509.200 491.700 ;
        RECT 509.800 490.200 510.400 493.600 ;
        RECT 515.200 492.300 515.800 493.600 ;
        RECT 511.700 491.700 515.800 492.300 ;
        RECT 511.700 490.400 512.300 491.700 ;
        RECT 511.600 490.200 512.400 490.400 ;
        RECT 501.400 489.200 503.000 489.800 ;
        RECT 509.400 489.600 510.400 490.200 ;
        RECT 511.000 489.600 512.400 490.200 ;
        RECT 513.200 490.200 514.000 490.400 ;
        RECT 515.200 490.200 515.800 491.700 ;
        RECT 516.400 491.600 517.200 493.200 ;
        RECT 519.600 491.400 520.400 494.800 ;
        RECT 526.600 494.200 527.400 494.400 ;
        RECT 532.400 494.200 533.000 495.600 ;
        RECT 537.200 495.000 538.000 499.800 ;
        RECT 538.800 496.000 539.600 499.800 ;
        RECT 542.000 496.000 542.800 499.800 ;
        RECT 538.800 495.800 542.800 496.000 ;
        RECT 539.000 495.400 542.600 495.800 ;
        RECT 543.600 495.600 544.400 499.800 ;
        RECT 545.200 496.000 546.000 499.800 ;
        RECT 548.400 496.000 549.200 499.800 ;
        RECT 545.200 495.800 549.200 496.000 ;
        RECT 550.000 495.800 550.800 499.800 ;
        RECT 539.600 494.400 540.400 494.800 ;
        RECT 543.600 494.400 544.200 495.600 ;
        RECT 545.400 495.400 549.000 495.800 ;
        RECT 546.000 494.400 546.800 494.800 ;
        RECT 550.000 494.400 550.600 495.800 ;
        RECT 551.600 495.400 552.400 499.800 ;
        RECT 555.800 498.400 557.000 499.800 ;
        RECT 555.800 497.800 557.200 498.400 ;
        RECT 560.400 497.800 561.200 499.800 ;
        RECT 564.800 498.400 565.600 499.800 ;
        RECT 564.800 497.800 566.800 498.400 ;
        RECT 556.400 497.000 557.200 497.800 ;
        RECT 560.600 497.200 561.200 497.800 ;
        RECT 560.600 496.600 563.400 497.200 ;
        RECT 562.600 496.400 563.400 496.600 ;
        RECT 564.400 496.400 565.200 497.200 ;
        RECT 566.000 497.000 566.800 497.800 ;
        RECT 554.600 495.400 555.400 495.600 ;
        RECT 551.600 494.800 555.400 495.400 ;
        RECT 535.600 494.200 537.200 494.400 ;
        RECT 526.200 493.600 537.200 494.200 ;
        RECT 538.800 493.800 540.400 494.400 ;
        RECT 538.800 493.600 539.600 493.800 ;
        RECT 541.800 493.600 544.400 494.400 ;
        RECT 545.200 493.800 546.800 494.400 ;
        RECT 545.200 493.600 546.000 493.800 ;
        RECT 548.200 493.600 550.800 494.400 ;
        RECT 524.400 492.800 525.200 493.000 ;
        RECT 521.400 492.200 525.200 492.800 ;
        RECT 521.400 492.000 522.200 492.200 ;
        RECT 523.000 491.400 523.800 491.600 ;
        RECT 519.600 490.800 523.800 491.400 ;
        RECT 513.200 489.600 514.600 490.200 ;
        RECT 515.200 489.600 516.200 490.200 ;
        RECT 497.200 483.000 498.000 487.000 ;
        RECT 501.400 482.200 502.200 489.200 ;
        RECT 509.400 482.200 510.200 489.600 ;
        RECT 511.000 488.400 511.600 489.600 ;
        RECT 510.800 487.600 511.600 488.400 ;
        RECT 514.000 488.400 514.600 489.600 ;
        RECT 514.000 487.600 514.800 488.400 ;
        RECT 515.400 482.200 516.200 489.600 ;
        RECT 519.600 482.200 520.400 490.800 ;
        RECT 522.800 489.600 523.600 490.800 ;
        RECT 526.200 490.400 526.800 493.600 ;
        RECT 533.400 493.400 534.200 493.600 ;
        RECT 535.000 492.400 535.800 492.600 ;
        RECT 529.200 492.300 530.000 492.400 ;
        RECT 530.800 492.300 535.800 492.400 ;
        RECT 529.200 491.800 535.800 492.300 ;
        RECT 529.200 491.700 531.600 491.800 ;
        RECT 529.200 491.600 530.000 491.700 ;
        RECT 530.800 491.600 531.600 491.700 ;
        RECT 540.400 491.600 541.200 493.200 ;
        RECT 532.400 491.000 538.000 491.200 ;
        RECT 532.200 490.800 538.000 491.000 ;
        RECT 524.400 489.800 526.800 490.400 ;
        RECT 528.200 490.600 538.000 490.800 ;
        RECT 528.200 490.200 533.000 490.600 ;
        RECT 524.400 488.800 525.000 489.800 ;
        RECT 523.600 488.000 525.000 488.800 ;
        RECT 526.600 489.000 527.400 489.200 ;
        RECT 528.200 489.000 528.800 490.200 ;
        RECT 526.600 488.400 528.800 489.000 ;
        RECT 529.400 489.000 534.800 489.600 ;
        RECT 529.400 488.800 530.200 489.000 ;
        RECT 534.000 488.800 534.800 489.000 ;
        RECT 527.800 487.400 528.600 487.600 ;
        RECT 530.600 487.400 531.400 487.600 ;
        RECT 524.400 486.200 525.200 487.000 ;
        RECT 527.800 486.800 531.400 487.400 ;
        RECT 528.600 486.200 529.200 486.800 ;
        RECT 534.000 486.200 534.800 487.000 ;
        RECT 523.800 482.200 525.000 486.200 ;
        RECT 528.400 482.200 529.200 486.200 ;
        RECT 532.800 485.600 534.800 486.200 ;
        RECT 532.800 482.200 533.600 485.600 ;
        RECT 537.200 482.200 538.000 490.600 ;
        RECT 541.800 490.200 542.400 493.600 ;
        RECT 546.800 491.600 547.600 493.200 ;
        RECT 548.200 490.400 548.800 493.600 ;
        RECT 551.600 491.400 552.400 494.800 ;
        RECT 558.600 494.200 559.400 494.400 ;
        RECT 564.400 494.200 565.000 496.400 ;
        RECT 569.200 495.000 570.000 499.800 ;
        RECT 570.800 495.800 571.600 499.800 ;
        RECT 572.400 496.000 573.200 499.800 ;
        RECT 575.600 496.000 576.400 499.800 ;
        RECT 578.800 496.000 579.600 499.800 ;
        RECT 572.400 495.800 576.400 496.000 ;
        RECT 571.000 494.400 571.600 495.800 ;
        RECT 572.600 495.400 576.200 495.800 ;
        RECT 578.600 495.200 579.600 496.000 ;
        RECT 574.800 494.400 575.600 494.800 ;
        RECT 567.600 494.200 569.200 494.400 ;
        RECT 558.200 493.600 569.200 494.200 ;
        RECT 570.800 493.600 573.400 494.400 ;
        RECT 574.800 493.800 576.400 494.400 ;
        RECT 575.600 493.600 576.400 493.800 ;
        RECT 556.400 492.800 557.200 493.000 ;
        RECT 553.400 492.200 557.200 492.800 ;
        RECT 553.400 492.000 554.200 492.200 ;
        RECT 555.000 491.400 555.800 491.600 ;
        RECT 551.600 490.800 555.800 491.400 ;
        RECT 543.600 490.200 544.400 490.400 ;
        RECT 541.400 489.600 542.400 490.200 ;
        RECT 543.000 489.600 544.400 490.200 ;
        RECT 546.800 489.600 548.800 490.400 ;
        RECT 550.000 490.300 550.800 490.400 ;
        RECT 551.600 490.300 552.400 490.800 ;
        RECT 558.200 490.400 558.800 493.600 ;
        RECT 565.400 493.400 566.200 493.600 ;
        RECT 567.000 492.400 567.800 492.600 ;
        RECT 572.800 492.400 573.400 493.600 ;
        RECT 562.800 491.800 567.800 492.400 ;
        RECT 562.800 491.600 563.600 491.800 ;
        RECT 572.400 491.600 573.400 492.400 ;
        RECT 574.000 491.600 574.800 493.200 ;
        RECT 564.400 491.000 570.000 491.200 ;
        RECT 564.200 490.800 570.000 491.000 ;
        RECT 550.000 490.200 552.400 490.300 ;
        RECT 549.400 489.700 552.400 490.200 ;
        RECT 549.400 489.600 550.800 489.700 ;
        RECT 541.400 482.200 542.200 489.600 ;
        RECT 543.000 488.400 543.600 489.600 ;
        RECT 542.800 487.600 543.600 488.400 ;
        RECT 547.800 482.200 548.600 489.600 ;
        RECT 549.400 488.400 550.000 489.600 ;
        RECT 549.200 487.600 550.000 488.400 ;
        RECT 551.600 482.200 552.400 489.700 ;
        RECT 556.400 489.800 558.800 490.400 ;
        RECT 560.200 490.600 570.000 490.800 ;
        RECT 560.200 490.200 565.000 490.600 ;
        RECT 556.400 488.800 557.000 489.800 ;
        RECT 555.600 488.000 557.000 488.800 ;
        RECT 558.600 489.000 559.400 489.200 ;
        RECT 560.200 489.000 560.800 490.200 ;
        RECT 558.600 488.400 560.800 489.000 ;
        RECT 561.400 489.000 566.800 489.600 ;
        RECT 561.400 488.800 562.200 489.000 ;
        RECT 566.000 488.800 566.800 489.000 ;
        RECT 559.800 487.400 560.600 487.600 ;
        RECT 562.600 487.400 563.400 487.600 ;
        RECT 556.400 486.200 557.200 487.000 ;
        RECT 559.800 486.800 563.400 487.400 ;
        RECT 560.600 486.200 561.200 486.800 ;
        RECT 566.000 486.200 566.800 487.000 ;
        RECT 555.800 482.200 557.000 486.200 ;
        RECT 560.400 482.200 561.200 486.200 ;
        RECT 564.800 485.600 566.800 486.200 ;
        RECT 564.800 482.200 565.600 485.600 ;
        RECT 569.200 482.200 570.000 490.600 ;
        RECT 570.800 490.200 571.600 490.400 ;
        RECT 572.800 490.200 573.400 491.600 ;
        RECT 578.600 490.800 579.400 495.200 ;
        RECT 580.400 494.600 581.200 499.800 ;
        RECT 586.800 496.600 587.600 499.800 ;
        RECT 588.400 497.000 589.200 499.800 ;
        RECT 590.000 497.000 590.800 499.800 ;
        RECT 591.600 497.000 592.400 499.800 ;
        RECT 593.200 497.000 594.000 499.800 ;
        RECT 596.400 497.000 597.200 499.800 ;
        RECT 599.600 497.000 600.400 499.800 ;
        RECT 601.200 497.000 602.000 499.800 ;
        RECT 602.800 497.000 603.600 499.800 ;
        RECT 585.200 495.800 587.600 496.600 ;
        RECT 604.400 496.600 605.200 499.800 ;
        RECT 585.200 495.200 586.000 495.800 ;
        RECT 580.000 494.000 581.200 494.600 ;
        RECT 584.200 494.600 586.000 495.200 ;
        RECT 590.000 495.600 591.000 496.400 ;
        RECT 594.000 495.600 595.600 496.400 ;
        RECT 596.400 495.800 601.000 496.400 ;
        RECT 604.400 495.800 607.000 496.600 ;
        RECT 596.400 495.600 597.200 495.800 ;
        RECT 580.000 492.000 580.600 494.000 ;
        RECT 584.200 493.400 585.000 494.600 ;
        RECT 581.200 492.600 585.000 493.400 ;
        RECT 590.000 492.800 590.800 495.600 ;
        RECT 596.400 494.800 597.200 495.000 ;
        RECT 592.800 494.200 597.200 494.800 ;
        RECT 592.800 494.000 593.600 494.200 ;
        RECT 598.000 493.600 598.800 495.200 ;
        RECT 600.200 493.400 601.000 495.800 ;
        RECT 606.200 495.200 607.000 495.800 ;
        RECT 606.200 494.400 609.200 495.200 ;
        RECT 610.800 493.800 611.600 499.800 ;
        RECT 593.200 492.600 596.400 493.400 ;
        RECT 600.200 492.600 602.200 493.400 ;
        RECT 602.800 493.000 611.600 493.800 ;
        RECT 586.800 492.000 587.600 492.600 ;
        RECT 604.400 492.000 605.200 492.400 ;
        RECT 606.000 492.000 606.800 492.400 ;
        RECT 609.400 492.000 610.200 492.200 ;
        RECT 580.000 491.400 580.800 492.000 ;
        RECT 586.800 491.400 610.200 492.000 ;
        RECT 570.800 489.600 572.200 490.200 ;
        RECT 572.800 489.600 573.800 490.200 ;
        RECT 578.600 490.000 579.600 490.800 ;
        RECT 571.600 488.400 572.200 489.600 ;
        RECT 571.600 487.600 572.400 488.400 ;
        RECT 573.000 482.200 573.800 489.600 ;
        RECT 578.800 482.200 579.600 490.000 ;
        RECT 580.200 489.600 580.800 491.400 ;
        RECT 580.200 489.000 589.200 489.600 ;
        RECT 580.200 487.400 580.800 489.000 ;
        RECT 588.400 488.800 589.200 489.000 ;
        RECT 591.600 489.000 600.200 489.600 ;
        RECT 591.600 488.800 592.400 489.000 ;
        RECT 583.400 487.600 586.000 488.400 ;
        RECT 580.200 486.800 582.800 487.400 ;
        RECT 582.000 482.200 582.800 486.800 ;
        RECT 585.200 482.200 586.000 487.600 ;
        RECT 586.600 486.800 590.800 487.600 ;
        RECT 588.400 482.200 589.200 485.000 ;
        RECT 590.000 482.200 590.800 485.000 ;
        RECT 591.600 482.200 592.400 485.000 ;
        RECT 593.200 482.200 594.000 488.400 ;
        RECT 596.400 487.600 599.000 488.400 ;
        RECT 599.600 488.200 600.200 489.000 ;
        RECT 601.200 489.400 602.000 489.600 ;
        RECT 601.200 489.000 606.600 489.400 ;
        RECT 601.200 488.800 607.400 489.000 ;
        RECT 606.000 488.200 607.400 488.800 ;
        RECT 599.600 487.600 605.400 488.200 ;
        RECT 608.400 488.000 610.000 488.800 ;
        RECT 608.400 487.600 609.000 488.000 ;
        RECT 596.400 482.200 597.200 487.000 ;
        RECT 599.600 482.200 600.400 487.000 ;
        RECT 604.800 486.800 609.000 487.600 ;
        RECT 610.800 487.400 611.600 493.000 ;
        RECT 609.600 486.800 611.600 487.400 ;
        RECT 601.200 482.200 602.000 485.000 ;
        RECT 602.800 482.200 603.600 485.000 ;
        RECT 606.000 482.200 606.800 486.800 ;
        RECT 609.600 486.200 610.200 486.800 ;
        RECT 609.200 485.600 610.200 486.200 ;
        RECT 609.200 482.200 610.000 485.600 ;
        RECT 1.200 471.400 2.000 479.800 ;
        RECT 5.600 476.400 6.400 479.800 ;
        RECT 4.400 475.800 6.400 476.400 ;
        RECT 10.000 475.800 10.800 479.800 ;
        RECT 14.200 475.800 15.400 479.800 ;
        RECT 4.400 475.000 5.200 475.800 ;
        RECT 10.000 475.200 10.600 475.800 ;
        RECT 7.800 474.600 11.400 475.200 ;
        RECT 14.000 475.000 14.800 475.800 ;
        RECT 7.800 474.400 8.600 474.600 ;
        RECT 10.600 474.400 11.400 474.600 ;
        RECT 4.400 473.000 5.200 473.200 ;
        RECT 9.000 473.000 9.800 473.200 ;
        RECT 4.400 472.400 9.800 473.000 ;
        RECT 10.400 473.000 12.600 473.600 ;
        RECT 10.400 471.800 11.000 473.000 ;
        RECT 11.800 472.800 12.600 473.000 ;
        RECT 14.200 473.200 15.600 474.000 ;
        RECT 14.200 472.200 14.800 473.200 ;
        RECT 6.200 471.400 11.000 471.800 ;
        RECT 1.200 471.200 11.000 471.400 ;
        RECT 12.400 471.600 14.800 472.200 ;
        RECT 1.200 471.000 7.000 471.200 ;
        RECT 1.200 470.800 6.800 471.000 ;
        RECT 12.400 470.400 13.000 471.600 ;
        RECT 18.800 471.200 19.600 479.800 ;
        RECT 23.000 472.400 23.800 479.800 ;
        RECT 24.400 473.600 25.200 474.400 ;
        RECT 24.600 472.400 25.200 473.600 ;
        RECT 27.600 473.600 28.400 474.400 ;
        RECT 27.600 472.400 28.200 473.600 ;
        RECT 29.000 472.400 29.800 479.800 ;
        RECT 23.000 471.800 24.000 472.400 ;
        RECT 24.600 471.800 26.000 472.400 ;
        RECT 15.400 470.600 19.600 471.200 ;
        RECT 15.400 470.400 16.200 470.600 ;
        RECT 7.600 470.200 8.400 470.400 ;
        RECT 3.400 469.600 8.400 470.200 ;
        RECT 12.400 469.600 13.200 470.400 ;
        RECT 17.000 469.800 17.800 470.000 ;
        RECT 3.400 469.400 4.200 469.600 ;
        RECT 5.000 468.400 5.800 468.600 ;
        RECT 12.400 468.400 13.000 469.600 ;
        RECT 14.000 469.200 17.800 469.800 ;
        RECT 14.000 469.000 14.800 469.200 ;
        RECT 2.000 467.800 13.000 468.400 ;
        RECT 2.000 467.600 3.600 467.800 ;
        RECT 1.200 462.200 2.000 467.000 ;
        RECT 6.200 465.600 6.800 467.800 ;
        RECT 11.800 467.600 12.600 467.800 ;
        RECT 18.800 467.200 19.600 470.600 ;
        RECT 23.400 470.400 24.000 471.800 ;
        RECT 25.200 471.600 26.000 471.800 ;
        RECT 26.800 471.800 28.200 472.400 ;
        RECT 28.800 471.800 29.800 472.400 ;
        RECT 26.800 471.600 27.600 471.800 ;
        RECT 22.000 468.800 22.800 470.400 ;
        RECT 23.400 469.600 24.400 470.400 ;
        RECT 25.300 470.300 25.900 471.600 ;
        RECT 28.800 470.300 29.400 471.800 ;
        RECT 33.200 471.400 34.000 479.800 ;
        RECT 37.600 476.400 38.400 479.800 ;
        RECT 36.400 475.800 38.400 476.400 ;
        RECT 42.000 475.800 42.800 479.800 ;
        RECT 46.200 475.800 47.400 479.800 ;
        RECT 36.400 475.000 37.200 475.800 ;
        RECT 42.000 475.200 42.600 475.800 ;
        RECT 39.800 474.600 43.400 475.200 ;
        RECT 46.000 475.000 46.800 475.800 ;
        RECT 39.800 474.400 40.600 474.600 ;
        RECT 42.600 474.400 43.400 474.600 ;
        RECT 36.400 473.000 37.200 473.200 ;
        RECT 41.000 473.000 41.800 473.200 ;
        RECT 36.400 472.400 41.800 473.000 ;
        RECT 42.400 473.000 44.600 473.600 ;
        RECT 42.400 471.800 43.000 473.000 ;
        RECT 43.800 472.800 44.600 473.000 ;
        RECT 46.200 473.200 47.600 474.000 ;
        RECT 46.200 472.200 46.800 473.200 ;
        RECT 38.200 471.400 43.000 471.800 ;
        RECT 33.200 471.200 43.000 471.400 ;
        RECT 44.400 471.600 46.800 472.200 ;
        RECT 33.200 471.000 39.000 471.200 ;
        RECT 33.200 470.800 38.800 471.000 ;
        RECT 25.300 469.700 29.400 470.300 ;
        RECT 23.400 468.400 24.000 469.600 ;
        RECT 28.800 468.400 29.400 469.700 ;
        RECT 30.000 468.800 30.800 470.400 ;
        RECT 39.600 470.200 40.400 470.400 ;
        RECT 35.400 469.600 40.400 470.200 ;
        RECT 35.400 469.400 36.200 469.600 ;
        RECT 37.000 468.400 37.800 468.600 ;
        RECT 44.400 468.400 45.000 471.600 ;
        RECT 50.800 471.200 51.600 479.800 ;
        RECT 55.000 472.400 55.800 479.800 ;
        RECT 56.400 473.600 57.200 474.400 ;
        RECT 56.600 472.400 57.200 473.600 ;
        RECT 59.600 473.600 60.400 474.400 ;
        RECT 59.600 472.400 60.200 473.600 ;
        RECT 61.000 472.400 61.800 479.800 ;
        RECT 69.000 472.800 69.800 479.800 ;
        RECT 73.200 475.000 74.000 479.000 ;
        RECT 55.000 471.800 56.000 472.400 ;
        RECT 56.600 471.800 58.000 472.400 ;
        RECT 47.400 470.600 51.600 471.200 ;
        RECT 47.400 470.400 48.200 470.600 ;
        RECT 49.000 469.800 49.800 470.000 ;
        RECT 46.000 469.200 49.800 469.800 ;
        RECT 46.000 469.000 46.800 469.200 ;
        RECT 20.400 468.200 21.200 468.400 ;
        RECT 20.400 467.600 22.000 468.200 ;
        RECT 23.400 467.600 26.000 468.400 ;
        RECT 26.800 467.600 29.400 468.400 ;
        RECT 31.600 468.200 32.400 468.400 ;
        RECT 30.800 467.600 32.400 468.200 ;
        RECT 34.000 467.800 45.000 468.400 ;
        RECT 34.000 467.600 35.600 467.800 ;
        RECT 38.000 467.600 38.800 467.800 ;
        RECT 43.800 467.600 44.600 467.800 ;
        RECT 21.200 467.200 22.000 467.600 ;
        RECT 15.800 466.600 19.600 467.200 ;
        RECT 15.800 466.400 16.600 466.600 ;
        RECT 4.400 464.200 5.200 465.000 ;
        RECT 6.000 464.800 6.800 465.600 ;
        RECT 7.800 465.400 8.600 465.600 ;
        RECT 7.800 464.800 10.600 465.400 ;
        RECT 10.000 464.200 10.600 464.800 ;
        RECT 14.000 464.200 14.800 465.000 ;
        RECT 4.400 463.600 6.400 464.200 ;
        RECT 5.600 462.200 6.400 463.600 ;
        RECT 10.000 462.200 10.800 464.200 ;
        RECT 14.000 463.600 15.400 464.200 ;
        RECT 14.200 462.200 15.400 463.600 ;
        RECT 18.800 462.200 19.600 466.600 ;
        RECT 20.600 466.200 24.200 466.600 ;
        RECT 25.200 466.200 25.800 467.600 ;
        RECT 27.000 466.200 27.600 467.600 ;
        RECT 30.800 467.200 31.600 467.600 ;
        RECT 28.600 466.200 32.200 466.600 ;
        RECT 20.400 466.000 24.400 466.200 ;
        RECT 20.400 462.200 21.200 466.000 ;
        RECT 23.600 462.200 24.400 466.000 ;
        RECT 25.200 462.200 26.000 466.200 ;
        RECT 26.800 462.200 27.600 466.200 ;
        RECT 28.400 466.000 32.400 466.200 ;
        RECT 28.400 462.200 29.200 466.000 ;
        RECT 31.600 462.200 32.400 466.000 ;
        RECT 33.200 462.200 34.000 467.000 ;
        RECT 38.200 465.600 38.800 467.600 ;
        RECT 50.800 467.200 51.600 470.600 ;
        RECT 54.000 468.800 54.800 470.400 ;
        RECT 55.400 470.300 56.000 471.800 ;
        RECT 57.200 471.600 58.000 471.800 ;
        RECT 58.800 471.800 60.200 472.400 ;
        RECT 60.800 471.800 61.800 472.400 ;
        RECT 68.200 472.200 69.800 472.800 ;
        RECT 58.800 471.600 59.600 471.800 ;
        RECT 58.900 470.300 59.500 471.600 ;
        RECT 55.400 469.700 59.500 470.300 ;
        RECT 55.400 468.400 56.000 469.700 ;
        RECT 60.800 468.400 61.400 471.800 ;
        RECT 62.000 468.800 62.800 470.400 ;
        RECT 65.200 470.300 66.000 470.400 ;
        RECT 66.800 470.300 67.600 471.200 ;
        RECT 65.200 469.700 67.600 470.300 ;
        RECT 65.200 469.600 66.000 469.700 ;
        RECT 66.800 469.600 67.600 469.700 ;
        RECT 68.200 468.400 68.800 472.200 ;
        RECT 73.400 471.600 74.000 475.000 ;
        RECT 74.800 471.600 75.600 474.400 ;
        RECT 70.200 471.000 74.000 471.600 ;
        RECT 70.200 469.000 70.800 471.000 ;
        RECT 52.400 468.200 53.200 468.400 ;
        RECT 52.400 467.600 54.000 468.200 ;
        RECT 55.400 467.600 58.000 468.400 ;
        RECT 58.800 467.600 61.400 468.400 ;
        RECT 63.600 468.200 64.400 468.400 ;
        RECT 62.800 467.600 64.400 468.200 ;
        RECT 66.800 467.600 68.800 468.400 ;
        RECT 69.400 468.200 70.800 469.000 ;
        RECT 71.600 468.800 72.400 470.400 ;
        RECT 73.200 468.800 74.000 470.400 ;
        RECT 53.200 467.200 54.000 467.600 ;
        RECT 47.800 466.600 51.600 467.200 ;
        RECT 47.800 466.400 48.600 466.600 ;
        RECT 36.400 464.200 37.200 465.000 ;
        RECT 38.000 464.800 38.800 465.600 ;
        RECT 39.800 465.400 40.600 465.600 ;
        RECT 39.800 464.800 42.600 465.400 ;
        RECT 42.000 464.200 42.600 464.800 ;
        RECT 46.000 464.200 46.800 465.000 ;
        RECT 36.400 463.600 38.400 464.200 ;
        RECT 37.600 462.200 38.400 463.600 ;
        RECT 42.000 462.200 42.800 464.200 ;
        RECT 46.000 463.600 47.400 464.200 ;
        RECT 46.200 462.200 47.400 463.600 ;
        RECT 50.800 462.200 51.600 466.600 ;
        RECT 52.600 466.200 56.200 466.600 ;
        RECT 57.200 466.200 57.800 467.600 ;
        RECT 59.000 466.200 59.600 467.600 ;
        RECT 62.800 467.200 63.600 467.600 ;
        RECT 68.200 467.000 68.800 467.600 ;
        RECT 69.800 467.800 70.800 468.200 ;
        RECT 69.800 467.200 74.000 467.800 ;
        RECT 68.200 466.600 69.000 467.000 ;
        RECT 60.600 466.200 64.200 466.600 ;
        RECT 52.400 466.000 56.400 466.200 ;
        RECT 52.400 462.200 53.200 466.000 ;
        RECT 55.600 462.200 56.400 466.000 ;
        RECT 57.200 462.200 58.000 466.200 ;
        RECT 58.800 462.200 59.600 466.200 ;
        RECT 60.400 466.000 64.400 466.200 ;
        RECT 68.200 466.000 69.800 466.600 ;
        RECT 60.400 462.200 61.200 466.000 ;
        RECT 63.600 462.200 64.400 466.000 ;
        RECT 69.000 464.400 69.800 466.000 ;
        RECT 73.400 465.000 74.000 467.200 ;
        RECT 76.400 466.200 77.200 479.800 ;
        RECT 83.400 472.800 84.200 479.800 ;
        RECT 87.600 475.000 88.400 479.000 ;
        RECT 82.600 472.200 84.200 472.800 ;
        RECT 81.200 469.600 82.000 471.200 ;
        RECT 82.600 468.400 83.200 472.200 ;
        RECT 87.800 471.600 88.400 475.000 ;
        RECT 90.800 472.800 91.600 479.800 ;
        RECT 84.600 471.000 88.400 471.600 ;
        RECT 90.600 471.800 91.600 472.800 ;
        RECT 94.000 472.400 94.800 479.800 ;
        RECT 99.400 478.400 100.200 479.800 ;
        RECT 98.800 477.600 100.200 478.400 ;
        RECT 99.400 472.800 100.200 477.600 ;
        RECT 103.600 475.000 104.400 479.000 ;
        RECT 92.200 471.800 94.800 472.400 ;
        RECT 98.600 472.200 100.200 472.800 ;
        RECT 84.600 469.000 85.200 471.000 ;
        RECT 78.000 466.800 78.800 468.400 ;
        RECT 79.600 468.300 80.400 468.400 ;
        RECT 81.200 468.300 83.200 468.400 ;
        RECT 79.600 467.700 83.200 468.300 ;
        RECT 83.800 468.200 85.200 469.000 ;
        RECT 86.000 468.800 86.800 470.400 ;
        RECT 87.600 468.800 88.400 470.400 ;
        RECT 79.600 467.600 80.400 467.700 ;
        RECT 81.200 467.600 83.200 467.700 ;
        RECT 82.600 467.000 83.200 467.600 ;
        RECT 84.200 467.800 85.200 468.200 ;
        RECT 90.600 468.400 91.200 471.800 ;
        RECT 92.200 469.800 92.800 471.800 ;
        RECT 91.800 469.000 92.800 469.800 ;
        RECT 84.200 467.200 88.400 467.800 ;
        RECT 68.400 463.600 69.800 464.400 ;
        RECT 69.000 463.000 69.800 463.600 ;
        RECT 73.200 463.000 74.000 465.000 ;
        RECT 75.400 465.600 77.200 466.200 ;
        RECT 82.600 466.600 83.400 467.000 ;
        RECT 82.600 466.000 84.200 466.600 ;
        RECT 75.400 464.400 76.200 465.600 ;
        RECT 74.800 463.600 76.200 464.400 ;
        RECT 75.400 462.200 76.200 463.600 ;
        RECT 83.400 463.000 84.200 466.000 ;
        RECT 87.800 465.000 88.400 467.200 ;
        RECT 90.600 467.600 91.600 468.400 ;
        RECT 90.600 466.200 91.200 467.600 ;
        RECT 92.200 467.400 92.800 469.000 ;
        RECT 93.800 469.600 94.800 470.400 ;
        RECT 95.600 470.300 96.400 470.400 ;
        RECT 97.200 470.300 98.000 471.200 ;
        RECT 95.600 469.700 98.000 470.300 ;
        RECT 95.600 469.600 96.400 469.700 ;
        RECT 97.200 469.600 98.000 469.700 ;
        RECT 93.800 468.800 94.600 469.600 ;
        RECT 98.600 468.400 99.200 472.200 ;
        RECT 103.800 471.600 104.400 475.000 ;
        RECT 106.800 472.800 107.600 479.800 ;
        RECT 100.600 471.000 104.400 471.600 ;
        RECT 106.600 471.800 107.600 472.800 ;
        RECT 110.000 472.400 110.800 479.800 ;
        RECT 108.200 471.800 110.800 472.400 ;
        RECT 100.600 469.000 101.200 471.000 ;
        RECT 97.200 467.600 99.200 468.400 ;
        RECT 99.800 468.200 101.200 469.000 ;
        RECT 102.000 468.800 102.800 470.400 ;
        RECT 103.600 468.800 104.400 470.400 ;
        RECT 92.200 466.800 94.800 467.400 ;
        RECT 90.600 465.600 91.600 466.200 ;
        RECT 87.600 463.000 88.400 465.000 ;
        RECT 90.800 462.200 91.600 465.600 ;
        RECT 94.000 462.200 94.800 466.800 ;
        RECT 98.600 467.000 99.200 467.600 ;
        RECT 100.200 467.800 101.200 468.200 ;
        RECT 106.600 468.400 107.200 471.800 ;
        RECT 108.200 469.800 108.800 471.800 ;
        RECT 107.800 469.000 108.800 469.800 ;
        RECT 100.200 467.200 104.400 467.800 ;
        RECT 98.600 466.600 99.400 467.000 ;
        RECT 98.600 466.000 100.200 466.600 ;
        RECT 99.400 463.000 100.200 466.000 ;
        RECT 103.800 465.000 104.400 467.200 ;
        RECT 106.600 467.600 107.600 468.400 ;
        RECT 106.600 466.200 107.200 467.600 ;
        RECT 108.200 467.400 108.800 469.000 ;
        RECT 109.800 470.300 110.800 470.400 ;
        RECT 111.600 470.300 112.400 470.400 ;
        RECT 109.800 469.700 112.400 470.300 ;
        RECT 109.800 469.600 110.800 469.700 ;
        RECT 111.600 469.600 112.400 469.700 ;
        RECT 109.800 468.800 110.600 469.600 ;
        RECT 108.200 466.800 110.800 467.400 ;
        RECT 106.600 465.600 107.600 466.200 ;
        RECT 103.600 463.000 104.400 465.000 ;
        RECT 106.800 462.200 107.600 465.600 ;
        RECT 110.000 462.200 110.800 466.800 ;
        RECT 111.600 464.800 112.400 466.400 ;
        RECT 113.200 462.200 114.000 479.800 ;
        RECT 116.400 475.800 117.200 479.800 ;
        RECT 116.600 475.600 117.200 475.800 ;
        RECT 119.600 475.800 120.400 479.800 ;
        RECT 123.400 476.400 124.200 479.800 ;
        RECT 119.600 475.600 120.200 475.800 ;
        RECT 116.600 475.000 120.200 475.600 ;
        RECT 119.600 474.400 120.200 475.000 ;
        RECT 123.400 475.600 125.200 476.400 ;
        RECT 118.000 472.800 118.800 474.400 ;
        RECT 119.600 473.600 120.400 474.400 ;
        RECT 122.000 473.600 122.800 474.400 ;
        RECT 119.600 472.400 120.200 473.600 ;
        RECT 122.000 472.400 122.600 473.600 ;
        RECT 123.400 472.400 124.200 475.600 ;
        RECT 128.400 473.600 129.200 474.400 ;
        RECT 128.400 472.400 129.000 473.600 ;
        RECT 129.800 472.400 130.600 479.800 ;
        RECT 136.600 474.400 137.400 479.800 ;
        RECT 135.600 473.600 137.400 474.400 ;
        RECT 138.000 473.600 138.800 474.400 ;
        RECT 136.600 472.400 137.400 473.600 ;
        RECT 138.200 472.400 138.800 473.600 ;
        RECT 143.000 472.600 143.800 479.800 ;
        RECT 114.800 470.800 115.600 472.400 ;
        RECT 119.600 471.600 120.400 472.400 ;
        RECT 121.200 471.800 122.600 472.400 ;
        RECT 123.200 471.800 124.200 472.400 ;
        RECT 127.600 471.800 129.000 472.400 ;
        RECT 121.200 471.600 122.000 471.800 ;
        RECT 116.400 469.600 118.000 470.400 ;
        RECT 119.600 468.400 120.200 471.600 ;
        RECT 123.200 468.400 123.800 471.800 ;
        RECT 127.600 471.600 128.400 471.800 ;
        RECT 129.600 471.600 131.600 472.400 ;
        RECT 136.600 471.800 137.600 472.400 ;
        RECT 138.200 471.800 139.600 472.400 ;
        RECT 142.000 471.800 143.800 472.600 ;
        RECT 147.800 472.400 148.600 479.800 ;
        RECT 149.200 473.600 150.000 474.400 ;
        RECT 149.400 472.400 150.000 473.600 ;
        RECT 156.400 472.400 157.200 479.800 ;
        RECT 159.600 472.800 160.400 479.800 ;
        RECT 166.600 472.800 167.400 479.800 ;
        RECT 170.800 475.000 171.600 479.000 ;
        RECT 147.800 471.800 148.800 472.400 ;
        RECT 149.400 471.800 150.800 472.400 ;
        RECT 156.400 471.800 159.000 472.400 ;
        RECT 159.600 471.800 160.600 472.800 ;
        RECT 124.400 470.300 125.200 470.400 ;
        RECT 127.600 470.300 128.400 470.400 ;
        RECT 124.400 469.700 128.400 470.300 ;
        RECT 124.400 468.800 125.200 469.700 ;
        RECT 127.600 469.600 128.400 469.700 ;
        RECT 129.600 468.400 130.200 471.600 ;
        RECT 130.800 468.800 131.600 470.400 ;
        RECT 135.600 468.800 136.400 470.400 ;
        RECT 137.000 468.400 137.600 471.800 ;
        RECT 138.800 471.600 139.600 471.800 ;
        RECT 142.200 468.400 142.800 471.800 ;
        RECT 143.600 469.600 144.400 471.200 ;
        RECT 146.800 468.800 147.600 470.400 ;
        RECT 148.200 468.400 148.800 471.800 ;
        RECT 150.000 471.600 150.800 471.800 ;
        RECT 154.800 470.300 155.600 470.400 ;
        RECT 156.400 470.300 157.400 470.400 ;
        RECT 154.800 469.700 157.400 470.300 ;
        RECT 154.800 469.600 155.600 469.700 ;
        RECT 156.400 469.600 157.400 469.700 ;
        RECT 156.600 468.800 157.400 469.600 ;
        RECT 158.400 469.800 159.000 471.800 ;
        RECT 158.400 469.000 159.400 469.800 ;
        RECT 118.600 468.200 120.200 468.400 ;
        RECT 118.400 467.800 120.200 468.200 ;
        RECT 118.400 462.200 119.200 467.800 ;
        RECT 121.200 467.600 123.800 468.400 ;
        RECT 126.000 468.200 126.800 468.400 ;
        RECT 125.200 467.600 126.800 468.200 ;
        RECT 127.600 467.600 130.200 468.400 ;
        RECT 132.400 468.200 133.200 468.400 ;
        RECT 131.600 467.600 133.200 468.200 ;
        RECT 134.000 468.200 134.800 468.400 ;
        RECT 134.000 467.600 135.600 468.200 ;
        RECT 137.000 467.600 139.600 468.400 ;
        RECT 142.000 467.600 142.800 468.400 ;
        RECT 145.200 468.200 146.000 468.400 ;
        RECT 145.200 467.600 146.800 468.200 ;
        RECT 148.200 467.600 150.800 468.400 ;
        RECT 121.400 466.200 122.000 467.600 ;
        RECT 125.200 467.200 126.000 467.600 ;
        RECT 123.000 466.200 126.600 466.600 ;
        RECT 127.800 466.200 128.400 467.600 ;
        RECT 131.600 467.200 132.400 467.600 ;
        RECT 134.800 467.200 135.600 467.600 ;
        RECT 129.400 466.200 133.000 466.600 ;
        RECT 134.200 466.200 137.800 466.600 ;
        RECT 138.800 466.200 139.400 467.600 ;
        RECT 121.200 462.200 122.000 466.200 ;
        RECT 122.800 466.000 126.800 466.200 ;
        RECT 122.800 462.200 123.600 466.000 ;
        RECT 126.000 462.200 126.800 466.000 ;
        RECT 127.600 462.200 128.400 466.200 ;
        RECT 129.200 466.000 133.200 466.200 ;
        RECT 129.200 462.200 130.000 466.000 ;
        RECT 132.400 462.200 133.200 466.000 ;
        RECT 134.000 466.000 138.000 466.200 ;
        RECT 134.000 462.200 134.800 466.000 ;
        RECT 137.200 462.200 138.000 466.000 ;
        RECT 138.800 462.200 139.600 466.200 ;
        RECT 140.400 464.800 141.200 466.400 ;
        RECT 142.200 464.400 142.800 467.600 ;
        RECT 146.000 467.200 146.800 467.600 ;
        RECT 145.400 466.200 149.000 466.600 ;
        RECT 150.000 466.300 150.600 467.600 ;
        RECT 158.400 467.400 159.000 469.000 ;
        RECT 160.000 468.400 160.600 471.800 ;
        RECT 165.800 472.200 167.400 472.800 ;
        RECT 164.400 469.600 165.200 471.200 ;
        RECT 165.800 470.400 166.400 472.200 ;
        RECT 171.000 471.600 171.600 475.000 ;
        RECT 175.000 472.400 175.800 479.800 ;
        RECT 176.400 473.600 177.200 474.400 ;
        RECT 176.600 472.400 177.200 473.600 ;
        RECT 181.400 472.400 182.200 479.800 ;
        RECT 182.800 473.600 183.600 474.400 ;
        RECT 183.000 472.400 183.600 473.600 ;
        RECT 175.000 471.800 176.000 472.400 ;
        RECT 176.600 471.800 178.000 472.400 ;
        RECT 181.400 471.800 182.400 472.400 ;
        RECT 183.000 471.800 184.400 472.400 ;
        RECT 167.800 471.000 171.600 471.600 ;
        RECT 165.800 469.600 166.800 470.400 ;
        RECT 165.800 468.400 166.400 469.600 ;
        RECT 167.800 469.000 168.400 471.000 ;
        RECT 159.600 468.300 160.600 468.400 ;
        RECT 162.800 468.300 163.600 468.400 ;
        RECT 159.600 467.700 163.600 468.300 ;
        RECT 159.600 467.600 160.600 467.700 ;
        RECT 162.800 467.600 163.600 467.700 ;
        RECT 164.400 467.600 166.400 468.400 ;
        RECT 167.000 468.200 168.400 469.000 ;
        RECT 169.200 468.800 170.000 470.400 ;
        RECT 170.800 468.800 171.600 470.400 ;
        RECT 172.400 470.300 173.200 470.400 ;
        RECT 174.000 470.300 174.800 470.400 ;
        RECT 172.400 469.700 174.800 470.300 ;
        RECT 172.400 469.600 173.200 469.700 ;
        RECT 174.000 468.800 174.800 469.700 ;
        RECT 175.400 468.400 176.000 471.800 ;
        RECT 177.200 471.600 178.000 471.800 ;
        RECT 181.800 470.400 182.400 471.800 ;
        RECT 183.600 471.600 184.400 471.800 ;
        RECT 185.200 471.200 186.000 479.800 ;
        RECT 189.400 475.800 190.600 479.800 ;
        RECT 194.000 475.800 194.800 479.800 ;
        RECT 198.400 476.400 199.200 479.800 ;
        RECT 198.400 475.800 200.400 476.400 ;
        RECT 190.000 475.000 190.800 475.800 ;
        RECT 194.200 475.200 194.800 475.800 ;
        RECT 193.400 474.600 197.000 475.200 ;
        RECT 199.600 475.000 200.400 475.800 ;
        RECT 193.400 474.400 194.200 474.600 ;
        RECT 196.200 474.400 197.000 474.600 ;
        RECT 189.200 473.200 190.600 474.000 ;
        RECT 190.000 472.200 190.600 473.200 ;
        RECT 192.200 473.000 194.400 473.600 ;
        RECT 192.200 472.800 193.000 473.000 ;
        RECT 190.000 471.600 192.400 472.200 ;
        RECT 185.200 470.600 189.400 471.200 ;
        RECT 180.400 468.800 181.200 470.400 ;
        RECT 181.800 469.600 182.800 470.400 ;
        RECT 181.800 468.400 182.400 469.600 ;
        RECT 156.400 466.800 159.000 467.400 ;
        RECT 153.200 466.300 154.000 466.400 ;
        RECT 142.000 462.200 142.800 464.400 ;
        RECT 145.200 466.000 149.200 466.200 ;
        RECT 145.200 462.200 146.000 466.000 ;
        RECT 148.400 462.200 149.200 466.000 ;
        RECT 150.000 465.700 154.000 466.300 ;
        RECT 150.000 462.200 150.800 465.700 ;
        RECT 153.200 465.600 154.000 465.700 ;
        RECT 156.400 462.200 157.200 466.800 ;
        RECT 160.000 466.200 160.600 467.600 ;
        RECT 159.600 465.600 160.600 466.200 ;
        RECT 165.800 467.000 166.400 467.600 ;
        RECT 167.400 467.800 168.400 468.200 ;
        RECT 172.400 468.200 173.200 468.400 ;
        RECT 167.400 467.200 171.600 467.800 ;
        RECT 172.400 467.600 174.000 468.200 ;
        RECT 175.400 467.600 178.000 468.400 ;
        RECT 178.800 468.200 179.600 468.400 ;
        RECT 178.800 467.600 180.400 468.200 ;
        RECT 181.800 467.600 184.400 468.400 ;
        RECT 173.200 467.200 174.000 467.600 ;
        RECT 165.800 466.600 166.600 467.000 ;
        RECT 165.800 466.000 167.400 466.600 ;
        RECT 159.600 462.200 160.400 465.600 ;
        RECT 166.600 463.000 167.400 466.000 ;
        RECT 171.000 465.000 171.600 467.200 ;
        RECT 172.600 466.200 176.200 466.600 ;
        RECT 177.200 466.200 177.800 467.600 ;
        RECT 179.600 467.200 180.400 467.600 ;
        RECT 179.000 466.200 182.600 466.600 ;
        RECT 183.600 466.200 184.200 467.600 ;
        RECT 185.200 467.200 186.000 470.600 ;
        RECT 188.600 470.400 189.400 470.600 ;
        RECT 187.000 469.800 187.800 470.000 ;
        RECT 187.000 469.200 190.800 469.800 ;
        RECT 190.000 469.000 190.800 469.200 ;
        RECT 191.800 468.400 192.400 471.600 ;
        RECT 193.800 471.800 194.400 473.000 ;
        RECT 195.000 473.000 195.800 473.200 ;
        RECT 199.600 473.000 200.400 473.200 ;
        RECT 195.000 472.400 200.400 473.000 ;
        RECT 193.800 471.400 198.600 471.800 ;
        RECT 202.800 471.400 203.600 479.800 ;
        RECT 193.800 471.200 203.600 471.400 ;
        RECT 197.800 471.000 203.600 471.200 ;
        RECT 198.000 470.800 203.600 471.000 ;
        RECT 196.400 470.200 197.200 470.400 ;
        RECT 196.400 469.600 201.400 470.200 ;
        RECT 200.600 469.400 201.400 469.600 ;
        RECT 199.000 468.400 199.800 468.600 ;
        RECT 191.800 467.800 202.800 468.400 ;
        RECT 192.200 467.600 193.000 467.800 ;
        RECT 185.200 466.600 189.000 467.200 ;
        RECT 170.800 463.000 171.600 465.000 ;
        RECT 172.400 466.000 176.400 466.200 ;
        RECT 172.400 462.200 173.200 466.000 ;
        RECT 175.600 462.200 176.400 466.000 ;
        RECT 177.200 462.200 178.000 466.200 ;
        RECT 178.800 466.000 182.800 466.200 ;
        RECT 178.800 462.200 179.600 466.000 ;
        RECT 182.000 462.200 182.800 466.000 ;
        RECT 183.600 462.200 184.400 466.200 ;
        RECT 185.200 462.200 186.000 466.600 ;
        RECT 188.200 466.400 189.000 466.600 ;
        RECT 198.000 465.600 198.600 467.800 ;
        RECT 201.200 467.600 202.800 467.800 ;
        RECT 196.200 465.400 197.000 465.600 ;
        RECT 190.000 464.200 190.800 465.000 ;
        RECT 194.200 464.800 197.000 465.400 ;
        RECT 198.000 464.800 198.800 465.600 ;
        RECT 194.200 464.200 194.800 464.800 ;
        RECT 199.600 464.200 200.400 465.000 ;
        RECT 189.400 463.600 190.800 464.200 ;
        RECT 189.400 462.200 190.600 463.600 ;
        RECT 194.000 462.200 194.800 464.200 ;
        RECT 198.400 463.600 200.400 464.200 ;
        RECT 198.400 462.200 199.200 463.600 ;
        RECT 202.800 462.200 203.600 467.000 ;
        RECT 204.400 466.800 205.200 468.400 ;
        RECT 206.000 466.200 206.800 479.800 ;
        RECT 207.600 471.600 208.400 473.200 ;
        RECT 207.700 470.300 208.300 471.600 ;
        RECT 210.800 470.300 211.600 479.800 ;
        RECT 215.000 478.400 215.800 479.800 ;
        RECT 214.000 477.600 215.800 478.400 ;
        RECT 215.000 472.400 215.800 477.600 ;
        RECT 216.400 473.600 217.200 474.400 ;
        RECT 216.600 472.400 217.200 473.600 ;
        RECT 219.600 473.600 220.400 474.400 ;
        RECT 219.600 472.400 220.200 473.600 ;
        RECT 221.000 472.400 221.800 479.800 ;
        RECT 215.000 471.800 216.000 472.400 ;
        RECT 216.600 471.800 218.000 472.400 ;
        RECT 207.700 469.700 211.600 470.300 ;
        RECT 209.200 466.800 210.000 468.400 ;
        RECT 206.000 465.600 207.800 466.200 ;
        RECT 207.000 464.400 207.800 465.600 ;
        RECT 206.000 463.600 207.800 464.400 ;
        RECT 207.000 462.200 207.800 463.600 ;
        RECT 210.800 462.200 211.600 469.700 ;
        RECT 214.000 468.800 214.800 470.400 ;
        RECT 215.400 468.400 216.000 471.800 ;
        RECT 217.200 471.600 218.000 471.800 ;
        RECT 218.800 471.800 220.200 472.400 ;
        RECT 220.800 471.800 221.800 472.400 ;
        RECT 225.200 472.400 226.000 479.800 ;
        RECT 226.800 472.400 227.600 472.600 ;
        RECT 229.600 472.400 231.200 479.800 ;
        RECT 225.200 471.800 227.600 472.400 ;
        RECT 229.200 471.800 231.200 472.400 ;
        RECT 233.400 472.400 234.200 472.600 ;
        RECT 234.800 472.400 235.600 479.800 ;
        RECT 236.400 473.600 238.000 474.400 ;
        RECT 237.200 472.400 237.800 473.600 ;
        RECT 238.600 472.400 239.400 479.800 ;
        RECT 233.400 471.800 235.600 472.400 ;
        RECT 236.400 471.800 237.800 472.400 ;
        RECT 238.400 471.800 239.400 472.400 ;
        RECT 243.400 472.600 244.200 479.800 ;
        RECT 243.400 471.800 245.200 472.600 ;
        RECT 247.600 472.400 248.400 479.800 ;
        RECT 250.800 472.800 251.600 479.800 ;
        RECT 255.600 476.400 256.400 479.800 ;
        RECT 255.400 475.800 256.400 476.400 ;
        RECT 255.400 475.200 256.000 475.800 ;
        RECT 258.800 475.200 259.600 479.800 ;
        RECT 262.000 477.000 262.800 479.800 ;
        RECT 263.600 477.000 264.400 479.800 ;
        RECT 254.000 474.600 256.000 475.200 ;
        RECT 247.600 471.800 250.200 472.400 ;
        RECT 218.800 471.600 219.600 471.800 ;
        RECT 217.300 470.300 217.900 471.600 ;
        RECT 220.800 470.300 221.400 471.800 ;
        RECT 229.200 470.400 229.800 471.800 ;
        RECT 233.400 471.200 234.000 471.800 ;
        RECT 236.400 471.600 237.200 471.800 ;
        RECT 230.600 470.600 234.000 471.200 ;
        RECT 230.600 470.400 231.400 470.600 ;
        RECT 217.300 469.700 221.400 470.300 ;
        RECT 220.800 468.400 221.400 469.700 ;
        RECT 222.000 468.800 222.800 470.400 ;
        RECT 228.400 469.800 229.800 470.400 ;
        RECT 232.800 469.800 233.600 470.000 ;
        RECT 228.400 469.600 230.200 469.800 ;
        RECT 229.200 469.200 230.200 469.600 ;
        RECT 212.400 468.200 213.200 468.400 ;
        RECT 212.400 467.600 214.000 468.200 ;
        RECT 215.400 467.600 218.000 468.400 ;
        RECT 218.800 467.600 221.400 468.400 ;
        RECT 223.600 468.300 224.400 468.400 ;
        RECT 225.200 468.300 226.800 468.400 ;
        RECT 223.600 468.200 226.800 468.300 ;
        RECT 222.800 467.700 226.800 468.200 ;
        RECT 222.800 467.600 224.400 467.700 ;
        RECT 225.200 467.600 226.800 467.700 ;
        RECT 228.000 467.600 228.800 468.400 ;
        RECT 213.200 467.200 214.000 467.600 ;
        RECT 212.600 466.200 216.200 466.600 ;
        RECT 217.200 466.200 217.800 467.600 ;
        RECT 219.000 466.200 219.600 467.600 ;
        RECT 222.800 467.200 223.600 467.600 ;
        RECT 228.200 467.200 228.800 467.600 ;
        RECT 226.800 466.800 227.600 467.000 ;
        RECT 220.600 466.200 224.200 466.600 ;
        RECT 225.200 466.200 227.600 466.800 ;
        RECT 228.200 466.400 229.000 467.200 ;
        RECT 212.400 466.000 216.400 466.200 ;
        RECT 212.400 462.200 213.200 466.000 ;
        RECT 215.600 462.200 216.400 466.000 ;
        RECT 217.200 462.200 218.000 466.200 ;
        RECT 218.800 462.200 219.600 466.200 ;
        RECT 220.400 466.000 224.400 466.200 ;
        RECT 220.400 462.200 221.200 466.000 ;
        RECT 223.600 462.200 224.400 466.000 ;
        RECT 225.200 462.200 226.000 466.200 ;
        RECT 229.600 465.800 230.200 469.200 ;
        RECT 231.000 469.200 233.600 469.800 ;
        RECT 231.000 468.600 231.600 469.200 ;
        RECT 230.800 467.800 231.600 468.600 ;
        RECT 238.400 468.400 239.000 471.800 ;
        RECT 239.600 470.300 240.400 470.400 ;
        RECT 241.200 470.300 242.000 470.400 ;
        RECT 242.800 470.300 243.600 471.200 ;
        RECT 239.600 469.700 243.600 470.300 ;
        RECT 239.600 468.800 240.400 469.700 ;
        RECT 241.200 469.600 242.000 469.700 ;
        RECT 242.800 469.600 243.600 469.700 ;
        RECT 244.400 468.400 245.000 471.800 ;
        RECT 247.600 469.600 248.600 470.400 ;
        RECT 247.800 468.800 248.600 469.600 ;
        RECT 249.600 469.800 250.200 471.800 ;
        RECT 250.800 471.600 251.800 472.800 ;
        RECT 249.600 469.000 250.600 469.800 ;
        RECT 234.000 468.200 235.600 468.400 ;
        RECT 232.200 467.600 235.600 468.200 ;
        RECT 236.400 467.600 239.000 468.400 ;
        RECT 241.200 468.200 242.000 468.400 ;
        RECT 240.400 467.600 242.000 468.200 ;
        RECT 242.800 468.300 243.600 468.400 ;
        RECT 244.400 468.300 245.200 468.400 ;
        RECT 242.800 467.700 245.200 468.300 ;
        RECT 242.800 467.600 243.600 467.700 ;
        RECT 244.400 467.600 245.200 467.700 ;
        RECT 232.200 467.200 232.800 467.600 ;
        RECT 230.800 466.600 232.800 467.200 ;
        RECT 233.400 466.800 234.200 467.000 ;
        RECT 230.800 466.400 232.400 466.600 ;
        RECT 233.400 466.200 235.600 466.800 ;
        RECT 236.600 466.200 237.200 467.600 ;
        RECT 240.400 467.200 241.200 467.600 ;
        RECT 238.200 466.200 241.800 466.600 ;
        RECT 229.600 462.200 231.200 465.800 ;
        RECT 234.800 462.200 235.600 466.200 ;
        RECT 236.400 462.200 237.200 466.200 ;
        RECT 238.000 466.000 242.000 466.200 ;
        RECT 238.000 462.200 238.800 466.000 ;
        RECT 241.200 462.200 242.000 466.000 ;
        RECT 244.400 464.200 245.000 467.600 ;
        RECT 249.600 467.400 250.200 469.000 ;
        RECT 251.200 468.400 251.800 471.600 ;
        RECT 250.800 467.600 251.800 468.400 ;
        RECT 247.600 466.800 250.200 467.400 ;
        RECT 246.000 464.800 246.800 466.400 ;
        RECT 244.400 462.200 245.200 464.200 ;
        RECT 247.600 462.200 248.400 466.800 ;
        RECT 251.200 466.200 251.800 467.600 ;
        RECT 250.800 465.600 251.800 466.200 ;
        RECT 254.000 469.000 254.800 474.600 ;
        RECT 256.600 474.400 260.800 475.200 ;
        RECT 265.200 475.000 266.000 479.800 ;
        RECT 268.400 475.000 269.200 479.800 ;
        RECT 256.600 474.000 257.200 474.400 ;
        RECT 255.600 473.200 257.200 474.000 ;
        RECT 260.200 473.800 266.000 474.400 ;
        RECT 258.200 473.200 259.600 473.800 ;
        RECT 258.200 473.000 264.400 473.200 ;
        RECT 259.000 472.600 264.400 473.000 ;
        RECT 263.600 472.400 264.400 472.600 ;
        RECT 265.400 473.000 266.000 473.800 ;
        RECT 266.600 473.600 269.200 474.400 ;
        RECT 271.600 473.600 272.400 479.800 ;
        RECT 273.200 477.000 274.000 479.800 ;
        RECT 274.800 477.000 275.600 479.800 ;
        RECT 276.400 477.000 277.200 479.800 ;
        RECT 274.800 474.400 279.000 475.200 ;
        RECT 279.600 474.400 280.400 479.800 ;
        RECT 282.800 475.200 283.600 479.800 ;
        RECT 282.800 474.600 285.400 475.200 ;
        RECT 279.600 473.600 282.200 474.400 ;
        RECT 273.200 473.000 274.000 473.200 ;
        RECT 265.400 472.400 274.000 473.000 ;
        RECT 276.400 473.000 277.200 473.200 ;
        RECT 284.800 473.000 285.400 474.600 ;
        RECT 276.400 472.400 285.400 473.000 ;
        RECT 257.200 471.800 258.000 472.400 ;
        RECT 260.600 471.800 261.400 472.000 ;
        RECT 257.200 471.200 284.200 471.800 ;
        RECT 283.400 471.000 284.200 471.200 ;
        RECT 284.800 470.600 285.400 472.400 ;
        RECT 286.000 472.000 286.800 479.800 ;
        RECT 286.000 471.200 287.000 472.000 ;
        RECT 284.800 470.000 285.600 470.600 ;
        RECT 254.000 468.200 262.800 469.000 ;
        RECT 263.400 468.600 265.400 469.400 ;
        RECT 269.200 468.600 272.400 469.400 ;
        RECT 250.800 462.200 251.600 465.600 ;
        RECT 254.000 462.200 254.800 468.200 ;
        RECT 256.400 466.800 259.400 467.600 ;
        RECT 258.600 466.200 259.400 466.800 ;
        RECT 264.600 466.200 265.400 468.600 ;
        RECT 266.800 466.800 267.600 468.400 ;
        RECT 272.000 467.800 272.800 468.000 ;
        RECT 268.400 467.200 272.800 467.800 ;
        RECT 268.400 467.000 269.200 467.200 ;
        RECT 274.800 466.400 275.600 469.200 ;
        RECT 280.600 468.600 284.400 469.400 ;
        RECT 280.600 467.400 281.400 468.600 ;
        RECT 285.000 468.000 285.600 470.000 ;
        RECT 268.400 466.200 269.200 466.400 ;
        RECT 258.600 465.400 261.200 466.200 ;
        RECT 264.600 465.600 269.200 466.200 ;
        RECT 270.000 465.600 271.600 466.400 ;
        RECT 274.600 465.600 275.600 466.400 ;
        RECT 279.600 466.800 281.400 467.400 ;
        RECT 284.400 467.400 285.600 468.000 ;
        RECT 279.600 466.200 280.400 466.800 ;
        RECT 260.400 462.200 261.200 465.400 ;
        RECT 278.000 465.400 280.400 466.200 ;
        RECT 262.000 462.200 262.800 465.000 ;
        RECT 263.600 462.200 264.400 465.000 ;
        RECT 265.200 462.200 266.000 465.000 ;
        RECT 268.400 462.200 269.200 465.000 ;
        RECT 271.600 462.200 272.400 465.000 ;
        RECT 273.200 462.200 274.000 465.000 ;
        RECT 274.800 462.200 275.600 465.000 ;
        RECT 276.400 462.200 277.200 465.000 ;
        RECT 278.000 462.200 278.800 465.400 ;
        RECT 284.400 462.200 285.200 467.400 ;
        RECT 286.200 466.800 287.000 471.200 ;
        RECT 289.200 466.800 290.000 468.400 ;
        RECT 286.000 466.000 287.000 466.800 ;
        RECT 290.800 466.200 291.600 479.800 ;
        RECT 292.400 471.600 293.200 473.200 ;
        RECT 294.600 472.600 295.400 479.800 ;
        RECT 300.400 472.800 301.200 479.800 ;
        RECT 294.600 471.800 296.400 472.600 ;
        RECT 300.200 471.800 301.200 472.800 ;
        RECT 303.600 472.400 304.400 479.800 ;
        RECT 301.800 471.800 304.400 472.400 ;
        RECT 294.000 469.600 294.800 471.200 ;
        RECT 295.600 468.400 296.200 471.800 ;
        RECT 300.200 468.400 300.800 471.800 ;
        RECT 301.800 469.800 302.400 471.800 ;
        RECT 310.000 471.400 310.800 479.800 ;
        RECT 314.400 476.400 315.200 479.800 ;
        RECT 313.200 475.800 315.200 476.400 ;
        RECT 318.800 475.800 319.600 479.800 ;
        RECT 323.000 475.800 324.200 479.800 ;
        RECT 313.200 475.000 314.000 475.800 ;
        RECT 318.800 475.200 319.400 475.800 ;
        RECT 316.600 474.600 320.200 475.200 ;
        RECT 322.800 475.000 323.600 475.800 ;
        RECT 316.600 474.400 317.400 474.600 ;
        RECT 319.400 474.400 320.200 474.600 ;
        RECT 313.200 473.000 314.000 473.200 ;
        RECT 317.800 473.000 318.600 473.200 ;
        RECT 313.200 472.400 318.600 473.000 ;
        RECT 319.200 473.000 321.400 473.600 ;
        RECT 319.200 471.800 319.800 473.000 ;
        RECT 320.600 472.800 321.400 473.000 ;
        RECT 323.000 473.200 324.400 474.000 ;
        RECT 323.000 472.200 323.600 473.200 ;
        RECT 315.000 471.400 319.800 471.800 ;
        RECT 310.000 471.200 319.800 471.400 ;
        RECT 321.200 471.600 323.600 472.200 ;
        RECT 310.000 471.000 315.800 471.200 ;
        RECT 310.000 470.800 315.600 471.000 ;
        RECT 301.400 469.000 302.400 469.800 ;
        RECT 295.600 467.600 296.400 468.400 ;
        RECT 300.200 467.600 301.200 468.400 ;
        RECT 286.000 462.200 286.800 466.000 ;
        RECT 290.800 465.600 292.600 466.200 ;
        RECT 291.800 464.400 292.600 465.600 ;
        RECT 295.600 464.400 296.200 467.600 ;
        RECT 297.200 464.800 298.000 466.400 ;
        RECT 300.200 466.200 300.800 467.600 ;
        RECT 301.800 467.400 302.400 469.000 ;
        RECT 303.400 469.600 304.400 470.400 ;
        RECT 316.400 470.200 317.200 470.400 ;
        RECT 312.200 469.600 317.200 470.200 ;
        RECT 303.400 468.800 304.200 469.600 ;
        RECT 312.200 469.400 313.000 469.600 ;
        RECT 313.800 468.400 314.600 468.600 ;
        RECT 321.200 468.400 321.800 471.600 ;
        RECT 327.600 471.200 328.400 479.800 ;
        RECT 330.000 473.600 330.800 474.400 ;
        RECT 330.000 472.400 330.600 473.600 ;
        RECT 331.400 472.400 332.200 479.800 ;
        RECT 338.200 478.400 339.000 479.800 ;
        RECT 337.200 477.600 339.000 478.400 ;
        RECT 329.200 471.800 330.600 472.400 ;
        RECT 331.200 471.800 332.200 472.400 ;
        RECT 338.200 472.400 339.000 477.600 ;
        RECT 339.600 473.600 340.400 474.400 ;
        RECT 339.800 472.400 340.400 473.600 ;
        RECT 338.200 471.800 339.200 472.400 ;
        RECT 339.800 472.300 341.200 472.400 ;
        RECT 342.000 472.300 342.800 479.800 ;
        RECT 339.800 471.800 342.800 472.300 ;
        RECT 347.800 472.400 348.600 479.800 ;
        RECT 353.800 476.400 354.600 479.800 ;
        RECT 353.800 475.600 355.600 476.400 ;
        RECT 349.200 473.600 350.000 474.400 ;
        RECT 349.400 472.400 350.000 473.600 ;
        RECT 352.400 473.600 353.200 474.400 ;
        RECT 352.400 472.400 353.000 473.600 ;
        RECT 353.800 472.400 354.600 475.600 ;
        RECT 361.800 474.400 362.600 479.800 ;
        RECT 366.000 475.000 366.800 479.000 ;
        RECT 361.200 473.600 362.600 474.400 ;
        RECT 361.800 472.800 362.600 473.600 ;
        RECT 347.800 471.800 348.800 472.400 ;
        RECT 349.400 471.800 350.800 472.400 ;
        RECT 329.200 471.600 330.000 471.800 ;
        RECT 324.200 470.600 328.400 471.200 ;
        RECT 324.200 470.400 325.000 470.600 ;
        RECT 325.800 469.800 326.600 470.000 ;
        RECT 322.800 469.200 326.600 469.800 ;
        RECT 322.800 469.000 323.600 469.200 ;
        RECT 310.800 467.800 321.800 468.400 ;
        RECT 310.800 467.600 312.400 467.800 ;
        RECT 301.800 466.800 304.400 467.400 ;
        RECT 300.200 465.600 301.200 466.200 ;
        RECT 291.800 463.600 293.200 464.400 ;
        RECT 291.800 462.200 292.600 463.600 ;
        RECT 295.600 462.200 296.400 464.400 ;
        RECT 300.400 462.200 301.200 465.600 ;
        RECT 303.600 462.200 304.400 466.800 ;
        RECT 310.000 462.200 310.800 467.000 ;
        RECT 315.000 466.400 315.600 467.800 ;
        RECT 320.600 467.600 321.400 467.800 ;
        RECT 327.600 467.200 328.400 470.600 ;
        RECT 331.200 470.400 331.800 471.800 ;
        RECT 330.800 469.600 331.800 470.400 ;
        RECT 331.200 468.400 331.800 469.600 ;
        RECT 332.400 468.800 333.200 470.400 ;
        RECT 334.000 470.300 334.800 470.400 ;
        RECT 337.200 470.300 338.000 470.400 ;
        RECT 334.000 469.700 338.000 470.300 ;
        RECT 334.000 469.600 334.800 469.700 ;
        RECT 334.100 468.400 334.700 469.600 ;
        RECT 337.200 468.800 338.000 469.700 ;
        RECT 338.600 468.400 339.200 471.800 ;
        RECT 340.400 471.700 342.800 471.800 ;
        RECT 340.400 471.600 341.200 471.700 ;
        RECT 329.200 467.600 331.800 468.400 ;
        RECT 334.000 468.200 334.800 468.400 ;
        RECT 333.200 467.600 334.800 468.200 ;
        RECT 335.600 468.200 336.400 468.400 ;
        RECT 335.600 467.600 337.200 468.200 ;
        RECT 338.600 467.600 341.200 468.400 ;
        RECT 324.600 466.600 328.400 467.200 ;
        RECT 324.600 466.400 325.400 466.600 ;
        RECT 313.200 464.200 314.000 465.000 ;
        RECT 314.800 464.800 315.600 466.400 ;
        RECT 316.600 465.400 317.400 465.600 ;
        RECT 316.600 464.800 319.400 465.400 ;
        RECT 318.800 464.200 319.400 464.800 ;
        RECT 322.800 464.200 323.600 465.000 ;
        RECT 313.200 463.600 315.200 464.200 ;
        RECT 314.400 462.200 315.200 463.600 ;
        RECT 318.800 462.200 319.600 464.200 ;
        RECT 322.800 463.600 324.200 464.200 ;
        RECT 323.000 462.200 324.200 463.600 ;
        RECT 327.600 462.200 328.400 466.600 ;
        RECT 329.400 466.200 330.000 467.600 ;
        RECT 333.200 467.200 334.000 467.600 ;
        RECT 336.400 467.200 337.200 467.600 ;
        RECT 331.000 466.200 334.600 466.600 ;
        RECT 335.800 466.200 339.400 466.600 ;
        RECT 340.400 466.200 341.000 467.600 ;
        RECT 329.200 462.200 330.000 466.200 ;
        RECT 330.800 466.000 334.800 466.200 ;
        RECT 330.800 462.200 331.600 466.000 ;
        RECT 334.000 462.200 334.800 466.000 ;
        RECT 335.600 466.000 339.600 466.200 ;
        RECT 335.600 462.200 336.400 466.000 ;
        RECT 338.800 462.200 339.600 466.000 ;
        RECT 340.400 462.200 341.200 466.200 ;
        RECT 342.000 462.200 342.800 471.700 ;
        RECT 346.800 468.800 347.600 470.400 ;
        RECT 348.200 470.300 348.800 471.800 ;
        RECT 350.000 471.600 350.800 471.800 ;
        RECT 351.600 471.800 353.000 472.400 ;
        RECT 353.600 471.800 354.600 472.400 ;
        RECT 361.000 472.200 362.600 472.800 ;
        RECT 351.600 471.600 352.400 471.800 ;
        RECT 351.700 470.300 352.300 471.600 ;
        RECT 348.200 469.700 352.300 470.300 ;
        RECT 348.200 468.400 348.800 469.700 ;
        RECT 353.600 468.400 354.200 471.800 ;
        RECT 354.800 468.800 355.600 470.400 ;
        RECT 356.400 470.300 357.200 470.400 ;
        RECT 359.600 470.300 360.400 471.200 ;
        RECT 356.400 469.700 360.400 470.300 ;
        RECT 356.400 469.600 357.200 469.700 ;
        RECT 359.600 469.600 360.400 469.700 ;
        RECT 361.000 468.400 361.600 472.200 ;
        RECT 366.200 471.600 366.800 475.000 ;
        RECT 363.000 471.000 366.800 471.600 ;
        RECT 367.600 471.400 368.400 479.800 ;
        RECT 372.000 476.400 372.800 479.800 ;
        RECT 370.800 475.800 372.800 476.400 ;
        RECT 376.400 475.800 377.200 479.800 ;
        RECT 380.600 475.800 381.800 479.800 ;
        RECT 370.800 475.000 371.600 475.800 ;
        RECT 376.400 475.200 377.000 475.800 ;
        RECT 374.200 474.600 377.800 475.200 ;
        RECT 380.400 475.000 381.200 475.800 ;
        RECT 374.200 474.400 375.000 474.600 ;
        RECT 377.000 474.400 377.800 474.600 ;
        RECT 370.800 473.000 371.600 473.200 ;
        RECT 375.400 473.000 376.200 473.200 ;
        RECT 370.800 472.400 376.200 473.000 ;
        RECT 376.800 473.000 379.000 473.600 ;
        RECT 376.800 471.800 377.400 473.000 ;
        RECT 378.200 472.800 379.000 473.000 ;
        RECT 380.600 473.200 382.000 474.000 ;
        RECT 380.600 472.200 381.200 473.200 ;
        RECT 372.600 471.400 377.400 471.800 ;
        RECT 367.600 471.200 377.400 471.400 ;
        RECT 378.800 471.600 381.200 472.200 ;
        RECT 367.600 471.000 373.400 471.200 ;
        RECT 363.000 469.000 363.600 471.000 ;
        RECT 367.600 470.800 373.200 471.000 ;
        RECT 345.200 468.300 346.000 468.400 ;
        RECT 343.700 468.200 346.000 468.300 ;
        RECT 343.700 467.700 346.800 468.200 ;
        RECT 343.700 466.400 344.300 467.700 ;
        RECT 345.200 467.600 346.800 467.700 ;
        RECT 348.200 467.600 350.800 468.400 ;
        RECT 351.600 467.600 354.200 468.400 ;
        RECT 356.400 468.300 357.200 468.400 ;
        RECT 358.000 468.300 358.800 468.400 ;
        RECT 356.400 468.200 358.800 468.300 ;
        RECT 355.600 467.700 358.800 468.200 ;
        RECT 355.600 467.600 357.200 467.700 ;
        RECT 358.000 467.600 358.800 467.700 ;
        RECT 359.600 467.600 361.600 468.400 ;
        RECT 362.200 468.200 363.600 469.000 ;
        RECT 364.400 468.800 365.200 470.400 ;
        RECT 366.000 468.800 366.800 470.400 ;
        RECT 374.000 470.200 374.800 470.400 ;
        RECT 369.800 469.600 374.800 470.200 ;
        RECT 369.800 469.400 370.600 469.600 ;
        RECT 371.400 468.400 372.200 468.600 ;
        RECT 378.800 468.400 379.400 471.600 ;
        RECT 385.200 471.200 386.000 479.800 ;
        RECT 388.400 472.800 389.200 479.800 ;
        RECT 381.800 470.600 386.000 471.200 ;
        RECT 381.800 470.400 382.600 470.600 ;
        RECT 383.400 469.800 384.200 470.000 ;
        RECT 380.400 469.200 384.200 469.800 ;
        RECT 380.400 469.000 381.200 469.200 ;
        RECT 346.000 467.200 346.800 467.600 ;
        RECT 343.600 464.800 344.400 466.400 ;
        RECT 345.400 466.200 349.000 466.600 ;
        RECT 350.000 466.200 350.600 467.600 ;
        RECT 351.800 466.200 352.400 467.600 ;
        RECT 355.600 467.200 356.400 467.600 ;
        RECT 361.000 467.000 361.600 467.600 ;
        RECT 362.600 467.800 363.600 468.200 ;
        RECT 368.400 467.800 379.400 468.400 ;
        RECT 362.600 467.200 366.800 467.800 ;
        RECT 368.400 467.600 370.000 467.800 ;
        RECT 372.400 467.600 373.200 467.800 ;
        RECT 378.200 467.600 379.000 467.800 ;
        RECT 361.000 466.600 361.800 467.000 ;
        RECT 353.400 466.200 357.000 466.600 ;
        RECT 345.200 466.000 349.200 466.200 ;
        RECT 345.200 462.200 346.000 466.000 ;
        RECT 348.400 462.200 349.200 466.000 ;
        RECT 350.000 462.200 350.800 466.200 ;
        RECT 351.600 462.200 352.400 466.200 ;
        RECT 353.200 466.000 357.200 466.200 ;
        RECT 361.000 466.000 362.600 466.600 ;
        RECT 353.200 462.200 354.000 466.000 ;
        RECT 356.400 462.200 357.200 466.000 ;
        RECT 361.800 463.000 362.600 466.000 ;
        RECT 366.200 465.000 366.800 467.200 ;
        RECT 366.000 463.000 366.800 465.000 ;
        RECT 367.600 462.200 368.400 467.000 ;
        RECT 372.600 465.600 373.200 467.600 ;
        RECT 385.200 467.200 386.000 470.600 ;
        RECT 382.200 466.600 386.000 467.200 ;
        RECT 382.200 466.400 383.000 466.600 ;
        RECT 370.800 464.200 371.600 465.000 ;
        RECT 372.400 464.800 373.200 465.600 ;
        RECT 374.200 465.400 375.000 465.600 ;
        RECT 374.200 464.800 377.000 465.400 ;
        RECT 376.400 464.200 377.000 464.800 ;
        RECT 380.400 464.200 381.200 465.000 ;
        RECT 370.800 463.600 372.800 464.200 ;
        RECT 372.000 462.200 372.800 463.600 ;
        RECT 376.400 462.200 377.200 464.200 ;
        RECT 380.400 463.600 381.800 464.200 ;
        RECT 380.600 462.200 381.800 463.600 ;
        RECT 385.200 462.200 386.000 466.600 ;
        RECT 388.200 471.800 389.200 472.800 ;
        RECT 391.600 472.400 392.400 479.800 ;
        RECT 394.000 473.600 394.800 474.400 ;
        RECT 394.000 472.400 394.600 473.600 ;
        RECT 395.400 472.400 396.200 479.800 ;
        RECT 389.800 471.800 392.400 472.400 ;
        RECT 393.200 471.800 394.600 472.400 ;
        RECT 395.200 471.800 396.200 472.400 ;
        RECT 388.200 468.400 388.800 471.800 ;
        RECT 389.800 469.800 390.400 471.800 ;
        RECT 393.200 471.600 394.000 471.800 ;
        RECT 389.400 469.000 390.400 469.800 ;
        RECT 388.200 467.600 389.200 468.400 ;
        RECT 388.200 466.200 388.800 467.600 ;
        RECT 389.800 467.400 390.400 469.000 ;
        RECT 391.400 469.600 392.400 470.400 ;
        RECT 391.400 468.800 392.200 469.600 ;
        RECT 395.200 468.400 395.800 471.800 ;
        RECT 396.400 468.800 397.200 470.400 ;
        RECT 393.200 467.600 395.800 468.400 ;
        RECT 398.000 468.200 398.800 468.400 ;
        RECT 397.200 467.600 398.800 468.200 ;
        RECT 389.800 466.800 392.400 467.400 ;
        RECT 388.200 465.600 389.200 466.200 ;
        RECT 388.400 462.200 389.200 465.600 ;
        RECT 391.600 462.200 392.400 466.800 ;
        RECT 393.400 466.200 394.000 467.600 ;
        RECT 397.200 467.200 398.000 467.600 ;
        RECT 395.000 466.200 398.600 466.600 ;
        RECT 393.200 462.200 394.000 466.200 ;
        RECT 394.800 466.000 398.800 466.200 ;
        RECT 394.800 462.200 395.600 466.000 ;
        RECT 398.000 462.200 398.800 466.000 ;
        RECT 399.600 464.800 400.400 466.400 ;
        RECT 401.200 462.200 402.000 479.800 ;
        RECT 402.800 471.400 403.600 479.800 ;
        RECT 407.200 476.400 408.000 479.800 ;
        RECT 406.000 475.800 408.000 476.400 ;
        RECT 411.600 475.800 412.400 479.800 ;
        RECT 415.800 475.800 417.000 479.800 ;
        RECT 406.000 475.000 406.800 475.800 ;
        RECT 411.600 475.200 412.200 475.800 ;
        RECT 409.400 474.600 413.000 475.200 ;
        RECT 415.600 475.000 416.400 475.800 ;
        RECT 409.400 474.400 410.200 474.600 ;
        RECT 412.200 474.400 413.000 474.600 ;
        RECT 406.000 473.000 406.800 473.200 ;
        RECT 410.600 473.000 411.400 473.200 ;
        RECT 406.000 472.400 411.400 473.000 ;
        RECT 412.000 473.000 414.200 473.600 ;
        RECT 412.000 471.800 412.600 473.000 ;
        RECT 413.400 472.800 414.200 473.000 ;
        RECT 415.800 473.200 417.200 474.000 ;
        RECT 415.800 472.200 416.400 473.200 ;
        RECT 407.800 471.400 412.600 471.800 ;
        RECT 402.800 471.200 412.600 471.400 ;
        RECT 414.000 471.600 416.400 472.200 ;
        RECT 402.800 471.000 408.600 471.200 ;
        RECT 402.800 470.800 408.400 471.000 ;
        RECT 409.200 470.200 410.000 470.400 ;
        RECT 405.000 469.600 410.000 470.200 ;
        RECT 405.000 469.400 405.800 469.600 ;
        RECT 406.600 468.400 407.400 468.600 ;
        RECT 414.000 468.400 414.600 471.600 ;
        RECT 420.400 471.200 421.200 479.800 ;
        RECT 417.000 470.600 421.200 471.200 ;
        RECT 417.000 470.400 417.800 470.600 ;
        RECT 418.600 469.800 419.400 470.000 ;
        RECT 415.600 469.200 419.400 469.800 ;
        RECT 415.600 469.000 416.400 469.200 ;
        RECT 403.600 467.800 414.600 468.400 ;
        RECT 403.600 467.600 405.200 467.800 ;
        RECT 402.800 462.200 403.600 467.000 ;
        RECT 407.800 465.600 408.400 467.800 ;
        RECT 413.400 467.600 414.200 467.800 ;
        RECT 420.400 467.200 421.200 470.600 ;
        RECT 417.400 466.600 421.200 467.200 ;
        RECT 422.000 466.800 422.800 468.400 ;
        RECT 417.400 466.400 418.200 466.600 ;
        RECT 406.000 464.200 406.800 465.000 ;
        RECT 407.600 464.800 408.400 465.600 ;
        RECT 409.400 465.400 410.200 465.600 ;
        RECT 409.400 464.800 412.200 465.400 ;
        RECT 411.600 464.200 412.200 464.800 ;
        RECT 415.600 464.200 416.400 465.000 ;
        RECT 406.000 463.600 408.000 464.200 ;
        RECT 407.200 462.200 408.000 463.600 ;
        RECT 411.600 462.200 412.400 464.200 ;
        RECT 415.600 463.600 417.000 464.200 ;
        RECT 415.800 462.200 417.000 463.600 ;
        RECT 420.400 462.200 421.200 466.600 ;
        RECT 423.600 466.200 424.400 479.800 ;
        RECT 425.200 472.300 426.000 473.200 ;
        RECT 426.800 472.300 427.600 472.400 ;
        RECT 425.200 471.700 427.600 472.300 ;
        RECT 425.200 471.600 426.000 471.700 ;
        RECT 426.800 471.600 427.600 471.700 ;
        RECT 425.200 468.300 426.000 468.400 ;
        RECT 426.800 468.300 427.600 468.400 ;
        RECT 425.200 467.700 427.600 468.300 ;
        RECT 425.200 467.600 426.000 467.700 ;
        RECT 426.800 466.800 427.600 467.700 ;
        RECT 428.400 466.200 429.200 479.800 ;
        RECT 430.000 471.600 430.800 473.200 ;
        RECT 434.200 472.400 435.000 479.800 ;
        RECT 435.600 473.600 436.400 474.400 ;
        RECT 435.800 472.400 436.400 473.600 ;
        RECT 438.800 473.600 439.600 474.400 ;
        RECT 438.800 472.400 439.400 473.600 ;
        RECT 440.200 472.400 441.000 479.800 ;
        RECT 434.200 471.800 435.200 472.400 ;
        RECT 435.800 471.800 437.200 472.400 ;
        RECT 434.600 470.400 435.200 471.800 ;
        RECT 436.400 471.600 437.200 471.800 ;
        RECT 438.000 471.800 439.400 472.400 ;
        RECT 440.000 471.800 441.000 472.400 ;
        RECT 444.400 475.000 445.200 479.000 ;
        RECT 448.600 478.400 449.400 479.800 ;
        RECT 447.600 477.600 449.400 478.400 ;
        RECT 438.000 471.600 438.800 471.800 ;
        RECT 433.200 468.800 434.000 470.400 ;
        RECT 434.600 469.600 435.600 470.400 ;
        RECT 436.500 470.300 437.100 471.600 ;
        RECT 440.000 470.300 440.600 471.800 ;
        RECT 444.400 471.600 445.000 475.000 ;
        RECT 448.600 472.800 449.400 477.600 ;
        RECT 462.600 472.800 463.400 479.800 ;
        RECT 466.800 475.000 467.600 479.000 ;
        RECT 448.600 472.200 450.200 472.800 ;
        RECT 444.400 471.000 448.200 471.600 ;
        RECT 436.500 469.700 440.600 470.300 ;
        RECT 434.600 468.400 435.200 469.600 ;
        RECT 440.000 468.400 440.600 469.700 ;
        RECT 441.200 468.800 442.000 470.400 ;
        RECT 444.400 468.800 445.200 470.400 ;
        RECT 446.000 468.800 446.800 470.400 ;
        RECT 447.600 469.000 448.200 471.000 ;
        RECT 431.600 468.200 432.400 468.400 ;
        RECT 431.600 467.600 433.200 468.200 ;
        RECT 434.600 467.600 437.200 468.400 ;
        RECT 438.000 467.600 440.600 468.400 ;
        RECT 442.800 468.200 443.600 468.400 ;
        RECT 442.000 467.600 443.600 468.200 ;
        RECT 447.600 468.200 449.000 469.000 ;
        RECT 449.600 468.400 450.200 472.200 ;
        RECT 461.800 472.200 463.400 472.800 ;
        RECT 450.800 470.300 451.600 471.200 ;
        RECT 460.400 470.300 461.200 471.200 ;
        RECT 450.800 469.700 461.200 470.300 ;
        RECT 450.800 469.600 451.600 469.700 ;
        RECT 460.400 469.600 461.200 469.700 ;
        RECT 461.800 468.400 462.400 472.200 ;
        RECT 467.000 471.600 467.600 475.000 ;
        RECT 463.800 471.000 467.600 471.600 ;
        RECT 463.800 469.000 464.400 471.000 ;
        RECT 447.600 467.800 448.600 468.200 ;
        RECT 432.400 467.200 433.200 467.600 ;
        RECT 431.800 466.200 435.400 466.600 ;
        RECT 436.400 466.200 437.000 467.600 ;
        RECT 438.200 466.200 438.800 467.600 ;
        RECT 442.000 467.200 442.800 467.600 ;
        RECT 444.400 467.200 448.600 467.800 ;
        RECT 449.600 467.600 451.600 468.400 ;
        RECT 452.400 468.300 453.200 468.400 ;
        RECT 460.400 468.300 462.400 468.400 ;
        RECT 452.400 467.700 462.400 468.300 ;
        RECT 463.000 468.200 464.400 469.000 ;
        RECT 465.200 468.800 466.000 470.400 ;
        RECT 466.800 468.800 467.600 470.400 ;
        RECT 452.400 467.600 453.200 467.700 ;
        RECT 460.400 467.600 462.400 467.700 ;
        RECT 439.800 466.200 443.400 466.600 ;
        RECT 423.600 465.600 425.400 466.200 ;
        RECT 428.400 465.600 430.200 466.200 ;
        RECT 424.600 464.400 425.400 465.600 ;
        RECT 423.600 463.600 425.400 464.400 ;
        RECT 424.600 462.200 425.400 463.600 ;
        RECT 429.400 464.400 430.200 465.600 ;
        RECT 431.600 466.000 435.600 466.200 ;
        RECT 429.400 463.600 430.800 464.400 ;
        RECT 429.400 462.200 430.200 463.600 ;
        RECT 431.600 462.200 432.400 466.000 ;
        RECT 434.800 462.200 435.600 466.000 ;
        RECT 436.400 462.200 437.200 466.200 ;
        RECT 438.000 462.200 438.800 466.200 ;
        RECT 439.600 466.000 443.600 466.200 ;
        RECT 439.600 462.200 440.400 466.000 ;
        RECT 442.800 462.200 443.600 466.000 ;
        RECT 444.400 465.000 445.000 467.200 ;
        RECT 449.600 467.000 450.200 467.600 ;
        RECT 449.400 466.600 450.200 467.000 ;
        RECT 448.600 466.000 450.200 466.600 ;
        RECT 461.800 467.000 462.400 467.600 ;
        RECT 463.400 467.800 464.400 468.200 ;
        RECT 463.400 467.200 467.600 467.800 ;
        RECT 461.800 466.600 462.600 467.000 ;
        RECT 461.800 466.000 463.400 466.600 ;
        RECT 444.400 463.000 445.200 465.000 ;
        RECT 448.600 463.000 449.400 466.000 ;
        RECT 462.600 463.000 463.400 466.000 ;
        RECT 467.000 465.000 467.600 467.200 ;
        RECT 468.400 466.800 469.200 468.400 ;
        RECT 470.000 466.200 470.800 479.800 ;
        RECT 471.600 471.600 472.400 473.200 ;
        RECT 475.800 472.400 476.600 479.800 ;
        RECT 477.200 473.600 478.000 474.400 ;
        RECT 477.400 472.400 478.000 473.600 ;
        RECT 481.200 472.800 482.000 479.800 ;
        RECT 475.800 471.800 476.800 472.400 ;
        RECT 477.400 471.800 478.800 472.400 ;
        RECT 474.800 468.800 475.600 470.400 ;
        RECT 476.200 468.400 476.800 471.800 ;
        RECT 478.000 471.600 478.800 471.800 ;
        RECT 481.000 471.600 482.000 472.800 ;
        RECT 484.400 472.400 485.200 479.800 ;
        RECT 482.600 471.800 485.200 472.400 ;
        RECT 486.000 475.000 486.800 479.000 ;
        RECT 490.200 478.400 491.000 479.800 ;
        RECT 489.200 477.600 491.000 478.400 ;
        RECT 481.000 468.400 481.600 471.600 ;
        RECT 482.600 469.800 483.200 471.800 ;
        RECT 486.000 471.600 486.600 475.000 ;
        RECT 490.200 472.800 491.000 477.600 ;
        RECT 490.200 472.200 491.800 472.800 ;
        RECT 486.000 471.000 489.800 471.600 ;
        RECT 482.200 469.000 483.200 469.800 ;
        RECT 473.200 468.200 474.000 468.400 ;
        RECT 473.200 467.600 474.800 468.200 ;
        RECT 476.200 467.600 478.800 468.400 ;
        RECT 481.000 467.600 482.000 468.400 ;
        RECT 474.000 467.200 474.800 467.600 ;
        RECT 473.400 466.200 477.000 466.600 ;
        RECT 478.000 466.200 478.600 467.600 ;
        RECT 481.000 466.200 481.600 467.600 ;
        RECT 482.600 467.400 483.200 469.000 ;
        RECT 484.200 469.600 485.200 470.400 ;
        RECT 484.200 468.800 485.000 469.600 ;
        RECT 486.000 468.800 486.800 470.400 ;
        RECT 487.600 468.800 488.400 470.400 ;
        RECT 489.200 469.000 489.800 471.000 ;
        RECT 489.200 468.200 490.600 469.000 ;
        RECT 491.200 468.400 491.800 472.200 ;
        RECT 492.400 470.300 493.200 471.200 ;
        RECT 495.600 470.300 496.400 470.400 ;
        RECT 492.400 469.700 496.400 470.300 ;
        RECT 492.400 469.600 493.200 469.700 ;
        RECT 495.600 469.600 496.400 469.700 ;
        RECT 489.200 467.800 490.200 468.200 ;
        RECT 482.600 466.800 485.200 467.400 ;
        RECT 470.000 465.600 471.800 466.200 ;
        RECT 466.800 463.000 467.600 465.000 ;
        RECT 471.000 464.400 471.800 465.600 ;
        RECT 470.000 463.600 471.800 464.400 ;
        RECT 471.000 462.200 471.800 463.600 ;
        RECT 473.200 466.000 477.200 466.200 ;
        RECT 473.200 462.200 474.000 466.000 ;
        RECT 476.400 462.200 477.200 466.000 ;
        RECT 478.000 462.200 478.800 466.200 ;
        RECT 481.000 465.600 482.000 466.200 ;
        RECT 481.200 462.200 482.000 465.600 ;
        RECT 484.400 462.200 485.200 466.800 ;
        RECT 486.000 467.200 490.200 467.800 ;
        RECT 491.200 467.600 493.200 468.400 ;
        RECT 486.000 465.000 486.600 467.200 ;
        RECT 491.200 467.000 491.800 467.600 ;
        RECT 491.000 466.600 491.800 467.000 ;
        RECT 490.200 466.000 491.800 466.600 ;
        RECT 486.000 463.000 486.800 465.000 ;
        RECT 490.200 463.000 491.000 466.000 ;
        RECT 495.600 464.800 496.400 466.400 ;
        RECT 497.200 462.200 498.000 479.800 ;
        RECT 501.400 472.400 502.200 479.800 ;
        RECT 502.800 473.600 503.600 474.400 ;
        RECT 503.000 472.400 503.600 473.600 ;
        RECT 501.400 471.800 502.400 472.400 ;
        RECT 503.000 471.800 504.400 472.400 ;
        RECT 501.800 470.400 502.400 471.800 ;
        RECT 503.600 471.600 504.400 471.800 ;
        RECT 500.400 468.800 501.200 470.400 ;
        RECT 501.800 469.600 502.800 470.400 ;
        RECT 501.800 468.400 502.400 469.600 ;
        RECT 498.800 468.200 499.600 468.400 ;
        RECT 498.800 467.600 500.400 468.200 ;
        RECT 501.800 467.600 504.400 468.400 ;
        RECT 499.600 467.200 500.400 467.600 ;
        RECT 499.000 466.200 502.600 466.600 ;
        RECT 503.600 466.200 504.200 467.600 ;
        RECT 505.200 466.800 506.000 468.400 ;
        RECT 506.800 466.200 507.600 479.800 ;
        RECT 510.600 478.400 511.400 479.800 ;
        RECT 517.400 478.400 518.200 479.800 ;
        RECT 510.600 477.600 512.400 478.400 ;
        RECT 516.400 477.600 518.200 478.400 ;
        RECT 508.400 471.600 509.200 473.200 ;
        RECT 510.600 472.600 511.400 477.600 ;
        RECT 517.400 472.600 518.200 477.600 ;
        RECT 510.600 471.800 512.400 472.600 ;
        RECT 516.400 471.800 518.200 472.600 ;
        RECT 519.600 475.000 520.400 479.000 ;
        RECT 523.800 478.400 524.600 479.800 ;
        RECT 523.800 477.600 525.200 478.400 ;
        RECT 508.500 470.300 509.100 471.600 ;
        RECT 510.000 470.300 510.800 471.200 ;
        RECT 508.500 469.700 510.800 470.300 ;
        RECT 510.000 469.600 510.800 469.700 ;
        RECT 511.600 468.400 512.200 471.800 ;
        RECT 516.600 468.400 517.200 471.800 ;
        RECT 519.600 471.600 520.200 475.000 ;
        RECT 523.800 472.800 524.600 477.600 ;
        RECT 523.800 472.200 525.400 472.800 ;
        RECT 518.000 469.600 518.800 471.200 ;
        RECT 519.600 471.000 523.400 471.600 ;
        RECT 519.600 468.800 520.400 470.400 ;
        RECT 521.200 468.800 522.000 470.400 ;
        RECT 522.800 469.000 523.400 471.000 ;
        RECT 511.600 467.600 512.400 468.400 ;
        RECT 516.400 467.600 517.200 468.400 ;
        RECT 522.800 468.200 524.200 469.000 ;
        RECT 524.800 468.400 525.400 472.200 ;
        RECT 529.800 472.600 530.600 479.800 ;
        RECT 529.800 471.800 531.600 472.600 ;
        RECT 526.000 469.600 526.800 471.200 ;
        RECT 529.200 469.600 530.000 471.200 ;
        RECT 530.800 470.400 531.400 471.800 ;
        RECT 530.800 469.600 531.600 470.400 ;
        RECT 530.800 468.400 531.400 469.600 ;
        RECT 522.800 467.800 523.800 468.200 ;
        RECT 498.800 466.000 502.800 466.200 ;
        RECT 498.800 462.200 499.600 466.000 ;
        RECT 502.000 462.200 502.800 466.000 ;
        RECT 503.600 462.200 504.400 466.200 ;
        RECT 506.800 465.600 508.600 466.200 ;
        RECT 507.800 462.200 508.600 465.600 ;
        RECT 511.600 464.200 512.200 467.600 ;
        RECT 513.200 466.300 514.000 466.400 ;
        RECT 514.800 466.300 515.600 466.400 ;
        RECT 513.200 465.700 515.600 466.300 ;
        RECT 513.200 464.800 514.000 465.700 ;
        RECT 514.800 464.800 515.600 465.700 ;
        RECT 516.600 464.200 517.200 467.600 ;
        RECT 511.600 462.200 512.400 464.200 ;
        RECT 516.400 462.200 517.200 464.200 ;
        RECT 519.600 467.200 523.800 467.800 ;
        RECT 524.800 467.600 526.800 468.400 ;
        RECT 530.800 467.600 531.600 468.400 ;
        RECT 534.000 468.300 534.800 479.800 ;
        RECT 537.200 472.400 538.000 479.800 ;
        RECT 538.800 472.400 539.600 472.600 ;
        RECT 541.600 472.400 543.200 479.800 ;
        RECT 537.200 471.800 539.600 472.400 ;
        RECT 541.200 471.800 543.200 472.400 ;
        RECT 545.400 472.400 546.200 472.600 ;
        RECT 546.800 472.400 547.600 479.800 ;
        RECT 545.400 471.800 547.600 472.400 ;
        RECT 549.000 472.600 549.800 479.800 ;
        RECT 549.000 471.800 550.800 472.600 ;
        RECT 541.200 470.400 541.800 471.800 ;
        RECT 545.400 471.200 546.000 471.800 ;
        RECT 542.600 470.600 546.000 471.200 ;
        RECT 542.600 470.400 543.400 470.600 ;
        RECT 540.400 469.800 541.800 470.400 ;
        RECT 544.800 469.800 545.600 470.000 ;
        RECT 540.400 469.600 542.200 469.800 ;
        RECT 541.200 469.200 542.200 469.600 ;
        RECT 537.200 468.300 538.800 468.400 ;
        RECT 534.000 467.700 538.800 468.300 ;
        RECT 519.600 465.000 520.200 467.200 ;
        RECT 524.800 467.000 525.400 467.600 ;
        RECT 524.600 466.600 525.400 467.000 ;
        RECT 523.800 466.000 525.400 466.600 ;
        RECT 519.600 463.000 520.400 465.000 ;
        RECT 523.800 463.000 524.600 466.000 ;
        RECT 530.800 464.200 531.400 467.600 ;
        RECT 532.400 466.300 533.200 466.400 ;
        RECT 534.000 466.300 534.800 467.700 ;
        RECT 537.200 467.600 538.800 467.700 ;
        RECT 540.000 467.600 540.800 468.400 ;
        RECT 540.200 467.200 540.800 467.600 ;
        RECT 538.800 466.800 539.600 467.000 ;
        RECT 532.400 465.700 534.800 466.300 ;
        RECT 532.400 464.800 533.200 465.700 ;
        RECT 530.800 462.200 531.600 464.200 ;
        RECT 534.000 462.200 534.800 465.700 ;
        RECT 535.600 464.800 536.400 466.400 ;
        RECT 537.200 466.200 539.600 466.800 ;
        RECT 540.200 466.400 541.000 467.200 ;
        RECT 537.200 462.200 538.000 466.200 ;
        RECT 541.600 465.800 542.200 469.200 ;
        RECT 543.000 469.200 545.600 469.800 ;
        RECT 548.400 469.600 549.200 471.200 ;
        RECT 543.000 468.600 543.600 469.200 ;
        RECT 542.800 467.800 543.600 468.600 ;
        RECT 550.000 468.400 550.600 471.800 ;
        RECT 546.000 468.300 547.600 468.400 ;
        RECT 550.000 468.300 550.800 468.400 ;
        RECT 546.000 468.200 550.800 468.300 ;
        RECT 544.200 467.700 550.800 468.200 ;
        RECT 544.200 467.600 547.600 467.700 ;
        RECT 550.000 467.600 550.800 467.700 ;
        RECT 544.200 467.200 544.800 467.600 ;
        RECT 542.800 466.600 544.800 467.200 ;
        RECT 545.400 466.800 546.200 467.000 ;
        RECT 542.800 466.400 544.400 466.600 ;
        RECT 545.400 466.200 547.600 466.800 ;
        RECT 541.600 464.400 543.200 465.800 ;
        RECT 541.600 463.600 544.400 464.400 ;
        RECT 541.600 462.200 543.200 463.600 ;
        RECT 546.800 462.200 547.600 466.200 ;
        RECT 550.000 464.200 550.600 467.600 ;
        RECT 551.600 466.300 552.400 466.400 ;
        RECT 553.200 466.300 554.000 479.800 ;
        RECT 556.400 472.400 557.200 479.800 ;
        RECT 557.800 472.400 558.600 472.600 ;
        RECT 556.400 471.800 558.600 472.400 ;
        RECT 560.800 472.400 562.400 479.800 ;
        RECT 564.400 472.400 565.200 472.600 ;
        RECT 566.000 472.400 566.800 479.800 ;
        RECT 560.800 471.800 562.800 472.400 ;
        RECT 564.400 471.800 566.800 472.400 ;
        RECT 567.600 472.400 568.400 479.800 ;
        RECT 569.000 472.400 569.800 472.600 ;
        RECT 567.600 471.800 569.800 472.400 ;
        RECT 572.000 472.400 573.600 479.800 ;
        RECT 575.600 472.400 576.400 472.600 ;
        RECT 577.200 472.400 578.000 479.800 ;
        RECT 572.000 471.800 574.000 472.400 ;
        RECT 575.600 471.800 578.000 472.400 ;
        RECT 580.400 472.000 581.200 479.800 ;
        RECT 583.600 475.200 584.400 479.800 ;
        RECT 558.000 471.200 558.600 471.800 ;
        RECT 558.000 470.600 561.400 471.200 ;
        RECT 560.600 470.400 561.400 470.600 ;
        RECT 562.200 470.400 562.800 471.800 ;
        RECT 569.200 471.200 569.800 471.800 ;
        RECT 569.200 470.600 572.600 471.200 ;
        RECT 571.800 470.400 572.600 470.600 ;
        RECT 573.400 470.400 574.000 471.800 ;
        RECT 580.200 471.200 581.200 472.000 ;
        RECT 581.800 474.600 584.400 475.200 ;
        RECT 581.800 473.000 582.400 474.600 ;
        RECT 586.800 474.400 587.600 479.800 ;
        RECT 590.000 477.000 590.800 479.800 ;
        RECT 591.600 477.000 592.400 479.800 ;
        RECT 593.200 477.000 594.000 479.800 ;
        RECT 588.200 474.400 592.400 475.200 ;
        RECT 585.000 473.600 587.600 474.400 ;
        RECT 594.800 473.600 595.600 479.800 ;
        RECT 598.000 475.000 598.800 479.800 ;
        RECT 601.200 475.000 602.000 479.800 ;
        RECT 602.800 477.000 603.600 479.800 ;
        RECT 604.400 477.000 605.200 479.800 ;
        RECT 607.600 475.200 608.400 479.800 ;
        RECT 610.800 476.400 611.600 479.800 ;
        RECT 610.800 475.800 611.800 476.400 ;
        RECT 611.200 475.200 611.800 475.800 ;
        RECT 606.400 474.400 610.600 475.200 ;
        RECT 611.200 474.600 613.200 475.200 ;
        RECT 598.000 473.600 600.600 474.400 ;
        RECT 601.200 473.800 607.000 474.400 ;
        RECT 610.000 474.000 610.600 474.400 ;
        RECT 590.000 473.000 590.800 473.200 ;
        RECT 581.800 472.400 590.800 473.000 ;
        RECT 593.200 473.000 594.000 473.200 ;
        RECT 601.200 473.000 601.800 473.800 ;
        RECT 607.600 473.200 609.000 473.800 ;
        RECT 610.000 473.200 611.600 474.000 ;
        RECT 593.200 472.400 601.800 473.000 ;
        RECT 602.800 473.000 609.000 473.200 ;
        RECT 602.800 472.600 608.200 473.000 ;
        RECT 602.800 472.400 603.600 472.600 ;
        RECT 558.400 469.800 559.200 470.000 ;
        RECT 562.200 469.800 563.600 470.400 ;
        RECT 573.400 470.300 574.800 470.400 ;
        RECT 578.800 470.300 579.600 470.400 ;
        RECT 558.400 469.200 561.000 469.800 ;
        RECT 560.400 468.600 561.000 469.200 ;
        RECT 561.800 469.600 563.600 469.800 ;
        RECT 569.600 469.800 570.400 470.000 ;
        RECT 573.400 469.800 579.600 470.300 ;
        RECT 561.800 469.200 562.800 469.600 ;
        RECT 569.600 469.200 572.200 469.800 ;
        RECT 556.400 468.200 558.000 468.400 ;
        RECT 556.400 467.600 559.800 468.200 ;
        RECT 560.400 467.800 561.200 468.600 ;
        RECT 559.200 467.200 559.800 467.600 ;
        RECT 557.800 466.800 558.600 467.000 ;
        RECT 551.600 465.700 554.000 466.300 ;
        RECT 551.600 464.800 552.400 465.700 ;
        RECT 550.000 462.200 550.800 464.200 ;
        RECT 553.200 462.200 554.000 465.700 ;
        RECT 554.800 464.800 555.600 466.400 ;
        RECT 556.400 466.200 558.600 466.800 ;
        RECT 559.200 466.600 561.200 467.200 ;
        RECT 559.600 466.400 561.200 466.600 ;
        RECT 556.400 462.200 557.200 466.200 ;
        RECT 561.800 465.800 562.400 469.200 ;
        RECT 571.600 468.600 572.200 469.200 ;
        RECT 573.000 469.700 579.600 469.800 ;
        RECT 573.000 469.600 574.800 469.700 ;
        RECT 578.800 469.600 579.600 469.700 ;
        RECT 573.000 469.200 574.000 469.600 ;
        RECT 563.200 467.600 564.000 468.400 ;
        RECT 565.200 467.600 566.800 468.400 ;
        RECT 567.600 468.200 569.200 468.400 ;
        RECT 567.600 467.600 571.000 468.200 ;
        RECT 571.600 467.800 572.400 468.600 ;
        RECT 563.200 467.200 563.800 467.600 ;
        RECT 563.000 466.400 563.800 467.200 ;
        RECT 570.400 467.200 571.000 467.600 ;
        RECT 564.400 466.800 565.200 467.000 ;
        RECT 569.000 466.800 569.800 467.000 ;
        RECT 564.400 466.200 566.800 466.800 ;
        RECT 560.800 464.400 562.400 465.800 ;
        RECT 560.800 463.600 563.600 464.400 ;
        RECT 560.800 462.200 562.400 463.600 ;
        RECT 566.000 462.200 566.800 466.200 ;
        RECT 567.600 466.200 569.800 466.800 ;
        RECT 570.400 466.600 572.400 467.200 ;
        RECT 570.800 466.400 572.400 466.600 ;
        RECT 567.600 462.200 568.400 466.200 ;
        RECT 573.000 465.800 573.600 469.200 ;
        RECT 574.400 467.600 575.200 468.400 ;
        RECT 576.400 468.300 578.000 468.400 ;
        RECT 580.200 468.300 581.000 471.200 ;
        RECT 581.800 470.600 582.400 472.400 ;
        RECT 576.400 467.700 581.000 468.300 ;
        RECT 576.400 467.600 578.000 467.700 ;
        RECT 574.400 467.200 575.000 467.600 ;
        RECT 574.200 466.400 575.000 467.200 ;
        RECT 575.600 466.800 576.400 467.000 ;
        RECT 580.200 466.800 581.000 467.700 ;
        RECT 581.600 470.000 582.400 470.600 ;
        RECT 588.400 470.000 611.800 470.600 ;
        RECT 581.600 468.000 582.200 470.000 ;
        RECT 588.400 469.400 589.200 470.000 ;
        RECT 606.000 469.600 606.800 470.000 ;
        RECT 611.000 469.800 611.800 470.000 ;
        RECT 582.800 468.600 586.600 469.400 ;
        RECT 581.600 467.400 582.800 468.000 ;
        RECT 575.600 466.200 578.000 466.800 ;
        RECT 572.000 462.200 573.600 465.800 ;
        RECT 577.200 462.200 578.000 466.200 ;
        RECT 580.200 466.000 581.200 466.800 ;
        RECT 580.400 462.200 581.200 466.000 ;
        RECT 582.000 462.200 582.800 467.400 ;
        RECT 585.800 467.400 586.600 468.600 ;
        RECT 585.800 466.800 587.600 467.400 ;
        RECT 586.800 466.200 587.600 466.800 ;
        RECT 591.600 466.400 592.400 469.200 ;
        RECT 594.800 468.600 598.000 469.400 ;
        RECT 601.800 468.600 603.800 469.400 ;
        RECT 612.400 469.000 613.200 474.600 ;
        RECT 594.400 467.800 595.200 468.000 ;
        RECT 594.400 467.200 598.800 467.800 ;
        RECT 598.000 467.000 598.800 467.200 ;
        RECT 599.600 466.800 600.400 468.400 ;
        RECT 586.800 465.400 589.200 466.200 ;
        RECT 591.600 465.600 592.600 466.400 ;
        RECT 595.600 465.600 597.200 466.400 ;
        RECT 598.000 466.200 598.800 466.400 ;
        RECT 601.800 466.200 602.600 468.600 ;
        RECT 604.400 468.200 613.200 469.000 ;
        RECT 607.800 466.800 610.800 467.600 ;
        RECT 607.800 466.200 608.600 466.800 ;
        RECT 598.000 465.600 602.600 466.200 ;
        RECT 588.400 462.200 589.200 465.400 ;
        RECT 606.000 465.400 608.600 466.200 ;
        RECT 590.000 462.200 590.800 465.000 ;
        RECT 591.600 462.200 592.400 465.000 ;
        RECT 593.200 462.200 594.000 465.000 ;
        RECT 594.800 462.200 595.600 465.000 ;
        RECT 598.000 462.200 598.800 465.000 ;
        RECT 601.200 462.200 602.000 465.000 ;
        RECT 602.800 462.200 603.600 465.000 ;
        RECT 604.400 462.200 605.200 465.000 ;
        RECT 606.000 462.200 606.800 465.400 ;
        RECT 612.400 462.200 613.200 468.200 ;
        RECT 1.200 455.400 2.000 459.800 ;
        RECT 5.400 458.400 6.600 459.800 ;
        RECT 5.400 457.800 6.800 458.400 ;
        RECT 10.000 457.800 10.800 459.800 ;
        RECT 14.400 458.400 15.200 459.800 ;
        RECT 14.400 457.800 16.400 458.400 ;
        RECT 6.000 457.000 6.800 457.800 ;
        RECT 10.200 457.200 10.800 457.800 ;
        RECT 10.200 456.600 13.000 457.200 ;
        RECT 12.200 456.400 13.000 456.600 ;
        RECT 14.000 456.400 14.800 457.200 ;
        RECT 15.600 457.000 16.400 457.800 ;
        RECT 4.200 455.400 5.000 455.600 ;
        RECT 1.200 454.800 5.000 455.400 ;
        RECT 1.200 451.400 2.000 454.800 ;
        RECT 8.200 454.200 9.000 454.400 ;
        RECT 14.000 454.200 14.600 456.400 ;
        RECT 18.800 455.000 19.600 459.800 ;
        RECT 20.400 456.000 21.200 459.800 ;
        RECT 23.600 456.000 24.400 459.800 ;
        RECT 20.400 455.800 24.400 456.000 ;
        RECT 25.200 455.800 26.000 459.800 ;
        RECT 30.600 456.000 31.400 459.000 ;
        RECT 34.800 457.000 35.600 459.000 ;
        RECT 20.600 455.400 24.200 455.800 ;
        RECT 21.200 454.400 22.000 454.800 ;
        RECT 25.200 454.400 25.800 455.800 ;
        RECT 29.800 455.400 31.400 456.000 ;
        RECT 29.800 455.000 30.600 455.400 ;
        RECT 29.800 454.400 30.400 455.000 ;
        RECT 35.000 454.800 35.600 457.000 ;
        RECT 36.400 455.600 37.200 457.200 ;
        RECT 17.200 454.200 18.800 454.400 ;
        RECT 7.800 453.600 18.800 454.200 ;
        RECT 20.400 453.800 22.000 454.400 ;
        RECT 20.400 453.600 21.200 453.800 ;
        RECT 23.400 453.600 26.000 454.400 ;
        RECT 26.800 454.300 27.600 454.400 ;
        RECT 28.400 454.300 30.400 454.400 ;
        RECT 26.800 453.700 30.400 454.300 ;
        RECT 31.400 454.200 35.600 454.800 ;
        RECT 31.400 453.800 32.400 454.200 ;
        RECT 26.800 453.600 27.600 453.700 ;
        RECT 28.400 453.600 30.400 453.700 ;
        RECT 6.000 452.800 6.800 453.000 ;
        RECT 3.000 452.200 6.800 452.800 ;
        RECT 3.000 452.000 3.800 452.200 ;
        RECT 4.600 451.400 5.400 451.600 ;
        RECT 1.200 450.800 5.400 451.400 ;
        RECT 1.200 442.200 2.000 450.800 ;
        RECT 7.800 450.400 8.400 453.600 ;
        RECT 15.000 453.400 15.800 453.600 ;
        RECT 14.000 452.400 14.800 452.600 ;
        RECT 16.600 452.400 17.400 452.600 ;
        RECT 12.400 451.800 17.400 452.400 ;
        RECT 12.400 451.600 13.200 451.800 ;
        RECT 22.000 451.600 22.800 453.200 ;
        RECT 23.400 452.400 24.000 453.600 ;
        RECT 23.400 451.600 24.400 452.400 ;
        RECT 14.000 451.000 19.600 451.200 ;
        RECT 13.800 450.800 19.600 451.000 ;
        RECT 6.000 449.800 8.400 450.400 ;
        RECT 9.800 450.600 19.600 450.800 ;
        RECT 9.800 450.200 14.600 450.600 ;
        RECT 6.000 448.800 6.600 449.800 ;
        RECT 5.200 448.000 6.600 448.800 ;
        RECT 8.200 449.000 9.000 449.200 ;
        RECT 9.800 449.000 10.400 450.200 ;
        RECT 8.200 448.400 10.400 449.000 ;
        RECT 11.000 449.000 16.400 449.600 ;
        RECT 11.000 448.800 11.800 449.000 ;
        RECT 15.600 448.800 16.400 449.000 ;
        RECT 9.400 447.400 10.200 447.600 ;
        RECT 12.200 447.400 13.000 447.600 ;
        RECT 6.000 446.200 6.800 447.000 ;
        RECT 9.400 446.800 13.000 447.400 ;
        RECT 10.200 446.200 10.800 446.800 ;
        RECT 15.600 446.200 16.400 447.000 ;
        RECT 5.400 442.200 6.600 446.200 ;
        RECT 10.000 442.200 10.800 446.200 ;
        RECT 14.400 445.600 16.400 446.200 ;
        RECT 14.400 442.200 15.200 445.600 ;
        RECT 18.800 442.200 19.600 450.600 ;
        RECT 23.400 450.200 24.000 451.600 ;
        RECT 28.400 450.800 29.200 452.400 ;
        RECT 25.200 450.200 26.000 450.400 ;
        RECT 23.000 449.600 24.000 450.200 ;
        RECT 24.600 449.600 26.000 450.200 ;
        RECT 29.800 449.800 30.400 453.600 ;
        RECT 31.000 453.000 32.400 453.800 ;
        RECT 31.800 451.000 32.400 453.000 ;
        RECT 33.200 451.600 34.000 453.200 ;
        RECT 34.800 451.600 35.600 453.200 ;
        RECT 31.800 450.400 35.600 451.000 ;
        RECT 23.000 442.200 23.800 449.600 ;
        RECT 24.600 448.400 25.200 449.600 ;
        RECT 29.800 449.200 31.400 449.800 ;
        RECT 24.400 447.600 25.200 448.400 ;
        RECT 30.600 442.200 31.400 449.200 ;
        RECT 35.000 447.000 35.600 450.400 ;
        RECT 34.800 443.000 35.600 447.000 ;
        RECT 38.000 442.200 38.800 459.800 ;
        RECT 41.200 456.400 42.000 459.800 ;
        RECT 41.000 455.800 42.000 456.400 ;
        RECT 41.000 454.400 41.600 455.800 ;
        RECT 44.400 455.200 45.200 459.800 ;
        RECT 46.000 455.800 46.800 459.800 ;
        RECT 47.600 456.000 48.400 459.800 ;
        RECT 50.800 456.000 51.600 459.800 ;
        RECT 47.600 455.800 51.600 456.000 ;
        RECT 42.600 454.600 45.200 455.200 ;
        RECT 41.000 453.600 42.000 454.400 ;
        RECT 41.000 450.200 41.600 453.600 ;
        RECT 42.600 453.000 43.200 454.600 ;
        RECT 46.200 454.400 46.800 455.800 ;
        RECT 47.800 455.400 51.400 455.800 ;
        RECT 52.400 455.000 53.200 459.800 ;
        RECT 56.800 458.400 57.600 459.800 ;
        RECT 55.600 457.800 57.600 458.400 ;
        RECT 61.200 457.800 62.000 459.800 ;
        RECT 65.400 458.400 66.600 459.800 ;
        RECT 65.200 457.800 66.600 458.400 ;
        RECT 55.600 457.000 56.400 457.800 ;
        RECT 61.200 457.200 61.800 457.800 ;
        RECT 57.200 456.400 58.000 457.200 ;
        RECT 59.000 456.600 61.800 457.200 ;
        RECT 65.200 457.000 66.000 457.800 ;
        RECT 59.000 456.400 59.800 456.600 ;
        RECT 50.000 454.400 50.800 454.800 ;
        RECT 46.000 453.600 48.600 454.400 ;
        RECT 50.000 453.800 51.600 454.400 ;
        RECT 50.800 453.600 51.600 453.800 ;
        RECT 53.200 454.200 54.800 454.400 ;
        RECT 57.400 454.200 58.000 456.400 ;
        RECT 67.000 455.400 67.800 455.600 ;
        RECT 70.000 455.400 70.800 459.800 ;
        RECT 67.000 454.800 70.800 455.400 ;
        RECT 63.000 454.200 63.800 454.400 ;
        RECT 53.200 453.600 64.200 454.200 ;
        RECT 42.200 452.200 43.200 453.000 ;
        RECT 42.600 450.200 43.200 452.200 ;
        RECT 44.200 452.400 45.000 453.200 ;
        RECT 44.200 451.600 45.200 452.400 ;
        RECT 46.000 450.200 46.800 450.400 ;
        RECT 48.000 450.200 48.600 453.600 ;
        RECT 56.200 453.400 57.000 453.600 ;
        RECT 49.200 451.600 50.000 453.200 ;
        RECT 54.600 452.400 55.400 452.600 ;
        RECT 54.600 451.800 59.600 452.400 ;
        RECT 58.800 451.600 59.600 451.800 ;
        RECT 52.400 451.000 58.000 451.200 ;
        RECT 52.400 450.800 58.200 451.000 ;
        RECT 52.400 450.600 62.200 450.800 ;
        RECT 41.000 449.200 42.000 450.200 ;
        RECT 42.600 449.600 45.200 450.200 ;
        RECT 46.000 449.600 47.400 450.200 ;
        RECT 48.000 449.600 49.000 450.200 ;
        RECT 41.200 442.200 42.000 449.200 ;
        RECT 44.400 442.200 45.200 449.600 ;
        RECT 46.800 448.400 47.400 449.600 ;
        RECT 46.800 447.600 47.600 448.400 ;
        RECT 48.200 442.200 49.000 449.600 ;
        RECT 52.400 442.200 53.200 450.600 ;
        RECT 57.400 450.200 62.200 450.600 ;
        RECT 55.600 449.000 61.000 449.600 ;
        RECT 55.600 448.800 56.400 449.000 ;
        RECT 60.200 448.800 61.000 449.000 ;
        RECT 61.600 449.000 62.200 450.200 ;
        RECT 63.600 450.400 64.200 453.600 ;
        RECT 65.200 452.800 66.000 453.000 ;
        RECT 65.200 452.200 69.000 452.800 ;
        RECT 68.200 452.000 69.000 452.200 ;
        RECT 66.600 451.400 67.400 451.600 ;
        RECT 70.000 451.400 70.800 454.800 ;
        RECT 71.600 457.000 72.400 459.000 ;
        RECT 71.600 454.800 72.200 457.000 ;
        RECT 75.800 456.000 76.600 459.000 ;
        RECT 81.200 456.000 82.000 459.800 ;
        RECT 84.400 456.000 85.200 459.800 ;
        RECT 75.800 455.400 77.400 456.000 ;
        RECT 81.200 455.800 85.200 456.000 ;
        RECT 86.000 455.800 86.800 459.800 ;
        RECT 87.600 455.800 88.400 459.800 ;
        RECT 89.200 456.000 90.000 459.800 ;
        RECT 92.400 456.000 93.200 459.800 ;
        RECT 95.600 456.400 96.400 459.800 ;
        RECT 89.200 455.800 93.200 456.000 ;
        RECT 95.400 455.800 96.400 456.400 ;
        RECT 81.400 455.400 85.000 455.800 ;
        RECT 76.600 455.000 77.400 455.400 ;
        RECT 71.600 454.200 75.800 454.800 ;
        RECT 74.800 453.800 75.800 454.200 ;
        RECT 76.800 454.400 77.400 455.000 ;
        RECT 82.000 454.400 82.800 454.800 ;
        RECT 86.000 454.400 86.600 455.800 ;
        RECT 87.800 454.400 88.400 455.800 ;
        RECT 89.400 455.400 93.000 455.800 ;
        RECT 91.600 454.400 92.400 454.800 ;
        RECT 95.400 454.400 96.000 455.800 ;
        RECT 98.800 455.200 99.600 459.800 ;
        RECT 100.400 456.000 101.200 459.800 ;
        RECT 103.600 456.000 104.400 459.800 ;
        RECT 100.400 455.800 104.400 456.000 ;
        RECT 100.600 455.400 104.200 455.800 ;
        RECT 105.200 455.600 106.000 459.800 ;
        RECT 97.000 454.600 99.600 455.200 ;
        RECT 76.800 454.300 78.800 454.400 ;
        RECT 79.600 454.300 80.400 454.400 ;
        RECT 71.600 451.600 72.400 453.200 ;
        RECT 73.200 451.600 74.000 453.200 ;
        RECT 74.800 453.000 76.200 453.800 ;
        RECT 76.800 453.700 80.400 454.300 ;
        RECT 76.800 453.600 78.800 453.700 ;
        RECT 79.600 453.600 80.400 453.700 ;
        RECT 81.200 453.800 82.800 454.400 ;
        RECT 81.200 453.600 82.000 453.800 ;
        RECT 84.200 453.600 86.800 454.400 ;
        RECT 87.600 453.600 90.200 454.400 ;
        RECT 91.600 454.300 93.200 454.400 ;
        RECT 95.400 454.300 96.400 454.400 ;
        RECT 91.600 453.800 96.400 454.300 ;
        RECT 92.400 453.700 96.400 453.800 ;
        RECT 92.400 453.600 93.200 453.700 ;
        RECT 95.400 453.600 96.400 453.700 ;
        RECT 66.600 450.800 70.800 451.400 ;
        RECT 74.800 451.000 75.400 453.000 ;
        RECT 63.600 449.800 66.000 450.400 ;
        RECT 63.000 449.000 63.800 449.200 ;
        RECT 61.600 448.400 63.800 449.000 ;
        RECT 65.400 448.800 66.000 449.800 ;
        RECT 65.400 448.000 66.800 448.800 ;
        RECT 59.000 447.400 59.800 447.600 ;
        RECT 61.800 447.400 62.600 447.600 ;
        RECT 55.600 446.200 56.400 447.000 ;
        RECT 59.000 446.800 62.600 447.400 ;
        RECT 61.200 446.200 61.800 446.800 ;
        RECT 65.200 446.200 66.000 447.000 ;
        RECT 55.600 445.600 57.600 446.200 ;
        RECT 56.800 442.200 57.600 445.600 ;
        RECT 61.200 442.200 62.000 446.200 ;
        RECT 65.400 442.200 66.600 446.200 ;
        RECT 70.000 442.200 70.800 450.800 ;
        RECT 71.600 450.400 75.400 451.000 ;
        RECT 71.600 447.000 72.200 450.400 ;
        RECT 76.800 449.800 77.400 453.600 ;
        RECT 78.000 452.300 78.800 452.400 ;
        RECT 79.600 452.300 80.400 452.400 ;
        RECT 78.000 451.700 80.400 452.300 ;
        RECT 78.000 450.800 78.800 451.700 ;
        RECT 79.600 451.600 80.400 451.700 ;
        RECT 82.800 451.600 83.600 453.200 ;
        RECT 84.200 450.400 84.800 453.600 ;
        RECT 89.600 452.300 90.200 453.600 ;
        RECT 86.100 451.700 90.200 452.300 ;
        RECT 86.100 450.400 86.700 451.700 ;
        RECT 75.800 449.200 77.400 449.800 ;
        RECT 82.800 449.600 84.800 450.400 ;
        RECT 86.000 450.200 86.800 450.400 ;
        RECT 85.400 449.600 86.800 450.200 ;
        RECT 87.600 450.200 88.400 450.400 ;
        RECT 89.600 450.200 90.200 451.700 ;
        RECT 90.800 451.600 91.600 453.200 ;
        RECT 95.400 450.200 96.000 453.600 ;
        RECT 97.000 453.000 97.600 454.600 ;
        RECT 101.200 454.400 102.000 454.800 ;
        RECT 105.200 454.400 105.800 455.600 ;
        RECT 100.400 453.800 102.000 454.400 ;
        RECT 100.400 453.600 101.200 453.800 ;
        RECT 103.400 453.600 106.000 454.400 ;
        RECT 110.400 454.200 111.200 459.800 ;
        RECT 116.800 454.200 117.600 459.800 ;
        RECT 123.400 456.000 124.200 459.000 ;
        RECT 127.600 457.000 128.400 459.000 ;
        RECT 122.600 455.400 124.200 456.000 ;
        RECT 122.600 455.000 123.400 455.400 ;
        RECT 122.600 454.400 123.200 455.000 ;
        RECT 127.800 454.800 128.400 457.000 ;
        RECT 129.200 455.600 130.000 457.200 ;
        RECT 110.400 453.800 112.200 454.200 ;
        RECT 116.800 453.800 118.600 454.200 ;
        RECT 110.600 453.600 112.200 453.800 ;
        RECT 117.000 453.600 118.600 453.800 ;
        RECT 121.200 453.600 123.200 454.400 ;
        RECT 124.200 454.200 128.400 454.800 ;
        RECT 124.200 453.800 125.200 454.200 ;
        RECT 96.600 452.200 97.600 453.000 ;
        RECT 97.000 450.200 97.600 452.200 ;
        RECT 98.600 452.400 99.400 453.200 ;
        RECT 98.600 451.600 99.600 452.400 ;
        RECT 100.400 452.300 101.200 452.400 ;
        RECT 102.000 452.300 102.800 453.200 ;
        RECT 100.400 451.700 102.800 452.300 ;
        RECT 100.400 451.600 101.200 451.700 ;
        RECT 102.000 451.600 102.800 451.700 ;
        RECT 103.400 450.200 104.000 453.600 ;
        RECT 108.400 451.600 110.000 452.400 ;
        RECT 105.200 450.200 106.000 450.400 ;
        RECT 87.600 449.600 89.000 450.200 ;
        RECT 89.600 449.600 90.600 450.200 ;
        RECT 71.600 443.000 72.400 447.000 ;
        RECT 75.800 442.200 76.600 449.200 ;
        RECT 83.800 442.200 84.600 449.600 ;
        RECT 85.400 448.400 86.000 449.600 ;
        RECT 85.200 447.600 86.000 448.400 ;
        RECT 88.400 448.400 89.000 449.600 ;
        RECT 88.400 447.600 89.200 448.400 ;
        RECT 89.800 442.200 90.600 449.600 ;
        RECT 95.400 449.200 96.400 450.200 ;
        RECT 97.000 449.600 99.600 450.200 ;
        RECT 95.600 442.200 96.400 449.200 ;
        RECT 98.800 442.200 99.600 449.600 ;
        RECT 103.000 449.600 104.000 450.200 ;
        RECT 104.600 449.600 106.000 450.200 ;
        RECT 106.800 449.600 107.600 451.200 ;
        RECT 111.600 450.400 112.200 453.600 ;
        RECT 114.800 451.600 116.400 452.400 ;
        RECT 111.600 449.600 112.400 450.400 ;
        RECT 113.200 449.600 114.000 451.200 ;
        RECT 118.000 450.400 118.600 453.600 ;
        RECT 121.200 450.800 122.000 452.400 ;
        RECT 118.000 449.600 118.800 450.400 ;
        RECT 122.600 449.800 123.200 453.600 ;
        RECT 123.800 453.000 125.200 453.800 ;
        RECT 124.600 451.000 125.200 453.000 ;
        RECT 126.000 451.600 126.800 453.200 ;
        RECT 127.600 451.600 128.400 453.200 ;
        RECT 124.600 450.400 128.400 451.000 ;
        RECT 103.000 442.200 103.800 449.600 ;
        RECT 104.600 448.400 105.200 449.600 ;
        RECT 104.400 447.600 105.200 448.400 ;
        RECT 110.000 447.600 110.800 449.200 ;
        RECT 111.600 448.300 112.200 449.600 ;
        RECT 114.800 448.300 115.600 448.400 ;
        RECT 111.600 447.700 115.600 448.300 ;
        RECT 111.600 447.000 112.200 447.700 ;
        RECT 114.800 447.600 115.600 447.700 ;
        RECT 116.400 447.600 117.200 449.200 ;
        RECT 118.000 447.000 118.600 449.600 ;
        RECT 122.600 449.200 124.200 449.800 ;
        RECT 108.600 446.400 112.200 447.000 ;
        RECT 108.600 446.200 109.200 446.400 ;
        RECT 108.400 442.200 109.200 446.200 ;
        RECT 111.600 446.200 112.200 446.400 ;
        RECT 115.000 446.400 118.600 447.000 ;
        RECT 115.000 446.200 115.600 446.400 ;
        RECT 111.600 442.200 112.400 446.200 ;
        RECT 114.800 442.200 115.600 446.200 ;
        RECT 118.000 446.200 118.600 446.400 ;
        RECT 118.000 442.200 118.800 446.200 ;
        RECT 123.400 444.400 124.200 449.200 ;
        RECT 127.800 447.000 128.400 450.400 ;
        RECT 122.800 443.600 124.200 444.400 ;
        RECT 123.400 442.200 124.200 443.600 ;
        RECT 127.600 443.000 128.400 447.000 ;
        RECT 130.800 442.200 131.600 459.800 ;
        RECT 132.400 456.000 133.200 459.800 ;
        RECT 135.600 456.000 136.400 459.800 ;
        RECT 132.400 455.800 136.400 456.000 ;
        RECT 137.200 455.800 138.000 459.800 ;
        RECT 138.800 456.000 139.600 459.800 ;
        RECT 142.000 456.000 142.800 459.800 ;
        RECT 138.800 455.800 142.800 456.000 ;
        RECT 143.600 455.800 144.400 459.800 ;
        RECT 147.800 458.300 148.600 459.800 ;
        RECT 150.000 458.300 150.800 458.400 ;
        RECT 147.800 457.700 150.800 458.300 ;
        RECT 147.800 456.400 148.600 457.700 ;
        RECT 150.000 457.600 150.800 457.700 ;
        RECT 146.800 455.800 148.600 456.400 ;
        RECT 158.600 456.000 159.400 459.000 ;
        RECT 162.800 457.000 163.600 459.000 ;
        RECT 132.600 455.400 136.200 455.800 ;
        RECT 133.200 454.400 134.000 454.800 ;
        RECT 137.200 454.400 137.800 455.800 ;
        RECT 139.000 455.400 142.600 455.800 ;
        RECT 139.600 454.400 140.400 454.800 ;
        RECT 143.600 454.400 144.200 455.800 ;
        RECT 132.400 453.800 134.000 454.400 ;
        RECT 135.400 454.300 138.000 454.400 ;
        RECT 138.800 454.300 140.400 454.400 ;
        RECT 135.400 453.800 140.400 454.300 ;
        RECT 132.400 453.600 133.200 453.800 ;
        RECT 135.400 453.700 139.600 453.800 ;
        RECT 135.400 453.600 138.000 453.700 ;
        RECT 138.800 453.600 139.600 453.700 ;
        RECT 141.800 453.600 144.400 454.400 ;
        RECT 145.200 453.600 146.000 455.200 ;
        RECT 134.000 451.600 134.800 453.200 ;
        RECT 135.400 450.200 136.000 453.600 ;
        RECT 138.800 452.300 139.600 452.400 ;
        RECT 137.300 451.700 139.600 452.300 ;
        RECT 137.300 450.400 137.900 451.700 ;
        RECT 138.800 451.600 139.600 451.700 ;
        RECT 140.400 451.600 141.200 453.200 ;
        RECT 137.200 450.200 138.000 450.400 ;
        RECT 141.800 450.200 142.400 453.600 ;
        RECT 143.600 450.200 144.400 450.400 ;
        RECT 135.000 449.600 136.000 450.200 ;
        RECT 136.600 449.600 138.000 450.200 ;
        RECT 141.400 449.600 142.400 450.200 ;
        RECT 143.000 449.600 144.400 450.200 ;
        RECT 135.000 442.200 135.800 449.600 ;
        RECT 136.600 448.400 137.200 449.600 ;
        RECT 136.400 447.600 137.200 448.400 ;
        RECT 141.400 444.400 142.200 449.600 ;
        RECT 143.000 448.400 143.600 449.600 ;
        RECT 142.800 447.600 143.600 448.400 ;
        RECT 140.400 443.600 142.200 444.400 ;
        RECT 141.400 442.200 142.200 443.600 ;
        RECT 146.800 442.200 147.600 455.800 ;
        RECT 157.800 455.400 159.400 456.000 ;
        RECT 157.800 455.000 158.600 455.400 ;
        RECT 157.800 454.400 158.400 455.000 ;
        RECT 163.000 454.800 163.600 457.000 ;
        RECT 156.400 453.600 158.400 454.400 ;
        RECT 159.400 454.200 163.600 454.800 ;
        RECT 165.600 454.200 166.400 459.800 ;
        RECT 170.800 456.000 171.600 459.800 ;
        RECT 174.000 456.000 174.800 459.800 ;
        RECT 170.800 455.800 174.800 456.000 ;
        RECT 175.600 455.800 176.400 459.800 ;
        RECT 171.000 455.400 174.600 455.800 ;
        RECT 171.600 454.400 172.400 454.800 ;
        RECT 175.600 454.400 176.200 455.800 ;
        RECT 177.200 455.400 178.000 459.800 ;
        RECT 181.400 458.400 182.600 459.800 ;
        RECT 181.400 457.800 182.800 458.400 ;
        RECT 186.000 457.800 186.800 459.800 ;
        RECT 190.400 458.400 191.200 459.800 ;
        RECT 190.400 457.800 192.400 458.400 ;
        RECT 182.000 457.000 182.800 457.800 ;
        RECT 186.200 457.200 186.800 457.800 ;
        RECT 186.200 456.600 189.000 457.200 ;
        RECT 188.200 456.400 189.000 456.600 ;
        RECT 190.000 456.400 190.800 457.200 ;
        RECT 191.600 457.000 192.400 457.800 ;
        RECT 180.200 455.400 181.000 455.600 ;
        RECT 177.200 454.800 181.000 455.400 ;
        RECT 159.400 453.800 160.400 454.200 ;
        RECT 156.400 450.800 157.200 452.400 ;
        RECT 148.400 448.800 149.200 450.400 ;
        RECT 157.800 449.800 158.400 453.600 ;
        RECT 159.000 453.000 160.400 453.800 ;
        RECT 164.600 453.800 166.400 454.200 ;
        RECT 170.800 453.800 172.400 454.400 ;
        RECT 164.600 453.600 166.200 453.800 ;
        RECT 170.800 453.600 171.600 453.800 ;
        RECT 173.800 453.600 176.400 454.400 ;
        RECT 159.800 451.000 160.400 453.000 ;
        RECT 161.200 451.600 162.000 453.200 ;
        RECT 162.800 451.600 163.600 453.200 ;
        RECT 159.800 450.400 163.600 451.000 ;
        RECT 164.600 450.400 165.200 453.600 ;
        RECT 166.800 451.600 168.400 452.400 ;
        RECT 172.400 451.600 173.200 453.200 ;
        RECT 157.800 449.200 159.400 449.800 ;
        RECT 158.600 444.400 159.400 449.200 ;
        RECT 163.000 447.000 163.600 450.400 ;
        RECT 164.400 449.600 165.200 450.400 ;
        RECT 169.200 449.600 170.000 451.200 ;
        RECT 173.800 450.200 174.400 453.600 ;
        RECT 177.200 451.400 178.000 454.800 ;
        RECT 184.200 454.200 185.000 454.400 ;
        RECT 190.000 454.200 190.600 456.400 ;
        RECT 194.800 455.000 195.600 459.800 ;
        RECT 193.200 454.200 194.800 454.400 ;
        RECT 183.800 453.600 194.800 454.200 ;
        RECT 200.000 454.200 200.800 459.800 ;
        RECT 202.800 455.600 203.600 457.200 ;
        RECT 200.000 453.800 201.800 454.200 ;
        RECT 200.200 453.600 201.800 453.800 ;
        RECT 182.000 452.800 182.800 453.000 ;
        RECT 179.000 452.200 182.800 452.800 ;
        RECT 179.000 452.000 179.800 452.200 ;
        RECT 180.600 451.400 181.400 451.600 ;
        RECT 177.200 450.800 181.400 451.400 ;
        RECT 175.600 450.200 176.400 450.400 ;
        RECT 173.400 449.600 174.400 450.200 ;
        RECT 175.000 449.600 176.400 450.200 ;
        RECT 158.000 443.600 159.400 444.400 ;
        RECT 158.600 442.200 159.400 443.600 ;
        RECT 162.800 443.000 163.600 447.000 ;
        RECT 164.600 447.000 165.200 449.600 ;
        RECT 166.000 447.600 166.800 449.200 ;
        RECT 164.600 446.400 168.200 447.000 ;
        RECT 164.600 446.200 165.200 446.400 ;
        RECT 164.400 442.200 165.200 446.200 ;
        RECT 167.600 446.200 168.200 446.400 ;
        RECT 167.600 442.200 168.400 446.200 ;
        RECT 173.400 442.200 174.200 449.600 ;
        RECT 175.000 448.400 175.600 449.600 ;
        RECT 174.800 447.600 175.600 448.400 ;
        RECT 177.200 442.200 178.000 450.800 ;
        RECT 183.800 450.400 184.400 453.600 ;
        RECT 191.000 453.400 191.800 453.600 ;
        RECT 192.600 452.400 193.400 452.600 ;
        RECT 188.400 451.800 193.400 452.400 ;
        RECT 188.400 451.600 189.200 451.800 ;
        RECT 198.000 451.600 199.600 452.400 ;
        RECT 190.000 451.000 195.600 451.200 ;
        RECT 189.800 450.800 195.600 451.000 ;
        RECT 182.000 449.800 184.400 450.400 ;
        RECT 185.800 450.600 195.600 450.800 ;
        RECT 185.800 450.200 190.600 450.600 ;
        RECT 182.000 448.800 182.600 449.800 ;
        RECT 181.200 448.000 182.600 448.800 ;
        RECT 184.200 449.000 185.000 449.200 ;
        RECT 185.800 449.000 186.400 450.200 ;
        RECT 184.200 448.400 186.400 449.000 ;
        RECT 187.000 449.000 192.400 449.600 ;
        RECT 187.000 448.800 187.800 449.000 ;
        RECT 191.600 448.800 192.400 449.000 ;
        RECT 185.400 447.400 186.200 447.600 ;
        RECT 188.200 447.400 189.000 447.600 ;
        RECT 182.000 446.200 182.800 447.000 ;
        RECT 185.400 446.800 189.000 447.400 ;
        RECT 186.200 446.200 186.800 446.800 ;
        RECT 191.600 446.200 192.400 447.000 ;
        RECT 181.400 442.200 182.600 446.200 ;
        RECT 186.000 442.200 186.800 446.200 ;
        RECT 190.400 445.600 192.400 446.200 ;
        RECT 190.400 442.200 191.200 445.600 ;
        RECT 194.800 442.200 195.600 450.600 ;
        RECT 196.400 449.600 197.200 451.200 ;
        RECT 201.200 450.400 201.800 453.600 ;
        RECT 201.200 449.600 202.000 450.400 ;
        RECT 204.400 450.300 205.200 459.800 ;
        RECT 206.600 458.400 207.400 459.800 ;
        RECT 206.600 457.600 208.400 458.400 ;
        RECT 206.600 456.400 207.400 457.600 ;
        RECT 206.600 455.800 208.400 456.400 ;
        RECT 206.000 450.300 206.800 450.400 ;
        RECT 204.400 449.700 206.800 450.300 ;
        RECT 199.600 447.600 200.400 449.200 ;
        RECT 201.200 447.000 201.800 449.600 ;
        RECT 198.200 446.400 201.800 447.000 ;
        RECT 198.200 446.200 198.800 446.400 ;
        RECT 198.000 442.200 198.800 446.200 ;
        RECT 201.200 446.200 201.800 446.400 ;
        RECT 201.200 442.200 202.000 446.200 ;
        RECT 204.400 442.200 205.200 449.700 ;
        RECT 206.000 448.800 206.800 449.700 ;
        RECT 207.600 442.200 208.400 455.800 ;
        RECT 212.400 455.200 213.200 459.800 ;
        RECT 215.600 455.200 216.400 459.800 ;
        RECT 218.800 455.200 219.600 459.800 ;
        RECT 222.000 455.200 222.800 459.800 ;
        RECT 225.800 458.400 226.600 459.800 ;
        RECT 225.200 457.600 226.600 458.400 ;
        RECT 225.800 456.400 226.600 457.600 ;
        RECT 225.800 455.800 227.600 456.400 ;
        RECT 209.200 453.600 210.000 455.200 ;
        RECT 212.400 454.400 214.200 455.200 ;
        RECT 215.600 454.400 217.800 455.200 ;
        RECT 218.800 454.400 221.000 455.200 ;
        RECT 222.000 454.400 224.400 455.200 ;
        RECT 210.800 453.800 211.600 454.400 ;
        RECT 213.400 453.800 214.200 454.400 ;
        RECT 217.000 453.800 217.800 454.400 ;
        RECT 220.200 453.800 221.000 454.400 ;
        RECT 210.800 453.000 212.600 453.800 ;
        RECT 213.400 453.000 216.000 453.800 ;
        RECT 217.000 453.000 219.400 453.800 ;
        RECT 220.200 453.000 222.800 453.800 ;
        RECT 213.400 451.600 214.200 453.000 ;
        RECT 217.000 451.600 217.800 453.000 ;
        RECT 220.200 451.600 221.000 453.000 ;
        RECT 223.600 451.600 224.400 454.400 ;
        RECT 212.400 450.800 214.200 451.600 ;
        RECT 215.600 450.800 217.800 451.600 ;
        RECT 218.800 450.800 221.000 451.600 ;
        RECT 222.000 450.800 224.400 451.600 ;
        RECT 212.400 442.200 213.200 450.800 ;
        RECT 215.600 442.200 216.400 450.800 ;
        RECT 218.800 442.200 219.600 450.800 ;
        RECT 222.000 442.200 222.800 450.800 ;
        RECT 225.200 448.800 226.000 450.400 ;
        RECT 226.800 442.200 227.600 455.800 ;
        RECT 230.000 455.200 230.800 459.800 ;
        RECT 233.200 456.400 234.000 459.800 ;
        RECT 233.200 455.800 234.200 456.400 ;
        RECT 238.000 456.000 238.800 459.800 ;
        RECT 228.400 453.600 229.200 455.200 ;
        RECT 230.000 454.600 232.600 455.200 ;
        RECT 230.200 452.400 231.000 453.200 ;
        RECT 230.000 451.600 231.000 452.400 ;
        RECT 232.000 453.000 232.600 454.600 ;
        RECT 233.600 454.400 234.200 455.800 ;
        RECT 233.200 453.600 234.200 454.400 ;
        RECT 232.000 452.200 233.000 453.000 ;
        RECT 232.000 450.200 232.600 452.200 ;
        RECT 233.600 450.200 234.200 453.600 ;
        RECT 230.000 449.600 232.600 450.200 ;
        RECT 230.000 442.200 230.800 449.600 ;
        RECT 233.200 449.200 234.200 450.200 ;
        RECT 237.800 455.200 238.800 456.000 ;
        RECT 237.800 450.800 238.600 455.200 ;
        RECT 239.600 454.600 240.400 459.800 ;
        RECT 246.000 456.600 246.800 459.800 ;
        RECT 247.600 457.000 248.400 459.800 ;
        RECT 249.200 457.000 250.000 459.800 ;
        RECT 250.800 457.000 251.600 459.800 ;
        RECT 252.400 457.000 253.200 459.800 ;
        RECT 255.600 457.000 256.400 459.800 ;
        RECT 258.800 457.000 259.600 459.800 ;
        RECT 260.400 457.000 261.200 459.800 ;
        RECT 262.000 457.000 262.800 459.800 ;
        RECT 244.400 455.800 246.800 456.600 ;
        RECT 263.600 456.600 264.400 459.800 ;
        RECT 244.400 455.200 245.200 455.800 ;
        RECT 239.200 454.000 240.400 454.600 ;
        RECT 243.400 454.600 245.200 455.200 ;
        RECT 249.200 455.600 250.200 456.400 ;
        RECT 253.200 455.600 254.800 456.400 ;
        RECT 255.600 455.800 260.200 456.400 ;
        RECT 263.600 455.800 266.200 456.600 ;
        RECT 255.600 455.600 256.400 455.800 ;
        RECT 239.200 452.000 239.800 454.000 ;
        RECT 243.400 453.400 244.200 454.600 ;
        RECT 240.400 452.600 244.200 453.400 ;
        RECT 249.200 452.800 250.000 455.600 ;
        RECT 255.600 454.800 256.400 455.000 ;
        RECT 252.000 454.200 256.400 454.800 ;
        RECT 252.000 454.000 252.800 454.200 ;
        RECT 257.200 453.600 258.000 455.200 ;
        RECT 259.400 453.400 260.200 455.800 ;
        RECT 265.400 455.200 266.200 455.800 ;
        RECT 265.400 454.400 268.400 455.200 ;
        RECT 270.000 453.800 270.800 459.800 ;
        RECT 252.400 452.600 255.600 453.400 ;
        RECT 259.400 452.600 261.400 453.400 ;
        RECT 262.000 453.000 270.800 453.800 ;
        RECT 246.000 452.000 246.800 452.600 ;
        RECT 263.600 452.000 264.400 452.400 ;
        RECT 268.600 452.000 269.400 452.200 ;
        RECT 239.200 451.400 240.000 452.000 ;
        RECT 246.000 451.400 269.400 452.000 ;
        RECT 237.800 450.000 238.800 450.800 ;
        RECT 233.200 442.200 234.000 449.200 ;
        RECT 238.000 442.200 238.800 450.000 ;
        RECT 239.400 449.600 240.000 451.400 ;
        RECT 239.400 449.000 248.400 449.600 ;
        RECT 239.400 447.400 240.000 449.000 ;
        RECT 247.600 448.800 248.400 449.000 ;
        RECT 250.800 449.000 259.400 449.600 ;
        RECT 250.800 448.800 251.600 449.000 ;
        RECT 242.600 447.600 245.200 448.400 ;
        RECT 239.400 446.800 242.000 447.400 ;
        RECT 241.200 442.200 242.000 446.800 ;
        RECT 244.400 442.200 245.200 447.600 ;
        RECT 245.800 446.800 250.000 447.600 ;
        RECT 247.600 442.200 248.400 445.000 ;
        RECT 249.200 442.200 250.000 445.000 ;
        RECT 250.800 442.200 251.600 445.000 ;
        RECT 252.400 442.200 253.200 448.400 ;
        RECT 255.600 447.600 258.200 448.400 ;
        RECT 258.800 448.200 259.400 449.000 ;
        RECT 260.400 449.400 261.200 449.600 ;
        RECT 260.400 449.000 265.800 449.400 ;
        RECT 260.400 448.800 266.600 449.000 ;
        RECT 265.200 448.200 266.600 448.800 ;
        RECT 258.800 447.600 264.600 448.200 ;
        RECT 267.600 448.000 269.200 448.800 ;
        RECT 267.600 447.600 268.200 448.000 ;
        RECT 255.600 442.200 256.400 447.000 ;
        RECT 258.800 442.200 259.600 447.000 ;
        RECT 264.000 446.800 268.200 447.600 ;
        RECT 270.000 447.400 270.800 453.000 ;
        RECT 271.600 455.800 272.400 459.800 ;
        RECT 274.800 457.800 275.600 459.800 ;
        RECT 271.600 452.400 272.200 455.800 ;
        RECT 274.800 455.600 275.400 457.800 ;
        RECT 276.400 455.600 277.200 457.200 ;
        RECT 273.000 455.000 275.400 455.600 ;
        RECT 278.000 455.200 278.800 459.800 ;
        RECT 281.200 456.400 282.000 459.800 ;
        RECT 281.200 455.600 282.200 456.400 ;
        RECT 284.400 456.000 285.200 459.800 ;
        RECT 287.600 456.000 288.400 459.800 ;
        RECT 284.400 455.800 288.400 456.000 ;
        RECT 289.200 455.800 290.000 459.800 ;
        RECT 297.200 456.000 298.000 459.800 ;
        RECT 271.600 451.600 272.400 452.400 ;
        RECT 273.000 452.000 273.600 455.000 ;
        RECT 278.000 454.600 280.600 455.200 ;
        RECT 274.600 453.600 275.600 454.400 ;
        RECT 274.400 452.800 275.200 453.600 ;
        RECT 278.200 452.400 279.000 453.200 ;
        RECT 271.600 450.200 272.200 451.600 ;
        RECT 273.000 451.400 273.800 452.000 ;
        RECT 278.000 451.600 279.000 452.400 ;
        RECT 280.000 453.000 280.600 454.600 ;
        RECT 281.600 454.400 282.200 455.600 ;
        RECT 284.600 455.400 288.200 455.800 ;
        RECT 285.200 454.400 286.000 454.800 ;
        RECT 289.200 454.400 289.800 455.800 ;
        RECT 297.000 455.200 298.000 456.000 ;
        RECT 281.200 454.300 282.200 454.400 ;
        RECT 284.400 454.300 286.000 454.400 ;
        RECT 281.200 453.800 286.000 454.300 ;
        RECT 281.200 453.700 285.200 453.800 ;
        RECT 281.200 453.600 282.200 453.700 ;
        RECT 284.400 453.600 285.200 453.700 ;
        RECT 287.400 453.600 290.000 454.400 ;
        RECT 280.000 452.200 281.000 453.000 ;
        RECT 273.000 451.200 277.200 451.400 ;
        RECT 273.200 450.800 277.200 451.200 ;
        RECT 271.600 449.600 273.000 450.200 ;
        RECT 268.800 446.800 270.800 447.400 ;
        RECT 260.400 442.200 261.200 445.000 ;
        RECT 262.000 442.200 262.800 445.000 ;
        RECT 265.200 442.200 266.000 446.800 ;
        RECT 268.800 446.200 269.400 446.800 ;
        RECT 268.400 445.600 269.400 446.200 ;
        RECT 268.400 442.200 269.200 445.600 ;
        RECT 272.200 444.400 273.000 449.600 ;
        RECT 271.600 443.600 273.000 444.400 ;
        RECT 272.200 442.200 273.000 443.600 ;
        RECT 276.400 442.200 277.200 450.800 ;
        RECT 280.000 450.200 280.600 452.200 ;
        RECT 281.600 450.200 282.200 453.600 ;
        RECT 286.000 451.600 286.800 453.200 ;
        RECT 287.400 450.200 288.000 453.600 ;
        RECT 297.000 450.800 297.800 455.200 ;
        RECT 298.800 454.600 299.600 459.800 ;
        RECT 305.200 456.600 306.000 459.800 ;
        RECT 306.800 457.000 307.600 459.800 ;
        RECT 308.400 457.000 309.200 459.800 ;
        RECT 310.000 457.000 310.800 459.800 ;
        RECT 311.600 457.000 312.400 459.800 ;
        RECT 314.800 457.000 315.600 459.800 ;
        RECT 318.000 457.000 318.800 459.800 ;
        RECT 319.600 457.000 320.400 459.800 ;
        RECT 321.200 457.000 322.000 459.800 ;
        RECT 303.600 455.800 306.000 456.600 ;
        RECT 322.800 456.600 323.600 459.800 ;
        RECT 303.600 455.200 304.400 455.800 ;
        RECT 298.400 454.000 299.600 454.600 ;
        RECT 302.600 454.600 304.400 455.200 ;
        RECT 308.400 455.600 309.400 456.400 ;
        RECT 312.400 455.600 314.000 456.400 ;
        RECT 314.800 455.800 319.400 456.400 ;
        RECT 322.800 455.800 325.400 456.600 ;
        RECT 314.800 455.600 315.600 455.800 ;
        RECT 298.400 452.000 299.000 454.000 ;
        RECT 302.600 453.400 303.400 454.600 ;
        RECT 299.600 452.600 303.400 453.400 ;
        RECT 308.400 452.800 309.200 455.600 ;
        RECT 314.800 454.800 315.600 455.000 ;
        RECT 311.200 454.200 315.600 454.800 ;
        RECT 311.200 454.000 312.000 454.200 ;
        RECT 316.400 453.600 317.200 455.200 ;
        RECT 318.600 453.400 319.400 455.800 ;
        RECT 324.600 455.200 325.400 455.800 ;
        RECT 324.600 454.400 327.600 455.200 ;
        RECT 329.200 453.800 330.000 459.800 ;
        RECT 311.600 452.600 314.800 453.400 ;
        RECT 318.600 452.600 320.600 453.400 ;
        RECT 321.200 453.000 330.000 453.800 ;
        RECT 305.200 452.000 306.000 452.600 ;
        RECT 322.800 452.000 323.600 452.400 ;
        RECT 327.800 452.000 328.600 452.200 ;
        RECT 298.400 451.400 299.200 452.000 ;
        RECT 305.200 451.400 328.600 452.000 ;
        RECT 289.200 450.300 290.000 450.400 ;
        RECT 297.000 450.300 298.000 450.800 ;
        RECT 289.200 450.200 298.000 450.300 ;
        RECT 278.000 449.600 280.600 450.200 ;
        RECT 278.000 442.200 278.800 449.600 ;
        RECT 281.200 449.200 282.200 450.200 ;
        RECT 287.000 449.600 288.000 450.200 ;
        RECT 288.600 449.700 298.000 450.200 ;
        RECT 288.600 449.600 290.000 449.700 ;
        RECT 281.200 442.200 282.000 449.200 ;
        RECT 287.000 442.200 287.800 449.600 ;
        RECT 288.600 448.400 289.200 449.600 ;
        RECT 288.400 447.600 289.200 448.400 ;
        RECT 297.200 442.200 298.000 449.700 ;
        RECT 298.600 449.600 299.200 451.400 ;
        RECT 298.600 449.000 307.600 449.600 ;
        RECT 298.600 447.400 299.200 449.000 ;
        RECT 306.800 448.800 307.600 449.000 ;
        RECT 310.000 449.000 318.600 449.600 ;
        RECT 310.000 448.800 310.800 449.000 ;
        RECT 301.800 447.600 304.400 448.400 ;
        RECT 298.600 446.800 301.200 447.400 ;
        RECT 300.400 442.200 301.200 446.800 ;
        RECT 303.600 442.200 304.400 447.600 ;
        RECT 305.000 446.800 309.200 447.600 ;
        RECT 306.800 442.200 307.600 445.000 ;
        RECT 308.400 442.200 309.200 445.000 ;
        RECT 310.000 442.200 310.800 445.000 ;
        RECT 311.600 442.200 312.400 448.400 ;
        RECT 314.800 447.600 317.400 448.400 ;
        RECT 318.000 448.200 318.600 449.000 ;
        RECT 319.600 449.400 320.400 449.600 ;
        RECT 319.600 449.000 325.000 449.400 ;
        RECT 319.600 448.800 325.800 449.000 ;
        RECT 324.400 448.200 325.800 448.800 ;
        RECT 318.000 447.600 323.800 448.200 ;
        RECT 326.800 448.000 328.400 448.800 ;
        RECT 326.800 447.600 327.400 448.000 ;
        RECT 314.800 442.200 315.600 447.000 ;
        RECT 318.000 442.200 318.800 447.000 ;
        RECT 323.200 446.800 327.400 447.600 ;
        RECT 329.200 447.400 330.000 453.000 ;
        RECT 328.000 446.800 330.000 447.400 ;
        RECT 330.800 455.400 331.600 459.800 ;
        RECT 335.000 458.400 336.200 459.800 ;
        RECT 335.000 457.800 336.400 458.400 ;
        RECT 339.600 457.800 340.400 459.800 ;
        RECT 344.000 458.400 344.800 459.800 ;
        RECT 344.000 457.800 346.000 458.400 ;
        RECT 335.600 457.000 336.400 457.800 ;
        RECT 339.800 457.200 340.400 457.800 ;
        RECT 339.800 456.600 342.600 457.200 ;
        RECT 341.800 456.400 342.600 456.600 ;
        RECT 343.600 455.600 344.400 457.200 ;
        RECT 345.200 457.000 346.000 457.800 ;
        RECT 333.800 455.400 334.600 455.600 ;
        RECT 330.800 454.800 334.600 455.400 ;
        RECT 330.800 451.400 331.600 454.800 ;
        RECT 337.800 454.200 338.600 454.400 ;
        RECT 343.600 454.200 344.200 455.600 ;
        RECT 348.400 455.000 349.200 459.800 ;
        RECT 350.000 455.600 350.800 457.200 ;
        RECT 346.800 454.200 348.400 454.400 ;
        RECT 337.400 453.600 348.400 454.200 ;
        RECT 335.600 452.800 336.400 453.000 ;
        RECT 332.600 452.200 336.400 452.800 ;
        RECT 332.600 452.000 333.400 452.200 ;
        RECT 334.200 451.400 335.000 451.600 ;
        RECT 330.800 450.800 335.000 451.400 ;
        RECT 319.600 442.200 320.400 445.000 ;
        RECT 321.200 442.200 322.000 445.000 ;
        RECT 324.400 442.200 325.200 446.800 ;
        RECT 328.000 446.200 328.600 446.800 ;
        RECT 327.600 445.600 328.600 446.200 ;
        RECT 327.600 442.200 328.400 445.600 ;
        RECT 330.800 442.200 331.600 450.800 ;
        RECT 337.400 450.400 338.000 453.600 ;
        RECT 344.600 453.400 345.400 453.600 ;
        RECT 343.600 452.400 344.400 452.600 ;
        RECT 346.200 452.400 347.000 452.600 ;
        RECT 342.000 451.800 347.000 452.400 ;
        RECT 342.000 451.600 342.800 451.800 ;
        RECT 343.600 451.000 349.200 451.200 ;
        RECT 343.400 450.800 349.200 451.000 ;
        RECT 335.600 449.800 338.000 450.400 ;
        RECT 339.400 450.600 349.200 450.800 ;
        RECT 339.400 450.200 344.200 450.600 ;
        RECT 335.600 448.800 336.200 449.800 ;
        RECT 334.800 448.000 336.200 448.800 ;
        RECT 337.800 449.000 338.600 449.200 ;
        RECT 339.400 449.000 340.000 450.200 ;
        RECT 337.800 448.400 340.000 449.000 ;
        RECT 340.600 449.000 346.000 449.600 ;
        RECT 340.600 448.800 341.400 449.000 ;
        RECT 345.200 448.800 346.000 449.000 ;
        RECT 339.000 447.400 339.800 447.600 ;
        RECT 341.800 447.400 342.600 447.600 ;
        RECT 335.600 446.200 336.400 447.000 ;
        RECT 339.000 446.800 342.600 447.400 ;
        RECT 339.800 446.200 340.400 446.800 ;
        RECT 345.200 446.200 346.000 447.000 ;
        RECT 335.000 442.200 336.200 446.200 ;
        RECT 339.600 442.200 340.400 446.200 ;
        RECT 344.000 445.600 346.000 446.200 ;
        RECT 344.000 442.200 344.800 445.600 ;
        RECT 348.400 442.200 349.200 450.600 ;
        RECT 351.600 442.200 352.400 459.800 ;
        RECT 353.200 455.200 354.000 459.800 ;
        RECT 356.400 456.400 357.200 459.800 ;
        RECT 356.400 455.800 357.400 456.400 ;
        RECT 359.600 456.000 360.400 459.800 ;
        RECT 362.800 456.000 363.600 459.800 ;
        RECT 359.600 455.800 363.600 456.000 ;
        RECT 364.400 455.800 365.200 459.800 ;
        RECT 366.000 457.000 366.800 459.000 ;
        RECT 353.200 454.600 355.800 455.200 ;
        RECT 353.400 452.400 354.200 453.200 ;
        RECT 353.200 451.600 354.200 452.400 ;
        RECT 355.200 453.000 355.800 454.600 ;
        RECT 356.800 454.400 357.400 455.800 ;
        RECT 359.800 455.400 363.400 455.800 ;
        RECT 360.400 454.400 361.200 454.800 ;
        RECT 364.400 454.400 365.000 455.800 ;
        RECT 366.000 454.800 366.600 457.000 ;
        RECT 370.200 456.400 371.000 459.000 ;
        RECT 369.200 456.000 371.000 456.400 ;
        RECT 375.600 457.000 376.400 459.000 ;
        RECT 369.200 455.600 371.800 456.000 ;
        RECT 370.200 455.400 371.800 455.600 ;
        RECT 371.000 455.000 371.800 455.400 ;
        RECT 356.400 454.300 357.400 454.400 ;
        RECT 358.000 454.300 358.800 454.400 ;
        RECT 359.600 454.300 361.200 454.400 ;
        RECT 356.400 453.800 361.200 454.300 ;
        RECT 356.400 453.700 360.400 453.800 ;
        RECT 356.400 453.600 357.400 453.700 ;
        RECT 358.000 453.600 358.800 453.700 ;
        RECT 359.600 453.600 360.400 453.700 ;
        RECT 362.600 453.600 365.200 454.400 ;
        RECT 366.000 454.200 370.200 454.800 ;
        RECT 369.200 453.800 370.200 454.200 ;
        RECT 371.200 454.400 371.800 455.000 ;
        RECT 375.600 454.800 376.200 457.000 ;
        RECT 379.800 456.000 380.600 459.000 ;
        RECT 385.200 456.000 386.000 459.800 ;
        RECT 388.400 456.000 389.200 459.800 ;
        RECT 379.800 455.400 381.400 456.000 ;
        RECT 385.200 455.800 389.200 456.000 ;
        RECT 390.000 455.800 390.800 459.800 ;
        RECT 385.400 455.400 389.000 455.800 ;
        RECT 380.600 455.000 381.400 455.400 ;
        RECT 355.200 452.200 356.200 453.000 ;
        RECT 355.200 450.200 355.800 452.200 ;
        RECT 356.800 450.200 357.400 453.600 ;
        RECT 361.200 451.600 362.000 453.200 ;
        RECT 362.600 452.400 363.200 453.600 ;
        RECT 362.600 451.600 363.600 452.400 ;
        RECT 366.000 451.600 366.800 453.200 ;
        RECT 367.600 451.600 368.400 453.200 ;
        RECT 369.200 453.000 370.600 453.800 ;
        RECT 371.200 453.600 373.200 454.400 ;
        RECT 375.600 454.200 379.800 454.800 ;
        RECT 378.800 453.800 379.800 454.200 ;
        RECT 380.800 454.400 381.400 455.000 ;
        RECT 386.000 454.400 386.800 454.800 ;
        RECT 390.000 454.400 390.600 455.800 ;
        RECT 391.600 455.000 392.400 459.800 ;
        RECT 396.000 458.400 396.800 459.800 ;
        RECT 394.800 457.800 396.800 458.400 ;
        RECT 400.400 457.800 401.200 459.800 ;
        RECT 404.600 458.400 405.800 459.800 ;
        RECT 404.400 457.800 405.800 458.400 ;
        RECT 394.800 457.000 395.600 457.800 ;
        RECT 400.400 457.200 401.000 457.800 ;
        RECT 396.400 456.400 397.200 457.200 ;
        RECT 398.200 456.600 401.000 457.200 ;
        RECT 404.400 457.000 405.200 457.800 ;
        RECT 398.200 456.400 399.000 456.600 ;
        RECT 362.600 450.200 363.200 451.600 ;
        RECT 369.200 451.000 369.800 453.000 ;
        RECT 366.000 450.400 369.800 451.000 ;
        RECT 364.400 450.200 365.200 450.400 ;
        RECT 353.200 449.600 355.800 450.200 ;
        RECT 353.200 442.200 354.000 449.600 ;
        RECT 356.400 449.200 357.400 450.200 ;
        RECT 362.200 449.600 363.200 450.200 ;
        RECT 363.800 449.600 365.200 450.200 ;
        RECT 356.400 442.200 357.200 449.200 ;
        RECT 362.200 442.200 363.000 449.600 ;
        RECT 363.800 448.400 364.400 449.600 ;
        RECT 363.600 447.600 364.400 448.400 ;
        RECT 366.000 447.000 366.600 450.400 ;
        RECT 371.200 449.800 371.800 453.600 ;
        RECT 372.400 450.800 373.200 452.400 ;
        RECT 375.600 451.600 376.400 453.200 ;
        RECT 377.200 451.600 378.000 453.200 ;
        RECT 378.800 453.000 380.200 453.800 ;
        RECT 380.800 453.600 382.800 454.400 ;
        RECT 383.600 454.300 384.400 454.400 ;
        RECT 385.200 454.300 386.800 454.400 ;
        RECT 383.600 453.800 386.800 454.300 ;
        RECT 383.600 453.700 386.000 453.800 ;
        RECT 383.600 453.600 384.400 453.700 ;
        RECT 385.200 453.600 386.000 453.700 ;
        RECT 388.200 453.600 390.800 454.400 ;
        RECT 392.400 454.200 394.000 454.400 ;
        RECT 396.600 454.200 397.200 456.400 ;
        RECT 406.200 455.400 407.000 455.600 ;
        RECT 409.200 455.400 410.000 459.800 ;
        RECT 410.800 455.600 411.600 459.800 ;
        RECT 412.400 456.000 413.200 459.800 ;
        RECT 415.600 456.000 416.400 459.800 ;
        RECT 412.400 455.800 416.400 456.000 ;
        RECT 417.200 455.800 418.000 459.800 ;
        RECT 418.800 456.000 419.600 459.800 ;
        RECT 422.000 456.000 422.800 459.800 ;
        RECT 418.800 455.800 422.800 456.000 ;
        RECT 423.600 455.800 424.400 459.800 ;
        RECT 425.200 456.000 426.000 459.800 ;
        RECT 428.400 456.000 429.200 459.800 ;
        RECT 425.200 455.800 429.200 456.000 ;
        RECT 430.000 456.000 430.800 459.800 ;
        RECT 433.200 456.000 434.000 459.800 ;
        RECT 430.000 455.800 434.000 456.000 ;
        RECT 434.800 455.800 435.600 459.800 ;
        RECT 436.400 456.000 437.200 459.800 ;
        RECT 439.600 456.000 440.400 459.800 ;
        RECT 436.400 455.800 440.400 456.000 ;
        RECT 441.200 455.800 442.000 459.800 ;
        RECT 406.200 454.800 410.000 455.400 ;
        RECT 398.000 454.200 398.800 454.400 ;
        RECT 402.200 454.200 403.000 454.400 ;
        RECT 392.400 453.600 403.400 454.200 ;
        RECT 378.800 451.000 379.400 453.000 ;
        RECT 370.200 449.200 371.800 449.800 ;
        RECT 375.600 450.400 379.400 451.000 ;
        RECT 366.000 443.000 366.800 447.000 ;
        RECT 370.200 442.200 371.000 449.200 ;
        RECT 375.600 447.000 376.200 450.400 ;
        RECT 380.800 449.800 381.400 453.600 ;
        RECT 382.000 452.300 382.800 452.400 ;
        RECT 385.200 452.300 386.000 452.400 ;
        RECT 382.000 451.700 386.000 452.300 ;
        RECT 382.000 450.800 382.800 451.700 ;
        RECT 385.200 451.600 386.000 451.700 ;
        RECT 386.800 451.600 387.600 453.200 ;
        RECT 388.200 450.200 388.800 453.600 ;
        RECT 395.400 453.400 396.200 453.600 ;
        RECT 393.800 452.400 394.600 452.600 ;
        RECT 393.800 452.300 398.800 452.400 ;
        RECT 399.600 452.300 400.400 452.400 ;
        RECT 393.800 451.800 400.400 452.300 ;
        RECT 398.000 451.700 400.400 451.800 ;
        RECT 398.000 451.600 398.800 451.700 ;
        RECT 399.600 451.600 400.400 451.700 ;
        RECT 391.600 451.000 397.200 451.200 ;
        RECT 391.600 450.800 397.400 451.000 ;
        RECT 391.600 450.600 401.400 450.800 ;
        RECT 390.000 450.200 390.800 450.400 ;
        RECT 379.800 449.200 381.400 449.800 ;
        RECT 387.800 449.600 388.800 450.200 ;
        RECT 389.400 449.600 390.800 450.200 ;
        RECT 375.600 443.000 376.400 447.000 ;
        RECT 379.800 442.200 380.600 449.200 ;
        RECT 387.800 442.200 388.600 449.600 ;
        RECT 389.400 448.400 390.000 449.600 ;
        RECT 389.200 447.600 390.000 448.400 ;
        RECT 391.600 442.200 392.400 450.600 ;
        RECT 396.600 450.200 401.400 450.600 ;
        RECT 394.800 449.000 400.200 449.600 ;
        RECT 394.800 448.800 395.600 449.000 ;
        RECT 399.400 448.800 400.200 449.000 ;
        RECT 400.800 449.000 401.400 450.200 ;
        RECT 402.800 450.400 403.400 453.600 ;
        RECT 404.400 452.800 405.200 453.000 ;
        RECT 404.400 452.200 408.200 452.800 ;
        RECT 407.400 452.000 408.200 452.200 ;
        RECT 405.800 451.400 406.600 451.600 ;
        RECT 409.200 451.400 410.000 454.800 ;
        RECT 411.000 454.400 411.600 455.600 ;
        RECT 412.600 455.400 416.200 455.800 ;
        RECT 414.800 454.400 415.600 454.800 ;
        RECT 417.400 454.400 418.000 455.800 ;
        RECT 419.000 455.400 422.600 455.800 ;
        RECT 421.200 454.400 422.000 454.800 ;
        RECT 423.800 454.400 424.400 455.800 ;
        RECT 425.400 455.400 429.000 455.800 ;
        RECT 430.200 455.400 433.800 455.800 ;
        RECT 427.600 454.400 428.400 454.800 ;
        RECT 430.800 454.400 431.600 454.800 ;
        RECT 434.800 454.400 435.400 455.800 ;
        RECT 436.600 455.400 440.200 455.800 ;
        RECT 437.200 454.400 438.000 454.800 ;
        RECT 441.200 454.400 441.800 455.800 ;
        RECT 410.800 453.600 413.400 454.400 ;
        RECT 414.800 453.800 416.400 454.400 ;
        RECT 415.600 453.600 416.400 453.800 ;
        RECT 417.200 453.600 419.800 454.400 ;
        RECT 421.200 453.800 422.800 454.400 ;
        RECT 422.000 453.600 422.800 453.800 ;
        RECT 423.600 453.600 426.200 454.400 ;
        RECT 427.600 453.800 429.200 454.400 ;
        RECT 428.400 453.600 429.200 453.800 ;
        RECT 430.000 453.800 431.600 454.400 ;
        RECT 430.000 453.600 430.800 453.800 ;
        RECT 433.000 453.600 435.600 454.400 ;
        RECT 436.400 453.800 438.000 454.400 ;
        RECT 436.400 453.600 437.200 453.800 ;
        RECT 439.400 453.600 442.000 454.400 ;
        RECT 446.400 454.200 447.200 459.800 ;
        RECT 452.800 454.200 453.600 459.800 ;
        RECT 455.600 455.600 456.400 457.200 ;
        RECT 457.200 454.300 458.000 459.800 ;
        RECT 463.600 456.000 464.400 459.800 ;
        RECT 466.800 456.000 467.600 459.800 ;
        RECT 463.600 455.800 467.600 456.000 ;
        RECT 468.400 455.800 469.200 459.800 ;
        RECT 470.000 456.000 470.800 459.800 ;
        RECT 473.200 456.000 474.000 459.800 ;
        RECT 470.000 455.800 474.000 456.000 ;
        RECT 474.800 455.800 475.600 459.800 ;
        RECT 476.400 455.800 477.200 459.800 ;
        RECT 478.000 456.000 478.800 459.800 ;
        RECT 481.200 456.000 482.000 459.800 ;
        RECT 478.000 455.800 482.000 456.000 ;
        RECT 482.800 457.000 483.600 459.000 ;
        RECT 463.800 455.400 467.400 455.800 ;
        RECT 464.400 454.400 465.200 454.800 ;
        RECT 468.400 454.400 469.000 455.800 ;
        RECT 470.200 455.400 473.800 455.800 ;
        RECT 470.800 454.400 471.600 454.800 ;
        RECT 474.800 454.400 475.400 455.800 ;
        RECT 476.600 454.400 477.200 455.800 ;
        RECT 478.200 455.400 481.800 455.800 ;
        RECT 482.800 454.800 483.400 457.000 ;
        RECT 487.000 456.400 487.800 459.000 ;
        RECT 486.000 456.000 487.800 456.400 ;
        RECT 486.000 455.600 488.600 456.000 ;
        RECT 492.400 455.800 493.200 459.800 ;
        RECT 494.000 456.000 494.800 459.800 ;
        RECT 497.200 456.000 498.000 459.800 ;
        RECT 494.000 455.800 498.000 456.000 ;
        RECT 498.800 456.000 499.600 459.800 ;
        RECT 502.000 456.000 502.800 459.800 ;
        RECT 498.800 455.800 502.800 456.000 ;
        RECT 503.600 455.800 504.400 459.800 ;
        RECT 506.800 457.600 507.600 459.800 ;
        RECT 487.000 455.400 488.600 455.600 ;
        RECT 487.800 455.000 488.600 455.400 ;
        RECT 480.400 454.400 481.200 454.800 ;
        RECT 463.600 454.300 465.200 454.400 ;
        RECT 446.400 453.800 448.200 454.200 ;
        RECT 452.800 453.800 454.600 454.200 ;
        RECT 446.600 453.600 448.200 453.800 ;
        RECT 453.000 453.600 454.600 453.800 ;
        RECT 405.800 450.800 410.000 451.400 ;
        RECT 402.800 449.800 405.200 450.400 ;
        RECT 402.200 449.000 403.000 449.200 ;
        RECT 400.800 448.400 403.000 449.000 ;
        RECT 404.600 448.800 405.200 449.800 ;
        RECT 404.600 448.000 406.000 448.800 ;
        RECT 398.200 447.400 399.000 447.600 ;
        RECT 401.000 447.400 401.800 447.600 ;
        RECT 394.800 446.200 395.600 447.000 ;
        RECT 398.200 446.800 401.800 447.400 ;
        RECT 400.400 446.200 401.000 446.800 ;
        RECT 404.400 446.200 405.200 447.000 ;
        RECT 394.800 445.600 396.800 446.200 ;
        RECT 396.000 442.200 396.800 445.600 ;
        RECT 400.400 442.200 401.200 446.200 ;
        RECT 404.600 442.200 405.800 446.200 ;
        RECT 409.200 442.200 410.000 450.800 ;
        RECT 410.800 450.200 411.600 450.400 ;
        RECT 412.800 450.200 413.400 453.600 ;
        RECT 414.000 451.600 414.800 453.200 ;
        RECT 417.200 450.200 418.000 450.400 ;
        RECT 419.200 450.200 419.800 453.600 ;
        RECT 420.400 451.600 421.200 453.200 ;
        RECT 423.600 450.200 424.400 450.400 ;
        RECT 425.600 450.200 426.200 453.600 ;
        RECT 426.800 451.600 427.600 453.200 ;
        RECT 431.600 451.600 432.400 453.200 ;
        RECT 433.000 450.200 433.600 453.600 ;
        RECT 438.000 451.600 438.800 453.200 ;
        RECT 434.800 450.200 435.600 450.400 ;
        RECT 439.400 450.200 440.000 453.600 ;
        RECT 444.400 451.600 446.000 452.400 ;
        RECT 441.200 450.200 442.000 450.400 ;
        RECT 410.800 449.600 412.200 450.200 ;
        RECT 412.800 449.600 413.800 450.200 ;
        RECT 417.200 449.600 418.600 450.200 ;
        RECT 419.200 449.600 420.200 450.200 ;
        RECT 423.600 449.600 425.000 450.200 ;
        RECT 425.600 449.600 426.600 450.200 ;
        RECT 411.600 448.400 412.200 449.600 ;
        RECT 411.600 447.600 412.400 448.400 ;
        RECT 413.000 442.200 413.800 449.600 ;
        RECT 418.000 448.400 418.600 449.600 ;
        RECT 418.000 447.600 418.800 448.400 ;
        RECT 419.400 444.400 420.200 449.600 ;
        RECT 424.400 448.400 425.000 449.600 ;
        RECT 424.400 447.600 425.200 448.400 ;
        RECT 425.800 444.400 426.600 449.600 ;
        RECT 432.600 449.600 433.600 450.200 ;
        RECT 434.200 449.600 435.600 450.200 ;
        RECT 439.000 449.600 440.000 450.200 ;
        RECT 440.600 449.600 442.000 450.200 ;
        RECT 442.800 450.300 443.600 451.200 ;
        RECT 447.600 450.400 448.200 453.600 ;
        RECT 450.800 451.600 452.400 452.400 ;
        RECT 444.400 450.300 445.200 450.400 ;
        RECT 442.800 449.700 445.200 450.300 ;
        RECT 442.800 449.600 443.600 449.700 ;
        RECT 444.400 449.600 445.200 449.700 ;
        RECT 447.600 449.600 448.400 450.400 ;
        RECT 449.200 449.600 450.000 451.200 ;
        RECT 454.000 450.400 454.600 453.600 ;
        RECT 457.200 453.800 465.200 454.300 ;
        RECT 457.200 453.700 464.400 453.800 ;
        RECT 454.000 449.600 454.800 450.400 ;
        RECT 432.600 444.400 433.400 449.600 ;
        RECT 434.200 448.400 434.800 449.600 ;
        RECT 434.000 447.600 434.800 448.400 ;
        RECT 419.400 443.600 421.200 444.400 ;
        RECT 425.800 443.600 427.600 444.400 ;
        RECT 431.600 443.600 433.400 444.400 ;
        RECT 419.400 442.200 420.200 443.600 ;
        RECT 425.800 442.200 426.600 443.600 ;
        RECT 432.600 442.200 433.400 443.600 ;
        RECT 439.000 442.200 439.800 449.600 ;
        RECT 440.600 448.400 441.200 449.600 ;
        RECT 440.400 447.600 441.200 448.400 ;
        RECT 446.000 447.600 446.800 449.200 ;
        RECT 447.600 447.000 448.200 449.600 ;
        RECT 452.400 447.600 453.200 449.200 ;
        RECT 454.000 447.000 454.600 449.600 ;
        RECT 444.600 446.400 448.200 447.000 ;
        RECT 444.600 446.200 445.200 446.400 ;
        RECT 444.400 442.200 445.200 446.200 ;
        RECT 447.600 446.200 448.200 446.400 ;
        RECT 451.000 446.400 454.600 447.000 ;
        RECT 451.000 446.200 451.600 446.400 ;
        RECT 447.600 442.200 448.400 446.200 ;
        RECT 450.800 442.200 451.600 446.200 ;
        RECT 454.000 446.200 454.600 446.400 ;
        RECT 454.000 442.200 454.800 446.200 ;
        RECT 457.200 442.200 458.000 453.700 ;
        RECT 463.600 453.600 464.400 453.700 ;
        RECT 466.600 453.600 469.200 454.400 ;
        RECT 470.000 453.800 471.600 454.400 ;
        RECT 470.000 453.600 470.800 453.800 ;
        RECT 473.000 453.600 475.600 454.400 ;
        RECT 476.400 453.600 479.000 454.400 ;
        RECT 480.400 453.800 482.000 454.400 ;
        RECT 482.800 454.200 487.000 454.800 ;
        RECT 481.200 453.600 482.000 453.800 ;
        RECT 486.000 453.800 487.000 454.200 ;
        RECT 488.000 454.400 488.600 455.000 ;
        RECT 492.600 454.400 493.200 455.800 ;
        RECT 494.200 455.400 497.800 455.800 ;
        RECT 499.000 455.400 502.600 455.800 ;
        RECT 496.400 454.400 497.200 454.800 ;
        RECT 499.600 454.400 500.400 454.800 ;
        RECT 503.600 454.400 504.200 455.800 ;
        RECT 506.800 454.400 507.400 457.600 ;
        RECT 508.400 455.600 509.200 457.200 ;
        RECT 463.600 452.300 464.400 452.400 ;
        RECT 465.200 452.300 466.000 453.200 ;
        RECT 463.600 451.700 466.000 452.300 ;
        RECT 463.600 451.600 464.400 451.700 ;
        RECT 465.200 451.600 466.000 451.700 ;
        RECT 466.600 450.200 467.200 453.600 ;
        RECT 471.600 451.600 472.400 453.200 ;
        RECT 473.000 452.300 473.600 453.600 ;
        RECT 473.000 451.700 477.100 452.300 ;
        RECT 468.400 450.200 469.200 450.400 ;
        RECT 473.000 450.200 473.600 451.700 ;
        RECT 476.500 450.400 477.100 451.700 ;
        RECT 474.800 450.200 475.600 450.400 ;
        RECT 466.200 449.600 467.200 450.200 ;
        RECT 467.800 449.600 469.200 450.200 ;
        RECT 472.600 449.600 473.600 450.200 ;
        RECT 474.200 449.600 475.600 450.200 ;
        RECT 476.400 450.200 477.200 450.400 ;
        RECT 478.400 450.200 479.000 453.600 ;
        RECT 479.600 451.600 480.400 453.200 ;
        RECT 482.800 451.600 483.600 453.200 ;
        RECT 484.400 451.600 485.200 453.200 ;
        RECT 486.000 453.000 487.400 453.800 ;
        RECT 488.000 453.600 490.000 454.400 ;
        RECT 492.400 453.600 495.000 454.400 ;
        RECT 496.400 453.800 498.000 454.400 ;
        RECT 497.200 453.600 498.000 453.800 ;
        RECT 498.800 453.800 500.400 454.400 ;
        RECT 501.800 454.300 504.400 454.400 ;
        RECT 505.200 454.300 506.000 454.400 ;
        RECT 498.800 453.600 499.600 453.800 ;
        RECT 501.800 453.700 506.000 454.300 ;
        RECT 501.800 453.600 504.400 453.700 ;
        RECT 505.200 453.600 506.000 453.700 ;
        RECT 506.800 453.600 507.600 454.400 ;
        RECT 511.200 454.200 512.000 459.800 ;
        RECT 516.400 455.800 517.200 459.800 ;
        RECT 518.000 456.000 518.800 459.800 ;
        RECT 521.200 456.000 522.000 459.800 ;
        RECT 518.000 455.800 522.000 456.000 ;
        RECT 516.600 454.400 517.200 455.800 ;
        RECT 518.200 455.400 521.800 455.800 ;
        RECT 522.800 455.600 523.600 457.200 ;
        RECT 520.400 454.400 521.200 454.800 ;
        RECT 510.200 453.800 512.000 454.200 ;
        RECT 510.200 453.600 511.800 453.800 ;
        RECT 516.400 453.600 519.000 454.400 ;
        RECT 520.400 454.300 522.000 454.400 ;
        RECT 524.400 454.300 525.200 459.800 ;
        RECT 526.000 455.800 526.800 459.800 ;
        RECT 527.600 456.000 528.400 459.800 ;
        RECT 530.800 456.000 531.600 459.800 ;
        RECT 527.600 455.800 531.600 456.000 ;
        RECT 526.200 454.400 526.800 455.800 ;
        RECT 527.800 455.400 531.400 455.800 ;
        RECT 532.400 455.200 533.200 459.800 ;
        RECT 535.600 456.400 536.400 459.800 ;
        RECT 535.600 455.800 536.600 456.400 ;
        RECT 540.400 456.000 541.200 459.800 ;
        RECT 530.000 454.400 530.800 454.800 ;
        RECT 532.400 454.600 535.000 455.200 ;
        RECT 520.400 453.800 525.200 454.300 ;
        RECT 521.200 453.700 525.200 453.800 ;
        RECT 521.200 453.600 522.000 453.700 ;
        RECT 486.000 451.000 486.600 453.000 ;
        RECT 482.800 450.400 486.600 451.000 ;
        RECT 476.400 449.600 477.800 450.200 ;
        RECT 478.400 449.600 479.400 450.200 ;
        RECT 466.200 444.400 467.000 449.600 ;
        RECT 467.800 448.400 468.400 449.600 ;
        RECT 467.600 447.600 468.400 448.400 ;
        RECT 465.200 443.600 467.000 444.400 ;
        RECT 466.200 442.200 467.000 443.600 ;
        RECT 472.600 442.200 473.400 449.600 ;
        RECT 474.200 448.400 474.800 449.600 ;
        RECT 474.000 447.600 474.800 448.400 ;
        RECT 477.200 448.400 477.800 449.600 ;
        RECT 477.200 447.600 478.000 448.400 ;
        RECT 478.600 442.200 479.400 449.600 ;
        RECT 482.800 447.000 483.400 450.400 ;
        RECT 488.000 449.800 488.600 453.600 ;
        RECT 489.200 450.800 490.000 452.400 ;
        RECT 487.000 449.200 488.600 449.800 ;
        RECT 492.400 450.200 493.200 450.400 ;
        RECT 494.400 450.200 495.000 453.600 ;
        RECT 495.600 451.600 496.400 453.200 ;
        RECT 500.400 451.600 501.200 453.200 ;
        RECT 501.800 450.200 502.400 453.600 ;
        RECT 505.200 450.800 506.000 452.400 ;
        RECT 503.600 450.200 504.400 450.400 ;
        RECT 506.800 450.200 507.400 453.600 ;
        RECT 510.200 450.400 510.800 453.600 ;
        RECT 518.400 452.400 519.000 453.600 ;
        RECT 512.400 451.600 514.000 452.400 ;
        RECT 518.000 451.600 519.000 452.400 ;
        RECT 519.600 451.600 520.400 453.200 ;
        RECT 492.400 449.600 493.800 450.200 ;
        RECT 494.400 449.600 495.400 450.200 ;
        RECT 482.800 443.000 483.600 447.000 ;
        RECT 487.000 442.200 487.800 449.200 ;
        RECT 493.200 448.400 493.800 449.600 ;
        RECT 493.200 447.600 494.000 448.400 ;
        RECT 494.600 442.200 495.400 449.600 ;
        RECT 501.400 449.600 502.400 450.200 ;
        RECT 503.000 449.600 504.400 450.200 ;
        RECT 501.400 442.200 502.200 449.600 ;
        RECT 503.000 448.400 503.600 449.600 ;
        RECT 502.800 447.600 503.600 448.400 ;
        RECT 505.800 449.400 507.600 450.200 ;
        RECT 510.000 449.600 510.800 450.400 ;
        RECT 514.800 449.600 515.600 451.200 ;
        RECT 516.400 450.200 517.200 450.400 ;
        RECT 518.400 450.200 519.000 451.600 ;
        RECT 516.400 449.600 517.800 450.200 ;
        RECT 518.400 449.600 519.400 450.200 ;
        RECT 505.800 442.200 506.600 449.400 ;
        RECT 510.200 447.000 510.800 449.600 ;
        RECT 511.600 447.600 512.400 449.200 ;
        RECT 517.200 448.400 517.800 449.600 ;
        RECT 517.200 447.600 518.000 448.400 ;
        RECT 510.200 446.400 513.800 447.000 ;
        RECT 510.200 446.200 510.800 446.400 ;
        RECT 510.000 442.200 510.800 446.200 ;
        RECT 513.200 442.200 514.000 446.400 ;
        RECT 518.600 442.200 519.400 449.600 ;
        RECT 524.400 442.200 525.200 453.700 ;
        RECT 526.000 453.600 528.600 454.400 ;
        RECT 530.000 453.800 531.600 454.400 ;
        RECT 530.800 453.600 531.600 453.800 ;
        RECT 526.000 450.200 526.800 450.400 ;
        RECT 528.000 450.200 528.600 453.600 ;
        RECT 529.200 451.600 530.000 453.200 ;
        RECT 532.600 452.400 533.400 453.200 ;
        RECT 532.400 451.600 533.400 452.400 ;
        RECT 534.400 453.000 535.000 454.600 ;
        RECT 536.000 454.400 536.600 455.800 ;
        RECT 535.600 453.600 536.600 454.400 ;
        RECT 534.400 452.200 535.400 453.000 ;
        RECT 534.400 450.200 535.000 452.200 ;
        RECT 536.000 450.200 536.600 453.600 ;
        RECT 526.000 449.600 527.400 450.200 ;
        RECT 528.000 449.600 529.000 450.200 ;
        RECT 526.800 448.400 527.400 449.600 ;
        RECT 526.800 447.600 527.600 448.400 ;
        RECT 528.200 444.400 529.000 449.600 ;
        RECT 532.400 449.600 535.000 450.200 ;
        RECT 528.200 443.600 530.000 444.400 ;
        RECT 528.200 442.200 529.000 443.600 ;
        RECT 532.400 442.200 533.200 449.600 ;
        RECT 535.600 449.200 536.600 450.200 ;
        RECT 540.200 455.200 541.200 456.000 ;
        RECT 540.200 450.800 541.000 455.200 ;
        RECT 542.000 454.600 542.800 459.800 ;
        RECT 548.400 456.600 549.200 459.800 ;
        RECT 550.000 457.000 550.800 459.800 ;
        RECT 551.600 457.000 552.400 459.800 ;
        RECT 553.200 457.000 554.000 459.800 ;
        RECT 554.800 457.000 555.600 459.800 ;
        RECT 558.000 457.000 558.800 459.800 ;
        RECT 561.200 457.000 562.000 459.800 ;
        RECT 562.800 457.000 563.600 459.800 ;
        RECT 564.400 457.000 565.200 459.800 ;
        RECT 546.800 455.800 549.200 456.600 ;
        RECT 566.000 456.600 566.800 459.800 ;
        RECT 546.800 455.200 547.600 455.800 ;
        RECT 541.600 454.000 542.800 454.600 ;
        RECT 545.800 454.600 547.600 455.200 ;
        RECT 551.600 455.600 552.600 456.400 ;
        RECT 555.600 455.600 557.200 456.400 ;
        RECT 558.000 455.800 562.600 456.400 ;
        RECT 566.000 455.800 568.600 456.600 ;
        RECT 558.000 455.600 558.800 455.800 ;
        RECT 541.600 452.000 542.200 454.000 ;
        RECT 545.800 453.400 546.600 454.600 ;
        RECT 542.800 452.600 546.600 453.400 ;
        RECT 551.600 452.800 552.400 455.600 ;
        RECT 558.000 454.800 558.800 455.000 ;
        RECT 554.400 454.200 558.800 454.800 ;
        RECT 554.400 454.000 555.200 454.200 ;
        RECT 559.600 453.600 560.400 455.200 ;
        RECT 561.800 453.400 562.600 455.800 ;
        RECT 567.800 455.200 568.600 455.800 ;
        RECT 567.800 454.400 570.800 455.200 ;
        RECT 572.400 453.800 573.200 459.800 ;
        RECT 575.600 456.000 576.400 459.800 ;
        RECT 554.800 452.600 558.000 453.400 ;
        RECT 561.800 452.600 563.800 453.400 ;
        RECT 564.400 453.000 573.200 453.800 ;
        RECT 548.400 452.000 549.200 452.600 ;
        RECT 559.600 452.000 560.400 452.400 ;
        RECT 566.000 452.000 566.800 452.400 ;
        RECT 571.000 452.000 571.800 452.200 ;
        RECT 541.600 451.400 542.400 452.000 ;
        RECT 548.400 451.400 571.800 452.000 ;
        RECT 540.200 450.000 541.200 450.800 ;
        RECT 535.600 442.200 536.400 449.200 ;
        RECT 540.400 442.200 541.200 450.000 ;
        RECT 541.800 449.600 542.400 451.400 ;
        RECT 541.800 449.000 550.800 449.600 ;
        RECT 541.800 447.400 542.400 449.000 ;
        RECT 550.000 448.800 550.800 449.000 ;
        RECT 553.200 449.000 561.800 449.600 ;
        RECT 553.200 448.800 554.000 449.000 ;
        RECT 545.000 447.600 547.600 448.400 ;
        RECT 541.800 446.800 544.400 447.400 ;
        RECT 543.600 442.200 544.400 446.800 ;
        RECT 546.800 442.200 547.600 447.600 ;
        RECT 548.200 446.800 552.400 447.600 ;
        RECT 550.000 442.200 550.800 445.000 ;
        RECT 551.600 442.200 552.400 445.000 ;
        RECT 553.200 442.200 554.000 445.000 ;
        RECT 554.800 442.200 555.600 448.400 ;
        RECT 558.000 447.600 560.600 448.400 ;
        RECT 561.200 448.200 561.800 449.000 ;
        RECT 562.800 449.400 563.600 449.600 ;
        RECT 562.800 449.000 568.200 449.400 ;
        RECT 562.800 448.800 569.000 449.000 ;
        RECT 567.600 448.200 569.000 448.800 ;
        RECT 561.200 447.600 567.000 448.200 ;
        RECT 570.000 448.000 571.600 448.800 ;
        RECT 570.000 447.600 570.600 448.000 ;
        RECT 558.000 442.200 558.800 447.000 ;
        RECT 561.200 442.200 562.000 447.000 ;
        RECT 566.400 446.800 570.600 447.600 ;
        RECT 572.400 447.400 573.200 453.000 ;
        RECT 575.400 455.200 576.400 456.000 ;
        RECT 575.400 450.800 576.200 455.200 ;
        RECT 577.200 454.600 578.000 459.800 ;
        RECT 583.600 456.600 584.400 459.800 ;
        RECT 585.200 457.000 586.000 459.800 ;
        RECT 586.800 457.000 587.600 459.800 ;
        RECT 588.400 457.000 589.200 459.800 ;
        RECT 590.000 457.000 590.800 459.800 ;
        RECT 593.200 457.000 594.000 459.800 ;
        RECT 596.400 457.000 597.200 459.800 ;
        RECT 598.000 457.000 598.800 459.800 ;
        RECT 599.600 457.000 600.400 459.800 ;
        RECT 582.000 455.800 584.400 456.600 ;
        RECT 601.200 456.600 602.000 459.800 ;
        RECT 582.000 455.200 582.800 455.800 ;
        RECT 576.800 454.000 578.000 454.600 ;
        RECT 581.000 454.600 582.800 455.200 ;
        RECT 586.800 455.600 587.800 456.400 ;
        RECT 590.800 455.600 592.400 456.400 ;
        RECT 593.200 455.800 597.800 456.400 ;
        RECT 601.200 455.800 603.800 456.600 ;
        RECT 593.200 455.600 594.000 455.800 ;
        RECT 576.800 452.000 577.400 454.000 ;
        RECT 581.000 453.400 581.800 454.600 ;
        RECT 578.000 452.600 581.800 453.400 ;
        RECT 586.800 452.800 587.600 455.600 ;
        RECT 593.200 454.800 594.000 455.000 ;
        RECT 589.600 454.200 594.000 454.800 ;
        RECT 589.600 454.000 590.400 454.200 ;
        RECT 594.800 453.600 595.600 455.200 ;
        RECT 597.000 453.400 597.800 455.800 ;
        RECT 603.000 455.200 603.800 455.800 ;
        RECT 603.000 454.400 606.000 455.200 ;
        RECT 607.600 453.800 608.400 459.800 ;
        RECT 590.000 452.600 593.200 453.400 ;
        RECT 597.000 452.600 599.000 453.400 ;
        RECT 599.600 453.000 608.400 453.800 ;
        RECT 583.600 452.000 584.400 452.600 ;
        RECT 601.200 452.000 602.000 452.400 ;
        RECT 606.200 452.000 607.000 452.200 ;
        RECT 576.800 451.400 577.600 452.000 ;
        RECT 583.600 451.400 607.000 452.000 ;
        RECT 575.400 450.000 576.400 450.800 ;
        RECT 571.200 446.800 573.200 447.400 ;
        RECT 562.800 442.200 563.600 445.000 ;
        RECT 564.400 442.200 565.200 445.000 ;
        RECT 567.600 442.200 568.400 446.800 ;
        RECT 571.200 446.200 571.800 446.800 ;
        RECT 570.800 445.600 571.800 446.200 ;
        RECT 570.800 442.200 571.600 445.600 ;
        RECT 575.600 442.200 576.400 450.000 ;
        RECT 577.000 449.600 577.600 451.400 ;
        RECT 577.000 449.000 586.000 449.600 ;
        RECT 577.000 447.400 577.600 449.000 ;
        RECT 585.200 448.800 586.000 449.000 ;
        RECT 588.400 449.000 597.000 449.600 ;
        RECT 588.400 448.800 589.200 449.000 ;
        RECT 580.200 447.600 582.800 448.400 ;
        RECT 577.000 446.800 579.600 447.400 ;
        RECT 578.800 442.200 579.600 446.800 ;
        RECT 582.000 442.200 582.800 447.600 ;
        RECT 583.400 446.800 587.600 447.600 ;
        RECT 585.200 442.200 586.000 445.000 ;
        RECT 586.800 442.200 587.600 445.000 ;
        RECT 588.400 442.200 589.200 445.000 ;
        RECT 590.000 442.200 590.800 448.400 ;
        RECT 593.200 447.600 595.800 448.400 ;
        RECT 596.400 448.200 597.000 449.000 ;
        RECT 598.000 449.400 598.800 449.600 ;
        RECT 598.000 449.000 603.400 449.400 ;
        RECT 598.000 448.800 604.200 449.000 ;
        RECT 602.800 448.200 604.200 448.800 ;
        RECT 596.400 447.600 602.200 448.200 ;
        RECT 605.200 448.000 606.800 448.800 ;
        RECT 605.200 447.600 605.800 448.000 ;
        RECT 593.200 442.200 594.000 447.000 ;
        RECT 596.400 442.200 597.200 447.000 ;
        RECT 601.600 446.800 605.800 447.600 ;
        RECT 607.600 447.400 608.400 453.000 ;
        RECT 606.400 446.800 608.400 447.400 ;
        RECT 598.000 442.200 598.800 445.000 ;
        RECT 599.600 442.200 600.400 445.000 ;
        RECT 602.800 442.200 603.600 446.800 ;
        RECT 606.400 446.200 607.000 446.800 ;
        RECT 606.000 445.600 607.000 446.200 ;
        RECT 606.000 442.200 606.800 445.600 ;
        RECT 2.800 428.300 3.600 439.800 ;
        RECT 7.000 432.400 7.800 439.800 ;
        RECT 8.400 433.600 9.200 434.400 ;
        RECT 8.600 432.400 9.200 433.600 ;
        RECT 7.000 431.800 8.000 432.400 ;
        RECT 8.600 431.800 10.000 432.400 ;
        RECT 6.000 428.800 6.800 430.400 ;
        RECT 7.400 428.400 8.000 431.800 ;
        RECT 9.200 431.600 10.000 431.800 ;
        RECT 12.400 431.200 13.200 439.800 ;
        RECT 15.600 431.200 16.400 439.800 ;
        RECT 18.800 431.200 19.600 439.800 ;
        RECT 22.000 431.200 22.800 439.800 ;
        RECT 27.400 438.400 28.200 439.800 ;
        RECT 27.400 437.600 29.200 438.400 ;
        RECT 26.000 433.600 26.800 434.400 ;
        RECT 26.000 432.400 26.600 433.600 ;
        RECT 27.400 432.400 28.200 437.600 ;
        RECT 25.200 431.800 26.600 432.400 ;
        RECT 27.200 431.800 28.200 432.400 ;
        RECT 25.200 431.600 26.000 431.800 ;
        RECT 12.400 430.400 14.200 431.200 ;
        RECT 15.600 430.400 17.800 431.200 ;
        RECT 18.800 430.400 21.000 431.200 ;
        RECT 22.000 430.400 24.400 431.200 ;
        RECT 13.400 429.000 14.200 430.400 ;
        RECT 17.000 429.000 17.800 430.400 ;
        RECT 20.200 429.000 21.000 430.400 ;
        RECT 4.400 428.300 5.200 428.400 ;
        RECT 2.800 428.200 5.200 428.300 ;
        RECT 2.800 427.700 6.000 428.200 ;
        RECT 2.800 422.200 3.600 427.700 ;
        RECT 4.400 427.600 6.000 427.700 ;
        RECT 7.400 427.600 10.000 428.400 ;
        RECT 10.800 428.200 12.600 429.000 ;
        RECT 13.400 428.200 16.000 429.000 ;
        RECT 17.000 428.200 19.400 429.000 ;
        RECT 20.200 428.200 22.800 429.000 ;
        RECT 10.800 427.600 11.600 428.200 ;
        RECT 13.400 427.600 14.200 428.200 ;
        RECT 17.000 427.600 17.800 428.200 ;
        RECT 20.200 427.600 21.000 428.200 ;
        RECT 23.600 427.600 24.400 430.400 ;
        RECT 27.200 428.400 27.800 431.800 ;
        RECT 31.600 431.200 32.400 439.800 ;
        RECT 35.800 432.400 36.600 439.800 ;
        RECT 35.800 431.800 37.200 432.400 ;
        RECT 31.600 430.800 35.600 431.200 ;
        RECT 31.600 430.600 35.800 430.800 ;
        RECT 28.400 428.800 29.200 430.400 ;
        RECT 35.000 430.000 35.800 430.600 ;
        RECT 36.600 430.400 37.200 431.800 ;
        RECT 39.600 431.200 40.400 439.800 ;
        RECT 42.800 431.200 43.600 439.800 ;
        RECT 46.000 431.200 46.800 439.800 ;
        RECT 49.200 431.200 50.000 439.800 ;
        RECT 52.400 431.400 53.200 439.800 ;
        RECT 56.800 436.400 57.600 439.800 ;
        RECT 55.600 435.800 57.600 436.400 ;
        RECT 61.200 435.800 62.000 439.800 ;
        RECT 65.400 435.800 66.600 439.800 ;
        RECT 55.600 435.000 56.400 435.800 ;
        RECT 61.200 435.200 61.800 435.800 ;
        RECT 59.000 434.600 62.600 435.200 ;
        RECT 65.200 435.000 66.000 435.800 ;
        RECT 59.000 434.400 59.800 434.600 ;
        RECT 61.800 434.400 62.600 434.600 ;
        RECT 66.200 434.000 67.600 434.400 ;
        RECT 65.400 433.600 67.600 434.000 ;
        RECT 55.600 433.000 56.400 433.200 ;
        RECT 60.200 433.000 61.000 433.200 ;
        RECT 55.600 432.400 61.000 433.000 ;
        RECT 61.600 433.000 63.800 433.600 ;
        RECT 61.600 431.800 62.200 433.000 ;
        RECT 63.000 432.800 63.800 433.000 ;
        RECT 65.400 433.200 66.800 433.600 ;
        RECT 65.400 432.200 66.000 433.200 ;
        RECT 57.400 431.400 62.200 431.800 ;
        RECT 52.400 431.200 62.200 431.400 ;
        RECT 63.600 431.600 66.000 432.200 ;
        RECT 39.600 430.400 41.400 431.200 ;
        RECT 42.800 430.400 45.000 431.200 ;
        RECT 46.000 430.400 48.200 431.200 ;
        RECT 49.200 430.400 51.600 431.200 ;
        RECT 52.400 431.000 58.200 431.200 ;
        RECT 52.400 430.800 58.000 431.000 ;
        RECT 33.600 428.400 34.400 429.200 ;
        RECT 25.200 427.600 27.800 428.400 ;
        RECT 30.000 428.300 30.800 428.400 ;
        RECT 30.000 428.200 32.300 428.300 ;
        RECT 29.200 427.700 32.300 428.200 ;
        RECT 29.200 427.600 30.800 427.700 ;
        RECT 5.200 427.200 6.000 427.600 ;
        RECT 4.600 426.200 8.200 426.600 ;
        RECT 9.200 426.200 9.800 427.600 ;
        RECT 12.400 426.800 14.200 427.600 ;
        RECT 15.600 426.800 17.800 427.600 ;
        RECT 18.800 426.800 21.000 427.600 ;
        RECT 22.000 426.800 24.400 427.600 ;
        RECT 4.400 426.000 8.400 426.200 ;
        RECT 4.400 422.200 5.200 426.000 ;
        RECT 7.600 422.200 8.400 426.000 ;
        RECT 9.200 422.200 10.000 426.200 ;
        RECT 12.400 422.200 13.200 426.800 ;
        RECT 15.600 422.200 16.400 426.800 ;
        RECT 18.800 422.200 19.600 426.800 ;
        RECT 22.000 422.200 22.800 426.800 ;
        RECT 25.400 426.200 26.000 427.600 ;
        RECT 29.200 427.200 30.000 427.600 ;
        RECT 27.000 426.200 30.600 426.600 ;
        RECT 31.700 426.400 32.300 427.700 ;
        RECT 33.200 427.600 34.200 428.400 ;
        RECT 35.200 427.000 35.800 430.000 ;
        RECT 36.400 429.600 37.200 430.400 ;
        RECT 33.400 426.400 35.800 427.000 ;
        RECT 25.200 422.200 26.000 426.200 ;
        RECT 26.800 426.000 30.800 426.200 ;
        RECT 26.800 422.200 27.600 426.000 ;
        RECT 30.000 422.200 30.800 426.000 ;
        RECT 31.600 424.800 32.400 426.400 ;
        RECT 33.400 424.200 34.000 426.400 ;
        RECT 36.600 426.200 37.200 429.600 ;
        RECT 40.600 429.000 41.400 430.400 ;
        RECT 44.200 429.000 45.000 430.400 ;
        RECT 47.400 429.000 48.200 430.400 ;
        RECT 38.000 428.200 39.800 429.000 ;
        RECT 40.600 428.200 43.200 429.000 ;
        RECT 44.200 428.200 46.600 429.000 ;
        RECT 47.400 428.200 50.000 429.000 ;
        RECT 38.000 427.600 38.800 428.200 ;
        RECT 40.600 427.600 41.400 428.200 ;
        RECT 44.200 427.600 45.000 428.200 ;
        RECT 47.400 427.600 48.200 428.200 ;
        RECT 50.800 427.600 51.600 430.400 ;
        RECT 58.800 430.300 59.600 430.400 ;
        RECT 60.400 430.300 61.200 430.400 ;
        RECT 58.800 430.200 61.200 430.300 ;
        RECT 54.600 429.700 61.200 430.200 ;
        RECT 54.600 429.600 59.600 429.700 ;
        RECT 60.400 429.600 61.200 429.700 ;
        RECT 54.600 429.400 55.400 429.600 ;
        RECT 56.200 428.400 57.000 428.600 ;
        RECT 63.600 428.400 64.200 431.600 ;
        RECT 70.000 431.200 70.800 439.800 ;
        RECT 66.600 430.600 70.800 431.200 ;
        RECT 71.600 435.000 72.400 439.000 ;
        RECT 71.600 431.600 72.200 435.000 ;
        RECT 75.800 432.800 76.600 439.800 ;
        RECT 75.800 432.200 77.400 432.800 ;
        RECT 71.600 431.000 75.400 431.600 ;
        RECT 66.600 430.400 67.400 430.600 ;
        RECT 68.200 429.800 69.000 430.000 ;
        RECT 65.200 429.200 69.000 429.800 ;
        RECT 65.200 429.000 66.000 429.200 ;
        RECT 53.200 427.800 64.200 428.400 ;
        RECT 53.200 427.600 54.800 427.800 ;
        RECT 33.200 422.200 34.000 424.200 ;
        RECT 36.400 422.200 37.200 426.200 ;
        RECT 39.600 426.800 41.400 427.600 ;
        RECT 42.800 426.800 45.000 427.600 ;
        RECT 46.000 426.800 48.200 427.600 ;
        RECT 49.200 426.800 51.600 427.600 ;
        RECT 39.600 422.200 40.400 426.800 ;
        RECT 42.800 422.200 43.600 426.800 ;
        RECT 46.000 422.200 46.800 426.800 ;
        RECT 49.200 422.200 50.000 426.800 ;
        RECT 52.400 422.200 53.200 427.000 ;
        RECT 57.400 426.400 58.000 427.800 ;
        RECT 63.000 427.600 63.800 427.800 ;
        RECT 70.000 427.200 70.800 430.600 ;
        RECT 71.600 428.800 72.400 430.400 ;
        RECT 73.200 428.800 74.000 430.400 ;
        RECT 74.800 429.000 75.400 431.000 ;
        RECT 74.800 428.200 76.200 429.000 ;
        RECT 76.800 428.400 77.400 432.200 ;
        RECT 83.800 432.400 84.600 439.800 ;
        RECT 85.200 433.600 86.000 434.400 ;
        RECT 85.400 432.400 86.000 433.600 ;
        RECT 88.400 433.600 89.200 434.400 ;
        RECT 88.400 432.400 89.000 433.600 ;
        RECT 89.800 432.400 90.600 439.800 ;
        RECT 83.800 431.800 84.800 432.400 ;
        RECT 85.400 431.800 86.800 432.400 ;
        RECT 78.000 429.600 78.800 431.200 ;
        RECT 84.200 430.400 84.800 431.800 ;
        RECT 86.000 431.600 86.800 431.800 ;
        RECT 87.600 431.800 89.000 432.400 ;
        RECT 89.600 431.800 90.600 432.400 ;
        RECT 87.600 431.600 88.400 431.800 ;
        RECT 82.800 430.300 83.600 430.400 ;
        RECT 79.700 429.700 83.600 430.300 ;
        RECT 76.800 428.300 78.800 428.400 ;
        RECT 79.700 428.300 80.300 429.700 ;
        RECT 82.800 428.800 83.600 429.700 ;
        RECT 84.200 429.600 85.200 430.400 ;
        RECT 86.100 430.300 86.700 431.600 ;
        RECT 89.600 430.300 90.200 431.800 ;
        RECT 86.100 429.700 90.200 430.300 ;
        RECT 84.200 428.400 84.800 429.600 ;
        RECT 89.600 428.400 90.200 429.700 ;
        RECT 90.800 428.800 91.600 430.400 ;
        RECT 74.800 427.800 75.800 428.200 ;
        RECT 67.000 426.600 70.800 427.200 ;
        RECT 67.000 426.400 67.800 426.600 ;
        RECT 55.600 424.200 56.400 425.000 ;
        RECT 57.200 424.800 58.000 426.400 ;
        RECT 59.000 425.400 59.800 425.600 ;
        RECT 59.000 424.800 61.800 425.400 ;
        RECT 61.200 424.200 61.800 424.800 ;
        RECT 65.200 424.200 66.000 425.000 ;
        RECT 55.600 423.600 57.600 424.200 ;
        RECT 56.800 422.200 57.600 423.600 ;
        RECT 61.200 422.200 62.000 424.200 ;
        RECT 65.200 423.600 66.600 424.200 ;
        RECT 65.400 422.200 66.600 423.600 ;
        RECT 70.000 422.200 70.800 426.600 ;
        RECT 71.600 427.200 75.800 427.800 ;
        RECT 76.800 427.700 80.300 428.300 ;
        RECT 81.200 428.200 82.000 428.400 ;
        RECT 76.800 427.600 78.800 427.700 ;
        RECT 81.200 427.600 82.800 428.200 ;
        RECT 84.200 427.600 86.800 428.400 ;
        RECT 87.600 427.600 90.200 428.400 ;
        RECT 92.400 428.200 93.200 428.400 ;
        RECT 91.600 427.600 93.200 428.200 ;
        RECT 71.600 425.000 72.200 427.200 ;
        RECT 76.800 427.000 77.400 427.600 ;
        RECT 82.000 427.200 82.800 427.600 ;
        RECT 76.600 426.600 77.400 427.000 ;
        RECT 75.800 426.000 77.400 426.600 ;
        RECT 81.400 426.200 85.000 426.600 ;
        RECT 86.000 426.200 86.600 427.600 ;
        RECT 87.800 426.200 88.400 427.600 ;
        RECT 91.600 427.200 92.400 427.600 ;
        RECT 94.000 426.800 94.800 428.400 ;
        RECT 89.400 426.200 93.000 426.600 ;
        RECT 95.600 426.200 96.400 439.800 ;
        RECT 98.800 435.000 99.600 439.000 ;
        RECT 97.200 431.600 98.000 433.200 ;
        RECT 98.800 431.600 99.400 435.000 ;
        RECT 103.000 432.800 103.800 439.800 ;
        RECT 103.000 432.200 104.600 432.800 ;
        RECT 98.800 431.000 102.600 431.600 ;
        RECT 98.800 428.800 99.600 430.400 ;
        RECT 100.400 428.800 101.200 430.400 ;
        RECT 102.000 429.000 102.600 431.000 ;
        RECT 102.000 428.200 103.400 429.000 ;
        RECT 104.000 428.400 104.600 432.200 ;
        RECT 111.000 432.400 111.800 439.800 ;
        RECT 112.400 433.600 113.200 434.400 ;
        RECT 112.600 432.400 113.200 433.600 ;
        RECT 115.600 433.600 116.400 434.400 ;
        RECT 115.600 432.400 116.200 433.600 ;
        RECT 117.000 432.400 117.800 439.800 ;
        RECT 111.000 431.800 112.000 432.400 ;
        RECT 112.600 431.800 114.000 432.400 ;
        RECT 105.200 430.300 106.000 431.200 ;
        RECT 106.800 430.300 107.600 430.400 ;
        RECT 105.200 429.700 107.600 430.300 ;
        RECT 105.200 429.600 106.000 429.700 ;
        RECT 106.800 429.600 107.600 429.700 ;
        RECT 110.000 428.800 110.800 430.400 ;
        RECT 111.400 428.400 112.000 431.800 ;
        RECT 113.200 431.600 114.000 431.800 ;
        RECT 114.800 431.800 116.200 432.400 ;
        RECT 116.800 431.800 117.800 432.400 ;
        RECT 114.800 431.600 115.600 431.800 ;
        RECT 113.300 430.300 113.900 431.600 ;
        RECT 116.800 430.300 117.400 431.800 ;
        RECT 113.300 429.700 117.400 430.300 ;
        RECT 116.800 428.400 117.400 429.700 ;
        RECT 118.000 428.800 118.800 430.400 ;
        RECT 104.000 428.300 106.000 428.400 ;
        RECT 106.800 428.300 107.600 428.400 ;
        RECT 102.000 427.800 103.000 428.200 ;
        RECT 98.800 427.200 103.000 427.800 ;
        RECT 104.000 427.700 107.600 428.300 ;
        RECT 104.000 427.600 106.000 427.700 ;
        RECT 106.800 427.600 107.600 427.700 ;
        RECT 108.400 428.200 109.200 428.400 ;
        RECT 108.400 427.600 110.000 428.200 ;
        RECT 111.400 427.600 114.000 428.400 ;
        RECT 114.800 427.600 117.400 428.400 ;
        RECT 119.600 428.200 120.400 428.400 ;
        RECT 118.800 427.600 120.400 428.200 ;
        RECT 122.800 428.300 123.600 439.800 ;
        RECT 127.000 432.400 127.800 439.800 ;
        RECT 128.400 433.600 129.200 434.400 ;
        RECT 128.600 432.400 129.200 433.600 ;
        RECT 127.000 431.800 128.000 432.400 ;
        RECT 128.600 431.800 130.000 432.400 ;
        RECT 126.000 428.800 126.800 430.400 ;
        RECT 127.400 428.400 128.000 431.800 ;
        RECT 129.200 431.600 130.000 431.800 ;
        RECT 124.400 428.300 125.200 428.400 ;
        RECT 122.800 428.200 125.200 428.300 ;
        RECT 122.800 427.700 126.000 428.200 ;
        RECT 81.200 426.000 85.200 426.200 ;
        RECT 71.600 423.000 72.400 425.000 ;
        RECT 75.800 423.000 76.600 426.000 ;
        RECT 81.200 422.200 82.000 426.000 ;
        RECT 84.400 422.200 85.200 426.000 ;
        RECT 86.000 422.200 86.800 426.200 ;
        RECT 87.600 422.200 88.400 426.200 ;
        RECT 89.200 426.000 93.200 426.200 ;
        RECT 89.200 422.200 90.000 426.000 ;
        RECT 92.400 422.200 93.200 426.000 ;
        RECT 95.600 425.600 97.400 426.200 ;
        RECT 96.600 424.400 97.400 425.600 ;
        RECT 95.600 423.600 97.400 424.400 ;
        RECT 96.600 422.200 97.400 423.600 ;
        RECT 98.800 425.000 99.400 427.200 ;
        RECT 104.000 427.000 104.600 427.600 ;
        RECT 109.200 427.200 110.000 427.600 ;
        RECT 103.800 426.600 104.600 427.000 ;
        RECT 103.000 426.000 104.600 426.600 ;
        RECT 108.600 426.200 112.200 426.600 ;
        RECT 113.200 426.200 113.800 427.600 ;
        RECT 115.000 426.200 115.600 427.600 ;
        RECT 118.800 427.200 119.600 427.600 ;
        RECT 116.600 426.200 120.200 426.600 ;
        RECT 108.400 426.000 112.400 426.200 ;
        RECT 98.800 423.000 99.600 425.000 ;
        RECT 103.000 423.000 103.800 426.000 ;
        RECT 108.400 422.200 109.200 426.000 ;
        RECT 111.600 422.200 112.400 426.000 ;
        RECT 113.200 422.200 114.000 426.200 ;
        RECT 114.800 422.200 115.600 426.200 ;
        RECT 116.400 426.000 120.400 426.200 ;
        RECT 116.400 422.200 117.200 426.000 ;
        RECT 119.600 422.200 120.400 426.000 ;
        RECT 121.200 424.800 122.000 426.400 ;
        RECT 122.800 422.200 123.600 427.700 ;
        RECT 124.400 427.600 126.000 427.700 ;
        RECT 127.400 427.600 130.000 428.400 ;
        RECT 125.200 427.200 126.000 427.600 ;
        RECT 124.600 426.200 128.200 426.600 ;
        RECT 129.200 426.200 129.800 427.600 ;
        RECT 124.400 426.000 128.400 426.200 ;
        RECT 124.400 422.200 125.200 426.000 ;
        RECT 127.600 422.200 128.400 426.000 ;
        RECT 129.200 422.200 130.000 426.200 ;
        RECT 130.800 424.800 131.600 426.400 ;
        RECT 132.400 422.200 133.200 439.800 ;
        RECT 134.000 431.200 134.800 439.800 ;
        RECT 138.200 435.800 139.400 439.800 ;
        RECT 142.800 435.800 143.600 439.800 ;
        RECT 147.200 436.400 148.000 439.800 ;
        RECT 147.200 435.800 149.200 436.400 ;
        RECT 138.800 435.000 139.600 435.800 ;
        RECT 143.000 435.200 143.600 435.800 ;
        RECT 142.200 434.600 145.800 435.200 ;
        RECT 148.400 435.000 149.200 435.800 ;
        RECT 142.200 434.400 143.000 434.600 ;
        RECT 145.000 434.400 145.800 434.600 ;
        RECT 138.000 433.200 139.400 434.000 ;
        RECT 138.800 432.200 139.400 433.200 ;
        RECT 141.000 433.000 143.200 433.600 ;
        RECT 141.000 432.800 141.800 433.000 ;
        RECT 138.800 431.600 141.200 432.200 ;
        RECT 134.000 430.600 138.200 431.200 ;
        RECT 134.000 427.200 134.800 430.600 ;
        RECT 137.400 430.400 138.200 430.600 ;
        RECT 135.800 429.800 136.600 430.000 ;
        RECT 135.800 429.200 139.600 429.800 ;
        RECT 138.800 429.000 139.600 429.200 ;
        RECT 140.600 428.400 141.200 431.600 ;
        RECT 142.600 431.800 143.200 433.000 ;
        RECT 143.800 433.000 144.600 433.200 ;
        RECT 148.400 433.000 149.200 433.200 ;
        RECT 143.800 432.400 149.200 433.000 ;
        RECT 142.600 431.400 147.400 431.800 ;
        RECT 151.600 431.400 152.400 439.800 ;
        RECT 160.600 432.400 161.400 439.800 ;
        RECT 166.600 434.400 167.400 439.800 ;
        RECT 162.000 433.600 162.800 434.400 ;
        RECT 162.200 432.400 162.800 433.600 ;
        RECT 165.200 433.600 166.000 434.400 ;
        RECT 166.600 433.600 168.400 434.400 ;
        RECT 165.200 432.400 165.800 433.600 ;
        RECT 166.600 432.400 167.400 433.600 ;
        RECT 160.600 431.800 161.600 432.400 ;
        RECT 162.200 431.800 163.600 432.400 ;
        RECT 142.600 431.200 152.400 431.400 ;
        RECT 146.600 431.000 152.400 431.200 ;
        RECT 146.800 430.800 152.400 431.000 ;
        RECT 145.200 430.200 146.000 430.400 ;
        RECT 156.400 430.300 157.200 430.400 ;
        RECT 159.600 430.300 160.400 430.400 ;
        RECT 145.200 429.600 150.200 430.200 ;
        RECT 156.400 429.700 160.400 430.300 ;
        RECT 156.400 429.600 157.200 429.700 ;
        RECT 149.400 429.400 150.200 429.600 ;
        RECT 159.600 428.800 160.400 429.700 ;
        RECT 161.000 430.300 161.600 431.800 ;
        RECT 162.800 431.600 163.600 431.800 ;
        RECT 164.400 431.800 165.800 432.400 ;
        RECT 166.400 431.800 167.400 432.400 ;
        RECT 173.400 432.400 174.200 439.800 ;
        RECT 179.400 438.400 180.200 439.800 ;
        RECT 179.400 437.600 181.200 438.400 ;
        RECT 174.800 433.600 175.600 434.400 ;
        RECT 175.000 432.400 175.600 433.600 ;
        RECT 178.000 433.600 178.800 434.400 ;
        RECT 178.000 432.400 178.600 433.600 ;
        RECT 179.400 432.400 180.200 437.600 ;
        RECT 173.400 431.800 174.400 432.400 ;
        RECT 175.000 431.800 176.400 432.400 ;
        RECT 164.400 431.600 165.200 431.800 ;
        RECT 164.500 430.300 165.100 431.600 ;
        RECT 161.000 429.700 165.100 430.300 ;
        RECT 147.800 428.400 148.600 428.600 ;
        RECT 161.000 428.400 161.600 429.700 ;
        RECT 166.400 428.400 167.000 431.800 ;
        RECT 167.600 428.800 168.400 430.400 ;
        RECT 172.400 428.800 173.200 430.400 ;
        RECT 173.800 430.300 174.400 431.800 ;
        RECT 175.600 431.600 176.400 431.800 ;
        RECT 177.200 431.800 178.600 432.400 ;
        RECT 179.200 431.800 180.200 432.400 ;
        RECT 177.200 431.600 178.000 431.800 ;
        RECT 177.300 430.300 177.900 431.600 ;
        RECT 173.800 429.700 177.900 430.300 ;
        RECT 173.800 428.400 174.400 429.700 ;
        RECT 179.200 428.400 179.800 431.800 ;
        RECT 183.600 431.200 184.400 439.800 ;
        RECT 187.800 435.800 189.000 439.800 ;
        RECT 192.400 435.800 193.200 439.800 ;
        RECT 196.800 436.400 197.600 439.800 ;
        RECT 196.800 435.800 198.800 436.400 ;
        RECT 188.400 435.000 189.200 435.800 ;
        RECT 192.600 435.200 193.200 435.800 ;
        RECT 191.800 434.600 195.400 435.200 ;
        RECT 198.000 435.000 198.800 435.800 ;
        RECT 191.800 434.400 192.600 434.600 ;
        RECT 194.600 434.400 195.400 434.600 ;
        RECT 187.600 433.200 189.000 434.000 ;
        RECT 188.400 432.200 189.000 433.200 ;
        RECT 190.600 433.000 192.800 433.600 ;
        RECT 190.600 432.800 191.400 433.000 ;
        RECT 188.400 431.600 190.800 432.200 ;
        RECT 183.600 430.600 187.800 431.200 ;
        RECT 180.400 428.800 181.200 430.400 ;
        RECT 140.600 427.800 151.600 428.400 ;
        RECT 141.000 427.600 141.800 427.800 ;
        RECT 134.000 426.600 137.800 427.200 ;
        RECT 134.000 422.200 134.800 426.600 ;
        RECT 137.000 426.400 137.800 426.600 ;
        RECT 146.800 425.600 147.400 427.800 ;
        RECT 150.000 427.600 151.600 427.800 ;
        RECT 158.000 428.200 158.800 428.400 ;
        RECT 158.000 427.600 159.600 428.200 ;
        RECT 161.000 427.600 163.600 428.400 ;
        RECT 164.400 427.600 167.000 428.400 ;
        RECT 169.200 428.200 170.000 428.400 ;
        RECT 168.400 427.600 170.000 428.200 ;
        RECT 170.800 428.200 171.600 428.400 ;
        RECT 170.800 427.600 172.400 428.200 ;
        RECT 173.800 427.600 176.400 428.400 ;
        RECT 177.200 427.600 179.800 428.400 ;
        RECT 182.000 428.200 182.800 428.400 ;
        RECT 181.200 427.600 182.800 428.200 ;
        RECT 158.800 427.200 159.600 427.600 ;
        RECT 145.000 425.400 145.800 425.600 ;
        RECT 138.800 424.200 139.600 425.000 ;
        RECT 143.000 424.800 145.800 425.400 ;
        RECT 146.800 424.800 147.600 425.600 ;
        RECT 143.000 424.200 143.600 424.800 ;
        RECT 148.400 424.200 149.200 425.000 ;
        RECT 138.200 423.600 139.600 424.200 ;
        RECT 138.200 422.200 139.400 423.600 ;
        RECT 142.800 422.200 143.600 424.200 ;
        RECT 147.200 423.600 149.200 424.200 ;
        RECT 147.200 422.200 148.000 423.600 ;
        RECT 151.600 422.200 152.400 427.000 ;
        RECT 158.200 426.200 161.800 426.600 ;
        RECT 162.800 426.200 163.400 427.600 ;
        RECT 164.600 426.200 165.200 427.600 ;
        RECT 168.400 427.200 169.200 427.600 ;
        RECT 171.600 427.200 172.400 427.600 ;
        RECT 166.200 426.200 169.800 426.600 ;
        RECT 171.000 426.200 174.600 426.600 ;
        RECT 175.600 426.200 176.200 427.600 ;
        RECT 177.400 426.200 178.000 427.600 ;
        RECT 181.200 427.200 182.000 427.600 ;
        RECT 183.600 427.200 184.400 430.600 ;
        RECT 187.000 430.400 187.800 430.600 ;
        RECT 185.400 429.800 186.200 430.000 ;
        RECT 185.400 429.200 189.200 429.800 ;
        RECT 188.400 429.000 189.200 429.200 ;
        RECT 190.200 428.400 190.800 431.600 ;
        RECT 192.200 431.800 192.800 433.000 ;
        RECT 193.400 433.000 194.200 433.200 ;
        RECT 198.000 433.000 198.800 433.200 ;
        RECT 193.400 432.400 198.800 433.000 ;
        RECT 192.200 431.400 197.000 431.800 ;
        RECT 201.200 431.400 202.000 439.800 ;
        RECT 205.400 432.400 206.200 439.800 ;
        RECT 206.800 433.600 207.600 434.400 ;
        RECT 207.000 432.400 207.600 433.600 ;
        RECT 211.800 432.400 212.600 439.800 ;
        RECT 213.200 433.600 214.000 434.400 ;
        RECT 213.400 432.400 214.000 433.600 ;
        RECT 205.400 431.800 206.400 432.400 ;
        RECT 207.000 431.800 208.400 432.400 ;
        RECT 211.800 431.800 212.800 432.400 ;
        RECT 213.400 431.800 214.800 432.400 ;
        RECT 192.200 431.200 202.000 431.400 ;
        RECT 196.200 431.000 202.000 431.200 ;
        RECT 196.400 430.800 202.000 431.000 ;
        RECT 194.800 430.200 195.600 430.400 ;
        RECT 194.800 429.600 199.800 430.200 ;
        RECT 199.000 429.400 199.800 429.600 ;
        RECT 204.400 428.800 205.200 430.400 ;
        RECT 197.400 428.400 198.200 428.600 ;
        RECT 205.800 428.400 206.400 431.800 ;
        RECT 207.600 431.600 208.400 431.800 ;
        RECT 210.800 428.800 211.600 430.400 ;
        RECT 212.200 428.400 212.800 431.800 ;
        RECT 214.000 431.600 214.800 431.800 ;
        RECT 215.600 431.600 216.400 433.200 ;
        RECT 190.200 427.800 201.200 428.400 ;
        RECT 190.600 427.600 191.400 427.800 ;
        RECT 193.200 427.600 194.000 427.800 ;
        RECT 183.600 426.600 187.400 427.200 ;
        RECT 179.000 426.200 182.600 426.600 ;
        RECT 158.000 426.000 162.000 426.200 ;
        RECT 158.000 422.200 158.800 426.000 ;
        RECT 161.200 422.200 162.000 426.000 ;
        RECT 162.800 422.200 163.600 426.200 ;
        RECT 164.400 422.200 165.200 426.200 ;
        RECT 166.000 426.000 170.000 426.200 ;
        RECT 166.000 422.200 166.800 426.000 ;
        RECT 169.200 422.200 170.000 426.000 ;
        RECT 170.800 426.000 174.800 426.200 ;
        RECT 170.800 422.200 171.600 426.000 ;
        RECT 174.000 422.200 174.800 426.000 ;
        RECT 175.600 422.200 176.400 426.200 ;
        RECT 177.200 422.200 178.000 426.200 ;
        RECT 178.800 426.000 182.800 426.200 ;
        RECT 178.800 422.200 179.600 426.000 ;
        RECT 182.000 422.200 182.800 426.000 ;
        RECT 183.600 422.200 184.400 426.600 ;
        RECT 186.600 426.400 187.400 426.600 ;
        RECT 196.400 425.600 197.000 427.800 ;
        RECT 199.600 427.600 201.200 427.800 ;
        RECT 202.800 428.200 203.600 428.400 ;
        RECT 205.800 428.300 208.400 428.400 ;
        RECT 209.200 428.300 210.000 428.400 ;
        RECT 205.800 428.200 210.000 428.300 ;
        RECT 202.800 427.600 204.400 428.200 ;
        RECT 205.800 427.700 210.800 428.200 ;
        RECT 205.800 427.600 208.400 427.700 ;
        RECT 209.200 427.600 210.800 427.700 ;
        RECT 212.200 427.600 214.800 428.400 ;
        RECT 203.600 427.200 204.400 427.600 ;
        RECT 194.600 425.400 195.400 425.600 ;
        RECT 188.400 424.200 189.200 425.000 ;
        RECT 192.600 424.800 195.400 425.400 ;
        RECT 196.400 424.800 197.200 425.600 ;
        RECT 192.600 424.200 193.200 424.800 ;
        RECT 198.000 424.200 198.800 425.000 ;
        RECT 187.800 423.600 189.200 424.200 ;
        RECT 187.800 422.200 189.000 423.600 ;
        RECT 192.400 422.200 193.200 424.200 ;
        RECT 196.800 423.600 198.800 424.200 ;
        RECT 196.800 422.200 197.600 423.600 ;
        RECT 201.200 422.200 202.000 427.000 ;
        RECT 203.000 426.200 206.600 426.600 ;
        RECT 207.600 426.200 208.200 427.600 ;
        RECT 210.000 427.200 210.800 427.600 ;
        RECT 209.400 426.200 213.000 426.600 ;
        RECT 214.000 426.200 214.600 427.600 ;
        RECT 217.200 426.200 218.000 439.800 ;
        RECT 221.200 433.600 222.000 434.400 ;
        RECT 221.200 432.400 221.800 433.600 ;
        RECT 222.600 432.400 223.400 439.800 ;
        RECT 220.400 431.800 221.800 432.400 ;
        RECT 222.400 431.800 223.400 432.400 ;
        RECT 226.800 431.800 227.600 439.800 ;
        RECT 230.000 435.800 230.800 439.800 ;
        RECT 220.400 431.600 221.200 431.800 ;
        RECT 218.800 430.300 219.600 430.400 ;
        RECT 222.400 430.300 223.000 431.800 ;
        RECT 226.800 430.400 227.400 431.800 ;
        RECT 230.000 431.600 230.600 435.800 ;
        RECT 228.200 431.000 230.600 431.600 ;
        RECT 218.800 429.700 223.000 430.300 ;
        RECT 218.800 429.600 219.600 429.700 ;
        RECT 222.400 428.400 223.000 429.700 ;
        RECT 223.600 428.800 224.400 430.400 ;
        RECT 226.800 430.300 227.600 430.400 ;
        RECT 225.300 429.700 227.600 430.300 ;
        RECT 225.300 428.400 225.900 429.700 ;
        RECT 226.800 429.600 227.600 429.700 ;
        RECT 218.800 426.800 219.600 428.400 ;
        RECT 220.400 427.600 223.000 428.400 ;
        RECT 225.200 428.200 226.000 428.400 ;
        RECT 224.400 427.600 226.000 428.200 ;
        RECT 220.600 426.200 221.200 427.600 ;
        RECT 224.400 427.200 225.200 427.600 ;
        RECT 222.200 426.200 225.800 426.600 ;
        RECT 226.800 426.200 227.400 429.600 ;
        RECT 228.200 427.600 228.800 431.000 ;
        RECT 230.000 429.600 230.800 430.400 ;
        RECT 230.000 428.800 230.600 429.600 ;
        RECT 229.600 428.200 230.600 428.800 ;
        RECT 229.600 428.000 230.400 428.200 ;
        RECT 231.600 427.600 232.400 429.200 ;
        RECT 228.000 427.400 228.800 427.600 ;
        RECT 228.000 427.000 231.000 427.400 ;
        RECT 228.000 426.800 232.200 427.000 ;
        RECT 233.200 426.800 234.000 428.400 ;
        RECT 230.400 426.400 232.200 426.800 ;
        RECT 231.600 426.200 232.200 426.400 ;
        RECT 234.800 426.200 235.600 439.800 ;
        RECT 236.400 432.300 237.200 433.200 ;
        RECT 239.600 432.300 240.400 439.800 ;
        RECT 243.600 433.600 244.400 434.400 ;
        RECT 236.400 431.700 240.400 432.300 ;
        RECT 236.400 431.600 237.200 431.700 ;
        RECT 238.000 426.800 238.800 428.400 ;
        RECT 239.600 426.200 240.400 431.700 ;
        RECT 241.200 431.600 242.000 433.200 ;
        RECT 243.600 432.400 244.200 433.600 ;
        RECT 245.000 432.400 245.800 439.800 ;
        RECT 242.800 431.800 244.200 432.400 ;
        RECT 244.800 431.800 245.800 432.400 ;
        RECT 242.800 431.600 243.600 431.800 ;
        RECT 242.800 430.300 243.600 430.400 ;
        RECT 244.800 430.300 245.400 431.800 ;
        RECT 242.800 429.700 245.400 430.300 ;
        RECT 242.800 429.600 243.600 429.700 ;
        RECT 244.800 428.400 245.400 429.700 ;
        RECT 246.000 428.800 246.800 430.400 ;
        RECT 242.800 427.600 245.400 428.400 ;
        RECT 247.600 428.300 248.400 428.400 ;
        RECT 249.200 428.300 250.000 439.800 ;
        RECT 253.200 433.600 254.000 434.400 ;
        RECT 253.200 432.400 253.800 433.600 ;
        RECT 254.600 432.400 255.400 439.800 ;
        RECT 252.400 431.800 253.800 432.400 ;
        RECT 254.400 431.800 255.400 432.400 ;
        RECT 258.800 435.000 259.600 439.000 ;
        RECT 252.400 431.600 253.200 431.800 ;
        RECT 254.400 428.400 255.000 431.800 ;
        RECT 258.800 431.600 259.400 435.000 ;
        RECT 263.000 432.800 263.800 439.800 ;
        RECT 268.400 435.000 269.200 439.000 ;
        RECT 272.600 438.400 273.400 439.800 ;
        RECT 272.600 437.600 274.000 438.400 ;
        RECT 263.000 432.200 264.600 432.800 ;
        RECT 258.800 431.000 262.600 431.600 ;
        RECT 255.600 428.800 256.400 430.400 ;
        RECT 258.800 428.800 259.600 430.400 ;
        RECT 260.400 428.800 261.200 430.400 ;
        RECT 262.000 429.000 262.600 431.000 ;
        RECT 247.600 428.200 250.000 428.300 ;
        RECT 246.800 427.700 250.000 428.200 ;
        RECT 246.800 427.600 248.400 427.700 ;
        RECT 243.000 426.200 243.600 427.600 ;
        RECT 246.800 427.200 247.600 427.600 ;
        RECT 244.600 426.200 248.200 426.600 ;
        RECT 202.800 426.000 206.800 426.200 ;
        RECT 202.800 422.200 203.600 426.000 ;
        RECT 206.000 422.200 206.800 426.000 ;
        RECT 207.600 422.200 208.400 426.200 ;
        RECT 209.200 426.000 213.200 426.200 ;
        RECT 209.200 422.200 210.000 426.000 ;
        RECT 212.400 422.200 213.200 426.000 ;
        RECT 214.000 422.200 214.800 426.200 ;
        RECT 216.200 425.600 218.000 426.200 ;
        RECT 216.200 424.400 217.000 425.600 ;
        RECT 215.600 423.600 217.000 424.400 ;
        RECT 216.200 422.200 217.000 423.600 ;
        RECT 220.400 422.200 221.200 426.200 ;
        RECT 222.000 426.000 226.000 426.200 ;
        RECT 222.000 422.200 222.800 426.000 ;
        RECT 225.200 422.200 226.000 426.000 ;
        RECT 226.800 425.200 228.200 426.200 ;
        RECT 227.400 422.200 228.200 425.200 ;
        RECT 231.600 422.200 232.400 426.200 ;
        RECT 234.800 425.600 236.600 426.200 ;
        RECT 239.600 425.600 241.400 426.200 ;
        RECT 235.800 424.400 236.600 425.600 ;
        RECT 234.800 423.600 236.600 424.400 ;
        RECT 235.800 422.200 236.600 423.600 ;
        RECT 240.600 422.200 241.400 425.600 ;
        RECT 242.800 422.200 243.600 426.200 ;
        RECT 244.400 426.000 248.400 426.200 ;
        RECT 244.400 422.200 245.200 426.000 ;
        RECT 247.600 422.200 248.400 426.000 ;
        RECT 249.200 422.200 250.000 427.700 ;
        RECT 252.400 427.600 255.000 428.400 ;
        RECT 257.200 428.200 258.000 428.400 ;
        RECT 256.400 427.600 258.000 428.200 ;
        RECT 262.000 428.200 263.400 429.000 ;
        RECT 264.000 428.400 264.600 432.200 ;
        RECT 268.400 431.600 269.000 435.000 ;
        RECT 272.600 432.800 273.400 437.600 ;
        RECT 272.600 432.200 274.200 432.800 ;
        RECT 265.200 430.300 266.000 431.200 ;
        RECT 268.400 431.000 272.200 431.600 ;
        RECT 266.800 430.300 267.600 430.400 ;
        RECT 265.200 429.700 267.600 430.300 ;
        RECT 265.200 429.600 266.000 429.700 ;
        RECT 266.800 429.600 267.600 429.700 ;
        RECT 268.400 428.800 269.200 430.400 ;
        RECT 270.000 428.800 270.800 430.400 ;
        RECT 271.600 429.000 272.200 431.000 ;
        RECT 262.000 427.800 263.000 428.200 ;
        RECT 250.800 426.300 251.600 426.400 ;
        RECT 252.600 426.300 253.200 427.600 ;
        RECT 256.400 427.200 257.200 427.600 ;
        RECT 258.800 427.200 263.000 427.800 ;
        RECT 264.000 427.600 266.000 428.400 ;
        RECT 271.600 428.200 273.000 429.000 ;
        RECT 273.600 428.400 274.200 432.200 ;
        RECT 278.000 431.600 278.800 433.200 ;
        RECT 274.800 429.600 275.600 431.200 ;
        RECT 271.600 427.800 272.600 428.200 ;
        RECT 250.800 425.700 253.200 426.300 ;
        RECT 254.200 426.200 257.800 426.600 ;
        RECT 250.800 424.800 251.600 425.700 ;
        RECT 252.400 422.200 253.200 425.700 ;
        RECT 254.000 426.000 258.000 426.200 ;
        RECT 254.000 422.200 254.800 426.000 ;
        RECT 257.200 422.200 258.000 426.000 ;
        RECT 258.800 425.000 259.400 427.200 ;
        RECT 264.000 427.000 264.600 427.600 ;
        RECT 263.800 426.600 264.600 427.000 ;
        RECT 263.000 426.000 264.600 426.600 ;
        RECT 268.400 427.200 272.600 427.800 ;
        RECT 273.600 427.600 275.600 428.400 ;
        RECT 258.800 423.000 259.600 425.000 ;
        RECT 263.000 423.000 263.800 426.000 ;
        RECT 268.400 425.000 269.000 427.200 ;
        RECT 273.600 427.000 274.200 427.600 ;
        RECT 273.400 426.600 274.200 427.000 ;
        RECT 272.600 426.000 274.200 426.600 ;
        RECT 279.600 426.200 280.400 439.800 ;
        RECT 281.200 426.800 282.000 428.400 ;
        RECT 268.400 423.000 269.200 425.000 ;
        RECT 272.600 423.000 273.400 426.000 ;
        RECT 278.600 425.600 280.400 426.200 ;
        RECT 278.600 424.400 279.400 425.600 ;
        RECT 282.800 424.800 283.600 426.400 ;
        RECT 278.600 423.600 280.400 424.400 ;
        RECT 278.600 422.200 279.400 423.600 ;
        RECT 284.400 422.200 285.200 439.800 ;
        RECT 287.600 432.000 288.400 439.800 ;
        RECT 290.800 435.200 291.600 439.800 ;
        RECT 287.400 431.200 288.400 432.000 ;
        RECT 289.000 434.600 291.600 435.200 ;
        RECT 289.000 433.000 289.600 434.600 ;
        RECT 294.000 434.400 294.800 439.800 ;
        RECT 297.200 437.000 298.000 439.800 ;
        RECT 298.800 437.000 299.600 439.800 ;
        RECT 300.400 437.000 301.200 439.800 ;
        RECT 295.400 434.400 299.600 435.200 ;
        RECT 292.200 433.600 294.800 434.400 ;
        RECT 302.000 433.600 302.800 439.800 ;
        RECT 305.200 435.000 306.000 439.800 ;
        RECT 308.400 435.000 309.200 439.800 ;
        RECT 310.000 437.000 310.800 439.800 ;
        RECT 311.600 437.000 312.400 439.800 ;
        RECT 314.800 435.200 315.600 439.800 ;
        RECT 318.000 436.400 318.800 439.800 ;
        RECT 318.000 435.800 319.000 436.400 ;
        RECT 318.400 435.200 319.000 435.800 ;
        RECT 313.600 434.400 317.800 435.200 ;
        RECT 318.400 434.600 320.400 435.200 ;
        RECT 305.200 433.600 307.800 434.400 ;
        RECT 308.400 433.800 314.200 434.400 ;
        RECT 317.200 434.000 317.800 434.400 ;
        RECT 297.200 433.000 298.000 433.200 ;
        RECT 289.000 432.400 298.000 433.000 ;
        RECT 300.400 433.000 301.200 433.200 ;
        RECT 308.400 433.000 309.000 433.800 ;
        RECT 314.800 433.200 316.200 433.800 ;
        RECT 317.200 433.200 318.800 434.000 ;
        RECT 300.400 432.400 309.000 433.000 ;
        RECT 310.000 433.000 316.200 433.200 ;
        RECT 310.000 432.600 315.400 433.000 ;
        RECT 310.000 432.400 310.800 432.600 ;
        RECT 287.400 426.800 288.200 431.200 ;
        RECT 289.000 430.600 289.600 432.400 ;
        RECT 288.800 430.000 289.600 430.600 ;
        RECT 295.600 430.000 319.000 430.600 ;
        RECT 288.800 428.000 289.400 430.000 ;
        RECT 295.600 429.400 296.400 430.000 ;
        RECT 313.200 429.600 314.000 430.000 ;
        RECT 318.200 429.800 319.000 430.000 ;
        RECT 290.000 428.600 293.800 429.400 ;
        RECT 288.800 427.400 290.000 428.000 ;
        RECT 287.400 426.000 288.400 426.800 ;
        RECT 287.600 422.200 288.400 426.000 ;
        RECT 289.200 422.200 290.000 427.400 ;
        RECT 293.000 427.400 293.800 428.600 ;
        RECT 293.000 426.800 294.800 427.400 ;
        RECT 294.000 426.200 294.800 426.800 ;
        RECT 298.800 426.400 299.600 429.200 ;
        RECT 302.000 428.600 305.200 429.400 ;
        RECT 309.000 428.600 311.000 429.400 ;
        RECT 319.600 429.000 320.400 434.600 ;
        RECT 301.600 427.800 302.400 428.000 ;
        RECT 301.600 427.200 306.000 427.800 ;
        RECT 305.200 427.000 306.000 427.200 ;
        RECT 306.800 426.800 307.600 428.400 ;
        RECT 294.000 425.400 296.400 426.200 ;
        RECT 298.800 425.600 299.800 426.400 ;
        RECT 302.800 425.600 304.400 426.400 ;
        RECT 305.200 426.200 306.000 426.400 ;
        RECT 309.000 426.200 309.800 428.600 ;
        RECT 311.600 428.200 320.400 429.000 ;
        RECT 315.000 426.800 318.000 427.600 ;
        RECT 315.000 426.200 315.800 426.800 ;
        RECT 305.200 425.600 309.800 426.200 ;
        RECT 295.600 422.200 296.400 425.400 ;
        RECT 313.200 425.400 315.800 426.200 ;
        RECT 297.200 422.200 298.000 425.000 ;
        RECT 298.800 422.200 299.600 425.000 ;
        RECT 300.400 422.200 301.200 425.000 ;
        RECT 302.000 422.200 302.800 425.000 ;
        RECT 305.200 422.200 306.000 425.000 ;
        RECT 308.400 422.200 309.200 425.000 ;
        RECT 310.000 422.200 310.800 425.000 ;
        RECT 311.600 422.200 312.400 425.000 ;
        RECT 313.200 422.200 314.000 425.400 ;
        RECT 319.600 422.200 320.400 428.200 ;
        RECT 326.000 424.800 326.800 426.400 ;
        RECT 327.600 422.200 328.400 439.800 ;
        RECT 329.200 431.400 330.000 439.800 ;
        RECT 333.600 436.400 334.400 439.800 ;
        RECT 332.400 435.800 334.400 436.400 ;
        RECT 338.000 435.800 338.800 439.800 ;
        RECT 342.200 435.800 343.400 439.800 ;
        RECT 332.400 435.000 333.200 435.800 ;
        RECT 338.000 435.200 338.600 435.800 ;
        RECT 335.800 434.600 339.400 435.200 ;
        RECT 342.000 435.000 342.800 435.800 ;
        RECT 335.800 434.400 336.600 434.600 ;
        RECT 338.600 434.400 339.400 434.600 ;
        RECT 332.400 433.000 333.200 433.200 ;
        RECT 337.000 433.000 337.800 433.200 ;
        RECT 332.400 432.400 337.800 433.000 ;
        RECT 338.400 433.000 340.600 433.600 ;
        RECT 338.400 431.800 339.000 433.000 ;
        RECT 339.800 432.800 340.600 433.000 ;
        RECT 342.200 433.200 343.600 434.000 ;
        RECT 342.200 432.200 342.800 433.200 ;
        RECT 334.200 431.400 339.000 431.800 ;
        RECT 329.200 431.200 339.000 431.400 ;
        RECT 340.400 431.600 342.800 432.200 ;
        RECT 329.200 431.000 335.000 431.200 ;
        RECT 329.200 430.800 334.800 431.000 ;
        RECT 335.600 430.200 336.400 430.400 ;
        RECT 331.400 429.600 336.400 430.200 ;
        RECT 331.400 429.400 332.200 429.600 ;
        RECT 333.000 428.400 333.800 428.600 ;
        RECT 340.400 428.400 341.000 431.600 ;
        RECT 346.800 431.200 347.600 439.800 ;
        RECT 343.400 430.600 347.600 431.200 ;
        RECT 348.400 435.000 349.200 439.000 ;
        RECT 348.400 431.600 349.000 435.000 ;
        RECT 352.600 432.800 353.400 439.800 ;
        RECT 352.600 432.200 354.200 432.800 ;
        RECT 348.400 431.000 352.200 431.600 ;
        RECT 343.400 430.400 344.200 430.600 ;
        RECT 345.000 429.800 345.800 430.000 ;
        RECT 342.000 429.200 345.800 429.800 ;
        RECT 342.000 429.000 342.800 429.200 ;
        RECT 330.000 427.800 341.000 428.400 ;
        RECT 330.000 427.600 331.600 427.800 ;
        RECT 329.200 422.200 330.000 427.000 ;
        RECT 334.200 425.600 334.800 427.800 ;
        RECT 337.200 427.600 338.000 427.800 ;
        RECT 339.800 427.600 340.600 427.800 ;
        RECT 346.800 427.200 347.600 430.600 ;
        RECT 348.400 428.800 349.200 430.400 ;
        RECT 350.000 428.800 350.800 430.400 ;
        RECT 351.600 429.000 352.200 431.000 ;
        RECT 351.600 428.200 353.000 429.000 ;
        RECT 353.600 428.400 354.200 432.200 ;
        RECT 360.600 432.400 361.400 439.800 ;
        RECT 362.000 433.600 362.800 434.400 ;
        RECT 362.200 432.400 362.800 433.600 ;
        RECT 365.200 433.600 366.000 434.400 ;
        RECT 365.200 432.400 365.800 433.600 ;
        RECT 366.600 432.400 367.400 439.800 ;
        RECT 374.600 432.800 375.400 439.800 ;
        RECT 378.800 435.000 379.600 439.000 ;
        RECT 383.000 438.400 383.800 439.800 ;
        RECT 382.000 437.600 383.800 438.400 ;
        RECT 360.600 431.800 361.600 432.400 ;
        RECT 362.200 431.800 363.600 432.400 ;
        RECT 354.800 429.600 355.600 431.200 ;
        RECT 361.000 430.400 361.600 431.800 ;
        RECT 362.800 431.600 363.600 431.800 ;
        RECT 364.400 431.800 365.800 432.400 ;
        RECT 366.400 431.800 367.400 432.400 ;
        RECT 373.800 432.200 375.400 432.800 ;
        RECT 364.400 431.600 365.200 431.800 ;
        RECT 359.600 430.300 360.400 430.400 ;
        RECT 356.500 429.700 360.400 430.300 ;
        RECT 353.600 428.300 355.600 428.400 ;
        RECT 356.500 428.300 357.100 429.700 ;
        RECT 359.600 428.800 360.400 429.700 ;
        RECT 361.000 429.600 362.000 430.400 ;
        RECT 362.900 430.300 363.500 431.600 ;
        RECT 366.400 430.300 367.000 431.800 ;
        RECT 362.900 429.700 367.000 430.300 ;
        RECT 361.000 428.400 361.600 429.600 ;
        RECT 366.400 428.400 367.000 429.700 ;
        RECT 367.600 428.800 368.400 430.400 ;
        RECT 372.400 429.600 373.200 431.200 ;
        RECT 373.800 428.400 374.400 432.200 ;
        RECT 379.000 431.600 379.600 435.000 ;
        RECT 383.000 432.400 383.800 437.600 ;
        RECT 384.400 433.600 385.200 434.400 ;
        RECT 384.600 432.400 385.200 433.600 ;
        RECT 390.600 432.800 391.400 439.800 ;
        RECT 394.800 435.000 395.600 439.000 ;
        RECT 383.000 431.800 384.000 432.400 ;
        RECT 384.600 431.800 386.000 432.400 ;
        RECT 375.800 431.000 379.600 431.600 ;
        RECT 375.800 429.000 376.400 431.000 ;
        RECT 351.600 427.800 352.600 428.200 ;
        RECT 343.800 426.600 347.600 427.200 ;
        RECT 343.800 426.400 344.600 426.600 ;
        RECT 332.400 424.200 333.200 425.000 ;
        RECT 334.000 424.800 334.800 425.600 ;
        RECT 335.800 425.400 336.600 425.600 ;
        RECT 335.800 424.800 338.600 425.400 ;
        RECT 338.000 424.200 338.600 424.800 ;
        RECT 342.000 424.200 342.800 425.000 ;
        RECT 332.400 423.600 334.400 424.200 ;
        RECT 333.600 422.200 334.400 423.600 ;
        RECT 338.000 422.200 338.800 424.200 ;
        RECT 342.000 423.600 343.400 424.200 ;
        RECT 342.200 422.200 343.400 423.600 ;
        RECT 346.800 422.200 347.600 426.600 ;
        RECT 348.400 427.200 352.600 427.800 ;
        RECT 353.600 427.700 357.100 428.300 ;
        RECT 358.000 428.200 358.800 428.400 ;
        RECT 353.600 427.600 355.600 427.700 ;
        RECT 358.000 427.600 359.600 428.200 ;
        RECT 361.000 427.600 363.600 428.400 ;
        RECT 364.400 427.600 367.000 428.400 ;
        RECT 369.200 428.200 370.000 428.400 ;
        RECT 368.400 427.600 370.000 428.200 ;
        RECT 372.400 427.600 374.400 428.400 ;
        RECT 375.000 428.200 376.400 429.000 ;
        RECT 377.200 428.800 378.000 430.400 ;
        RECT 378.800 428.800 379.600 430.400 ;
        RECT 382.000 428.800 382.800 430.400 ;
        RECT 383.400 428.400 384.000 431.800 ;
        RECT 385.200 431.600 386.000 431.800 ;
        RECT 389.800 432.200 391.400 432.800 ;
        RECT 385.200 430.300 386.000 430.400 ;
        RECT 388.400 430.300 389.200 431.200 ;
        RECT 385.200 429.700 389.200 430.300 ;
        RECT 385.200 429.600 386.000 429.700 ;
        RECT 388.400 429.600 389.200 429.700 ;
        RECT 389.800 428.400 390.400 432.200 ;
        RECT 395.000 431.600 395.600 435.000 ;
        RECT 391.800 431.000 395.600 431.600 ;
        RECT 391.800 429.000 392.400 431.000 ;
        RECT 348.400 425.000 349.000 427.200 ;
        RECT 353.600 427.000 354.200 427.600 ;
        RECT 358.800 427.200 359.600 427.600 ;
        RECT 353.400 426.600 354.200 427.000 ;
        RECT 352.600 426.000 354.200 426.600 ;
        RECT 358.200 426.200 361.800 426.600 ;
        RECT 362.800 426.200 363.400 427.600 ;
        RECT 364.600 426.200 365.200 427.600 ;
        RECT 368.400 427.200 369.200 427.600 ;
        RECT 373.800 427.000 374.400 427.600 ;
        RECT 375.400 427.800 376.400 428.200 ;
        RECT 380.400 428.200 381.200 428.400 ;
        RECT 375.400 427.200 379.600 427.800 ;
        RECT 380.400 427.600 382.000 428.200 ;
        RECT 383.400 427.600 386.000 428.400 ;
        RECT 388.400 427.600 390.400 428.400 ;
        RECT 391.000 428.200 392.400 429.000 ;
        RECT 393.200 428.800 394.000 430.400 ;
        RECT 394.800 430.300 395.600 430.400 ;
        RECT 396.400 430.300 397.200 430.400 ;
        RECT 394.800 429.700 397.200 430.300 ;
        RECT 394.800 428.800 395.600 429.700 ;
        RECT 396.400 429.600 397.200 429.700 ;
        RECT 381.200 427.200 382.000 427.600 ;
        RECT 373.800 426.600 374.600 427.000 ;
        RECT 366.200 426.200 369.800 426.600 ;
        RECT 358.000 426.000 362.000 426.200 ;
        RECT 348.400 423.000 349.200 425.000 ;
        RECT 352.600 423.000 353.400 426.000 ;
        RECT 358.000 422.200 358.800 426.000 ;
        RECT 361.200 422.200 362.000 426.000 ;
        RECT 362.800 422.200 363.600 426.200 ;
        RECT 364.400 422.200 365.200 426.200 ;
        RECT 366.000 426.000 370.000 426.200 ;
        RECT 373.800 426.000 375.400 426.600 ;
        RECT 366.000 422.200 366.800 426.000 ;
        RECT 369.200 422.200 370.000 426.000 ;
        RECT 374.600 424.400 375.400 426.000 ;
        RECT 379.000 425.000 379.600 427.200 ;
        RECT 380.600 426.200 384.200 426.600 ;
        RECT 385.200 426.200 385.800 427.600 ;
        RECT 389.800 427.000 390.400 427.600 ;
        RECT 391.400 427.800 392.400 428.200 ;
        RECT 391.400 427.200 395.600 427.800 ;
        RECT 389.800 426.600 390.600 427.000 ;
        RECT 374.000 423.600 375.400 424.400 ;
        RECT 374.600 423.000 375.400 423.600 ;
        RECT 378.800 423.000 379.600 425.000 ;
        RECT 380.400 426.000 384.400 426.200 ;
        RECT 380.400 422.200 381.200 426.000 ;
        RECT 383.600 422.200 384.400 426.000 ;
        RECT 385.200 422.200 386.000 426.200 ;
        RECT 389.800 426.000 391.400 426.600 ;
        RECT 390.600 424.400 391.400 426.000 ;
        RECT 395.000 425.000 395.600 427.200 ;
        RECT 390.000 423.600 391.400 424.400 ;
        RECT 390.600 423.000 391.400 423.600 ;
        RECT 394.800 423.000 395.600 425.000 ;
        RECT 396.400 424.800 397.200 426.400 ;
        RECT 398.000 422.200 398.800 439.800 ;
        RECT 403.400 432.800 404.200 439.800 ;
        RECT 407.600 435.000 408.400 439.000 ;
        RECT 402.600 432.200 404.200 432.800 ;
        RECT 401.200 429.600 402.000 431.200 ;
        RECT 402.600 430.400 403.200 432.200 ;
        RECT 407.800 431.600 408.400 435.000 ;
        RECT 411.800 432.400 412.600 439.800 ;
        RECT 413.200 433.600 414.000 434.400 ;
        RECT 413.400 432.400 414.000 433.600 ;
        RECT 411.800 431.800 412.800 432.400 ;
        RECT 413.400 431.800 414.800 432.400 ;
        RECT 404.600 431.000 408.400 431.600 ;
        RECT 402.600 429.600 403.600 430.400 ;
        RECT 402.600 428.400 403.200 429.600 ;
        RECT 404.600 429.000 405.200 431.000 ;
        RECT 401.200 427.600 403.200 428.400 ;
        RECT 403.800 428.200 405.200 429.000 ;
        RECT 406.000 428.800 406.800 430.400 ;
        RECT 407.600 428.800 408.400 430.400 ;
        RECT 410.800 428.800 411.600 430.400 ;
        RECT 412.200 430.300 412.800 431.800 ;
        RECT 414.000 431.600 414.800 431.800 ;
        RECT 415.600 431.200 416.400 439.800 ;
        RECT 419.800 435.800 421.000 439.800 ;
        RECT 424.400 435.800 425.200 439.800 ;
        RECT 428.800 436.400 429.600 439.800 ;
        RECT 428.800 435.800 430.800 436.400 ;
        RECT 420.400 435.000 421.200 435.800 ;
        RECT 424.600 435.200 425.200 435.800 ;
        RECT 423.800 434.600 427.400 435.200 ;
        RECT 430.000 435.000 430.800 435.800 ;
        RECT 423.800 434.400 424.600 434.600 ;
        RECT 426.600 434.400 427.400 434.600 ;
        RECT 419.600 433.200 421.000 434.000 ;
        RECT 420.400 432.200 421.000 433.200 ;
        RECT 422.600 433.000 424.800 433.600 ;
        RECT 422.600 432.800 423.400 433.000 ;
        RECT 420.400 431.600 422.800 432.200 ;
        RECT 415.600 430.600 419.800 431.200 ;
        RECT 414.000 430.300 414.800 430.400 ;
        RECT 412.200 429.700 414.800 430.300 ;
        RECT 412.200 428.400 412.800 429.700 ;
        RECT 414.000 429.600 414.800 429.700 ;
        RECT 402.600 427.000 403.200 427.600 ;
        RECT 404.200 427.800 405.200 428.200 ;
        RECT 409.200 428.200 410.000 428.400 ;
        RECT 404.200 427.200 408.400 427.800 ;
        RECT 409.200 427.600 410.800 428.200 ;
        RECT 412.200 427.600 414.800 428.400 ;
        RECT 410.000 427.200 410.800 427.600 ;
        RECT 402.600 426.600 403.400 427.000 ;
        RECT 402.600 426.000 404.200 426.600 ;
        RECT 403.400 423.000 404.200 426.000 ;
        RECT 407.800 425.000 408.400 427.200 ;
        RECT 409.400 426.200 413.000 426.600 ;
        RECT 414.000 426.200 414.600 427.600 ;
        RECT 415.600 427.200 416.400 430.600 ;
        RECT 419.000 430.400 419.800 430.600 ;
        RECT 417.400 429.800 418.200 430.000 ;
        RECT 417.400 429.200 421.200 429.800 ;
        RECT 420.400 429.000 421.200 429.200 ;
        RECT 422.200 428.400 422.800 431.600 ;
        RECT 424.200 431.800 424.800 433.000 ;
        RECT 425.400 433.000 426.200 433.200 ;
        RECT 430.000 433.000 430.800 433.200 ;
        RECT 425.400 432.400 430.800 433.000 ;
        RECT 424.200 431.400 429.000 431.800 ;
        RECT 433.200 431.400 434.000 439.800 ;
        RECT 424.200 431.200 434.000 431.400 ;
        RECT 428.200 431.000 434.000 431.200 ;
        RECT 428.400 430.800 434.000 431.000 ;
        RECT 425.200 430.300 426.000 430.400 ;
        RECT 426.800 430.300 427.600 430.400 ;
        RECT 425.200 430.200 427.600 430.300 ;
        RECT 425.200 429.700 431.800 430.200 ;
        RECT 425.200 429.600 426.000 429.700 ;
        RECT 426.800 429.600 431.800 429.700 ;
        RECT 431.000 429.400 431.800 429.600 ;
        RECT 429.400 428.400 430.200 428.600 ;
        RECT 422.200 427.800 433.200 428.400 ;
        RECT 422.600 427.600 423.400 427.800 ;
        RECT 425.200 427.600 426.000 427.800 ;
        RECT 415.600 426.600 419.400 427.200 ;
        RECT 407.600 423.000 408.400 425.000 ;
        RECT 409.200 426.000 413.200 426.200 ;
        RECT 409.200 422.200 410.000 426.000 ;
        RECT 412.400 422.200 413.200 426.000 ;
        RECT 414.000 422.200 414.800 426.200 ;
        RECT 415.600 422.200 416.400 426.600 ;
        RECT 418.600 426.400 419.400 426.600 ;
        RECT 428.400 425.600 429.000 427.800 ;
        RECT 431.600 427.600 433.200 427.800 ;
        RECT 436.400 428.300 437.200 439.800 ;
        RECT 440.600 432.400 441.400 439.800 ;
        RECT 442.000 433.600 442.800 434.400 ;
        RECT 442.200 432.400 442.800 433.600 ;
        RECT 440.600 431.800 441.600 432.400 ;
        RECT 442.200 431.800 443.600 432.400 ;
        RECT 439.600 430.300 440.400 430.400 ;
        RECT 438.100 429.700 440.400 430.300 ;
        RECT 439.600 428.800 440.400 429.700 ;
        RECT 441.000 428.400 441.600 431.800 ;
        RECT 442.800 431.600 443.600 431.800 ;
        RECT 444.400 431.400 445.200 439.800 ;
        RECT 448.800 436.400 449.600 439.800 ;
        RECT 447.600 435.800 449.600 436.400 ;
        RECT 453.200 435.800 454.000 439.800 ;
        RECT 457.400 435.800 458.600 439.800 ;
        RECT 447.600 435.000 448.400 435.800 ;
        RECT 453.200 435.200 453.800 435.800 ;
        RECT 451.000 434.600 454.600 435.200 ;
        RECT 457.200 435.000 458.000 435.800 ;
        RECT 451.000 434.400 451.800 434.600 ;
        RECT 453.800 434.400 454.600 434.600 ;
        RECT 447.600 433.000 448.400 433.200 ;
        RECT 452.200 433.000 453.000 433.200 ;
        RECT 447.600 432.400 453.000 433.000 ;
        RECT 453.600 433.000 455.800 433.600 ;
        RECT 453.600 431.800 454.200 433.000 ;
        RECT 455.000 432.800 455.800 433.000 ;
        RECT 457.400 433.200 458.800 434.000 ;
        RECT 457.400 432.200 458.000 433.200 ;
        RECT 449.400 431.400 454.200 431.800 ;
        RECT 444.400 431.200 454.200 431.400 ;
        RECT 455.600 431.600 458.000 432.200 ;
        RECT 444.400 431.000 450.200 431.200 ;
        RECT 444.400 430.800 450.000 431.000 ;
        RECT 450.800 430.300 451.600 430.400 ;
        RECT 454.000 430.300 454.800 430.400 ;
        RECT 450.800 430.200 454.800 430.300 ;
        RECT 446.600 429.700 454.800 430.200 ;
        RECT 446.600 429.600 451.600 429.700 ;
        RECT 454.000 429.600 454.800 429.700 ;
        RECT 446.600 429.400 447.400 429.600 ;
        RECT 448.200 428.400 449.000 428.600 ;
        RECT 455.600 428.400 456.200 431.600 ;
        RECT 462.000 431.200 462.800 439.800 ;
        RECT 468.400 435.800 469.200 439.800 ;
        RECT 468.600 435.600 469.200 435.800 ;
        RECT 471.600 435.800 472.400 439.800 ;
        RECT 471.600 435.600 472.200 435.800 ;
        RECT 468.600 435.000 472.200 435.600 ;
        RECT 468.600 432.400 469.200 435.000 ;
        RECT 470.000 434.300 470.800 434.400 ;
        RECT 476.400 434.300 477.200 439.800 ;
        RECT 479.600 435.200 480.400 439.800 ;
        RECT 470.000 433.700 477.200 434.300 ;
        RECT 470.000 432.800 470.800 433.700 ;
        RECT 468.400 431.600 469.200 432.400 ;
        RECT 458.600 430.600 462.800 431.200 ;
        RECT 458.600 430.400 459.400 430.600 ;
        RECT 460.200 429.800 461.000 430.000 ;
        RECT 457.200 429.200 461.000 429.800 ;
        RECT 457.200 429.000 458.000 429.200 ;
        RECT 438.000 428.300 438.800 428.400 ;
        RECT 436.400 428.200 438.800 428.300 ;
        RECT 436.400 427.700 439.600 428.200 ;
        RECT 426.600 425.400 427.400 425.600 ;
        RECT 420.400 424.200 421.200 425.000 ;
        RECT 424.600 424.800 427.400 425.400 ;
        RECT 428.400 424.800 429.200 425.600 ;
        RECT 424.600 424.200 425.200 424.800 ;
        RECT 430.000 424.200 430.800 425.000 ;
        RECT 419.800 423.600 421.200 424.200 ;
        RECT 419.800 422.200 421.000 423.600 ;
        RECT 424.400 422.200 425.200 424.200 ;
        RECT 428.800 423.600 430.800 424.200 ;
        RECT 428.800 422.200 429.600 423.600 ;
        RECT 433.200 422.200 434.000 427.000 ;
        RECT 434.800 424.800 435.600 426.400 ;
        RECT 436.400 422.200 437.200 427.700 ;
        RECT 438.000 427.600 439.600 427.700 ;
        RECT 441.000 427.600 443.600 428.400 ;
        RECT 445.200 427.800 456.200 428.400 ;
        RECT 445.200 427.600 446.800 427.800 ;
        RECT 438.800 427.200 439.600 427.600 ;
        RECT 438.200 426.200 441.800 426.600 ;
        RECT 442.800 426.200 443.400 427.600 ;
        RECT 438.000 426.000 442.000 426.200 ;
        RECT 438.000 422.200 438.800 426.000 ;
        RECT 441.200 422.200 442.000 426.000 ;
        RECT 442.800 422.200 443.600 426.200 ;
        RECT 444.400 422.200 445.200 427.000 ;
        RECT 449.400 425.600 450.000 427.800 ;
        RECT 455.000 427.600 455.800 427.800 ;
        RECT 462.000 427.200 462.800 430.600 ;
        RECT 468.600 428.400 469.200 431.600 ;
        RECT 473.200 432.300 474.000 432.400 ;
        RECT 474.800 432.300 475.600 432.400 ;
        RECT 473.200 431.700 475.600 432.300 ;
        RECT 476.400 432.000 477.200 433.700 ;
        RECT 473.200 430.800 474.000 431.700 ;
        RECT 474.800 431.600 475.600 431.700 ;
        RECT 476.200 431.200 477.200 432.000 ;
        RECT 477.800 434.600 480.400 435.200 ;
        RECT 477.800 433.000 478.400 434.600 ;
        RECT 482.800 434.400 483.600 439.800 ;
        RECT 486.000 437.000 486.800 439.800 ;
        RECT 487.600 437.000 488.400 439.800 ;
        RECT 489.200 437.000 490.000 439.800 ;
        RECT 484.200 434.400 488.400 435.200 ;
        RECT 481.000 433.600 483.600 434.400 ;
        RECT 490.800 433.600 491.600 439.800 ;
        RECT 494.000 435.000 494.800 439.800 ;
        RECT 497.200 435.000 498.000 439.800 ;
        RECT 498.800 437.000 499.600 439.800 ;
        RECT 500.400 437.000 501.200 439.800 ;
        RECT 503.600 435.200 504.400 439.800 ;
        RECT 506.800 436.400 507.600 439.800 ;
        RECT 506.800 435.800 507.800 436.400 ;
        RECT 507.200 435.200 507.800 435.800 ;
        RECT 502.400 434.400 506.600 435.200 ;
        RECT 507.200 434.600 509.200 435.200 ;
        RECT 494.000 433.600 496.600 434.400 ;
        RECT 497.200 433.800 503.000 434.400 ;
        RECT 506.000 434.000 506.600 434.400 ;
        RECT 486.000 433.000 486.800 433.200 ;
        RECT 477.800 432.400 486.800 433.000 ;
        RECT 489.200 433.000 490.000 433.200 ;
        RECT 497.200 433.000 497.800 433.800 ;
        RECT 503.600 433.200 505.000 433.800 ;
        RECT 506.000 433.200 507.600 434.000 ;
        RECT 489.200 432.400 497.800 433.000 ;
        RECT 498.800 433.000 505.000 433.200 ;
        RECT 498.800 432.600 504.200 433.000 ;
        RECT 498.800 432.400 499.600 432.600 ;
        RECT 470.800 429.600 472.400 430.400 ;
        RECT 468.600 428.200 470.200 428.400 ;
        RECT 468.600 427.800 470.400 428.200 ;
        RECT 459.000 426.600 462.800 427.200 ;
        RECT 459.000 426.400 459.800 426.600 ;
        RECT 447.600 424.200 448.400 425.000 ;
        RECT 449.200 424.800 450.000 425.600 ;
        RECT 451.000 425.400 451.800 425.600 ;
        RECT 451.000 424.800 453.800 425.400 ;
        RECT 453.200 424.200 453.800 424.800 ;
        RECT 457.200 424.200 458.000 425.000 ;
        RECT 447.600 423.600 449.600 424.200 ;
        RECT 448.800 422.200 449.600 423.600 ;
        RECT 453.200 422.200 454.000 424.200 ;
        RECT 457.200 423.600 458.600 424.200 ;
        RECT 457.400 422.200 458.600 423.600 ;
        RECT 462.000 422.200 462.800 426.600 ;
        RECT 469.600 422.200 470.400 427.800 ;
        RECT 476.200 426.800 477.000 431.200 ;
        RECT 477.800 430.600 478.400 432.400 ;
        RECT 477.600 430.000 478.400 430.600 ;
        RECT 484.400 430.000 507.800 430.600 ;
        RECT 477.600 428.000 478.200 430.000 ;
        RECT 484.400 429.400 485.200 430.000 ;
        RECT 502.000 429.600 502.800 430.000 ;
        RECT 505.200 429.600 506.000 430.000 ;
        RECT 507.000 429.800 507.800 430.000 ;
        RECT 478.800 428.600 482.600 429.400 ;
        RECT 477.600 427.400 478.800 428.000 ;
        RECT 476.200 426.000 477.200 426.800 ;
        RECT 476.400 422.200 477.200 426.000 ;
        RECT 478.000 422.200 478.800 427.400 ;
        RECT 481.800 427.400 482.600 428.600 ;
        RECT 481.800 426.800 483.600 427.400 ;
        RECT 482.800 426.200 483.600 426.800 ;
        RECT 487.600 426.400 488.400 429.200 ;
        RECT 490.800 428.600 494.000 429.400 ;
        RECT 497.800 428.600 499.800 429.400 ;
        RECT 508.400 429.000 509.200 434.600 ;
        RECT 511.600 432.000 512.400 439.800 ;
        RECT 514.800 435.200 515.600 439.800 ;
        RECT 490.400 427.800 491.200 428.000 ;
        RECT 490.400 427.200 494.800 427.800 ;
        RECT 494.000 427.000 494.800 427.200 ;
        RECT 495.600 426.800 496.400 428.400 ;
        RECT 482.800 425.400 485.200 426.200 ;
        RECT 487.600 425.600 488.600 426.400 ;
        RECT 491.600 425.600 493.200 426.400 ;
        RECT 494.000 426.200 494.800 426.400 ;
        RECT 497.800 426.200 498.600 428.600 ;
        RECT 500.400 428.200 509.200 429.000 ;
        RECT 503.800 426.800 506.800 427.600 ;
        RECT 503.800 426.200 504.600 426.800 ;
        RECT 494.000 425.600 498.600 426.200 ;
        RECT 484.400 422.200 485.200 425.400 ;
        RECT 502.000 425.400 504.600 426.200 ;
        RECT 486.000 422.200 486.800 425.000 ;
        RECT 487.600 422.200 488.400 425.000 ;
        RECT 489.200 422.200 490.000 425.000 ;
        RECT 490.800 422.200 491.600 425.000 ;
        RECT 494.000 422.200 494.800 425.000 ;
        RECT 497.200 422.200 498.000 425.000 ;
        RECT 498.800 422.200 499.600 425.000 ;
        RECT 500.400 422.200 501.200 425.000 ;
        RECT 502.000 422.200 502.800 425.400 ;
        RECT 508.400 422.200 509.200 428.200 ;
        RECT 511.400 431.200 512.400 432.000 ;
        RECT 513.000 434.600 515.600 435.200 ;
        RECT 513.000 433.000 513.600 434.600 ;
        RECT 518.000 434.400 518.800 439.800 ;
        RECT 521.200 437.000 522.000 439.800 ;
        RECT 522.800 437.000 523.600 439.800 ;
        RECT 524.400 437.000 525.200 439.800 ;
        RECT 519.400 434.400 523.600 435.200 ;
        RECT 516.200 433.600 518.800 434.400 ;
        RECT 526.000 433.600 526.800 439.800 ;
        RECT 529.200 435.000 530.000 439.800 ;
        RECT 532.400 435.000 533.200 439.800 ;
        RECT 534.000 437.000 534.800 439.800 ;
        RECT 535.600 437.000 536.400 439.800 ;
        RECT 538.800 435.200 539.600 439.800 ;
        RECT 542.000 436.400 542.800 439.800 ;
        RECT 542.000 435.800 543.000 436.400 ;
        RECT 542.400 435.200 543.000 435.800 ;
        RECT 537.600 434.400 541.800 435.200 ;
        RECT 542.400 434.600 544.400 435.200 ;
        RECT 529.200 433.600 531.800 434.400 ;
        RECT 532.400 433.800 538.200 434.400 ;
        RECT 541.200 434.000 541.800 434.400 ;
        RECT 521.200 433.000 522.000 433.200 ;
        RECT 513.000 432.400 522.000 433.000 ;
        RECT 524.400 433.000 525.200 433.200 ;
        RECT 532.400 433.000 533.000 433.800 ;
        RECT 538.800 433.200 540.200 433.800 ;
        RECT 541.200 433.200 542.800 434.000 ;
        RECT 524.400 432.400 533.000 433.000 ;
        RECT 534.000 433.000 540.200 433.200 ;
        RECT 534.000 432.600 539.400 433.000 ;
        RECT 534.000 432.400 534.800 432.600 ;
        RECT 511.400 426.800 512.200 431.200 ;
        RECT 513.000 430.600 513.600 432.400 ;
        RECT 512.800 430.000 513.600 430.600 ;
        RECT 519.600 430.000 543.000 430.600 ;
        RECT 512.800 428.000 513.400 430.000 ;
        RECT 519.600 429.400 520.400 430.000 ;
        RECT 537.200 429.600 538.000 430.000 ;
        RECT 542.000 429.800 543.000 430.000 ;
        RECT 542.000 429.600 542.800 429.800 ;
        RECT 514.000 428.600 517.800 429.400 ;
        RECT 512.800 427.400 514.000 428.000 ;
        RECT 511.400 426.000 512.400 426.800 ;
        RECT 511.600 422.200 512.400 426.000 ;
        RECT 513.200 422.200 514.000 427.400 ;
        RECT 517.000 427.400 517.800 428.600 ;
        RECT 517.000 426.800 518.800 427.400 ;
        RECT 518.000 426.200 518.800 426.800 ;
        RECT 522.800 426.400 523.600 429.200 ;
        RECT 526.000 428.600 529.200 429.400 ;
        RECT 533.000 428.600 535.000 429.400 ;
        RECT 543.600 429.000 544.400 434.600 ;
        RECT 545.200 435.000 546.000 439.000 ;
        RECT 545.200 431.600 545.800 435.000 ;
        RECT 549.400 432.800 550.200 439.800 ;
        RECT 554.800 435.000 555.600 439.000 ;
        RECT 559.000 438.400 559.800 439.800 ;
        RECT 559.000 437.600 560.400 438.400 ;
        RECT 549.400 432.200 551.000 432.800 ;
        RECT 545.200 431.000 549.000 431.600 ;
        RECT 525.600 427.800 526.400 428.000 ;
        RECT 525.600 427.200 530.000 427.800 ;
        RECT 529.200 427.000 530.000 427.200 ;
        RECT 530.800 426.800 531.600 428.400 ;
        RECT 518.000 425.400 520.400 426.200 ;
        RECT 522.800 425.600 523.800 426.400 ;
        RECT 526.800 425.600 528.400 426.400 ;
        RECT 529.200 426.200 530.000 426.400 ;
        RECT 533.000 426.200 533.800 428.600 ;
        RECT 535.600 428.200 544.400 429.000 ;
        RECT 545.200 428.800 546.000 430.400 ;
        RECT 546.800 428.800 547.600 430.400 ;
        RECT 548.400 429.000 549.000 431.000 ;
        RECT 539.000 426.800 542.000 427.600 ;
        RECT 539.000 426.200 539.800 426.800 ;
        RECT 529.200 425.600 533.800 426.200 ;
        RECT 519.600 422.200 520.400 425.400 ;
        RECT 537.200 425.400 539.800 426.200 ;
        RECT 521.200 422.200 522.000 425.000 ;
        RECT 522.800 422.200 523.600 425.000 ;
        RECT 524.400 422.200 525.200 425.000 ;
        RECT 526.000 422.200 526.800 425.000 ;
        RECT 529.200 422.200 530.000 425.000 ;
        RECT 532.400 422.200 533.200 425.000 ;
        RECT 534.000 422.200 534.800 425.000 ;
        RECT 535.600 422.200 536.400 425.000 ;
        RECT 537.200 422.200 538.000 425.400 ;
        RECT 543.600 422.200 544.400 428.200 ;
        RECT 548.400 428.200 549.800 429.000 ;
        RECT 550.400 428.400 551.000 432.200 ;
        RECT 554.800 431.600 555.400 435.000 ;
        RECT 559.000 432.800 559.800 437.600 ;
        RECT 559.000 432.200 560.600 432.800 ;
        RECT 551.600 429.600 552.400 431.200 ;
        RECT 554.800 431.000 558.600 431.600 ;
        RECT 554.800 428.800 555.600 430.400 ;
        RECT 556.400 428.800 557.200 430.400 ;
        RECT 558.000 429.000 558.600 431.000 ;
        RECT 550.400 428.300 552.400 428.400 ;
        RECT 553.200 428.300 554.000 428.400 ;
        RECT 548.400 427.800 549.400 428.200 ;
        RECT 545.200 427.200 549.400 427.800 ;
        RECT 550.400 427.700 554.000 428.300 ;
        RECT 558.000 428.200 559.400 429.000 ;
        RECT 560.000 428.400 560.600 432.200 ;
        RECT 566.000 432.000 566.800 439.800 ;
        RECT 569.200 435.200 570.000 439.800 ;
        RECT 565.800 431.200 566.800 432.000 ;
        RECT 567.400 434.600 570.000 435.200 ;
        RECT 567.400 433.000 568.000 434.600 ;
        RECT 572.400 434.400 573.200 439.800 ;
        RECT 575.600 437.000 576.400 439.800 ;
        RECT 577.200 437.000 578.000 439.800 ;
        RECT 578.800 437.000 579.600 439.800 ;
        RECT 573.800 434.400 578.000 435.200 ;
        RECT 570.600 433.600 573.200 434.400 ;
        RECT 580.400 433.600 581.200 439.800 ;
        RECT 583.600 435.000 584.400 439.800 ;
        RECT 586.800 435.000 587.600 439.800 ;
        RECT 588.400 437.000 589.200 439.800 ;
        RECT 590.000 437.000 590.800 439.800 ;
        RECT 593.200 435.200 594.000 439.800 ;
        RECT 596.400 436.400 597.200 439.800 ;
        RECT 596.400 435.800 597.400 436.400 ;
        RECT 596.800 435.200 597.400 435.800 ;
        RECT 592.000 434.400 596.200 435.200 ;
        RECT 596.800 434.600 598.800 435.200 ;
        RECT 583.600 433.600 586.200 434.400 ;
        RECT 586.800 433.800 592.600 434.400 ;
        RECT 595.600 434.000 596.200 434.400 ;
        RECT 575.600 433.000 576.400 433.200 ;
        RECT 567.400 432.400 576.400 433.000 ;
        RECT 578.800 433.000 579.600 433.200 ;
        RECT 586.800 433.000 587.400 433.800 ;
        RECT 593.200 433.200 594.600 433.800 ;
        RECT 595.600 433.200 597.200 434.000 ;
        RECT 578.800 432.400 587.400 433.000 ;
        RECT 588.400 433.000 594.600 433.200 ;
        RECT 588.400 432.600 593.800 433.000 ;
        RECT 588.400 432.400 589.200 432.600 ;
        RECT 561.200 429.600 562.000 431.200 ;
        RECT 558.000 427.800 559.000 428.200 ;
        RECT 550.400 427.600 552.400 427.700 ;
        RECT 553.200 427.600 554.000 427.700 ;
        RECT 545.200 425.000 545.800 427.200 ;
        RECT 550.400 427.000 551.000 427.600 ;
        RECT 550.200 426.600 551.000 427.000 ;
        RECT 549.400 426.000 551.000 426.600 ;
        RECT 554.800 427.200 559.000 427.800 ;
        RECT 560.000 427.600 562.000 428.400 ;
        RECT 545.200 423.000 546.000 425.000 ;
        RECT 549.400 423.000 550.200 426.000 ;
        RECT 554.800 425.000 555.400 427.200 ;
        RECT 560.000 427.000 560.600 427.600 ;
        RECT 559.800 426.600 560.600 427.000 ;
        RECT 559.000 426.000 560.600 426.600 ;
        RECT 565.800 426.800 566.600 431.200 ;
        RECT 567.400 430.600 568.000 432.400 ;
        RECT 567.200 430.000 568.000 430.600 ;
        RECT 574.000 430.000 597.400 430.600 ;
        RECT 567.200 428.000 567.800 430.000 ;
        RECT 574.000 429.400 574.800 430.000 ;
        RECT 585.200 429.600 586.000 430.000 ;
        RECT 591.600 429.600 592.400 430.000 ;
        RECT 596.600 429.800 597.400 430.000 ;
        RECT 568.400 428.600 572.200 429.400 ;
        RECT 567.200 427.400 568.400 428.000 ;
        RECT 565.800 426.000 566.800 426.800 ;
        RECT 554.800 423.000 555.600 425.000 ;
        RECT 559.000 423.000 559.800 426.000 ;
        RECT 566.000 422.200 566.800 426.000 ;
        RECT 567.600 422.200 568.400 427.400 ;
        RECT 571.400 427.400 572.200 428.600 ;
        RECT 571.400 426.800 573.200 427.400 ;
        RECT 572.400 426.200 573.200 426.800 ;
        RECT 577.200 426.400 578.000 429.200 ;
        RECT 580.400 428.600 583.600 429.400 ;
        RECT 587.400 428.600 589.400 429.400 ;
        RECT 598.000 429.000 598.800 434.600 ;
        RECT 601.200 431.200 602.000 439.800 ;
        RECT 604.400 431.200 605.200 439.800 ;
        RECT 607.600 431.200 608.400 439.800 ;
        RECT 610.800 431.200 611.600 439.800 ;
        RECT 580.000 427.800 580.800 428.000 ;
        RECT 580.000 427.200 584.400 427.800 ;
        RECT 583.600 427.000 584.400 427.200 ;
        RECT 585.200 426.800 586.000 428.400 ;
        RECT 572.400 425.400 574.800 426.200 ;
        RECT 577.200 425.600 578.200 426.400 ;
        RECT 581.200 425.600 582.800 426.400 ;
        RECT 583.600 426.200 584.400 426.400 ;
        RECT 587.400 426.200 588.200 428.600 ;
        RECT 590.000 428.200 598.800 429.000 ;
        RECT 593.400 426.800 596.400 427.600 ;
        RECT 593.400 426.200 594.200 426.800 ;
        RECT 583.600 425.600 588.200 426.200 ;
        RECT 574.000 422.200 574.800 425.400 ;
        RECT 591.600 425.400 594.200 426.200 ;
        RECT 575.600 422.200 576.400 425.000 ;
        RECT 577.200 422.200 578.000 425.000 ;
        RECT 578.800 422.200 579.600 425.000 ;
        RECT 580.400 422.200 581.200 425.000 ;
        RECT 583.600 422.200 584.400 425.000 ;
        RECT 586.800 422.200 587.600 425.000 ;
        RECT 588.400 422.200 589.200 425.000 ;
        RECT 590.000 422.200 590.800 425.000 ;
        RECT 591.600 422.200 592.400 425.400 ;
        RECT 598.000 422.200 598.800 428.200 ;
        RECT 599.600 430.400 602.000 431.200 ;
        RECT 603.000 430.400 605.200 431.200 ;
        RECT 606.200 430.400 608.400 431.200 ;
        RECT 609.800 430.400 611.600 431.200 ;
        RECT 599.600 427.600 600.400 430.400 ;
        RECT 603.000 429.000 603.800 430.400 ;
        RECT 606.200 429.000 607.000 430.400 ;
        RECT 609.800 429.000 610.600 430.400 ;
        RECT 601.200 428.200 603.800 429.000 ;
        RECT 604.600 428.200 607.000 429.000 ;
        RECT 608.000 428.200 610.600 429.000 ;
        RECT 611.400 428.200 613.200 429.000 ;
        RECT 603.000 427.600 603.800 428.200 ;
        RECT 606.200 427.600 607.000 428.200 ;
        RECT 609.800 427.600 610.600 428.200 ;
        RECT 612.400 427.600 613.200 428.200 ;
        RECT 599.600 426.800 602.000 427.600 ;
        RECT 603.000 426.800 605.200 427.600 ;
        RECT 606.200 426.800 608.400 427.600 ;
        RECT 609.800 426.800 611.600 427.600 ;
        RECT 601.200 422.200 602.000 426.800 ;
        RECT 604.400 422.200 605.200 426.800 ;
        RECT 607.600 422.200 608.400 426.800 ;
        RECT 610.800 422.200 611.600 426.800 ;
        RECT 1.200 413.800 2.000 419.800 ;
        RECT 7.600 416.600 8.400 419.800 ;
        RECT 9.200 417.000 10.000 419.800 ;
        RECT 10.800 417.000 11.600 419.800 ;
        RECT 12.400 417.000 13.200 419.800 ;
        RECT 15.600 417.000 16.400 419.800 ;
        RECT 18.800 417.000 19.600 419.800 ;
        RECT 20.400 417.000 21.200 419.800 ;
        RECT 22.000 417.000 22.800 419.800 ;
        RECT 23.600 417.000 24.400 419.800 ;
        RECT 5.800 415.800 8.400 416.600 ;
        RECT 25.200 416.600 26.000 419.800 ;
        RECT 11.800 415.800 16.400 416.400 ;
        RECT 5.800 415.200 6.600 415.800 ;
        RECT 3.600 414.400 6.600 415.200 ;
        RECT 1.200 413.000 10.000 413.800 ;
        RECT 11.800 413.400 12.600 415.800 ;
        RECT 15.600 415.600 16.400 415.800 ;
        RECT 17.200 415.600 18.800 416.400 ;
        RECT 21.800 415.600 22.800 416.400 ;
        RECT 25.200 415.800 27.600 416.600 ;
        RECT 14.000 413.600 14.800 415.200 ;
        RECT 15.600 414.800 16.400 415.000 ;
        RECT 15.600 414.200 20.000 414.800 ;
        RECT 19.200 414.000 20.000 414.200 ;
        RECT 1.200 407.400 2.000 413.000 ;
        RECT 10.600 412.600 12.600 413.400 ;
        RECT 16.400 412.600 19.600 413.400 ;
        RECT 22.000 412.800 22.800 415.600 ;
        RECT 26.800 415.200 27.600 415.800 ;
        RECT 26.800 414.600 28.600 415.200 ;
        RECT 27.800 413.400 28.600 414.600 ;
        RECT 31.600 414.600 32.400 419.800 ;
        RECT 33.200 416.000 34.000 419.800 ;
        RECT 33.200 415.200 34.200 416.000 ;
        RECT 36.400 415.800 37.200 419.800 ;
        RECT 38.000 416.000 38.800 419.800 ;
        RECT 41.200 416.000 42.000 419.800 ;
        RECT 38.000 415.800 42.000 416.000 ;
        RECT 42.800 416.000 43.600 419.800 ;
        RECT 46.000 416.000 46.800 419.800 ;
        RECT 42.800 415.800 46.800 416.000 ;
        RECT 47.600 415.800 48.400 419.800 ;
        RECT 49.200 417.000 50.000 419.000 ;
        RECT 31.600 414.000 32.800 414.600 ;
        RECT 27.800 412.600 31.600 413.400 ;
        RECT 2.600 412.000 3.400 412.200 ;
        RECT 7.600 412.000 8.400 412.400 ;
        RECT 25.200 412.000 26.000 412.600 ;
        RECT 32.200 412.000 32.800 414.000 ;
        RECT 2.600 411.400 26.000 412.000 ;
        RECT 32.000 411.400 32.800 412.000 ;
        RECT 32.000 409.600 32.600 411.400 ;
        RECT 33.400 410.800 34.200 415.200 ;
        RECT 36.600 414.400 37.200 415.800 ;
        RECT 38.200 415.400 41.800 415.800 ;
        RECT 43.000 415.400 46.600 415.800 ;
        RECT 40.400 414.400 41.200 414.800 ;
        RECT 43.600 414.400 44.400 414.800 ;
        RECT 47.600 414.400 48.200 415.800 ;
        RECT 49.200 414.800 49.800 417.000 ;
        RECT 53.400 416.000 54.200 419.000 ;
        RECT 53.400 415.400 55.000 416.000 ;
        RECT 58.800 415.800 59.600 419.800 ;
        RECT 60.400 416.000 61.200 419.800 ;
        RECT 63.600 416.000 64.400 419.800 ;
        RECT 60.400 415.800 64.400 416.000 ;
        RECT 54.200 415.000 55.000 415.400 ;
        RECT 36.400 413.600 39.000 414.400 ;
        RECT 40.400 414.300 42.000 414.400 ;
        RECT 42.800 414.300 44.400 414.400 ;
        RECT 40.400 413.800 44.400 414.300 ;
        RECT 41.200 413.700 43.600 413.800 ;
        RECT 41.200 413.600 42.000 413.700 ;
        RECT 42.800 413.600 43.600 413.700 ;
        RECT 45.800 413.600 48.400 414.400 ;
        RECT 49.200 414.200 53.400 414.800 ;
        RECT 52.400 413.800 53.400 414.200 ;
        RECT 54.400 414.400 55.000 415.000 ;
        RECT 59.000 414.400 59.600 415.800 ;
        RECT 60.600 415.400 64.200 415.800 ;
        RECT 65.200 415.000 66.000 419.800 ;
        RECT 69.600 418.400 70.400 419.800 ;
        RECT 68.400 417.800 70.400 418.400 ;
        RECT 74.000 417.800 74.800 419.800 ;
        RECT 78.200 418.400 79.400 419.800 ;
        RECT 78.000 417.800 79.400 418.400 ;
        RECT 68.400 417.000 69.200 417.800 ;
        RECT 74.000 417.200 74.600 417.800 ;
        RECT 70.000 416.400 70.800 417.200 ;
        RECT 71.800 416.600 74.600 417.200 ;
        RECT 78.000 417.000 78.800 417.800 ;
        RECT 71.800 416.400 72.600 416.600 ;
        RECT 62.800 414.400 63.600 414.800 ;
        RECT 10.800 409.400 11.600 409.600 ;
        RECT 6.200 409.000 11.600 409.400 ;
        RECT 5.400 408.800 11.600 409.000 ;
        RECT 12.600 409.000 21.200 409.600 ;
        RECT 2.800 408.000 4.400 408.800 ;
        RECT 5.400 408.200 6.800 408.800 ;
        RECT 12.600 408.200 13.200 409.000 ;
        RECT 20.400 408.800 21.200 409.000 ;
        RECT 23.600 409.000 32.600 409.600 ;
        RECT 23.600 408.800 24.400 409.000 ;
        RECT 3.800 407.600 4.400 408.000 ;
        RECT 7.400 407.600 13.200 408.200 ;
        RECT 13.800 407.600 16.400 408.400 ;
        RECT 1.200 406.800 3.200 407.400 ;
        RECT 3.800 406.800 8.000 407.600 ;
        RECT 2.600 406.200 3.200 406.800 ;
        RECT 2.600 405.600 3.600 406.200 ;
        RECT 2.800 402.200 3.600 405.600 ;
        RECT 6.000 402.200 6.800 406.800 ;
        RECT 9.200 402.200 10.000 405.000 ;
        RECT 10.800 402.200 11.600 405.000 ;
        RECT 12.400 402.200 13.200 407.000 ;
        RECT 15.600 402.200 16.400 407.000 ;
        RECT 18.800 402.200 19.600 408.400 ;
        RECT 26.800 407.600 29.400 408.400 ;
        RECT 22.000 406.800 26.200 407.600 ;
        RECT 20.400 402.200 21.200 405.000 ;
        RECT 22.000 402.200 22.800 405.000 ;
        RECT 23.600 402.200 24.400 405.000 ;
        RECT 26.800 402.200 27.600 407.600 ;
        RECT 32.000 407.400 32.600 409.000 ;
        RECT 30.000 406.800 32.600 407.400 ;
        RECT 33.200 410.300 34.200 410.800 ;
        RECT 36.400 410.300 37.200 410.400 ;
        RECT 33.200 410.200 37.200 410.300 ;
        RECT 38.400 410.200 39.000 413.600 ;
        RECT 39.600 411.600 40.400 413.200 ;
        RECT 44.400 411.600 45.200 413.200 ;
        RECT 45.800 412.300 46.400 413.600 ;
        RECT 47.600 412.300 48.400 412.400 ;
        RECT 45.800 411.700 48.400 412.300 ;
        RECT 45.800 410.200 46.400 411.700 ;
        RECT 47.600 411.600 48.400 411.700 ;
        RECT 49.200 411.600 50.000 413.200 ;
        RECT 50.800 411.600 51.600 413.200 ;
        RECT 52.400 413.000 53.800 413.800 ;
        RECT 54.400 413.600 56.400 414.400 ;
        RECT 58.800 413.600 61.400 414.400 ;
        RECT 62.800 413.800 64.400 414.400 ;
        RECT 63.600 413.600 64.400 413.800 ;
        RECT 66.000 414.200 67.600 414.400 ;
        RECT 70.200 414.200 70.800 416.400 ;
        RECT 79.800 415.400 80.600 415.600 ;
        RECT 82.800 415.400 83.600 419.800 ;
        RECT 84.400 416.000 85.200 419.800 ;
        RECT 87.600 416.000 88.400 419.800 ;
        RECT 84.400 415.800 88.400 416.000 ;
        RECT 89.200 415.800 90.000 419.800 ;
        RECT 90.800 415.800 91.600 419.800 ;
        RECT 92.400 416.000 93.200 419.800 ;
        RECT 95.600 416.000 96.400 419.800 ;
        RECT 99.800 418.400 100.600 419.800 ;
        RECT 99.800 417.600 101.200 418.400 ;
        RECT 99.800 416.400 100.600 417.600 ;
        RECT 92.400 415.800 96.400 416.000 ;
        RECT 98.800 415.800 100.600 416.400 ;
        RECT 102.000 416.000 102.800 419.800 ;
        RECT 105.200 416.000 106.000 419.800 ;
        RECT 102.000 415.800 106.000 416.000 ;
        RECT 106.800 415.800 107.600 419.800 ;
        RECT 110.000 416.400 110.800 419.800 ;
        RECT 109.800 415.800 110.800 416.400 ;
        RECT 84.600 415.400 88.200 415.800 ;
        RECT 79.800 414.800 83.600 415.400 ;
        RECT 75.800 414.200 76.600 414.400 ;
        RECT 66.000 413.600 77.000 414.200 ;
        RECT 52.400 411.000 53.000 413.000 ;
        RECT 49.200 410.400 53.000 411.000 ;
        RECT 47.600 410.200 48.400 410.400 ;
        RECT 33.200 409.700 37.800 410.200 ;
        RECT 30.000 402.200 30.800 406.800 ;
        RECT 33.200 402.200 34.000 409.700 ;
        RECT 36.400 409.600 37.800 409.700 ;
        RECT 38.400 409.600 39.400 410.200 ;
        RECT 37.200 408.400 37.800 409.600 ;
        RECT 37.200 407.600 38.000 408.400 ;
        RECT 38.600 402.200 39.400 409.600 ;
        RECT 45.400 409.600 46.400 410.200 ;
        RECT 47.000 409.600 48.400 410.200 ;
        RECT 45.400 402.200 46.200 409.600 ;
        RECT 47.000 408.400 47.600 409.600 ;
        RECT 46.800 407.600 47.600 408.400 ;
        RECT 49.200 407.000 49.800 410.400 ;
        RECT 54.400 409.800 55.000 413.600 ;
        RECT 60.800 412.400 61.400 413.600 ;
        RECT 69.000 413.400 69.800 413.600 ;
        RECT 55.600 410.800 56.400 412.400 ;
        RECT 60.400 411.600 61.400 412.400 ;
        RECT 62.000 411.600 62.800 413.200 ;
        RECT 67.400 412.400 68.200 412.600 ;
        RECT 70.000 412.400 70.800 412.600 ;
        RECT 67.400 411.800 72.400 412.400 ;
        RECT 71.600 411.600 72.400 411.800 ;
        RECT 53.400 409.200 55.000 409.800 ;
        RECT 58.800 410.200 59.600 410.400 ;
        RECT 60.800 410.200 61.400 411.600 ;
        RECT 65.200 411.000 70.800 411.200 ;
        RECT 65.200 410.800 71.000 411.000 ;
        RECT 65.200 410.600 75.000 410.800 ;
        RECT 58.800 409.600 60.200 410.200 ;
        RECT 60.800 409.600 61.800 410.200 ;
        RECT 49.200 403.000 50.000 407.000 ;
        RECT 53.400 402.200 54.200 409.200 ;
        RECT 59.600 408.400 60.200 409.600 ;
        RECT 59.600 407.600 60.400 408.400 ;
        RECT 61.000 402.200 61.800 409.600 ;
        RECT 65.200 402.200 66.000 410.600 ;
        RECT 70.200 410.200 75.000 410.600 ;
        RECT 68.400 409.000 73.800 409.600 ;
        RECT 68.400 408.800 69.200 409.000 ;
        RECT 73.000 408.800 73.800 409.000 ;
        RECT 74.400 409.000 75.000 410.200 ;
        RECT 76.400 410.400 77.000 413.600 ;
        RECT 78.000 412.800 78.800 413.000 ;
        RECT 78.000 412.200 81.800 412.800 ;
        RECT 81.000 412.000 81.800 412.200 ;
        RECT 79.400 411.400 80.200 411.600 ;
        RECT 82.800 411.400 83.600 414.800 ;
        RECT 85.200 414.400 86.000 414.800 ;
        RECT 89.200 414.400 89.800 415.800 ;
        RECT 91.000 414.400 91.600 415.800 ;
        RECT 92.600 415.400 96.200 415.800 ;
        RECT 94.800 414.400 95.600 414.800 ;
        RECT 84.400 413.800 86.000 414.400 ;
        RECT 84.400 413.600 85.200 413.800 ;
        RECT 87.400 413.600 90.000 414.400 ;
        RECT 90.800 413.600 93.400 414.400 ;
        RECT 94.800 413.800 96.400 414.400 ;
        RECT 95.600 413.600 96.400 413.800 ;
        RECT 97.200 413.600 98.000 415.200 ;
        RECT 86.000 411.600 86.800 413.200 ;
        RECT 79.400 410.800 83.600 411.400 ;
        RECT 76.400 409.800 78.800 410.400 ;
        RECT 75.800 409.000 76.600 409.200 ;
        RECT 74.400 408.400 76.600 409.000 ;
        RECT 78.200 408.800 78.800 409.800 ;
        RECT 78.200 408.000 79.600 408.800 ;
        RECT 71.800 407.400 72.600 407.600 ;
        RECT 74.600 407.400 75.400 407.600 ;
        RECT 68.400 406.200 69.200 407.000 ;
        RECT 71.800 406.800 75.400 407.400 ;
        RECT 74.000 406.200 74.600 406.800 ;
        RECT 78.000 406.200 78.800 407.000 ;
        RECT 68.400 405.600 70.400 406.200 ;
        RECT 69.600 402.200 70.400 405.600 ;
        RECT 74.000 402.200 74.800 406.200 ;
        RECT 78.200 402.200 79.400 406.200 ;
        RECT 82.800 402.200 83.600 410.800 ;
        RECT 87.400 410.200 88.000 413.600 ;
        RECT 92.800 412.300 93.400 413.600 ;
        RECT 89.300 411.700 93.400 412.300 ;
        RECT 89.300 410.400 89.900 411.700 ;
        RECT 89.200 410.200 90.000 410.400 ;
        RECT 87.000 409.600 88.000 410.200 ;
        RECT 88.600 409.600 90.000 410.200 ;
        RECT 90.800 410.200 91.600 410.400 ;
        RECT 92.800 410.200 93.400 411.700 ;
        RECT 94.000 411.600 94.800 413.200 ;
        RECT 90.800 409.600 92.200 410.200 ;
        RECT 92.800 409.600 93.800 410.200 ;
        RECT 87.000 404.400 87.800 409.600 ;
        RECT 88.600 408.400 89.200 409.600 ;
        RECT 88.400 407.600 89.200 408.400 ;
        RECT 91.600 408.400 92.200 409.600 ;
        RECT 91.600 407.600 92.400 408.400 ;
        RECT 86.000 403.600 87.800 404.400 ;
        RECT 87.000 402.200 87.800 403.600 ;
        RECT 93.000 402.200 93.800 409.600 ;
        RECT 98.800 402.200 99.600 415.800 ;
        RECT 102.200 415.400 105.800 415.800 ;
        RECT 102.800 414.400 103.600 414.800 ;
        RECT 106.800 414.400 107.400 415.800 ;
        RECT 109.800 414.400 110.400 415.800 ;
        RECT 113.200 415.200 114.000 419.800 ;
        RECT 116.400 416.400 117.200 419.800 ;
        RECT 111.400 414.600 114.000 415.200 ;
        RECT 116.200 415.800 117.200 416.400 ;
        RECT 100.400 414.300 101.200 414.400 ;
        RECT 102.000 414.300 103.600 414.400 ;
        RECT 100.400 413.800 103.600 414.300 ;
        RECT 105.000 414.300 107.600 414.400 ;
        RECT 108.400 414.300 109.200 414.400 ;
        RECT 100.400 413.700 102.800 413.800 ;
        RECT 100.400 413.600 101.200 413.700 ;
        RECT 102.000 413.600 102.800 413.700 ;
        RECT 105.000 413.700 109.200 414.300 ;
        RECT 105.000 413.600 107.600 413.700 ;
        RECT 108.400 413.600 109.200 413.700 ;
        RECT 109.800 413.600 110.800 414.400 ;
        RECT 102.000 412.300 102.800 412.400 ;
        RECT 103.600 412.300 104.400 413.200 ;
        RECT 102.000 411.700 104.400 412.300 ;
        RECT 102.000 411.600 102.800 411.700 ;
        RECT 103.600 411.600 104.400 411.700 ;
        RECT 100.400 408.800 101.200 410.400 ;
        RECT 105.000 410.200 105.600 413.600 ;
        RECT 106.800 410.200 107.600 410.400 ;
        RECT 104.600 409.600 105.600 410.200 ;
        RECT 106.200 409.600 107.600 410.200 ;
        RECT 109.800 410.200 110.400 413.600 ;
        RECT 111.400 413.000 112.000 414.600 ;
        RECT 116.200 414.400 116.800 415.800 ;
        RECT 119.600 415.200 120.400 419.800 ;
        RECT 117.800 414.600 120.400 415.200 ;
        RECT 121.200 415.200 122.000 419.800 ;
        RECT 124.400 416.400 125.200 419.800 ;
        RECT 124.400 415.800 125.400 416.400 ;
        RECT 121.200 414.600 123.800 415.200 ;
        RECT 116.200 413.600 117.200 414.400 ;
        RECT 111.000 412.200 112.000 413.000 ;
        RECT 111.400 410.200 112.000 412.200 ;
        RECT 113.000 412.400 113.800 413.200 ;
        RECT 113.000 411.600 114.000 412.400 ;
        RECT 116.200 410.200 116.800 413.600 ;
        RECT 117.800 413.000 118.400 414.600 ;
        RECT 117.400 412.200 118.400 413.000 ;
        RECT 117.800 410.200 118.400 412.200 ;
        RECT 119.400 412.400 120.200 413.200 ;
        RECT 121.400 412.400 122.200 413.200 ;
        RECT 119.400 412.300 120.400 412.400 ;
        RECT 121.200 412.300 122.200 412.400 ;
        RECT 119.400 411.700 122.200 412.300 ;
        RECT 119.400 411.600 120.400 411.700 ;
        RECT 121.200 411.600 122.200 411.700 ;
        RECT 123.200 413.000 123.800 414.600 ;
        RECT 124.800 414.400 125.400 415.800 ;
        RECT 127.600 415.600 128.400 417.200 ;
        RECT 124.400 413.600 125.400 414.400 ;
        RECT 123.200 412.200 124.200 413.000 ;
        RECT 123.200 410.200 123.800 412.200 ;
        RECT 124.800 410.200 125.400 413.600 ;
        RECT 104.600 402.200 105.400 409.600 ;
        RECT 106.200 408.400 106.800 409.600 ;
        RECT 109.800 409.200 110.800 410.200 ;
        RECT 111.400 409.600 114.000 410.200 ;
        RECT 106.000 407.600 106.800 408.400 ;
        RECT 110.000 402.200 110.800 409.200 ;
        RECT 113.200 402.200 114.000 409.600 ;
        RECT 116.200 409.200 117.200 410.200 ;
        RECT 117.800 409.600 120.400 410.200 ;
        RECT 116.400 402.200 117.200 409.200 ;
        RECT 119.600 402.200 120.400 409.600 ;
        RECT 121.200 409.600 123.800 410.200 ;
        RECT 121.200 402.200 122.000 409.600 ;
        RECT 124.400 409.200 125.400 410.200 ;
        RECT 124.400 402.200 125.200 409.200 ;
        RECT 129.200 402.200 130.000 419.800 ;
        RECT 130.800 416.000 131.600 419.800 ;
        RECT 134.000 416.000 134.800 419.800 ;
        RECT 130.800 415.800 134.800 416.000 ;
        RECT 135.600 415.800 136.400 419.800 ;
        RECT 137.200 417.000 138.000 419.000 ;
        RECT 131.000 415.400 134.600 415.800 ;
        RECT 131.600 414.400 132.400 414.800 ;
        RECT 135.600 414.400 136.200 415.800 ;
        RECT 137.200 414.800 137.800 417.000 ;
        RECT 141.400 416.000 142.200 419.000 ;
        RECT 149.400 416.400 150.200 419.800 ;
        RECT 141.400 415.400 143.000 416.000 ;
        RECT 142.200 415.000 143.000 415.400 ;
        RECT 148.400 415.800 150.200 416.400 ;
        RECT 156.400 416.000 157.200 419.800 ;
        RECT 159.600 416.000 160.400 419.800 ;
        RECT 156.400 415.800 160.400 416.000 ;
        RECT 130.800 413.800 132.400 414.400 ;
        RECT 130.800 413.600 131.600 413.800 ;
        RECT 133.800 413.600 136.400 414.400 ;
        RECT 137.200 414.200 141.400 414.800 ;
        RECT 140.400 413.800 141.400 414.200 ;
        RECT 142.400 414.400 143.000 415.000 ;
        RECT 132.400 411.600 133.200 413.200 ;
        RECT 133.800 410.200 134.400 413.600 ;
        RECT 137.200 411.600 138.000 413.200 ;
        RECT 138.800 411.600 139.600 413.200 ;
        RECT 140.400 413.000 141.800 413.800 ;
        RECT 142.400 413.600 144.400 414.400 ;
        RECT 145.200 414.300 146.000 414.400 ;
        RECT 146.800 414.300 147.600 415.200 ;
        RECT 145.200 413.700 147.600 414.300 ;
        RECT 145.200 413.600 146.000 413.700 ;
        RECT 146.800 413.600 147.600 413.700 ;
        RECT 140.400 411.000 141.000 413.000 ;
        RECT 137.200 410.400 141.000 411.000 ;
        RECT 135.600 410.200 136.400 410.400 ;
        RECT 133.400 409.600 134.400 410.200 ;
        RECT 135.000 409.600 136.400 410.200 ;
        RECT 133.400 404.400 134.200 409.600 ;
        RECT 135.000 408.400 135.600 409.600 ;
        RECT 134.800 407.600 135.600 408.400 ;
        RECT 132.400 403.600 134.200 404.400 ;
        RECT 133.400 402.200 134.200 403.600 ;
        RECT 137.200 407.000 137.800 410.400 ;
        RECT 142.400 409.800 143.000 413.600 ;
        RECT 143.600 412.300 144.400 412.400 ;
        RECT 146.800 412.300 147.600 412.400 ;
        RECT 143.600 411.700 147.600 412.300 ;
        RECT 143.600 410.800 144.400 411.700 ;
        RECT 146.800 411.600 147.600 411.700 ;
        RECT 141.400 409.200 143.000 409.800 ;
        RECT 137.200 403.000 138.000 407.000 ;
        RECT 141.400 404.400 142.200 409.200 ;
        RECT 141.400 403.600 142.800 404.400 ;
        RECT 141.400 402.200 142.200 403.600 ;
        RECT 148.400 402.200 149.200 415.800 ;
        RECT 156.600 415.400 160.200 415.800 ;
        RECT 161.200 415.600 162.000 419.800 ;
        RECT 162.800 416.000 163.600 419.800 ;
        RECT 166.000 416.000 166.800 419.800 ;
        RECT 162.800 415.800 166.800 416.000 ;
        RECT 167.600 415.800 168.400 419.800 ;
        RECT 157.200 414.400 158.000 414.800 ;
        RECT 161.200 414.400 161.800 415.600 ;
        RECT 163.000 415.400 166.600 415.800 ;
        RECT 163.600 414.400 164.400 414.800 ;
        RECT 167.600 414.400 168.200 415.800 ;
        RECT 169.200 415.200 170.000 419.800 ;
        RECT 172.400 416.400 173.200 419.800 ;
        RECT 172.400 415.800 173.400 416.400 ;
        RECT 175.600 416.000 176.400 419.800 ;
        RECT 178.800 416.000 179.600 419.800 ;
        RECT 175.600 415.800 179.600 416.000 ;
        RECT 180.400 415.800 181.200 419.800 ;
        RECT 169.200 414.600 171.800 415.200 ;
        RECT 156.400 413.800 158.000 414.400 ;
        RECT 156.400 413.600 157.200 413.800 ;
        RECT 159.400 413.600 162.000 414.400 ;
        RECT 162.800 413.800 164.400 414.400 ;
        RECT 162.800 413.600 163.600 413.800 ;
        RECT 165.800 413.600 168.400 414.400 ;
        RECT 158.000 411.600 158.800 413.200 ;
        RECT 150.000 408.800 150.800 410.400 ;
        RECT 159.400 410.200 160.000 413.600 ;
        RECT 164.400 411.600 165.200 413.200 ;
        RECT 161.200 410.200 162.000 410.400 ;
        RECT 165.800 410.200 166.400 413.600 ;
        RECT 169.400 412.400 170.200 413.200 ;
        RECT 169.200 411.600 170.200 412.400 ;
        RECT 171.200 413.000 171.800 414.600 ;
        RECT 172.800 414.400 173.400 415.800 ;
        RECT 175.800 415.400 179.400 415.800 ;
        RECT 176.400 414.400 177.200 414.800 ;
        RECT 180.400 414.400 181.000 415.800 ;
        RECT 172.400 413.600 173.400 414.400 ;
        RECT 175.600 413.800 177.200 414.400 ;
        RECT 175.600 413.600 176.400 413.800 ;
        RECT 178.600 413.600 181.200 414.400 ;
        RECT 182.000 413.800 182.800 419.800 ;
        RECT 188.400 416.600 189.200 419.800 ;
        RECT 190.000 417.000 190.800 419.800 ;
        RECT 191.600 417.000 192.400 419.800 ;
        RECT 193.200 417.000 194.000 419.800 ;
        RECT 196.400 417.000 197.200 419.800 ;
        RECT 199.600 417.000 200.400 419.800 ;
        RECT 201.200 417.000 202.000 419.800 ;
        RECT 202.800 417.000 203.600 419.800 ;
        RECT 204.400 417.000 205.200 419.800 ;
        RECT 186.600 415.800 189.200 416.600 ;
        RECT 206.000 416.600 206.800 419.800 ;
        RECT 192.600 415.800 197.200 416.400 ;
        RECT 186.600 415.200 187.400 415.800 ;
        RECT 184.400 414.400 187.400 415.200 ;
        RECT 171.200 412.200 172.200 413.000 ;
        RECT 167.600 410.200 168.400 410.400 ;
        RECT 171.200 410.200 171.800 412.200 ;
        RECT 172.800 410.200 173.400 413.600 ;
        RECT 174.000 412.300 174.800 412.400 ;
        RECT 177.200 412.300 178.000 413.200 ;
        RECT 174.000 411.700 178.000 412.300 ;
        RECT 174.000 411.600 174.800 411.700 ;
        RECT 177.200 411.600 178.000 411.700 ;
        RECT 178.600 410.200 179.200 413.600 ;
        RECT 182.000 413.000 190.800 413.800 ;
        RECT 192.600 413.400 193.400 415.800 ;
        RECT 196.400 415.600 197.200 415.800 ;
        RECT 198.000 415.600 199.600 416.400 ;
        RECT 202.600 415.600 203.600 416.400 ;
        RECT 206.000 415.800 208.400 416.600 ;
        RECT 194.800 413.600 195.600 415.200 ;
        RECT 196.400 414.800 197.200 415.000 ;
        RECT 196.400 414.200 200.800 414.800 ;
        RECT 200.000 414.000 200.800 414.200 ;
        RECT 180.400 410.200 181.200 410.400 ;
        RECT 159.000 409.600 160.000 410.200 ;
        RECT 160.600 409.600 162.000 410.200 ;
        RECT 165.400 409.600 166.400 410.200 ;
        RECT 167.000 409.600 168.400 410.200 ;
        RECT 169.200 409.600 171.800 410.200 ;
        RECT 159.000 402.200 159.800 409.600 ;
        RECT 160.600 408.400 161.200 409.600 ;
        RECT 160.400 407.600 161.200 408.400 ;
        RECT 165.400 402.200 166.200 409.600 ;
        RECT 167.000 408.400 167.600 409.600 ;
        RECT 166.800 407.600 167.600 408.400 ;
        RECT 169.200 402.200 170.000 409.600 ;
        RECT 172.400 409.200 173.400 410.200 ;
        RECT 178.200 409.600 179.200 410.200 ;
        RECT 179.800 409.600 181.200 410.200 ;
        RECT 172.400 402.200 173.200 409.200 ;
        RECT 178.200 404.400 179.000 409.600 ;
        RECT 179.800 408.400 180.400 409.600 ;
        RECT 179.600 407.600 180.400 408.400 ;
        RECT 182.000 407.400 182.800 413.000 ;
        RECT 191.400 412.600 193.400 413.400 ;
        RECT 197.200 412.600 200.400 413.400 ;
        RECT 202.800 412.800 203.600 415.600 ;
        RECT 207.600 415.200 208.400 415.800 ;
        RECT 207.600 414.600 209.400 415.200 ;
        RECT 208.600 413.400 209.400 414.600 ;
        RECT 212.400 414.600 213.200 419.800 ;
        RECT 214.000 416.300 214.800 419.800 ;
        RECT 217.200 416.300 218.000 417.200 ;
        RECT 214.000 415.700 218.000 416.300 ;
        RECT 214.000 415.200 215.000 415.700 ;
        RECT 217.200 415.600 218.000 415.700 ;
        RECT 218.800 416.300 219.600 419.800 ;
        RECT 222.000 417.800 222.800 419.800 ;
        RECT 220.400 416.300 221.200 417.200 ;
        RECT 218.800 415.700 221.200 416.300 ;
        RECT 212.400 414.000 213.600 414.600 ;
        RECT 208.600 412.600 212.400 413.400 ;
        RECT 183.400 412.000 184.200 412.200 ;
        RECT 188.400 412.000 189.200 412.400 ;
        RECT 194.800 412.000 195.600 412.400 ;
        RECT 206.000 412.000 206.800 412.600 ;
        RECT 213.000 412.000 213.600 414.000 ;
        RECT 183.400 411.400 206.800 412.000 ;
        RECT 212.800 411.400 213.600 412.000 ;
        RECT 212.800 409.600 213.400 411.400 ;
        RECT 214.200 410.800 215.000 415.200 ;
        RECT 191.600 409.400 192.400 409.600 ;
        RECT 187.000 409.000 192.400 409.400 ;
        RECT 186.200 408.800 192.400 409.000 ;
        RECT 193.400 409.000 202.000 409.600 ;
        RECT 183.600 408.000 185.200 408.800 ;
        RECT 186.200 408.200 187.600 408.800 ;
        RECT 193.400 408.200 194.000 409.000 ;
        RECT 201.200 408.800 202.000 409.000 ;
        RECT 204.400 409.000 213.400 409.600 ;
        RECT 204.400 408.800 205.200 409.000 ;
        RECT 184.600 407.600 185.200 408.000 ;
        RECT 188.200 407.600 194.000 408.200 ;
        RECT 194.600 407.600 197.200 408.400 ;
        RECT 182.000 406.800 184.000 407.400 ;
        RECT 184.600 406.800 188.800 407.600 ;
        RECT 183.400 406.200 184.000 406.800 ;
        RECT 183.400 405.600 184.400 406.200 ;
        RECT 177.200 403.600 179.000 404.400 ;
        RECT 178.200 402.200 179.000 403.600 ;
        RECT 183.600 402.200 184.400 405.600 ;
        RECT 186.800 402.200 187.600 406.800 ;
        RECT 190.000 402.200 190.800 405.000 ;
        RECT 191.600 402.200 192.400 405.000 ;
        RECT 193.200 402.200 194.000 407.000 ;
        RECT 196.400 402.200 197.200 407.000 ;
        RECT 199.600 402.200 200.400 408.400 ;
        RECT 207.600 407.600 210.200 408.400 ;
        RECT 202.800 406.800 207.000 407.600 ;
        RECT 201.200 402.200 202.000 405.000 ;
        RECT 202.800 402.200 203.600 405.000 ;
        RECT 204.400 402.200 205.200 405.000 ;
        RECT 207.600 402.200 208.400 407.600 ;
        RECT 212.800 407.400 213.400 409.000 ;
        RECT 210.800 406.800 213.400 407.400 ;
        RECT 214.000 410.000 215.000 410.800 ;
        RECT 210.800 402.200 211.600 406.800 ;
        RECT 214.000 402.200 214.800 410.000 ;
        RECT 218.800 402.200 219.600 415.700 ;
        RECT 220.400 415.600 221.200 415.700 ;
        RECT 222.200 414.400 222.800 417.800 ;
        RECT 225.400 416.400 226.200 417.200 ;
        RECT 225.200 415.600 226.000 416.400 ;
        RECT 226.800 415.800 227.600 419.800 ;
        RECT 222.000 413.600 222.800 414.400 ;
        RECT 222.200 410.200 222.800 413.600 ;
        RECT 223.600 410.800 224.400 412.400 ;
        RECT 225.200 412.200 226.000 412.400 ;
        RECT 227.000 412.200 227.600 415.800 ;
        RECT 228.400 414.300 229.200 414.400 ;
        RECT 232.800 414.300 233.600 419.800 ;
        RECT 239.600 417.800 240.400 419.800 ;
        RECT 238.000 415.600 238.800 417.200 ;
        RECT 239.800 415.600 240.400 417.800 ;
        RECT 242.800 415.800 243.600 419.800 ;
        RECT 239.800 415.000 242.200 415.600 ;
        RECT 228.400 413.800 233.600 414.300 ;
        RECT 228.400 413.700 233.400 413.800 ;
        RECT 228.400 412.800 229.200 413.700 ;
        RECT 231.800 413.600 233.400 413.700 ;
        RECT 239.600 413.600 240.600 414.400 ;
        RECT 230.000 412.200 230.800 412.400 ;
        RECT 225.200 411.600 227.600 412.200 ;
        RECT 229.200 411.600 230.800 412.200 ;
        RECT 225.400 410.200 226.000 411.600 ;
        RECT 229.200 411.200 230.000 411.600 ;
        RECT 231.800 410.400 232.400 413.600 ;
        RECT 240.000 412.800 240.800 413.600 ;
        RECT 234.000 411.600 235.600 412.400 ;
        RECT 241.600 412.000 242.200 415.000 ;
        RECT 243.000 412.400 243.600 415.800 ;
        RECT 246.000 417.600 246.800 419.800 ;
        RECT 246.000 414.400 246.600 417.600 ;
        RECT 247.600 415.600 248.400 417.200 ;
        RECT 249.200 415.800 250.000 419.800 ;
        RECT 253.600 416.200 255.200 419.800 ;
        RECT 249.200 415.200 251.800 415.800 ;
        RECT 251.000 415.000 251.800 415.200 ;
        RECT 252.400 414.800 254.000 415.600 ;
        RECT 246.000 413.600 246.800 414.400 ;
        RECT 247.600 414.300 248.400 414.400 ;
        RECT 249.200 414.300 250.800 414.400 ;
        RECT 247.600 414.200 250.800 414.300 ;
        RECT 254.600 414.200 255.200 416.200 ;
        RECT 258.800 415.800 259.600 419.800 ;
        RECT 260.400 415.800 261.200 419.800 ;
        RECT 262.000 416.000 262.800 419.800 ;
        RECT 265.200 416.000 266.000 419.800 ;
        RECT 262.000 415.800 266.000 416.000 ;
        RECT 266.800 415.800 267.600 419.800 ;
        RECT 271.200 418.400 272.800 419.800 ;
        RECT 271.200 417.600 274.000 418.400 ;
        RECT 271.200 416.200 272.800 417.600 ;
        RECT 255.800 414.800 256.600 415.600 ;
        RECT 257.200 415.200 259.600 415.800 ;
        RECT 257.200 415.000 258.000 415.200 ;
        RECT 247.600 414.000 251.400 414.200 ;
        RECT 247.600 413.700 253.600 414.000 ;
        RECT 247.600 413.600 248.400 413.700 ;
        RECT 249.200 413.600 253.600 413.700 ;
        RECT 241.400 411.400 242.200 412.000 ;
        RECT 242.800 412.300 243.600 412.400 ;
        RECT 244.400 412.300 245.200 412.400 ;
        RECT 242.800 411.700 245.200 412.300 ;
        RECT 242.800 411.600 243.600 411.700 ;
        RECT 238.000 411.200 242.200 411.400 ;
        RECT 222.000 409.400 223.800 410.200 ;
        RECT 223.000 404.400 223.800 409.400 ;
        RECT 222.000 403.600 223.800 404.400 ;
        RECT 223.000 402.200 223.800 403.600 ;
        RECT 225.200 402.200 226.000 410.200 ;
        RECT 226.800 409.600 230.800 410.200 ;
        RECT 231.600 409.600 232.400 410.400 ;
        RECT 236.400 409.600 237.200 411.200 ;
        RECT 238.000 410.800 242.000 411.200 ;
        RECT 226.800 402.200 227.600 409.600 ;
        RECT 230.000 402.200 230.800 409.600 ;
        RECT 231.800 407.000 232.400 409.600 ;
        RECT 233.200 407.600 234.000 409.200 ;
        RECT 231.800 406.400 235.400 407.000 ;
        RECT 231.800 406.200 232.400 406.400 ;
        RECT 231.600 402.200 232.400 406.200 ;
        RECT 234.800 406.200 235.400 406.400 ;
        RECT 234.800 402.200 235.600 406.200 ;
        RECT 238.000 402.200 238.800 410.800 ;
        RECT 243.000 410.400 243.600 411.600 ;
        RECT 244.400 410.800 245.200 411.700 ;
        RECT 242.800 410.200 243.600 410.400 ;
        RECT 246.000 410.200 246.600 413.600 ;
        RECT 250.800 413.400 253.600 413.600 ;
        RECT 252.800 413.200 253.600 413.400 ;
        RECT 254.200 413.600 255.200 414.200 ;
        RECT 256.000 414.400 256.600 414.800 ;
        RECT 260.600 414.400 261.200 415.800 ;
        RECT 262.200 415.400 265.800 415.800 ;
        RECT 266.800 415.200 269.400 415.800 ;
        RECT 268.600 415.000 269.400 415.200 ;
        RECT 270.000 414.800 271.600 415.600 ;
        RECT 264.400 414.400 265.200 414.800 ;
        RECT 256.000 413.600 256.800 414.400 ;
        RECT 258.000 413.600 259.600 414.400 ;
        RECT 260.400 413.600 263.000 414.400 ;
        RECT 264.400 413.800 266.000 414.400 ;
        RECT 265.200 413.600 266.000 413.800 ;
        RECT 266.800 414.200 268.400 414.400 ;
        RECT 272.200 414.200 272.800 416.200 ;
        RECT 276.400 415.800 277.200 419.800 ;
        RECT 278.000 416.000 278.800 419.800 ;
        RECT 281.200 416.000 282.000 419.800 ;
        RECT 278.000 415.800 282.000 416.000 ;
        RECT 282.800 415.800 283.600 419.800 ;
        RECT 284.400 416.000 285.200 419.800 ;
        RECT 287.600 416.000 288.400 419.800 ;
        RECT 284.400 415.800 288.400 416.000 ;
        RECT 289.200 415.800 290.000 419.800 ;
        RECT 293.400 416.400 294.200 419.800 ;
        RECT 292.400 415.800 294.200 416.400 ;
        RECT 273.400 414.800 274.200 415.600 ;
        RECT 274.800 415.200 277.200 415.800 ;
        RECT 278.200 415.400 281.800 415.800 ;
        RECT 274.800 415.000 275.600 415.200 ;
        RECT 266.800 414.000 269.000 414.200 ;
        RECT 266.800 413.600 271.200 414.000 ;
        RECT 254.200 412.400 254.800 413.600 ;
        RECT 251.400 412.200 252.200 412.400 ;
        RECT 251.400 411.600 253.000 412.200 ;
        RECT 254.000 411.600 254.800 412.400 ;
        RECT 252.200 411.400 253.000 411.600 ;
        RECT 254.200 410.200 254.800 411.600 ;
        RECT 260.400 410.200 261.200 410.400 ;
        RECT 262.400 410.200 263.000 413.600 ;
        RECT 268.400 413.400 271.200 413.600 ;
        RECT 270.400 413.200 271.200 413.400 ;
        RECT 271.800 413.600 272.800 414.200 ;
        RECT 273.600 414.400 274.200 414.800 ;
        RECT 278.800 414.400 279.600 414.800 ;
        RECT 282.800 414.400 283.400 415.800 ;
        RECT 284.600 415.400 288.200 415.800 ;
        RECT 285.200 414.400 286.000 414.800 ;
        RECT 289.200 414.400 289.800 415.800 ;
        RECT 273.600 413.600 274.400 414.400 ;
        RECT 275.600 413.600 277.200 414.400 ;
        RECT 278.000 413.800 279.600 414.400 ;
        RECT 278.000 413.600 278.800 413.800 ;
        RECT 281.000 413.600 283.600 414.400 ;
        RECT 284.400 413.800 286.000 414.400 ;
        RECT 287.400 414.300 290.000 414.400 ;
        RECT 290.800 414.300 291.600 415.200 ;
        RECT 284.400 413.600 285.200 413.800 ;
        RECT 287.400 413.700 291.600 414.300 ;
        RECT 287.400 413.600 290.000 413.700 ;
        RECT 290.800 413.600 291.600 413.700 ;
        RECT 292.400 414.300 293.200 415.800 ;
        RECT 298.800 414.300 299.600 414.400 ;
        RECT 292.400 413.700 299.600 414.300 ;
        RECT 263.600 411.600 264.400 413.200 ;
        RECT 271.800 412.400 272.400 413.600 ;
        RECT 269.000 412.200 269.800 412.400 ;
        RECT 269.000 411.600 270.600 412.200 ;
        RECT 271.600 411.600 272.400 412.400 ;
        RECT 279.600 411.600 280.400 413.200 ;
        RECT 269.800 411.400 270.600 411.600 ;
        RECT 271.800 410.200 272.400 411.600 ;
        RECT 281.000 410.200 281.600 413.600 ;
        RECT 286.000 411.600 286.800 413.200 ;
        RECT 282.800 410.200 283.600 410.400 ;
        RECT 287.400 410.200 288.000 413.600 ;
        RECT 289.200 410.200 290.000 410.400 ;
        RECT 242.200 409.600 243.600 410.200 ;
        RECT 242.200 402.200 243.000 409.600 ;
        RECT 245.000 409.400 246.800 410.200 ;
        RECT 249.200 409.600 251.800 410.200 ;
        RECT 245.000 402.200 245.800 409.400 ;
        RECT 249.200 402.200 250.000 409.600 ;
        RECT 251.000 409.400 251.800 409.600 ;
        RECT 253.600 402.200 255.200 410.200 ;
        RECT 257.200 409.600 259.600 410.200 ;
        RECT 260.400 409.600 261.800 410.200 ;
        RECT 262.400 409.600 263.400 410.200 ;
        RECT 257.200 409.400 258.000 409.600 ;
        RECT 258.800 402.200 259.600 409.600 ;
        RECT 261.200 408.400 261.800 409.600 ;
        RECT 261.200 407.600 262.000 408.400 ;
        RECT 262.600 402.200 263.400 409.600 ;
        RECT 266.800 409.600 269.400 410.200 ;
        RECT 266.800 402.200 267.600 409.600 ;
        RECT 268.600 409.400 269.400 409.600 ;
        RECT 271.200 402.200 272.800 410.200 ;
        RECT 274.800 409.600 277.200 410.200 ;
        RECT 274.800 409.400 275.600 409.600 ;
        RECT 276.400 402.200 277.200 409.600 ;
        RECT 280.600 409.600 281.600 410.200 ;
        RECT 282.200 409.600 283.600 410.200 ;
        RECT 287.000 409.600 288.000 410.200 ;
        RECT 288.600 409.600 290.000 410.200 ;
        RECT 280.600 402.200 281.400 409.600 ;
        RECT 282.200 408.400 282.800 409.600 ;
        RECT 282.000 407.600 283.600 408.400 ;
        RECT 287.000 402.200 287.800 409.600 ;
        RECT 288.600 408.400 289.200 409.600 ;
        RECT 288.400 408.300 289.200 408.400 ;
        RECT 290.800 408.300 291.600 408.400 ;
        RECT 288.400 407.700 291.600 408.300 ;
        RECT 288.400 407.600 289.200 407.700 ;
        RECT 290.800 407.600 291.600 407.700 ;
        RECT 292.400 402.200 293.200 413.700 ;
        RECT 298.800 413.600 299.600 413.700 ;
        RECT 300.400 413.800 301.200 419.800 ;
        RECT 306.800 416.600 307.600 419.800 ;
        RECT 308.400 417.000 309.200 419.800 ;
        RECT 310.000 417.000 310.800 419.800 ;
        RECT 311.600 417.000 312.400 419.800 ;
        RECT 314.800 417.000 315.600 419.800 ;
        RECT 318.000 417.000 318.800 419.800 ;
        RECT 319.600 417.000 320.400 419.800 ;
        RECT 321.200 417.000 322.000 419.800 ;
        RECT 322.800 417.000 323.600 419.800 ;
        RECT 305.000 415.800 307.600 416.600 ;
        RECT 324.400 416.600 325.200 419.800 ;
        RECT 311.000 415.800 315.600 416.400 ;
        RECT 305.000 415.200 305.800 415.800 ;
        RECT 302.800 414.400 305.800 415.200 ;
        RECT 300.400 413.000 309.200 413.800 ;
        RECT 311.000 413.400 311.800 415.800 ;
        RECT 314.800 415.600 315.600 415.800 ;
        RECT 316.400 415.600 318.000 416.400 ;
        RECT 321.000 415.600 322.000 416.400 ;
        RECT 324.400 415.800 326.800 416.600 ;
        RECT 313.200 413.600 314.000 415.200 ;
        RECT 314.800 414.800 315.600 415.000 ;
        RECT 314.800 414.200 319.200 414.800 ;
        RECT 318.400 414.000 319.200 414.200 ;
        RECT 294.000 408.800 294.800 410.400 ;
        RECT 300.400 407.400 301.200 413.000 ;
        RECT 309.800 412.600 311.800 413.400 ;
        RECT 315.600 412.600 318.800 413.400 ;
        RECT 321.200 412.800 322.000 415.600 ;
        RECT 326.000 415.200 326.800 415.800 ;
        RECT 326.000 414.600 327.800 415.200 ;
        RECT 327.000 413.400 327.800 414.600 ;
        RECT 330.800 414.600 331.600 419.800 ;
        RECT 332.400 416.000 333.200 419.800 ;
        RECT 332.400 415.200 333.400 416.000 ;
        RECT 330.800 414.000 332.000 414.600 ;
        RECT 327.000 412.600 330.800 413.400 ;
        RECT 301.800 412.000 302.600 412.200 ;
        RECT 303.600 412.000 304.400 412.400 ;
        RECT 306.800 412.000 307.600 412.400 ;
        RECT 324.400 412.000 325.200 412.600 ;
        RECT 331.400 412.000 332.000 414.000 ;
        RECT 301.800 411.400 325.200 412.000 ;
        RECT 331.200 411.400 332.000 412.000 ;
        RECT 331.200 409.600 331.800 411.400 ;
        RECT 332.600 410.800 333.400 415.200 ;
        RECT 335.600 415.000 336.400 419.800 ;
        RECT 340.000 418.400 340.800 419.800 ;
        RECT 338.800 417.800 340.800 418.400 ;
        RECT 344.400 417.800 345.200 419.800 ;
        RECT 348.600 418.400 349.800 419.800 ;
        RECT 348.400 417.800 349.800 418.400 ;
        RECT 338.800 417.000 339.600 417.800 ;
        RECT 344.400 417.200 345.000 417.800 ;
        RECT 340.400 416.400 341.200 417.200 ;
        RECT 342.200 416.600 345.000 417.200 ;
        RECT 348.400 417.000 349.200 417.800 ;
        RECT 342.200 416.400 343.000 416.600 ;
        RECT 336.400 414.200 338.000 414.400 ;
        RECT 340.600 414.200 341.200 416.400 ;
        RECT 350.200 415.400 351.000 415.600 ;
        RECT 353.200 415.400 354.000 419.800 ;
        RECT 354.800 416.000 355.600 419.800 ;
        RECT 358.000 416.000 358.800 419.800 ;
        RECT 354.800 415.800 358.800 416.000 ;
        RECT 359.600 415.800 360.400 419.800 ;
        RECT 355.000 415.400 358.600 415.800 ;
        RECT 350.200 414.800 354.000 415.400 ;
        RECT 346.200 414.200 347.000 414.400 ;
        RECT 336.400 413.600 347.400 414.200 ;
        RECT 339.400 413.400 340.200 413.600 ;
        RECT 337.800 412.400 338.600 412.600 ;
        RECT 337.800 411.800 342.800 412.400 ;
        RECT 342.000 411.600 342.800 411.800 ;
        RECT 310.000 409.400 310.800 409.600 ;
        RECT 305.400 409.000 310.800 409.400 ;
        RECT 304.600 408.800 310.800 409.000 ;
        RECT 311.800 409.000 320.400 409.600 ;
        RECT 302.000 408.000 303.600 408.800 ;
        RECT 304.600 408.200 306.000 408.800 ;
        RECT 311.800 408.200 312.400 409.000 ;
        RECT 319.600 408.800 320.400 409.000 ;
        RECT 322.800 409.000 331.800 409.600 ;
        RECT 322.800 408.800 323.600 409.000 ;
        RECT 303.000 407.600 303.600 408.000 ;
        RECT 306.600 407.600 312.400 408.200 ;
        RECT 313.000 407.600 315.600 408.400 ;
        RECT 300.400 406.800 302.400 407.400 ;
        RECT 303.000 406.800 307.200 407.600 ;
        RECT 301.800 406.200 302.400 406.800 ;
        RECT 301.800 405.600 302.800 406.200 ;
        RECT 302.000 402.200 302.800 405.600 ;
        RECT 305.200 402.200 306.000 406.800 ;
        RECT 308.400 402.200 309.200 405.000 ;
        RECT 310.000 402.200 310.800 405.000 ;
        RECT 311.600 402.200 312.400 407.000 ;
        RECT 314.800 402.200 315.600 407.000 ;
        RECT 318.000 402.200 318.800 408.400 ;
        RECT 326.000 407.600 328.600 408.400 ;
        RECT 321.200 406.800 325.400 407.600 ;
        RECT 319.600 402.200 320.400 405.000 ;
        RECT 321.200 402.200 322.000 405.000 ;
        RECT 322.800 402.200 323.600 405.000 ;
        RECT 326.000 402.200 326.800 407.600 ;
        RECT 331.200 407.400 331.800 409.000 ;
        RECT 329.200 406.800 331.800 407.400 ;
        RECT 332.400 410.000 333.400 410.800 ;
        RECT 335.600 411.000 341.200 411.200 ;
        RECT 335.600 410.800 341.400 411.000 ;
        RECT 335.600 410.600 345.400 410.800 ;
        RECT 329.200 402.200 330.000 406.800 ;
        RECT 332.400 402.200 333.200 410.000 ;
        RECT 335.600 402.200 336.400 410.600 ;
        RECT 340.600 410.200 345.400 410.600 ;
        RECT 338.800 409.000 344.200 409.600 ;
        RECT 338.800 408.800 339.600 409.000 ;
        RECT 343.400 408.800 344.200 409.000 ;
        RECT 344.800 409.000 345.400 410.200 ;
        RECT 346.800 410.400 347.400 413.600 ;
        RECT 348.400 412.800 349.200 413.000 ;
        RECT 348.400 412.200 352.200 412.800 ;
        RECT 351.400 412.000 352.200 412.200 ;
        RECT 349.800 411.400 350.600 411.600 ;
        RECT 353.200 411.400 354.000 414.800 ;
        RECT 355.600 414.400 356.400 414.800 ;
        RECT 359.600 414.400 360.200 415.800 ;
        RECT 361.200 415.600 362.000 419.800 ;
        RECT 362.800 416.000 363.600 419.800 ;
        RECT 366.000 416.000 366.800 419.800 ;
        RECT 362.800 415.800 366.800 416.000 ;
        RECT 361.400 414.400 362.000 415.600 ;
        RECT 363.000 415.400 366.600 415.800 ;
        RECT 367.600 415.600 368.400 417.200 ;
        RECT 365.200 414.400 366.000 414.800 ;
        RECT 354.800 413.800 356.400 414.400 ;
        RECT 354.800 413.600 355.600 413.800 ;
        RECT 357.800 413.600 360.400 414.400 ;
        RECT 361.200 413.600 363.800 414.400 ;
        RECT 365.200 413.800 366.800 414.400 ;
        RECT 366.000 413.600 366.800 413.800 ;
        RECT 356.400 411.600 357.200 413.200 ;
        RECT 357.800 412.300 358.400 413.600 ;
        RECT 357.800 411.700 361.900 412.300 ;
        RECT 349.800 410.800 354.000 411.400 ;
        RECT 346.800 409.800 349.200 410.400 ;
        RECT 346.200 409.000 347.000 409.200 ;
        RECT 344.800 408.400 347.000 409.000 ;
        RECT 348.600 408.800 349.200 409.800 ;
        RECT 348.600 408.400 350.000 408.800 ;
        RECT 348.600 408.000 350.800 408.400 ;
        RECT 349.400 407.600 350.800 408.000 ;
        RECT 342.200 407.400 343.000 407.600 ;
        RECT 345.000 407.400 345.800 407.600 ;
        RECT 338.800 406.200 339.600 407.000 ;
        RECT 342.200 406.800 345.800 407.400 ;
        RECT 344.400 406.200 345.000 406.800 ;
        RECT 348.400 406.200 349.200 407.000 ;
        RECT 338.800 405.600 340.800 406.200 ;
        RECT 340.000 402.200 340.800 405.600 ;
        RECT 344.400 402.200 345.200 406.200 ;
        RECT 348.600 402.200 349.800 406.200 ;
        RECT 353.200 402.200 354.000 410.800 ;
        RECT 357.800 410.200 358.400 411.700 ;
        RECT 361.300 410.400 361.900 411.700 ;
        RECT 359.600 410.200 360.400 410.400 ;
        RECT 357.400 409.600 358.400 410.200 ;
        RECT 359.000 409.600 360.400 410.200 ;
        RECT 361.200 410.200 362.000 410.400 ;
        RECT 363.200 410.200 363.800 413.600 ;
        RECT 364.400 411.600 365.200 413.200 ;
        RECT 361.200 409.600 362.600 410.200 ;
        RECT 363.200 409.600 364.200 410.200 ;
        RECT 357.400 402.200 358.200 409.600 ;
        RECT 359.000 408.400 359.600 409.600 ;
        RECT 358.800 407.600 359.600 408.400 ;
        RECT 362.000 408.400 362.600 409.600 ;
        RECT 362.000 407.600 362.800 408.400 ;
        RECT 363.400 402.200 364.200 409.600 ;
        RECT 369.200 402.200 370.000 419.800 ;
        RECT 370.800 416.000 371.600 419.800 ;
        RECT 374.000 416.000 374.800 419.800 ;
        RECT 370.800 415.800 374.800 416.000 ;
        RECT 375.600 415.800 376.400 419.800 ;
        RECT 377.200 415.800 378.000 419.800 ;
        RECT 378.800 416.000 379.600 419.800 ;
        RECT 382.000 416.000 382.800 419.800 ;
        RECT 378.800 415.800 382.800 416.000 ;
        RECT 371.000 415.400 374.600 415.800 ;
        RECT 371.600 414.400 372.400 414.800 ;
        RECT 375.600 414.400 376.200 415.800 ;
        RECT 377.400 414.400 378.000 415.800 ;
        RECT 379.000 415.400 382.600 415.800 ;
        RECT 383.600 415.600 384.400 417.200 ;
        RECT 381.200 414.400 382.000 414.800 ;
        RECT 370.800 413.800 372.400 414.400 ;
        RECT 370.800 413.600 371.600 413.800 ;
        RECT 373.800 413.600 376.400 414.400 ;
        RECT 377.200 413.600 379.800 414.400 ;
        RECT 381.200 413.800 382.800 414.400 ;
        RECT 382.000 413.600 382.800 413.800 ;
        RECT 385.200 414.300 386.000 419.800 ;
        RECT 386.800 416.000 387.600 419.800 ;
        RECT 390.000 416.000 390.800 419.800 ;
        RECT 386.800 415.800 390.800 416.000 ;
        RECT 387.000 415.400 390.600 415.800 ;
        RECT 391.600 415.600 392.400 419.800 ;
        RECT 387.600 414.400 388.400 414.800 ;
        RECT 391.600 414.400 392.200 415.600 ;
        RECT 386.800 414.300 388.400 414.400 ;
        RECT 385.200 413.800 388.400 414.300 ;
        RECT 385.200 413.700 387.600 413.800 ;
        RECT 372.400 411.600 373.200 413.200 ;
        RECT 373.800 412.300 374.400 413.600 ;
        RECT 373.800 411.700 377.900 412.300 ;
        RECT 373.800 410.200 374.400 411.700 ;
        RECT 377.300 410.400 377.900 411.700 ;
        RECT 375.600 410.200 376.400 410.400 ;
        RECT 373.400 409.600 374.400 410.200 ;
        RECT 375.000 409.600 376.400 410.200 ;
        RECT 377.200 410.200 378.000 410.400 ;
        RECT 379.200 410.200 379.800 413.600 ;
        RECT 380.400 411.600 381.200 413.200 ;
        RECT 377.200 409.600 378.600 410.200 ;
        RECT 379.200 409.600 380.200 410.200 ;
        RECT 373.400 402.200 374.200 409.600 ;
        RECT 375.000 408.400 375.600 409.600 ;
        RECT 374.800 407.600 375.600 408.400 ;
        RECT 378.000 408.400 378.600 409.600 ;
        RECT 378.000 407.600 378.800 408.400 ;
        RECT 379.400 404.400 380.200 409.600 ;
        RECT 379.400 403.600 381.200 404.400 ;
        RECT 379.400 402.200 380.200 403.600 ;
        RECT 385.200 402.200 386.000 413.700 ;
        RECT 386.800 413.600 387.600 413.700 ;
        RECT 389.800 413.600 392.400 414.400 ;
        RECT 396.800 414.200 397.600 419.800 ;
        RECT 403.200 414.200 404.000 419.800 ;
        RECT 406.000 416.000 406.800 419.800 ;
        RECT 409.200 416.000 410.000 419.800 ;
        RECT 406.000 415.800 410.000 416.000 ;
        RECT 410.800 415.800 411.600 419.800 ;
        RECT 406.200 415.400 409.800 415.800 ;
        RECT 406.800 414.400 407.600 414.800 ;
        RECT 410.800 414.400 411.400 415.800 ;
        RECT 412.400 415.600 413.200 417.200 ;
        RECT 396.800 413.800 398.600 414.200 ;
        RECT 403.200 413.800 405.000 414.200 ;
        RECT 397.000 413.600 398.600 413.800 ;
        RECT 403.400 413.600 405.000 413.800 ;
        RECT 406.000 413.800 407.600 414.400 ;
        RECT 406.000 413.600 406.800 413.800 ;
        RECT 409.000 413.600 411.600 414.400 ;
        RECT 414.000 414.300 414.800 419.800 ;
        RECT 415.600 416.000 416.400 419.800 ;
        RECT 418.800 416.000 419.600 419.800 ;
        RECT 415.600 415.800 419.600 416.000 ;
        RECT 420.400 415.800 421.200 419.800 ;
        RECT 422.000 416.000 422.800 419.800 ;
        RECT 425.200 416.000 426.000 419.800 ;
        RECT 422.000 415.800 426.000 416.000 ;
        RECT 426.800 415.800 427.600 419.800 ;
        RECT 428.400 416.000 429.200 419.800 ;
        RECT 431.600 416.000 432.400 419.800 ;
        RECT 428.400 415.800 432.400 416.000 ;
        RECT 433.200 415.800 434.000 419.800 ;
        RECT 437.400 416.400 438.200 419.800 ;
        RECT 436.400 415.800 438.200 416.400 ;
        RECT 415.800 415.400 419.400 415.800 ;
        RECT 416.400 414.400 417.200 414.800 ;
        RECT 420.400 414.400 421.000 415.800 ;
        RECT 422.200 415.400 425.800 415.800 ;
        RECT 422.800 414.400 423.600 414.800 ;
        RECT 426.800 414.400 427.400 415.800 ;
        RECT 428.600 415.400 432.200 415.800 ;
        RECT 429.200 414.400 430.000 414.800 ;
        RECT 433.200 414.400 433.800 415.800 ;
        RECT 415.600 414.300 417.200 414.400 ;
        RECT 414.000 413.800 417.200 414.300 ;
        RECT 414.000 413.700 416.400 413.800 ;
        RECT 388.400 411.600 389.200 413.200 ;
        RECT 389.800 410.200 390.400 413.600 ;
        RECT 394.800 411.600 396.400 412.400 ;
        RECT 391.600 410.200 392.400 410.400 ;
        RECT 389.400 409.600 390.400 410.200 ;
        RECT 391.000 409.600 392.400 410.200 ;
        RECT 393.200 409.600 394.000 411.200 ;
        RECT 398.000 410.400 398.600 413.600 ;
        RECT 401.200 411.600 402.800 412.400 ;
        RECT 404.400 412.300 405.000 413.600 ;
        RECT 406.000 412.300 406.800 412.400 ;
        RECT 404.400 411.700 406.800 412.300 ;
        RECT 398.000 409.600 398.800 410.400 ;
        RECT 399.600 409.600 400.400 411.200 ;
        RECT 404.400 410.400 405.000 411.700 ;
        RECT 406.000 411.600 406.800 411.700 ;
        RECT 407.600 411.600 408.400 413.200 ;
        RECT 404.400 409.600 405.200 410.400 ;
        RECT 409.000 410.200 409.600 413.600 ;
        RECT 410.800 410.200 411.600 410.400 ;
        RECT 408.600 409.600 409.600 410.200 ;
        RECT 410.200 409.600 411.600 410.200 ;
        RECT 389.400 402.200 390.200 409.600 ;
        RECT 391.000 408.400 391.600 409.600 ;
        RECT 390.800 407.600 391.600 408.400 ;
        RECT 396.400 407.600 397.200 409.200 ;
        RECT 398.000 407.000 398.600 409.600 ;
        RECT 402.800 407.600 403.600 409.200 ;
        RECT 404.400 407.000 405.000 409.600 ;
        RECT 395.000 406.400 398.600 407.000 ;
        RECT 394.800 402.200 395.600 406.400 ;
        RECT 398.000 406.200 398.600 406.400 ;
        RECT 401.400 406.400 405.000 407.000 ;
        RECT 401.400 406.200 402.000 406.400 ;
        RECT 398.000 402.200 398.800 406.200 ;
        RECT 401.200 402.200 402.000 406.200 ;
        RECT 404.400 406.200 405.000 406.400 ;
        RECT 404.400 402.200 405.200 406.200 ;
        RECT 408.600 402.200 409.400 409.600 ;
        RECT 410.200 408.400 410.800 409.600 ;
        RECT 410.000 407.600 410.800 408.400 ;
        RECT 414.000 402.200 414.800 413.700 ;
        RECT 415.600 413.600 416.400 413.700 ;
        RECT 418.600 413.600 421.200 414.400 ;
        RECT 422.000 413.800 423.600 414.400 ;
        RECT 422.000 413.600 422.800 413.800 ;
        RECT 425.000 413.600 427.600 414.400 ;
        RECT 428.400 413.800 430.000 414.400 ;
        RECT 428.400 413.600 429.200 413.800 ;
        RECT 431.400 413.600 434.000 414.400 ;
        RECT 434.800 413.600 435.600 415.200 ;
        RECT 417.200 411.600 418.000 413.200 ;
        RECT 418.600 412.300 419.200 413.600 ;
        RECT 423.600 412.300 424.400 413.200 ;
        RECT 418.600 411.700 424.400 412.300 ;
        RECT 418.600 410.200 419.200 411.700 ;
        RECT 423.600 411.600 424.400 411.700 ;
        RECT 420.400 410.200 421.200 410.400 ;
        RECT 425.000 410.200 425.600 413.600 ;
        RECT 430.000 411.600 430.800 413.200 ;
        RECT 426.800 410.200 427.600 410.400 ;
        RECT 431.400 410.200 432.000 413.600 ;
        RECT 433.200 410.200 434.000 410.400 ;
        RECT 418.200 409.600 419.200 410.200 ;
        RECT 419.800 409.600 421.200 410.200 ;
        RECT 424.600 409.600 425.600 410.200 ;
        RECT 426.200 409.600 427.600 410.200 ;
        RECT 431.000 409.600 432.000 410.200 ;
        RECT 432.600 409.600 434.000 410.200 ;
        RECT 418.200 402.200 419.000 409.600 ;
        RECT 419.800 408.400 420.400 409.600 ;
        RECT 419.600 407.600 420.400 408.400 ;
        RECT 424.600 404.400 425.400 409.600 ;
        RECT 426.200 408.400 426.800 409.600 ;
        RECT 426.000 407.600 426.800 408.400 ;
        RECT 431.000 404.400 431.800 409.600 ;
        RECT 432.600 408.400 433.200 409.600 ;
        RECT 432.400 407.600 433.200 408.400 ;
        RECT 423.600 403.600 425.400 404.400 ;
        RECT 430.000 403.600 431.800 404.400 ;
        RECT 424.600 402.200 425.400 403.600 ;
        RECT 431.000 402.200 431.800 403.600 ;
        RECT 436.400 402.200 437.200 415.800 ;
        RECT 438.000 410.300 438.800 410.400 ;
        RECT 439.600 410.300 440.400 419.800 ;
        RECT 441.200 415.600 442.000 417.200 ;
        RECT 442.800 416.000 443.600 419.800 ;
        RECT 446.000 416.000 446.800 419.800 ;
        RECT 442.800 415.800 446.800 416.000 ;
        RECT 447.600 415.800 448.400 419.800 ;
        RECT 451.800 418.400 452.600 419.800 ;
        RECT 450.800 417.600 452.600 418.400 ;
        RECT 451.800 416.400 452.600 417.600 ;
        RECT 450.800 415.800 452.600 416.400 ;
        RECT 443.000 415.400 446.600 415.800 ;
        RECT 443.600 414.400 444.400 414.800 ;
        RECT 447.600 414.400 448.200 415.800 ;
        RECT 442.800 413.800 444.400 414.400 ;
        RECT 442.800 413.600 443.600 413.800 ;
        RECT 445.800 413.600 448.400 414.400 ;
        RECT 449.200 413.600 450.000 415.200 ;
        RECT 444.400 411.600 445.200 413.200 ;
        RECT 438.000 409.700 440.400 410.300 ;
        RECT 445.800 410.200 446.400 413.600 ;
        RECT 447.600 410.200 448.400 410.400 ;
        RECT 438.000 408.800 438.800 409.700 ;
        RECT 439.600 402.200 440.400 409.700 ;
        RECT 445.400 409.600 446.400 410.200 ;
        RECT 447.000 409.600 448.400 410.200 ;
        RECT 445.400 404.400 446.200 409.600 ;
        RECT 447.000 408.400 447.600 409.600 ;
        RECT 446.800 407.600 447.600 408.400 ;
        RECT 444.400 403.600 446.200 404.400 ;
        RECT 445.400 402.200 446.200 403.600 ;
        RECT 450.800 402.200 451.600 415.800 ;
        RECT 452.400 414.300 453.200 414.400 ;
        RECT 454.000 414.300 454.800 415.200 ;
        RECT 452.400 413.700 454.800 414.300 ;
        RECT 452.400 413.600 453.200 413.700 ;
        RECT 454.000 413.600 454.800 413.700 ;
        RECT 455.600 414.300 456.400 419.800 ;
        RECT 462.000 415.800 462.800 419.800 ;
        RECT 463.600 416.000 464.400 419.800 ;
        RECT 466.800 416.000 467.600 419.800 ;
        RECT 463.600 415.800 467.600 416.000 ;
        RECT 468.400 415.800 469.200 419.800 ;
        RECT 470.000 416.000 470.800 419.800 ;
        RECT 473.200 416.000 474.000 419.800 ;
        RECT 470.000 415.800 474.000 416.000 ;
        RECT 474.800 415.800 475.600 419.800 ;
        RECT 479.200 418.400 480.800 419.800 ;
        RECT 479.200 417.600 482.000 418.400 ;
        RECT 479.200 416.200 480.800 417.600 ;
        RECT 462.200 414.400 462.800 415.800 ;
        RECT 463.800 415.400 467.400 415.800 ;
        RECT 466.000 414.400 466.800 414.800 ;
        RECT 468.600 414.400 469.200 415.800 ;
        RECT 470.200 415.400 473.800 415.800 ;
        RECT 474.800 415.200 477.200 415.800 ;
        RECT 476.400 415.000 477.200 415.200 ;
        RECT 477.800 414.800 478.600 415.600 ;
        RECT 472.400 414.400 473.200 414.800 ;
        RECT 477.800 414.400 478.400 414.800 ;
        RECT 460.400 414.300 461.200 414.400 ;
        RECT 455.600 413.700 461.200 414.300 ;
        RECT 455.600 412.300 456.400 413.700 ;
        RECT 460.400 413.600 461.200 413.700 ;
        RECT 462.000 413.600 464.600 414.400 ;
        RECT 466.000 413.800 467.600 414.400 ;
        RECT 466.800 413.600 467.600 413.800 ;
        RECT 468.400 413.600 471.000 414.400 ;
        RECT 472.400 413.800 474.000 414.400 ;
        RECT 473.200 413.600 474.000 413.800 ;
        RECT 474.800 413.600 476.400 414.400 ;
        RECT 477.600 413.600 478.400 414.400 ;
        RECT 452.500 411.700 456.400 412.300 ;
        RECT 452.500 410.400 453.100 411.700 ;
        RECT 452.400 408.800 453.200 410.400 ;
        RECT 455.600 402.200 456.400 411.700 ;
        RECT 457.200 410.300 458.000 410.400 ;
        RECT 462.000 410.300 462.800 410.400 ;
        RECT 457.200 410.200 462.800 410.300 ;
        RECT 464.000 410.200 464.600 413.600 ;
        RECT 465.200 411.600 466.000 413.200 ;
        RECT 468.400 410.200 469.200 410.400 ;
        RECT 470.400 410.200 471.000 413.600 ;
        RECT 471.600 411.600 472.400 413.200 ;
        RECT 479.200 412.800 479.800 416.200 ;
        RECT 484.400 415.800 485.200 419.800 ;
        RECT 486.000 415.800 486.800 419.800 ;
        RECT 487.600 416.000 488.400 419.800 ;
        RECT 490.800 416.000 491.600 419.800 ;
        RECT 493.000 416.800 493.800 419.800 ;
        RECT 487.600 415.800 491.600 416.000 ;
        RECT 492.400 415.800 493.800 416.800 ;
        RECT 497.200 415.800 498.000 419.800 ;
        RECT 499.000 416.400 499.800 417.200 ;
        RECT 480.400 415.400 482.000 415.600 ;
        RECT 480.400 414.800 482.400 415.400 ;
        RECT 483.000 415.200 485.200 415.800 ;
        RECT 483.000 415.000 483.800 415.200 ;
        RECT 481.800 414.400 482.400 414.800 ;
        RECT 486.200 414.400 486.800 415.800 ;
        RECT 487.800 415.400 491.400 415.800 ;
        RECT 490.000 414.400 490.800 414.800 ;
        RECT 480.400 413.400 481.200 414.200 ;
        RECT 481.800 413.800 485.200 414.400 ;
        RECT 483.600 413.600 485.200 413.800 ;
        RECT 486.000 413.600 488.600 414.400 ;
        RECT 490.000 413.800 491.600 414.400 ;
        RECT 490.800 413.600 491.600 413.800 ;
        RECT 478.800 412.400 479.800 412.800 ;
        RECT 478.000 412.200 479.800 412.400 ;
        RECT 480.600 412.800 481.200 413.400 ;
        RECT 480.600 412.200 483.200 412.800 ;
        RECT 478.000 411.600 479.400 412.200 ;
        RECT 482.400 412.000 483.200 412.200 ;
        RECT 478.800 410.200 479.400 411.600 ;
        RECT 480.200 411.400 481.000 411.600 ;
        RECT 480.200 410.800 483.600 411.400 ;
        RECT 483.000 410.200 483.600 410.800 ;
        RECT 486.000 410.200 486.800 410.400 ;
        RECT 488.000 410.200 488.600 413.600 ;
        RECT 489.200 411.600 490.000 413.200 ;
        RECT 490.900 412.300 491.500 413.600 ;
        RECT 492.400 412.400 493.000 415.800 ;
        RECT 497.200 415.600 497.800 415.800 ;
        RECT 498.800 415.600 499.600 416.400 ;
        RECT 500.400 415.800 501.200 419.800 ;
        RECT 507.800 416.400 508.600 419.800 ;
        RECT 512.600 416.400 513.400 419.800 ;
        RECT 496.000 415.200 497.800 415.600 ;
        RECT 493.600 415.000 497.800 415.200 ;
        RECT 493.600 414.600 496.600 415.000 ;
        RECT 493.600 414.400 494.400 414.600 ;
        RECT 492.400 412.300 493.200 412.400 ;
        RECT 490.900 411.700 493.200 412.300 ;
        RECT 492.400 411.600 493.200 411.700 ;
        RECT 492.400 410.200 493.000 411.600 ;
        RECT 493.800 411.000 494.400 414.400 ;
        RECT 497.200 414.300 498.000 414.400 ;
        RECT 498.900 414.300 499.500 415.600 ;
        RECT 495.200 413.200 496.400 414.000 ;
        RECT 497.200 413.700 499.500 414.300 ;
        RECT 495.600 412.400 496.200 413.200 ;
        RECT 497.200 412.800 498.000 413.700 ;
        RECT 495.600 411.600 496.400 412.400 ;
        RECT 498.800 412.200 499.600 412.400 ;
        RECT 500.600 412.200 501.200 415.800 ;
        RECT 506.800 415.800 508.600 416.400 ;
        RECT 511.600 415.800 513.400 416.400 ;
        RECT 502.000 412.800 502.800 414.400 ;
        RECT 505.200 413.600 506.000 415.200 ;
        RECT 503.600 412.300 504.400 412.400 ;
        RECT 506.800 412.300 507.600 415.800 ;
        RECT 510.000 413.600 510.800 415.200 ;
        RECT 503.600 412.200 507.600 412.300 ;
        RECT 498.800 411.600 501.200 412.200 ;
        RECT 502.800 411.700 507.600 412.200 ;
        RECT 502.800 411.600 504.400 411.700 ;
        RECT 493.800 410.400 496.200 411.000 ;
        RECT 457.200 409.700 463.400 410.200 ;
        RECT 457.200 409.600 458.000 409.700 ;
        RECT 462.000 409.600 463.400 409.700 ;
        RECT 464.000 409.600 465.000 410.200 ;
        RECT 468.400 409.600 469.800 410.200 ;
        RECT 470.400 409.600 471.400 410.200 ;
        RECT 462.800 408.400 463.400 409.600 ;
        RECT 462.800 407.600 463.600 408.400 ;
        RECT 464.200 406.400 465.000 409.600 ;
        RECT 469.200 408.400 469.800 409.600 ;
        RECT 469.200 407.600 470.000 408.400 ;
        RECT 464.200 405.600 466.000 406.400 ;
        RECT 464.200 402.200 465.000 405.600 ;
        RECT 470.600 404.400 471.400 409.600 ;
        RECT 474.800 409.600 477.200 410.200 ;
        RECT 478.800 409.600 480.800 410.200 ;
        RECT 470.600 403.600 472.400 404.400 ;
        RECT 470.600 402.200 471.400 403.600 ;
        RECT 474.800 402.200 475.600 409.600 ;
        RECT 476.400 409.400 477.200 409.600 ;
        RECT 479.200 402.200 480.800 409.600 ;
        RECT 483.000 409.600 485.200 410.200 ;
        RECT 486.000 409.600 487.400 410.200 ;
        RECT 488.000 409.600 489.000 410.200 ;
        RECT 483.000 409.400 483.800 409.600 ;
        RECT 484.400 402.200 485.200 409.600 ;
        RECT 486.800 408.400 487.400 409.600 ;
        RECT 486.800 407.600 487.600 408.400 ;
        RECT 488.200 404.400 489.000 409.600 ;
        RECT 488.200 403.600 490.000 404.400 ;
        RECT 488.200 402.200 489.000 403.600 ;
        RECT 492.400 402.200 493.200 410.200 ;
        RECT 495.600 406.200 496.200 410.400 ;
        RECT 499.000 410.200 499.600 411.600 ;
        RECT 502.800 411.200 503.600 411.600 ;
        RECT 495.600 402.200 496.400 406.200 ;
        RECT 498.800 402.200 499.600 410.200 ;
        RECT 500.400 409.600 504.400 410.200 ;
        RECT 500.400 402.200 501.200 409.600 ;
        RECT 503.600 402.200 504.400 409.600 ;
        RECT 506.800 402.200 507.600 411.700 ;
        RECT 508.400 410.300 509.200 410.400 ;
        RECT 511.600 410.300 512.400 415.800 ;
        RECT 518.400 414.200 519.200 419.800 ;
        RECT 521.200 415.600 522.000 417.200 ;
        RECT 522.800 416.300 523.600 419.800 ;
        RECT 526.000 417.600 526.800 419.800 ;
        RECT 524.400 416.300 525.200 417.200 ;
        RECT 522.800 415.700 525.200 416.300 ;
        RECT 518.400 413.800 520.200 414.200 ;
        RECT 518.600 413.600 520.200 413.800 ;
        RECT 516.400 411.600 518.000 412.400 ;
        RECT 508.400 409.700 512.400 410.300 ;
        RECT 508.400 408.800 509.200 409.700 ;
        RECT 511.600 402.200 512.400 409.700 ;
        RECT 513.200 408.800 514.000 410.400 ;
        RECT 514.800 409.600 515.600 411.200 ;
        RECT 519.600 410.400 520.200 413.600 ;
        RECT 519.600 409.600 520.400 410.400 ;
        RECT 521.200 410.300 522.000 410.400 ;
        RECT 522.800 410.300 523.600 415.700 ;
        RECT 524.400 415.600 525.200 415.700 ;
        RECT 526.200 414.400 526.800 417.600 ;
        RECT 526.000 413.600 526.800 414.400 ;
        RECT 521.200 409.700 523.600 410.300 ;
        RECT 526.200 410.200 526.800 413.600 ;
        RECT 529.200 415.800 530.000 419.800 ;
        RECT 532.400 417.800 533.200 419.800 ;
        RECT 529.200 412.400 529.800 415.800 ;
        RECT 532.400 415.600 533.000 417.800 ;
        RECT 534.000 415.600 534.800 417.200 ;
        RECT 535.600 415.800 536.400 419.800 ;
        RECT 540.000 418.400 541.600 419.800 ;
        RECT 540.000 417.600 542.800 418.400 ;
        RECT 540.000 416.200 541.600 417.600 ;
        RECT 530.600 415.000 533.000 415.600 ;
        RECT 527.600 412.300 528.400 412.400 ;
        RECT 529.200 412.300 530.000 412.400 ;
        RECT 527.600 411.700 530.000 412.300 ;
        RECT 527.600 410.800 528.400 411.700 ;
        RECT 529.200 411.600 530.000 411.700 ;
        RECT 530.600 412.000 531.200 415.000 ;
        RECT 532.200 413.600 533.200 414.400 ;
        RECT 534.100 414.300 534.700 415.600 ;
        RECT 535.600 415.200 538.200 415.800 ;
        RECT 537.400 415.000 538.200 415.200 ;
        RECT 538.800 414.800 540.400 415.600 ;
        RECT 535.600 414.300 537.200 414.400 ;
        RECT 534.100 414.200 537.200 414.300 ;
        RECT 541.000 414.200 541.600 416.200 ;
        RECT 545.200 415.800 546.000 419.800 ;
        RECT 546.800 416.000 547.600 419.800 ;
        RECT 550.000 416.000 550.800 419.800 ;
        RECT 546.800 415.800 550.800 416.000 ;
        RECT 551.600 415.800 552.400 419.800 ;
        RECT 553.200 416.000 554.000 419.800 ;
        RECT 556.400 416.000 557.200 419.800 ;
        RECT 553.200 415.800 557.200 416.000 ;
        RECT 558.000 415.800 558.800 419.800 ;
        RECT 559.600 415.800 560.400 419.800 ;
        RECT 564.000 418.400 565.600 419.800 ;
        RECT 564.000 417.600 566.800 418.400 ;
        RECT 564.000 416.200 565.600 417.600 ;
        RECT 542.200 414.800 543.000 415.600 ;
        RECT 543.600 415.200 546.000 415.800 ;
        RECT 547.000 415.400 550.600 415.800 ;
        RECT 543.600 415.000 544.400 415.200 ;
        RECT 534.100 414.000 537.800 414.200 ;
        RECT 534.100 413.700 540.000 414.000 ;
        RECT 535.600 413.600 540.000 413.700 ;
        RECT 532.000 412.800 532.800 413.600 ;
        RECT 537.200 413.400 540.000 413.600 ;
        RECT 539.200 413.200 540.000 413.400 ;
        RECT 540.600 413.600 541.600 414.200 ;
        RECT 542.400 414.400 543.000 414.800 ;
        RECT 547.600 414.400 548.400 414.800 ;
        RECT 551.600 414.400 552.200 415.800 ;
        RECT 553.400 415.400 557.000 415.800 ;
        RECT 554.000 414.400 554.800 414.800 ;
        RECT 558.000 414.400 558.600 415.800 ;
        RECT 559.600 415.200 562.200 415.800 ;
        RECT 561.400 415.000 562.200 415.200 ;
        RECT 562.800 414.800 564.400 415.600 ;
        RECT 542.400 413.600 543.200 414.400 ;
        RECT 544.400 413.600 546.000 414.400 ;
        RECT 546.800 413.800 548.400 414.400 ;
        RECT 546.800 413.600 547.600 413.800 ;
        RECT 549.800 413.600 552.400 414.400 ;
        RECT 553.200 413.800 554.800 414.400 ;
        RECT 556.200 414.300 558.800 414.400 ;
        RECT 559.600 414.300 561.200 414.400 ;
        RECT 556.200 414.200 561.200 414.300 ;
        RECT 565.000 414.200 565.600 416.200 ;
        RECT 569.200 415.800 570.000 419.800 ;
        RECT 573.400 416.400 574.200 419.800 ;
        RECT 566.200 414.800 567.000 415.600 ;
        RECT 567.600 415.200 570.000 415.800 ;
        RECT 572.400 415.800 574.200 416.400 ;
        RECT 567.600 415.000 568.400 415.200 ;
        RECT 556.200 414.000 561.800 414.200 ;
        RECT 553.200 413.600 554.000 413.800 ;
        RECT 556.200 413.700 564.000 414.000 ;
        RECT 556.200 413.600 558.800 413.700 ;
        RECT 559.600 413.600 564.000 413.700 ;
        RECT 540.600 412.400 541.200 413.600 ;
        RECT 537.800 412.200 538.600 412.400 ;
        RECT 529.200 410.200 529.800 411.600 ;
        RECT 530.600 411.400 531.400 412.000 ;
        RECT 537.800 411.600 539.400 412.200 ;
        RECT 540.400 411.600 541.200 412.400 ;
        RECT 545.200 412.300 546.000 412.400 ;
        RECT 548.400 412.300 549.200 413.200 ;
        RECT 545.200 411.700 549.200 412.300 ;
        RECT 545.200 411.600 546.000 411.700 ;
        RECT 548.400 411.600 549.200 411.700 ;
        RECT 538.600 411.400 539.400 411.600 ;
        RECT 530.600 411.200 534.800 411.400 ;
        RECT 530.800 410.800 534.800 411.200 ;
        RECT 521.200 409.600 522.000 409.700 ;
        RECT 518.000 407.600 518.800 409.200 ;
        RECT 519.600 407.000 520.200 409.600 ;
        RECT 516.600 406.400 520.200 407.000 ;
        RECT 516.400 402.200 517.200 406.400 ;
        RECT 519.600 406.200 520.200 406.400 ;
        RECT 519.600 402.200 520.400 406.200 ;
        RECT 522.800 402.200 523.600 409.700 ;
        RECT 526.000 409.400 527.800 410.200 ;
        RECT 529.200 409.600 530.600 410.200 ;
        RECT 527.000 402.200 527.800 409.400 ;
        RECT 529.800 404.400 530.600 409.600 ;
        RECT 529.200 403.600 530.600 404.400 ;
        RECT 529.800 402.200 530.600 403.600 ;
        RECT 534.000 402.200 534.800 410.800 ;
        RECT 540.600 410.200 541.200 411.600 ;
        RECT 549.800 410.200 550.400 413.600 ;
        RECT 554.800 411.600 555.600 413.200 ;
        RECT 551.600 410.200 552.400 410.400 ;
        RECT 556.200 410.200 556.800 413.600 ;
        RECT 561.200 413.400 564.000 413.600 ;
        RECT 563.200 413.200 564.000 413.400 ;
        RECT 564.600 413.600 565.600 414.200 ;
        RECT 566.400 414.400 567.000 414.800 ;
        RECT 566.400 413.600 567.200 414.400 ;
        RECT 568.400 413.600 570.000 414.400 ;
        RECT 570.800 413.600 571.600 415.200 ;
        RECT 564.600 412.400 565.200 413.600 ;
        RECT 561.800 412.200 562.600 412.400 ;
        RECT 561.800 411.600 563.400 412.200 ;
        RECT 564.400 411.600 565.200 412.400 ;
        RECT 562.600 411.400 563.400 411.600 ;
        RECT 558.000 410.200 558.800 410.400 ;
        RECT 564.600 410.200 565.200 411.600 ;
        RECT 535.600 409.600 538.200 410.200 ;
        RECT 535.600 402.200 536.400 409.600 ;
        RECT 537.400 409.400 538.200 409.600 ;
        RECT 540.000 402.200 541.600 410.200 ;
        RECT 543.600 409.600 546.000 410.200 ;
        RECT 543.600 409.400 544.400 409.600 ;
        RECT 545.200 402.200 546.000 409.600 ;
        RECT 549.400 409.600 550.400 410.200 ;
        RECT 551.000 409.600 552.400 410.200 ;
        RECT 555.800 409.600 556.800 410.200 ;
        RECT 557.400 409.600 558.800 410.200 ;
        RECT 559.600 409.600 562.200 410.200 ;
        RECT 549.400 404.400 550.200 409.600 ;
        RECT 551.000 408.400 551.600 409.600 ;
        RECT 550.800 407.600 551.600 408.400 ;
        RECT 548.400 403.600 550.200 404.400 ;
        RECT 549.400 402.200 550.200 403.600 ;
        RECT 555.800 402.200 556.600 409.600 ;
        RECT 557.400 408.400 558.000 409.600 ;
        RECT 557.200 407.600 558.000 408.400 ;
        RECT 559.600 402.200 560.400 409.600 ;
        RECT 561.400 409.400 562.200 409.600 ;
        RECT 564.000 402.200 565.600 410.200 ;
        RECT 567.600 409.600 570.000 410.200 ;
        RECT 567.600 409.400 568.400 409.600 ;
        RECT 569.200 402.200 570.000 409.600 ;
        RECT 572.400 402.200 573.200 415.800 ;
        RECT 575.600 413.800 576.400 419.800 ;
        RECT 582.000 416.600 582.800 419.800 ;
        RECT 583.600 417.000 584.400 419.800 ;
        RECT 585.200 417.000 586.000 419.800 ;
        RECT 586.800 417.000 587.600 419.800 ;
        RECT 590.000 417.000 590.800 419.800 ;
        RECT 593.200 417.000 594.000 419.800 ;
        RECT 594.800 417.000 595.600 419.800 ;
        RECT 596.400 417.000 597.200 419.800 ;
        RECT 598.000 417.000 598.800 419.800 ;
        RECT 580.200 415.800 582.800 416.600 ;
        RECT 599.600 416.600 600.400 419.800 ;
        RECT 586.200 415.800 590.800 416.400 ;
        RECT 580.200 415.200 581.000 415.800 ;
        RECT 578.000 414.400 581.000 415.200 ;
        RECT 575.600 413.000 584.400 413.800 ;
        RECT 586.200 413.400 587.000 415.800 ;
        RECT 590.000 415.600 590.800 415.800 ;
        RECT 591.600 415.600 593.200 416.400 ;
        RECT 596.200 415.600 597.200 416.400 ;
        RECT 599.600 415.800 602.000 416.600 ;
        RECT 588.400 413.600 589.200 415.200 ;
        RECT 590.000 414.800 590.800 415.000 ;
        RECT 590.000 414.200 594.400 414.800 ;
        RECT 593.600 414.000 594.400 414.200 ;
        RECT 574.000 408.800 574.800 410.400 ;
        RECT 575.600 407.400 576.400 413.000 ;
        RECT 585.000 412.600 587.000 413.400 ;
        RECT 590.800 412.600 594.000 413.400 ;
        RECT 596.400 412.800 597.200 415.600 ;
        RECT 601.200 415.200 602.000 415.800 ;
        RECT 601.200 414.600 603.000 415.200 ;
        RECT 602.200 413.400 603.000 414.600 ;
        RECT 606.000 414.600 606.800 419.800 ;
        RECT 607.600 416.000 608.400 419.800 ;
        RECT 607.600 415.200 608.600 416.000 ;
        RECT 606.000 414.000 607.200 414.600 ;
        RECT 602.200 412.600 606.000 413.400 ;
        RECT 577.000 412.000 577.800 412.200 ;
        RECT 578.800 412.000 579.600 412.400 ;
        RECT 582.000 412.000 582.800 412.400 ;
        RECT 599.600 412.000 600.400 412.600 ;
        RECT 606.600 412.000 607.200 414.000 ;
        RECT 577.000 411.400 600.400 412.000 ;
        RECT 606.400 411.400 607.200 412.000 ;
        RECT 606.400 409.600 607.000 411.400 ;
        RECT 607.800 410.800 608.600 415.200 ;
        RECT 585.200 409.400 586.000 409.600 ;
        RECT 580.600 409.000 586.000 409.400 ;
        RECT 579.800 408.800 586.000 409.000 ;
        RECT 587.000 409.000 595.600 409.600 ;
        RECT 577.200 408.000 578.800 408.800 ;
        RECT 579.800 408.200 581.200 408.800 ;
        RECT 587.000 408.200 587.600 409.000 ;
        RECT 594.800 408.800 595.600 409.000 ;
        RECT 598.000 409.000 607.000 409.600 ;
        RECT 598.000 408.800 598.800 409.000 ;
        RECT 578.200 407.600 578.800 408.000 ;
        RECT 581.800 407.600 587.600 408.200 ;
        RECT 588.200 407.600 590.800 408.400 ;
        RECT 575.600 406.800 577.600 407.400 ;
        RECT 578.200 406.800 582.400 407.600 ;
        RECT 577.000 406.200 577.600 406.800 ;
        RECT 577.000 405.600 578.000 406.200 ;
        RECT 577.200 402.200 578.000 405.600 ;
        RECT 580.400 402.200 581.200 406.800 ;
        RECT 583.600 402.200 584.400 405.000 ;
        RECT 585.200 402.200 586.000 405.000 ;
        RECT 586.800 402.200 587.600 407.000 ;
        RECT 590.000 402.200 590.800 407.000 ;
        RECT 593.200 402.200 594.000 408.400 ;
        RECT 601.200 407.600 603.800 408.400 ;
        RECT 596.400 406.800 600.600 407.600 ;
        RECT 594.800 402.200 595.600 405.000 ;
        RECT 596.400 402.200 597.200 405.000 ;
        RECT 598.000 402.200 598.800 405.000 ;
        RECT 601.200 402.200 602.000 407.600 ;
        RECT 606.400 407.400 607.000 409.000 ;
        RECT 604.400 406.800 607.000 407.400 ;
        RECT 607.600 410.000 608.600 410.800 ;
        RECT 604.400 402.200 605.200 406.800 ;
        RECT 607.600 402.200 608.400 410.000 ;
        RECT 2.800 396.400 3.600 399.800 ;
        RECT 2.600 395.800 3.600 396.400 ;
        RECT 2.600 395.200 3.200 395.800 ;
        RECT 6.000 395.200 6.800 399.800 ;
        RECT 9.200 397.000 10.000 399.800 ;
        RECT 10.800 397.000 11.600 399.800 ;
        RECT 1.200 394.600 3.200 395.200 ;
        RECT 1.200 389.000 2.000 394.600 ;
        RECT 3.800 394.400 8.000 395.200 ;
        RECT 12.400 395.000 13.200 399.800 ;
        RECT 15.600 395.000 16.400 399.800 ;
        RECT 3.800 394.000 4.400 394.400 ;
        RECT 2.800 393.200 4.400 394.000 ;
        RECT 7.400 393.800 13.200 394.400 ;
        RECT 5.400 393.200 6.800 393.800 ;
        RECT 5.400 393.000 11.600 393.200 ;
        RECT 6.200 392.600 11.600 393.000 ;
        RECT 10.800 392.400 11.600 392.600 ;
        RECT 12.600 393.000 13.200 393.800 ;
        RECT 13.800 393.600 16.400 394.400 ;
        RECT 18.800 393.600 19.600 399.800 ;
        RECT 20.400 397.000 21.200 399.800 ;
        RECT 22.000 397.000 22.800 399.800 ;
        RECT 23.600 397.000 24.400 399.800 ;
        RECT 22.000 394.400 26.200 395.200 ;
        RECT 26.800 394.400 27.600 399.800 ;
        RECT 30.000 395.200 30.800 399.800 ;
        RECT 30.000 394.600 32.600 395.200 ;
        RECT 26.800 393.600 29.400 394.400 ;
        RECT 20.400 393.000 21.200 393.200 ;
        RECT 12.600 392.400 21.200 393.000 ;
        RECT 23.600 393.000 24.400 393.200 ;
        RECT 32.000 393.000 32.600 394.600 ;
        RECT 23.600 392.400 32.600 393.000 ;
        RECT 32.000 390.600 32.600 392.400 ;
        RECT 33.200 392.000 34.000 399.800 ;
        RECT 33.200 391.200 34.200 392.000 ;
        RECT 36.400 391.600 37.200 394.400 ;
        RECT 2.600 390.000 26.000 390.600 ;
        RECT 32.000 390.000 32.800 390.600 ;
        RECT 2.600 389.800 3.400 390.000 ;
        RECT 7.600 389.600 8.400 390.000 ;
        RECT 25.200 389.400 26.000 390.000 ;
        RECT 1.200 388.200 10.000 389.000 ;
        RECT 10.600 388.600 12.600 389.400 ;
        RECT 16.400 388.600 19.600 389.400 ;
        RECT 1.200 382.200 2.000 388.200 ;
        RECT 3.600 386.800 6.600 387.600 ;
        RECT 5.800 386.200 6.600 386.800 ;
        RECT 11.800 386.200 12.600 388.600 ;
        RECT 14.000 386.800 14.800 388.400 ;
        RECT 19.200 387.800 20.000 388.000 ;
        RECT 15.600 387.200 20.000 387.800 ;
        RECT 15.600 387.000 16.400 387.200 ;
        RECT 22.000 386.400 22.800 389.200 ;
        RECT 27.800 388.600 31.600 389.400 ;
        RECT 27.800 387.400 28.600 388.600 ;
        RECT 32.200 388.000 32.800 390.000 ;
        RECT 15.600 386.200 16.400 386.400 ;
        RECT 5.800 385.400 8.400 386.200 ;
        RECT 11.800 385.600 16.400 386.200 ;
        RECT 17.200 385.600 18.800 386.400 ;
        RECT 21.800 385.600 22.800 386.400 ;
        RECT 26.800 386.800 28.600 387.400 ;
        RECT 31.600 387.400 32.800 388.000 ;
        RECT 26.800 386.200 27.600 386.800 ;
        RECT 7.600 382.200 8.400 385.400 ;
        RECT 25.200 385.400 27.600 386.200 ;
        RECT 9.200 382.200 10.000 385.000 ;
        RECT 10.800 382.200 11.600 385.000 ;
        RECT 12.400 382.200 13.200 385.000 ;
        RECT 15.600 382.200 16.400 385.000 ;
        RECT 18.800 382.200 19.600 385.000 ;
        RECT 20.400 382.200 21.200 385.000 ;
        RECT 22.000 382.200 22.800 385.000 ;
        RECT 23.600 382.200 24.400 385.000 ;
        RECT 25.200 382.200 26.000 385.400 ;
        RECT 31.600 382.200 32.400 387.400 ;
        RECT 33.400 386.800 34.200 391.200 ;
        RECT 33.200 386.300 34.200 386.800 ;
        RECT 34.800 386.300 35.600 386.400 ;
        RECT 33.200 385.700 35.600 386.300 ;
        RECT 38.000 386.200 38.800 399.800 ;
        RECT 42.800 392.800 43.600 399.800 ;
        RECT 42.600 391.800 43.600 392.800 ;
        RECT 46.000 392.400 46.800 399.800 ;
        RECT 44.200 391.800 46.800 392.400 ;
        RECT 42.600 388.400 43.200 391.800 ;
        RECT 44.200 389.800 44.800 391.800 ;
        RECT 47.600 391.400 48.400 399.800 ;
        RECT 52.000 396.400 52.800 399.800 ;
        RECT 50.800 395.800 52.800 396.400 ;
        RECT 56.400 395.800 57.200 399.800 ;
        RECT 60.600 395.800 61.800 399.800 ;
        RECT 50.800 395.000 51.600 395.800 ;
        RECT 56.400 395.200 57.000 395.800 ;
        RECT 54.200 394.600 57.800 395.200 ;
        RECT 60.400 395.000 61.200 395.800 ;
        RECT 54.200 394.400 55.000 394.600 ;
        RECT 57.000 394.400 57.800 394.600 ;
        RECT 50.800 393.000 51.600 393.200 ;
        RECT 55.400 393.000 56.200 393.200 ;
        RECT 50.800 392.400 56.200 393.000 ;
        RECT 56.800 393.000 59.000 393.600 ;
        RECT 56.800 391.800 57.400 393.000 ;
        RECT 58.200 392.800 59.000 393.000 ;
        RECT 60.600 393.200 62.000 394.000 ;
        RECT 60.600 392.200 61.200 393.200 ;
        RECT 52.600 391.400 57.400 391.800 ;
        RECT 47.600 391.200 57.400 391.400 ;
        RECT 58.800 391.600 61.200 392.200 ;
        RECT 47.600 391.000 53.400 391.200 ;
        RECT 47.600 390.800 53.200 391.000 ;
        RECT 43.800 389.000 44.800 389.800 ;
        RECT 39.600 386.800 40.400 388.400 ;
        RECT 42.600 387.600 43.600 388.400 ;
        RECT 33.200 382.200 34.000 385.700 ;
        RECT 34.800 385.600 35.600 385.700 ;
        RECT 37.000 385.600 38.800 386.200 ;
        RECT 42.600 386.200 43.200 387.600 ;
        RECT 44.200 387.400 44.800 389.000 ;
        RECT 45.800 389.600 46.800 390.400 ;
        RECT 54.000 390.200 54.800 390.400 ;
        RECT 49.800 389.600 54.800 390.200 ;
        RECT 57.200 390.300 58.000 390.400 ;
        RECT 58.800 390.300 59.400 391.600 ;
        RECT 65.200 391.200 66.000 399.800 ;
        RECT 66.800 392.400 67.600 399.800 ;
        RECT 70.000 392.800 70.800 399.800 ;
        RECT 74.000 393.600 74.800 394.400 ;
        RECT 66.800 391.800 69.400 392.400 ;
        RECT 70.000 391.800 71.000 392.800 ;
        RECT 74.000 392.400 74.600 393.600 ;
        RECT 75.400 392.400 76.200 399.800 ;
        RECT 83.400 392.800 84.200 399.800 ;
        RECT 87.600 395.000 88.400 399.000 ;
        RECT 93.000 398.400 93.800 399.800 ;
        RECT 92.400 397.600 93.800 398.400 ;
        RECT 61.800 390.600 66.000 391.200 ;
        RECT 61.800 390.400 62.600 390.600 ;
        RECT 57.200 389.700 59.500 390.300 ;
        RECT 63.400 389.800 64.200 390.000 ;
        RECT 57.200 389.600 58.000 389.700 ;
        RECT 45.800 388.800 46.600 389.600 ;
        RECT 49.800 389.400 50.600 389.600 ;
        RECT 51.400 388.400 52.200 388.600 ;
        RECT 58.800 388.400 59.400 389.700 ;
        RECT 60.400 389.200 64.200 389.800 ;
        RECT 60.400 389.000 61.200 389.200 ;
        RECT 48.400 387.800 59.400 388.400 ;
        RECT 48.400 387.600 50.000 387.800 ;
        RECT 44.200 386.800 46.800 387.400 ;
        RECT 42.600 385.600 43.600 386.200 ;
        RECT 37.000 384.400 37.800 385.600 ;
        RECT 37.000 383.600 38.800 384.400 ;
        RECT 37.000 382.200 37.800 383.600 ;
        RECT 42.800 382.200 43.600 385.600 ;
        RECT 46.000 382.200 46.800 386.800 ;
        RECT 47.600 382.200 48.400 387.000 ;
        RECT 52.600 385.600 53.200 387.800 ;
        RECT 58.200 387.600 59.000 387.800 ;
        RECT 65.200 387.200 66.000 390.600 ;
        RECT 66.800 389.600 67.800 390.400 ;
        RECT 67.000 388.800 67.800 389.600 ;
        RECT 68.800 389.800 69.400 391.800 ;
        RECT 68.800 389.000 69.800 389.800 ;
        RECT 68.800 387.400 69.400 389.000 ;
        RECT 70.400 388.400 71.000 391.800 ;
        RECT 73.200 391.800 74.600 392.400 ;
        RECT 75.200 391.800 76.200 392.400 ;
        RECT 82.600 392.200 84.200 392.800 ;
        RECT 73.200 391.600 74.000 391.800 ;
        RECT 75.200 390.400 75.800 391.800 ;
        RECT 74.800 389.600 75.800 390.400 ;
        RECT 75.200 388.400 75.800 389.600 ;
        RECT 76.400 390.300 77.200 390.400 ;
        RECT 79.600 390.300 80.400 390.400 ;
        RECT 76.400 389.700 80.400 390.300 ;
        RECT 76.400 388.800 77.200 389.700 ;
        RECT 79.600 389.600 80.400 389.700 ;
        RECT 81.200 389.600 82.000 391.200 ;
        RECT 82.600 388.400 83.200 392.200 ;
        RECT 87.800 391.600 88.400 395.000 ;
        RECT 93.000 392.800 93.800 397.600 ;
        RECT 97.200 395.000 98.000 399.000 ;
        RECT 84.600 391.000 88.400 391.600 ;
        RECT 92.200 392.200 93.800 392.800 ;
        RECT 84.600 389.000 85.200 391.000 ;
        RECT 70.000 387.600 71.000 388.400 ;
        RECT 73.200 387.600 75.800 388.400 ;
        RECT 78.000 388.200 78.800 388.400 ;
        RECT 77.200 387.600 78.800 388.200 ;
        RECT 81.200 387.600 83.200 388.400 ;
        RECT 83.800 388.200 85.200 389.000 ;
        RECT 86.000 388.800 86.800 390.400 ;
        RECT 87.600 390.300 88.400 390.400 ;
        RECT 89.200 390.300 90.000 390.400 ;
        RECT 87.600 389.700 90.000 390.300 ;
        RECT 87.600 388.800 88.400 389.700 ;
        RECT 89.200 389.600 90.000 389.700 ;
        RECT 90.800 389.600 91.600 391.200 ;
        RECT 92.200 388.400 92.800 392.200 ;
        RECT 97.400 391.600 98.000 395.000 ;
        RECT 94.200 391.000 98.000 391.600 ;
        RECT 94.200 389.000 94.800 391.000 ;
        RECT 62.200 386.600 66.000 387.200 ;
        RECT 62.200 386.400 63.000 386.600 ;
        RECT 50.800 384.200 51.600 385.000 ;
        RECT 52.400 384.800 53.200 385.600 ;
        RECT 54.200 385.400 55.000 385.600 ;
        RECT 54.200 384.800 57.000 385.400 ;
        RECT 56.400 384.200 57.000 384.800 ;
        RECT 60.400 384.200 61.200 385.000 ;
        RECT 50.800 383.600 52.800 384.200 ;
        RECT 52.000 382.200 52.800 383.600 ;
        RECT 56.400 382.200 57.200 384.200 ;
        RECT 60.400 383.600 61.800 384.200 ;
        RECT 60.600 382.200 61.800 383.600 ;
        RECT 65.200 382.200 66.000 386.600 ;
        RECT 66.800 386.800 69.400 387.400 ;
        RECT 66.800 382.200 67.600 386.800 ;
        RECT 70.400 386.200 71.000 387.600 ;
        RECT 73.400 386.200 74.000 387.600 ;
        RECT 77.200 387.200 78.000 387.600 ;
        RECT 82.600 387.000 83.200 387.600 ;
        RECT 84.200 387.800 85.200 388.200 ;
        RECT 84.200 387.200 88.400 387.800 ;
        RECT 90.800 387.600 92.800 388.400 ;
        RECT 93.400 388.200 94.800 389.000 ;
        RECT 95.600 388.800 96.400 390.400 ;
        RECT 97.200 388.800 98.000 390.400 ;
        RECT 82.600 386.600 83.400 387.000 ;
        RECT 75.000 386.200 78.600 386.600 ;
        RECT 70.000 385.600 71.000 386.200 ;
        RECT 70.000 382.200 70.800 385.600 ;
        RECT 73.200 382.200 74.000 386.200 ;
        RECT 74.800 386.000 78.800 386.200 ;
        RECT 82.600 386.000 84.200 386.600 ;
        RECT 74.800 382.200 75.600 386.000 ;
        RECT 78.000 382.200 78.800 386.000 ;
        RECT 83.400 384.400 84.200 386.000 ;
        RECT 87.800 385.000 88.400 387.200 ;
        RECT 92.200 387.000 92.800 387.600 ;
        RECT 93.800 387.800 94.800 388.200 ;
        RECT 93.800 387.200 98.000 387.800 ;
        RECT 92.200 386.600 93.000 387.000 ;
        RECT 92.200 386.000 93.800 386.600 ;
        RECT 82.800 383.600 84.200 384.400 ;
        RECT 83.400 383.000 84.200 383.600 ;
        RECT 87.600 383.000 88.400 385.000 ;
        RECT 93.000 383.000 93.800 386.000 ;
        RECT 97.400 385.000 98.000 387.200 ;
        RECT 97.200 383.000 98.000 385.000 ;
        RECT 98.800 382.200 99.600 399.800 ;
        RECT 103.600 392.800 104.400 399.800 ;
        RECT 103.400 391.800 104.400 392.800 ;
        RECT 106.800 392.400 107.600 399.800 ;
        RECT 105.000 391.800 107.600 392.400 ;
        RECT 109.000 392.600 109.800 399.800 ;
        RECT 109.000 391.800 110.800 392.600 ;
        RECT 103.400 388.400 104.000 391.800 ;
        RECT 105.000 389.800 105.600 391.800 ;
        RECT 104.600 389.000 105.600 389.800 ;
        RECT 103.400 387.600 104.400 388.400 ;
        RECT 100.400 384.800 101.200 386.400 ;
        RECT 103.400 386.200 104.000 387.600 ;
        RECT 105.000 387.400 105.600 389.000 ;
        RECT 106.600 389.600 107.600 390.400 ;
        RECT 108.400 389.600 109.200 391.200 ;
        RECT 110.000 390.300 110.600 391.800 ;
        RECT 113.200 391.400 114.000 399.800 ;
        RECT 117.600 396.400 118.400 399.800 ;
        RECT 116.400 395.800 118.400 396.400 ;
        RECT 122.000 395.800 122.800 399.800 ;
        RECT 126.200 395.800 127.400 399.800 ;
        RECT 116.400 395.000 117.200 395.800 ;
        RECT 122.000 395.200 122.600 395.800 ;
        RECT 119.800 394.600 123.400 395.200 ;
        RECT 126.000 395.000 126.800 395.800 ;
        RECT 119.800 394.400 120.600 394.600 ;
        RECT 122.600 394.400 123.400 394.600 ;
        RECT 116.400 393.000 117.200 393.200 ;
        RECT 121.000 393.000 121.800 393.200 ;
        RECT 116.400 392.400 121.800 393.000 ;
        RECT 122.400 393.000 124.600 393.600 ;
        RECT 122.400 391.800 123.000 393.000 ;
        RECT 123.800 392.800 124.600 393.000 ;
        RECT 126.200 393.200 127.600 394.000 ;
        RECT 126.200 392.200 126.800 393.200 ;
        RECT 118.200 391.400 123.000 391.800 ;
        RECT 113.200 391.200 123.000 391.400 ;
        RECT 124.400 391.600 126.800 392.200 ;
        RECT 113.200 391.000 119.000 391.200 ;
        RECT 113.200 390.800 118.800 391.000 ;
        RECT 111.600 390.300 112.400 390.400 ;
        RECT 110.000 389.700 112.400 390.300 ;
        RECT 119.600 390.200 120.400 390.400 ;
        RECT 106.600 388.800 107.400 389.600 ;
        RECT 110.000 388.400 110.600 389.700 ;
        RECT 111.600 389.600 112.400 389.700 ;
        RECT 115.400 389.600 120.400 390.200 ;
        RECT 115.400 389.400 116.200 389.600 ;
        RECT 117.000 388.400 117.800 388.600 ;
        RECT 124.400 388.400 125.000 391.600 ;
        RECT 130.800 391.200 131.600 399.800 ;
        RECT 135.000 392.400 135.800 399.800 ;
        RECT 136.400 393.600 137.200 394.400 ;
        RECT 136.600 392.400 137.200 393.600 ;
        RECT 139.600 393.600 140.400 394.400 ;
        RECT 139.600 392.400 140.200 393.600 ;
        RECT 141.000 392.400 141.800 399.800 ;
        RECT 146.800 392.800 147.600 399.800 ;
        RECT 135.000 391.800 136.000 392.400 ;
        RECT 136.600 391.800 138.000 392.400 ;
        RECT 127.400 390.600 131.600 391.200 ;
        RECT 127.400 390.400 128.200 390.600 ;
        RECT 129.000 389.800 129.800 390.000 ;
        RECT 126.000 389.200 129.800 389.800 ;
        RECT 126.000 389.000 126.800 389.200 ;
        RECT 110.000 387.600 110.800 388.400 ;
        RECT 114.000 387.800 125.000 388.400 ;
        RECT 114.000 387.600 115.600 387.800 ;
        RECT 105.000 386.800 107.600 387.400 ;
        RECT 103.400 385.600 104.400 386.200 ;
        RECT 103.600 382.200 104.400 385.600 ;
        RECT 106.800 382.200 107.600 386.800 ;
        RECT 110.000 384.200 110.600 387.600 ;
        RECT 111.600 384.800 112.400 386.400 ;
        RECT 110.000 382.200 110.800 384.200 ;
        RECT 113.200 382.200 114.000 387.000 ;
        RECT 118.200 385.600 118.800 387.800 ;
        RECT 121.200 387.600 122.000 387.800 ;
        RECT 123.800 387.600 124.600 387.800 ;
        RECT 130.800 387.200 131.600 390.600 ;
        RECT 134.000 388.800 134.800 390.400 ;
        RECT 135.400 390.300 136.000 391.800 ;
        RECT 137.200 391.600 138.000 391.800 ;
        RECT 138.800 391.800 140.200 392.400 ;
        RECT 140.800 391.800 141.800 392.400 ;
        RECT 146.600 391.800 147.600 392.800 ;
        RECT 150.000 392.400 150.800 399.800 ;
        RECT 148.200 391.800 150.800 392.400 ;
        RECT 138.800 391.600 139.600 391.800 ;
        RECT 138.900 390.300 139.500 391.600 ;
        RECT 135.400 389.700 139.500 390.300 ;
        RECT 135.400 388.400 136.000 389.700 ;
        RECT 140.800 388.400 141.400 391.800 ;
        RECT 142.000 388.800 142.800 390.400 ;
        RECT 146.600 388.400 147.200 391.800 ;
        RECT 148.200 389.800 148.800 391.800 ;
        RECT 147.800 389.000 148.800 389.800 ;
        RECT 132.400 388.200 133.200 388.400 ;
        RECT 132.400 387.600 134.000 388.200 ;
        RECT 135.400 387.600 138.000 388.400 ;
        RECT 138.800 387.600 141.400 388.400 ;
        RECT 143.600 388.300 144.400 388.400 ;
        RECT 146.600 388.300 147.600 388.400 ;
        RECT 143.600 388.200 147.600 388.300 ;
        RECT 142.800 387.700 147.600 388.200 ;
        RECT 142.800 387.600 144.400 387.700 ;
        RECT 146.600 387.600 147.600 387.700 ;
        RECT 133.200 387.200 134.000 387.600 ;
        RECT 127.800 386.600 131.600 387.200 ;
        RECT 127.800 386.400 128.600 386.600 ;
        RECT 116.400 384.200 117.200 385.000 ;
        RECT 118.000 384.800 118.800 385.600 ;
        RECT 119.800 385.400 120.600 385.600 ;
        RECT 119.800 384.800 122.600 385.400 ;
        RECT 122.000 384.200 122.600 384.800 ;
        RECT 126.000 384.200 126.800 385.000 ;
        RECT 116.400 383.600 118.400 384.200 ;
        RECT 117.600 382.200 118.400 383.600 ;
        RECT 122.000 382.200 122.800 384.200 ;
        RECT 126.000 383.600 127.400 384.200 ;
        RECT 126.200 382.200 127.400 383.600 ;
        RECT 130.800 382.200 131.600 386.600 ;
        RECT 132.600 386.200 136.200 386.600 ;
        RECT 137.200 386.200 137.800 387.600 ;
        RECT 139.000 386.200 139.600 387.600 ;
        RECT 142.800 387.200 143.600 387.600 ;
        RECT 140.600 386.200 144.200 386.600 ;
        RECT 146.600 386.200 147.200 387.600 ;
        RECT 148.200 387.400 148.800 389.000 ;
        RECT 149.800 390.300 150.800 390.400 ;
        RECT 156.400 390.300 157.200 390.400 ;
        RECT 149.800 389.700 157.200 390.300 ;
        RECT 149.800 389.600 150.800 389.700 ;
        RECT 156.400 389.600 157.200 389.700 ;
        RECT 149.800 388.800 150.600 389.600 ;
        RECT 148.200 386.800 150.800 387.400 ;
        RECT 132.400 386.000 136.400 386.200 ;
        RECT 132.400 382.200 133.200 386.000 ;
        RECT 135.600 382.200 136.400 386.000 ;
        RECT 137.200 382.200 138.000 386.200 ;
        RECT 138.800 382.200 139.600 386.200 ;
        RECT 140.400 386.000 144.400 386.200 ;
        RECT 140.400 382.200 141.200 386.000 ;
        RECT 143.600 382.200 144.400 386.000 ;
        RECT 146.600 385.600 147.600 386.200 ;
        RECT 146.800 382.200 147.600 385.600 ;
        RECT 150.000 382.200 150.800 386.800 ;
        RECT 151.600 386.300 152.400 386.400 ;
        RECT 156.400 386.300 157.200 386.400 ;
        RECT 151.600 385.700 157.200 386.300 ;
        RECT 151.600 385.600 152.400 385.700 ;
        RECT 156.400 384.800 157.200 385.700 ;
        RECT 158.000 382.200 158.800 399.800 ;
        RECT 161.200 392.800 162.000 399.800 ;
        RECT 161.000 391.800 162.000 392.800 ;
        RECT 164.400 392.400 165.200 399.800 ;
        RECT 162.600 391.800 165.200 392.400 ;
        RECT 167.600 392.000 168.400 399.800 ;
        RECT 170.800 395.200 171.600 399.800 ;
        RECT 161.000 388.400 161.600 391.800 ;
        RECT 162.600 389.800 163.200 391.800 ;
        RECT 167.400 391.200 168.400 392.000 ;
        RECT 169.000 394.600 171.600 395.200 ;
        RECT 169.000 393.000 169.600 394.600 ;
        RECT 174.000 394.400 174.800 399.800 ;
        RECT 177.200 397.000 178.000 399.800 ;
        RECT 178.800 397.000 179.600 399.800 ;
        RECT 180.400 397.000 181.200 399.800 ;
        RECT 175.400 394.400 179.600 395.200 ;
        RECT 172.200 393.600 174.800 394.400 ;
        RECT 182.000 393.600 182.800 399.800 ;
        RECT 185.200 395.000 186.000 399.800 ;
        RECT 188.400 395.000 189.200 399.800 ;
        RECT 190.000 397.000 190.800 399.800 ;
        RECT 191.600 397.000 192.400 399.800 ;
        RECT 194.800 395.200 195.600 399.800 ;
        RECT 198.000 396.400 198.800 399.800 ;
        RECT 198.000 395.800 199.000 396.400 ;
        RECT 198.400 395.200 199.000 395.800 ;
        RECT 193.600 394.400 197.800 395.200 ;
        RECT 198.400 394.600 200.400 395.200 ;
        RECT 185.200 393.600 187.800 394.400 ;
        RECT 188.400 393.800 194.200 394.400 ;
        RECT 197.200 394.000 197.800 394.400 ;
        RECT 177.200 393.000 178.000 393.200 ;
        RECT 169.000 392.400 178.000 393.000 ;
        RECT 180.400 393.000 181.200 393.200 ;
        RECT 188.400 393.000 189.000 393.800 ;
        RECT 194.800 393.200 196.200 393.800 ;
        RECT 197.200 393.200 198.800 394.000 ;
        RECT 180.400 392.400 189.000 393.000 ;
        RECT 190.000 393.000 196.200 393.200 ;
        RECT 190.000 392.600 195.400 393.000 ;
        RECT 190.000 392.400 190.800 392.600 ;
        RECT 162.200 389.000 163.200 389.800 ;
        RECT 161.000 387.600 162.000 388.400 ;
        RECT 161.000 386.200 161.600 387.600 ;
        RECT 162.600 387.400 163.200 389.000 ;
        RECT 164.200 390.300 165.200 390.400 ;
        RECT 167.400 390.300 168.200 391.200 ;
        RECT 169.000 390.600 169.600 392.400 ;
        RECT 164.200 389.700 168.200 390.300 ;
        RECT 164.200 389.600 165.200 389.700 ;
        RECT 164.200 388.800 165.000 389.600 ;
        RECT 162.600 386.800 165.200 387.400 ;
        RECT 161.000 385.600 162.000 386.200 ;
        RECT 161.200 382.200 162.000 385.600 ;
        RECT 164.400 382.200 165.200 386.800 ;
        RECT 167.400 386.800 168.200 389.700 ;
        RECT 168.800 390.000 169.600 390.600 ;
        RECT 175.600 390.000 199.000 390.600 ;
        RECT 168.800 388.000 169.400 390.000 ;
        RECT 175.600 389.400 176.400 390.000 ;
        RECT 193.200 389.600 194.000 390.000 ;
        RECT 194.800 389.600 195.600 390.000 ;
        RECT 196.400 389.600 197.200 390.000 ;
        RECT 198.200 389.800 199.000 390.000 ;
        RECT 170.000 388.600 173.800 389.400 ;
        RECT 168.800 387.400 170.000 388.000 ;
        RECT 167.400 386.000 168.400 386.800 ;
        RECT 167.600 382.200 168.400 386.000 ;
        RECT 169.200 382.200 170.000 387.400 ;
        RECT 173.000 387.400 173.800 388.600 ;
        RECT 173.000 386.800 174.800 387.400 ;
        RECT 174.000 386.200 174.800 386.800 ;
        RECT 178.800 386.400 179.600 389.200 ;
        RECT 182.000 388.600 185.200 389.400 ;
        RECT 189.000 388.600 191.000 389.400 ;
        RECT 199.600 389.000 200.400 394.600 ;
        RECT 181.600 387.800 182.400 388.000 ;
        RECT 181.600 387.200 186.000 387.800 ;
        RECT 185.200 387.000 186.000 387.200 ;
        RECT 186.800 386.800 187.600 388.400 ;
        RECT 174.000 385.400 176.400 386.200 ;
        RECT 178.800 385.600 179.800 386.400 ;
        RECT 182.800 385.600 184.400 386.400 ;
        RECT 185.200 386.200 186.000 386.400 ;
        RECT 189.000 386.200 189.800 388.600 ;
        RECT 191.600 388.200 200.400 389.000 ;
        RECT 195.000 386.800 198.000 387.600 ;
        RECT 195.000 386.200 195.800 386.800 ;
        RECT 185.200 385.600 189.800 386.200 ;
        RECT 175.600 382.200 176.400 385.400 ;
        RECT 193.200 385.400 195.800 386.200 ;
        RECT 177.200 382.200 178.000 385.000 ;
        RECT 178.800 382.200 179.600 385.000 ;
        RECT 180.400 382.200 181.200 385.000 ;
        RECT 182.000 382.200 182.800 385.000 ;
        RECT 185.200 382.200 186.000 385.000 ;
        RECT 188.400 382.200 189.200 385.000 ;
        RECT 190.000 382.200 190.800 385.000 ;
        RECT 191.600 382.200 192.400 385.000 ;
        RECT 193.200 382.200 194.000 385.400 ;
        RECT 199.600 382.200 200.400 388.200 ;
        RECT 201.200 384.800 202.000 386.400 ;
        RECT 202.800 382.200 203.600 399.800 ;
        RECT 204.400 391.600 205.200 393.200 ;
        RECT 206.000 386.200 206.800 399.800 ;
        RECT 209.200 391.600 210.000 393.200 ;
        RECT 207.600 386.800 208.400 388.400 ;
        RECT 210.800 386.200 211.600 399.800 ;
        RECT 215.600 396.400 216.400 399.800 ;
        RECT 215.400 395.800 216.400 396.400 ;
        RECT 215.400 395.200 216.000 395.800 ;
        RECT 218.800 395.200 219.600 399.800 ;
        RECT 222.000 397.000 222.800 399.800 ;
        RECT 223.600 397.000 224.400 399.800 ;
        RECT 214.000 394.600 216.000 395.200 ;
        RECT 214.000 389.000 214.800 394.600 ;
        RECT 216.600 394.400 220.800 395.200 ;
        RECT 225.200 395.000 226.000 399.800 ;
        RECT 228.400 395.000 229.200 399.800 ;
        RECT 216.600 394.000 217.200 394.400 ;
        RECT 215.600 393.200 217.200 394.000 ;
        RECT 220.200 393.800 226.000 394.400 ;
        RECT 218.200 393.200 219.600 393.800 ;
        RECT 218.200 393.000 224.400 393.200 ;
        RECT 219.000 392.600 224.400 393.000 ;
        RECT 223.600 392.400 224.400 392.600 ;
        RECT 225.400 393.000 226.000 393.800 ;
        RECT 226.600 393.600 229.200 394.400 ;
        RECT 231.600 393.600 232.400 399.800 ;
        RECT 233.200 397.000 234.000 399.800 ;
        RECT 234.800 397.000 235.600 399.800 ;
        RECT 236.400 397.000 237.200 399.800 ;
        RECT 234.800 394.400 239.000 395.200 ;
        RECT 239.600 394.400 240.400 399.800 ;
        RECT 242.800 395.200 243.600 399.800 ;
        RECT 242.800 394.600 245.400 395.200 ;
        RECT 239.600 393.600 242.200 394.400 ;
        RECT 233.200 393.000 234.000 393.200 ;
        RECT 225.400 392.400 234.000 393.000 ;
        RECT 236.400 393.000 237.200 393.200 ;
        RECT 244.800 393.000 245.400 394.600 ;
        RECT 236.400 392.400 245.400 393.000 ;
        RECT 244.800 390.600 245.400 392.400 ;
        RECT 246.000 392.000 246.800 399.800 ;
        RECT 246.000 391.200 247.000 392.000 ;
        RECT 215.400 390.000 238.800 390.600 ;
        RECT 244.800 390.000 245.600 390.600 ;
        RECT 215.400 389.800 216.200 390.000 ;
        RECT 217.200 389.600 218.000 390.000 ;
        RECT 220.400 389.600 221.200 390.000 ;
        RECT 238.000 389.400 238.800 390.000 ;
        RECT 212.400 386.800 213.200 388.400 ;
        RECT 214.000 388.200 222.800 389.000 ;
        RECT 223.400 388.600 225.400 389.400 ;
        RECT 229.200 388.600 232.400 389.400 ;
        RECT 205.000 385.600 206.800 386.200 ;
        RECT 209.800 385.600 211.600 386.200 ;
        RECT 205.000 384.400 205.800 385.600 ;
        RECT 204.400 383.600 205.800 384.400 ;
        RECT 205.000 382.200 205.800 383.600 ;
        RECT 209.800 382.200 210.600 385.600 ;
        RECT 214.000 382.200 214.800 388.200 ;
        RECT 216.400 386.800 219.400 387.600 ;
        RECT 218.600 386.200 219.400 386.800 ;
        RECT 224.600 386.200 225.400 388.600 ;
        RECT 226.800 386.800 227.600 388.400 ;
        RECT 232.000 387.800 232.800 388.000 ;
        RECT 228.400 387.200 232.800 387.800 ;
        RECT 228.400 387.000 229.200 387.200 ;
        RECT 234.800 386.400 235.600 389.200 ;
        RECT 240.600 388.600 244.400 389.400 ;
        RECT 240.600 387.400 241.400 388.600 ;
        RECT 245.000 388.000 245.600 390.000 ;
        RECT 228.400 386.200 229.200 386.400 ;
        RECT 218.600 385.400 221.200 386.200 ;
        RECT 224.600 385.600 229.200 386.200 ;
        RECT 230.000 385.600 231.600 386.400 ;
        RECT 234.600 385.600 235.600 386.400 ;
        RECT 239.600 386.800 241.400 387.400 ;
        RECT 244.400 387.400 245.600 388.000 ;
        RECT 239.600 386.200 240.400 386.800 ;
        RECT 220.400 382.200 221.200 385.400 ;
        RECT 238.000 385.400 240.400 386.200 ;
        RECT 222.000 382.200 222.800 385.000 ;
        RECT 223.600 382.200 224.400 385.000 ;
        RECT 225.200 382.200 226.000 385.000 ;
        RECT 228.400 382.200 229.200 385.000 ;
        RECT 231.600 382.200 232.400 385.000 ;
        RECT 233.200 382.200 234.000 385.000 ;
        RECT 234.800 382.200 235.600 385.000 ;
        RECT 236.400 382.200 237.200 385.000 ;
        RECT 238.000 382.200 238.800 385.400 ;
        RECT 244.400 382.200 245.200 387.400 ;
        RECT 246.200 386.800 247.000 391.200 ;
        RECT 249.200 386.800 250.000 388.400 ;
        RECT 246.000 386.000 247.000 386.800 ;
        RECT 250.800 386.200 251.600 399.800 ;
        RECT 254.000 393.600 255.600 394.400 ;
        RECT 252.400 391.600 253.200 393.200 ;
        RECT 254.800 392.400 255.400 393.600 ;
        RECT 256.200 392.400 257.000 399.800 ;
        RECT 254.000 391.800 255.400 392.400 ;
        RECT 256.000 391.800 257.000 392.400 ;
        RECT 260.400 391.800 261.200 399.800 ;
        RECT 263.600 392.400 264.400 399.800 ;
        RECT 266.800 396.400 267.600 399.800 ;
        RECT 266.600 395.800 267.600 396.400 ;
        RECT 266.600 395.200 267.200 395.800 ;
        RECT 270.000 395.200 270.800 399.800 ;
        RECT 273.200 397.000 274.000 399.800 ;
        RECT 274.800 397.000 275.600 399.800 ;
        RECT 262.200 391.800 264.400 392.400 ;
        RECT 265.200 394.600 267.200 395.200 ;
        RECT 254.000 391.600 254.800 391.800 ;
        RECT 252.400 390.300 253.200 390.400 ;
        RECT 256.000 390.300 256.600 391.800 ;
        RECT 252.400 389.700 256.600 390.300 ;
        RECT 252.400 389.600 253.200 389.700 ;
        RECT 256.000 388.400 256.600 389.700 ;
        RECT 257.200 388.800 258.000 390.400 ;
        RECT 260.400 389.600 261.000 391.800 ;
        RECT 262.200 391.200 262.800 391.800 ;
        RECT 261.600 390.400 262.800 391.200 ;
        RECT 254.000 387.600 256.600 388.400 ;
        RECT 258.800 388.300 259.600 388.400 ;
        RECT 260.400 388.300 261.200 389.600 ;
        RECT 258.800 388.200 261.200 388.300 ;
        RECT 258.000 387.700 261.200 388.200 ;
        RECT 258.000 387.600 259.600 387.700 ;
        RECT 254.200 386.200 254.800 387.600 ;
        RECT 258.000 387.200 258.800 387.600 ;
        RECT 255.800 386.200 259.400 386.600 ;
        RECT 246.000 382.200 246.800 386.000 ;
        RECT 250.800 385.600 252.600 386.200 ;
        RECT 251.800 384.400 252.600 385.600 ;
        RECT 251.800 383.600 253.200 384.400 ;
        RECT 251.800 382.200 252.600 383.600 ;
        RECT 254.000 382.200 254.800 386.200 ;
        RECT 255.600 386.000 259.600 386.200 ;
        RECT 255.600 382.200 256.400 386.000 ;
        RECT 258.800 382.200 259.600 386.000 ;
        RECT 260.400 382.200 261.200 387.700 ;
        RECT 262.200 387.400 262.800 390.400 ;
        RECT 263.600 388.800 264.400 390.400 ;
        RECT 265.200 389.000 266.000 394.600 ;
        RECT 267.800 394.400 272.000 395.200 ;
        RECT 276.400 395.000 277.200 399.800 ;
        RECT 279.600 395.000 280.400 399.800 ;
        RECT 267.800 394.000 268.400 394.400 ;
        RECT 266.800 393.200 268.400 394.000 ;
        RECT 271.400 393.800 277.200 394.400 ;
        RECT 269.400 393.200 270.800 393.800 ;
        RECT 269.400 393.000 275.600 393.200 ;
        RECT 270.200 392.600 275.600 393.000 ;
        RECT 274.800 392.400 275.600 392.600 ;
        RECT 276.600 393.000 277.200 393.800 ;
        RECT 277.800 393.600 280.400 394.400 ;
        RECT 282.800 393.600 283.600 399.800 ;
        RECT 284.400 397.000 285.200 399.800 ;
        RECT 286.000 397.000 286.800 399.800 ;
        RECT 287.600 397.000 288.400 399.800 ;
        RECT 286.000 394.400 290.200 395.200 ;
        RECT 290.800 394.400 291.600 399.800 ;
        RECT 294.000 395.200 294.800 399.800 ;
        RECT 294.000 394.600 296.600 395.200 ;
        RECT 290.800 393.600 293.400 394.400 ;
        RECT 284.400 393.000 285.200 393.200 ;
        RECT 276.600 392.400 285.200 393.000 ;
        RECT 287.600 393.000 288.400 393.200 ;
        RECT 296.000 393.000 296.600 394.600 ;
        RECT 287.600 392.400 296.600 393.000 ;
        RECT 296.000 390.600 296.600 392.400 ;
        RECT 297.200 392.000 298.000 399.800 ;
        RECT 306.800 396.400 307.600 399.800 ;
        RECT 306.600 395.800 307.600 396.400 ;
        RECT 306.600 395.200 307.200 395.800 ;
        RECT 310.000 395.200 310.800 399.800 ;
        RECT 313.200 397.000 314.000 399.800 ;
        RECT 314.800 397.000 315.600 399.800 ;
        RECT 305.200 394.600 307.200 395.200 ;
        RECT 297.200 391.200 298.200 392.000 ;
        RECT 266.600 390.000 290.000 390.600 ;
        RECT 296.000 390.000 296.800 390.600 ;
        RECT 266.600 389.800 267.600 390.000 ;
        RECT 266.800 389.600 267.600 389.800 ;
        RECT 271.600 389.600 272.400 390.000 ;
        RECT 289.200 389.400 290.000 390.000 ;
        RECT 265.200 388.200 274.000 389.000 ;
        RECT 274.600 388.600 276.600 389.400 ;
        RECT 280.400 388.600 283.600 389.400 ;
        RECT 262.200 386.800 264.400 387.400 ;
        RECT 263.600 382.200 264.400 386.800 ;
        RECT 265.200 382.200 266.000 388.200 ;
        RECT 267.600 386.800 270.600 387.600 ;
        RECT 269.800 386.200 270.600 386.800 ;
        RECT 275.800 386.200 276.600 388.600 ;
        RECT 278.000 386.800 278.800 388.400 ;
        RECT 283.200 387.800 284.000 388.000 ;
        RECT 279.600 387.200 284.000 387.800 ;
        RECT 279.600 387.000 280.400 387.200 ;
        RECT 286.000 386.400 286.800 389.200 ;
        RECT 291.800 388.600 295.600 389.400 ;
        RECT 291.800 387.400 292.600 388.600 ;
        RECT 296.200 388.000 296.800 390.000 ;
        RECT 279.600 386.200 280.400 386.400 ;
        RECT 269.800 385.400 272.400 386.200 ;
        RECT 275.800 385.600 280.400 386.200 ;
        RECT 281.200 385.600 282.800 386.400 ;
        RECT 285.800 385.600 286.800 386.400 ;
        RECT 290.800 386.800 292.600 387.400 ;
        RECT 295.600 387.400 296.800 388.000 ;
        RECT 290.800 386.200 291.600 386.800 ;
        RECT 271.600 382.200 272.400 385.400 ;
        RECT 289.200 385.400 291.600 386.200 ;
        RECT 273.200 382.200 274.000 385.000 ;
        RECT 274.800 382.200 275.600 385.000 ;
        RECT 276.400 382.200 277.200 385.000 ;
        RECT 279.600 382.200 280.400 385.000 ;
        RECT 282.800 382.200 283.600 385.000 ;
        RECT 284.400 382.200 285.200 385.000 ;
        RECT 286.000 382.200 286.800 385.000 ;
        RECT 287.600 382.200 288.400 385.000 ;
        RECT 289.200 382.200 290.000 385.400 ;
        RECT 295.600 382.200 296.400 387.400 ;
        RECT 297.400 386.800 298.200 391.200 ;
        RECT 297.200 386.000 298.200 386.800 ;
        RECT 305.200 389.000 306.000 394.600 ;
        RECT 307.800 394.400 312.000 395.200 ;
        RECT 316.400 395.000 317.200 399.800 ;
        RECT 319.600 395.000 320.400 399.800 ;
        RECT 307.800 394.000 308.400 394.400 ;
        RECT 306.800 393.200 308.400 394.000 ;
        RECT 311.400 393.800 317.200 394.400 ;
        RECT 309.400 393.200 310.800 393.800 ;
        RECT 309.400 393.000 315.600 393.200 ;
        RECT 310.200 392.600 315.600 393.000 ;
        RECT 314.800 392.400 315.600 392.600 ;
        RECT 316.600 393.000 317.200 393.800 ;
        RECT 317.800 393.600 320.400 394.400 ;
        RECT 322.800 393.600 323.600 399.800 ;
        RECT 324.400 397.000 325.200 399.800 ;
        RECT 326.000 397.000 326.800 399.800 ;
        RECT 327.600 397.000 328.400 399.800 ;
        RECT 326.000 394.400 330.200 395.200 ;
        RECT 330.800 394.400 331.600 399.800 ;
        RECT 334.000 395.200 334.800 399.800 ;
        RECT 334.000 394.600 336.600 395.200 ;
        RECT 330.800 393.600 333.400 394.400 ;
        RECT 324.400 393.000 325.200 393.200 ;
        RECT 316.600 392.400 325.200 393.000 ;
        RECT 327.600 393.000 328.400 393.200 ;
        RECT 336.000 393.000 336.600 394.600 ;
        RECT 327.600 392.400 336.600 393.000 ;
        RECT 336.000 390.600 336.600 392.400 ;
        RECT 337.200 392.000 338.000 399.800 ;
        RECT 342.000 392.000 342.800 399.800 ;
        RECT 345.200 395.200 346.000 399.800 ;
        RECT 337.200 391.200 338.200 392.000 ;
        RECT 306.600 390.000 330.000 390.600 ;
        RECT 336.000 390.000 336.800 390.600 ;
        RECT 306.600 389.800 307.400 390.000 ;
        RECT 311.600 389.600 312.400 390.000 ;
        RECT 329.200 389.400 330.000 390.000 ;
        RECT 305.200 388.200 314.000 389.000 ;
        RECT 314.600 388.600 316.600 389.400 ;
        RECT 320.400 388.600 323.600 389.400 ;
        RECT 297.200 382.200 298.000 386.000 ;
        RECT 305.200 382.200 306.000 388.200 ;
        RECT 307.600 386.800 310.600 387.600 ;
        RECT 309.800 386.200 310.600 386.800 ;
        RECT 315.800 386.200 316.600 388.600 ;
        RECT 318.000 386.800 318.800 388.400 ;
        RECT 323.200 387.800 324.000 388.000 ;
        RECT 319.600 387.200 324.000 387.800 ;
        RECT 319.600 387.000 320.400 387.200 ;
        RECT 326.000 386.400 326.800 389.200 ;
        RECT 331.800 388.600 335.600 389.400 ;
        RECT 331.800 387.400 332.600 388.600 ;
        RECT 336.200 388.000 336.800 390.000 ;
        RECT 319.600 386.200 320.400 386.400 ;
        RECT 309.800 385.400 312.400 386.200 ;
        RECT 315.800 385.600 320.400 386.200 ;
        RECT 321.200 385.600 322.800 386.400 ;
        RECT 325.800 385.600 326.800 386.400 ;
        RECT 330.800 386.800 332.600 387.400 ;
        RECT 335.600 387.400 336.800 388.000 ;
        RECT 330.800 386.200 331.600 386.800 ;
        RECT 311.600 382.200 312.400 385.400 ;
        RECT 329.200 385.400 331.600 386.200 ;
        RECT 313.200 382.200 314.000 385.000 ;
        RECT 314.800 382.200 315.600 385.000 ;
        RECT 316.400 382.200 317.200 385.000 ;
        RECT 319.600 382.200 320.400 385.000 ;
        RECT 322.800 382.200 323.600 385.000 ;
        RECT 324.400 382.200 325.200 385.000 ;
        RECT 326.000 382.200 326.800 385.000 ;
        RECT 327.600 382.200 328.400 385.000 ;
        RECT 329.200 382.200 330.000 385.400 ;
        RECT 335.600 382.200 336.400 387.400 ;
        RECT 337.400 386.800 338.200 391.200 ;
        RECT 337.200 386.000 338.200 386.800 ;
        RECT 341.800 391.200 342.800 392.000 ;
        RECT 343.400 394.600 346.000 395.200 ;
        RECT 343.400 393.000 344.000 394.600 ;
        RECT 348.400 394.400 349.200 399.800 ;
        RECT 351.600 397.000 352.400 399.800 ;
        RECT 353.200 397.000 354.000 399.800 ;
        RECT 354.800 397.000 355.600 399.800 ;
        RECT 349.800 394.400 354.000 395.200 ;
        RECT 346.600 393.600 349.200 394.400 ;
        RECT 356.400 393.600 357.200 399.800 ;
        RECT 359.600 395.000 360.400 399.800 ;
        RECT 362.800 395.000 363.600 399.800 ;
        RECT 364.400 397.000 365.200 399.800 ;
        RECT 366.000 397.000 366.800 399.800 ;
        RECT 369.200 395.200 370.000 399.800 ;
        RECT 372.400 396.400 373.200 399.800 ;
        RECT 372.400 395.800 373.400 396.400 ;
        RECT 372.800 395.200 373.400 395.800 ;
        RECT 368.000 394.400 372.200 395.200 ;
        RECT 372.800 394.600 374.800 395.200 ;
        RECT 359.600 393.600 362.200 394.400 ;
        RECT 362.800 393.800 368.600 394.400 ;
        RECT 371.600 394.000 372.200 394.400 ;
        RECT 351.600 393.000 352.400 393.200 ;
        RECT 343.400 392.400 352.400 393.000 ;
        RECT 354.800 393.000 355.600 393.200 ;
        RECT 362.800 393.000 363.400 393.800 ;
        RECT 369.200 393.200 370.600 393.800 ;
        RECT 371.600 393.200 373.200 394.000 ;
        RECT 354.800 392.400 363.400 393.000 ;
        RECT 364.400 393.000 370.600 393.200 ;
        RECT 364.400 392.600 369.800 393.000 ;
        RECT 364.400 392.400 365.200 392.600 ;
        RECT 341.800 386.800 342.600 391.200 ;
        RECT 343.400 390.600 344.000 392.400 ;
        RECT 343.200 390.000 344.000 390.600 ;
        RECT 350.000 390.000 373.400 390.600 ;
        RECT 343.200 388.000 343.800 390.000 ;
        RECT 350.000 389.400 350.800 390.000 ;
        RECT 367.600 389.600 368.400 390.000 ;
        RECT 372.600 389.800 373.400 390.000 ;
        RECT 344.400 388.600 348.200 389.400 ;
        RECT 343.200 387.400 344.400 388.000 ;
        RECT 341.800 386.000 342.800 386.800 ;
        RECT 337.200 382.200 338.000 386.000 ;
        RECT 342.000 382.200 342.800 386.000 ;
        RECT 343.600 382.200 344.400 387.400 ;
        RECT 347.400 387.400 348.200 388.600 ;
        RECT 347.400 386.800 349.200 387.400 ;
        RECT 348.400 386.200 349.200 386.800 ;
        RECT 353.200 386.400 354.000 389.200 ;
        RECT 356.400 388.600 359.600 389.400 ;
        RECT 363.400 388.600 365.400 389.400 ;
        RECT 374.000 389.000 374.800 394.600 ;
        RECT 375.600 391.400 376.400 399.800 ;
        RECT 380.000 396.400 380.800 399.800 ;
        RECT 378.800 395.800 380.800 396.400 ;
        RECT 384.400 395.800 385.200 399.800 ;
        RECT 388.600 395.800 389.800 399.800 ;
        RECT 378.800 395.000 379.600 395.800 ;
        RECT 384.400 395.200 385.000 395.800 ;
        RECT 382.200 394.600 385.800 395.200 ;
        RECT 388.400 395.000 389.200 395.800 ;
        RECT 382.200 394.400 383.000 394.600 ;
        RECT 385.000 394.400 385.800 394.600 ;
        RECT 378.800 393.000 379.600 393.200 ;
        RECT 383.400 393.000 384.200 393.200 ;
        RECT 378.800 392.400 384.200 393.000 ;
        RECT 384.800 393.000 387.000 393.600 ;
        RECT 384.800 391.800 385.400 393.000 ;
        RECT 386.200 392.800 387.000 393.000 ;
        RECT 388.600 393.200 390.000 394.000 ;
        RECT 388.600 392.200 389.200 393.200 ;
        RECT 380.600 391.400 385.400 391.800 ;
        RECT 375.600 391.200 385.400 391.400 ;
        RECT 386.800 391.600 389.200 392.200 ;
        RECT 375.600 391.000 381.400 391.200 ;
        RECT 375.600 390.800 381.200 391.000 ;
        RECT 386.800 390.400 387.400 391.600 ;
        RECT 393.200 391.200 394.000 399.800 ;
        RECT 389.800 390.600 394.000 391.200 ;
        RECT 389.800 390.400 390.600 390.600 ;
        RECT 382.000 390.200 382.800 390.400 ;
        RECT 377.800 389.600 382.800 390.200 ;
        RECT 386.800 389.600 387.600 390.400 ;
        RECT 391.400 389.800 392.200 390.000 ;
        RECT 377.800 389.400 378.600 389.600 ;
        RECT 380.400 389.400 381.200 389.600 ;
        RECT 356.000 387.800 356.800 388.000 ;
        RECT 356.000 387.200 360.400 387.800 ;
        RECT 359.600 387.000 360.400 387.200 ;
        RECT 361.200 386.800 362.000 388.400 ;
        RECT 348.400 385.400 350.800 386.200 ;
        RECT 353.200 385.600 354.200 386.400 ;
        RECT 357.200 385.600 358.800 386.400 ;
        RECT 359.600 386.200 360.400 386.400 ;
        RECT 363.400 386.200 364.200 388.600 ;
        RECT 366.000 388.200 374.800 389.000 ;
        RECT 379.400 388.400 380.200 388.600 ;
        RECT 386.800 388.400 387.400 389.600 ;
        RECT 388.400 389.200 392.200 389.800 ;
        RECT 388.400 389.000 389.200 389.200 ;
        RECT 369.400 386.800 372.400 387.600 ;
        RECT 369.400 386.200 370.200 386.800 ;
        RECT 359.600 385.600 364.200 386.200 ;
        RECT 350.000 382.200 350.800 385.400 ;
        RECT 367.600 385.400 370.200 386.200 ;
        RECT 351.600 382.200 352.400 385.000 ;
        RECT 353.200 382.200 354.000 385.000 ;
        RECT 354.800 382.200 355.600 385.000 ;
        RECT 356.400 382.200 357.200 385.000 ;
        RECT 359.600 382.200 360.400 385.000 ;
        RECT 362.800 382.200 363.600 385.000 ;
        RECT 364.400 382.200 365.200 385.000 ;
        RECT 366.000 382.200 366.800 385.000 ;
        RECT 367.600 382.200 368.400 385.400 ;
        RECT 374.000 382.200 374.800 388.200 ;
        RECT 376.400 387.800 387.400 388.400 ;
        RECT 376.400 387.600 378.000 387.800 ;
        RECT 375.600 382.200 376.400 387.000 ;
        RECT 380.600 385.600 381.200 387.800 ;
        RECT 386.200 387.600 387.000 387.800 ;
        RECT 393.200 387.200 394.000 390.600 ;
        RECT 390.200 386.600 394.000 387.200 ;
        RECT 390.200 386.400 391.000 386.600 ;
        RECT 378.800 384.200 379.600 385.000 ;
        RECT 380.400 384.800 381.200 385.600 ;
        RECT 382.200 385.400 383.000 385.600 ;
        RECT 382.200 384.800 385.000 385.400 ;
        RECT 384.400 384.200 385.000 384.800 ;
        RECT 388.400 384.200 389.200 385.000 ;
        RECT 378.800 383.600 380.800 384.200 ;
        RECT 380.000 382.200 380.800 383.600 ;
        RECT 384.400 382.200 385.200 384.200 ;
        RECT 388.400 383.600 389.800 384.200 ;
        RECT 388.600 382.200 389.800 383.600 ;
        RECT 393.200 382.200 394.000 386.600 ;
        RECT 394.800 384.800 395.600 386.400 ;
        RECT 396.400 382.200 397.200 399.800 ;
        RECT 398.000 384.800 398.800 386.400 ;
        RECT 399.600 382.200 400.400 399.800 ;
        RECT 401.200 392.400 402.000 399.800 ;
        RECT 404.400 392.800 405.200 399.800 ;
        RECT 401.200 391.800 403.800 392.400 ;
        RECT 404.400 391.800 405.400 392.800 ;
        RECT 409.200 392.000 410.000 399.800 ;
        RECT 412.400 395.200 413.200 399.800 ;
        RECT 401.200 389.600 402.200 390.400 ;
        RECT 401.400 388.800 402.200 389.600 ;
        RECT 403.200 389.800 403.800 391.800 ;
        RECT 403.200 389.000 404.200 389.800 ;
        RECT 403.200 387.400 403.800 389.000 ;
        RECT 404.800 388.400 405.400 391.800 ;
        RECT 404.400 387.600 405.400 388.400 ;
        RECT 401.200 386.800 403.800 387.400 ;
        RECT 401.200 382.200 402.000 386.800 ;
        RECT 404.800 386.200 405.400 387.600 ;
        RECT 404.400 385.600 405.400 386.200 ;
        RECT 409.000 391.200 410.000 392.000 ;
        RECT 410.600 394.600 413.200 395.200 ;
        RECT 410.600 393.000 411.200 394.600 ;
        RECT 415.600 394.400 416.400 399.800 ;
        RECT 418.800 397.000 419.600 399.800 ;
        RECT 420.400 397.000 421.200 399.800 ;
        RECT 422.000 397.000 422.800 399.800 ;
        RECT 417.000 394.400 421.200 395.200 ;
        RECT 413.800 393.600 416.400 394.400 ;
        RECT 423.600 393.600 424.400 399.800 ;
        RECT 426.800 395.000 427.600 399.800 ;
        RECT 430.000 395.000 430.800 399.800 ;
        RECT 431.600 397.000 432.400 399.800 ;
        RECT 433.200 397.000 434.000 399.800 ;
        RECT 436.400 395.200 437.200 399.800 ;
        RECT 439.600 396.400 440.400 399.800 ;
        RECT 439.600 395.800 440.600 396.400 ;
        RECT 440.000 395.200 440.600 395.800 ;
        RECT 435.200 394.400 439.400 395.200 ;
        RECT 440.000 394.600 442.000 395.200 ;
        RECT 426.800 393.600 429.400 394.400 ;
        RECT 430.000 393.800 435.800 394.400 ;
        RECT 438.800 394.000 439.400 394.400 ;
        RECT 418.800 393.000 419.600 393.200 ;
        RECT 410.600 392.400 419.600 393.000 ;
        RECT 422.000 393.000 422.800 393.200 ;
        RECT 430.000 393.000 430.600 393.800 ;
        RECT 436.400 393.200 437.800 393.800 ;
        RECT 438.800 393.200 440.400 394.000 ;
        RECT 422.000 392.400 430.600 393.000 ;
        RECT 431.600 393.000 437.800 393.200 ;
        RECT 431.600 392.600 437.000 393.000 ;
        RECT 431.600 392.400 432.400 392.600 ;
        RECT 409.000 386.800 409.800 391.200 ;
        RECT 410.600 390.600 411.200 392.400 ;
        RECT 410.400 390.000 411.200 390.600 ;
        RECT 417.200 390.000 440.600 390.600 ;
        RECT 410.400 388.000 411.000 390.000 ;
        RECT 417.200 389.400 418.000 390.000 ;
        RECT 434.800 389.600 435.600 390.000 ;
        RECT 438.000 389.600 438.800 390.000 ;
        RECT 439.800 389.800 440.600 390.000 ;
        RECT 411.600 388.600 415.400 389.400 ;
        RECT 410.400 387.400 411.600 388.000 ;
        RECT 409.000 386.000 410.000 386.800 ;
        RECT 404.400 382.200 405.200 385.600 ;
        RECT 409.200 382.200 410.000 386.000 ;
        RECT 410.800 382.200 411.600 387.400 ;
        RECT 414.600 387.400 415.400 388.600 ;
        RECT 414.600 386.800 416.400 387.400 ;
        RECT 415.600 386.200 416.400 386.800 ;
        RECT 420.400 386.400 421.200 389.200 ;
        RECT 423.600 388.600 426.800 389.400 ;
        RECT 430.600 388.600 432.600 389.400 ;
        RECT 441.200 389.000 442.000 394.600 ;
        RECT 442.800 391.600 443.600 393.200 ;
        RECT 423.200 387.800 424.000 388.000 ;
        RECT 423.200 387.200 427.600 387.800 ;
        RECT 426.800 387.000 427.600 387.200 ;
        RECT 428.400 386.800 429.200 388.400 ;
        RECT 415.600 385.400 418.000 386.200 ;
        RECT 420.400 385.600 421.400 386.400 ;
        RECT 424.400 385.600 426.000 386.400 ;
        RECT 426.800 386.200 427.600 386.400 ;
        RECT 430.600 386.200 431.400 388.600 ;
        RECT 433.200 388.200 442.000 389.000 ;
        RECT 436.600 386.800 439.600 387.600 ;
        RECT 436.600 386.200 437.400 386.800 ;
        RECT 426.800 385.600 431.400 386.200 ;
        RECT 417.200 382.200 418.000 385.400 ;
        RECT 434.800 385.400 437.400 386.200 ;
        RECT 418.800 382.200 419.600 385.000 ;
        RECT 420.400 382.200 421.200 385.000 ;
        RECT 422.000 382.200 422.800 385.000 ;
        RECT 423.600 382.200 424.400 385.000 ;
        RECT 426.800 382.200 427.600 385.000 ;
        RECT 430.000 382.200 430.800 385.000 ;
        RECT 431.600 382.200 432.400 385.000 ;
        RECT 433.200 382.200 434.000 385.000 ;
        RECT 434.800 382.200 435.600 385.400 ;
        RECT 441.200 382.200 442.000 388.200 ;
        RECT 442.800 388.300 443.600 388.400 ;
        RECT 444.400 388.300 445.200 399.800 ;
        RECT 446.000 394.300 446.800 394.400 ;
        RECT 448.400 394.300 449.200 394.400 ;
        RECT 446.000 393.700 449.200 394.300 ;
        RECT 446.000 393.600 446.800 393.700 ;
        RECT 448.400 393.600 449.200 393.700 ;
        RECT 448.400 392.400 449.000 393.600 ;
        RECT 449.800 392.400 450.600 399.800 ;
        RECT 460.400 396.400 461.200 399.800 ;
        RECT 460.200 395.800 461.200 396.400 ;
        RECT 460.200 395.200 460.800 395.800 ;
        RECT 463.600 395.200 464.400 399.800 ;
        RECT 466.800 397.000 467.600 399.800 ;
        RECT 468.400 397.000 469.200 399.800 ;
        RECT 447.600 391.800 449.000 392.400 ;
        RECT 449.600 391.800 450.600 392.400 ;
        RECT 458.800 394.600 460.800 395.200 ;
        RECT 447.600 391.600 448.400 391.800 ;
        RECT 449.600 388.400 450.200 391.800 ;
        RECT 450.800 388.800 451.600 390.400 ;
        RECT 458.800 389.000 459.600 394.600 ;
        RECT 461.400 394.400 465.600 395.200 ;
        RECT 470.000 395.000 470.800 399.800 ;
        RECT 473.200 395.000 474.000 399.800 ;
        RECT 461.400 394.000 462.000 394.400 ;
        RECT 460.400 393.200 462.000 394.000 ;
        RECT 465.000 393.800 470.800 394.400 ;
        RECT 463.000 393.200 464.400 393.800 ;
        RECT 463.000 393.000 469.200 393.200 ;
        RECT 463.800 392.600 469.200 393.000 ;
        RECT 468.400 392.400 469.200 392.600 ;
        RECT 470.200 393.000 470.800 393.800 ;
        RECT 471.400 393.600 474.000 394.400 ;
        RECT 476.400 393.600 477.200 399.800 ;
        RECT 478.000 397.000 478.800 399.800 ;
        RECT 479.600 397.000 480.400 399.800 ;
        RECT 481.200 397.000 482.000 399.800 ;
        RECT 479.600 394.400 483.800 395.200 ;
        RECT 484.400 394.400 485.200 399.800 ;
        RECT 487.600 395.200 488.400 399.800 ;
        RECT 487.600 394.600 490.200 395.200 ;
        RECT 484.400 393.600 487.000 394.400 ;
        RECT 478.000 393.000 478.800 393.200 ;
        RECT 470.200 392.400 478.800 393.000 ;
        RECT 481.200 393.000 482.000 393.200 ;
        RECT 489.600 393.000 490.200 394.600 ;
        RECT 481.200 392.400 490.200 393.000 ;
        RECT 489.600 390.600 490.200 392.400 ;
        RECT 490.800 392.000 491.600 399.800 ;
        RECT 490.800 391.200 491.800 392.000 ;
        RECT 495.600 391.200 496.400 399.800 ;
        RECT 498.800 391.200 499.600 399.800 ;
        RECT 502.000 391.200 502.800 399.800 ;
        RECT 505.200 391.200 506.000 399.800 ;
        RECT 509.000 398.400 509.800 399.800 ;
        RECT 509.000 397.600 510.800 398.400 ;
        RECT 509.000 392.600 509.800 397.600 ;
        RECT 509.000 391.800 510.800 392.600 ;
        RECT 460.200 390.000 483.600 390.600 ;
        RECT 489.600 390.000 490.400 390.600 ;
        RECT 460.200 389.800 461.000 390.000 ;
        RECT 465.200 389.600 466.000 390.000 ;
        RECT 482.800 389.400 483.600 390.000 ;
        RECT 442.800 387.700 445.200 388.300 ;
        RECT 442.800 387.600 443.600 387.700 ;
        RECT 444.400 386.200 445.200 387.700 ;
        RECT 446.000 388.300 446.800 388.400 ;
        RECT 447.600 388.300 450.200 388.400 ;
        RECT 446.000 387.700 450.200 388.300 ;
        RECT 452.400 388.200 453.200 388.400 ;
        RECT 446.000 386.800 446.800 387.700 ;
        RECT 447.600 387.600 450.200 387.700 ;
        RECT 451.600 387.600 453.200 388.200 ;
        RECT 458.800 388.200 467.600 389.000 ;
        RECT 468.200 388.600 470.200 389.400 ;
        RECT 474.000 388.600 477.200 389.400 ;
        RECT 447.800 386.200 448.400 387.600 ;
        RECT 451.600 387.200 452.400 387.600 ;
        RECT 449.400 386.200 453.000 386.600 ;
        RECT 443.400 385.600 445.200 386.200 ;
        RECT 443.400 382.200 444.200 385.600 ;
        RECT 447.600 382.200 448.400 386.200 ;
        RECT 449.200 386.000 453.200 386.200 ;
        RECT 449.200 382.200 450.000 386.000 ;
        RECT 452.400 382.200 453.200 386.000 ;
        RECT 458.800 382.200 459.600 388.200 ;
        RECT 461.200 386.800 464.200 387.600 ;
        RECT 463.400 386.200 464.200 386.800 ;
        RECT 469.400 386.200 470.200 388.600 ;
        RECT 471.600 386.800 472.400 388.400 ;
        RECT 476.800 387.800 477.600 388.000 ;
        RECT 473.200 387.200 477.600 387.800 ;
        RECT 473.200 387.000 474.000 387.200 ;
        RECT 479.600 386.400 480.400 389.200 ;
        RECT 485.400 388.600 489.200 389.400 ;
        RECT 485.400 387.400 486.200 388.600 ;
        RECT 489.800 388.000 490.400 390.000 ;
        RECT 473.200 386.200 474.000 386.400 ;
        RECT 463.400 385.400 466.000 386.200 ;
        RECT 469.400 385.600 474.000 386.200 ;
        RECT 474.800 385.600 476.400 386.400 ;
        RECT 479.400 385.600 480.400 386.400 ;
        RECT 484.400 386.800 486.200 387.400 ;
        RECT 489.200 387.400 490.400 388.000 ;
        RECT 484.400 386.200 485.200 386.800 ;
        RECT 465.200 382.200 466.000 385.400 ;
        RECT 482.800 385.400 485.200 386.200 ;
        RECT 466.800 382.200 467.600 385.000 ;
        RECT 468.400 382.200 469.200 385.000 ;
        RECT 470.000 382.200 470.800 385.000 ;
        RECT 473.200 382.200 474.000 385.000 ;
        RECT 476.400 382.200 477.200 385.000 ;
        RECT 478.000 382.200 478.800 385.000 ;
        RECT 479.600 382.200 480.400 385.000 ;
        RECT 481.200 382.200 482.000 385.000 ;
        RECT 482.800 382.200 483.600 385.400 ;
        RECT 489.200 382.200 490.000 387.400 ;
        RECT 491.000 386.800 491.800 391.200 ;
        RECT 494.000 390.400 496.400 391.200 ;
        RECT 497.400 390.400 499.600 391.200 ;
        RECT 500.600 390.400 502.800 391.200 ;
        RECT 504.200 390.400 506.000 391.200 ;
        RECT 494.000 387.600 494.800 390.400 ;
        RECT 497.400 389.000 498.200 390.400 ;
        RECT 500.600 389.000 501.400 390.400 ;
        RECT 504.200 389.000 505.000 390.400 ;
        RECT 508.400 389.600 509.200 391.200 ;
        RECT 495.600 388.200 498.200 389.000 ;
        RECT 499.000 388.200 501.400 389.000 ;
        RECT 502.400 388.200 505.000 389.000 ;
        RECT 505.800 388.200 507.600 389.000 ;
        RECT 497.400 387.600 498.200 388.200 ;
        RECT 500.600 387.600 501.400 388.200 ;
        RECT 504.200 387.600 505.000 388.200 ;
        RECT 506.800 387.600 507.600 388.200 ;
        RECT 510.000 388.400 510.600 391.800 ;
        RECT 513.200 391.600 514.000 393.200 ;
        RECT 510.000 387.600 510.800 388.400 ;
        RECT 494.000 386.800 496.400 387.600 ;
        RECT 497.400 386.800 499.600 387.600 ;
        RECT 500.600 386.800 502.800 387.600 ;
        RECT 504.200 386.800 506.000 387.600 ;
        RECT 490.800 386.000 491.800 386.800 ;
        RECT 490.800 382.200 491.600 386.000 ;
        RECT 495.600 382.200 496.400 386.800 ;
        RECT 498.800 382.200 499.600 386.800 ;
        RECT 502.000 382.200 502.800 386.800 ;
        RECT 505.200 382.200 506.000 386.800 ;
        RECT 510.000 384.200 510.600 387.600 ;
        RECT 511.600 384.800 512.400 386.400 ;
        RECT 514.800 386.200 515.600 399.800 ;
        RECT 519.600 396.400 520.400 399.800 ;
        RECT 519.400 395.800 520.400 396.400 ;
        RECT 519.400 395.200 520.000 395.800 ;
        RECT 522.800 395.200 523.600 399.800 ;
        RECT 526.000 397.000 526.800 399.800 ;
        RECT 527.600 397.000 528.400 399.800 ;
        RECT 518.000 394.600 520.000 395.200 ;
        RECT 518.000 389.000 518.800 394.600 ;
        RECT 520.600 394.400 524.800 395.200 ;
        RECT 529.200 395.000 530.000 399.800 ;
        RECT 532.400 395.000 533.200 399.800 ;
        RECT 520.600 394.000 521.200 394.400 ;
        RECT 519.600 393.200 521.200 394.000 ;
        RECT 524.200 393.800 530.000 394.400 ;
        RECT 522.200 393.200 523.600 393.800 ;
        RECT 522.200 393.000 528.400 393.200 ;
        RECT 523.000 392.600 528.400 393.000 ;
        RECT 527.600 392.400 528.400 392.600 ;
        RECT 529.400 393.000 530.000 393.800 ;
        RECT 530.600 393.600 533.200 394.400 ;
        RECT 535.600 393.600 536.400 399.800 ;
        RECT 537.200 397.000 538.000 399.800 ;
        RECT 538.800 397.000 539.600 399.800 ;
        RECT 540.400 397.000 541.200 399.800 ;
        RECT 538.800 394.400 543.000 395.200 ;
        RECT 543.600 394.400 544.400 399.800 ;
        RECT 546.800 395.200 547.600 399.800 ;
        RECT 546.800 394.600 549.400 395.200 ;
        RECT 543.600 393.600 546.200 394.400 ;
        RECT 537.200 393.000 538.000 393.200 ;
        RECT 529.400 392.400 538.000 393.000 ;
        RECT 540.400 393.000 541.200 393.200 ;
        RECT 548.800 393.000 549.400 394.600 ;
        RECT 540.400 392.400 549.400 393.000 ;
        RECT 548.800 390.600 549.400 392.400 ;
        RECT 550.000 392.000 550.800 399.800 ;
        RECT 553.800 392.600 554.600 399.800 ;
        RECT 560.200 394.400 561.000 399.800 ;
        RECT 558.800 393.600 559.600 394.400 ;
        RECT 560.200 393.600 562.000 394.400 ;
        RECT 550.000 391.200 551.000 392.000 ;
        RECT 553.800 391.800 555.600 392.600 ;
        RECT 558.800 392.400 559.400 393.600 ;
        RECT 560.200 392.400 561.000 393.600 ;
        RECT 558.000 391.800 559.400 392.400 ;
        RECT 560.000 391.800 561.000 392.400 ;
        RECT 519.400 390.000 542.800 390.600 ;
        RECT 548.800 390.000 549.600 390.600 ;
        RECT 519.400 389.800 520.400 390.000 ;
        RECT 519.600 389.600 520.400 389.800 ;
        RECT 521.200 389.600 522.000 390.000 ;
        RECT 524.400 389.600 525.200 390.000 ;
        RECT 542.000 389.400 542.800 390.000 ;
        RECT 516.400 386.800 517.200 388.400 ;
        RECT 518.000 388.200 526.800 389.000 ;
        RECT 527.400 388.600 529.400 389.400 ;
        RECT 533.200 388.600 536.400 389.400 ;
        RECT 513.800 385.600 515.600 386.200 ;
        RECT 510.000 382.200 510.800 384.200 ;
        RECT 513.800 382.200 514.600 385.600 ;
        RECT 518.000 382.200 518.800 388.200 ;
        RECT 520.400 386.800 523.400 387.600 ;
        RECT 522.600 386.200 523.400 386.800 ;
        RECT 528.600 386.200 529.400 388.600 ;
        RECT 530.800 386.800 531.600 388.400 ;
        RECT 536.000 387.800 536.800 388.000 ;
        RECT 532.400 387.200 536.800 387.800 ;
        RECT 532.400 387.000 533.200 387.200 ;
        RECT 538.800 386.400 539.600 389.200 ;
        RECT 544.600 388.600 548.400 389.400 ;
        RECT 544.600 387.400 545.400 388.600 ;
        RECT 549.000 388.000 549.600 390.000 ;
        RECT 532.400 386.200 533.200 386.400 ;
        RECT 522.600 385.400 525.200 386.200 ;
        RECT 528.600 385.600 533.200 386.200 ;
        RECT 534.000 385.600 535.600 386.400 ;
        RECT 538.600 385.600 539.600 386.400 ;
        RECT 543.600 386.800 545.400 387.400 ;
        RECT 548.400 387.400 549.600 388.000 ;
        RECT 543.600 386.200 544.400 386.800 ;
        RECT 524.400 382.200 525.200 385.400 ;
        RECT 542.000 385.400 544.400 386.200 ;
        RECT 526.000 382.200 526.800 385.000 ;
        RECT 527.600 382.200 528.400 385.000 ;
        RECT 529.200 382.200 530.000 385.000 ;
        RECT 532.400 382.200 533.200 385.000 ;
        RECT 535.600 382.200 536.400 385.000 ;
        RECT 537.200 382.200 538.000 385.000 ;
        RECT 538.800 382.200 539.600 385.000 ;
        RECT 540.400 382.200 541.200 385.000 ;
        RECT 542.000 382.200 542.800 385.400 ;
        RECT 548.400 382.200 549.200 387.400 ;
        RECT 550.200 386.800 551.000 391.200 ;
        RECT 551.600 390.300 552.400 390.400 ;
        RECT 553.200 390.300 554.000 391.200 ;
        RECT 551.600 389.700 554.000 390.300 ;
        RECT 551.600 389.600 552.400 389.700 ;
        RECT 553.200 389.600 554.000 389.700 ;
        RECT 554.800 390.300 555.400 391.800 ;
        RECT 558.000 391.600 558.800 391.800 ;
        RECT 558.000 390.300 558.800 390.400 ;
        RECT 554.800 389.700 558.800 390.300 ;
        RECT 550.000 386.000 551.000 386.800 ;
        RECT 554.800 388.400 555.400 389.700 ;
        RECT 558.000 389.600 558.800 389.700 ;
        RECT 560.000 388.400 560.600 391.800 ;
        RECT 561.200 388.800 562.000 390.400 ;
        RECT 554.800 387.600 555.600 388.400 ;
        RECT 558.000 387.600 560.600 388.400 ;
        RECT 562.800 388.300 563.600 388.400 ;
        RECT 564.400 388.300 565.200 399.800 ;
        RECT 568.200 398.400 569.000 399.800 ;
        RECT 567.600 397.600 569.000 398.400 ;
        RECT 568.200 392.400 569.000 397.600 ;
        RECT 562.800 388.200 565.200 388.300 ;
        RECT 562.000 387.700 565.200 388.200 ;
        RECT 562.000 387.600 563.600 387.700 ;
        RECT 550.000 382.200 550.800 386.000 ;
        RECT 554.800 384.400 555.400 387.600 ;
        RECT 556.400 384.800 557.200 386.400 ;
        RECT 558.200 386.200 558.800 387.600 ;
        RECT 562.000 387.200 562.800 387.600 ;
        RECT 559.800 386.200 563.400 386.600 ;
        RECT 554.800 382.200 555.600 384.400 ;
        RECT 558.000 382.200 558.800 386.200 ;
        RECT 559.600 386.000 563.600 386.200 ;
        RECT 559.600 382.200 560.400 386.000 ;
        RECT 562.800 382.200 563.600 386.000 ;
        RECT 564.400 382.200 565.200 387.700 ;
        RECT 567.600 391.800 569.000 392.400 ;
        RECT 567.600 390.400 568.200 391.800 ;
        RECT 572.400 391.200 573.200 399.800 ;
        RECT 575.600 396.400 576.400 399.800 ;
        RECT 575.400 395.800 576.400 396.400 ;
        RECT 575.400 395.200 576.000 395.800 ;
        RECT 578.800 395.200 579.600 399.800 ;
        RECT 582.000 397.000 582.800 399.800 ;
        RECT 583.600 397.000 584.400 399.800 ;
        RECT 569.200 390.800 573.200 391.200 ;
        RECT 569.000 390.600 573.200 390.800 ;
        RECT 574.000 394.600 576.000 395.200 ;
        RECT 567.600 389.600 568.400 390.400 ;
        RECT 569.000 390.000 569.800 390.600 ;
        RECT 566.000 384.800 566.800 386.400 ;
        RECT 567.600 386.200 568.200 389.600 ;
        RECT 569.000 387.000 569.600 390.000 ;
        RECT 570.400 388.400 571.200 389.200 ;
        RECT 574.000 389.000 574.800 394.600 ;
        RECT 576.600 394.400 580.800 395.200 ;
        RECT 585.200 395.000 586.000 399.800 ;
        RECT 588.400 395.000 589.200 399.800 ;
        RECT 576.600 394.000 577.200 394.400 ;
        RECT 575.600 393.200 577.200 394.000 ;
        RECT 580.200 393.800 586.000 394.400 ;
        RECT 578.200 393.200 579.600 393.800 ;
        RECT 578.200 393.000 584.400 393.200 ;
        RECT 579.000 392.600 584.400 393.000 ;
        RECT 583.600 392.400 584.400 392.600 ;
        RECT 585.400 393.000 586.000 393.800 ;
        RECT 586.600 393.600 589.200 394.400 ;
        RECT 591.600 393.600 592.400 399.800 ;
        RECT 593.200 397.000 594.000 399.800 ;
        RECT 594.800 397.000 595.600 399.800 ;
        RECT 596.400 397.000 597.200 399.800 ;
        RECT 594.800 394.400 599.000 395.200 ;
        RECT 599.600 394.400 600.400 399.800 ;
        RECT 602.800 395.200 603.600 399.800 ;
        RECT 602.800 394.600 605.400 395.200 ;
        RECT 599.600 393.600 602.200 394.400 ;
        RECT 593.200 393.000 594.000 393.200 ;
        RECT 585.400 392.400 594.000 393.000 ;
        RECT 596.400 393.000 597.200 393.200 ;
        RECT 604.800 393.000 605.400 394.600 ;
        RECT 596.400 392.400 605.400 393.000 ;
        RECT 604.800 390.600 605.400 392.400 ;
        RECT 606.000 392.000 606.800 399.800 ;
        RECT 606.000 391.200 607.000 392.000 ;
        RECT 575.400 390.000 598.800 390.600 ;
        RECT 604.800 390.000 605.600 390.600 ;
        RECT 575.400 389.800 576.400 390.000 ;
        RECT 575.600 389.600 576.400 389.800 ;
        RECT 577.200 389.600 578.000 390.000 ;
        RECT 580.400 389.600 581.200 390.000 ;
        RECT 598.000 389.400 598.800 390.000 ;
        RECT 570.600 387.600 571.600 388.400 ;
        RECT 574.000 388.200 582.800 389.000 ;
        RECT 583.400 388.600 585.400 389.400 ;
        RECT 589.200 388.600 592.400 389.400 ;
        RECT 569.000 386.400 571.400 387.000 ;
        RECT 567.600 382.200 568.400 386.200 ;
        RECT 570.800 384.200 571.400 386.400 ;
        RECT 572.400 384.800 573.200 386.400 ;
        RECT 570.800 382.200 571.600 384.200 ;
        RECT 574.000 382.200 574.800 388.200 ;
        RECT 576.400 386.800 579.400 387.600 ;
        RECT 578.600 386.200 579.400 386.800 ;
        RECT 584.600 386.200 585.400 388.600 ;
        RECT 586.800 386.800 587.600 388.400 ;
        RECT 592.000 387.800 592.800 388.000 ;
        RECT 588.400 387.200 592.800 387.800 ;
        RECT 588.400 387.000 589.200 387.200 ;
        RECT 594.800 386.400 595.600 389.200 ;
        RECT 600.600 388.600 604.400 389.400 ;
        RECT 600.600 387.400 601.400 388.600 ;
        RECT 605.000 388.000 605.600 390.000 ;
        RECT 588.400 386.200 589.200 386.400 ;
        RECT 578.600 385.400 581.200 386.200 ;
        RECT 584.600 385.600 589.200 386.200 ;
        RECT 590.000 385.600 591.600 386.400 ;
        RECT 594.600 385.600 595.600 386.400 ;
        RECT 599.600 386.800 601.400 387.400 ;
        RECT 604.400 387.400 605.600 388.000 ;
        RECT 599.600 386.200 600.400 386.800 ;
        RECT 580.400 382.200 581.200 385.400 ;
        RECT 598.000 385.400 600.400 386.200 ;
        RECT 582.000 382.200 582.800 385.000 ;
        RECT 583.600 382.200 584.400 385.000 ;
        RECT 585.200 382.200 586.000 385.000 ;
        RECT 588.400 382.200 589.200 385.000 ;
        RECT 591.600 382.200 592.400 385.000 ;
        RECT 593.200 382.200 594.000 385.000 ;
        RECT 594.800 382.200 595.600 385.000 ;
        RECT 596.400 382.200 597.200 385.000 ;
        RECT 598.000 382.200 598.800 385.400 ;
        RECT 604.400 382.200 605.200 387.400 ;
        RECT 606.200 386.800 607.000 391.200 ;
        RECT 606.000 386.000 607.000 386.800 ;
        RECT 606.000 382.200 606.800 386.000 ;
        RECT 2.800 372.300 3.600 379.800 ;
        RECT 4.400 372.300 5.200 372.400 ;
        RECT 2.800 371.700 5.200 372.300 ;
        RECT 2.800 362.200 3.600 371.700 ;
        RECT 4.400 371.600 5.200 371.700 ;
        RECT 6.000 362.200 6.800 379.800 ;
        RECT 7.600 376.000 8.400 379.800 ;
        RECT 10.800 376.000 11.600 379.800 ;
        RECT 7.600 375.800 11.600 376.000 ;
        RECT 12.400 375.800 13.200 379.800 ;
        RECT 14.000 376.000 14.800 379.800 ;
        RECT 17.200 376.000 18.000 379.800 ;
        RECT 14.000 375.800 18.000 376.000 ;
        RECT 18.800 375.800 19.600 379.800 ;
        RECT 20.400 375.800 21.200 379.800 ;
        RECT 22.000 376.000 22.800 379.800 ;
        RECT 25.200 376.000 26.000 379.800 ;
        RECT 22.000 375.800 26.000 376.000 ;
        RECT 26.800 376.000 27.600 379.800 ;
        RECT 30.000 376.000 30.800 379.800 ;
        RECT 26.800 375.800 30.800 376.000 ;
        RECT 31.600 375.800 32.400 379.800 ;
        RECT 7.800 375.400 11.400 375.800 ;
        RECT 8.400 374.400 9.200 374.800 ;
        RECT 12.400 374.400 13.000 375.800 ;
        RECT 14.200 375.400 17.800 375.800 ;
        RECT 14.800 374.400 15.600 374.800 ;
        RECT 18.800 374.400 19.400 375.800 ;
        RECT 20.600 374.400 21.200 375.800 ;
        RECT 22.200 375.400 25.800 375.800 ;
        RECT 27.000 375.400 30.600 375.800 ;
        RECT 24.400 374.400 25.200 374.800 ;
        RECT 27.600 374.400 28.400 374.800 ;
        RECT 31.600 374.400 32.200 375.800 ;
        RECT 33.200 375.600 34.000 379.800 ;
        RECT 34.800 376.000 35.600 379.800 ;
        RECT 38.000 376.000 38.800 379.800 ;
        RECT 34.800 375.800 38.800 376.000 ;
        RECT 39.600 375.800 40.400 379.800 ;
        RECT 41.200 376.000 42.000 379.800 ;
        RECT 44.400 376.000 45.200 379.800 ;
        RECT 41.200 375.800 45.200 376.000 ;
        RECT 46.600 376.400 47.400 379.800 ;
        RECT 46.600 375.800 48.400 376.400 ;
        RECT 50.800 375.800 51.600 379.800 ;
        RECT 52.400 376.000 53.200 379.800 ;
        RECT 55.600 376.000 56.400 379.800 ;
        RECT 52.400 375.800 56.400 376.000 ;
        RECT 57.200 377.000 58.000 379.000 ;
        RECT 33.400 374.400 34.000 375.600 ;
        RECT 35.000 375.400 38.600 375.800 ;
        RECT 37.200 374.400 38.000 374.800 ;
        RECT 39.800 374.400 40.400 375.800 ;
        RECT 41.400 375.400 45.000 375.800 ;
        RECT 43.600 374.400 44.400 374.800 ;
        RECT 7.600 373.800 9.200 374.400 ;
        RECT 7.600 373.600 8.400 373.800 ;
        RECT 10.600 373.600 13.200 374.400 ;
        RECT 14.000 373.800 15.600 374.400 ;
        RECT 14.000 373.600 14.800 373.800 ;
        RECT 17.000 373.600 19.600 374.400 ;
        RECT 20.400 373.600 23.000 374.400 ;
        RECT 24.400 374.300 26.000 374.400 ;
        RECT 26.800 374.300 28.400 374.400 ;
        RECT 24.400 373.800 28.400 374.300 ;
        RECT 25.200 373.700 27.600 373.800 ;
        RECT 25.200 373.600 26.000 373.700 ;
        RECT 26.800 373.600 27.600 373.700 ;
        RECT 29.800 373.600 32.400 374.400 ;
        RECT 33.200 373.600 35.800 374.400 ;
        RECT 37.200 373.800 38.800 374.400 ;
        RECT 38.000 373.600 38.800 373.800 ;
        RECT 39.600 373.600 42.200 374.400 ;
        RECT 43.600 373.800 45.200 374.400 ;
        RECT 44.400 373.600 45.200 373.800 ;
        RECT 9.200 371.600 10.000 373.200 ;
        RECT 10.600 370.200 11.200 373.600 ;
        RECT 15.600 371.600 16.400 373.200 ;
        RECT 12.400 370.200 13.200 370.400 ;
        RECT 17.000 370.200 17.600 373.600 ;
        RECT 22.400 372.300 23.000 373.600 ;
        RECT 18.900 371.700 23.000 372.300 ;
        RECT 18.900 370.400 19.500 371.700 ;
        RECT 18.800 370.200 19.600 370.400 ;
        RECT 10.200 369.600 11.200 370.200 ;
        RECT 11.800 369.600 13.200 370.200 ;
        RECT 16.600 369.600 17.600 370.200 ;
        RECT 18.200 369.600 19.600 370.200 ;
        RECT 20.400 370.200 21.200 370.400 ;
        RECT 22.400 370.200 23.000 371.700 ;
        RECT 23.600 372.300 24.400 373.200 ;
        RECT 28.400 372.300 29.200 373.200 ;
        RECT 23.600 371.700 29.200 372.300 ;
        RECT 23.600 371.600 24.400 371.700 ;
        RECT 28.400 371.600 29.200 371.700 ;
        RECT 29.800 370.200 30.400 373.600 ;
        RECT 31.600 370.200 32.400 370.400 ;
        RECT 20.400 369.600 21.800 370.200 ;
        RECT 22.400 369.600 23.400 370.200 ;
        RECT 10.200 362.200 11.000 369.600 ;
        RECT 11.800 368.400 12.400 369.600 ;
        RECT 11.600 367.600 12.400 368.400 ;
        RECT 16.600 364.400 17.400 369.600 ;
        RECT 18.200 368.400 18.800 369.600 ;
        RECT 18.000 367.600 18.800 368.400 ;
        RECT 21.200 368.400 21.800 369.600 ;
        RECT 21.200 367.600 22.000 368.400 ;
        RECT 15.600 363.600 17.400 364.400 ;
        RECT 16.600 362.200 17.400 363.600 ;
        RECT 22.600 362.200 23.400 369.600 ;
        RECT 29.400 369.600 30.400 370.200 ;
        RECT 31.000 369.600 32.400 370.200 ;
        RECT 33.200 370.200 34.000 370.400 ;
        RECT 35.200 370.200 35.800 373.600 ;
        RECT 36.400 371.600 37.200 373.200 ;
        RECT 39.600 370.200 40.400 370.400 ;
        RECT 41.600 370.200 42.200 373.600 ;
        RECT 42.800 371.600 43.600 373.200 ;
        RECT 33.200 369.600 34.600 370.200 ;
        RECT 35.200 369.600 36.200 370.200 ;
        RECT 39.600 369.600 41.000 370.200 ;
        RECT 41.600 369.600 42.600 370.200 ;
        RECT 29.400 364.400 30.200 369.600 ;
        RECT 31.000 368.400 31.600 369.600 ;
        RECT 30.800 367.600 31.600 368.400 ;
        RECT 34.000 368.400 34.600 369.600 ;
        RECT 34.000 367.600 34.800 368.400 ;
        RECT 28.400 363.600 30.200 364.400 ;
        RECT 29.400 362.200 30.200 363.600 ;
        RECT 35.400 362.200 36.200 369.600 ;
        RECT 40.400 368.400 41.000 369.600 ;
        RECT 40.400 367.600 41.200 368.400 ;
        RECT 41.800 362.200 42.600 369.600 ;
        RECT 46.000 368.800 46.800 370.400 ;
        RECT 47.600 370.300 48.400 375.800 ;
        RECT 49.200 373.600 50.000 375.200 ;
        RECT 51.000 374.400 51.600 375.800 ;
        RECT 52.600 375.400 56.200 375.800 ;
        RECT 57.200 374.800 57.800 377.000 ;
        RECT 61.400 376.000 62.200 379.000 ;
        RECT 66.800 376.000 67.600 379.800 ;
        RECT 70.000 376.000 70.800 379.800 ;
        RECT 61.400 375.400 63.000 376.000 ;
        RECT 66.800 375.800 70.800 376.000 ;
        RECT 71.600 375.800 72.400 379.800 ;
        RECT 73.200 375.800 74.000 379.800 ;
        RECT 74.800 376.000 75.600 379.800 ;
        RECT 78.000 376.000 78.800 379.800 ;
        RECT 74.800 375.800 78.800 376.000 ;
        RECT 79.600 376.000 80.400 379.800 ;
        RECT 82.800 376.000 83.600 379.800 ;
        RECT 79.600 375.800 83.600 376.000 ;
        RECT 84.400 375.800 85.200 379.800 ;
        RECT 86.000 375.800 86.800 379.800 ;
        RECT 87.600 376.000 88.400 379.800 ;
        RECT 90.800 376.000 91.600 379.800 ;
        RECT 87.600 375.800 91.600 376.000 ;
        RECT 67.000 375.400 70.600 375.800 ;
        RECT 62.200 375.000 63.000 375.400 ;
        RECT 54.800 374.400 55.600 374.800 ;
        RECT 50.800 373.600 53.400 374.400 ;
        RECT 54.800 373.800 56.400 374.400 ;
        RECT 57.200 374.200 61.400 374.800 ;
        RECT 55.600 373.600 56.400 373.800 ;
        RECT 60.400 373.800 61.400 374.200 ;
        RECT 62.400 374.400 63.000 375.000 ;
        RECT 67.600 374.400 68.400 374.800 ;
        RECT 71.600 374.400 72.200 375.800 ;
        RECT 73.400 374.400 74.000 375.800 ;
        RECT 75.000 375.400 78.600 375.800 ;
        RECT 79.800 375.400 83.400 375.800 ;
        RECT 77.200 374.400 78.000 374.800 ;
        RECT 80.400 374.400 81.200 374.800 ;
        RECT 84.400 374.400 85.000 375.800 ;
        RECT 86.200 374.400 86.800 375.800 ;
        RECT 87.800 375.400 91.400 375.800 ;
        RECT 92.400 375.400 93.200 379.800 ;
        RECT 96.600 378.400 97.800 379.800 ;
        RECT 96.600 377.800 98.000 378.400 ;
        RECT 101.200 377.800 102.000 379.800 ;
        RECT 105.600 378.400 106.400 379.800 ;
        RECT 105.600 377.800 107.600 378.400 ;
        RECT 97.200 377.000 98.000 377.800 ;
        RECT 101.400 377.200 102.000 377.800 ;
        RECT 101.400 376.600 104.200 377.200 ;
        RECT 103.400 376.400 104.200 376.600 ;
        RECT 105.200 376.400 106.000 377.200 ;
        RECT 106.800 377.000 107.600 377.800 ;
        RECT 95.400 375.400 96.200 375.600 ;
        RECT 92.400 374.800 96.200 375.400 ;
        RECT 90.000 374.400 90.800 374.800 ;
        RECT 62.400 374.300 64.400 374.400 ;
        RECT 50.800 370.300 51.600 370.400 ;
        RECT 47.600 370.200 51.600 370.300 ;
        RECT 52.800 370.200 53.400 373.600 ;
        RECT 54.000 372.300 54.800 373.200 ;
        RECT 55.600 372.300 56.400 372.400 ;
        RECT 54.000 371.700 56.400 372.300 ;
        RECT 54.000 371.600 54.800 371.700 ;
        RECT 55.600 371.600 56.400 371.700 ;
        RECT 57.200 371.600 58.000 373.200 ;
        RECT 58.800 371.600 59.600 373.200 ;
        RECT 60.400 373.000 61.800 373.800 ;
        RECT 62.400 373.700 65.900 374.300 ;
        RECT 62.400 373.600 64.400 373.700 ;
        RECT 60.400 371.000 61.000 373.000 ;
        RECT 57.200 370.400 61.000 371.000 ;
        RECT 47.600 369.700 52.200 370.200 ;
        RECT 47.600 362.200 48.400 369.700 ;
        RECT 50.800 369.600 52.200 369.700 ;
        RECT 52.800 369.600 53.800 370.200 ;
        RECT 51.600 368.400 52.200 369.600 ;
        RECT 51.600 367.600 52.400 368.400 ;
        RECT 53.000 362.200 53.800 369.600 ;
        RECT 57.200 367.000 57.800 370.400 ;
        RECT 62.400 369.800 63.000 373.600 ;
        RECT 63.600 370.800 64.400 372.400 ;
        RECT 65.300 372.300 65.900 373.700 ;
        RECT 66.800 373.800 68.400 374.400 ;
        RECT 66.800 373.600 67.600 373.800 ;
        RECT 69.800 373.600 72.400 374.400 ;
        RECT 73.200 373.600 75.800 374.400 ;
        RECT 77.200 374.300 78.800 374.400 ;
        RECT 79.600 374.300 81.200 374.400 ;
        RECT 77.200 373.800 81.200 374.300 ;
        RECT 78.000 373.700 80.400 373.800 ;
        RECT 78.000 373.600 78.800 373.700 ;
        RECT 79.600 373.600 80.400 373.700 ;
        RECT 82.600 373.600 85.200 374.400 ;
        RECT 86.000 373.600 88.600 374.400 ;
        RECT 90.000 373.800 91.600 374.400 ;
        RECT 90.800 373.600 91.600 373.800 ;
        RECT 68.400 372.300 69.200 373.200 ;
        RECT 65.300 371.700 69.200 372.300 ;
        RECT 68.400 371.600 69.200 371.700 ;
        RECT 69.800 370.200 70.400 373.600 ;
        RECT 75.200 372.300 75.800 373.600 ;
        RECT 71.700 371.700 75.800 372.300 ;
        RECT 71.700 370.400 72.300 371.700 ;
        RECT 71.600 370.200 72.400 370.400 ;
        RECT 61.400 369.200 63.000 369.800 ;
        RECT 69.400 369.600 70.400 370.200 ;
        RECT 71.000 369.600 72.400 370.200 ;
        RECT 73.200 370.200 74.000 370.400 ;
        RECT 75.200 370.200 75.800 371.700 ;
        RECT 76.400 372.300 77.200 373.200 ;
        RECT 81.200 372.300 82.000 373.200 ;
        RECT 76.400 371.700 82.000 372.300 ;
        RECT 76.400 371.600 77.200 371.700 ;
        RECT 81.200 371.600 82.000 371.700 ;
        RECT 82.600 372.300 83.200 373.600 ;
        RECT 82.600 371.700 86.700 372.300 ;
        RECT 82.600 370.200 83.200 371.700 ;
        RECT 86.100 370.400 86.700 371.700 ;
        RECT 88.000 370.400 88.600 373.600 ;
        RECT 89.200 371.600 90.000 373.200 ;
        RECT 92.400 371.400 93.200 374.800 ;
        RECT 99.400 374.200 100.200 374.400 ;
        RECT 105.200 374.200 105.800 376.400 ;
        RECT 110.000 375.000 110.800 379.800 ;
        RECT 111.600 375.600 112.400 377.200 ;
        RECT 108.400 374.200 110.000 374.400 ;
        RECT 99.000 373.600 110.000 374.200 ;
        RECT 97.200 372.800 98.000 373.000 ;
        RECT 94.200 372.200 98.000 372.800 ;
        RECT 94.200 372.000 95.000 372.200 ;
        RECT 95.800 371.400 96.600 371.600 ;
        RECT 92.400 370.800 96.600 371.400 ;
        RECT 84.400 370.200 85.200 370.400 ;
        RECT 73.200 369.600 74.600 370.200 ;
        RECT 75.200 369.600 76.200 370.200 ;
        RECT 57.200 363.000 58.000 367.000 ;
        RECT 61.400 362.200 62.200 369.200 ;
        RECT 69.400 364.400 70.200 369.600 ;
        RECT 71.000 368.400 71.600 369.600 ;
        RECT 70.800 367.600 71.600 368.400 ;
        RECT 74.000 368.400 74.600 369.600 ;
        RECT 74.000 367.600 74.800 368.400 ;
        RECT 68.400 363.600 70.200 364.400 ;
        RECT 69.400 362.200 70.200 363.600 ;
        RECT 75.400 362.200 76.200 369.600 ;
        RECT 82.200 369.600 83.200 370.200 ;
        RECT 83.800 369.600 85.200 370.200 ;
        RECT 86.000 370.200 86.800 370.400 ;
        RECT 86.000 369.600 87.400 370.200 ;
        RECT 88.000 369.600 90.000 370.400 ;
        RECT 82.200 362.200 83.000 369.600 ;
        RECT 83.800 368.400 84.400 369.600 ;
        RECT 83.600 367.600 84.400 368.400 ;
        RECT 86.800 368.400 87.400 369.600 ;
        RECT 86.800 367.600 87.600 368.400 ;
        RECT 88.200 362.200 89.000 369.600 ;
        RECT 92.400 362.200 93.200 370.800 ;
        RECT 99.000 370.400 99.600 373.600 ;
        RECT 106.200 373.400 107.000 373.600 ;
        RECT 107.800 372.400 108.600 372.600 ;
        RECT 102.000 372.300 102.800 372.400 ;
        RECT 103.600 372.300 108.600 372.400 ;
        RECT 102.000 371.800 108.600 372.300 ;
        RECT 102.000 371.700 104.400 371.800 ;
        RECT 102.000 371.600 102.800 371.700 ;
        RECT 103.600 371.600 104.400 371.700 ;
        RECT 105.200 371.000 110.800 371.200 ;
        RECT 105.000 370.800 110.800 371.000 ;
        RECT 97.200 369.800 99.600 370.400 ;
        RECT 101.000 370.600 110.800 370.800 ;
        RECT 101.000 370.200 105.800 370.600 ;
        RECT 97.200 368.800 97.800 369.800 ;
        RECT 96.400 368.000 97.800 368.800 ;
        RECT 99.400 369.000 100.200 369.200 ;
        RECT 101.000 369.000 101.600 370.200 ;
        RECT 99.400 368.400 101.600 369.000 ;
        RECT 102.200 369.000 107.600 369.600 ;
        RECT 102.200 368.800 103.000 369.000 ;
        RECT 106.800 368.800 107.600 369.000 ;
        RECT 100.600 367.400 101.400 367.600 ;
        RECT 103.400 367.400 104.200 367.600 ;
        RECT 97.200 366.200 98.000 367.000 ;
        RECT 100.600 366.800 104.200 367.400 ;
        RECT 101.400 366.200 102.000 366.800 ;
        RECT 106.800 366.200 107.600 367.000 ;
        RECT 96.600 362.200 97.800 366.200 ;
        RECT 101.200 362.200 102.000 366.200 ;
        RECT 105.600 365.600 107.600 366.200 ;
        RECT 105.600 362.200 106.400 365.600 ;
        RECT 110.000 362.200 110.800 370.600 ;
        RECT 113.200 370.300 114.000 379.800 ;
        RECT 114.800 375.800 115.600 379.800 ;
        RECT 116.400 376.000 117.200 379.800 ;
        RECT 119.600 376.000 120.400 379.800 ;
        RECT 116.400 375.800 120.400 376.000 ;
        RECT 121.200 376.000 122.000 379.800 ;
        RECT 124.400 376.000 125.200 379.800 ;
        RECT 121.200 375.800 125.200 376.000 ;
        RECT 126.000 375.800 126.800 379.800 ;
        RECT 127.600 377.000 128.400 379.000 ;
        RECT 115.000 374.400 115.600 375.800 ;
        RECT 116.600 375.400 120.200 375.800 ;
        RECT 121.400 375.400 125.000 375.800 ;
        RECT 118.800 374.400 119.600 374.800 ;
        RECT 122.000 374.400 122.800 374.800 ;
        RECT 126.000 374.400 126.600 375.800 ;
        RECT 127.600 374.800 128.200 377.000 ;
        RECT 131.800 376.000 132.600 379.000 ;
        RECT 137.200 376.000 138.000 379.800 ;
        RECT 140.400 376.000 141.200 379.800 ;
        RECT 131.800 375.400 133.400 376.000 ;
        RECT 137.200 375.800 141.200 376.000 ;
        RECT 142.000 375.800 142.800 379.800 ;
        RECT 143.600 376.000 144.400 379.800 ;
        RECT 146.800 376.000 147.600 379.800 ;
        RECT 143.600 375.800 147.600 376.000 ;
        RECT 148.400 375.800 149.200 379.800 ;
        RECT 137.400 375.400 141.000 375.800 ;
        RECT 132.600 375.000 133.400 375.400 ;
        RECT 114.800 373.600 117.400 374.400 ;
        RECT 118.800 373.800 120.400 374.400 ;
        RECT 119.600 373.600 120.400 373.800 ;
        RECT 121.200 373.800 122.800 374.400 ;
        RECT 121.200 373.600 122.000 373.800 ;
        RECT 124.200 373.600 126.800 374.400 ;
        RECT 127.600 374.200 131.800 374.800 ;
        RECT 130.800 373.800 131.800 374.200 ;
        RECT 132.800 374.400 133.400 375.000 ;
        RECT 138.000 374.400 138.800 374.800 ;
        RECT 142.000 374.400 142.600 375.800 ;
        RECT 143.800 375.400 147.400 375.800 ;
        RECT 144.400 374.400 145.200 374.800 ;
        RECT 148.400 374.400 149.000 375.800 ;
        RECT 154.800 375.000 155.600 379.800 ;
        RECT 159.200 378.400 160.000 379.800 ;
        RECT 158.000 377.800 160.000 378.400 ;
        RECT 163.600 377.800 164.400 379.800 ;
        RECT 167.800 378.400 169.000 379.800 ;
        RECT 167.600 377.800 169.000 378.400 ;
        RECT 158.000 377.000 158.800 377.800 ;
        RECT 163.600 377.200 164.200 377.800 ;
        RECT 159.600 376.400 160.400 377.200 ;
        RECT 161.400 376.600 164.200 377.200 ;
        RECT 167.600 377.000 168.400 377.800 ;
        RECT 161.400 376.400 162.200 376.600 ;
        RECT 114.800 370.300 115.600 370.400 ;
        RECT 113.200 370.200 115.600 370.300 ;
        RECT 116.800 370.200 117.400 373.600 ;
        RECT 118.000 371.600 118.800 373.200 ;
        RECT 122.800 371.600 123.600 373.200 ;
        RECT 124.200 370.200 124.800 373.600 ;
        RECT 127.600 371.600 128.400 373.200 ;
        RECT 129.200 371.600 130.000 373.200 ;
        RECT 130.800 373.000 132.200 373.800 ;
        RECT 132.800 373.600 134.800 374.400 ;
        RECT 137.200 373.800 138.800 374.400 ;
        RECT 137.200 373.600 138.000 373.800 ;
        RECT 140.200 373.600 142.800 374.400 ;
        RECT 143.600 373.800 145.200 374.400 ;
        RECT 143.600 373.600 144.400 373.800 ;
        RECT 146.600 373.600 149.200 374.400 ;
        RECT 155.600 374.200 157.200 374.400 ;
        RECT 159.800 374.200 160.400 376.400 ;
        RECT 169.400 375.400 170.200 375.600 ;
        RECT 172.400 375.400 173.200 379.800 ;
        RECT 169.400 374.800 173.200 375.400 ;
        RECT 165.400 374.200 166.800 374.400 ;
        RECT 155.600 373.600 166.800 374.200 ;
        RECT 130.800 371.000 131.400 373.000 ;
        RECT 127.600 370.400 131.400 371.000 ;
        RECT 126.000 370.200 126.800 370.400 ;
        RECT 113.200 369.700 116.200 370.200 ;
        RECT 113.200 362.200 114.000 369.700 ;
        RECT 114.800 369.600 116.200 369.700 ;
        RECT 116.800 369.600 117.800 370.200 ;
        RECT 115.600 368.400 116.200 369.600 ;
        RECT 115.600 367.600 116.400 368.400 ;
        RECT 117.000 362.200 117.800 369.600 ;
        RECT 123.800 369.600 124.800 370.200 ;
        RECT 125.400 369.600 126.800 370.200 ;
        RECT 123.800 364.400 124.600 369.600 ;
        RECT 125.400 368.400 126.000 369.600 ;
        RECT 125.200 367.600 126.000 368.400 ;
        RECT 122.800 363.600 124.600 364.400 ;
        RECT 123.800 362.200 124.600 363.600 ;
        RECT 127.600 367.000 128.200 370.400 ;
        RECT 132.800 369.800 133.400 373.600 ;
        RECT 134.000 372.300 134.800 372.400 ;
        RECT 137.200 372.300 138.000 372.400 ;
        RECT 134.000 371.700 138.000 372.300 ;
        RECT 134.000 370.800 134.800 371.700 ;
        RECT 137.200 371.600 138.000 371.700 ;
        RECT 138.800 371.600 139.600 373.200 ;
        RECT 140.200 370.200 140.800 373.600 ;
        RECT 145.200 371.600 146.000 373.200 ;
        RECT 146.600 372.300 147.200 373.600 ;
        RECT 158.600 373.400 159.400 373.600 ;
        RECT 157.000 372.400 157.800 372.600 ;
        RECT 159.600 372.400 160.400 372.600 ;
        RECT 153.200 372.300 154.000 372.400 ;
        RECT 146.600 371.700 154.000 372.300 ;
        RECT 157.000 371.800 162.000 372.400 ;
        RECT 142.000 370.200 142.800 370.400 ;
        RECT 146.600 370.200 147.200 371.700 ;
        RECT 153.200 371.600 154.000 371.700 ;
        RECT 161.200 371.600 162.000 371.800 ;
        RECT 154.800 371.000 160.400 371.200 ;
        RECT 154.800 370.800 160.600 371.000 ;
        RECT 154.800 370.600 164.600 370.800 ;
        RECT 148.400 370.200 149.200 370.400 ;
        RECT 131.800 369.200 133.400 369.800 ;
        RECT 139.800 369.600 140.800 370.200 ;
        RECT 141.400 369.600 142.800 370.200 ;
        RECT 146.200 369.600 147.200 370.200 ;
        RECT 147.800 369.600 149.200 370.200 ;
        RECT 131.800 368.400 132.600 369.200 ;
        RECT 131.800 367.600 133.200 368.400 ;
        RECT 127.600 363.000 128.400 367.000 ;
        RECT 131.800 362.200 132.600 367.600 ;
        RECT 139.800 362.200 140.600 369.600 ;
        RECT 141.400 368.400 142.000 369.600 ;
        RECT 141.200 367.600 142.000 368.400 ;
        RECT 146.200 362.200 147.000 369.600 ;
        RECT 147.800 368.400 148.400 369.600 ;
        RECT 147.600 367.600 148.400 368.400 ;
        RECT 154.800 362.200 155.600 370.600 ;
        RECT 159.800 370.200 164.600 370.600 ;
        RECT 158.000 369.000 163.400 369.600 ;
        RECT 158.000 368.800 158.800 369.000 ;
        RECT 162.600 368.800 163.400 369.000 ;
        RECT 164.000 369.000 164.600 370.200 ;
        RECT 166.000 370.400 166.600 373.600 ;
        RECT 167.600 372.800 168.400 373.000 ;
        RECT 167.600 372.200 171.400 372.800 ;
        RECT 170.600 372.000 171.400 372.200 ;
        RECT 169.000 371.400 169.800 371.600 ;
        RECT 172.400 371.400 173.200 374.800 ;
        RECT 169.000 370.800 173.200 371.400 ;
        RECT 166.000 369.800 168.400 370.400 ;
        RECT 165.400 369.000 166.200 369.200 ;
        RECT 164.000 368.400 166.200 369.000 ;
        RECT 167.800 368.800 168.400 369.800 ;
        RECT 167.800 368.000 169.200 368.800 ;
        RECT 161.400 367.400 162.200 367.600 ;
        RECT 164.200 367.400 165.000 367.600 ;
        RECT 158.000 366.200 158.800 367.000 ;
        RECT 161.400 366.800 165.000 367.400 ;
        RECT 163.600 366.200 164.200 366.800 ;
        RECT 167.600 366.200 168.400 367.000 ;
        RECT 158.000 365.600 160.000 366.200 ;
        RECT 159.200 362.200 160.000 365.600 ;
        RECT 163.600 362.200 164.400 366.200 ;
        RECT 167.800 362.200 169.000 366.200 ;
        RECT 172.400 362.200 173.200 370.800 ;
        RECT 174.000 373.800 174.800 379.800 ;
        RECT 180.400 376.600 181.200 379.800 ;
        RECT 182.000 377.000 182.800 379.800 ;
        RECT 183.600 377.000 184.400 379.800 ;
        RECT 185.200 377.000 186.000 379.800 ;
        RECT 188.400 377.000 189.200 379.800 ;
        RECT 191.600 377.000 192.400 379.800 ;
        RECT 193.200 377.000 194.000 379.800 ;
        RECT 194.800 377.000 195.600 379.800 ;
        RECT 196.400 377.000 197.200 379.800 ;
        RECT 178.600 375.800 181.200 376.600 ;
        RECT 198.000 376.600 198.800 379.800 ;
        RECT 184.600 375.800 189.200 376.400 ;
        RECT 178.600 375.200 179.400 375.800 ;
        RECT 176.400 374.400 179.400 375.200 ;
        RECT 174.000 373.000 182.800 373.800 ;
        RECT 184.600 373.400 185.400 375.800 ;
        RECT 188.400 375.600 189.200 375.800 ;
        RECT 190.000 375.600 191.600 376.400 ;
        RECT 194.600 375.600 195.600 376.400 ;
        RECT 198.000 375.800 200.400 376.600 ;
        RECT 186.800 373.600 187.600 375.200 ;
        RECT 188.400 374.800 189.200 375.000 ;
        RECT 188.400 374.200 192.800 374.800 ;
        RECT 192.000 374.000 192.800 374.200 ;
        RECT 174.000 367.400 174.800 373.000 ;
        RECT 183.400 372.600 185.400 373.400 ;
        RECT 189.200 372.600 192.400 373.400 ;
        RECT 194.800 372.800 195.600 375.600 ;
        RECT 199.600 375.200 200.400 375.800 ;
        RECT 199.600 374.600 201.400 375.200 ;
        RECT 200.600 373.400 201.400 374.600 ;
        RECT 204.400 374.600 205.200 379.800 ;
        RECT 206.000 376.000 206.800 379.800 ;
        RECT 209.800 376.400 210.600 379.800 ;
        RECT 206.000 375.200 207.000 376.000 ;
        RECT 209.800 375.800 211.600 376.400 ;
        RECT 214.000 375.800 214.800 379.800 ;
        RECT 215.600 376.000 216.400 379.800 ;
        RECT 218.800 376.000 219.600 379.800 ;
        RECT 215.600 375.800 219.600 376.000 ;
        RECT 220.400 375.800 221.200 379.800 ;
        RECT 222.000 376.000 222.800 379.800 ;
        RECT 225.200 376.000 226.000 379.800 ;
        RECT 222.000 375.800 226.000 376.000 ;
        RECT 226.800 376.000 227.600 379.800 ;
        RECT 230.000 376.000 230.800 379.800 ;
        RECT 226.800 375.800 230.800 376.000 ;
        RECT 231.600 375.800 232.400 379.800 ;
        RECT 234.800 376.000 235.600 379.800 ;
        RECT 204.400 374.000 205.600 374.600 ;
        RECT 200.600 372.600 204.400 373.400 ;
        RECT 175.400 372.000 176.200 372.200 ;
        RECT 180.400 372.000 181.200 372.400 ;
        RECT 198.000 372.000 198.800 372.600 ;
        RECT 205.000 372.000 205.600 374.000 ;
        RECT 175.400 371.400 198.800 372.000 ;
        RECT 204.800 371.400 205.600 372.000 ;
        RECT 204.800 369.600 205.400 371.400 ;
        RECT 206.200 370.800 207.000 375.200 ;
        RECT 183.600 369.400 184.400 369.600 ;
        RECT 179.000 369.000 184.400 369.400 ;
        RECT 178.200 368.800 184.400 369.000 ;
        RECT 185.400 369.000 194.000 369.600 ;
        RECT 175.600 368.000 177.200 368.800 ;
        RECT 178.200 368.200 179.600 368.800 ;
        RECT 185.400 368.200 186.000 369.000 ;
        RECT 193.200 368.800 194.000 369.000 ;
        RECT 196.400 369.000 205.400 369.600 ;
        RECT 196.400 368.800 197.200 369.000 ;
        RECT 176.600 367.600 177.200 368.000 ;
        RECT 180.200 367.600 186.000 368.200 ;
        RECT 186.600 367.600 189.200 368.400 ;
        RECT 174.000 366.800 176.000 367.400 ;
        RECT 176.600 366.800 180.800 367.600 ;
        RECT 175.400 366.200 176.000 366.800 ;
        RECT 175.400 365.600 176.400 366.200 ;
        RECT 175.600 362.200 176.400 365.600 ;
        RECT 178.800 362.200 179.600 366.800 ;
        RECT 182.000 362.200 182.800 365.000 ;
        RECT 183.600 362.200 184.400 365.000 ;
        RECT 185.200 362.200 186.000 367.000 ;
        RECT 188.400 362.200 189.200 367.000 ;
        RECT 191.600 362.200 192.400 368.400 ;
        RECT 199.600 367.600 202.200 368.400 ;
        RECT 194.800 366.800 199.000 367.600 ;
        RECT 193.200 362.200 194.000 365.000 ;
        RECT 194.800 362.200 195.600 365.000 ;
        RECT 196.400 362.200 197.200 365.000 ;
        RECT 199.600 362.200 200.400 367.600 ;
        RECT 204.800 367.400 205.400 369.000 ;
        RECT 202.800 366.800 205.400 367.400 ;
        RECT 206.000 370.000 207.000 370.800 ;
        RECT 202.800 362.200 203.600 366.800 ;
        RECT 206.000 362.200 206.800 370.000 ;
        RECT 209.200 368.800 210.000 370.400 ;
        RECT 210.800 362.200 211.600 375.800 ;
        RECT 212.400 373.600 213.200 375.200 ;
        RECT 214.200 374.400 214.800 375.800 ;
        RECT 215.800 375.400 219.400 375.800 ;
        RECT 218.000 374.400 218.800 374.800 ;
        RECT 220.600 374.400 221.200 375.800 ;
        RECT 222.200 375.400 225.800 375.800 ;
        RECT 227.000 375.400 230.600 375.800 ;
        RECT 224.400 374.400 225.200 374.800 ;
        RECT 227.600 374.400 228.400 374.800 ;
        RECT 231.600 374.400 232.200 375.800 ;
        RECT 234.600 375.200 235.600 376.000 ;
        RECT 214.000 373.600 216.600 374.400 ;
        RECT 218.000 373.800 219.600 374.400 ;
        RECT 218.800 373.600 219.600 373.800 ;
        RECT 220.400 373.600 223.000 374.400 ;
        RECT 224.400 374.300 226.000 374.400 ;
        RECT 226.800 374.300 228.400 374.400 ;
        RECT 224.400 373.800 228.400 374.300 ;
        RECT 225.200 373.700 227.600 373.800 ;
        RECT 225.200 373.600 226.000 373.700 ;
        RECT 226.800 373.600 227.600 373.700 ;
        RECT 229.800 373.600 232.400 374.400 ;
        RECT 212.400 370.300 213.200 370.400 ;
        RECT 214.000 370.300 214.800 370.400 ;
        RECT 212.400 370.200 214.800 370.300 ;
        RECT 216.000 370.200 216.600 373.600 ;
        RECT 217.200 372.300 218.000 373.200 ;
        RECT 218.800 372.300 219.600 372.400 ;
        RECT 217.200 371.700 219.600 372.300 ;
        RECT 217.200 371.600 218.000 371.700 ;
        RECT 218.800 371.600 219.600 371.700 ;
        RECT 220.400 370.200 221.200 370.400 ;
        RECT 222.400 370.200 223.000 373.600 ;
        RECT 223.600 372.300 224.400 373.200 ;
        RECT 228.400 372.300 229.200 373.200 ;
        RECT 223.600 371.700 229.200 372.300 ;
        RECT 223.600 371.600 224.400 371.700 ;
        RECT 228.400 371.600 229.200 371.700 ;
        RECT 229.800 370.200 230.400 373.600 ;
        RECT 234.600 370.800 235.400 375.200 ;
        RECT 236.400 374.600 237.200 379.800 ;
        RECT 242.800 376.600 243.600 379.800 ;
        RECT 244.400 377.000 245.200 379.800 ;
        RECT 246.000 377.000 246.800 379.800 ;
        RECT 247.600 377.000 248.400 379.800 ;
        RECT 249.200 377.000 250.000 379.800 ;
        RECT 252.400 377.000 253.200 379.800 ;
        RECT 255.600 377.000 256.400 379.800 ;
        RECT 257.200 377.000 258.000 379.800 ;
        RECT 258.800 377.000 259.600 379.800 ;
        RECT 241.200 375.800 243.600 376.600 ;
        RECT 260.400 376.600 261.200 379.800 ;
        RECT 241.200 375.200 242.000 375.800 ;
        RECT 236.000 374.000 237.200 374.600 ;
        RECT 240.200 374.600 242.000 375.200 ;
        RECT 246.000 375.600 247.000 376.400 ;
        RECT 250.000 375.600 251.600 376.400 ;
        RECT 252.400 375.800 257.000 376.400 ;
        RECT 260.400 375.800 263.000 376.600 ;
        RECT 252.400 375.600 253.200 375.800 ;
        RECT 236.000 372.000 236.600 374.000 ;
        RECT 240.200 373.400 241.000 374.600 ;
        RECT 237.200 372.600 241.000 373.400 ;
        RECT 246.000 372.800 246.800 375.600 ;
        RECT 252.400 374.800 253.200 375.000 ;
        RECT 248.800 374.200 253.200 374.800 ;
        RECT 248.800 374.000 249.600 374.200 ;
        RECT 254.000 373.600 254.800 375.200 ;
        RECT 256.200 373.400 257.000 375.800 ;
        RECT 262.200 375.200 263.000 375.800 ;
        RECT 262.200 374.400 265.200 375.200 ;
        RECT 266.800 373.800 267.600 379.800 ;
        RECT 270.000 376.400 270.800 379.800 ;
        RECT 249.200 372.600 252.400 373.400 ;
        RECT 256.200 372.600 258.200 373.400 ;
        RECT 258.800 373.000 267.600 373.800 ;
        RECT 242.800 372.000 243.600 372.600 ;
        RECT 260.400 372.000 261.200 372.400 ;
        RECT 263.600 372.000 264.400 372.400 ;
        RECT 265.400 372.000 266.200 372.200 ;
        RECT 236.000 371.400 236.800 372.000 ;
        RECT 242.800 371.400 266.200 372.000 ;
        RECT 231.600 370.300 232.400 370.400 ;
        RECT 234.600 370.300 235.600 370.800 ;
        RECT 231.600 370.200 235.600 370.300 ;
        RECT 212.400 369.700 215.400 370.200 ;
        RECT 212.400 369.600 213.200 369.700 ;
        RECT 214.000 369.600 215.400 369.700 ;
        RECT 216.000 369.600 217.000 370.200 ;
        RECT 220.400 369.600 221.800 370.200 ;
        RECT 222.400 369.600 223.400 370.200 ;
        RECT 214.800 368.400 215.400 369.600 ;
        RECT 214.800 367.600 215.600 368.400 ;
        RECT 216.200 362.200 217.000 369.600 ;
        RECT 221.200 368.400 221.800 369.600 ;
        RECT 220.400 367.600 222.000 368.400 ;
        RECT 222.600 362.200 223.400 369.600 ;
        RECT 229.400 369.600 230.400 370.200 ;
        RECT 231.000 369.700 235.600 370.200 ;
        RECT 231.000 369.600 232.400 369.700 ;
        RECT 229.400 362.200 230.200 369.600 ;
        RECT 231.000 368.400 231.600 369.600 ;
        RECT 230.800 367.600 232.400 368.400 ;
        RECT 234.800 362.200 235.600 369.700 ;
        RECT 236.200 369.600 236.800 371.400 ;
        RECT 236.200 369.000 245.200 369.600 ;
        RECT 236.200 367.400 236.800 369.000 ;
        RECT 244.400 368.800 245.200 369.000 ;
        RECT 247.600 369.000 256.200 369.600 ;
        RECT 247.600 368.800 248.400 369.000 ;
        RECT 239.400 367.600 242.000 368.400 ;
        RECT 236.200 366.800 238.800 367.400 ;
        RECT 238.000 362.200 238.800 366.800 ;
        RECT 241.200 362.200 242.000 367.600 ;
        RECT 242.600 366.800 246.800 367.600 ;
        RECT 244.400 362.200 245.200 365.000 ;
        RECT 246.000 362.200 246.800 365.000 ;
        RECT 247.600 362.200 248.400 365.000 ;
        RECT 249.200 362.200 250.000 368.400 ;
        RECT 252.400 367.600 255.000 368.400 ;
        RECT 255.600 368.200 256.200 369.000 ;
        RECT 257.200 369.400 258.000 369.600 ;
        RECT 257.200 369.000 262.600 369.400 ;
        RECT 257.200 368.800 263.400 369.000 ;
        RECT 262.000 368.200 263.400 368.800 ;
        RECT 255.600 367.600 261.400 368.200 ;
        RECT 264.400 368.000 266.000 368.800 ;
        RECT 264.400 367.600 265.000 368.000 ;
        RECT 252.400 362.200 253.200 367.000 ;
        RECT 255.600 362.200 256.400 367.000 ;
        RECT 260.800 366.800 265.000 367.600 ;
        RECT 266.800 367.400 267.600 373.000 ;
        RECT 269.800 375.800 270.800 376.400 ;
        RECT 269.800 374.400 270.400 375.800 ;
        RECT 273.200 375.200 274.000 379.800 ;
        RECT 271.400 374.600 274.000 375.200 ;
        RECT 276.400 375.200 277.200 379.800 ;
        RECT 279.600 375.200 280.400 379.800 ;
        RECT 282.800 375.200 283.600 379.800 ;
        RECT 286.000 375.200 286.800 379.800 ;
        RECT 290.800 375.200 291.600 379.800 ;
        RECT 294.000 375.200 294.800 379.800 ;
        RECT 297.200 375.200 298.000 379.800 ;
        RECT 300.400 375.200 301.200 379.800 ;
        RECT 308.400 377.000 309.200 379.000 ;
        RECT 312.600 378.400 313.400 379.000 ;
        RECT 312.600 377.600 314.000 378.400 ;
        RECT 269.800 373.600 270.800 374.400 ;
        RECT 269.800 370.200 270.400 373.600 ;
        RECT 271.400 373.000 272.000 374.600 ;
        RECT 276.400 374.400 278.200 375.200 ;
        RECT 279.600 374.400 281.800 375.200 ;
        RECT 282.800 374.400 285.000 375.200 ;
        RECT 286.000 374.400 288.400 375.200 ;
        RECT 290.800 374.400 292.600 375.200 ;
        RECT 294.000 374.400 296.200 375.200 ;
        RECT 297.200 374.400 299.400 375.200 ;
        RECT 300.400 374.400 302.800 375.200 ;
        RECT 274.800 373.800 275.600 374.400 ;
        RECT 277.400 373.800 278.200 374.400 ;
        RECT 281.000 373.800 281.800 374.400 ;
        RECT 284.200 373.800 285.000 374.400 ;
        RECT 274.800 373.000 276.600 373.800 ;
        RECT 277.400 373.000 280.000 373.800 ;
        RECT 281.000 373.000 283.400 373.800 ;
        RECT 284.200 373.000 286.800 373.800 ;
        RECT 271.000 372.200 272.000 373.000 ;
        RECT 271.400 370.200 272.000 372.200 ;
        RECT 277.400 371.600 278.200 373.000 ;
        RECT 281.000 371.600 281.800 373.000 ;
        RECT 284.200 371.600 285.000 373.000 ;
        RECT 287.600 371.600 288.400 374.400 ;
        RECT 289.200 373.800 290.000 374.400 ;
        RECT 291.800 373.800 292.600 374.400 ;
        RECT 295.400 373.800 296.200 374.400 ;
        RECT 298.600 373.800 299.400 374.400 ;
        RECT 289.200 373.000 291.000 373.800 ;
        RECT 291.800 373.000 294.400 373.800 ;
        RECT 295.400 373.000 297.800 373.800 ;
        RECT 298.600 373.000 301.200 373.800 ;
        RECT 291.800 371.600 292.600 373.000 ;
        RECT 295.400 371.600 296.200 373.000 ;
        RECT 298.600 371.600 299.400 373.000 ;
        RECT 302.000 371.600 302.800 374.400 ;
        RECT 308.400 374.800 309.000 377.000 ;
        RECT 312.600 376.000 313.400 377.600 ;
        RECT 312.600 375.400 314.200 376.000 ;
        RECT 313.400 375.000 314.200 375.400 ;
        RECT 308.400 374.200 312.600 374.800 ;
        RECT 311.600 373.800 312.600 374.200 ;
        RECT 313.600 374.400 314.200 375.000 ;
        RECT 308.400 371.600 309.200 373.200 ;
        RECT 310.000 371.600 310.800 373.200 ;
        RECT 311.600 373.000 313.000 373.800 ;
        RECT 313.600 373.600 315.600 374.400 ;
        RECT 276.400 370.800 278.200 371.600 ;
        RECT 279.600 370.800 281.800 371.600 ;
        RECT 282.800 370.800 285.000 371.600 ;
        RECT 286.000 370.800 288.400 371.600 ;
        RECT 290.800 370.800 292.600 371.600 ;
        RECT 294.000 370.800 296.200 371.600 ;
        RECT 297.200 370.800 299.400 371.600 ;
        RECT 300.400 370.800 302.800 371.600 ;
        RECT 311.600 371.000 312.200 373.000 ;
        RECT 269.800 369.200 270.800 370.200 ;
        RECT 271.400 369.600 274.000 370.200 ;
        RECT 265.600 366.800 267.600 367.400 ;
        RECT 257.200 362.200 258.000 365.000 ;
        RECT 258.800 362.200 259.600 365.000 ;
        RECT 262.000 362.200 262.800 366.800 ;
        RECT 265.600 366.200 266.200 366.800 ;
        RECT 265.200 365.600 266.200 366.200 ;
        RECT 265.200 362.200 266.000 365.600 ;
        RECT 270.000 362.200 270.800 369.200 ;
        RECT 273.200 362.200 274.000 369.600 ;
        RECT 276.400 362.200 277.200 370.800 ;
        RECT 279.600 362.200 280.400 370.800 ;
        RECT 282.800 362.200 283.600 370.800 ;
        RECT 286.000 362.200 286.800 370.800 ;
        RECT 290.800 362.200 291.600 370.800 ;
        RECT 294.000 362.200 294.800 370.800 ;
        RECT 297.200 362.200 298.000 370.800 ;
        RECT 300.400 362.200 301.200 370.800 ;
        RECT 308.400 370.400 312.200 371.000 ;
        RECT 308.400 367.000 309.000 370.400 ;
        RECT 313.600 369.800 314.200 373.600 ;
        RECT 314.800 372.300 315.600 372.400 ;
        RECT 318.000 372.300 318.800 379.800 ;
        RECT 319.600 375.600 320.400 377.200 ;
        RECT 321.200 375.800 322.000 379.800 ;
        RECT 322.800 376.000 323.600 379.800 ;
        RECT 326.000 376.000 326.800 379.800 ;
        RECT 322.800 375.800 326.800 376.000 ;
        RECT 321.400 374.400 322.000 375.800 ;
        RECT 323.000 375.400 326.600 375.800 ;
        RECT 325.200 374.400 326.000 374.800 ;
        RECT 321.200 373.600 323.800 374.400 ;
        RECT 325.200 374.300 326.800 374.400 ;
        RECT 327.600 374.300 328.400 379.800 ;
        RECT 329.200 375.600 330.000 377.200 ;
        RECT 330.800 377.000 331.600 379.000 ;
        RECT 325.200 373.800 328.400 374.300 ;
        RECT 330.800 374.800 331.400 377.000 ;
        RECT 335.000 376.000 335.800 379.000 ;
        RECT 335.000 375.400 336.600 376.000 ;
        RECT 335.800 375.000 336.600 375.400 ;
        RECT 330.800 374.200 335.000 374.800 ;
        RECT 326.000 373.700 328.400 373.800 ;
        RECT 326.000 373.600 326.800 373.700 ;
        RECT 314.800 371.700 318.800 372.300 ;
        RECT 314.800 370.800 315.600 371.700 ;
        RECT 312.600 369.200 314.200 369.800 ;
        RECT 308.400 363.000 309.200 367.000 ;
        RECT 312.600 362.200 313.400 369.200 ;
        RECT 318.000 362.200 318.800 371.700 ;
        RECT 321.200 370.200 322.000 370.400 ;
        RECT 323.200 370.200 323.800 373.600 ;
        RECT 324.400 372.300 325.200 373.200 ;
        RECT 326.000 372.300 326.800 372.400 ;
        RECT 324.400 371.700 326.800 372.300 ;
        RECT 324.400 371.600 325.200 371.700 ;
        RECT 326.000 371.600 326.800 371.700 ;
        RECT 321.200 369.600 322.600 370.200 ;
        RECT 323.200 369.600 324.200 370.200 ;
        RECT 322.000 368.400 322.600 369.600 ;
        RECT 322.000 367.600 322.800 368.400 ;
        RECT 323.400 362.200 324.200 369.600 ;
        RECT 327.600 362.200 328.400 373.700 ;
        RECT 334.000 373.800 335.000 374.200 ;
        RECT 336.000 374.400 336.600 375.000 ;
        RECT 336.000 374.300 338.000 374.400 ;
        RECT 338.800 374.300 339.600 374.400 ;
        RECT 330.800 371.600 331.600 373.200 ;
        RECT 332.400 371.600 333.200 373.200 ;
        RECT 334.000 373.000 335.400 373.800 ;
        RECT 336.000 373.700 339.600 374.300 ;
        RECT 336.000 373.600 338.000 373.700 ;
        RECT 338.800 373.600 339.600 373.700 ;
        RECT 334.000 371.000 334.600 373.000 ;
        RECT 330.800 370.400 334.600 371.000 ;
        RECT 330.800 367.000 331.400 370.400 ;
        RECT 336.000 369.800 336.600 373.600 ;
        RECT 337.200 372.300 338.000 372.400 ;
        RECT 340.400 372.300 341.200 379.800 ;
        RECT 342.000 375.600 342.800 377.200 ;
        RECT 337.200 371.700 341.200 372.300 ;
        RECT 337.200 370.800 338.000 371.700 ;
        RECT 335.000 369.200 336.600 369.800 ;
        RECT 330.800 363.000 331.600 367.000 ;
        RECT 335.000 362.200 335.800 369.200 ;
        RECT 340.400 362.200 341.200 371.700 ;
        RECT 343.600 373.800 344.400 379.800 ;
        RECT 350.000 376.600 350.800 379.800 ;
        RECT 351.600 377.000 352.400 379.800 ;
        RECT 353.200 377.000 354.000 379.800 ;
        RECT 354.800 377.000 355.600 379.800 ;
        RECT 358.000 377.000 358.800 379.800 ;
        RECT 361.200 377.000 362.000 379.800 ;
        RECT 362.800 377.000 363.600 379.800 ;
        RECT 364.400 377.000 365.200 379.800 ;
        RECT 366.000 377.000 366.800 379.800 ;
        RECT 348.200 375.800 350.800 376.600 ;
        RECT 367.600 376.600 368.400 379.800 ;
        RECT 354.200 375.800 358.800 376.400 ;
        RECT 348.200 375.200 349.000 375.800 ;
        RECT 346.000 374.400 349.000 375.200 ;
        RECT 343.600 373.000 352.400 373.800 ;
        RECT 354.200 373.400 355.000 375.800 ;
        RECT 358.000 375.600 358.800 375.800 ;
        RECT 359.600 375.600 361.200 376.400 ;
        RECT 364.200 375.600 365.200 376.400 ;
        RECT 367.600 375.800 370.000 376.600 ;
        RECT 356.400 373.600 357.200 375.200 ;
        RECT 358.000 374.800 358.800 375.000 ;
        RECT 358.000 374.200 362.400 374.800 ;
        RECT 361.600 374.000 362.400 374.200 ;
        RECT 343.600 367.400 344.400 373.000 ;
        RECT 353.000 372.600 355.000 373.400 ;
        RECT 358.800 372.600 362.000 373.400 ;
        RECT 364.400 372.800 365.200 375.600 ;
        RECT 369.200 375.200 370.000 375.800 ;
        RECT 369.200 374.600 371.000 375.200 ;
        RECT 370.200 373.400 371.000 374.600 ;
        RECT 374.000 374.600 374.800 379.800 ;
        RECT 375.600 376.000 376.400 379.800 ;
        RECT 380.400 376.000 381.200 379.800 ;
        RECT 375.600 375.200 376.600 376.000 ;
        RECT 374.000 374.000 375.200 374.600 ;
        RECT 370.200 372.600 374.000 373.400 ;
        RECT 345.000 372.000 345.800 372.200 ;
        RECT 346.800 372.000 347.600 372.400 ;
        RECT 350.000 372.000 350.800 372.400 ;
        RECT 367.600 372.000 368.400 372.600 ;
        RECT 374.600 372.000 375.200 374.000 ;
        RECT 345.000 371.400 368.400 372.000 ;
        RECT 374.400 371.400 375.200 372.000 ;
        RECT 374.400 369.600 375.000 371.400 ;
        RECT 375.800 370.800 376.600 375.200 ;
        RECT 353.200 369.400 354.000 369.600 ;
        RECT 348.600 369.000 354.000 369.400 ;
        RECT 347.800 368.800 354.000 369.000 ;
        RECT 355.000 369.000 363.600 369.600 ;
        RECT 345.200 368.000 346.800 368.800 ;
        RECT 347.800 368.200 349.200 368.800 ;
        RECT 355.000 368.200 355.600 369.000 ;
        RECT 362.800 368.800 363.600 369.000 ;
        RECT 366.000 369.000 375.000 369.600 ;
        RECT 366.000 368.800 366.800 369.000 ;
        RECT 346.200 367.600 346.800 368.000 ;
        RECT 349.800 367.600 355.600 368.200 ;
        RECT 356.200 367.600 358.800 368.400 ;
        RECT 343.600 366.800 345.600 367.400 ;
        RECT 346.200 366.800 350.400 367.600 ;
        RECT 345.000 366.200 345.600 366.800 ;
        RECT 345.000 365.600 346.000 366.200 ;
        RECT 345.200 362.200 346.000 365.600 ;
        RECT 348.400 362.200 349.200 366.800 ;
        RECT 351.600 362.200 352.400 365.000 ;
        RECT 353.200 362.200 354.000 365.000 ;
        RECT 354.800 362.200 355.600 367.000 ;
        RECT 358.000 362.200 358.800 367.000 ;
        RECT 361.200 362.200 362.000 368.400 ;
        RECT 369.200 367.600 371.800 368.400 ;
        RECT 364.400 366.800 368.600 367.600 ;
        RECT 362.800 362.200 363.600 365.000 ;
        RECT 364.400 362.200 365.200 365.000 ;
        RECT 366.000 362.200 366.800 365.000 ;
        RECT 369.200 362.200 370.000 367.600 ;
        RECT 374.400 367.400 375.000 369.000 ;
        RECT 372.400 366.800 375.000 367.400 ;
        RECT 375.600 370.000 376.600 370.800 ;
        RECT 380.200 375.200 381.200 376.000 ;
        RECT 380.200 370.800 381.000 375.200 ;
        RECT 382.000 374.600 382.800 379.800 ;
        RECT 388.400 376.600 389.200 379.800 ;
        RECT 390.000 377.000 390.800 379.800 ;
        RECT 391.600 377.000 392.400 379.800 ;
        RECT 393.200 377.000 394.000 379.800 ;
        RECT 394.800 377.000 395.600 379.800 ;
        RECT 398.000 377.000 398.800 379.800 ;
        RECT 401.200 377.000 402.000 379.800 ;
        RECT 402.800 377.000 403.600 379.800 ;
        RECT 404.400 377.000 405.200 379.800 ;
        RECT 386.800 375.800 389.200 376.600 ;
        RECT 406.000 376.600 406.800 379.800 ;
        RECT 386.800 375.200 387.600 375.800 ;
        RECT 381.600 374.000 382.800 374.600 ;
        RECT 385.800 374.600 387.600 375.200 ;
        RECT 391.600 375.600 392.600 376.400 ;
        RECT 395.600 375.600 397.200 376.400 ;
        RECT 398.000 375.800 402.600 376.400 ;
        RECT 406.000 375.800 408.600 376.600 ;
        RECT 398.000 375.600 398.800 375.800 ;
        RECT 381.600 372.000 382.200 374.000 ;
        RECT 385.800 373.400 386.600 374.600 ;
        RECT 382.800 372.600 386.600 373.400 ;
        RECT 391.600 372.800 392.400 375.600 ;
        RECT 398.000 374.800 398.800 375.000 ;
        RECT 394.400 374.200 398.800 374.800 ;
        RECT 394.400 374.000 395.200 374.200 ;
        RECT 399.600 373.600 400.400 375.200 ;
        RECT 401.800 373.400 402.600 375.800 ;
        RECT 407.800 375.200 408.600 375.800 ;
        RECT 407.800 374.400 410.800 375.200 ;
        RECT 412.400 373.800 413.200 379.800 ;
        RECT 414.000 375.200 414.800 379.800 ;
        RECT 417.200 376.400 418.000 379.800 ;
        RECT 421.000 376.400 421.800 379.800 ;
        RECT 417.200 375.600 418.200 376.400 ;
        RECT 421.000 375.800 422.800 376.400 ;
        RECT 425.200 375.800 426.000 379.800 ;
        RECT 426.800 376.000 427.600 379.800 ;
        RECT 430.000 376.000 430.800 379.800 ;
        RECT 426.800 375.800 430.800 376.000 ;
        RECT 431.600 376.000 432.400 379.800 ;
        RECT 434.800 376.000 435.600 379.800 ;
        RECT 431.600 375.800 435.600 376.000 ;
        RECT 436.400 375.800 437.200 379.800 ;
        RECT 440.600 376.400 441.400 379.800 ;
        RECT 439.600 375.800 441.400 376.400 ;
        RECT 449.200 376.000 450.000 379.800 ;
        RECT 414.000 374.600 416.600 375.200 ;
        RECT 394.800 372.600 398.000 373.400 ;
        RECT 401.800 372.600 403.800 373.400 ;
        RECT 404.400 373.000 413.200 373.800 ;
        RECT 388.400 372.000 389.200 372.600 ;
        RECT 406.000 372.000 406.800 372.400 ;
        RECT 407.600 372.000 408.400 372.400 ;
        RECT 411.000 372.000 411.800 372.200 ;
        RECT 381.600 371.400 382.400 372.000 ;
        RECT 388.400 371.400 411.800 372.000 ;
        RECT 380.200 370.000 381.200 370.800 ;
        RECT 372.400 362.200 373.200 366.800 ;
        RECT 375.600 362.200 376.400 370.000 ;
        RECT 380.400 362.200 381.200 370.000 ;
        RECT 381.800 369.600 382.400 371.400 ;
        RECT 381.800 369.000 390.800 369.600 ;
        RECT 381.800 367.400 382.400 369.000 ;
        RECT 390.000 368.800 390.800 369.000 ;
        RECT 393.200 369.000 401.800 369.600 ;
        RECT 393.200 368.800 394.000 369.000 ;
        RECT 385.000 367.600 387.600 368.400 ;
        RECT 381.800 366.800 384.400 367.400 ;
        RECT 383.600 362.200 384.400 366.800 ;
        RECT 386.800 362.200 387.600 367.600 ;
        RECT 388.200 366.800 392.400 367.600 ;
        RECT 390.000 362.200 390.800 365.000 ;
        RECT 391.600 362.200 392.400 365.000 ;
        RECT 393.200 362.200 394.000 365.000 ;
        RECT 394.800 362.200 395.600 368.400 ;
        RECT 398.000 367.600 400.600 368.400 ;
        RECT 401.200 368.200 401.800 369.000 ;
        RECT 402.800 369.400 403.600 369.600 ;
        RECT 402.800 369.000 408.200 369.400 ;
        RECT 402.800 368.800 409.000 369.000 ;
        RECT 407.600 368.200 409.000 368.800 ;
        RECT 401.200 367.600 407.000 368.200 ;
        RECT 410.000 368.000 411.600 368.800 ;
        RECT 410.000 367.600 410.600 368.000 ;
        RECT 398.000 362.200 398.800 367.000 ;
        RECT 401.200 362.200 402.000 367.000 ;
        RECT 406.400 366.800 410.600 367.600 ;
        RECT 412.400 367.400 413.200 373.000 ;
        RECT 416.000 373.000 416.600 374.600 ;
        RECT 417.600 374.400 418.200 375.600 ;
        RECT 417.200 373.600 418.200 374.400 ;
        RECT 418.800 374.300 419.600 374.400 ;
        RECT 422.000 374.300 422.800 375.800 ;
        RECT 418.800 373.700 422.800 374.300 ;
        RECT 418.800 373.600 419.600 373.700 ;
        RECT 416.000 372.200 417.000 373.000 ;
        RECT 416.000 370.200 416.600 372.200 ;
        RECT 417.600 370.200 418.200 373.600 ;
        RECT 411.200 366.800 413.200 367.400 ;
        RECT 414.000 369.600 416.600 370.200 ;
        RECT 402.800 362.200 403.600 365.000 ;
        RECT 404.400 362.200 405.200 365.000 ;
        RECT 407.600 362.200 408.400 366.800 ;
        RECT 411.200 366.200 411.800 366.800 ;
        RECT 410.800 365.600 411.800 366.200 ;
        RECT 410.800 362.200 411.600 365.600 ;
        RECT 414.000 362.200 414.800 369.600 ;
        RECT 417.200 369.200 418.200 370.200 ;
        RECT 417.200 362.200 418.000 369.200 ;
        RECT 420.400 368.800 421.200 370.400 ;
        RECT 422.000 362.200 422.800 373.700 ;
        RECT 423.600 374.300 424.400 375.200 ;
        RECT 425.400 374.400 426.000 375.800 ;
        RECT 427.000 375.400 430.600 375.800 ;
        RECT 431.800 375.400 435.400 375.800 ;
        RECT 429.200 374.400 430.000 374.800 ;
        RECT 432.400 374.400 433.200 374.800 ;
        RECT 436.400 374.400 437.000 375.800 ;
        RECT 425.200 374.300 427.800 374.400 ;
        RECT 423.600 373.700 427.800 374.300 ;
        RECT 429.200 374.300 430.800 374.400 ;
        RECT 431.600 374.300 433.200 374.400 ;
        RECT 429.200 373.800 433.200 374.300 ;
        RECT 434.600 374.300 437.200 374.400 ;
        RECT 438.000 374.300 438.800 375.200 ;
        RECT 423.600 373.600 424.400 373.700 ;
        RECT 425.200 373.600 427.800 373.700 ;
        RECT 430.000 373.700 432.400 373.800 ;
        RECT 430.000 373.600 430.800 373.700 ;
        RECT 431.600 373.600 432.400 373.700 ;
        RECT 434.600 373.700 438.800 374.300 ;
        RECT 434.600 373.600 437.200 373.700 ;
        RECT 438.000 373.600 438.800 373.700 ;
        RECT 439.600 374.300 440.400 375.800 ;
        RECT 449.000 375.200 450.000 376.000 ;
        RECT 447.600 374.300 448.400 374.400 ;
        RECT 439.600 373.700 448.400 374.300 ;
        RECT 423.600 370.300 424.400 370.400 ;
        RECT 425.200 370.300 426.000 370.400 ;
        RECT 423.600 370.200 426.000 370.300 ;
        RECT 427.200 370.200 427.800 373.600 ;
        RECT 428.400 372.300 429.200 373.200 ;
        RECT 433.200 372.300 434.000 373.200 ;
        RECT 428.400 371.700 434.000 372.300 ;
        RECT 428.400 371.600 429.200 371.700 ;
        RECT 433.200 371.600 434.000 371.700 ;
        RECT 434.600 370.200 435.200 373.600 ;
        RECT 436.400 370.300 437.200 370.400 ;
        RECT 438.000 370.300 438.800 370.400 ;
        RECT 436.400 370.200 438.800 370.300 ;
        RECT 423.600 369.700 426.600 370.200 ;
        RECT 423.600 369.600 424.400 369.700 ;
        RECT 425.200 369.600 426.600 369.700 ;
        RECT 427.200 369.600 428.200 370.200 ;
        RECT 426.000 368.400 426.600 369.600 ;
        RECT 426.000 367.600 426.800 368.400 ;
        RECT 427.400 362.200 428.200 369.600 ;
        RECT 434.200 369.600 435.200 370.200 ;
        RECT 435.800 369.700 438.800 370.200 ;
        RECT 435.800 369.600 437.200 369.700 ;
        RECT 438.000 369.600 438.800 369.700 ;
        RECT 434.200 362.200 435.000 369.600 ;
        RECT 435.800 368.400 436.400 369.600 ;
        RECT 435.600 367.600 436.400 368.400 ;
        RECT 439.600 362.200 440.400 373.700 ;
        RECT 447.600 373.600 448.400 373.700 ;
        RECT 449.000 370.800 449.800 375.200 ;
        RECT 450.800 374.600 451.600 379.800 ;
        RECT 457.200 376.600 458.000 379.800 ;
        RECT 458.800 377.000 459.600 379.800 ;
        RECT 460.400 377.000 461.200 379.800 ;
        RECT 462.000 377.000 462.800 379.800 ;
        RECT 463.600 377.000 464.400 379.800 ;
        RECT 466.800 377.000 467.600 379.800 ;
        RECT 470.000 377.000 470.800 379.800 ;
        RECT 471.600 377.000 472.400 379.800 ;
        RECT 473.200 377.000 474.000 379.800 ;
        RECT 455.600 375.800 458.000 376.600 ;
        RECT 474.800 376.600 475.600 379.800 ;
        RECT 455.600 375.200 456.400 375.800 ;
        RECT 450.400 374.000 451.600 374.600 ;
        RECT 454.600 374.600 456.400 375.200 ;
        RECT 460.400 375.600 461.400 376.400 ;
        RECT 464.400 375.600 466.000 376.400 ;
        RECT 466.800 375.800 471.400 376.400 ;
        RECT 474.800 375.800 477.400 376.600 ;
        RECT 466.800 375.600 467.600 375.800 ;
        RECT 450.400 372.000 451.000 374.000 ;
        RECT 454.600 373.400 455.400 374.600 ;
        RECT 451.600 372.600 455.400 373.400 ;
        RECT 460.400 372.800 461.200 375.600 ;
        RECT 466.800 374.800 467.600 375.000 ;
        RECT 463.200 374.200 467.600 374.800 ;
        RECT 463.200 374.000 464.000 374.200 ;
        RECT 468.400 373.600 469.200 375.200 ;
        RECT 470.600 373.400 471.400 375.800 ;
        RECT 476.600 375.200 477.400 375.800 ;
        RECT 476.600 374.400 479.600 375.200 ;
        RECT 481.200 373.800 482.000 379.800 ;
        RECT 463.600 372.600 466.800 373.400 ;
        RECT 470.600 372.600 472.600 373.400 ;
        RECT 473.200 373.000 482.000 373.800 ;
        RECT 457.200 372.000 458.000 372.600 ;
        RECT 474.800 372.000 475.600 372.400 ;
        RECT 478.000 372.000 478.800 372.400 ;
        RECT 479.800 372.000 480.600 372.200 ;
        RECT 450.400 371.400 451.200 372.000 ;
        RECT 457.200 371.400 480.600 372.000 ;
        RECT 441.200 370.300 442.000 370.400 ;
        RECT 444.400 370.300 445.200 370.400 ;
        RECT 441.200 369.700 445.200 370.300 ;
        RECT 449.000 370.000 450.000 370.800 ;
        RECT 441.200 368.800 442.000 369.700 ;
        RECT 444.400 369.600 445.200 369.700 ;
        RECT 449.200 362.200 450.000 370.000 ;
        RECT 450.600 369.600 451.200 371.400 ;
        RECT 450.600 369.000 459.600 369.600 ;
        RECT 450.600 367.400 451.200 369.000 ;
        RECT 458.800 368.800 459.600 369.000 ;
        RECT 462.000 369.000 470.600 369.600 ;
        RECT 462.000 368.800 462.800 369.000 ;
        RECT 453.800 367.600 456.400 368.400 ;
        RECT 450.600 366.800 453.200 367.400 ;
        RECT 452.400 362.200 453.200 366.800 ;
        RECT 455.600 362.200 456.400 367.600 ;
        RECT 457.000 366.800 461.200 367.600 ;
        RECT 458.800 362.200 459.600 365.000 ;
        RECT 460.400 362.200 461.200 365.000 ;
        RECT 462.000 362.200 462.800 365.000 ;
        RECT 463.600 362.200 464.400 368.400 ;
        RECT 466.800 367.600 469.400 368.400 ;
        RECT 470.000 368.200 470.600 369.000 ;
        RECT 471.600 369.400 472.400 369.600 ;
        RECT 471.600 369.000 477.000 369.400 ;
        RECT 471.600 368.800 477.800 369.000 ;
        RECT 476.400 368.200 477.800 368.800 ;
        RECT 470.000 367.600 475.800 368.200 ;
        RECT 478.800 368.000 480.400 368.800 ;
        RECT 478.800 367.600 479.400 368.000 ;
        RECT 466.800 362.200 467.600 367.000 ;
        RECT 470.000 362.200 470.800 367.000 ;
        RECT 475.200 366.800 479.400 367.600 ;
        RECT 481.200 367.400 482.000 373.000 ;
        RECT 480.000 366.800 482.000 367.400 ;
        RECT 471.600 362.200 472.400 365.000 ;
        RECT 473.200 362.200 474.000 365.000 ;
        RECT 476.400 362.200 477.200 366.800 ;
        RECT 480.000 366.200 480.600 366.800 ;
        RECT 479.600 365.600 480.600 366.200 ;
        RECT 479.600 362.200 480.400 365.600 ;
        RECT 482.800 362.200 483.600 379.800 ;
        RECT 484.400 375.600 485.200 377.200 ;
        RECT 487.600 375.200 488.400 379.800 ;
        RECT 490.800 375.200 491.600 379.800 ;
        RECT 494.000 375.200 494.800 379.800 ;
        RECT 497.200 375.200 498.000 379.800 ;
        RECT 502.000 376.400 502.800 379.800 ;
        RECT 486.000 374.400 488.400 375.200 ;
        RECT 489.400 374.400 491.600 375.200 ;
        RECT 492.600 374.400 494.800 375.200 ;
        RECT 496.200 374.400 498.000 375.200 ;
        RECT 501.800 375.800 502.800 376.400 ;
        RECT 501.800 374.400 502.400 375.800 ;
        RECT 505.200 375.200 506.000 379.800 ;
        RECT 508.400 376.400 509.200 379.800 ;
        RECT 503.400 374.600 506.000 375.200 ;
        RECT 508.200 375.800 509.200 376.400 ;
        RECT 486.000 371.600 486.800 374.400 ;
        RECT 489.400 373.800 490.200 374.400 ;
        RECT 492.600 373.800 493.400 374.400 ;
        RECT 496.200 373.800 497.000 374.400 ;
        RECT 498.800 373.800 499.600 374.400 ;
        RECT 487.600 373.000 490.200 373.800 ;
        RECT 491.000 373.000 493.400 373.800 ;
        RECT 494.400 373.000 497.000 373.800 ;
        RECT 497.800 373.000 499.600 373.800 ;
        RECT 500.400 374.300 501.200 374.400 ;
        RECT 501.800 374.300 502.800 374.400 ;
        RECT 500.400 373.700 502.800 374.300 ;
        RECT 500.400 373.600 501.200 373.700 ;
        RECT 501.800 373.600 502.800 373.700 ;
        RECT 489.400 371.600 490.200 373.000 ;
        RECT 492.600 371.600 493.400 373.000 ;
        RECT 496.200 371.600 497.000 373.000 ;
        RECT 486.000 370.800 488.400 371.600 ;
        RECT 489.400 370.800 491.600 371.600 ;
        RECT 492.600 370.800 494.800 371.600 ;
        RECT 496.200 370.800 498.000 371.600 ;
        RECT 487.600 362.200 488.400 370.800 ;
        RECT 490.800 362.200 491.600 370.800 ;
        RECT 494.000 362.200 494.800 370.800 ;
        RECT 497.200 362.200 498.000 370.800 ;
        RECT 501.800 370.200 502.400 373.600 ;
        RECT 503.400 373.000 504.000 374.600 ;
        RECT 508.200 374.400 508.800 375.800 ;
        RECT 511.600 375.200 512.400 379.800 ;
        RECT 514.800 376.400 515.600 379.800 ;
        RECT 509.800 374.600 512.400 375.200 ;
        RECT 514.600 375.800 515.600 376.400 ;
        RECT 508.200 373.600 509.200 374.400 ;
        RECT 503.000 372.200 504.000 373.000 ;
        RECT 503.400 370.200 504.000 372.200 ;
        RECT 505.000 372.400 505.800 373.200 ;
        RECT 505.000 371.600 506.000 372.400 ;
        RECT 508.200 370.200 508.800 373.600 ;
        RECT 509.800 373.000 510.400 374.600 ;
        RECT 514.600 374.400 515.200 375.800 ;
        RECT 518.000 375.200 518.800 379.800 ;
        RECT 521.200 376.000 522.000 379.800 ;
        RECT 516.200 374.600 518.800 375.200 ;
        RECT 521.000 375.200 522.000 376.000 ;
        RECT 514.600 373.600 515.600 374.400 ;
        RECT 509.400 372.200 510.400 373.000 ;
        RECT 509.800 370.200 510.400 372.200 ;
        RECT 511.400 372.400 512.200 373.200 ;
        RECT 511.400 371.600 512.400 372.400 ;
        RECT 514.600 370.200 515.200 373.600 ;
        RECT 516.200 373.000 516.800 374.600 ;
        RECT 515.800 372.200 516.800 373.000 ;
        RECT 516.200 370.200 516.800 372.200 ;
        RECT 517.800 372.400 518.600 373.200 ;
        RECT 517.800 372.300 518.800 372.400 ;
        RECT 521.000 372.300 521.800 375.200 ;
        RECT 522.800 374.600 523.600 379.800 ;
        RECT 529.200 376.600 530.000 379.800 ;
        RECT 530.800 377.000 531.600 379.800 ;
        RECT 532.400 377.000 533.200 379.800 ;
        RECT 534.000 377.000 534.800 379.800 ;
        RECT 535.600 377.000 536.400 379.800 ;
        RECT 538.800 377.000 539.600 379.800 ;
        RECT 542.000 377.000 542.800 379.800 ;
        RECT 543.600 377.000 544.400 379.800 ;
        RECT 545.200 377.000 546.000 379.800 ;
        RECT 527.600 375.800 530.000 376.600 ;
        RECT 546.800 376.600 547.600 379.800 ;
        RECT 527.600 375.200 528.400 375.800 ;
        RECT 517.800 371.700 521.800 372.300 ;
        RECT 517.800 371.600 518.800 371.700 ;
        RECT 521.000 370.800 521.800 371.700 ;
        RECT 522.400 374.000 523.600 374.600 ;
        RECT 526.600 374.600 528.400 375.200 ;
        RECT 532.400 375.600 533.400 376.400 ;
        RECT 536.400 375.600 538.000 376.400 ;
        RECT 538.800 375.800 543.400 376.400 ;
        RECT 546.800 375.800 549.400 376.600 ;
        RECT 538.800 375.600 539.600 375.800 ;
        RECT 522.400 372.000 523.000 374.000 ;
        RECT 526.600 373.400 527.400 374.600 ;
        RECT 523.600 372.600 527.400 373.400 ;
        RECT 532.400 372.800 533.200 375.600 ;
        RECT 538.800 374.800 539.600 375.000 ;
        RECT 535.200 374.200 539.600 374.800 ;
        RECT 535.200 374.000 536.000 374.200 ;
        RECT 540.400 373.600 541.200 375.200 ;
        RECT 542.600 373.400 543.400 375.800 ;
        RECT 548.600 375.200 549.400 375.800 ;
        RECT 548.600 374.400 551.600 375.200 ;
        RECT 553.200 373.800 554.000 379.800 ;
        RECT 554.800 375.200 555.600 379.800 ;
        RECT 558.000 376.400 558.800 379.800 ;
        RECT 561.800 376.400 562.600 379.800 ;
        RECT 558.000 375.800 559.000 376.400 ;
        RECT 561.800 375.800 563.600 376.400 ;
        RECT 566.000 376.000 566.800 379.800 ;
        RECT 569.200 376.000 570.000 379.800 ;
        RECT 566.000 375.800 570.000 376.000 ;
        RECT 570.800 375.800 571.600 379.800 ;
        RECT 574.000 376.000 574.800 379.800 ;
        RECT 554.800 374.600 557.400 375.200 ;
        RECT 535.600 372.600 538.800 373.400 ;
        RECT 542.600 372.600 544.600 373.400 ;
        RECT 545.200 373.000 554.000 373.800 ;
        RECT 522.400 371.400 523.200 372.000 ;
        RECT 501.800 369.200 502.800 370.200 ;
        RECT 503.400 369.600 506.000 370.200 ;
        RECT 502.000 362.200 502.800 369.200 ;
        RECT 505.200 362.200 506.000 369.600 ;
        RECT 508.200 369.200 509.200 370.200 ;
        RECT 509.800 369.600 512.400 370.200 ;
        RECT 508.400 362.200 509.200 369.200 ;
        RECT 511.600 362.200 512.400 369.600 ;
        RECT 514.600 369.200 515.600 370.200 ;
        RECT 516.200 369.600 518.800 370.200 ;
        RECT 521.000 370.000 522.000 370.800 ;
        RECT 514.800 362.200 515.600 369.200 ;
        RECT 518.000 362.200 518.800 369.600 ;
        RECT 521.200 362.200 522.000 370.000 ;
        RECT 522.600 369.600 523.200 371.400 ;
        RECT 523.800 370.800 524.600 371.000 ;
        RECT 523.800 370.200 550.800 370.800 ;
        RECT 546.600 370.000 547.600 370.200 ;
        RECT 550.000 369.600 550.800 370.200 ;
        RECT 522.600 369.000 531.600 369.600 ;
        RECT 522.600 367.400 523.200 369.000 ;
        RECT 530.800 368.800 531.600 369.000 ;
        RECT 534.000 369.000 542.600 369.600 ;
        RECT 534.000 368.800 534.800 369.000 ;
        RECT 525.800 367.600 528.400 368.400 ;
        RECT 522.600 366.800 525.200 367.400 ;
        RECT 524.400 362.200 525.200 366.800 ;
        RECT 527.600 362.200 528.400 367.600 ;
        RECT 529.000 366.800 533.200 367.600 ;
        RECT 530.800 362.200 531.600 365.000 ;
        RECT 532.400 362.200 533.200 365.000 ;
        RECT 534.000 362.200 534.800 365.000 ;
        RECT 535.600 362.200 536.400 368.400 ;
        RECT 538.800 367.600 541.400 368.400 ;
        RECT 542.000 368.200 542.600 369.000 ;
        RECT 543.600 369.400 544.400 369.600 ;
        RECT 543.600 369.000 549.000 369.400 ;
        RECT 543.600 368.800 549.800 369.000 ;
        RECT 548.400 368.200 549.800 368.800 ;
        RECT 542.000 367.600 547.800 368.200 ;
        RECT 550.800 368.000 552.400 368.800 ;
        RECT 550.800 367.600 551.400 368.000 ;
        RECT 538.800 362.200 539.600 367.000 ;
        RECT 542.000 362.200 542.800 367.000 ;
        RECT 547.200 366.800 551.400 367.600 ;
        RECT 553.200 367.400 554.000 373.000 ;
        RECT 555.000 372.400 555.800 373.200 ;
        RECT 554.800 371.600 555.800 372.400 ;
        RECT 556.800 373.000 557.400 374.600 ;
        RECT 558.400 374.400 559.000 375.800 ;
        RECT 558.000 373.600 559.000 374.400 ;
        RECT 556.800 372.200 557.800 373.000 ;
        RECT 556.800 370.200 557.400 372.200 ;
        RECT 558.400 370.200 559.000 373.600 ;
        RECT 552.000 366.800 554.000 367.400 ;
        RECT 554.800 369.600 557.400 370.200 ;
        RECT 543.600 362.200 544.400 365.000 ;
        RECT 545.200 362.200 546.000 365.000 ;
        RECT 548.400 362.200 549.200 366.800 ;
        RECT 552.000 366.200 552.600 366.800 ;
        RECT 551.600 365.600 552.600 366.200 ;
        RECT 551.600 362.200 552.400 365.600 ;
        RECT 554.800 362.200 555.600 369.600 ;
        RECT 558.000 369.200 559.000 370.200 ;
        RECT 558.000 362.200 558.800 369.200 ;
        RECT 561.200 368.800 562.000 370.400 ;
        RECT 562.800 362.200 563.600 375.800 ;
        RECT 566.200 375.400 569.800 375.800 ;
        RECT 564.400 373.600 565.200 375.200 ;
        RECT 566.800 374.400 567.600 374.800 ;
        RECT 570.800 374.400 571.400 375.800 ;
        RECT 573.800 375.200 574.800 376.000 ;
        RECT 566.000 373.800 567.600 374.400 ;
        RECT 566.000 373.600 566.800 373.800 ;
        RECT 569.000 373.600 571.600 374.400 ;
        RECT 567.600 371.600 568.400 373.200 ;
        RECT 569.000 370.200 569.600 373.600 ;
        RECT 573.800 370.800 574.600 375.200 ;
        RECT 575.600 374.600 576.400 379.800 ;
        RECT 582.000 376.600 582.800 379.800 ;
        RECT 583.600 377.000 584.400 379.800 ;
        RECT 585.200 377.000 586.000 379.800 ;
        RECT 586.800 377.000 587.600 379.800 ;
        RECT 588.400 377.000 589.200 379.800 ;
        RECT 591.600 377.000 592.400 379.800 ;
        RECT 594.800 377.000 595.600 379.800 ;
        RECT 596.400 377.000 597.200 379.800 ;
        RECT 598.000 377.000 598.800 379.800 ;
        RECT 580.400 375.800 582.800 376.600 ;
        RECT 599.600 376.600 600.400 379.800 ;
        RECT 580.400 375.200 581.200 375.800 ;
        RECT 575.200 374.000 576.400 374.600 ;
        RECT 579.400 374.600 581.200 375.200 ;
        RECT 585.200 375.600 586.200 376.400 ;
        RECT 589.200 375.600 590.800 376.400 ;
        RECT 591.600 375.800 596.200 376.400 ;
        RECT 599.600 375.800 602.200 376.600 ;
        RECT 591.600 375.600 592.400 375.800 ;
        RECT 575.200 372.000 575.800 374.000 ;
        RECT 579.400 373.400 580.200 374.600 ;
        RECT 576.400 372.600 580.200 373.400 ;
        RECT 585.200 372.800 586.000 375.600 ;
        RECT 591.600 374.800 592.400 375.000 ;
        RECT 588.000 374.200 592.400 374.800 ;
        RECT 588.000 374.000 588.800 374.200 ;
        RECT 593.200 373.600 594.000 375.200 ;
        RECT 595.400 373.400 596.200 375.800 ;
        RECT 601.400 375.200 602.200 375.800 ;
        RECT 601.400 374.400 604.400 375.200 ;
        RECT 606.000 373.800 606.800 379.800 ;
        RECT 607.600 375.200 608.400 379.800 ;
        RECT 607.600 374.600 609.800 375.200 ;
        RECT 588.400 372.600 591.600 373.400 ;
        RECT 595.400 372.600 597.400 373.400 ;
        RECT 598.000 373.000 606.800 373.800 ;
        RECT 582.000 372.000 582.800 372.600 ;
        RECT 599.600 372.000 600.400 372.400 ;
        RECT 604.600 372.000 605.400 372.200 ;
        RECT 575.200 371.400 576.000 372.000 ;
        RECT 582.000 371.400 605.400 372.000 ;
        RECT 570.800 370.300 571.600 370.400 ;
        RECT 573.800 370.300 574.800 370.800 ;
        RECT 570.800 370.200 574.800 370.300 ;
        RECT 568.600 369.600 569.600 370.200 ;
        RECT 570.200 369.700 574.800 370.200 ;
        RECT 570.200 369.600 571.600 369.700 ;
        RECT 568.600 362.200 569.400 369.600 ;
        RECT 570.200 368.400 570.800 369.600 ;
        RECT 570.000 367.600 571.600 368.400 ;
        RECT 574.000 362.200 574.800 369.700 ;
        RECT 575.400 369.600 576.000 371.400 ;
        RECT 575.400 369.000 584.400 369.600 ;
        RECT 575.400 367.400 576.000 369.000 ;
        RECT 583.600 368.800 584.400 369.000 ;
        RECT 586.800 369.000 595.400 369.600 ;
        RECT 586.800 368.800 587.600 369.000 ;
        RECT 578.600 367.600 581.200 368.400 ;
        RECT 575.400 366.800 578.000 367.400 ;
        RECT 577.200 362.200 578.000 366.800 ;
        RECT 580.400 362.200 581.200 367.600 ;
        RECT 581.800 366.800 586.000 367.600 ;
        RECT 583.600 362.200 584.400 365.000 ;
        RECT 585.200 362.200 586.000 365.000 ;
        RECT 586.800 362.200 587.600 365.000 ;
        RECT 588.400 362.200 589.200 368.400 ;
        RECT 591.600 367.600 594.200 368.400 ;
        RECT 594.800 368.200 595.400 369.000 ;
        RECT 596.400 369.400 597.200 369.600 ;
        RECT 596.400 369.000 601.800 369.400 ;
        RECT 596.400 368.800 602.600 369.000 ;
        RECT 601.200 368.200 602.600 368.800 ;
        RECT 594.800 367.600 600.600 368.200 ;
        RECT 603.600 368.000 605.200 368.800 ;
        RECT 603.600 367.600 604.200 368.000 ;
        RECT 591.600 362.200 592.400 367.000 ;
        RECT 594.800 362.200 595.600 367.000 ;
        RECT 600.000 366.800 604.200 367.600 ;
        RECT 606.000 367.400 606.800 373.000 ;
        RECT 607.600 371.600 608.400 373.200 ;
        RECT 609.200 371.600 609.800 374.600 ;
        RECT 609.200 370.800 610.400 371.600 ;
        RECT 609.200 370.200 609.800 370.800 ;
        RECT 604.800 366.800 606.800 367.400 ;
        RECT 607.600 369.600 609.800 370.200 ;
        RECT 596.400 362.200 597.200 365.000 ;
        RECT 598.000 362.200 598.800 365.000 ;
        RECT 601.200 362.200 602.000 366.800 ;
        RECT 604.800 366.200 605.400 366.800 ;
        RECT 604.400 365.600 605.400 366.200 ;
        RECT 604.400 362.200 605.200 365.600 ;
        RECT 607.600 362.200 608.400 369.600 ;
        RECT 2.800 348.300 3.600 359.800 ;
        RECT 7.000 352.400 7.800 359.800 ;
        RECT 12.400 356.400 13.200 359.800 ;
        RECT 12.200 355.800 13.200 356.400 ;
        RECT 12.200 355.200 12.800 355.800 ;
        RECT 15.600 355.200 16.400 359.800 ;
        RECT 18.800 357.000 19.600 359.800 ;
        RECT 20.400 357.000 21.200 359.800 ;
        RECT 10.800 354.600 12.800 355.200 ;
        RECT 8.400 353.600 9.200 354.400 ;
        RECT 8.600 352.400 9.200 353.600 ;
        RECT 7.000 351.800 8.000 352.400 ;
        RECT 8.600 351.800 10.000 352.400 ;
        RECT 6.000 348.800 6.800 350.400 ;
        RECT 7.400 348.400 8.000 351.800 ;
        RECT 9.200 351.600 10.000 351.800 ;
        RECT 10.800 349.000 11.600 354.600 ;
        RECT 13.400 354.400 17.600 355.200 ;
        RECT 22.000 355.000 22.800 359.800 ;
        RECT 25.200 355.000 26.000 359.800 ;
        RECT 13.400 354.000 14.000 354.400 ;
        RECT 12.400 353.200 14.000 354.000 ;
        RECT 17.000 353.800 22.800 354.400 ;
        RECT 15.000 353.200 16.400 353.800 ;
        RECT 15.000 353.000 21.200 353.200 ;
        RECT 15.800 352.600 21.200 353.000 ;
        RECT 20.400 352.400 21.200 352.600 ;
        RECT 22.200 353.000 22.800 353.800 ;
        RECT 23.400 353.600 26.000 354.400 ;
        RECT 28.400 353.600 29.200 359.800 ;
        RECT 30.000 357.000 30.800 359.800 ;
        RECT 31.600 357.000 32.400 359.800 ;
        RECT 33.200 357.000 34.000 359.800 ;
        RECT 31.600 354.400 35.800 355.200 ;
        RECT 36.400 354.400 37.200 359.800 ;
        RECT 39.600 355.200 40.400 359.800 ;
        RECT 39.600 354.600 42.200 355.200 ;
        RECT 36.400 353.600 39.000 354.400 ;
        RECT 30.000 353.000 30.800 353.200 ;
        RECT 22.200 352.400 30.800 353.000 ;
        RECT 33.200 353.000 34.000 353.200 ;
        RECT 41.600 353.000 42.200 354.600 ;
        RECT 33.200 352.400 42.200 353.000 ;
        RECT 41.600 350.600 42.200 352.400 ;
        RECT 42.800 352.000 43.600 359.800 ;
        RECT 42.800 351.200 43.800 352.000 ;
        RECT 12.200 350.000 35.600 350.600 ;
        RECT 41.600 350.000 42.400 350.600 ;
        RECT 12.200 349.800 13.200 350.000 ;
        RECT 12.400 349.600 13.200 349.800 ;
        RECT 17.200 349.600 18.000 350.000 ;
        RECT 23.600 349.600 24.400 350.000 ;
        RECT 34.800 349.400 35.600 350.000 ;
        RECT 4.400 348.300 5.200 348.400 ;
        RECT 2.800 348.200 5.200 348.300 ;
        RECT 2.800 347.700 6.000 348.200 ;
        RECT 2.800 342.200 3.600 347.700 ;
        RECT 4.400 347.600 6.000 347.700 ;
        RECT 7.400 347.600 10.000 348.400 ;
        RECT 10.800 348.200 19.600 349.000 ;
        RECT 20.200 348.600 22.200 349.400 ;
        RECT 26.000 348.600 29.200 349.400 ;
        RECT 5.200 347.200 6.000 347.600 ;
        RECT 4.600 346.200 8.200 346.600 ;
        RECT 9.200 346.200 9.800 347.600 ;
        RECT 4.400 346.000 8.400 346.200 ;
        RECT 4.400 342.200 5.200 346.000 ;
        RECT 7.600 342.200 8.400 346.000 ;
        RECT 9.200 342.200 10.000 346.200 ;
        RECT 10.800 342.200 11.600 348.200 ;
        RECT 13.200 346.800 16.200 347.600 ;
        RECT 15.400 346.200 16.200 346.800 ;
        RECT 21.400 346.200 22.200 348.600 ;
        RECT 23.600 346.800 24.400 348.400 ;
        RECT 28.800 347.800 29.600 348.000 ;
        RECT 25.200 347.200 29.600 347.800 ;
        RECT 25.200 347.000 26.000 347.200 ;
        RECT 31.600 346.400 32.400 349.200 ;
        RECT 37.400 348.600 41.200 349.400 ;
        RECT 37.400 347.400 38.200 348.600 ;
        RECT 41.800 348.000 42.400 350.000 ;
        RECT 25.200 346.200 26.000 346.400 ;
        RECT 15.400 345.400 18.000 346.200 ;
        RECT 21.400 345.600 26.000 346.200 ;
        RECT 26.800 345.600 28.400 346.400 ;
        RECT 31.400 345.600 32.400 346.400 ;
        RECT 36.400 346.800 38.200 347.400 ;
        RECT 41.200 347.400 42.400 348.000 ;
        RECT 36.400 346.200 37.200 346.800 ;
        RECT 17.200 342.200 18.000 345.400 ;
        RECT 34.800 345.400 37.200 346.200 ;
        RECT 18.800 342.200 19.600 345.000 ;
        RECT 20.400 342.200 21.200 345.000 ;
        RECT 22.000 342.200 22.800 345.000 ;
        RECT 25.200 342.200 26.000 345.000 ;
        RECT 28.400 342.200 29.200 345.000 ;
        RECT 30.000 342.200 30.800 345.000 ;
        RECT 31.600 342.200 32.400 345.000 ;
        RECT 33.200 342.200 34.000 345.000 ;
        RECT 34.800 342.200 35.600 345.400 ;
        RECT 41.200 342.200 42.000 347.400 ;
        RECT 43.000 346.800 43.800 351.200 ;
        RECT 42.800 346.000 43.800 346.800 ;
        RECT 44.400 346.300 45.200 346.400 ;
        RECT 46.000 346.300 46.800 346.400 ;
        RECT 42.800 342.200 43.600 346.000 ;
        RECT 44.400 345.700 46.800 346.300 ;
        RECT 44.400 345.600 45.200 345.700 ;
        RECT 46.000 344.800 46.800 345.700 ;
        RECT 47.600 342.200 48.400 359.800 ;
        RECT 49.200 342.200 50.000 359.800 ;
        RECT 54.000 354.300 54.800 359.800 ;
        RECT 55.600 354.300 56.400 354.400 ;
        RECT 54.000 353.700 56.400 354.300 ;
        RECT 50.800 352.300 51.600 352.400 ;
        RECT 52.400 352.300 53.200 353.200 ;
        RECT 50.800 351.700 53.200 352.300 ;
        RECT 50.800 351.600 51.600 351.700 ;
        RECT 52.400 351.600 53.200 351.700 ;
        RECT 50.800 344.800 51.600 346.400 ;
        RECT 54.000 346.200 54.800 353.700 ;
        RECT 55.600 353.600 56.400 353.700 ;
        RECT 55.600 346.800 56.400 348.400 ;
        RECT 53.000 345.600 54.800 346.200 ;
        RECT 53.000 342.200 53.800 345.600 ;
        RECT 57.200 342.200 58.000 359.800 ;
        RECT 60.400 351.400 61.200 359.800 ;
        RECT 64.800 356.400 65.600 359.800 ;
        RECT 63.600 355.800 65.600 356.400 ;
        RECT 69.200 355.800 70.000 359.800 ;
        RECT 73.400 355.800 74.600 359.800 ;
        RECT 63.600 355.000 64.400 355.800 ;
        RECT 69.200 355.200 69.800 355.800 ;
        RECT 67.000 354.600 70.600 355.200 ;
        RECT 73.200 355.000 74.000 355.800 ;
        RECT 67.000 354.400 67.800 354.600 ;
        RECT 69.800 354.400 70.600 354.600 ;
        RECT 63.600 353.000 64.400 353.200 ;
        RECT 68.200 353.000 69.000 353.200 ;
        RECT 63.600 352.400 69.000 353.000 ;
        RECT 69.600 353.000 71.800 353.600 ;
        RECT 69.600 351.800 70.200 353.000 ;
        RECT 71.000 352.800 71.800 353.000 ;
        RECT 73.400 353.200 74.800 354.000 ;
        RECT 73.400 352.200 74.000 353.200 ;
        RECT 65.400 351.400 70.200 351.800 ;
        RECT 60.400 351.200 70.200 351.400 ;
        RECT 71.600 351.600 74.000 352.200 ;
        RECT 60.400 351.000 66.200 351.200 ;
        RECT 60.400 350.800 66.000 351.000 ;
        RECT 66.800 350.300 67.600 350.400 ;
        RECT 68.400 350.300 69.200 350.400 ;
        RECT 66.800 350.200 69.200 350.300 ;
        RECT 62.600 349.700 69.200 350.200 ;
        RECT 62.600 349.600 67.600 349.700 ;
        RECT 68.400 349.600 69.200 349.700 ;
        RECT 62.600 349.400 63.400 349.600 ;
        RECT 64.200 348.400 65.000 348.600 ;
        RECT 71.600 348.400 72.200 351.600 ;
        RECT 78.000 351.200 78.800 359.800 ;
        RECT 74.600 350.600 78.800 351.200 ;
        RECT 74.600 350.400 75.400 350.600 ;
        RECT 76.200 349.800 77.000 350.000 ;
        RECT 73.200 349.200 77.000 349.800 ;
        RECT 73.200 349.000 74.000 349.200 ;
        RECT 61.200 347.800 72.200 348.400 ;
        RECT 61.200 347.600 62.800 347.800 ;
        RECT 58.800 344.800 59.600 346.400 ;
        RECT 60.400 342.200 61.200 347.000 ;
        RECT 65.400 345.600 66.000 347.800 ;
        RECT 68.400 347.600 69.200 347.800 ;
        RECT 71.000 347.600 71.800 347.800 ;
        RECT 78.000 347.200 78.800 350.600 ;
        RECT 75.000 346.600 78.800 347.200 ;
        RECT 75.000 346.400 75.800 346.600 ;
        RECT 63.600 344.200 64.400 345.000 ;
        RECT 65.200 344.800 66.000 345.600 ;
        RECT 67.000 345.400 67.800 345.600 ;
        RECT 67.000 344.800 69.800 345.400 ;
        RECT 69.200 344.200 69.800 344.800 ;
        RECT 73.200 344.200 74.000 345.000 ;
        RECT 63.600 343.600 65.600 344.200 ;
        RECT 64.800 342.200 65.600 343.600 ;
        RECT 69.200 342.200 70.000 344.200 ;
        RECT 73.200 343.600 74.600 344.200 ;
        RECT 73.400 342.200 74.600 343.600 ;
        RECT 78.000 342.200 78.800 346.600 ;
        RECT 79.600 342.200 80.400 359.800 ;
        RECT 81.200 352.300 82.000 352.400 ;
        RECT 82.800 352.300 83.600 353.200 ;
        RECT 81.200 351.700 83.600 352.300 ;
        RECT 81.200 351.600 82.000 351.700 ;
        RECT 82.800 351.600 83.600 351.700 ;
        RECT 84.400 352.300 85.200 359.800 ;
        RECT 88.400 353.600 89.200 354.400 ;
        RECT 88.400 352.400 89.000 353.600 ;
        RECT 89.800 352.400 90.600 359.800 ;
        RECT 96.200 354.400 97.000 359.800 ;
        RECT 94.800 353.600 95.600 354.400 ;
        RECT 96.200 353.600 98.000 354.400 ;
        RECT 94.800 352.400 95.400 353.600 ;
        RECT 96.200 352.400 97.000 353.600 ;
        RECT 87.600 352.300 89.000 352.400 ;
        RECT 84.400 351.800 89.000 352.300 ;
        RECT 84.400 351.700 88.400 351.800 ;
        RECT 81.200 344.800 82.000 346.400 ;
        RECT 84.400 346.200 85.200 351.700 ;
        RECT 87.600 351.600 88.400 351.700 ;
        RECT 89.600 351.600 91.600 352.400 ;
        RECT 94.000 351.800 95.400 352.400 ;
        RECT 96.000 351.800 97.000 352.400 ;
        RECT 94.000 351.600 94.800 351.800 ;
        RECT 89.600 348.400 90.200 351.600 ;
        RECT 90.800 348.800 91.600 350.400 ;
        RECT 92.400 350.300 93.200 350.400 ;
        RECT 96.000 350.300 96.600 351.800 ;
        RECT 92.400 349.700 96.600 350.300 ;
        RECT 92.400 349.600 93.200 349.700 ;
        RECT 96.000 348.400 96.600 349.700 ;
        RECT 97.200 350.300 98.000 350.400 ;
        RECT 100.400 350.300 101.200 359.800 ;
        RECT 103.600 355.000 104.400 359.000 ;
        RECT 103.600 351.600 104.200 355.000 ;
        RECT 107.800 352.800 108.600 359.800 ;
        RECT 107.800 352.200 109.400 352.800 ;
        RECT 103.600 351.000 107.400 351.600 ;
        RECT 97.200 349.700 101.200 350.300 ;
        RECT 97.200 348.800 98.000 349.700 ;
        RECT 86.000 346.800 86.800 348.400 ;
        RECT 87.600 347.600 90.200 348.400 ;
        RECT 92.400 348.200 93.200 348.400 ;
        RECT 91.600 347.600 93.200 348.200 ;
        RECT 94.000 347.600 96.600 348.400 ;
        RECT 98.800 348.200 99.600 348.400 ;
        RECT 98.000 347.600 99.600 348.200 ;
        RECT 87.800 346.200 88.400 347.600 ;
        RECT 91.600 347.200 92.400 347.600 ;
        RECT 89.400 346.200 93.000 346.600 ;
        RECT 94.200 346.200 94.800 347.600 ;
        RECT 98.000 347.200 98.800 347.600 ;
        RECT 95.800 346.200 99.400 346.600 ;
        RECT 83.400 345.600 85.200 346.200 ;
        RECT 83.400 342.200 84.200 345.600 ;
        RECT 87.600 342.200 88.400 346.200 ;
        RECT 89.200 346.000 93.200 346.200 ;
        RECT 89.200 342.200 90.000 346.000 ;
        RECT 92.400 342.200 93.200 346.000 ;
        RECT 94.000 342.200 94.800 346.200 ;
        RECT 95.600 346.000 99.600 346.200 ;
        RECT 95.600 342.200 96.400 346.000 ;
        RECT 98.800 342.200 99.600 346.000 ;
        RECT 100.400 342.200 101.200 349.700 ;
        RECT 103.600 348.800 104.400 350.400 ;
        RECT 105.200 348.800 106.000 350.400 ;
        RECT 106.800 349.000 107.400 351.000 ;
        RECT 106.800 348.200 108.200 349.000 ;
        RECT 108.800 348.400 109.400 352.200 ;
        RECT 115.800 352.400 116.600 359.800 ;
        RECT 117.200 353.600 118.000 354.400 ;
        RECT 117.400 352.400 118.000 353.600 ;
        RECT 120.400 353.600 121.200 354.400 ;
        RECT 120.400 352.400 121.000 353.600 ;
        RECT 121.800 352.400 122.600 359.800 ;
        RECT 126.800 353.600 127.600 354.400 ;
        RECT 126.800 352.400 127.400 353.600 ;
        RECT 128.200 352.400 129.000 359.800 ;
        RECT 115.800 351.800 116.800 352.400 ;
        RECT 117.400 351.800 118.800 352.400 ;
        RECT 110.000 350.300 110.800 351.200 ;
        RECT 113.200 350.300 114.000 350.400 ;
        RECT 110.000 349.700 114.000 350.300 ;
        RECT 110.000 349.600 110.800 349.700 ;
        RECT 113.200 349.600 114.000 349.700 ;
        RECT 114.800 348.800 115.600 350.400 ;
        RECT 116.200 348.400 116.800 351.800 ;
        RECT 118.000 351.600 118.800 351.800 ;
        RECT 119.600 351.800 121.000 352.400 ;
        RECT 121.600 351.800 122.600 352.400 ;
        RECT 126.000 351.800 127.400 352.400 ;
        RECT 128.000 351.800 129.000 352.400 ;
        RECT 132.400 355.000 133.200 359.000 ;
        RECT 119.600 351.600 120.400 351.800 ;
        RECT 118.100 350.300 118.700 351.600 ;
        RECT 121.600 350.300 122.200 351.800 ;
        RECT 126.000 351.600 126.800 351.800 ;
        RECT 118.100 349.700 122.200 350.300 ;
        RECT 121.600 348.400 122.200 349.700 ;
        RECT 122.800 348.800 123.600 350.400 ;
        RECT 128.000 348.400 128.600 351.800 ;
        RECT 132.400 351.600 133.000 355.000 ;
        RECT 136.600 352.800 137.400 359.800 ;
        RECT 136.600 352.200 138.200 352.800 ;
        RECT 132.400 351.000 136.200 351.600 ;
        RECT 129.200 348.800 130.000 350.400 ;
        RECT 132.400 348.800 133.200 350.400 ;
        RECT 134.000 348.800 134.800 350.400 ;
        RECT 135.600 349.000 136.200 351.000 ;
        RECT 108.800 348.300 110.800 348.400 ;
        RECT 111.600 348.300 112.400 348.400 ;
        RECT 106.800 347.800 107.800 348.200 ;
        RECT 103.600 347.200 107.800 347.800 ;
        RECT 108.800 347.700 112.400 348.300 ;
        RECT 108.800 347.600 110.800 347.700 ;
        RECT 111.600 347.600 112.400 347.700 ;
        RECT 113.200 348.200 114.000 348.400 ;
        RECT 113.200 347.600 114.800 348.200 ;
        RECT 116.200 347.600 118.800 348.400 ;
        RECT 119.600 347.600 122.200 348.400 ;
        RECT 124.400 348.200 125.200 348.400 ;
        RECT 123.600 347.600 125.200 348.200 ;
        RECT 126.000 347.600 128.600 348.400 ;
        RECT 130.800 348.200 131.600 348.400 ;
        RECT 130.000 347.600 131.600 348.200 ;
        RECT 135.600 348.200 137.000 349.000 ;
        RECT 137.600 348.400 138.200 352.200 ;
        RECT 143.600 351.200 144.400 359.800 ;
        RECT 146.800 351.200 147.600 359.800 ;
        RECT 150.000 351.200 150.800 359.800 ;
        RECT 153.200 351.200 154.000 359.800 ;
        RECT 138.800 350.300 139.600 351.200 ;
        RECT 143.600 350.400 145.400 351.200 ;
        RECT 146.800 350.400 149.000 351.200 ;
        RECT 150.000 350.400 152.200 351.200 ;
        RECT 153.200 350.400 155.600 351.200 ;
        RECT 142.000 350.300 142.800 350.400 ;
        RECT 138.800 349.700 142.800 350.300 ;
        RECT 138.800 349.600 139.600 349.700 ;
        RECT 142.000 349.600 142.800 349.700 ;
        RECT 144.600 349.000 145.400 350.400 ;
        RECT 148.200 349.000 149.000 350.400 ;
        RECT 151.400 349.000 152.200 350.400 ;
        RECT 135.600 347.800 136.600 348.200 ;
        RECT 102.000 344.800 102.800 346.400 ;
        RECT 103.600 345.000 104.200 347.200 ;
        RECT 108.800 347.000 109.400 347.600 ;
        RECT 114.000 347.200 114.800 347.600 ;
        RECT 108.600 346.600 109.400 347.000 ;
        RECT 107.800 346.000 109.400 346.600 ;
        RECT 113.400 346.200 117.000 346.600 ;
        RECT 118.000 346.200 118.600 347.600 ;
        RECT 119.800 346.200 120.400 347.600 ;
        RECT 123.600 347.200 124.400 347.600 ;
        RECT 121.400 346.200 125.000 346.600 ;
        RECT 126.200 346.200 126.800 347.600 ;
        RECT 130.000 347.200 130.800 347.600 ;
        RECT 132.400 347.200 136.600 347.800 ;
        RECT 137.600 347.600 139.600 348.400 ;
        RECT 142.000 348.200 143.800 349.000 ;
        RECT 144.600 348.200 147.200 349.000 ;
        RECT 148.200 348.200 150.600 349.000 ;
        RECT 151.400 348.200 154.000 349.000 ;
        RECT 142.000 347.600 142.800 348.200 ;
        RECT 144.600 347.600 145.400 348.200 ;
        RECT 148.200 347.600 149.000 348.200 ;
        RECT 151.400 347.600 152.200 348.200 ;
        RECT 154.800 347.600 155.600 350.400 ;
        RECT 127.800 346.200 131.400 346.600 ;
        RECT 113.200 346.000 117.200 346.200 ;
        RECT 103.600 343.000 104.400 345.000 ;
        RECT 107.800 343.000 108.600 346.000 ;
        RECT 113.200 342.200 114.000 346.000 ;
        RECT 116.400 342.200 117.200 346.000 ;
        RECT 118.000 342.200 118.800 346.200 ;
        RECT 119.600 342.200 120.400 346.200 ;
        RECT 121.200 346.000 125.200 346.200 ;
        RECT 121.200 342.200 122.000 346.000 ;
        RECT 124.400 342.200 125.200 346.000 ;
        RECT 126.000 342.200 126.800 346.200 ;
        RECT 127.600 346.000 131.600 346.200 ;
        RECT 127.600 342.200 128.400 346.000 ;
        RECT 130.800 342.200 131.600 346.000 ;
        RECT 132.400 345.000 133.000 347.200 ;
        RECT 137.600 347.000 138.200 347.600 ;
        RECT 137.400 346.600 138.200 347.000 ;
        RECT 136.600 346.000 138.200 346.600 ;
        RECT 143.600 346.800 145.400 347.600 ;
        RECT 146.800 346.800 149.000 347.600 ;
        RECT 150.000 346.800 152.200 347.600 ;
        RECT 153.200 346.800 155.600 347.600 ;
        RECT 162.800 350.300 163.600 359.800 ;
        RECT 168.200 352.800 169.000 359.800 ;
        RECT 172.400 355.000 173.200 359.000 ;
        RECT 167.400 352.200 169.000 352.800 ;
        RECT 166.000 350.300 166.800 351.200 ;
        RECT 162.800 349.700 166.800 350.300 ;
        RECT 132.400 343.000 133.200 345.000 ;
        RECT 136.600 344.400 137.400 346.000 ;
        RECT 135.600 343.600 137.400 344.400 ;
        RECT 136.600 343.000 137.400 343.600 ;
        RECT 143.600 342.200 144.400 346.800 ;
        RECT 146.800 342.200 147.600 346.800 ;
        RECT 150.000 342.200 150.800 346.800 ;
        RECT 153.200 342.200 154.000 346.800 ;
        RECT 156.400 346.300 157.200 346.400 ;
        RECT 161.200 346.300 162.000 346.400 ;
        RECT 156.400 345.700 162.000 346.300 ;
        RECT 156.400 345.600 157.200 345.700 ;
        RECT 161.200 344.800 162.000 345.700 ;
        RECT 162.800 342.200 163.600 349.700 ;
        RECT 166.000 349.600 166.800 349.700 ;
        RECT 167.400 348.400 168.000 352.200 ;
        RECT 172.600 351.600 173.200 355.000 ;
        RECT 174.000 352.400 174.800 359.800 ;
        RECT 174.000 351.800 176.200 352.400 ;
        RECT 177.200 351.800 178.000 359.800 ;
        RECT 180.400 356.400 181.200 359.800 ;
        RECT 180.200 355.800 181.200 356.400 ;
        RECT 180.200 355.200 180.800 355.800 ;
        RECT 183.600 355.200 184.400 359.800 ;
        RECT 186.800 357.000 187.600 359.800 ;
        RECT 188.400 357.000 189.200 359.800 ;
        RECT 169.400 351.000 173.200 351.600 ;
        RECT 175.600 351.200 176.200 351.800 ;
        RECT 169.400 349.000 170.000 351.000 ;
        RECT 175.600 350.400 176.800 351.200 ;
        RECT 166.000 347.600 168.000 348.400 ;
        RECT 168.600 348.200 170.000 349.000 ;
        RECT 170.800 348.800 171.600 350.400 ;
        RECT 172.400 348.800 173.200 350.400 ;
        RECT 174.000 348.800 174.800 350.400 ;
        RECT 167.400 347.000 168.000 347.600 ;
        RECT 169.000 347.800 170.000 348.200 ;
        RECT 169.000 347.200 173.200 347.800 ;
        RECT 175.600 347.400 176.200 350.400 ;
        RECT 177.400 349.600 178.000 351.800 ;
        RECT 167.400 346.600 168.200 347.000 ;
        RECT 167.400 346.000 169.000 346.600 ;
        RECT 168.200 344.400 169.000 346.000 ;
        RECT 172.600 345.000 173.200 347.200 ;
        RECT 168.200 343.600 170.000 344.400 ;
        RECT 168.200 343.000 169.000 343.600 ;
        RECT 172.400 343.000 173.200 345.000 ;
        RECT 174.000 346.800 176.200 347.400 ;
        RECT 174.000 342.200 174.800 346.800 ;
        RECT 177.200 342.200 178.000 349.600 ;
        RECT 178.800 354.600 180.800 355.200 ;
        RECT 178.800 349.000 179.600 354.600 ;
        RECT 181.400 354.400 185.600 355.200 ;
        RECT 190.000 355.000 190.800 359.800 ;
        RECT 193.200 355.000 194.000 359.800 ;
        RECT 181.400 354.000 182.000 354.400 ;
        RECT 180.400 353.200 182.000 354.000 ;
        RECT 185.000 353.800 190.800 354.400 ;
        RECT 183.000 353.200 184.400 353.800 ;
        RECT 183.000 353.000 189.200 353.200 ;
        RECT 183.800 352.600 189.200 353.000 ;
        RECT 188.400 352.400 189.200 352.600 ;
        RECT 190.200 353.000 190.800 353.800 ;
        RECT 191.400 353.600 194.000 354.400 ;
        RECT 196.400 353.600 197.200 359.800 ;
        RECT 198.000 357.000 198.800 359.800 ;
        RECT 199.600 357.000 200.400 359.800 ;
        RECT 201.200 357.000 202.000 359.800 ;
        RECT 199.600 354.400 203.800 355.200 ;
        RECT 204.400 354.400 205.200 359.800 ;
        RECT 207.600 355.200 208.400 359.800 ;
        RECT 207.600 354.600 210.200 355.200 ;
        RECT 204.400 353.600 207.000 354.400 ;
        RECT 198.000 353.000 198.800 353.200 ;
        RECT 190.200 352.400 198.800 353.000 ;
        RECT 201.200 353.000 202.000 353.200 ;
        RECT 209.600 353.000 210.200 354.600 ;
        RECT 201.200 352.400 210.200 353.000 ;
        RECT 209.600 350.600 210.200 352.400 ;
        RECT 210.800 352.000 211.600 359.800 ;
        RECT 215.600 352.800 216.400 359.800 ;
        RECT 210.800 351.200 211.800 352.000 ;
        RECT 180.200 350.000 203.600 350.600 ;
        RECT 209.600 350.000 210.400 350.600 ;
        RECT 180.200 349.800 181.000 350.000 ;
        RECT 185.200 349.600 186.000 350.000 ;
        RECT 202.800 349.400 203.600 350.000 ;
        RECT 178.800 348.200 187.600 349.000 ;
        RECT 188.200 348.600 190.200 349.400 ;
        RECT 194.000 348.600 197.200 349.400 ;
        RECT 178.800 342.200 179.600 348.200 ;
        RECT 181.200 346.800 184.200 347.600 ;
        RECT 183.400 346.200 184.200 346.800 ;
        RECT 189.400 346.200 190.200 348.600 ;
        RECT 191.600 346.800 192.400 348.400 ;
        RECT 196.800 347.800 197.600 348.000 ;
        RECT 193.200 347.200 197.600 347.800 ;
        RECT 193.200 347.000 194.000 347.200 ;
        RECT 199.600 346.400 200.400 349.200 ;
        RECT 205.400 348.600 209.200 349.400 ;
        RECT 205.400 347.400 206.200 348.600 ;
        RECT 209.800 348.000 210.400 350.000 ;
        RECT 193.200 346.200 194.000 346.400 ;
        RECT 183.400 345.400 186.000 346.200 ;
        RECT 189.400 345.600 194.000 346.200 ;
        RECT 194.800 345.600 196.400 346.400 ;
        RECT 199.400 345.600 200.400 346.400 ;
        RECT 204.400 346.800 206.200 347.400 ;
        RECT 209.200 347.400 210.400 348.000 ;
        RECT 204.400 346.200 205.200 346.800 ;
        RECT 185.200 342.200 186.000 345.400 ;
        RECT 202.800 345.400 205.200 346.200 ;
        RECT 186.800 342.200 187.600 345.000 ;
        RECT 188.400 342.200 189.200 345.000 ;
        RECT 190.000 342.200 190.800 345.000 ;
        RECT 193.200 342.200 194.000 345.000 ;
        RECT 196.400 342.200 197.200 345.000 ;
        RECT 198.000 342.200 198.800 345.000 ;
        RECT 199.600 342.200 200.400 345.000 ;
        RECT 201.200 342.200 202.000 345.000 ;
        RECT 202.800 342.200 203.600 345.400 ;
        RECT 209.200 342.200 210.000 347.400 ;
        RECT 211.000 346.800 211.800 351.200 ;
        RECT 215.400 351.800 216.400 352.800 ;
        RECT 218.800 352.400 219.600 359.800 ;
        RECT 217.000 351.800 219.600 352.400 ;
        RECT 215.400 348.400 216.000 351.800 ;
        RECT 217.000 349.800 217.600 351.800 ;
        RECT 222.000 351.200 222.800 359.800 ;
        RECT 225.200 351.200 226.000 359.800 ;
        RECT 228.400 352.400 229.200 359.800 ;
        RECT 231.600 352.800 232.400 359.800 ;
        RECT 236.400 356.400 237.200 359.800 ;
        RECT 236.200 355.800 237.200 356.400 ;
        RECT 236.200 355.200 236.800 355.800 ;
        RECT 239.600 355.200 240.400 359.800 ;
        RECT 242.800 357.000 243.600 359.800 ;
        RECT 244.400 357.000 245.200 359.800 ;
        RECT 234.800 354.600 236.800 355.200 ;
        RECT 228.400 351.800 231.000 352.400 ;
        RECT 231.600 351.800 232.600 352.800 ;
        RECT 222.000 350.400 226.000 351.200 ;
        RECT 216.600 349.000 217.600 349.800 ;
        RECT 212.400 348.300 213.200 348.400 ;
        RECT 215.400 348.300 216.400 348.400 ;
        RECT 212.400 347.700 216.400 348.300 ;
        RECT 212.400 347.600 213.200 347.700 ;
        RECT 215.400 347.600 216.400 347.700 ;
        RECT 210.800 346.000 211.800 346.800 ;
        RECT 215.400 346.200 216.000 347.600 ;
        RECT 217.000 347.400 217.600 349.000 ;
        RECT 218.600 349.600 219.600 350.400 ;
        RECT 218.600 348.800 219.400 349.600 ;
        RECT 222.000 347.600 222.800 350.400 ;
        RECT 228.400 349.600 229.400 350.400 ;
        RECT 228.600 348.800 229.400 349.600 ;
        RECT 230.400 349.800 231.000 351.800 ;
        RECT 230.400 349.000 231.400 349.800 ;
        RECT 217.000 346.800 219.600 347.400 ;
        RECT 210.800 342.200 211.600 346.000 ;
        RECT 215.400 345.600 216.400 346.200 ;
        RECT 215.600 342.200 216.400 345.600 ;
        RECT 218.800 342.200 219.600 346.800 ;
        RECT 222.000 346.800 226.000 347.600 ;
        RECT 230.400 347.400 231.000 349.000 ;
        RECT 232.000 348.400 232.600 351.800 ;
        RECT 234.800 349.000 235.600 354.600 ;
        RECT 237.400 354.400 241.600 355.200 ;
        RECT 246.000 355.000 246.800 359.800 ;
        RECT 249.200 355.000 250.000 359.800 ;
        RECT 237.400 354.000 238.000 354.400 ;
        RECT 236.400 353.200 238.000 354.000 ;
        RECT 241.000 353.800 246.800 354.400 ;
        RECT 239.000 353.200 240.400 353.800 ;
        RECT 239.000 353.000 245.200 353.200 ;
        RECT 239.800 352.600 245.200 353.000 ;
        RECT 244.400 352.400 245.200 352.600 ;
        RECT 246.200 353.000 246.800 353.800 ;
        RECT 247.400 353.600 250.000 354.400 ;
        RECT 252.400 353.600 253.200 359.800 ;
        RECT 254.000 357.000 254.800 359.800 ;
        RECT 255.600 357.000 256.400 359.800 ;
        RECT 257.200 357.000 258.000 359.800 ;
        RECT 255.600 354.400 259.800 355.200 ;
        RECT 260.400 354.400 261.200 359.800 ;
        RECT 263.600 355.200 264.400 359.800 ;
        RECT 263.600 354.600 266.200 355.200 ;
        RECT 260.400 353.600 263.000 354.400 ;
        RECT 254.000 353.000 254.800 353.200 ;
        RECT 246.200 352.400 254.800 353.000 ;
        RECT 257.200 353.000 258.000 353.200 ;
        RECT 265.600 353.000 266.200 354.600 ;
        RECT 257.200 352.400 266.200 353.000 ;
        RECT 265.600 350.600 266.200 352.400 ;
        RECT 266.800 352.000 267.600 359.800 ;
        RECT 270.000 355.000 270.800 359.000 ;
        RECT 266.800 351.200 267.800 352.000 ;
        RECT 236.200 350.000 259.600 350.600 ;
        RECT 265.600 350.000 266.400 350.600 ;
        RECT 236.200 349.800 237.000 350.000 ;
        RECT 238.000 349.600 238.800 350.000 ;
        RECT 241.200 349.600 242.000 350.000 ;
        RECT 258.800 349.400 259.600 350.000 ;
        RECT 231.600 348.300 232.600 348.400 ;
        RECT 233.200 348.300 234.000 348.400 ;
        RECT 231.600 347.700 234.000 348.300 ;
        RECT 231.600 347.600 232.600 347.700 ;
        RECT 233.200 347.600 234.000 347.700 ;
        RECT 234.800 348.200 243.600 349.000 ;
        RECT 244.200 348.600 246.200 349.400 ;
        RECT 250.000 348.600 253.200 349.400 ;
        RECT 222.000 342.200 222.800 346.800 ;
        RECT 225.200 342.200 226.000 346.800 ;
        RECT 228.400 346.800 231.000 347.400 ;
        RECT 228.400 342.200 229.200 346.800 ;
        RECT 232.000 346.200 232.600 347.600 ;
        RECT 231.600 345.600 232.600 346.200 ;
        RECT 231.600 342.200 232.400 345.600 ;
        RECT 234.800 342.200 235.600 348.200 ;
        RECT 237.200 346.800 240.200 347.600 ;
        RECT 239.400 346.200 240.200 346.800 ;
        RECT 245.400 346.200 246.200 348.600 ;
        RECT 247.600 346.800 248.400 348.400 ;
        RECT 252.800 347.800 253.600 348.000 ;
        RECT 249.200 347.200 253.600 347.800 ;
        RECT 249.200 347.000 250.000 347.200 ;
        RECT 255.600 346.400 256.400 349.200 ;
        RECT 261.400 348.600 265.200 349.400 ;
        RECT 261.400 347.400 262.200 348.600 ;
        RECT 265.800 348.000 266.400 350.000 ;
        RECT 249.200 346.200 250.000 346.400 ;
        RECT 239.400 345.400 242.000 346.200 ;
        RECT 245.400 345.600 250.000 346.200 ;
        RECT 250.800 345.600 252.400 346.400 ;
        RECT 255.400 345.600 256.400 346.400 ;
        RECT 260.400 346.800 262.200 347.400 ;
        RECT 265.200 347.400 266.400 348.000 ;
        RECT 260.400 346.200 261.200 346.800 ;
        RECT 241.200 342.200 242.000 345.400 ;
        RECT 258.800 345.400 261.200 346.200 ;
        RECT 242.800 342.200 243.600 345.000 ;
        RECT 244.400 342.200 245.200 345.000 ;
        RECT 246.000 342.200 246.800 345.000 ;
        RECT 249.200 342.200 250.000 345.000 ;
        RECT 252.400 342.200 253.200 345.000 ;
        RECT 254.000 342.200 254.800 345.000 ;
        RECT 255.600 342.200 256.400 345.000 ;
        RECT 257.200 342.200 258.000 345.000 ;
        RECT 258.800 342.200 259.600 345.400 ;
        RECT 265.200 342.200 266.000 347.400 ;
        RECT 267.000 346.800 267.800 351.200 ;
        RECT 270.000 351.600 270.600 355.000 ;
        RECT 274.200 352.800 275.000 359.800 ;
        RECT 274.200 352.200 275.800 352.800 ;
        RECT 270.000 351.000 273.800 351.600 ;
        RECT 270.000 348.800 270.800 350.400 ;
        RECT 271.600 348.800 272.400 350.400 ;
        RECT 273.200 349.000 273.800 351.000 ;
        RECT 273.200 348.200 274.600 349.000 ;
        RECT 275.200 348.400 275.800 352.200 ;
        RECT 276.400 350.300 277.200 351.200 ;
        RECT 279.600 350.300 280.400 359.800 ;
        RECT 276.400 349.700 280.400 350.300 ;
        RECT 276.400 349.600 277.200 349.700 ;
        RECT 273.200 347.800 274.200 348.200 ;
        RECT 266.800 346.000 267.800 346.800 ;
        RECT 270.000 347.200 274.200 347.800 ;
        RECT 275.200 347.600 277.200 348.400 ;
        RECT 266.800 342.200 267.600 346.000 ;
        RECT 270.000 345.000 270.600 347.200 ;
        RECT 275.200 347.000 275.800 347.600 ;
        RECT 275.000 346.600 275.800 347.000 ;
        RECT 274.200 346.400 275.800 346.600 ;
        RECT 273.200 346.000 275.800 346.400 ;
        RECT 273.200 345.600 275.000 346.000 ;
        RECT 270.000 343.000 270.800 345.000 ;
        RECT 274.200 343.000 275.000 345.600 ;
        RECT 279.600 342.200 280.400 349.700 ;
        RECT 281.200 344.800 282.000 346.400 ;
        RECT 282.800 344.800 283.600 346.400 ;
        RECT 284.400 342.200 285.200 359.800 ;
        RECT 287.600 356.400 288.400 359.800 ;
        RECT 287.400 355.800 288.400 356.400 ;
        RECT 287.400 355.200 288.000 355.800 ;
        RECT 290.800 355.200 291.600 359.800 ;
        RECT 294.000 357.000 294.800 359.800 ;
        RECT 295.600 357.000 296.400 359.800 ;
        RECT 286.000 354.600 288.000 355.200 ;
        RECT 286.000 349.000 286.800 354.600 ;
        RECT 288.600 354.400 292.800 355.200 ;
        RECT 297.200 355.000 298.000 359.800 ;
        RECT 300.400 355.000 301.200 359.800 ;
        RECT 288.600 354.000 289.200 354.400 ;
        RECT 287.600 353.200 289.200 354.000 ;
        RECT 292.200 353.800 298.000 354.400 ;
        RECT 290.200 353.200 291.600 353.800 ;
        RECT 290.200 353.000 296.400 353.200 ;
        RECT 291.000 352.600 296.400 353.000 ;
        RECT 295.600 352.400 296.400 352.600 ;
        RECT 297.400 353.000 298.000 353.800 ;
        RECT 298.600 353.600 301.200 354.400 ;
        RECT 303.600 353.600 304.400 359.800 ;
        RECT 305.200 357.000 306.000 359.800 ;
        RECT 306.800 357.000 307.600 359.800 ;
        RECT 308.400 357.000 309.200 359.800 ;
        RECT 306.800 354.400 311.000 355.200 ;
        RECT 311.600 354.400 312.400 359.800 ;
        RECT 314.800 355.200 315.600 359.800 ;
        RECT 314.800 354.600 317.400 355.200 ;
        RECT 311.600 353.600 314.200 354.400 ;
        RECT 305.200 353.000 306.000 353.200 ;
        RECT 297.400 352.400 306.000 353.000 ;
        RECT 308.400 353.000 309.200 353.200 ;
        RECT 316.800 353.000 317.400 354.600 ;
        RECT 308.400 352.400 317.400 353.000 ;
        RECT 316.800 350.600 317.400 352.400 ;
        RECT 318.000 352.000 318.800 359.800 ;
        RECT 326.000 355.000 326.800 359.000 ;
        RECT 318.000 351.200 319.000 352.000 ;
        RECT 287.400 350.000 310.800 350.600 ;
        RECT 316.800 350.000 317.600 350.600 ;
        RECT 287.400 349.800 288.200 350.000 ;
        RECT 289.200 349.600 290.000 350.000 ;
        RECT 292.400 349.600 293.200 350.000 ;
        RECT 310.000 349.400 310.800 350.000 ;
        RECT 286.000 348.200 294.800 349.000 ;
        RECT 295.400 348.600 297.400 349.400 ;
        RECT 301.200 348.600 304.400 349.400 ;
        RECT 286.000 342.200 286.800 348.200 ;
        RECT 288.400 346.800 291.400 347.600 ;
        RECT 290.600 346.200 291.400 346.800 ;
        RECT 296.600 346.200 297.400 348.600 ;
        RECT 298.800 346.800 299.600 348.400 ;
        RECT 304.000 347.800 304.800 348.000 ;
        RECT 300.400 347.200 304.800 347.800 ;
        RECT 300.400 347.000 301.200 347.200 ;
        RECT 306.800 346.400 307.600 349.200 ;
        RECT 312.600 348.600 316.400 349.400 ;
        RECT 312.600 347.400 313.400 348.600 ;
        RECT 317.000 348.000 317.600 350.000 ;
        RECT 300.400 346.200 301.200 346.400 ;
        RECT 290.600 345.400 293.200 346.200 ;
        RECT 296.600 345.600 301.200 346.200 ;
        RECT 302.000 345.600 303.600 346.400 ;
        RECT 306.600 345.600 307.600 346.400 ;
        RECT 311.600 346.800 313.400 347.400 ;
        RECT 316.400 347.400 317.600 348.000 ;
        RECT 311.600 346.200 312.400 346.800 ;
        RECT 292.400 342.200 293.200 345.400 ;
        RECT 310.000 345.400 312.400 346.200 ;
        RECT 294.000 342.200 294.800 345.000 ;
        RECT 295.600 342.200 296.400 345.000 ;
        RECT 297.200 342.200 298.000 345.000 ;
        RECT 300.400 342.200 301.200 345.000 ;
        RECT 303.600 342.200 304.400 345.000 ;
        RECT 305.200 342.200 306.000 345.000 ;
        RECT 306.800 342.200 307.600 345.000 ;
        RECT 308.400 342.200 309.200 345.000 ;
        RECT 310.000 342.200 310.800 345.400 ;
        RECT 316.400 342.200 317.200 347.400 ;
        RECT 318.200 346.800 319.000 351.200 ;
        RECT 326.000 351.600 326.600 355.000 ;
        RECT 330.200 352.800 331.000 359.800 ;
        RECT 330.200 352.200 331.800 352.800 ;
        RECT 326.000 351.000 329.800 351.600 ;
        RECT 321.200 350.300 322.000 350.400 ;
        RECT 324.400 350.300 325.200 350.400 ;
        RECT 326.000 350.300 326.800 350.400 ;
        RECT 321.200 349.700 326.800 350.300 ;
        RECT 321.200 349.600 322.000 349.700 ;
        RECT 324.400 349.600 325.200 349.700 ;
        RECT 326.000 348.800 326.800 349.700 ;
        RECT 327.600 348.800 328.400 350.400 ;
        RECT 329.200 349.000 329.800 351.000 ;
        RECT 329.200 348.200 330.600 349.000 ;
        RECT 331.200 348.400 331.800 352.200 ;
        RECT 332.400 350.300 333.200 351.200 ;
        RECT 335.600 350.300 336.400 359.800 ;
        RECT 340.400 356.400 341.200 359.800 ;
        RECT 340.200 355.800 341.200 356.400 ;
        RECT 340.200 355.200 340.800 355.800 ;
        RECT 343.600 355.200 344.400 359.800 ;
        RECT 346.800 357.000 347.600 359.800 ;
        RECT 348.400 357.000 349.200 359.800 ;
        RECT 332.400 349.700 336.400 350.300 ;
        RECT 332.400 349.600 333.200 349.700 ;
        RECT 329.200 347.800 330.200 348.200 ;
        RECT 318.000 346.000 319.000 346.800 ;
        RECT 326.000 347.200 330.200 347.800 ;
        RECT 331.200 347.600 333.200 348.400 ;
        RECT 318.000 342.200 318.800 346.000 ;
        RECT 326.000 345.000 326.600 347.200 ;
        RECT 331.200 347.000 331.800 347.600 ;
        RECT 331.000 346.600 331.800 347.000 ;
        RECT 330.200 346.400 331.800 346.600 ;
        RECT 329.200 346.000 331.800 346.400 ;
        RECT 329.200 345.600 331.000 346.000 ;
        RECT 326.000 343.000 326.800 345.000 ;
        RECT 330.200 343.000 331.000 345.600 ;
        RECT 335.600 342.200 336.400 349.700 ;
        RECT 338.800 354.600 340.800 355.200 ;
        RECT 338.800 349.000 339.600 354.600 ;
        RECT 341.400 354.400 345.600 355.200 ;
        RECT 350.000 355.000 350.800 359.800 ;
        RECT 353.200 355.000 354.000 359.800 ;
        RECT 341.400 354.000 342.000 354.400 ;
        RECT 340.400 353.200 342.000 354.000 ;
        RECT 345.000 353.800 350.800 354.400 ;
        RECT 343.000 353.200 344.400 353.800 ;
        RECT 343.000 353.000 349.200 353.200 ;
        RECT 343.800 352.600 349.200 353.000 ;
        RECT 348.400 352.400 349.200 352.600 ;
        RECT 350.200 353.000 350.800 353.800 ;
        RECT 351.400 353.600 354.000 354.400 ;
        RECT 356.400 353.600 357.200 359.800 ;
        RECT 358.000 357.000 358.800 359.800 ;
        RECT 359.600 357.000 360.400 359.800 ;
        RECT 361.200 357.000 362.000 359.800 ;
        RECT 359.600 354.400 363.800 355.200 ;
        RECT 364.400 354.400 365.200 359.800 ;
        RECT 367.600 355.200 368.400 359.800 ;
        RECT 367.600 354.600 370.200 355.200 ;
        RECT 364.400 353.600 367.000 354.400 ;
        RECT 358.000 353.000 358.800 353.200 ;
        RECT 350.200 352.400 358.800 353.000 ;
        RECT 361.200 353.000 362.000 353.200 ;
        RECT 369.600 353.000 370.200 354.600 ;
        RECT 361.200 352.400 370.200 353.000 ;
        RECT 369.600 350.600 370.200 352.400 ;
        RECT 370.800 352.000 371.600 359.800 ;
        RECT 370.800 351.200 371.800 352.000 ;
        RECT 340.200 350.000 363.600 350.600 ;
        RECT 369.600 350.000 370.400 350.600 ;
        RECT 340.200 349.800 341.000 350.000 ;
        RECT 343.600 349.600 344.400 350.000 ;
        RECT 345.200 349.600 346.000 350.000 ;
        RECT 362.800 349.400 363.600 350.000 ;
        RECT 338.800 348.200 347.600 349.000 ;
        RECT 348.200 348.600 350.200 349.400 ;
        RECT 354.000 348.600 357.200 349.400 ;
        RECT 337.200 344.800 338.000 346.400 ;
        RECT 338.800 342.200 339.600 348.200 ;
        RECT 341.200 346.800 344.200 347.600 ;
        RECT 343.400 346.200 344.200 346.800 ;
        RECT 349.400 346.200 350.200 348.600 ;
        RECT 351.600 346.800 352.400 348.400 ;
        RECT 356.800 347.800 357.600 348.000 ;
        RECT 353.200 347.200 357.600 347.800 ;
        RECT 353.200 347.000 354.000 347.200 ;
        RECT 359.600 346.400 360.400 349.200 ;
        RECT 365.400 348.600 369.200 349.400 ;
        RECT 365.400 347.400 366.200 348.600 ;
        RECT 369.800 348.000 370.400 350.000 ;
        RECT 353.200 346.200 354.000 346.400 ;
        RECT 343.400 345.400 346.000 346.200 ;
        RECT 349.400 345.600 354.000 346.200 ;
        RECT 354.800 345.600 356.400 346.400 ;
        RECT 359.400 345.600 360.400 346.400 ;
        RECT 364.400 346.800 366.200 347.400 ;
        RECT 369.200 347.400 370.400 348.000 ;
        RECT 364.400 346.200 365.200 346.800 ;
        RECT 345.200 342.200 346.000 345.400 ;
        RECT 362.800 345.400 365.200 346.200 ;
        RECT 346.800 342.200 347.600 345.000 ;
        RECT 348.400 342.200 349.200 345.000 ;
        RECT 350.000 342.200 350.800 345.000 ;
        RECT 353.200 342.200 354.000 345.000 ;
        RECT 356.400 342.200 357.200 345.000 ;
        RECT 358.000 342.200 358.800 345.000 ;
        RECT 359.600 342.200 360.400 345.000 ;
        RECT 361.200 342.200 362.000 345.000 ;
        RECT 362.800 342.200 363.600 345.400 ;
        RECT 369.200 342.200 370.000 347.400 ;
        RECT 371.000 346.800 371.800 351.200 ;
        RECT 370.800 346.000 371.800 346.800 ;
        RECT 375.600 348.300 376.400 359.800 ;
        RECT 377.200 348.300 378.000 348.400 ;
        RECT 375.600 347.700 378.000 348.300 ;
        RECT 370.800 342.200 371.600 346.000 ;
        RECT 374.000 344.800 374.800 346.400 ;
        RECT 375.600 342.200 376.400 347.700 ;
        RECT 377.200 346.800 378.000 347.700 ;
        RECT 378.800 346.200 379.600 359.800 ;
        RECT 380.400 351.600 381.200 353.200 ;
        RECT 385.800 352.800 386.600 359.800 ;
        RECT 390.000 355.000 390.800 359.000 ;
        RECT 385.000 352.200 386.600 352.800 ;
        RECT 382.000 350.300 382.800 350.400 ;
        RECT 383.600 350.300 384.400 351.200 ;
        RECT 382.000 349.700 384.400 350.300 ;
        RECT 382.000 349.600 382.800 349.700 ;
        RECT 383.600 349.600 384.400 349.700 ;
        RECT 385.000 348.400 385.600 352.200 ;
        RECT 390.200 351.600 390.800 355.000 ;
        RECT 395.400 352.800 396.200 359.800 ;
        RECT 399.600 355.000 400.400 359.000 ;
        RECT 387.000 351.000 390.800 351.600 ;
        RECT 394.600 352.200 396.200 352.800 ;
        RECT 394.600 351.600 395.600 352.200 ;
        RECT 399.800 351.600 400.400 355.000 ;
        RECT 401.200 351.600 402.000 353.200 ;
        RECT 387.000 349.000 387.600 351.000 ;
        RECT 380.400 348.300 381.200 348.400 ;
        RECT 383.600 348.300 385.600 348.400 ;
        RECT 380.400 347.700 385.600 348.300 ;
        RECT 386.200 348.200 387.600 349.000 ;
        RECT 388.400 348.800 389.200 350.400 ;
        RECT 390.000 348.800 390.800 350.400 ;
        RECT 393.200 349.600 394.000 351.200 ;
        RECT 394.600 348.400 395.200 351.600 ;
        RECT 396.600 351.000 400.400 351.600 ;
        RECT 396.600 349.000 397.200 351.000 ;
        RECT 380.400 347.600 381.200 347.700 ;
        RECT 383.600 347.600 385.600 347.700 ;
        RECT 385.000 347.000 385.600 347.600 ;
        RECT 386.600 347.800 387.600 348.200 ;
        RECT 386.600 347.200 390.800 347.800 ;
        RECT 393.200 347.600 395.200 348.400 ;
        RECT 395.800 348.200 397.200 349.000 ;
        RECT 398.000 348.800 398.800 350.400 ;
        RECT 399.600 348.800 400.400 350.400 ;
        RECT 385.000 346.600 385.800 347.000 ;
        RECT 378.800 345.600 380.600 346.200 ;
        RECT 385.000 346.000 386.600 346.600 ;
        RECT 379.800 344.400 380.600 345.600 ;
        RECT 379.800 343.600 381.200 344.400 ;
        RECT 379.800 342.200 380.600 343.600 ;
        RECT 385.800 343.000 386.600 346.000 ;
        RECT 390.200 345.000 390.800 347.200 ;
        RECT 394.600 347.000 395.200 347.600 ;
        RECT 396.200 347.800 397.200 348.200 ;
        RECT 396.200 347.200 400.400 347.800 ;
        RECT 394.600 346.600 395.400 347.000 ;
        RECT 394.600 346.000 396.200 346.600 ;
        RECT 390.000 343.000 390.800 345.000 ;
        RECT 395.400 343.000 396.200 346.000 ;
        RECT 399.800 345.000 400.400 347.200 ;
        RECT 402.800 346.200 403.600 359.800 ;
        RECT 406.000 352.300 406.800 359.800 ;
        RECT 407.600 352.300 408.400 352.400 ;
        RECT 406.000 351.700 408.400 352.300 ;
        RECT 404.400 346.800 405.200 348.400 ;
        RECT 399.600 343.000 400.400 345.000 ;
        RECT 401.800 345.600 403.600 346.200 ;
        RECT 401.800 344.400 402.600 345.600 ;
        RECT 401.800 343.600 403.600 344.400 ;
        RECT 401.800 342.200 402.600 343.600 ;
        RECT 406.000 342.200 406.800 351.700 ;
        RECT 407.600 351.600 408.400 351.700 ;
        RECT 409.200 346.800 410.000 348.400 ;
        RECT 407.600 344.800 408.400 346.400 ;
        RECT 410.800 346.200 411.600 359.800 ;
        RECT 412.400 351.600 413.200 353.200 ;
        RECT 415.600 352.000 416.400 359.800 ;
        RECT 418.800 355.200 419.600 359.800 ;
        RECT 415.400 351.200 416.400 352.000 ;
        RECT 417.000 354.600 419.600 355.200 ;
        RECT 417.000 353.000 417.600 354.600 ;
        RECT 422.000 354.400 422.800 359.800 ;
        RECT 425.200 357.000 426.000 359.800 ;
        RECT 426.800 357.000 427.600 359.800 ;
        RECT 428.400 357.000 429.200 359.800 ;
        RECT 423.400 354.400 427.600 355.200 ;
        RECT 420.200 353.600 422.800 354.400 ;
        RECT 430.000 353.600 430.800 359.800 ;
        RECT 433.200 355.000 434.000 359.800 ;
        RECT 436.400 355.000 437.200 359.800 ;
        RECT 438.000 357.000 438.800 359.800 ;
        RECT 439.600 357.000 440.400 359.800 ;
        RECT 442.800 355.200 443.600 359.800 ;
        RECT 446.000 356.400 446.800 359.800 ;
        RECT 451.800 358.400 452.600 359.800 ;
        RECT 450.800 357.600 452.600 358.400 ;
        RECT 446.000 355.800 447.000 356.400 ;
        RECT 446.400 355.200 447.000 355.800 ;
        RECT 441.600 354.400 445.800 355.200 ;
        RECT 446.400 354.600 448.400 355.200 ;
        RECT 433.200 353.600 435.800 354.400 ;
        RECT 436.400 353.800 442.200 354.400 ;
        RECT 445.200 354.000 445.800 354.400 ;
        RECT 425.200 353.000 426.000 353.200 ;
        RECT 417.000 352.400 426.000 353.000 ;
        RECT 428.400 353.000 429.200 353.200 ;
        RECT 436.400 353.000 437.000 353.800 ;
        RECT 442.800 353.200 444.200 353.800 ;
        RECT 445.200 353.200 446.800 354.000 ;
        RECT 428.400 352.400 437.000 353.000 ;
        RECT 438.000 353.000 444.200 353.200 ;
        RECT 438.000 352.600 443.400 353.000 ;
        RECT 438.000 352.400 438.800 352.600 ;
        RECT 415.400 346.800 416.200 351.200 ;
        RECT 417.000 350.600 417.600 352.400 ;
        RECT 416.800 350.000 417.600 350.600 ;
        RECT 423.600 350.000 447.000 350.600 ;
        RECT 416.800 348.000 417.400 350.000 ;
        RECT 423.600 349.400 424.400 350.000 ;
        RECT 441.200 349.600 442.000 350.000 ;
        RECT 442.800 349.600 443.600 350.000 ;
        RECT 446.200 349.800 447.000 350.000 ;
        RECT 418.000 348.600 421.800 349.400 ;
        RECT 416.800 347.400 418.000 348.000 ;
        RECT 410.800 345.600 412.600 346.200 ;
        RECT 415.400 346.000 416.400 346.800 ;
        RECT 411.800 344.400 412.600 345.600 ;
        RECT 410.800 343.600 412.600 344.400 ;
        RECT 411.800 342.200 412.600 343.600 ;
        RECT 415.600 342.200 416.400 346.000 ;
        RECT 417.200 342.200 418.000 347.400 ;
        RECT 421.000 347.400 421.800 348.600 ;
        RECT 421.000 346.800 422.800 347.400 ;
        RECT 422.000 346.200 422.800 346.800 ;
        RECT 426.800 346.400 427.600 349.200 ;
        RECT 430.000 348.600 433.200 349.400 ;
        RECT 437.000 348.600 439.000 349.400 ;
        RECT 447.600 349.000 448.400 354.600 ;
        RECT 451.800 352.600 452.600 357.600 ;
        RECT 450.800 351.800 452.600 352.600 ;
        RECT 460.400 352.000 461.200 359.800 ;
        RECT 463.600 355.200 464.400 359.800 ;
        RECT 429.600 347.800 430.400 348.000 ;
        RECT 429.600 347.200 434.000 347.800 ;
        RECT 433.200 347.000 434.000 347.200 ;
        RECT 434.800 346.800 435.600 348.400 ;
        RECT 422.000 345.400 424.400 346.200 ;
        RECT 426.800 345.600 427.800 346.400 ;
        RECT 430.800 345.600 432.400 346.400 ;
        RECT 433.200 346.200 434.000 346.400 ;
        RECT 437.000 346.200 437.800 348.600 ;
        RECT 439.600 348.200 448.400 349.000 ;
        RECT 451.000 348.400 451.600 351.800 ;
        RECT 460.200 351.200 461.200 352.000 ;
        RECT 461.800 354.600 464.400 355.200 ;
        RECT 461.800 353.000 462.400 354.600 ;
        RECT 466.800 354.400 467.600 359.800 ;
        RECT 470.000 357.000 470.800 359.800 ;
        RECT 471.600 357.000 472.400 359.800 ;
        RECT 473.200 357.000 474.000 359.800 ;
        RECT 468.200 354.400 472.400 355.200 ;
        RECT 465.000 353.600 467.600 354.400 ;
        RECT 474.800 353.600 475.600 359.800 ;
        RECT 478.000 355.000 478.800 359.800 ;
        RECT 481.200 355.000 482.000 359.800 ;
        RECT 482.800 357.000 483.600 359.800 ;
        RECT 484.400 357.000 485.200 359.800 ;
        RECT 487.600 355.200 488.400 359.800 ;
        RECT 490.800 356.400 491.600 359.800 ;
        RECT 495.600 356.400 496.400 359.800 ;
        RECT 490.800 355.800 491.800 356.400 ;
        RECT 491.200 355.200 491.800 355.800 ;
        RECT 495.400 355.800 496.400 356.400 ;
        RECT 495.400 355.200 496.000 355.800 ;
        RECT 498.800 355.200 499.600 359.800 ;
        RECT 502.000 357.000 502.800 359.800 ;
        RECT 503.600 357.000 504.400 359.800 ;
        RECT 486.400 354.400 490.600 355.200 ;
        RECT 491.200 354.600 493.200 355.200 ;
        RECT 478.000 353.600 480.600 354.400 ;
        RECT 481.200 353.800 487.000 354.400 ;
        RECT 490.000 354.000 490.600 354.400 ;
        RECT 470.000 353.000 470.800 353.200 ;
        RECT 461.800 352.400 470.800 353.000 ;
        RECT 473.200 353.000 474.000 353.200 ;
        RECT 481.200 353.000 481.800 353.800 ;
        RECT 487.600 353.200 489.000 353.800 ;
        RECT 490.000 353.200 491.600 354.000 ;
        RECT 473.200 352.400 481.800 353.000 ;
        RECT 482.800 353.000 489.000 353.200 ;
        RECT 482.800 352.600 488.200 353.000 ;
        RECT 482.800 352.400 483.600 352.600 ;
        RECT 452.400 350.300 453.200 351.200 ;
        RECT 460.200 350.300 461.000 351.200 ;
        RECT 461.800 350.600 462.400 352.400 ;
        RECT 452.400 349.700 461.000 350.300 ;
        RECT 452.400 349.600 453.200 349.700 ;
        RECT 443.000 346.800 446.000 347.600 ;
        RECT 443.000 346.200 443.800 346.800 ;
        RECT 433.200 345.600 437.800 346.200 ;
        RECT 423.600 342.200 424.400 345.400 ;
        RECT 441.200 345.400 443.800 346.200 ;
        RECT 425.200 342.200 426.000 345.000 ;
        RECT 426.800 342.200 427.600 345.000 ;
        RECT 428.400 342.200 429.200 345.000 ;
        RECT 430.000 342.200 430.800 345.000 ;
        RECT 433.200 342.200 434.000 345.000 ;
        RECT 436.400 342.200 437.200 345.000 ;
        RECT 438.000 342.200 438.800 345.000 ;
        RECT 439.600 342.200 440.400 345.000 ;
        RECT 441.200 342.200 442.000 345.400 ;
        RECT 447.600 342.200 448.400 348.200 ;
        RECT 450.800 347.600 451.600 348.400 ;
        RECT 449.200 344.800 450.000 346.400 ;
        RECT 451.000 344.200 451.600 347.600 ;
        RECT 460.200 346.800 461.000 349.700 ;
        RECT 461.600 350.000 462.400 350.600 ;
        RECT 468.400 350.000 491.800 350.600 ;
        RECT 461.600 348.000 462.200 350.000 ;
        RECT 468.400 349.400 469.200 350.000 ;
        RECT 486.000 349.600 486.800 350.000 ;
        RECT 489.200 349.600 490.000 350.000 ;
        RECT 491.000 349.800 491.800 350.000 ;
        RECT 462.800 348.600 466.600 349.400 ;
        RECT 461.600 347.400 462.800 348.000 ;
        RECT 460.200 346.000 461.200 346.800 ;
        RECT 450.800 342.200 451.600 344.200 ;
        RECT 460.400 342.200 461.200 346.000 ;
        RECT 462.000 342.200 462.800 347.400 ;
        RECT 465.800 347.400 466.600 348.600 ;
        RECT 465.800 346.800 467.600 347.400 ;
        RECT 466.800 346.200 467.600 346.800 ;
        RECT 471.600 346.400 472.400 349.200 ;
        RECT 474.800 348.600 478.000 349.400 ;
        RECT 481.800 348.600 483.800 349.400 ;
        RECT 492.400 349.000 493.200 354.600 ;
        RECT 474.400 347.800 475.200 348.000 ;
        RECT 474.400 347.200 478.800 347.800 ;
        RECT 478.000 347.000 478.800 347.200 ;
        RECT 479.600 346.800 480.400 348.400 ;
        RECT 466.800 345.400 469.200 346.200 ;
        RECT 471.600 345.600 472.600 346.400 ;
        RECT 475.600 345.600 477.200 346.400 ;
        RECT 478.000 346.200 478.800 346.400 ;
        RECT 481.800 346.200 482.600 348.600 ;
        RECT 484.400 348.200 493.200 349.000 ;
        RECT 487.800 346.800 490.800 347.600 ;
        RECT 487.800 346.200 488.600 346.800 ;
        RECT 478.000 345.600 482.600 346.200 ;
        RECT 468.400 342.200 469.200 345.400 ;
        RECT 486.000 345.400 488.600 346.200 ;
        RECT 470.000 342.200 470.800 345.000 ;
        RECT 471.600 342.200 472.400 345.000 ;
        RECT 473.200 342.200 474.000 345.000 ;
        RECT 474.800 342.200 475.600 345.000 ;
        RECT 478.000 342.200 478.800 345.000 ;
        RECT 481.200 342.200 482.000 345.000 ;
        RECT 482.800 342.200 483.600 345.000 ;
        RECT 484.400 342.200 485.200 345.000 ;
        RECT 486.000 342.200 486.800 345.400 ;
        RECT 492.400 342.200 493.200 348.200 ;
        RECT 494.000 354.600 496.000 355.200 ;
        RECT 494.000 349.000 494.800 354.600 ;
        RECT 496.600 354.400 500.800 355.200 ;
        RECT 505.200 355.000 506.000 359.800 ;
        RECT 508.400 355.000 509.200 359.800 ;
        RECT 496.600 354.000 497.200 354.400 ;
        RECT 495.600 353.200 497.200 354.000 ;
        RECT 500.200 353.800 506.000 354.400 ;
        RECT 498.200 353.200 499.600 353.800 ;
        RECT 498.200 353.000 504.400 353.200 ;
        RECT 499.000 352.600 504.400 353.000 ;
        RECT 503.600 352.400 504.400 352.600 ;
        RECT 505.400 353.000 506.000 353.800 ;
        RECT 506.600 353.600 509.200 354.400 ;
        RECT 511.600 353.600 512.400 359.800 ;
        RECT 513.200 357.000 514.000 359.800 ;
        RECT 514.800 357.000 515.600 359.800 ;
        RECT 516.400 357.000 517.200 359.800 ;
        RECT 514.800 354.400 519.000 355.200 ;
        RECT 519.600 354.400 520.400 359.800 ;
        RECT 522.800 355.200 523.600 359.800 ;
        RECT 522.800 354.600 525.400 355.200 ;
        RECT 519.600 353.600 522.200 354.400 ;
        RECT 513.200 353.000 514.000 353.200 ;
        RECT 505.400 352.400 514.000 353.000 ;
        RECT 516.400 353.000 517.200 353.200 ;
        RECT 524.800 353.000 525.400 354.600 ;
        RECT 516.400 352.400 525.400 353.000 ;
        RECT 524.800 350.600 525.400 352.400 ;
        RECT 526.000 352.000 526.800 359.800 ;
        RECT 526.000 351.200 527.000 352.000 ;
        RECT 495.400 350.000 518.800 350.600 ;
        RECT 524.800 350.000 525.600 350.600 ;
        RECT 495.400 349.800 496.400 350.000 ;
        RECT 495.600 349.600 496.400 349.800 ;
        RECT 500.400 349.600 501.200 350.000 ;
        RECT 518.000 349.400 518.800 350.000 ;
        RECT 494.000 348.200 502.800 349.000 ;
        RECT 503.400 348.600 505.400 349.400 ;
        RECT 509.200 348.600 512.400 349.400 ;
        RECT 494.000 342.200 494.800 348.200 ;
        RECT 496.400 346.800 499.400 347.600 ;
        RECT 498.600 346.200 499.400 346.800 ;
        RECT 504.600 346.200 505.400 348.600 ;
        RECT 506.800 346.800 507.600 348.400 ;
        RECT 512.000 347.800 512.800 348.000 ;
        RECT 508.400 347.200 512.800 347.800 ;
        RECT 508.400 347.000 509.200 347.200 ;
        RECT 514.800 346.400 515.600 349.200 ;
        RECT 520.600 348.600 524.400 349.400 ;
        RECT 520.600 347.400 521.400 348.600 ;
        RECT 525.000 348.000 525.600 350.000 ;
        RECT 508.400 346.200 509.200 346.400 ;
        RECT 498.600 345.400 501.200 346.200 ;
        RECT 504.600 345.600 509.200 346.200 ;
        RECT 510.000 345.600 511.600 346.400 ;
        RECT 514.600 345.600 515.600 346.400 ;
        RECT 519.600 346.800 521.400 347.400 ;
        RECT 524.400 347.400 525.600 348.000 ;
        RECT 519.600 346.200 520.400 346.800 ;
        RECT 500.400 342.200 501.200 345.400 ;
        RECT 518.000 345.400 520.400 346.200 ;
        RECT 502.000 342.200 502.800 345.000 ;
        RECT 503.600 342.200 504.400 345.000 ;
        RECT 505.200 342.200 506.000 345.000 ;
        RECT 508.400 342.200 509.200 345.000 ;
        RECT 511.600 342.200 512.400 345.000 ;
        RECT 513.200 342.200 514.000 345.000 ;
        RECT 514.800 342.200 515.600 345.000 ;
        RECT 516.400 342.200 517.200 345.000 ;
        RECT 518.000 342.200 518.800 345.400 ;
        RECT 524.400 342.200 525.200 347.400 ;
        RECT 526.200 346.800 527.000 351.200 ;
        RECT 529.200 346.800 530.000 348.400 ;
        RECT 526.000 346.000 527.000 346.800 ;
        RECT 530.800 346.200 531.600 359.800 ;
        RECT 532.400 351.600 533.200 353.200 ;
        RECT 535.600 352.800 536.400 359.800 ;
        RECT 535.400 351.800 536.400 352.800 ;
        RECT 538.800 352.400 539.600 359.800 ;
        RECT 537.000 351.800 539.600 352.400 ;
        RECT 540.400 352.400 541.200 359.800 ;
        RECT 543.600 352.800 544.400 359.800 ;
        RECT 540.400 351.800 543.000 352.400 ;
        RECT 543.600 351.800 544.600 352.800 ;
        RECT 535.400 348.400 536.000 351.800 ;
        RECT 537.000 349.800 537.600 351.800 ;
        RECT 536.600 349.000 537.600 349.800 ;
        RECT 535.400 347.600 536.400 348.400 ;
        RECT 535.400 346.200 536.000 347.600 ;
        RECT 537.000 347.400 537.600 349.000 ;
        RECT 538.600 349.600 539.600 350.400 ;
        RECT 540.400 349.600 541.400 350.400 ;
        RECT 538.600 348.800 539.400 349.600 ;
        RECT 540.600 348.800 541.400 349.600 ;
        RECT 542.400 349.800 543.000 351.800 ;
        RECT 542.400 349.000 543.400 349.800 ;
        RECT 542.400 347.400 543.000 349.000 ;
        RECT 544.000 348.400 544.600 351.800 ;
        RECT 548.400 351.200 549.200 359.800 ;
        RECT 551.600 351.200 552.400 359.800 ;
        RECT 554.800 351.600 555.600 353.200 ;
        RECT 548.400 350.400 552.400 351.200 ;
        RECT 543.600 347.600 544.600 348.400 ;
        RECT 551.600 347.600 552.400 350.400 ;
        RECT 537.000 346.800 539.600 347.400 ;
        RECT 526.000 342.200 526.800 346.000 ;
        RECT 530.800 345.600 532.600 346.200 ;
        RECT 535.400 345.600 536.400 346.200 ;
        RECT 531.800 344.400 532.600 345.600 ;
        RECT 530.800 343.600 532.600 344.400 ;
        RECT 531.800 342.200 532.600 343.600 ;
        RECT 535.600 342.200 536.400 345.600 ;
        RECT 538.800 342.200 539.600 346.800 ;
        RECT 540.400 346.800 543.000 347.400 ;
        RECT 540.400 342.200 541.200 346.800 ;
        RECT 544.000 346.200 544.600 347.600 ;
        RECT 543.600 345.600 544.600 346.200 ;
        RECT 548.400 346.800 552.400 347.600 ;
        RECT 543.600 342.200 544.400 345.600 ;
        RECT 548.400 342.200 549.200 346.800 ;
        RECT 551.600 342.200 552.400 346.800 ;
        RECT 556.400 346.200 557.200 359.800 ;
        RECT 562.200 352.400 563.000 359.800 ;
        RECT 567.600 356.400 568.400 359.800 ;
        RECT 567.400 355.800 568.400 356.400 ;
        RECT 567.400 355.200 568.000 355.800 ;
        RECT 570.800 355.200 571.600 359.800 ;
        RECT 574.000 357.000 574.800 359.800 ;
        RECT 575.600 357.000 576.400 359.800 ;
        RECT 566.000 354.600 568.000 355.200 ;
        RECT 563.600 353.600 564.400 354.400 ;
        RECT 563.800 352.400 564.400 353.600 ;
        RECT 561.200 351.600 563.200 352.400 ;
        RECT 563.800 351.800 565.200 352.400 ;
        RECT 564.400 351.600 565.200 351.800 ;
        RECT 559.600 350.300 560.400 350.400 ;
        RECT 561.200 350.300 562.000 350.400 ;
        RECT 559.600 349.700 562.000 350.300 ;
        RECT 559.600 349.600 560.400 349.700 ;
        RECT 561.200 348.800 562.000 349.700 ;
        RECT 562.600 348.400 563.200 351.600 ;
        RECT 566.000 349.000 566.800 354.600 ;
        RECT 568.600 354.400 572.800 355.200 ;
        RECT 577.200 355.000 578.000 359.800 ;
        RECT 580.400 355.000 581.200 359.800 ;
        RECT 568.600 354.000 569.200 354.400 ;
        RECT 567.600 353.200 569.200 354.000 ;
        RECT 572.200 353.800 578.000 354.400 ;
        RECT 570.200 353.200 571.600 353.800 ;
        RECT 570.200 353.000 576.400 353.200 ;
        RECT 571.000 352.600 576.400 353.000 ;
        RECT 575.600 352.400 576.400 352.600 ;
        RECT 577.400 353.000 578.000 353.800 ;
        RECT 578.600 353.600 581.200 354.400 ;
        RECT 583.600 353.600 584.400 359.800 ;
        RECT 585.200 357.000 586.000 359.800 ;
        RECT 586.800 357.000 587.600 359.800 ;
        RECT 588.400 357.000 589.200 359.800 ;
        RECT 586.800 354.400 591.000 355.200 ;
        RECT 591.600 354.400 592.400 359.800 ;
        RECT 594.800 355.200 595.600 359.800 ;
        RECT 594.800 354.600 597.400 355.200 ;
        RECT 591.600 353.600 594.200 354.400 ;
        RECT 585.200 353.000 586.000 353.200 ;
        RECT 577.400 352.400 586.000 353.000 ;
        RECT 588.400 353.000 589.200 353.200 ;
        RECT 596.800 353.000 597.400 354.600 ;
        RECT 588.400 352.400 597.400 353.000 ;
        RECT 596.800 350.600 597.400 352.400 ;
        RECT 598.000 352.000 598.800 359.800 ;
        RECT 598.000 351.200 599.000 352.000 ;
        RECT 567.400 350.000 590.800 350.600 ;
        RECT 596.800 350.000 597.600 350.600 ;
        RECT 567.400 349.800 568.400 350.000 ;
        RECT 567.600 349.600 568.400 349.800 ;
        RECT 572.400 349.600 573.200 350.000 ;
        RECT 578.800 349.600 579.600 350.000 ;
        RECT 590.000 349.400 590.800 350.000 ;
        RECT 558.000 346.800 558.800 348.400 ;
        RECT 559.600 348.200 560.400 348.400 ;
        RECT 559.600 347.600 561.200 348.200 ;
        RECT 562.600 347.600 565.200 348.400 ;
        RECT 566.000 348.200 574.800 349.000 ;
        RECT 575.400 348.600 577.400 349.400 ;
        RECT 581.200 348.600 584.400 349.400 ;
        RECT 560.400 347.200 561.200 347.600 ;
        RECT 559.800 346.200 563.400 346.600 ;
        RECT 564.400 346.200 565.000 347.600 ;
        RECT 555.400 345.600 557.200 346.200 ;
        RECT 559.600 346.000 563.600 346.200 ;
        RECT 555.400 344.400 556.200 345.600 ;
        RECT 554.800 343.600 556.200 344.400 ;
        RECT 555.400 342.200 556.200 343.600 ;
        RECT 559.600 342.200 560.400 346.000 ;
        RECT 562.800 342.200 563.600 346.000 ;
        RECT 564.400 342.200 565.200 346.200 ;
        RECT 566.000 342.200 566.800 348.200 ;
        RECT 568.400 346.800 571.400 347.600 ;
        RECT 570.600 346.200 571.400 346.800 ;
        RECT 576.600 346.200 577.400 348.600 ;
        RECT 578.800 346.800 579.600 348.400 ;
        RECT 584.000 347.800 584.800 348.000 ;
        RECT 580.400 347.200 584.800 347.800 ;
        RECT 580.400 347.000 581.200 347.200 ;
        RECT 586.800 346.400 587.600 349.200 ;
        RECT 592.600 348.600 596.400 349.400 ;
        RECT 592.600 347.400 593.400 348.600 ;
        RECT 597.000 348.000 597.600 350.000 ;
        RECT 580.400 346.200 581.200 346.400 ;
        RECT 570.600 345.400 573.200 346.200 ;
        RECT 576.600 345.600 581.200 346.200 ;
        RECT 582.000 345.600 583.600 346.400 ;
        RECT 586.600 345.600 587.600 346.400 ;
        RECT 591.600 346.800 593.400 347.400 ;
        RECT 596.400 347.400 597.600 348.000 ;
        RECT 591.600 346.200 592.400 346.800 ;
        RECT 572.400 342.200 573.200 345.400 ;
        RECT 590.000 345.400 592.400 346.200 ;
        RECT 574.000 342.200 574.800 345.000 ;
        RECT 575.600 342.200 576.400 345.000 ;
        RECT 577.200 342.200 578.000 345.000 ;
        RECT 580.400 342.200 581.200 345.000 ;
        RECT 583.600 342.200 584.400 345.000 ;
        RECT 585.200 342.200 586.000 345.000 ;
        RECT 586.800 342.200 587.600 345.000 ;
        RECT 588.400 342.200 589.200 345.000 ;
        RECT 590.000 342.200 590.800 345.400 ;
        RECT 596.400 342.200 597.200 347.400 ;
        RECT 598.200 346.800 599.000 351.200 ;
        RECT 599.600 348.300 600.400 348.400 ;
        RECT 601.200 348.300 602.000 348.400 ;
        RECT 599.600 347.700 602.000 348.300 ;
        RECT 599.600 347.600 600.400 347.700 ;
        RECT 601.200 346.800 602.000 347.700 ;
        RECT 598.000 346.000 599.000 346.800 ;
        RECT 602.800 346.200 603.600 359.800 ;
        RECT 604.400 351.600 605.200 353.200 ;
        RECT 606.000 352.400 606.800 359.800 ;
        RECT 606.000 351.800 608.200 352.400 ;
        RECT 607.600 351.200 608.200 351.800 ;
        RECT 607.600 350.400 608.800 351.200 ;
        RECT 604.400 350.300 605.200 350.400 ;
        RECT 606.000 350.300 606.800 350.400 ;
        RECT 604.400 349.700 606.800 350.300 ;
        RECT 604.400 349.600 605.200 349.700 ;
        RECT 606.000 348.800 606.800 349.700 ;
        RECT 607.600 347.400 608.200 350.400 ;
        RECT 606.000 346.800 608.200 347.400 ;
        RECT 598.000 342.200 598.800 346.000 ;
        RECT 602.800 345.600 604.600 346.200 ;
        RECT 603.800 344.400 604.600 345.600 ;
        RECT 602.800 343.600 604.600 344.400 ;
        RECT 603.800 342.200 604.600 343.600 ;
        RECT 606.000 342.200 606.800 346.800 ;
        RECT 1.200 333.800 2.000 339.800 ;
        RECT 7.600 336.600 8.400 339.800 ;
        RECT 9.200 337.000 10.000 339.800 ;
        RECT 10.800 337.000 11.600 339.800 ;
        RECT 12.400 337.000 13.200 339.800 ;
        RECT 15.600 337.000 16.400 339.800 ;
        RECT 18.800 337.000 19.600 339.800 ;
        RECT 20.400 337.000 21.200 339.800 ;
        RECT 22.000 337.000 22.800 339.800 ;
        RECT 23.600 337.000 24.400 339.800 ;
        RECT 5.800 335.800 8.400 336.600 ;
        RECT 25.200 336.600 26.000 339.800 ;
        RECT 11.800 335.800 16.400 336.400 ;
        RECT 5.800 335.200 6.600 335.800 ;
        RECT 3.600 334.400 6.600 335.200 ;
        RECT 1.200 333.000 10.000 333.800 ;
        RECT 11.800 333.400 12.600 335.800 ;
        RECT 15.600 335.600 16.400 335.800 ;
        RECT 17.200 335.600 18.800 336.400 ;
        RECT 21.800 335.600 22.800 336.400 ;
        RECT 25.200 335.800 27.600 336.600 ;
        RECT 14.000 333.600 14.800 335.200 ;
        RECT 15.600 334.800 16.400 335.000 ;
        RECT 15.600 334.200 20.000 334.800 ;
        RECT 19.200 334.000 20.000 334.200 ;
        RECT 1.200 327.400 2.000 333.000 ;
        RECT 10.600 332.600 12.600 333.400 ;
        RECT 16.400 332.600 19.600 333.400 ;
        RECT 22.000 332.800 22.800 335.600 ;
        RECT 26.800 335.200 27.600 335.800 ;
        RECT 26.800 334.600 28.600 335.200 ;
        RECT 27.800 333.400 28.600 334.600 ;
        RECT 31.600 334.600 32.400 339.800 ;
        RECT 33.200 336.300 34.000 339.800 ;
        RECT 38.000 336.400 38.800 339.800 ;
        RECT 34.800 336.300 35.600 336.400 ;
        RECT 33.200 335.700 35.600 336.300 ;
        RECT 33.200 335.200 34.200 335.700 ;
        RECT 34.800 335.600 35.600 335.700 ;
        RECT 37.800 335.800 38.800 336.400 ;
        RECT 31.600 334.000 32.800 334.600 ;
        RECT 27.800 332.600 31.600 333.400 ;
        RECT 2.600 332.000 3.400 332.200 ;
        RECT 7.600 332.000 8.400 332.400 ;
        RECT 25.200 332.000 26.000 332.600 ;
        RECT 32.200 332.000 32.800 334.000 ;
        RECT 2.600 331.400 26.000 332.000 ;
        RECT 32.000 331.400 32.800 332.000 ;
        RECT 32.000 329.600 32.600 331.400 ;
        RECT 33.400 330.800 34.200 335.200 ;
        RECT 10.800 329.400 11.600 329.600 ;
        RECT 6.200 329.000 11.600 329.400 ;
        RECT 5.400 328.800 11.600 329.000 ;
        RECT 12.600 329.000 21.200 329.600 ;
        RECT 2.800 328.000 4.400 328.800 ;
        RECT 5.400 328.200 6.800 328.800 ;
        RECT 12.600 328.200 13.200 329.000 ;
        RECT 20.400 328.800 21.200 329.000 ;
        RECT 23.600 329.000 32.600 329.600 ;
        RECT 23.600 328.800 24.400 329.000 ;
        RECT 3.800 327.600 4.400 328.000 ;
        RECT 7.400 327.600 13.200 328.200 ;
        RECT 13.800 327.600 16.400 328.400 ;
        RECT 1.200 326.800 3.200 327.400 ;
        RECT 3.800 326.800 8.000 327.600 ;
        RECT 2.600 326.200 3.200 326.800 ;
        RECT 2.600 325.600 3.600 326.200 ;
        RECT 2.800 322.200 3.600 325.600 ;
        RECT 6.000 322.200 6.800 326.800 ;
        RECT 9.200 322.200 10.000 325.000 ;
        RECT 10.800 322.200 11.600 325.000 ;
        RECT 12.400 322.200 13.200 327.000 ;
        RECT 15.600 322.200 16.400 327.000 ;
        RECT 18.800 322.200 19.600 328.400 ;
        RECT 26.800 327.600 29.400 328.400 ;
        RECT 22.000 326.800 26.200 327.600 ;
        RECT 20.400 322.200 21.200 325.000 ;
        RECT 22.000 322.200 22.800 325.000 ;
        RECT 23.600 322.200 24.400 325.000 ;
        RECT 26.800 322.200 27.600 327.600 ;
        RECT 32.000 327.400 32.600 329.000 ;
        RECT 30.000 326.800 32.600 327.400 ;
        RECT 33.200 330.000 34.200 330.800 ;
        RECT 37.800 334.400 38.400 335.800 ;
        RECT 41.200 335.200 42.000 339.800 ;
        RECT 39.400 334.600 42.000 335.200 ;
        RECT 37.800 333.600 38.800 334.400 ;
        RECT 37.800 330.200 38.400 333.600 ;
        RECT 39.400 333.000 40.000 334.600 ;
        RECT 39.000 332.200 40.000 333.000 ;
        RECT 39.400 330.200 40.000 332.200 ;
        RECT 42.800 332.300 43.600 339.800 ;
        RECT 44.400 335.600 45.200 337.200 ;
        RECT 49.800 336.000 50.600 339.000 ;
        RECT 54.000 337.000 54.800 339.000 ;
        RECT 49.000 335.400 50.600 336.000 ;
        RECT 49.000 335.000 49.800 335.400 ;
        RECT 49.000 334.400 49.600 335.000 ;
        RECT 54.200 334.800 54.800 337.000 ;
        RECT 55.600 335.600 56.400 337.200 ;
        RECT 47.600 333.600 49.600 334.400 ;
        RECT 50.600 334.200 54.800 334.800 ;
        RECT 50.600 333.800 51.600 334.200 ;
        RECT 47.600 332.300 48.400 332.400 ;
        RECT 42.800 331.700 48.400 332.300 ;
        RECT 30.000 322.200 30.800 326.800 ;
        RECT 33.200 322.200 34.000 330.000 ;
        RECT 37.800 329.200 38.800 330.200 ;
        RECT 39.400 329.600 42.000 330.200 ;
        RECT 38.000 322.200 38.800 329.200 ;
        RECT 41.200 322.200 42.000 329.600 ;
        RECT 42.800 322.200 43.600 331.700 ;
        RECT 47.600 330.800 48.400 331.700 ;
        RECT 49.000 329.800 49.600 333.600 ;
        RECT 50.200 333.000 51.600 333.800 ;
        RECT 51.000 331.000 51.600 333.000 ;
        RECT 52.400 331.600 53.200 333.200 ;
        RECT 54.000 331.600 54.800 333.200 ;
        RECT 51.000 330.400 54.800 331.000 ;
        RECT 49.000 329.200 50.600 329.800 ;
        RECT 49.800 324.400 50.600 329.200 ;
        RECT 54.200 327.000 54.800 330.400 ;
        RECT 49.200 323.600 50.600 324.400 ;
        RECT 49.800 322.200 50.600 323.600 ;
        RECT 54.000 323.000 54.800 327.000 ;
        RECT 57.200 322.200 58.000 339.800 ;
        RECT 60.400 336.000 61.200 339.800 ;
        RECT 60.200 335.200 61.200 336.000 ;
        RECT 60.200 330.800 61.000 335.200 ;
        RECT 62.000 334.600 62.800 339.800 ;
        RECT 68.400 336.600 69.200 339.800 ;
        RECT 70.000 337.000 70.800 339.800 ;
        RECT 71.600 337.000 72.400 339.800 ;
        RECT 73.200 337.000 74.000 339.800 ;
        RECT 74.800 337.000 75.600 339.800 ;
        RECT 78.000 337.000 78.800 339.800 ;
        RECT 81.200 337.000 82.000 339.800 ;
        RECT 82.800 337.000 83.600 339.800 ;
        RECT 84.400 337.000 85.200 339.800 ;
        RECT 66.800 335.800 69.200 336.600 ;
        RECT 86.000 336.600 86.800 339.800 ;
        RECT 66.800 335.200 67.600 335.800 ;
        RECT 61.600 334.000 62.800 334.600 ;
        RECT 65.800 334.600 67.600 335.200 ;
        RECT 71.600 335.600 72.600 336.400 ;
        RECT 75.600 335.600 77.200 336.400 ;
        RECT 78.000 335.800 82.600 336.400 ;
        RECT 86.000 335.800 88.600 336.600 ;
        RECT 78.000 335.600 78.800 335.800 ;
        RECT 61.600 332.000 62.200 334.000 ;
        RECT 65.800 333.400 66.600 334.600 ;
        RECT 62.800 332.600 66.600 333.400 ;
        RECT 71.600 332.800 72.400 335.600 ;
        RECT 78.000 334.800 78.800 335.000 ;
        RECT 74.400 334.200 78.800 334.800 ;
        RECT 74.400 334.000 75.200 334.200 ;
        RECT 79.600 333.600 80.400 335.200 ;
        RECT 81.800 333.400 82.600 335.800 ;
        RECT 87.800 335.200 88.600 335.800 ;
        RECT 87.800 334.400 90.800 335.200 ;
        RECT 92.400 333.800 93.200 339.800 ;
        RECT 94.000 335.600 94.800 337.200 ;
        RECT 74.800 332.600 78.000 333.400 ;
        RECT 81.800 332.600 83.800 333.400 ;
        RECT 84.400 333.000 93.200 333.800 ;
        RECT 68.400 332.000 69.200 332.600 ;
        RECT 79.600 332.000 80.400 332.400 ;
        RECT 86.000 332.000 86.800 332.400 ;
        RECT 91.000 332.000 91.800 332.200 ;
        RECT 61.600 331.400 62.400 332.000 ;
        RECT 68.400 331.400 91.800 332.000 ;
        RECT 60.200 330.000 61.200 330.800 ;
        RECT 60.400 322.200 61.200 330.000 ;
        RECT 61.800 329.600 62.400 331.400 ;
        RECT 61.800 329.000 70.800 329.600 ;
        RECT 61.800 327.400 62.400 329.000 ;
        RECT 70.000 328.800 70.800 329.000 ;
        RECT 73.200 329.000 81.800 329.600 ;
        RECT 73.200 328.800 74.000 329.000 ;
        RECT 65.000 327.600 67.600 328.400 ;
        RECT 61.800 326.800 64.400 327.400 ;
        RECT 63.600 322.200 64.400 326.800 ;
        RECT 66.800 322.200 67.600 327.600 ;
        RECT 68.200 326.800 72.400 327.600 ;
        RECT 70.000 322.200 70.800 325.000 ;
        RECT 71.600 322.200 72.400 325.000 ;
        RECT 73.200 322.200 74.000 325.000 ;
        RECT 74.800 322.200 75.600 328.400 ;
        RECT 78.000 327.600 80.600 328.400 ;
        RECT 81.200 328.200 81.800 329.000 ;
        RECT 82.800 329.400 83.600 329.600 ;
        RECT 82.800 329.000 88.200 329.400 ;
        RECT 82.800 328.800 89.000 329.000 ;
        RECT 87.600 328.200 89.000 328.800 ;
        RECT 81.200 327.600 87.000 328.200 ;
        RECT 90.000 328.000 91.600 328.800 ;
        RECT 90.000 327.600 90.600 328.000 ;
        RECT 78.000 322.200 78.800 327.000 ;
        RECT 81.200 322.200 82.000 327.000 ;
        RECT 86.400 326.800 90.600 327.600 ;
        RECT 92.400 327.400 93.200 333.000 ;
        RECT 91.200 326.800 93.200 327.400 ;
        RECT 95.600 332.300 96.400 339.800 ;
        RECT 101.000 336.000 101.800 339.000 ;
        RECT 105.200 337.000 106.000 339.000 ;
        RECT 100.200 335.400 101.800 336.000 ;
        RECT 100.200 335.000 101.000 335.400 ;
        RECT 100.200 334.400 100.800 335.000 ;
        RECT 105.400 334.800 106.000 337.000 ;
        RECT 106.800 335.000 107.600 339.800 ;
        RECT 111.200 338.400 112.000 339.800 ;
        RECT 110.000 337.800 112.000 338.400 ;
        RECT 115.600 337.800 116.400 339.800 ;
        RECT 119.800 338.400 121.000 339.800 ;
        RECT 119.600 337.800 121.000 338.400 ;
        RECT 110.000 337.000 110.800 337.800 ;
        RECT 115.600 337.200 116.200 337.800 ;
        RECT 111.600 336.400 112.400 337.200 ;
        RECT 113.400 336.600 116.200 337.200 ;
        RECT 119.600 337.000 120.400 337.800 ;
        RECT 113.400 336.400 114.200 336.600 ;
        RECT 97.200 334.300 98.000 334.400 ;
        RECT 98.800 334.300 100.800 334.400 ;
        RECT 97.200 333.700 100.800 334.300 ;
        RECT 101.800 334.200 106.000 334.800 ;
        RECT 107.600 334.200 109.200 334.400 ;
        RECT 111.800 334.200 112.400 336.400 ;
        RECT 121.400 335.400 122.200 335.600 ;
        RECT 124.400 335.400 125.200 339.800 ;
        RECT 121.400 334.800 125.200 335.400 ;
        RECT 126.000 335.000 126.800 339.800 ;
        RECT 130.400 338.400 131.200 339.800 ;
        RECT 129.200 337.800 131.200 338.400 ;
        RECT 134.800 337.800 135.600 339.800 ;
        RECT 139.000 338.400 140.200 339.800 ;
        RECT 138.800 337.800 140.200 338.400 ;
        RECT 129.200 337.000 130.000 337.800 ;
        RECT 134.800 337.200 135.400 337.800 ;
        RECT 130.800 336.400 131.600 337.200 ;
        RECT 132.600 336.600 135.400 337.200 ;
        RECT 138.800 337.000 139.600 337.800 ;
        RECT 132.600 336.400 133.400 336.600 ;
        RECT 117.400 334.200 118.200 334.400 ;
        RECT 101.800 333.800 102.800 334.200 ;
        RECT 97.200 333.600 98.000 333.700 ;
        RECT 98.800 333.600 100.800 333.700 ;
        RECT 98.800 332.300 99.600 332.400 ;
        RECT 95.600 331.700 99.600 332.300 ;
        RECT 82.800 322.200 83.600 325.000 ;
        RECT 84.400 322.200 85.200 325.000 ;
        RECT 87.600 322.200 88.400 326.800 ;
        RECT 91.200 326.200 91.800 326.800 ;
        RECT 90.800 325.600 91.800 326.200 ;
        RECT 90.800 322.200 91.600 325.600 ;
        RECT 95.600 322.200 96.400 331.700 ;
        RECT 98.800 330.800 99.600 331.700 ;
        RECT 100.200 329.800 100.800 333.600 ;
        RECT 101.400 333.000 102.800 333.800 ;
        RECT 107.600 333.600 118.600 334.200 ;
        RECT 110.600 333.400 111.400 333.600 ;
        RECT 102.200 331.000 102.800 333.000 ;
        RECT 103.600 331.600 104.400 333.200 ;
        RECT 105.200 331.600 106.000 333.200 ;
        RECT 109.000 332.400 109.800 332.600 ;
        RECT 109.000 332.300 114.000 332.400 ;
        RECT 116.400 332.300 117.200 332.400 ;
        RECT 109.000 331.800 117.200 332.300 ;
        RECT 113.200 331.700 117.200 331.800 ;
        RECT 113.200 331.600 114.000 331.700 ;
        RECT 116.400 331.600 117.200 331.700 ;
        RECT 106.800 331.000 112.400 331.200 ;
        RECT 102.200 330.400 106.000 331.000 ;
        RECT 100.200 329.200 101.800 329.800 ;
        RECT 101.000 322.200 101.800 329.200 ;
        RECT 105.400 327.000 106.000 330.400 ;
        RECT 105.200 323.000 106.000 327.000 ;
        RECT 106.800 330.800 112.600 331.000 ;
        RECT 106.800 330.600 116.600 330.800 ;
        RECT 106.800 322.200 107.600 330.600 ;
        RECT 111.800 330.200 116.600 330.600 ;
        RECT 110.000 329.000 115.400 329.600 ;
        RECT 110.000 328.800 110.800 329.000 ;
        RECT 114.600 328.800 115.400 329.000 ;
        RECT 116.000 329.000 116.600 330.200 ;
        RECT 118.000 330.400 118.600 333.600 ;
        RECT 119.600 332.800 120.400 333.000 ;
        RECT 119.600 332.200 123.400 332.800 ;
        RECT 122.600 332.000 123.400 332.200 ;
        RECT 121.000 331.400 121.800 331.600 ;
        RECT 124.400 331.400 125.200 334.800 ;
        RECT 126.800 334.200 128.400 334.400 ;
        RECT 131.000 334.200 131.600 336.400 ;
        RECT 140.600 335.400 141.400 335.600 ;
        RECT 143.600 335.400 144.400 339.800 ;
        RECT 140.600 334.800 144.400 335.400 ;
        RECT 134.000 334.200 134.800 334.400 ;
        RECT 136.600 334.200 137.400 334.400 ;
        RECT 126.800 333.600 137.800 334.200 ;
        RECT 129.800 333.400 130.600 333.600 ;
        RECT 128.200 332.400 129.000 332.600 ;
        RECT 130.800 332.400 131.600 332.600 ;
        RECT 128.200 331.800 133.200 332.400 ;
        RECT 132.400 331.600 133.200 331.800 ;
        RECT 121.000 330.800 125.200 331.400 ;
        RECT 118.000 329.800 120.400 330.400 ;
        RECT 117.400 329.000 118.200 329.200 ;
        RECT 116.000 328.400 118.200 329.000 ;
        RECT 119.800 328.800 120.400 329.800 ;
        RECT 119.800 328.000 121.200 328.800 ;
        RECT 113.400 327.400 114.200 327.600 ;
        RECT 116.200 327.400 117.000 327.600 ;
        RECT 110.000 326.200 110.800 327.000 ;
        RECT 113.400 326.800 117.000 327.400 ;
        RECT 115.600 326.200 116.200 326.800 ;
        RECT 119.600 326.200 120.400 327.000 ;
        RECT 110.000 325.600 112.000 326.200 ;
        RECT 111.200 322.200 112.000 325.600 ;
        RECT 115.600 322.200 116.400 326.200 ;
        RECT 119.800 322.200 121.000 326.200 ;
        RECT 124.400 322.200 125.200 330.800 ;
        RECT 126.000 331.000 131.600 331.200 ;
        RECT 126.000 330.800 131.800 331.000 ;
        RECT 126.000 330.600 135.800 330.800 ;
        RECT 126.000 322.200 126.800 330.600 ;
        RECT 131.000 330.200 135.800 330.600 ;
        RECT 129.200 329.000 134.600 329.600 ;
        RECT 129.200 328.800 130.000 329.000 ;
        RECT 133.800 328.800 134.600 329.000 ;
        RECT 135.200 329.000 135.800 330.200 ;
        RECT 137.200 330.400 137.800 333.600 ;
        RECT 138.800 332.800 139.600 333.000 ;
        RECT 138.800 332.200 142.600 332.800 ;
        RECT 141.800 332.000 142.600 332.200 ;
        RECT 140.200 331.400 141.000 331.600 ;
        RECT 143.600 331.400 144.400 334.800 ;
        RECT 140.200 330.800 144.400 331.400 ;
        RECT 137.200 329.800 139.600 330.400 ;
        RECT 136.600 329.000 137.400 329.200 ;
        RECT 135.200 328.400 137.400 329.000 ;
        RECT 139.000 328.800 139.600 329.800 ;
        RECT 139.000 328.000 140.400 328.800 ;
        RECT 132.600 327.400 133.400 327.600 ;
        RECT 135.400 327.400 136.200 327.600 ;
        RECT 129.200 326.200 130.000 327.000 ;
        RECT 132.600 326.800 136.200 327.400 ;
        RECT 134.800 326.200 135.400 326.800 ;
        RECT 138.800 326.200 139.600 327.000 ;
        RECT 129.200 325.600 131.200 326.200 ;
        RECT 130.400 322.200 131.200 325.600 ;
        RECT 134.800 322.200 135.600 326.200 ;
        RECT 139.000 322.200 140.200 326.200 ;
        RECT 143.600 322.200 144.400 330.800 ;
        RECT 145.200 322.200 146.000 339.800 ;
        RECT 146.800 336.300 147.600 337.200 ;
        RECT 154.800 336.300 155.600 339.800 ;
        RECT 146.800 335.700 155.600 336.300 ;
        RECT 146.800 335.600 147.600 335.700 ;
        RECT 154.600 335.200 155.600 335.700 ;
        RECT 154.600 330.800 155.400 335.200 ;
        RECT 156.400 334.600 157.200 339.800 ;
        RECT 162.800 336.600 163.600 339.800 ;
        RECT 164.400 337.000 165.200 339.800 ;
        RECT 166.000 337.000 166.800 339.800 ;
        RECT 167.600 337.000 168.400 339.800 ;
        RECT 169.200 337.000 170.000 339.800 ;
        RECT 172.400 337.000 173.200 339.800 ;
        RECT 175.600 337.000 176.400 339.800 ;
        RECT 177.200 337.000 178.000 339.800 ;
        RECT 178.800 337.000 179.600 339.800 ;
        RECT 161.200 335.800 163.600 336.600 ;
        RECT 180.400 336.600 181.200 339.800 ;
        RECT 161.200 335.200 162.000 335.800 ;
        RECT 156.000 334.000 157.200 334.600 ;
        RECT 160.200 334.600 162.000 335.200 ;
        RECT 166.000 335.600 167.000 336.400 ;
        RECT 170.000 335.600 171.600 336.400 ;
        RECT 172.400 335.800 177.000 336.400 ;
        RECT 180.400 335.800 183.000 336.600 ;
        RECT 172.400 335.600 173.200 335.800 ;
        RECT 156.000 332.000 156.600 334.000 ;
        RECT 160.200 333.400 161.000 334.600 ;
        RECT 157.200 332.600 161.000 333.400 ;
        RECT 166.000 332.800 166.800 335.600 ;
        RECT 172.400 334.800 173.200 335.000 ;
        RECT 168.800 334.200 173.200 334.800 ;
        RECT 168.800 334.000 169.600 334.200 ;
        RECT 174.000 333.600 174.800 335.200 ;
        RECT 176.200 333.400 177.000 335.800 ;
        RECT 182.200 335.200 183.000 335.800 ;
        RECT 182.200 334.400 185.200 335.200 ;
        RECT 186.800 333.800 187.600 339.800 ;
        RECT 188.400 335.200 189.200 339.800 ;
        RECT 191.600 336.400 192.400 339.800 ;
        RECT 191.600 335.800 192.600 336.400 ;
        RECT 188.400 334.600 191.000 335.200 ;
        RECT 169.200 332.600 172.400 333.400 ;
        RECT 176.200 332.600 178.200 333.400 ;
        RECT 178.800 333.000 187.600 333.800 ;
        RECT 162.800 332.000 163.600 332.600 ;
        RECT 180.400 332.000 181.200 332.400 ;
        RECT 183.600 332.000 184.400 332.400 ;
        RECT 185.400 332.000 186.200 332.200 ;
        RECT 156.000 331.400 156.800 332.000 ;
        RECT 162.800 331.400 186.200 332.000 ;
        RECT 154.600 330.000 155.600 330.800 ;
        RECT 154.800 322.200 155.600 330.000 ;
        RECT 156.200 329.600 156.800 331.400 ;
        RECT 156.200 329.000 165.200 329.600 ;
        RECT 156.200 327.400 156.800 329.000 ;
        RECT 164.400 328.800 165.200 329.000 ;
        RECT 167.600 329.000 176.200 329.600 ;
        RECT 167.600 328.800 168.400 329.000 ;
        RECT 159.400 327.600 162.000 328.400 ;
        RECT 156.200 326.800 158.800 327.400 ;
        RECT 158.000 322.200 158.800 326.800 ;
        RECT 161.200 322.200 162.000 327.600 ;
        RECT 162.600 326.800 166.800 327.600 ;
        RECT 164.400 322.200 165.200 325.000 ;
        RECT 166.000 322.200 166.800 325.000 ;
        RECT 167.600 322.200 168.400 325.000 ;
        RECT 169.200 322.200 170.000 328.400 ;
        RECT 172.400 327.600 175.000 328.400 ;
        RECT 175.600 328.200 176.200 329.000 ;
        RECT 177.200 329.400 178.000 329.600 ;
        RECT 177.200 329.000 182.600 329.400 ;
        RECT 177.200 328.800 183.400 329.000 ;
        RECT 182.000 328.200 183.400 328.800 ;
        RECT 175.600 327.600 181.400 328.200 ;
        RECT 184.400 328.000 186.000 328.800 ;
        RECT 184.400 327.600 185.000 328.000 ;
        RECT 172.400 322.200 173.200 327.000 ;
        RECT 175.600 322.200 176.400 327.000 ;
        RECT 180.800 326.800 185.000 327.600 ;
        RECT 186.800 327.400 187.600 333.000 ;
        RECT 188.600 332.400 189.400 333.200 ;
        RECT 188.400 331.600 189.400 332.400 ;
        RECT 190.400 333.000 191.000 334.600 ;
        RECT 192.000 334.400 192.600 335.800 ;
        RECT 191.600 333.600 192.600 334.400 ;
        RECT 190.400 332.200 191.400 333.000 ;
        RECT 190.400 330.200 191.000 332.200 ;
        RECT 192.000 330.200 192.600 333.600 ;
        RECT 185.600 326.800 187.600 327.400 ;
        RECT 188.400 329.600 191.000 330.200 ;
        RECT 177.200 322.200 178.000 325.000 ;
        RECT 178.800 322.200 179.600 325.000 ;
        RECT 182.000 322.200 182.800 326.800 ;
        RECT 185.600 326.200 186.200 326.800 ;
        RECT 185.200 325.600 186.200 326.200 ;
        RECT 185.200 322.200 186.000 325.600 ;
        RECT 188.400 322.200 189.200 329.600 ;
        RECT 191.600 329.200 192.600 330.200 ;
        RECT 194.800 333.800 195.600 339.800 ;
        RECT 201.200 336.600 202.000 339.800 ;
        RECT 202.800 337.000 203.600 339.800 ;
        RECT 204.400 337.000 205.200 339.800 ;
        RECT 206.000 337.000 206.800 339.800 ;
        RECT 209.200 337.000 210.000 339.800 ;
        RECT 212.400 337.000 213.200 339.800 ;
        RECT 214.000 337.000 214.800 339.800 ;
        RECT 215.600 337.000 216.400 339.800 ;
        RECT 217.200 337.000 218.000 339.800 ;
        RECT 199.400 335.800 202.000 336.600 ;
        RECT 218.800 336.600 219.600 339.800 ;
        RECT 205.400 335.800 210.000 336.400 ;
        RECT 199.400 335.200 200.200 335.800 ;
        RECT 197.200 334.400 200.200 335.200 ;
        RECT 194.800 333.000 203.600 333.800 ;
        RECT 205.400 333.400 206.200 335.800 ;
        RECT 209.200 335.600 210.000 335.800 ;
        RECT 210.800 335.600 212.400 336.400 ;
        RECT 215.400 335.600 216.400 336.400 ;
        RECT 218.800 335.800 221.200 336.600 ;
        RECT 207.600 333.600 208.400 335.200 ;
        RECT 209.200 334.800 210.000 335.000 ;
        RECT 209.200 334.200 213.600 334.800 ;
        RECT 212.800 334.000 213.600 334.200 ;
        RECT 191.600 322.200 192.400 329.200 ;
        RECT 194.800 327.400 195.600 333.000 ;
        RECT 204.200 332.600 206.200 333.400 ;
        RECT 210.000 332.600 213.200 333.400 ;
        RECT 215.600 332.800 216.400 335.600 ;
        RECT 220.400 335.200 221.200 335.800 ;
        RECT 220.400 334.600 222.200 335.200 ;
        RECT 221.400 333.400 222.200 334.600 ;
        RECT 225.200 334.600 226.000 339.800 ;
        RECT 226.800 336.000 227.600 339.800 ;
        RECT 226.800 335.200 227.800 336.000 ;
        RECT 225.200 334.000 226.400 334.600 ;
        RECT 221.400 332.600 225.200 333.400 ;
        RECT 196.200 332.000 197.000 332.200 ;
        RECT 201.200 332.000 202.000 332.400 ;
        RECT 218.800 332.000 219.600 332.600 ;
        RECT 225.800 332.000 226.400 334.000 ;
        RECT 196.200 331.400 219.600 332.000 ;
        RECT 225.600 331.400 226.400 332.000 ;
        RECT 225.600 329.600 226.200 331.400 ;
        RECT 227.000 330.800 227.800 335.200 ;
        RECT 231.600 335.200 232.400 339.800 ;
        RECT 234.800 335.200 235.600 339.800 ;
        RECT 238.000 335.600 238.800 337.200 ;
        RECT 231.600 334.400 235.600 335.200 ;
        RECT 234.800 331.600 235.600 334.400 ;
        RECT 204.400 329.400 205.200 329.600 ;
        RECT 199.800 329.000 205.200 329.400 ;
        RECT 199.000 328.800 205.200 329.000 ;
        RECT 206.200 329.000 214.800 329.600 ;
        RECT 196.400 328.000 198.000 328.800 ;
        RECT 199.000 328.200 200.400 328.800 ;
        RECT 206.200 328.200 206.800 329.000 ;
        RECT 214.000 328.800 214.800 329.000 ;
        RECT 217.200 329.000 226.200 329.600 ;
        RECT 217.200 328.800 218.000 329.000 ;
        RECT 197.400 327.600 198.000 328.000 ;
        RECT 201.000 327.600 206.800 328.200 ;
        RECT 207.400 327.600 210.000 328.400 ;
        RECT 194.800 326.800 196.800 327.400 ;
        RECT 197.400 326.800 201.600 327.600 ;
        RECT 196.200 326.200 196.800 326.800 ;
        RECT 196.200 325.600 197.200 326.200 ;
        RECT 196.400 322.200 197.200 325.600 ;
        RECT 199.600 322.200 200.400 326.800 ;
        RECT 202.800 322.200 203.600 325.000 ;
        RECT 204.400 322.200 205.200 325.000 ;
        RECT 206.000 322.200 206.800 327.000 ;
        RECT 209.200 322.200 210.000 327.000 ;
        RECT 212.400 322.200 213.200 328.400 ;
        RECT 220.400 327.600 223.000 328.400 ;
        RECT 215.600 326.800 219.800 327.600 ;
        RECT 214.000 322.200 214.800 325.000 ;
        RECT 215.600 322.200 216.400 325.000 ;
        RECT 217.200 322.200 218.000 325.000 ;
        RECT 220.400 322.200 221.200 327.600 ;
        RECT 225.600 327.400 226.200 329.000 ;
        RECT 223.600 326.800 226.200 327.400 ;
        RECT 226.800 330.000 227.800 330.800 ;
        RECT 231.600 330.800 235.600 331.600 ;
        RECT 223.600 322.200 224.400 326.800 ;
        RECT 226.800 322.200 227.600 330.000 ;
        RECT 231.600 322.200 232.400 330.800 ;
        RECT 234.800 322.200 235.600 330.800 ;
        RECT 239.600 322.200 240.400 339.800 ;
        RECT 241.200 333.800 242.000 339.800 ;
        RECT 247.600 336.600 248.400 339.800 ;
        RECT 249.200 337.000 250.000 339.800 ;
        RECT 250.800 337.000 251.600 339.800 ;
        RECT 252.400 337.000 253.200 339.800 ;
        RECT 255.600 337.000 256.400 339.800 ;
        RECT 258.800 337.000 259.600 339.800 ;
        RECT 260.400 337.000 261.200 339.800 ;
        RECT 262.000 337.000 262.800 339.800 ;
        RECT 263.600 337.000 264.400 339.800 ;
        RECT 245.800 335.800 248.400 336.600 ;
        RECT 265.200 336.600 266.000 339.800 ;
        RECT 251.800 335.800 256.400 336.400 ;
        RECT 245.800 335.200 246.600 335.800 ;
        RECT 243.600 334.400 246.600 335.200 ;
        RECT 241.200 333.000 250.000 333.800 ;
        RECT 251.800 333.400 252.600 335.800 ;
        RECT 255.600 335.600 256.400 335.800 ;
        RECT 257.200 335.600 258.800 336.400 ;
        RECT 261.800 335.600 262.800 336.400 ;
        RECT 265.200 335.800 267.600 336.600 ;
        RECT 254.000 333.600 254.800 335.200 ;
        RECT 255.600 334.800 256.400 335.000 ;
        RECT 255.600 334.200 260.000 334.800 ;
        RECT 259.200 334.000 260.000 334.200 ;
        RECT 241.200 327.400 242.000 333.000 ;
        RECT 250.600 332.600 252.600 333.400 ;
        RECT 256.400 332.600 259.600 333.400 ;
        RECT 262.000 332.800 262.800 335.600 ;
        RECT 266.800 335.200 267.600 335.800 ;
        RECT 266.800 334.600 268.600 335.200 ;
        RECT 267.800 333.400 268.600 334.600 ;
        RECT 271.600 334.600 272.400 339.800 ;
        RECT 273.200 336.000 274.000 339.800 ;
        RECT 273.200 335.200 274.200 336.000 ;
        RECT 271.600 334.000 272.800 334.600 ;
        RECT 267.800 332.600 271.600 333.400 ;
        RECT 242.600 332.000 243.400 332.200 ;
        RECT 247.600 332.000 248.400 332.400 ;
        RECT 254.000 332.000 254.800 332.400 ;
        RECT 265.200 332.000 266.000 332.600 ;
        RECT 272.200 332.000 272.800 334.000 ;
        RECT 242.600 331.400 266.000 332.000 ;
        RECT 272.000 331.400 272.800 332.000 ;
        RECT 272.000 329.600 272.600 331.400 ;
        RECT 273.400 330.800 274.200 335.200 ;
        RECT 250.800 329.400 251.600 329.600 ;
        RECT 246.200 329.000 251.600 329.400 ;
        RECT 245.400 328.800 251.600 329.000 ;
        RECT 252.600 329.000 261.200 329.600 ;
        RECT 242.800 328.000 244.400 328.800 ;
        RECT 245.400 328.200 246.800 328.800 ;
        RECT 252.600 328.200 253.200 329.000 ;
        RECT 260.400 328.800 261.200 329.000 ;
        RECT 263.600 329.000 272.600 329.600 ;
        RECT 263.600 328.800 264.400 329.000 ;
        RECT 243.800 327.600 244.400 328.000 ;
        RECT 247.400 327.600 253.200 328.200 ;
        RECT 253.800 327.600 256.400 328.400 ;
        RECT 241.200 326.800 243.200 327.400 ;
        RECT 243.800 326.800 248.000 327.600 ;
        RECT 242.600 326.200 243.200 326.800 ;
        RECT 242.600 325.600 243.600 326.200 ;
        RECT 242.800 322.200 243.600 325.600 ;
        RECT 246.000 322.200 246.800 326.800 ;
        RECT 249.200 322.200 250.000 325.000 ;
        RECT 250.800 322.200 251.600 325.000 ;
        RECT 252.400 322.200 253.200 327.000 ;
        RECT 255.600 322.200 256.400 327.000 ;
        RECT 258.800 322.200 259.600 328.400 ;
        RECT 266.800 327.600 269.400 328.400 ;
        RECT 262.000 326.800 266.200 327.600 ;
        RECT 260.400 322.200 261.200 325.000 ;
        RECT 262.000 322.200 262.800 325.000 ;
        RECT 263.600 322.200 264.400 325.000 ;
        RECT 266.800 322.200 267.600 327.600 ;
        RECT 272.000 327.400 272.600 329.000 ;
        RECT 270.000 326.800 272.600 327.400 ;
        RECT 273.200 330.000 274.200 330.800 ;
        RECT 270.000 322.200 270.800 326.800 ;
        RECT 273.200 322.200 274.000 330.000 ;
        RECT 276.400 322.200 277.200 339.800 ;
        RECT 278.000 335.600 278.800 337.200 ;
        RECT 280.800 334.200 281.600 339.800 ;
        RECT 287.200 334.200 288.000 339.800 ;
        RECT 293.600 334.200 294.400 339.800 ;
        RECT 300.000 334.200 300.800 339.800 ;
        RECT 311.600 336.400 312.400 339.800 ;
        RECT 311.400 335.800 312.400 336.400 ;
        RECT 311.400 334.400 312.000 335.800 ;
        RECT 314.800 335.200 315.600 339.800 ;
        RECT 319.000 336.400 319.800 339.800 ;
        RECT 318.000 335.800 319.800 336.400 ;
        RECT 321.200 336.000 322.000 339.800 ;
        RECT 324.400 339.200 328.400 339.800 ;
        RECT 324.400 336.000 325.200 339.200 ;
        RECT 321.200 335.800 325.200 336.000 ;
        RECT 313.000 334.600 315.600 335.200 ;
        RECT 279.800 333.800 281.600 334.200 ;
        RECT 286.200 333.800 288.000 334.200 ;
        RECT 292.600 333.800 294.400 334.200 ;
        RECT 299.000 333.800 300.800 334.200 ;
        RECT 305.200 334.300 306.000 334.400 ;
        RECT 311.400 334.300 312.400 334.400 ;
        RECT 279.800 333.600 281.400 333.800 ;
        RECT 286.200 333.600 287.800 333.800 ;
        RECT 292.600 333.600 294.200 333.800 ;
        RECT 299.000 333.600 300.600 333.800 ;
        RECT 305.200 333.700 312.400 334.300 ;
        RECT 305.200 333.600 306.000 333.700 ;
        RECT 311.400 333.600 312.400 333.700 ;
        RECT 279.800 330.400 280.400 333.600 ;
        RECT 279.600 329.600 280.400 330.400 ;
        RECT 284.400 329.600 285.200 331.200 ;
        RECT 286.200 330.400 286.800 333.600 ;
        RECT 286.000 329.600 286.800 330.400 ;
        RECT 290.800 329.600 291.600 331.200 ;
        RECT 292.600 330.400 293.200 333.600 ;
        RECT 292.400 329.600 293.200 330.400 ;
        RECT 297.200 329.600 298.000 331.200 ;
        RECT 299.000 330.400 299.600 333.600 ;
        RECT 298.800 329.600 299.600 330.400 ;
        RECT 303.600 330.300 304.400 331.200 ;
        RECT 305.200 330.300 306.000 330.400 ;
        RECT 303.600 329.700 306.000 330.300 ;
        RECT 303.600 329.600 304.400 329.700 ;
        RECT 305.200 329.600 306.000 329.700 ;
        RECT 311.400 330.200 312.000 333.600 ;
        RECT 313.000 333.000 313.600 334.600 ;
        RECT 316.400 333.600 317.200 335.200 ;
        RECT 312.600 332.200 313.600 333.000 ;
        RECT 313.000 330.200 313.600 332.200 ;
        RECT 314.600 332.400 315.400 333.200 ;
        RECT 314.600 331.600 315.600 332.400 ;
        RECT 318.000 332.300 318.800 335.800 ;
        RECT 321.400 335.400 325.000 335.800 ;
        RECT 326.000 335.600 326.800 338.600 ;
        RECT 327.600 335.800 328.400 339.200 ;
        RECT 329.200 335.800 330.000 339.800 ;
        RECT 330.800 336.000 331.600 339.800 ;
        RECT 334.000 336.000 334.800 339.800 ;
        RECT 337.200 336.000 338.000 339.800 ;
        RECT 330.800 335.800 334.800 336.000 ;
        RECT 322.000 334.400 322.800 334.800 ;
        RECT 326.200 334.400 326.800 335.600 ;
        RECT 329.400 334.400 330.000 335.800 ;
        RECT 331.000 335.400 334.600 335.800 ;
        RECT 337.000 335.200 338.000 336.000 ;
        RECT 333.200 334.400 334.000 334.800 ;
        RECT 321.200 333.800 322.800 334.400 ;
        RECT 324.400 333.800 326.800 334.400 ;
        RECT 321.200 333.600 322.000 333.800 ;
        RECT 324.400 333.600 325.200 333.800 ;
        RECT 322.800 332.300 323.600 333.200 ;
        RECT 318.000 331.700 323.600 332.300 ;
        RECT 279.800 327.000 280.400 329.600 ;
        RECT 281.200 327.600 282.000 329.200 ;
        RECT 286.200 327.000 286.800 329.600 ;
        RECT 287.600 327.600 288.400 329.200 ;
        RECT 292.600 327.000 293.200 329.600 ;
        RECT 294.000 327.600 294.800 329.200 ;
        RECT 299.000 327.000 299.600 329.600 ;
        RECT 311.400 329.200 312.400 330.200 ;
        RECT 313.000 329.600 315.600 330.200 ;
        RECT 300.400 327.600 301.200 329.200 ;
        RECT 279.800 326.400 283.400 327.000 ;
        RECT 279.800 326.200 280.400 326.400 ;
        RECT 279.600 322.200 280.400 326.200 ;
        RECT 282.800 326.200 283.400 326.400 ;
        RECT 286.200 326.400 289.800 327.000 ;
        RECT 286.200 326.200 286.800 326.400 ;
        RECT 282.800 322.200 283.600 326.200 ;
        RECT 286.000 322.200 286.800 326.200 ;
        RECT 289.200 326.200 289.800 326.400 ;
        RECT 292.600 326.400 296.200 327.000 ;
        RECT 292.600 326.200 293.200 326.400 ;
        RECT 289.200 322.200 290.000 326.200 ;
        RECT 292.400 322.200 293.200 326.200 ;
        RECT 295.600 326.200 296.200 326.400 ;
        RECT 299.000 326.400 302.600 327.000 ;
        RECT 299.000 326.200 299.600 326.400 ;
        RECT 295.600 322.200 296.400 326.200 ;
        RECT 298.800 322.200 299.600 326.200 ;
        RECT 302.000 326.200 302.600 326.400 ;
        RECT 302.000 322.200 302.800 326.200 ;
        RECT 311.600 322.200 312.400 329.200 ;
        RECT 314.800 322.200 315.600 329.600 ;
        RECT 318.000 322.200 318.800 331.700 ;
        RECT 322.800 331.600 323.600 331.700 ;
        RECT 324.400 330.200 325.000 333.600 ;
        RECT 326.000 331.600 326.800 333.200 ;
        RECT 327.600 332.800 328.400 334.400 ;
        RECT 329.200 333.600 331.800 334.400 ;
        RECT 333.200 333.800 334.800 334.400 ;
        RECT 334.000 333.600 334.800 333.800 ;
        RECT 329.200 330.200 330.000 330.400 ;
        RECT 331.200 330.200 331.800 333.600 ;
        RECT 332.400 331.600 333.200 333.200 ;
        RECT 337.000 330.800 337.800 335.200 ;
        RECT 338.800 334.600 339.600 339.800 ;
        RECT 345.200 336.600 346.000 339.800 ;
        RECT 346.800 337.000 347.600 339.800 ;
        RECT 348.400 337.000 349.200 339.800 ;
        RECT 350.000 337.000 350.800 339.800 ;
        RECT 351.600 337.000 352.400 339.800 ;
        RECT 354.800 337.000 355.600 339.800 ;
        RECT 358.000 337.000 358.800 339.800 ;
        RECT 359.600 337.000 360.400 339.800 ;
        RECT 361.200 337.000 362.000 339.800 ;
        RECT 343.600 335.800 346.000 336.600 ;
        RECT 362.800 336.600 363.600 339.800 ;
        RECT 343.600 335.200 344.400 335.800 ;
        RECT 338.400 334.000 339.600 334.600 ;
        RECT 342.600 334.600 344.400 335.200 ;
        RECT 348.400 335.600 349.400 336.400 ;
        RECT 352.400 335.600 354.000 336.400 ;
        RECT 354.800 335.800 359.400 336.400 ;
        RECT 362.800 335.800 365.400 336.600 ;
        RECT 354.800 335.600 355.600 335.800 ;
        RECT 338.400 332.000 339.000 334.000 ;
        RECT 342.600 333.400 343.400 334.600 ;
        RECT 339.600 332.600 343.400 333.400 ;
        RECT 348.400 332.800 349.200 335.600 ;
        RECT 354.800 334.800 355.600 335.000 ;
        RECT 351.200 334.200 355.600 334.800 ;
        RECT 351.200 334.000 352.000 334.200 ;
        RECT 356.400 333.600 357.200 335.200 ;
        RECT 358.600 333.400 359.400 335.800 ;
        RECT 364.600 335.200 365.400 335.800 ;
        RECT 364.600 334.400 367.600 335.200 ;
        RECT 369.200 333.800 370.000 339.800 ;
        RECT 370.800 335.800 371.600 339.800 ;
        RECT 372.400 336.000 373.200 339.800 ;
        RECT 375.600 336.000 376.400 339.800 ;
        RECT 372.400 335.800 376.400 336.000 ;
        RECT 377.200 339.200 381.200 339.800 ;
        RECT 377.200 335.800 378.000 339.200 ;
        RECT 378.800 335.800 379.600 338.600 ;
        RECT 380.400 336.000 381.200 339.200 ;
        RECT 383.600 336.000 384.400 339.800 ;
        RECT 380.400 335.800 384.400 336.000 ;
        RECT 385.800 336.400 386.600 339.800 ;
        RECT 391.600 336.400 392.400 339.800 ;
        RECT 385.800 335.800 387.600 336.400 ;
        RECT 371.000 334.400 371.600 335.800 ;
        RECT 372.600 335.400 376.200 335.800 ;
        RECT 374.800 334.400 375.600 334.800 ;
        RECT 378.800 334.400 379.400 335.800 ;
        RECT 380.600 335.400 384.200 335.800 ;
        RECT 382.800 334.400 383.600 334.800 ;
        RECT 351.600 332.600 354.800 333.400 ;
        RECT 358.600 332.600 360.600 333.400 ;
        RECT 361.200 333.000 370.000 333.800 ;
        RECT 370.800 333.600 373.400 334.400 ;
        RECT 374.800 333.800 376.400 334.400 ;
        RECT 375.600 333.600 376.400 333.800 ;
        RECT 345.200 332.000 346.000 332.600 ;
        RECT 362.800 332.000 363.600 332.400 ;
        RECT 367.800 332.000 368.600 332.200 ;
        RECT 338.400 331.400 339.200 332.000 ;
        RECT 345.200 331.400 368.600 332.000 ;
        RECT 323.800 322.200 325.800 330.200 ;
        RECT 329.200 329.600 330.600 330.200 ;
        RECT 331.200 329.600 332.200 330.200 ;
        RECT 337.000 330.000 338.000 330.800 ;
        RECT 330.000 328.400 330.600 329.600 ;
        RECT 330.000 327.600 330.800 328.400 ;
        RECT 331.400 322.200 332.200 329.600 ;
        RECT 337.200 322.200 338.000 330.000 ;
        RECT 338.600 329.600 339.200 331.400 ;
        RECT 338.600 329.000 347.600 329.600 ;
        RECT 338.600 327.400 339.200 329.000 ;
        RECT 346.800 328.800 347.600 329.000 ;
        RECT 350.000 329.000 358.600 329.600 ;
        RECT 350.000 328.800 350.800 329.000 ;
        RECT 341.800 327.600 344.400 328.400 ;
        RECT 338.600 326.800 341.200 327.400 ;
        RECT 340.400 322.200 341.200 326.800 ;
        RECT 343.600 322.200 344.400 327.600 ;
        RECT 345.000 326.800 349.200 327.600 ;
        RECT 346.800 322.200 347.600 325.000 ;
        RECT 348.400 322.200 349.200 325.000 ;
        RECT 350.000 322.200 350.800 325.000 ;
        RECT 351.600 322.200 352.400 328.400 ;
        RECT 354.800 327.600 357.400 328.400 ;
        RECT 358.000 328.200 358.600 329.000 ;
        RECT 359.600 329.400 360.400 329.600 ;
        RECT 359.600 329.000 365.000 329.400 ;
        RECT 359.600 328.800 365.800 329.000 ;
        RECT 364.400 328.200 365.800 328.800 ;
        RECT 358.000 327.600 363.800 328.200 ;
        RECT 366.800 328.000 368.400 328.800 ;
        RECT 366.800 327.600 367.400 328.000 ;
        RECT 354.800 322.200 355.600 327.000 ;
        RECT 358.000 322.200 358.800 327.000 ;
        RECT 363.200 326.800 367.400 327.600 ;
        RECT 369.200 327.400 370.000 333.000 ;
        RECT 370.800 330.200 371.600 330.400 ;
        RECT 372.800 330.200 373.400 333.600 ;
        RECT 374.000 331.600 374.800 333.200 ;
        RECT 377.200 332.800 378.000 334.400 ;
        RECT 378.800 333.800 381.200 334.400 ;
        RECT 382.800 333.800 384.400 334.400 ;
        RECT 380.400 333.600 381.200 333.800 ;
        RECT 383.600 333.600 384.400 333.800 ;
        RECT 378.800 331.600 379.600 333.200 ;
        RECT 380.600 330.200 381.200 333.600 ;
        RECT 382.000 332.300 382.800 333.200 ;
        RECT 386.800 332.300 387.600 335.800 ;
        RECT 382.000 331.700 387.600 332.300 ;
        RECT 382.000 331.600 382.800 331.700 ;
        RECT 370.800 329.600 372.200 330.200 ;
        RECT 372.800 329.600 373.800 330.200 ;
        RECT 371.600 328.400 372.200 329.600 ;
        RECT 373.000 328.400 373.800 329.600 ;
        RECT 371.600 327.600 372.400 328.400 ;
        RECT 373.000 327.600 374.800 328.400 ;
        RECT 368.000 326.800 370.000 327.400 ;
        RECT 359.600 322.200 360.400 325.000 ;
        RECT 361.200 322.200 362.000 325.000 ;
        RECT 364.400 322.200 365.200 326.800 ;
        RECT 368.000 326.200 368.600 326.800 ;
        RECT 367.600 325.600 368.600 326.200 ;
        RECT 367.600 322.200 368.400 325.600 ;
        RECT 373.000 322.200 373.800 327.600 ;
        RECT 379.800 322.200 381.800 330.200 ;
        RECT 385.200 328.800 386.000 330.400 ;
        RECT 386.800 322.200 387.600 331.700 ;
        RECT 391.400 335.800 392.400 336.400 ;
        RECT 391.400 334.400 392.000 335.800 ;
        RECT 394.800 335.200 395.600 339.800 ;
        RECT 398.000 336.000 398.800 339.800 ;
        RECT 393.000 334.600 395.600 335.200 ;
        RECT 397.800 335.200 398.800 336.000 ;
        RECT 391.400 333.600 392.400 334.400 ;
        RECT 391.400 330.200 392.000 333.600 ;
        RECT 393.000 333.000 393.600 334.600 ;
        RECT 392.600 332.200 393.600 333.000 ;
        RECT 393.000 330.200 393.600 332.200 ;
        RECT 394.600 332.400 395.400 333.200 ;
        RECT 394.600 332.300 395.600 332.400 ;
        RECT 397.800 332.300 398.600 335.200 ;
        RECT 399.600 334.600 400.400 339.800 ;
        RECT 406.000 336.600 406.800 339.800 ;
        RECT 407.600 337.000 408.400 339.800 ;
        RECT 409.200 337.000 410.000 339.800 ;
        RECT 410.800 337.000 411.600 339.800 ;
        RECT 412.400 337.000 413.200 339.800 ;
        RECT 415.600 337.000 416.400 339.800 ;
        RECT 418.800 337.000 419.600 339.800 ;
        RECT 420.400 337.000 421.200 339.800 ;
        RECT 422.000 337.000 422.800 339.800 ;
        RECT 404.400 335.800 406.800 336.600 ;
        RECT 423.600 336.600 424.400 339.800 ;
        RECT 404.400 335.200 405.200 335.800 ;
        RECT 394.600 331.700 398.600 332.300 ;
        RECT 394.600 331.600 395.600 331.700 ;
        RECT 397.800 330.800 398.600 331.700 ;
        RECT 399.200 334.000 400.400 334.600 ;
        RECT 403.400 334.600 405.200 335.200 ;
        RECT 409.200 335.600 410.200 336.400 ;
        RECT 413.200 335.600 414.800 336.400 ;
        RECT 415.600 335.800 420.200 336.400 ;
        RECT 423.600 335.800 426.200 336.600 ;
        RECT 415.600 335.600 416.400 335.800 ;
        RECT 399.200 332.000 399.800 334.000 ;
        RECT 403.400 333.400 404.200 334.600 ;
        RECT 400.400 332.600 404.200 333.400 ;
        RECT 409.200 332.800 410.000 335.600 ;
        RECT 415.600 334.800 416.400 335.000 ;
        RECT 412.000 334.200 416.400 334.800 ;
        RECT 412.000 334.000 412.800 334.200 ;
        RECT 417.200 333.600 418.000 335.200 ;
        RECT 419.400 333.400 420.200 335.800 ;
        RECT 425.400 335.200 426.200 335.800 ;
        RECT 425.400 334.400 428.400 335.200 ;
        RECT 430.000 333.800 430.800 339.800 ;
        RECT 432.200 336.400 433.000 339.800 ;
        RECT 432.200 335.800 434.000 336.400 ;
        RECT 412.400 332.600 415.600 333.400 ;
        RECT 419.400 332.600 421.400 333.400 ;
        RECT 422.000 333.000 430.800 333.800 ;
        RECT 406.000 332.000 406.800 332.600 ;
        RECT 423.600 332.000 424.400 332.400 ;
        RECT 428.600 332.000 429.400 332.200 ;
        RECT 399.200 331.400 400.000 332.000 ;
        RECT 406.000 331.400 429.400 332.000 ;
        RECT 391.400 329.200 392.400 330.200 ;
        RECT 393.000 329.600 395.600 330.200 ;
        RECT 397.800 330.000 398.800 330.800 ;
        RECT 391.600 322.200 392.400 329.200 ;
        RECT 394.800 322.200 395.600 329.600 ;
        RECT 398.000 322.200 398.800 330.000 ;
        RECT 399.400 329.600 400.000 331.400 ;
        RECT 399.400 329.000 408.400 329.600 ;
        RECT 399.400 327.400 400.000 329.000 ;
        RECT 407.600 328.800 408.400 329.000 ;
        RECT 410.800 329.000 419.400 329.600 ;
        RECT 410.800 328.800 411.600 329.000 ;
        RECT 402.600 327.600 405.200 328.400 ;
        RECT 399.400 326.800 402.000 327.400 ;
        RECT 401.200 322.200 402.000 326.800 ;
        RECT 404.400 322.200 405.200 327.600 ;
        RECT 405.800 326.800 410.000 327.600 ;
        RECT 407.600 322.200 408.400 325.000 ;
        RECT 409.200 322.200 410.000 325.000 ;
        RECT 410.800 322.200 411.600 325.000 ;
        RECT 412.400 322.200 413.200 328.400 ;
        RECT 415.600 327.600 418.200 328.400 ;
        RECT 418.800 328.200 419.400 329.000 ;
        RECT 420.400 329.400 421.200 329.600 ;
        RECT 420.400 329.000 425.800 329.400 ;
        RECT 420.400 328.800 426.600 329.000 ;
        RECT 425.200 328.200 426.600 328.800 ;
        RECT 418.800 327.600 424.600 328.200 ;
        RECT 427.600 328.000 429.200 328.800 ;
        RECT 427.600 327.600 428.200 328.000 ;
        RECT 415.600 322.200 416.400 327.000 ;
        RECT 418.800 322.200 419.600 327.000 ;
        RECT 424.000 326.800 428.200 327.600 ;
        RECT 430.000 327.400 430.800 333.000 ;
        RECT 431.600 328.800 432.400 330.400 ;
        RECT 428.800 326.800 430.800 327.400 ;
        RECT 420.400 322.200 421.200 325.000 ;
        RECT 422.000 322.200 422.800 325.000 ;
        RECT 425.200 322.200 426.000 326.800 ;
        RECT 428.800 326.200 429.400 326.800 ;
        RECT 428.400 325.600 429.400 326.200 ;
        RECT 428.400 322.200 429.200 325.600 ;
        RECT 433.200 322.200 434.000 335.800 ;
        RECT 436.400 335.600 437.200 337.200 ;
        RECT 434.800 333.600 435.600 335.200 ;
        RECT 438.000 332.300 438.800 339.800 ;
        RECT 439.600 336.000 440.400 339.800 ;
        RECT 442.800 336.000 443.600 339.800 ;
        RECT 439.600 335.800 443.600 336.000 ;
        RECT 444.400 335.800 445.200 339.800 ;
        RECT 446.000 336.000 446.800 339.800 ;
        RECT 449.200 336.000 450.000 339.800 ;
        RECT 446.000 335.800 450.000 336.000 ;
        RECT 450.800 335.800 451.600 339.800 ;
        RECT 455.000 336.400 455.800 339.800 ;
        RECT 454.000 335.800 455.800 336.400 ;
        RECT 465.200 335.800 466.000 339.800 ;
        RECT 470.000 337.800 470.800 339.800 ;
        RECT 466.600 336.400 467.400 337.200 ;
        RECT 439.800 335.400 443.400 335.800 ;
        RECT 440.400 334.400 441.200 334.800 ;
        RECT 444.400 334.400 445.000 335.800 ;
        RECT 446.200 335.400 449.800 335.800 ;
        RECT 446.800 334.400 447.600 334.800 ;
        RECT 450.800 334.400 451.400 335.800 ;
        RECT 439.600 333.800 441.200 334.400 ;
        RECT 439.600 333.600 440.400 333.800 ;
        RECT 442.600 333.600 445.200 334.400 ;
        RECT 446.000 333.800 447.600 334.400 ;
        RECT 446.000 333.600 446.800 333.800 ;
        RECT 449.000 333.600 451.600 334.400 ;
        RECT 452.400 333.600 453.200 335.200 ;
        RECT 441.200 332.300 442.000 333.200 ;
        RECT 438.000 331.700 442.000 332.300 ;
        RECT 438.000 322.200 438.800 331.700 ;
        RECT 441.200 331.600 442.000 331.700 ;
        RECT 442.600 330.400 443.200 333.600 ;
        RECT 447.600 331.600 448.400 333.200 ;
        RECT 441.200 329.600 443.200 330.400 ;
        RECT 444.400 330.200 445.200 330.400 ;
        RECT 449.000 330.200 449.600 333.600 ;
        RECT 454.000 332.300 454.800 335.800 ;
        RECT 455.600 334.300 456.400 334.400 ;
        RECT 463.600 334.300 464.400 334.400 ;
        RECT 455.600 333.700 464.400 334.300 ;
        RECT 455.600 333.600 456.400 333.700 ;
        RECT 463.600 332.800 464.400 333.700 ;
        RECT 460.400 332.300 461.200 332.400 ;
        RECT 454.000 331.700 461.200 332.300 ;
        RECT 450.800 330.200 451.600 330.400 ;
        RECT 443.800 329.600 445.200 330.200 ;
        RECT 448.600 329.600 449.600 330.200 ;
        RECT 450.200 329.600 451.600 330.200 ;
        RECT 442.200 322.200 443.000 329.600 ;
        RECT 443.800 328.400 444.400 329.600 ;
        RECT 443.600 327.600 444.400 328.400 ;
        RECT 448.600 322.200 449.400 329.600 ;
        RECT 450.200 328.400 450.800 329.600 ;
        RECT 450.000 327.600 450.800 328.400 ;
        RECT 454.000 322.200 454.800 331.700 ;
        RECT 460.400 331.600 461.200 331.700 ;
        RECT 462.000 332.200 462.800 332.400 ;
        RECT 465.200 332.200 465.800 335.800 ;
        RECT 466.800 335.600 467.600 336.400 ;
        RECT 468.400 335.600 469.200 337.200 ;
        RECT 470.200 334.400 470.800 337.800 ;
        RECT 470.000 334.300 470.800 334.400 ;
        RECT 474.800 337.800 475.600 339.800 ;
        RECT 474.800 334.400 475.400 337.800 ;
        RECT 476.400 336.300 477.200 337.200 ;
        RECT 478.000 336.300 478.800 339.800 ;
        RECT 476.400 335.700 478.800 336.300 ;
        RECT 479.600 336.000 480.400 339.800 ;
        RECT 482.800 336.000 483.600 339.800 ;
        RECT 487.000 336.400 487.800 339.800 ;
        RECT 479.600 335.800 483.600 336.000 ;
        RECT 486.000 335.800 487.800 336.400 ;
        RECT 476.400 335.600 477.200 335.700 ;
        RECT 478.200 334.400 478.800 335.700 ;
        RECT 479.800 335.400 483.400 335.800 ;
        RECT 482.000 334.400 482.800 334.800 ;
        RECT 470.000 333.700 473.900 334.300 ;
        RECT 470.000 333.600 470.800 333.700 ;
        RECT 466.800 332.200 467.600 332.400 ;
        RECT 462.000 331.600 463.600 332.200 ;
        RECT 465.200 331.600 467.600 332.200 ;
        RECT 462.800 331.200 463.600 331.600 ;
        RECT 455.600 328.800 456.400 330.400 ;
        RECT 466.800 330.200 467.400 331.600 ;
        RECT 470.200 330.200 470.800 333.600 ;
        RECT 473.300 332.400 473.900 333.700 ;
        RECT 474.800 333.600 475.600 334.400 ;
        RECT 478.000 333.600 480.600 334.400 ;
        RECT 482.000 333.800 483.600 334.400 ;
        RECT 482.800 333.600 483.600 333.800 ;
        RECT 484.400 333.600 485.200 335.200 ;
        RECT 471.600 330.800 472.400 332.400 ;
        RECT 473.200 330.800 474.000 332.400 ;
        RECT 474.800 330.200 475.400 333.600 ;
        RECT 478.000 330.200 478.800 330.400 ;
        RECT 480.000 330.200 480.600 333.600 ;
        RECT 481.200 331.600 482.000 333.200 ;
        RECT 462.000 329.600 466.000 330.200 ;
        RECT 462.000 322.200 462.800 329.600 ;
        RECT 465.200 322.200 466.000 329.600 ;
        RECT 466.800 322.200 467.600 330.200 ;
        RECT 470.000 329.400 471.800 330.200 ;
        RECT 471.000 322.200 471.800 329.400 ;
        RECT 473.800 329.400 475.600 330.200 ;
        RECT 478.000 329.600 479.400 330.200 ;
        RECT 480.000 329.600 481.000 330.200 ;
        RECT 473.800 324.400 474.600 329.400 ;
        RECT 478.800 328.400 479.400 329.600 ;
        RECT 478.800 327.600 479.600 328.400 ;
        RECT 473.800 323.600 475.600 324.400 ;
        RECT 473.800 322.200 474.600 323.600 ;
        RECT 480.200 322.200 481.000 329.600 ;
        RECT 486.000 322.200 486.800 335.800 ;
        RECT 489.200 333.600 490.000 335.200 ;
        RECT 487.600 328.800 488.400 330.400 ;
        RECT 490.800 322.200 491.600 339.800 ;
        RECT 497.600 334.200 498.400 339.800 ;
        RECT 502.000 337.800 502.800 339.800 ;
        RECT 502.000 334.400 502.600 337.800 ;
        RECT 503.600 336.300 504.400 337.200 ;
        RECT 505.200 336.300 506.000 336.400 ;
        RECT 503.600 335.700 506.000 336.300 ;
        RECT 506.800 336.000 507.600 339.800 ;
        RECT 503.600 335.600 504.400 335.700 ;
        RECT 505.200 335.600 506.000 335.700 ;
        RECT 506.600 335.200 507.600 336.000 ;
        RECT 497.600 333.800 499.400 334.200 ;
        RECT 497.800 333.600 499.400 333.800 ;
        RECT 495.600 331.600 497.200 332.400 ;
        RECT 494.000 329.600 494.800 331.200 ;
        RECT 498.800 330.400 499.400 333.600 ;
        RECT 502.000 333.600 502.800 334.400 ;
        RECT 500.400 330.800 501.200 332.400 ;
        RECT 498.800 329.600 499.600 330.400 ;
        RECT 502.000 330.200 502.600 333.600 ;
        RECT 506.600 330.800 507.400 335.200 ;
        RECT 508.400 334.600 509.200 339.800 ;
        RECT 514.800 336.600 515.600 339.800 ;
        RECT 516.400 337.000 517.200 339.800 ;
        RECT 518.000 337.000 518.800 339.800 ;
        RECT 519.600 337.000 520.400 339.800 ;
        RECT 521.200 337.000 522.000 339.800 ;
        RECT 524.400 337.000 525.200 339.800 ;
        RECT 527.600 337.000 528.400 339.800 ;
        RECT 529.200 337.000 530.000 339.800 ;
        RECT 530.800 337.000 531.600 339.800 ;
        RECT 513.200 335.800 515.600 336.600 ;
        RECT 532.400 336.600 533.200 339.800 ;
        RECT 513.200 335.200 514.000 335.800 ;
        RECT 508.000 334.000 509.200 334.600 ;
        RECT 512.200 334.600 514.000 335.200 ;
        RECT 518.000 335.600 519.000 336.400 ;
        RECT 522.000 335.600 523.600 336.400 ;
        RECT 524.400 335.800 529.000 336.400 ;
        RECT 532.400 335.800 535.000 336.600 ;
        RECT 524.400 335.600 525.200 335.800 ;
        RECT 508.000 332.000 508.600 334.000 ;
        RECT 512.200 333.400 513.000 334.600 ;
        RECT 509.200 332.600 513.000 333.400 ;
        RECT 518.000 332.800 518.800 335.600 ;
        RECT 524.400 334.800 525.200 335.000 ;
        RECT 520.800 334.200 525.200 334.800 ;
        RECT 520.800 334.000 521.600 334.200 ;
        RECT 526.000 333.600 526.800 335.200 ;
        RECT 528.200 333.400 529.000 335.800 ;
        RECT 534.200 335.200 535.000 335.800 ;
        RECT 534.200 334.400 537.200 335.200 ;
        RECT 538.800 333.800 539.600 339.800 ;
        RECT 521.200 332.600 524.400 333.400 ;
        RECT 528.200 332.600 530.200 333.400 ;
        RECT 530.800 333.000 539.600 333.800 ;
        RECT 514.800 332.000 515.600 332.600 ;
        RECT 532.400 332.000 533.200 332.400 ;
        RECT 535.600 332.000 536.400 332.400 ;
        RECT 537.400 332.000 538.200 332.200 ;
        RECT 508.000 331.400 508.800 332.000 ;
        RECT 514.800 331.400 538.200 332.000 ;
        RECT 495.600 328.300 496.400 328.400 ;
        RECT 497.200 328.300 498.000 329.200 ;
        RECT 495.600 327.700 498.000 328.300 ;
        RECT 495.600 327.600 496.400 327.700 ;
        RECT 497.200 327.600 498.000 327.700 ;
        RECT 498.800 327.000 499.400 329.600 ;
        RECT 495.800 326.400 499.400 327.000 ;
        RECT 495.800 326.200 496.400 326.400 ;
        RECT 495.600 322.200 496.400 326.200 ;
        RECT 498.800 326.200 499.400 326.400 ;
        RECT 501.000 329.400 502.800 330.200 ;
        RECT 506.600 330.000 507.600 330.800 ;
        RECT 498.800 322.200 499.600 326.200 ;
        RECT 501.000 324.400 501.800 329.400 ;
        RECT 501.000 323.600 502.800 324.400 ;
        RECT 501.000 322.200 501.800 323.600 ;
        RECT 506.800 322.200 507.600 330.000 ;
        RECT 508.200 329.600 508.800 331.400 ;
        RECT 508.200 329.000 517.200 329.600 ;
        RECT 508.200 327.400 508.800 329.000 ;
        RECT 516.400 328.800 517.200 329.000 ;
        RECT 519.600 329.000 528.200 329.600 ;
        RECT 519.600 328.800 520.400 329.000 ;
        RECT 511.400 327.600 514.000 328.400 ;
        RECT 508.200 326.800 510.800 327.400 ;
        RECT 510.000 322.200 510.800 326.800 ;
        RECT 513.200 322.200 514.000 327.600 ;
        RECT 514.600 326.800 518.800 327.600 ;
        RECT 516.400 322.200 517.200 325.000 ;
        RECT 518.000 322.200 518.800 325.000 ;
        RECT 519.600 322.200 520.400 325.000 ;
        RECT 521.200 322.200 522.000 328.400 ;
        RECT 524.400 327.600 527.000 328.400 ;
        RECT 527.600 328.200 528.200 329.000 ;
        RECT 529.200 329.400 530.000 329.600 ;
        RECT 529.200 329.000 534.600 329.400 ;
        RECT 529.200 328.800 535.400 329.000 ;
        RECT 534.000 328.200 535.400 328.800 ;
        RECT 527.600 327.600 533.400 328.200 ;
        RECT 536.400 328.000 538.000 328.800 ;
        RECT 536.400 327.600 537.000 328.000 ;
        RECT 524.400 322.200 525.200 327.000 ;
        RECT 527.600 322.200 528.400 327.000 ;
        RECT 532.800 326.800 537.000 327.600 ;
        RECT 538.800 327.400 539.600 333.000 ;
        RECT 537.600 326.800 539.600 327.400 ;
        RECT 540.400 333.800 541.200 339.800 ;
        RECT 546.800 336.600 547.600 339.800 ;
        RECT 548.400 337.000 549.200 339.800 ;
        RECT 550.000 337.000 550.800 339.800 ;
        RECT 551.600 337.000 552.400 339.800 ;
        RECT 554.800 337.000 555.600 339.800 ;
        RECT 558.000 337.000 558.800 339.800 ;
        RECT 559.600 337.000 560.400 339.800 ;
        RECT 561.200 337.000 562.000 339.800 ;
        RECT 562.800 337.000 563.600 339.800 ;
        RECT 545.000 335.800 547.600 336.600 ;
        RECT 564.400 336.600 565.200 339.800 ;
        RECT 551.000 335.800 555.600 336.400 ;
        RECT 545.000 335.200 545.800 335.800 ;
        RECT 542.800 334.400 545.800 335.200 ;
        RECT 540.400 333.000 549.200 333.800 ;
        RECT 551.000 333.400 551.800 335.800 ;
        RECT 554.800 335.600 555.600 335.800 ;
        RECT 556.400 335.600 558.000 336.400 ;
        RECT 561.000 335.600 562.000 336.400 ;
        RECT 564.400 335.800 566.800 336.600 ;
        RECT 553.200 333.600 554.000 335.200 ;
        RECT 554.800 334.800 555.600 335.000 ;
        RECT 554.800 334.200 559.200 334.800 ;
        RECT 558.400 334.000 559.200 334.200 ;
        RECT 540.400 327.400 541.200 333.000 ;
        RECT 549.800 332.600 551.800 333.400 ;
        RECT 555.600 332.600 558.800 333.400 ;
        RECT 561.200 332.800 562.000 335.600 ;
        RECT 566.000 335.200 566.800 335.800 ;
        RECT 566.000 334.600 567.800 335.200 ;
        RECT 567.000 333.400 567.800 334.600 ;
        RECT 570.800 334.600 571.600 339.800 ;
        RECT 572.400 336.000 573.200 339.800 ;
        RECT 576.200 336.400 577.000 339.800 ;
        RECT 572.400 335.200 573.400 336.000 ;
        RECT 576.200 335.800 578.000 336.400 ;
        RECT 580.400 335.800 581.200 339.800 ;
        RECT 582.000 336.000 582.800 339.800 ;
        RECT 585.200 336.000 586.000 339.800 ;
        RECT 582.000 335.800 586.000 336.000 ;
        RECT 570.800 334.000 572.000 334.600 ;
        RECT 567.000 332.600 570.800 333.400 ;
        RECT 541.800 332.000 542.600 332.200 ;
        RECT 543.600 332.000 544.400 332.400 ;
        RECT 546.800 332.000 547.600 332.400 ;
        RECT 564.400 332.000 565.200 332.600 ;
        RECT 571.400 332.000 572.000 334.000 ;
        RECT 541.800 331.400 565.200 332.000 ;
        RECT 571.200 331.400 572.000 332.000 ;
        RECT 571.200 329.600 571.800 331.400 ;
        RECT 572.600 330.800 573.400 335.200 ;
        RECT 550.000 329.400 550.800 329.600 ;
        RECT 545.400 329.000 550.800 329.400 ;
        RECT 544.600 328.800 550.800 329.000 ;
        RECT 551.800 329.000 560.400 329.600 ;
        RECT 542.000 328.000 543.600 328.800 ;
        RECT 544.600 328.200 546.000 328.800 ;
        RECT 551.800 328.200 552.400 329.000 ;
        RECT 559.600 328.800 560.400 329.000 ;
        RECT 562.800 329.000 571.800 329.600 ;
        RECT 562.800 328.800 563.600 329.000 ;
        RECT 543.000 327.600 543.600 328.000 ;
        RECT 546.600 327.600 552.400 328.200 ;
        RECT 553.000 327.600 555.600 328.400 ;
        RECT 540.400 326.800 542.400 327.400 ;
        RECT 543.000 326.800 547.200 327.600 ;
        RECT 529.200 322.200 530.000 325.000 ;
        RECT 530.800 322.200 531.600 325.000 ;
        RECT 534.000 322.200 534.800 326.800 ;
        RECT 537.600 326.200 538.200 326.800 ;
        RECT 537.200 325.600 538.200 326.200 ;
        RECT 541.800 326.200 542.400 326.800 ;
        RECT 541.800 325.600 542.800 326.200 ;
        RECT 537.200 322.200 538.000 325.600 ;
        RECT 542.000 322.200 542.800 325.600 ;
        RECT 545.200 322.200 546.000 326.800 ;
        RECT 548.400 322.200 549.200 325.000 ;
        RECT 550.000 322.200 550.800 325.000 ;
        RECT 551.600 322.200 552.400 327.000 ;
        RECT 554.800 322.200 555.600 327.000 ;
        RECT 558.000 322.200 558.800 328.400 ;
        RECT 566.000 327.600 568.600 328.400 ;
        RECT 561.200 326.800 565.400 327.600 ;
        RECT 559.600 322.200 560.400 325.000 ;
        RECT 561.200 322.200 562.000 325.000 ;
        RECT 562.800 322.200 563.600 325.000 ;
        RECT 566.000 322.200 566.800 327.600 ;
        RECT 571.200 327.400 571.800 329.000 ;
        RECT 569.200 326.800 571.800 327.400 ;
        RECT 572.400 330.300 573.400 330.800 ;
        RECT 575.600 330.300 576.400 330.400 ;
        RECT 572.400 329.700 576.400 330.300 ;
        RECT 569.200 322.200 570.000 326.800 ;
        RECT 572.400 322.200 573.200 329.700 ;
        RECT 575.600 328.800 576.400 329.700 ;
        RECT 577.200 330.300 578.000 335.800 ;
        RECT 578.800 333.600 579.600 335.200 ;
        RECT 580.600 334.400 581.200 335.800 ;
        RECT 582.200 335.400 585.800 335.800 ;
        RECT 584.400 334.400 585.200 334.800 ;
        RECT 580.400 333.600 583.000 334.400 ;
        RECT 584.400 333.800 586.000 334.400 ;
        RECT 585.200 333.600 586.000 333.800 ;
        RECT 580.400 330.300 581.200 330.400 ;
        RECT 577.200 330.200 581.200 330.300 ;
        RECT 582.400 330.200 583.000 333.600 ;
        RECT 583.600 332.300 584.400 333.200 ;
        RECT 586.800 332.300 587.600 339.800 ;
        RECT 588.400 335.600 589.200 337.200 ;
        RECT 592.600 336.400 593.400 339.800 ;
        RECT 591.600 335.800 593.400 336.400 ;
        RECT 594.800 335.800 595.600 339.800 ;
        RECT 596.400 336.000 597.200 339.800 ;
        RECT 599.600 336.000 600.400 339.800 ;
        RECT 596.400 335.800 600.400 336.000 ;
        RECT 590.000 333.600 590.800 335.200 ;
        RECT 583.600 331.700 587.600 332.300 ;
        RECT 583.600 331.600 584.400 331.700 ;
        RECT 577.200 329.700 581.800 330.200 ;
        RECT 577.200 322.200 578.000 329.700 ;
        RECT 580.400 329.600 581.800 329.700 ;
        RECT 582.400 329.600 583.400 330.200 ;
        RECT 581.200 328.400 581.800 329.600 ;
        RECT 581.200 327.600 582.000 328.400 ;
        RECT 582.600 322.200 583.400 329.600 ;
        RECT 586.800 322.200 587.600 331.700 ;
        RECT 591.600 322.200 592.400 335.800 ;
        RECT 595.000 334.400 595.600 335.800 ;
        RECT 596.600 335.400 600.200 335.800 ;
        RECT 598.800 334.400 599.600 334.800 ;
        RECT 593.200 334.300 594.000 334.400 ;
        RECT 594.800 334.300 597.400 334.400 ;
        RECT 593.200 333.700 597.400 334.300 ;
        RECT 598.800 333.800 600.400 334.400 ;
        RECT 593.200 333.600 594.000 333.700 ;
        RECT 594.800 333.600 597.400 333.700 ;
        RECT 599.600 333.600 600.400 333.800 ;
        RECT 593.200 328.800 594.000 330.400 ;
        RECT 594.800 330.200 595.600 330.400 ;
        RECT 596.800 330.200 597.400 333.600 ;
        RECT 598.000 332.300 598.800 333.200 ;
        RECT 601.200 332.300 602.000 339.800 ;
        RECT 602.800 335.600 603.600 337.200 ;
        RECT 598.000 331.700 602.000 332.300 ;
        RECT 598.000 331.600 598.800 331.700 ;
        RECT 594.800 329.600 596.200 330.200 ;
        RECT 596.800 329.600 597.800 330.200 ;
        RECT 595.600 328.400 596.200 329.600 ;
        RECT 595.600 327.600 596.400 328.400 ;
        RECT 597.000 322.200 597.800 329.600 ;
        RECT 601.200 322.200 602.000 331.700 ;
        RECT 606.000 335.200 606.800 339.800 ;
        RECT 609.200 335.200 610.000 339.800 ;
        RECT 606.000 334.400 610.000 335.200 ;
        RECT 606.000 331.600 606.800 334.400 ;
        RECT 606.000 330.800 610.000 331.600 ;
        RECT 606.000 322.200 606.800 330.800 ;
        RECT 609.200 322.200 610.000 330.800 ;
        RECT 2.800 311.200 3.600 319.800 ;
        RECT 6.000 311.200 6.800 319.800 ;
        RECT 9.200 311.200 10.000 319.800 ;
        RECT 12.400 311.200 13.200 319.800 ;
        RECT 17.200 316.400 18.000 319.800 ;
        RECT 17.000 315.800 18.000 316.400 ;
        RECT 17.000 315.200 17.600 315.800 ;
        RECT 20.400 315.200 21.200 319.800 ;
        RECT 23.600 317.000 24.400 319.800 ;
        RECT 25.200 317.000 26.000 319.800 ;
        RECT 15.600 314.600 17.600 315.200 ;
        RECT 2.800 310.400 4.600 311.200 ;
        RECT 6.000 310.400 8.200 311.200 ;
        RECT 9.200 310.400 11.400 311.200 ;
        RECT 12.400 310.400 14.800 311.200 ;
        RECT 3.800 309.000 4.600 310.400 ;
        RECT 7.400 309.000 8.200 310.400 ;
        RECT 10.600 309.000 11.400 310.400 ;
        RECT 1.200 308.200 3.000 309.000 ;
        RECT 3.800 308.200 6.400 309.000 ;
        RECT 7.400 308.200 9.800 309.000 ;
        RECT 10.600 308.200 13.200 309.000 ;
        RECT 1.200 307.600 2.000 308.200 ;
        RECT 3.800 307.600 4.600 308.200 ;
        RECT 7.400 307.600 8.200 308.200 ;
        RECT 10.600 307.600 11.400 308.200 ;
        RECT 14.000 307.600 14.800 310.400 ;
        RECT 2.800 306.800 4.600 307.600 ;
        RECT 6.000 306.800 8.200 307.600 ;
        RECT 9.200 306.800 11.400 307.600 ;
        RECT 12.400 306.800 14.800 307.600 ;
        RECT 15.600 309.000 16.400 314.600 ;
        RECT 18.200 314.400 22.400 315.200 ;
        RECT 26.800 315.000 27.600 319.800 ;
        RECT 30.000 315.000 30.800 319.800 ;
        RECT 18.200 314.000 18.800 314.400 ;
        RECT 17.200 313.200 18.800 314.000 ;
        RECT 21.800 313.800 27.600 314.400 ;
        RECT 19.800 313.200 21.200 313.800 ;
        RECT 19.800 313.000 26.000 313.200 ;
        RECT 20.600 312.600 26.000 313.000 ;
        RECT 25.200 312.400 26.000 312.600 ;
        RECT 27.000 313.000 27.600 313.800 ;
        RECT 28.200 313.600 30.800 314.400 ;
        RECT 33.200 313.600 34.000 319.800 ;
        RECT 34.800 317.000 35.600 319.800 ;
        RECT 36.400 317.000 37.200 319.800 ;
        RECT 38.000 317.000 38.800 319.800 ;
        RECT 36.400 314.400 40.600 315.200 ;
        RECT 41.200 314.400 42.000 319.800 ;
        RECT 44.400 315.200 45.200 319.800 ;
        RECT 44.400 314.600 47.000 315.200 ;
        RECT 41.200 313.600 43.800 314.400 ;
        RECT 34.800 313.000 35.600 313.200 ;
        RECT 27.000 312.400 35.600 313.000 ;
        RECT 38.000 313.000 38.800 313.200 ;
        RECT 46.400 313.000 47.000 314.600 ;
        RECT 38.000 312.400 47.000 313.000 ;
        RECT 46.400 310.600 47.000 312.400 ;
        RECT 47.600 312.000 48.400 319.800 ;
        RECT 52.400 312.000 53.200 319.800 ;
        RECT 55.600 315.200 56.400 319.800 ;
        RECT 47.600 311.200 48.600 312.000 ;
        RECT 17.000 310.000 40.400 310.600 ;
        RECT 46.400 310.000 47.200 310.600 ;
        RECT 17.000 309.800 17.800 310.000 ;
        RECT 18.800 309.600 19.600 310.000 ;
        RECT 22.000 309.600 22.800 310.000 ;
        RECT 39.600 309.400 40.400 310.000 ;
        RECT 15.600 308.200 24.400 309.000 ;
        RECT 25.000 308.600 27.000 309.400 ;
        RECT 30.800 308.600 34.000 309.400 ;
        RECT 2.800 302.200 3.600 306.800 ;
        RECT 6.000 302.200 6.800 306.800 ;
        RECT 9.200 302.200 10.000 306.800 ;
        RECT 12.400 302.200 13.200 306.800 ;
        RECT 15.600 302.200 16.400 308.200 ;
        RECT 18.000 306.800 21.000 307.600 ;
        RECT 20.200 306.200 21.000 306.800 ;
        RECT 26.200 306.200 27.000 308.600 ;
        RECT 28.400 306.800 29.200 308.400 ;
        RECT 33.600 307.800 34.400 308.000 ;
        RECT 30.000 307.200 34.400 307.800 ;
        RECT 30.000 307.000 30.800 307.200 ;
        RECT 36.400 306.400 37.200 309.200 ;
        RECT 42.200 308.600 46.000 309.400 ;
        RECT 42.200 307.400 43.000 308.600 ;
        RECT 46.600 308.000 47.200 310.000 ;
        RECT 30.000 306.200 30.800 306.400 ;
        RECT 20.200 305.400 22.800 306.200 ;
        RECT 26.200 305.600 30.800 306.200 ;
        RECT 31.600 305.600 33.200 306.400 ;
        RECT 36.200 305.600 37.200 306.400 ;
        RECT 41.200 306.800 43.000 307.400 ;
        RECT 46.000 307.400 47.200 308.000 ;
        RECT 41.200 306.200 42.000 306.800 ;
        RECT 22.000 302.200 22.800 305.400 ;
        RECT 39.600 305.400 42.000 306.200 ;
        RECT 23.600 302.200 24.400 305.000 ;
        RECT 25.200 302.200 26.000 305.000 ;
        RECT 26.800 302.200 27.600 305.000 ;
        RECT 30.000 302.200 30.800 305.000 ;
        RECT 33.200 302.200 34.000 305.000 ;
        RECT 34.800 302.200 35.600 305.000 ;
        RECT 36.400 302.200 37.200 305.000 ;
        RECT 38.000 302.200 38.800 305.000 ;
        RECT 39.600 302.200 40.400 305.400 ;
        RECT 46.000 302.200 46.800 307.400 ;
        RECT 47.800 306.800 48.600 311.200 ;
        RECT 47.600 306.000 48.600 306.800 ;
        RECT 52.200 311.200 53.200 312.000 ;
        RECT 53.800 314.600 56.400 315.200 ;
        RECT 53.800 313.000 54.400 314.600 ;
        RECT 58.800 314.400 59.600 319.800 ;
        RECT 62.000 317.000 62.800 319.800 ;
        RECT 63.600 317.000 64.400 319.800 ;
        RECT 65.200 317.000 66.000 319.800 ;
        RECT 60.200 314.400 64.400 315.200 ;
        RECT 57.000 313.600 59.600 314.400 ;
        RECT 66.800 313.600 67.600 319.800 ;
        RECT 70.000 315.000 70.800 319.800 ;
        RECT 73.200 315.000 74.000 319.800 ;
        RECT 74.800 317.000 75.600 319.800 ;
        RECT 76.400 317.000 77.200 319.800 ;
        RECT 79.600 315.200 80.400 319.800 ;
        RECT 82.800 316.400 83.600 319.800 ;
        RECT 82.800 315.800 83.800 316.400 ;
        RECT 83.200 315.200 83.800 315.800 ;
        RECT 78.400 314.400 82.600 315.200 ;
        RECT 83.200 314.600 85.200 315.200 ;
        RECT 70.000 313.600 72.600 314.400 ;
        RECT 73.200 313.800 79.000 314.400 ;
        RECT 82.000 314.000 82.600 314.400 ;
        RECT 62.000 313.000 62.800 313.200 ;
        RECT 53.800 312.400 62.800 313.000 ;
        RECT 65.200 313.000 66.000 313.200 ;
        RECT 73.200 313.000 73.800 313.800 ;
        RECT 79.600 313.200 81.000 313.800 ;
        RECT 82.000 313.200 83.600 314.000 ;
        RECT 65.200 312.400 73.800 313.000 ;
        RECT 74.800 313.000 81.000 313.200 ;
        RECT 74.800 312.600 80.200 313.000 ;
        RECT 74.800 312.400 75.600 312.600 ;
        RECT 52.200 306.800 53.000 311.200 ;
        RECT 53.800 310.600 54.400 312.400 ;
        RECT 53.600 310.000 54.400 310.600 ;
        RECT 60.400 310.000 83.800 310.600 ;
        RECT 53.600 308.000 54.200 310.000 ;
        RECT 60.400 309.400 61.200 310.000 ;
        RECT 78.000 309.600 78.800 310.000 ;
        RECT 79.600 309.600 80.400 310.000 ;
        RECT 83.000 309.800 83.800 310.000 ;
        RECT 54.800 308.600 58.600 309.400 ;
        RECT 53.600 307.400 54.800 308.000 ;
        RECT 52.200 306.000 53.200 306.800 ;
        RECT 47.600 302.200 48.400 306.000 ;
        RECT 52.400 302.200 53.200 306.000 ;
        RECT 54.000 302.200 54.800 307.400 ;
        RECT 57.800 307.400 58.600 308.600 ;
        RECT 57.800 306.800 59.600 307.400 ;
        RECT 58.800 306.200 59.600 306.800 ;
        RECT 63.600 306.400 64.400 309.200 ;
        RECT 66.800 308.600 70.000 309.400 ;
        RECT 73.800 308.600 75.800 309.400 ;
        RECT 84.400 309.000 85.200 314.600 ;
        RECT 89.800 312.800 90.600 319.800 ;
        RECT 94.000 315.000 94.800 319.000 ;
        RECT 89.000 312.200 90.600 312.800 ;
        RECT 87.600 309.600 88.400 311.200 ;
        RECT 66.400 307.800 67.200 308.000 ;
        RECT 66.400 307.200 70.800 307.800 ;
        RECT 70.000 307.000 70.800 307.200 ;
        RECT 71.600 306.800 72.400 308.400 ;
        RECT 58.800 305.400 61.200 306.200 ;
        RECT 63.600 305.600 64.600 306.400 ;
        RECT 67.600 305.600 69.200 306.400 ;
        RECT 70.000 306.200 70.800 306.400 ;
        RECT 73.800 306.200 74.600 308.600 ;
        RECT 76.400 308.200 85.200 309.000 ;
        RECT 89.000 308.400 89.600 312.200 ;
        RECT 94.200 311.600 94.800 315.000 ;
        RECT 91.000 311.000 94.800 311.600 ;
        RECT 95.600 315.000 96.400 319.000 ;
        RECT 95.600 311.600 96.200 315.000 ;
        RECT 99.800 312.800 100.600 319.800 ;
        RECT 99.800 312.200 101.400 312.800 ;
        RECT 95.600 311.000 99.400 311.600 ;
        RECT 91.000 309.000 91.600 311.000 ;
        RECT 79.800 306.800 82.800 307.600 ;
        RECT 79.800 306.200 80.600 306.800 ;
        RECT 70.000 305.600 74.600 306.200 ;
        RECT 60.400 302.200 61.200 305.400 ;
        RECT 78.000 305.400 80.600 306.200 ;
        RECT 62.000 302.200 62.800 305.000 ;
        RECT 63.600 302.200 64.400 305.000 ;
        RECT 65.200 302.200 66.000 305.000 ;
        RECT 66.800 302.200 67.600 305.000 ;
        RECT 70.000 302.200 70.800 305.000 ;
        RECT 73.200 302.200 74.000 305.000 ;
        RECT 74.800 302.200 75.600 305.000 ;
        RECT 76.400 302.200 77.200 305.000 ;
        RECT 78.000 302.200 78.800 305.400 ;
        RECT 84.400 302.200 85.200 308.200 ;
        RECT 86.000 308.300 86.800 308.400 ;
        RECT 87.600 308.300 89.600 308.400 ;
        RECT 86.000 307.700 89.600 308.300 ;
        RECT 90.200 308.200 91.600 309.000 ;
        RECT 92.400 308.800 93.200 310.400 ;
        RECT 94.000 310.300 94.800 310.400 ;
        RECT 95.600 310.300 96.400 310.400 ;
        RECT 94.000 309.700 96.400 310.300 ;
        RECT 94.000 308.800 94.800 309.700 ;
        RECT 95.600 308.800 96.400 309.700 ;
        RECT 97.200 308.800 98.000 310.400 ;
        RECT 98.800 309.000 99.400 311.000 ;
        RECT 86.000 307.600 86.800 307.700 ;
        RECT 87.600 307.600 89.600 307.700 ;
        RECT 89.000 307.000 89.600 307.600 ;
        RECT 90.600 307.800 91.600 308.200 ;
        RECT 98.800 308.200 100.200 309.000 ;
        RECT 100.800 308.400 101.400 312.200 ;
        RECT 102.000 310.300 102.800 311.200 ;
        RECT 105.200 310.300 106.000 319.800 ;
        RECT 110.000 312.000 110.800 319.800 ;
        RECT 113.200 315.200 114.000 319.800 ;
        RECT 102.000 309.700 106.000 310.300 ;
        RECT 102.000 309.600 102.800 309.700 ;
        RECT 100.800 308.300 102.800 308.400 ;
        RECT 103.600 308.300 104.400 308.400 ;
        RECT 98.800 307.800 99.800 308.200 ;
        RECT 90.600 307.200 94.800 307.800 ;
        RECT 89.000 306.600 89.800 307.000 ;
        RECT 89.000 306.000 90.600 306.600 ;
        RECT 89.800 303.000 90.600 306.000 ;
        RECT 94.200 305.000 94.800 307.200 ;
        RECT 94.000 303.000 94.800 305.000 ;
        RECT 95.600 307.200 99.800 307.800 ;
        RECT 100.800 307.700 104.400 308.300 ;
        RECT 100.800 307.600 102.800 307.700 ;
        RECT 103.600 307.600 104.400 307.700 ;
        RECT 95.600 305.000 96.200 307.200 ;
        RECT 100.800 307.000 101.400 307.600 ;
        RECT 100.600 306.600 101.400 307.000 ;
        RECT 99.800 306.000 101.400 306.600 ;
        RECT 95.600 303.000 96.400 305.000 ;
        RECT 99.800 303.000 100.600 306.000 ;
        RECT 105.200 302.200 106.000 309.700 ;
        RECT 109.800 311.200 110.800 312.000 ;
        RECT 111.400 314.600 114.000 315.200 ;
        RECT 111.400 313.000 112.000 314.600 ;
        RECT 116.400 314.400 117.200 319.800 ;
        RECT 119.600 317.000 120.400 319.800 ;
        RECT 121.200 317.000 122.000 319.800 ;
        RECT 122.800 317.000 123.600 319.800 ;
        RECT 117.800 314.400 122.000 315.200 ;
        RECT 114.600 313.600 117.200 314.400 ;
        RECT 124.400 313.600 125.200 319.800 ;
        RECT 127.600 315.000 128.400 319.800 ;
        RECT 130.800 315.000 131.600 319.800 ;
        RECT 132.400 317.000 133.200 319.800 ;
        RECT 134.000 317.000 134.800 319.800 ;
        RECT 137.200 315.200 138.000 319.800 ;
        RECT 140.400 316.400 141.200 319.800 ;
        RECT 140.400 315.800 141.400 316.400 ;
        RECT 140.800 315.200 141.400 315.800 ;
        RECT 136.000 314.400 140.200 315.200 ;
        RECT 140.800 314.600 142.800 315.200 ;
        RECT 127.600 313.600 130.200 314.400 ;
        RECT 130.800 313.800 136.600 314.400 ;
        RECT 139.600 314.000 140.200 314.400 ;
        RECT 119.600 313.000 120.400 313.200 ;
        RECT 111.400 312.400 120.400 313.000 ;
        RECT 122.800 313.000 123.600 313.200 ;
        RECT 130.800 313.000 131.400 313.800 ;
        RECT 137.200 313.200 138.600 313.800 ;
        RECT 139.600 313.200 141.200 314.000 ;
        RECT 122.800 312.400 131.400 313.000 ;
        RECT 132.400 313.000 138.600 313.200 ;
        RECT 132.400 312.600 137.800 313.000 ;
        RECT 132.400 312.400 133.200 312.600 ;
        RECT 109.800 306.800 110.600 311.200 ;
        RECT 111.400 310.600 112.000 312.400 ;
        RECT 111.200 310.000 112.000 310.600 ;
        RECT 118.000 310.000 141.400 310.600 ;
        RECT 111.200 308.000 111.800 310.000 ;
        RECT 118.000 309.400 118.800 310.000 ;
        RECT 135.600 309.600 136.400 310.000 ;
        RECT 137.200 309.600 138.000 310.000 ;
        RECT 140.600 309.800 141.400 310.000 ;
        RECT 112.400 308.600 116.200 309.400 ;
        RECT 111.200 307.400 112.400 308.000 ;
        RECT 106.800 306.300 107.600 306.400 ;
        RECT 109.800 306.300 110.800 306.800 ;
        RECT 106.800 305.700 110.800 306.300 ;
        RECT 106.800 304.800 107.600 305.700 ;
        RECT 110.000 302.200 110.800 305.700 ;
        RECT 111.600 302.200 112.400 307.400 ;
        RECT 115.400 307.400 116.200 308.600 ;
        RECT 115.400 306.800 117.200 307.400 ;
        RECT 116.400 306.200 117.200 306.800 ;
        RECT 121.200 306.400 122.000 309.200 ;
        RECT 124.400 308.600 127.600 309.400 ;
        RECT 131.400 308.600 133.400 309.400 ;
        RECT 142.000 309.000 142.800 314.600 ;
        RECT 146.200 312.600 147.000 319.800 ;
        RECT 145.200 311.800 147.000 312.600 ;
        RECT 153.200 311.800 154.000 319.800 ;
        RECT 154.800 312.400 155.600 319.800 ;
        RECT 158.000 312.400 158.800 319.800 ;
        RECT 154.800 311.800 158.800 312.400 ;
        RECT 161.200 312.000 162.000 319.800 ;
        RECT 164.400 315.200 165.200 319.800 ;
        RECT 124.000 307.800 124.800 308.000 ;
        RECT 124.000 307.200 128.400 307.800 ;
        RECT 127.600 307.000 128.400 307.200 ;
        RECT 129.200 306.800 130.000 308.400 ;
        RECT 116.400 305.400 118.800 306.200 ;
        RECT 121.200 305.600 122.200 306.400 ;
        RECT 125.200 305.600 126.800 306.400 ;
        RECT 127.600 306.200 128.400 306.400 ;
        RECT 131.400 306.200 132.200 308.600 ;
        RECT 134.000 308.200 142.800 309.000 ;
        RECT 145.400 308.400 146.000 311.800 ;
        RECT 146.800 309.600 147.600 311.200 ;
        RECT 153.400 310.400 154.000 311.800 ;
        RECT 161.000 311.200 162.000 312.000 ;
        RECT 162.600 314.600 165.200 315.200 ;
        RECT 162.600 313.000 163.200 314.600 ;
        RECT 167.600 314.400 168.400 319.800 ;
        RECT 170.800 317.000 171.600 319.800 ;
        RECT 172.400 317.000 173.200 319.800 ;
        RECT 174.000 317.000 174.800 319.800 ;
        RECT 169.000 314.400 173.200 315.200 ;
        RECT 165.800 313.600 168.400 314.400 ;
        RECT 175.600 313.600 176.400 319.800 ;
        RECT 178.800 315.000 179.600 319.800 ;
        RECT 182.000 315.000 182.800 319.800 ;
        RECT 183.600 317.000 184.400 319.800 ;
        RECT 185.200 317.000 186.000 319.800 ;
        RECT 188.400 315.200 189.200 319.800 ;
        RECT 191.600 316.400 192.400 319.800 ;
        RECT 191.600 315.800 192.600 316.400 ;
        RECT 196.400 315.800 197.200 319.800 ;
        RECT 192.000 315.200 192.600 315.800 ;
        RECT 196.600 315.600 197.200 315.800 ;
        RECT 199.600 315.800 200.400 319.800 ;
        RECT 202.800 316.400 203.600 319.800 ;
        RECT 202.600 315.800 203.600 316.400 ;
        RECT 199.600 315.600 200.200 315.800 ;
        RECT 187.200 314.400 191.400 315.200 ;
        RECT 192.000 314.600 194.000 315.200 ;
        RECT 196.600 315.000 200.200 315.600 ;
        RECT 202.600 315.200 203.200 315.800 ;
        RECT 206.000 315.200 206.800 319.800 ;
        RECT 209.200 317.000 210.000 319.800 ;
        RECT 210.800 317.000 211.600 319.800 ;
        RECT 178.800 313.600 181.400 314.400 ;
        RECT 182.000 313.800 187.800 314.400 ;
        RECT 190.800 314.000 191.400 314.400 ;
        RECT 170.800 313.000 171.600 313.200 ;
        RECT 162.600 312.400 171.600 313.000 ;
        RECT 174.000 313.000 174.800 313.200 ;
        RECT 182.000 313.000 182.600 313.800 ;
        RECT 188.400 313.200 189.800 313.800 ;
        RECT 190.800 313.200 192.400 314.000 ;
        RECT 174.000 312.400 182.600 313.000 ;
        RECT 183.600 313.000 189.800 313.200 ;
        RECT 183.600 312.600 189.000 313.000 ;
        RECT 183.600 312.400 184.400 312.600 ;
        RECT 157.200 310.400 158.000 310.800 ;
        RECT 153.200 309.800 155.600 310.400 ;
        RECT 157.200 309.800 158.800 310.400 ;
        RECT 153.200 309.600 154.000 309.800 ;
        RECT 137.400 306.800 140.400 307.600 ;
        RECT 137.400 306.200 138.200 306.800 ;
        RECT 127.600 305.600 132.200 306.200 ;
        RECT 118.000 302.200 118.800 305.400 ;
        RECT 135.600 305.400 138.200 306.200 ;
        RECT 119.600 302.200 120.400 305.000 ;
        RECT 121.200 302.200 122.000 305.000 ;
        RECT 122.800 302.200 123.600 305.000 ;
        RECT 124.400 302.200 125.200 305.000 ;
        RECT 127.600 302.200 128.400 305.000 ;
        RECT 130.800 302.200 131.600 305.000 ;
        RECT 132.400 302.200 133.200 305.000 ;
        RECT 134.000 302.200 134.800 305.000 ;
        RECT 135.600 302.200 136.400 305.400 ;
        RECT 142.000 302.200 142.800 308.200 ;
        RECT 145.200 307.600 146.000 308.400 ;
        RECT 143.600 304.800 144.400 306.400 ;
        RECT 145.400 306.300 146.000 307.600 ;
        RECT 153.200 306.300 154.000 306.400 ;
        RECT 145.300 305.700 154.000 306.300 ;
        RECT 155.000 306.200 155.600 309.800 ;
        RECT 158.000 309.600 158.800 309.800 ;
        RECT 156.400 307.600 157.200 309.200 ;
        RECT 145.400 304.200 146.000 305.700 ;
        RECT 153.200 305.600 154.000 305.700 ;
        RECT 153.400 304.800 154.200 305.600 ;
        RECT 145.200 302.200 146.000 304.200 ;
        RECT 154.800 302.200 155.600 306.200 ;
        RECT 161.000 306.800 161.800 311.200 ;
        RECT 162.600 310.600 163.200 312.400 ;
        RECT 162.400 310.000 163.200 310.600 ;
        RECT 169.200 310.000 192.600 310.600 ;
        RECT 162.400 308.000 163.000 310.000 ;
        RECT 169.200 309.400 170.000 310.000 ;
        RECT 180.400 309.600 181.200 310.000 ;
        RECT 186.800 309.600 187.600 310.000 ;
        RECT 191.600 309.800 192.600 310.000 ;
        RECT 191.600 309.600 192.400 309.800 ;
        RECT 163.600 308.600 167.400 309.400 ;
        RECT 162.400 307.400 163.600 308.000 ;
        RECT 161.000 306.000 162.000 306.800 ;
        RECT 161.200 302.200 162.000 306.000 ;
        RECT 162.800 302.200 163.600 307.400 ;
        RECT 166.600 307.400 167.400 308.600 ;
        RECT 166.600 306.800 168.400 307.400 ;
        RECT 167.600 306.200 168.400 306.800 ;
        RECT 172.400 306.400 173.200 309.200 ;
        RECT 175.600 308.600 178.800 309.400 ;
        RECT 182.600 308.600 184.600 309.400 ;
        RECT 193.200 309.000 194.000 314.600 ;
        RECT 199.600 312.400 200.200 315.000 ;
        RECT 201.200 314.600 203.200 315.200 ;
        RECT 194.800 310.800 195.600 312.400 ;
        RECT 199.600 311.600 200.400 312.400 ;
        RECT 196.400 309.600 198.000 310.400 ;
        RECT 175.200 307.800 176.000 308.000 ;
        RECT 175.200 307.200 179.600 307.800 ;
        RECT 178.800 307.000 179.600 307.200 ;
        RECT 180.400 306.800 181.200 308.400 ;
        RECT 167.600 305.400 170.000 306.200 ;
        RECT 172.400 305.600 173.400 306.400 ;
        RECT 176.400 305.600 178.000 306.400 ;
        RECT 178.800 306.200 179.600 306.400 ;
        RECT 182.600 306.200 183.400 308.600 ;
        RECT 185.200 308.200 194.000 309.000 ;
        RECT 199.600 308.400 200.200 311.600 ;
        RECT 198.600 308.200 200.200 308.400 ;
        RECT 188.600 306.800 191.600 307.600 ;
        RECT 188.600 306.200 189.400 306.800 ;
        RECT 178.800 305.600 183.400 306.200 ;
        RECT 169.200 302.200 170.000 305.400 ;
        RECT 186.800 305.400 189.400 306.200 ;
        RECT 170.800 302.200 171.600 305.000 ;
        RECT 172.400 302.200 173.200 305.000 ;
        RECT 174.000 302.200 174.800 305.000 ;
        RECT 175.600 302.200 176.400 305.000 ;
        RECT 178.800 302.200 179.600 305.000 ;
        RECT 182.000 302.200 182.800 305.000 ;
        RECT 183.600 302.200 184.400 305.000 ;
        RECT 185.200 302.200 186.000 305.000 ;
        RECT 186.800 302.200 187.600 305.400 ;
        RECT 193.200 302.200 194.000 308.200 ;
        RECT 198.400 307.800 200.200 308.200 ;
        RECT 201.200 309.000 202.000 314.600 ;
        RECT 203.800 314.400 208.000 315.200 ;
        RECT 212.400 315.000 213.200 319.800 ;
        RECT 215.600 315.000 216.400 319.800 ;
        RECT 203.800 314.000 204.400 314.400 ;
        RECT 202.800 313.200 204.400 314.000 ;
        RECT 207.400 313.800 213.200 314.400 ;
        RECT 205.400 313.200 206.800 313.800 ;
        RECT 205.400 313.000 211.600 313.200 ;
        RECT 206.200 312.600 211.600 313.000 ;
        RECT 210.800 312.400 211.600 312.600 ;
        RECT 212.600 313.000 213.200 313.800 ;
        RECT 213.800 313.600 216.400 314.400 ;
        RECT 218.800 313.600 219.600 319.800 ;
        RECT 220.400 317.000 221.200 319.800 ;
        RECT 222.000 317.000 222.800 319.800 ;
        RECT 223.600 317.000 224.400 319.800 ;
        RECT 222.000 314.400 226.200 315.200 ;
        RECT 226.800 314.400 227.600 319.800 ;
        RECT 230.000 315.200 230.800 319.800 ;
        RECT 230.000 314.600 232.600 315.200 ;
        RECT 226.800 313.600 229.400 314.400 ;
        RECT 220.400 313.000 221.200 313.200 ;
        RECT 212.600 312.400 221.200 313.000 ;
        RECT 223.600 313.000 224.400 313.200 ;
        RECT 232.000 313.000 232.600 314.600 ;
        RECT 223.600 312.400 232.600 313.000 ;
        RECT 232.000 310.600 232.600 312.400 ;
        RECT 233.200 312.000 234.000 319.800 ;
        RECT 233.200 311.200 234.200 312.000 ;
        RECT 202.600 310.000 226.000 310.600 ;
        RECT 232.000 310.000 232.800 310.600 ;
        RECT 202.600 309.800 203.400 310.000 ;
        RECT 204.400 309.600 205.200 310.000 ;
        RECT 207.600 309.600 208.400 310.000 ;
        RECT 225.200 309.400 226.000 310.000 ;
        RECT 201.200 308.200 210.000 309.000 ;
        RECT 210.600 308.600 212.600 309.400 ;
        RECT 216.400 308.600 219.600 309.400 ;
        RECT 196.400 304.300 197.200 304.400 ;
        RECT 198.400 304.300 199.200 307.800 ;
        RECT 196.400 303.700 199.200 304.300 ;
        RECT 196.400 303.600 197.200 303.700 ;
        RECT 198.400 302.200 199.200 303.700 ;
        RECT 201.200 302.200 202.000 308.200 ;
        RECT 203.600 306.800 206.600 307.600 ;
        RECT 205.800 306.200 206.600 306.800 ;
        RECT 211.800 306.200 212.600 308.600 ;
        RECT 214.000 306.800 214.800 308.400 ;
        RECT 219.200 307.800 220.000 308.000 ;
        RECT 215.600 307.200 220.000 307.800 ;
        RECT 215.600 307.000 216.400 307.200 ;
        RECT 222.000 306.400 222.800 309.200 ;
        RECT 227.800 308.600 231.600 309.400 ;
        RECT 227.800 307.400 228.600 308.600 ;
        RECT 232.200 308.000 232.800 310.000 ;
        RECT 215.600 306.200 216.400 306.400 ;
        RECT 205.800 305.400 208.400 306.200 ;
        RECT 211.800 305.600 216.400 306.200 ;
        RECT 217.200 305.600 218.800 306.400 ;
        RECT 221.800 305.600 222.800 306.400 ;
        RECT 226.800 306.800 228.600 307.400 ;
        RECT 231.600 307.400 232.800 308.000 ;
        RECT 226.800 306.200 227.600 306.800 ;
        RECT 207.600 302.200 208.400 305.400 ;
        RECT 225.200 305.400 227.600 306.200 ;
        RECT 209.200 302.200 210.000 305.000 ;
        RECT 210.800 302.200 211.600 305.000 ;
        RECT 212.400 302.200 213.200 305.000 ;
        RECT 215.600 302.200 216.400 305.000 ;
        RECT 218.800 302.200 219.600 305.000 ;
        RECT 220.400 302.200 221.200 305.000 ;
        RECT 222.000 302.200 222.800 305.000 ;
        RECT 223.600 302.200 224.400 305.000 ;
        RECT 225.200 302.200 226.000 305.400 ;
        RECT 231.600 302.200 232.400 307.400 ;
        RECT 233.400 306.800 234.200 311.200 ;
        RECT 233.200 306.000 234.200 306.800 ;
        RECT 233.200 302.200 234.000 306.000 ;
        RECT 236.400 302.200 237.200 319.800 ;
        RECT 238.000 308.300 238.800 308.400 ;
        RECT 239.600 308.300 240.400 308.400 ;
        RECT 238.000 307.700 240.400 308.300 ;
        RECT 238.000 306.800 238.800 307.700 ;
        RECT 239.600 306.800 240.400 307.700 ;
        RECT 241.200 308.300 242.000 319.800 ;
        RECT 242.800 311.600 243.600 313.200 ;
        RECT 244.400 308.300 245.200 308.400 ;
        RECT 241.200 307.700 245.200 308.300 ;
        RECT 241.200 306.200 242.000 307.700 ;
        RECT 244.400 306.800 245.200 307.700 ;
        RECT 246.000 306.200 246.800 319.800 ;
        RECT 247.600 311.600 248.400 313.200 ;
        RECT 249.200 312.400 250.000 319.800 ;
        RECT 252.400 312.800 253.200 319.800 ;
        RECT 259.400 318.400 260.200 319.800 ;
        RECT 258.800 317.600 260.200 318.400 ;
        RECT 259.400 312.800 260.200 317.600 ;
        RECT 263.600 315.000 264.400 319.000 ;
        RECT 249.200 311.800 251.800 312.400 ;
        RECT 252.400 311.800 253.400 312.800 ;
        RECT 249.200 309.600 250.200 310.400 ;
        RECT 249.400 308.800 250.200 309.600 ;
        RECT 251.200 309.800 251.800 311.800 ;
        RECT 251.200 309.000 252.200 309.800 ;
        RECT 251.200 307.400 251.800 309.000 ;
        RECT 252.800 308.400 253.400 311.800 ;
        RECT 258.600 312.200 260.200 312.800 ;
        RECT 257.200 309.600 258.000 311.200 ;
        RECT 258.600 308.400 259.200 312.200 ;
        RECT 263.800 311.600 264.400 315.000 ;
        RECT 260.600 311.000 264.400 311.600 ;
        RECT 265.200 315.000 266.000 319.000 ;
        RECT 269.400 318.400 270.200 319.800 ;
        RECT 268.400 317.600 270.200 318.400 ;
        RECT 265.200 311.600 265.800 315.000 ;
        RECT 269.400 312.800 270.200 317.600 ;
        RECT 275.600 313.600 276.400 314.400 ;
        RECT 269.400 312.200 271.000 312.800 ;
        RECT 275.600 312.400 276.200 313.600 ;
        RECT 277.000 312.400 277.800 319.800 ;
        RECT 265.200 311.000 269.000 311.600 ;
        RECT 260.600 309.000 261.200 311.000 ;
        RECT 252.400 308.300 253.400 308.400 ;
        RECT 254.000 308.300 254.800 308.400 ;
        RECT 252.400 307.700 254.800 308.300 ;
        RECT 252.400 307.600 253.400 307.700 ;
        RECT 254.000 307.600 254.800 307.700 ;
        RECT 257.200 307.600 259.200 308.400 ;
        RECT 259.800 308.200 261.200 309.000 ;
        RECT 262.000 308.800 262.800 310.400 ;
        RECT 263.600 310.300 264.400 310.400 ;
        RECT 265.200 310.300 266.000 310.400 ;
        RECT 263.600 309.700 266.000 310.300 ;
        RECT 263.600 308.800 264.400 309.700 ;
        RECT 265.200 308.800 266.000 309.700 ;
        RECT 266.800 308.800 267.600 310.400 ;
        RECT 268.400 309.000 269.000 311.000 ;
        RECT 249.200 306.800 251.800 307.400 ;
        RECT 241.200 305.600 243.000 306.200 ;
        RECT 246.000 305.600 247.800 306.200 ;
        RECT 242.200 302.200 243.000 305.600 ;
        RECT 247.000 302.200 247.800 305.600 ;
        RECT 249.200 302.200 250.000 306.800 ;
        RECT 252.800 306.200 253.400 307.600 ;
        RECT 252.400 305.600 253.400 306.200 ;
        RECT 258.600 307.000 259.200 307.600 ;
        RECT 260.200 307.800 261.200 308.200 ;
        RECT 268.400 308.200 269.800 309.000 ;
        RECT 270.400 308.400 271.000 312.200 ;
        RECT 274.800 311.800 276.200 312.400 ;
        RECT 276.800 311.800 277.800 312.400 ;
        RECT 274.800 311.600 275.600 311.800 ;
        RECT 271.600 310.300 272.400 311.200 ;
        RECT 274.800 310.300 275.600 310.400 ;
        RECT 271.600 309.700 275.600 310.300 ;
        RECT 271.600 309.600 272.400 309.700 ;
        RECT 274.800 309.600 275.600 309.700 ;
        RECT 276.800 308.400 277.400 311.800 ;
        RECT 278.000 308.800 278.800 310.400 ;
        RECT 279.600 310.300 280.400 310.400 ;
        RECT 279.600 309.700 281.900 310.300 ;
        RECT 279.600 309.600 280.400 309.700 ;
        RECT 281.300 308.400 281.900 309.700 ;
        RECT 268.400 307.800 269.400 308.200 ;
        RECT 260.200 307.200 264.400 307.800 ;
        RECT 258.600 306.600 259.400 307.000 ;
        RECT 258.600 306.000 260.200 306.600 ;
        RECT 252.400 302.200 253.200 305.600 ;
        RECT 259.400 303.000 260.200 306.000 ;
        RECT 263.800 305.000 264.400 307.200 ;
        RECT 263.600 303.000 264.400 305.000 ;
        RECT 265.200 307.200 269.400 307.800 ;
        RECT 270.400 307.600 272.400 308.400 ;
        RECT 273.200 308.300 274.000 308.400 ;
        RECT 274.800 308.300 277.400 308.400 ;
        RECT 273.200 307.700 277.400 308.300 ;
        RECT 279.600 308.200 280.400 308.400 ;
        RECT 273.200 307.600 274.000 307.700 ;
        RECT 274.800 307.600 277.400 307.700 ;
        RECT 278.800 307.600 280.400 308.200 ;
        RECT 265.200 305.000 265.800 307.200 ;
        RECT 270.400 307.000 271.000 307.600 ;
        RECT 270.200 306.600 271.000 307.000 ;
        RECT 269.400 306.000 271.000 306.600 ;
        RECT 275.000 306.200 275.600 307.600 ;
        RECT 278.800 307.200 279.600 307.600 ;
        RECT 281.200 306.800 282.000 308.400 ;
        RECT 276.600 306.200 280.200 306.600 ;
        RECT 282.800 306.200 283.600 319.800 ;
        RECT 284.400 311.600 285.200 313.200 ;
        RECT 284.400 310.300 285.200 310.400 ;
        RECT 286.000 310.300 286.800 319.800 ;
        RECT 284.400 309.700 286.800 310.300 ;
        RECT 284.400 309.600 285.200 309.700 ;
        RECT 265.200 303.000 266.000 305.000 ;
        RECT 269.400 303.000 270.200 306.000 ;
        RECT 274.800 302.200 275.600 306.200 ;
        RECT 276.400 306.000 280.400 306.200 ;
        RECT 276.400 302.200 277.200 306.000 ;
        RECT 279.600 302.200 280.400 306.000 ;
        RECT 282.800 305.600 284.600 306.200 ;
        RECT 283.800 302.200 284.600 305.600 ;
        RECT 286.000 302.200 286.800 309.700 ;
        RECT 289.200 310.300 290.000 319.800 ;
        RECT 298.800 312.000 299.600 319.800 ;
        RECT 302.000 315.200 302.800 319.800 ;
        RECT 298.600 311.200 299.600 312.000 ;
        RECT 300.200 314.600 302.800 315.200 ;
        RECT 300.200 313.000 300.800 314.600 ;
        RECT 305.200 314.400 306.000 319.800 ;
        RECT 308.400 317.000 309.200 319.800 ;
        RECT 310.000 317.000 310.800 319.800 ;
        RECT 311.600 317.000 312.400 319.800 ;
        RECT 306.600 314.400 310.800 315.200 ;
        RECT 303.400 313.600 306.000 314.400 ;
        RECT 313.200 313.600 314.000 319.800 ;
        RECT 316.400 315.000 317.200 319.800 ;
        RECT 319.600 315.000 320.400 319.800 ;
        RECT 321.200 317.000 322.000 319.800 ;
        RECT 322.800 317.000 323.600 319.800 ;
        RECT 326.000 315.200 326.800 319.800 ;
        RECT 329.200 316.400 330.000 319.800 ;
        RECT 329.200 315.800 330.200 316.400 ;
        RECT 329.600 315.200 330.200 315.800 ;
        RECT 324.800 314.400 329.000 315.200 ;
        RECT 329.600 314.600 331.600 315.200 ;
        RECT 316.400 313.600 319.000 314.400 ;
        RECT 319.600 313.800 325.400 314.400 ;
        RECT 328.400 314.000 329.000 314.400 ;
        RECT 308.400 313.000 309.200 313.200 ;
        RECT 300.200 312.400 309.200 313.000 ;
        RECT 311.600 313.000 312.400 313.200 ;
        RECT 319.600 313.000 320.200 313.800 ;
        RECT 326.000 313.200 327.400 313.800 ;
        RECT 328.400 313.200 330.000 314.000 ;
        RECT 311.600 312.400 320.200 313.000 ;
        RECT 321.200 313.000 327.400 313.200 ;
        RECT 321.200 312.600 326.600 313.000 ;
        RECT 321.200 312.400 322.000 312.600 ;
        RECT 292.400 310.300 293.200 310.400 ;
        RECT 289.200 309.700 293.200 310.300 ;
        RECT 287.600 306.800 288.400 308.400 ;
        RECT 289.200 302.200 290.000 309.700 ;
        RECT 292.400 309.600 293.200 309.700 ;
        RECT 290.800 308.300 291.600 308.400 ;
        RECT 294.000 308.300 294.800 308.400 ;
        RECT 290.800 307.700 294.800 308.300 ;
        RECT 290.800 306.800 291.600 307.700 ;
        RECT 294.000 307.600 294.800 307.700 ;
        RECT 298.600 306.800 299.400 311.200 ;
        RECT 300.200 310.600 300.800 312.400 ;
        RECT 300.000 310.000 300.800 310.600 ;
        RECT 306.800 310.000 330.200 310.600 ;
        RECT 300.000 308.000 300.600 310.000 ;
        RECT 306.800 309.400 307.600 310.000 ;
        RECT 324.400 309.600 325.200 310.000 ;
        RECT 329.400 309.800 330.200 310.000 ;
        RECT 301.200 308.600 305.000 309.400 ;
        RECT 300.000 307.400 301.200 308.000 ;
        RECT 298.600 306.000 299.600 306.800 ;
        RECT 298.800 302.200 299.600 306.000 ;
        RECT 300.400 302.200 301.200 307.400 ;
        RECT 304.200 307.400 305.000 308.600 ;
        RECT 304.200 306.800 306.000 307.400 ;
        RECT 305.200 306.200 306.000 306.800 ;
        RECT 310.000 306.400 310.800 309.200 ;
        RECT 313.200 308.600 316.400 309.400 ;
        RECT 320.200 308.600 322.200 309.400 ;
        RECT 330.800 309.000 331.600 314.600 ;
        RECT 312.800 307.800 313.600 308.000 ;
        RECT 312.800 307.200 317.200 307.800 ;
        RECT 316.400 307.000 317.200 307.200 ;
        RECT 318.000 306.800 318.800 308.400 ;
        RECT 305.200 305.400 307.600 306.200 ;
        RECT 310.000 305.600 311.000 306.400 ;
        RECT 314.000 305.600 315.600 306.400 ;
        RECT 316.400 306.200 317.200 306.400 ;
        RECT 320.200 306.200 321.000 308.600 ;
        RECT 322.800 308.200 331.600 309.000 ;
        RECT 326.200 306.800 329.200 307.600 ;
        RECT 326.200 306.200 327.000 306.800 ;
        RECT 316.400 305.600 321.000 306.200 ;
        RECT 306.800 302.200 307.600 305.400 ;
        RECT 324.400 305.400 327.000 306.200 ;
        RECT 308.400 302.200 309.200 305.000 ;
        RECT 310.000 302.200 310.800 305.000 ;
        RECT 311.600 302.200 312.400 305.000 ;
        RECT 313.200 302.200 314.000 305.000 ;
        RECT 316.400 302.200 317.200 305.000 ;
        RECT 319.600 302.200 320.400 305.000 ;
        RECT 321.200 302.200 322.000 305.000 ;
        RECT 322.800 302.200 323.600 305.000 ;
        RECT 324.400 302.200 325.200 305.400 ;
        RECT 330.800 302.200 331.600 308.200 ;
        RECT 332.400 306.800 333.200 308.400 ;
        RECT 334.000 308.300 334.800 319.800 ;
        RECT 335.600 312.300 336.400 313.200 ;
        RECT 337.200 312.300 338.000 312.400 ;
        RECT 335.600 311.700 338.000 312.300 ;
        RECT 335.600 311.600 336.400 311.700 ;
        RECT 337.200 311.600 338.000 311.700 ;
        RECT 337.200 308.300 338.000 308.400 ;
        RECT 334.000 307.700 338.000 308.300 ;
        RECT 334.000 306.200 334.800 307.700 ;
        RECT 337.200 306.800 338.000 307.700 ;
        RECT 338.800 306.200 339.600 319.800 ;
        RECT 342.800 313.600 343.600 314.400 ;
        RECT 340.400 311.600 341.200 313.200 ;
        RECT 342.800 312.400 343.400 313.600 ;
        RECT 344.200 312.400 345.000 319.800 ;
        RECT 349.200 313.600 350.000 314.400 ;
        RECT 349.200 312.400 349.800 313.600 ;
        RECT 350.600 312.400 351.400 319.800 ;
        RECT 342.000 311.800 343.400 312.400 ;
        RECT 344.000 311.800 345.000 312.400 ;
        RECT 348.400 311.800 349.800 312.400 ;
        RECT 350.400 311.800 351.400 312.400 ;
        RECT 342.000 311.600 342.800 311.800 ;
        RECT 340.500 310.300 341.100 311.600 ;
        RECT 344.000 310.300 344.600 311.800 ;
        RECT 348.400 311.600 349.200 311.800 ;
        RECT 340.500 309.700 344.600 310.300 ;
        RECT 344.000 308.400 344.600 309.700 ;
        RECT 345.200 310.300 346.000 310.400 ;
        RECT 350.400 310.300 351.000 311.800 ;
        RECT 345.200 309.700 351.000 310.300 ;
        RECT 345.200 308.800 346.000 309.700 ;
        RECT 350.400 308.400 351.000 309.700 ;
        RECT 351.600 308.800 352.400 310.400 ;
        RECT 342.000 307.600 344.600 308.400 ;
        RECT 346.800 308.200 347.600 308.400 ;
        RECT 346.000 307.600 347.600 308.200 ;
        RECT 348.400 307.600 351.000 308.400 ;
        RECT 353.200 308.300 354.000 308.400 ;
        RECT 354.800 308.300 355.600 319.800 ;
        RECT 359.600 315.800 360.400 319.800 ;
        RECT 359.800 315.600 360.400 315.800 ;
        RECT 362.800 315.800 363.600 319.800 ;
        RECT 362.800 315.600 363.400 315.800 ;
        RECT 359.800 315.000 363.400 315.600 ;
        RECT 358.000 314.300 358.800 314.400 ;
        RECT 361.200 314.300 362.000 314.400 ;
        RECT 358.000 313.700 362.000 314.300 ;
        RECT 358.000 313.600 358.800 313.700 ;
        RECT 361.200 312.800 362.000 313.700 ;
        RECT 362.800 312.400 363.400 315.000 ;
        RECT 362.800 311.600 363.600 312.400 ;
        RECT 359.600 309.600 361.200 310.400 ;
        RECT 362.800 308.400 363.400 311.600 ;
        RECT 364.400 310.300 365.200 310.400 ;
        RECT 366.000 310.300 366.800 319.800 ;
        RECT 370.800 315.600 371.600 319.800 ;
        RECT 374.000 315.800 374.800 319.800 ;
        RECT 375.600 319.200 379.600 319.800 ;
        RECT 374.000 315.600 374.600 315.800 ;
        RECT 371.000 315.000 374.600 315.600 ;
        RECT 372.400 312.800 373.200 314.400 ;
        RECT 374.000 312.400 374.600 315.000 ;
        RECT 374.000 311.600 374.800 312.400 ;
        RECT 375.600 311.800 376.400 319.200 ;
        RECT 377.200 311.800 378.000 318.600 ;
        RECT 378.800 312.400 379.600 319.200 ;
        RECT 382.000 312.400 382.800 319.800 ;
        RECT 378.800 311.800 382.800 312.400 ;
        RECT 364.400 309.700 366.800 310.300 ;
        RECT 364.400 309.600 365.200 309.700 ;
        RECT 353.200 308.200 355.600 308.300 ;
        RECT 361.800 308.200 363.400 308.400 ;
        RECT 352.400 307.700 355.600 308.200 ;
        RECT 352.400 307.600 354.000 307.700 ;
        RECT 342.200 306.200 342.800 307.600 ;
        RECT 346.000 307.200 346.800 307.600 ;
        RECT 343.800 306.200 347.400 306.600 ;
        RECT 348.600 306.200 349.200 307.600 ;
        RECT 352.400 307.200 353.200 307.600 ;
        RECT 350.200 306.200 353.800 306.600 ;
        RECT 334.000 305.600 335.800 306.200 ;
        RECT 338.800 305.600 340.600 306.200 ;
        RECT 335.000 302.200 335.800 305.600 ;
        RECT 339.800 304.400 340.600 305.600 ;
        RECT 338.800 303.600 340.600 304.400 ;
        RECT 339.800 302.200 340.600 303.600 ;
        RECT 342.000 302.200 342.800 306.200 ;
        RECT 343.600 306.000 347.600 306.200 ;
        RECT 343.600 302.200 344.400 306.000 ;
        RECT 346.800 302.200 347.600 306.000 ;
        RECT 348.400 302.200 349.200 306.200 ;
        RECT 350.000 306.000 354.000 306.200 ;
        RECT 350.000 302.200 350.800 306.000 ;
        RECT 353.200 302.200 354.000 306.000 ;
        RECT 354.800 302.200 355.600 307.700 ;
        RECT 361.600 307.800 363.400 308.200 ;
        RECT 356.400 304.800 357.200 306.400 ;
        RECT 359.600 304.300 360.400 304.400 ;
        RECT 361.600 304.300 362.400 307.800 ;
        RECT 359.600 303.700 362.400 304.300 ;
        RECT 359.600 303.600 360.400 303.700 ;
        RECT 361.600 302.200 362.400 303.700 ;
        RECT 366.000 302.200 366.800 309.700 ;
        RECT 370.800 309.600 372.400 310.400 ;
        RECT 374.000 308.400 374.600 311.600 ;
        RECT 377.400 311.200 378.000 311.800 ;
        RECT 375.600 309.600 376.400 311.200 ;
        RECT 377.400 310.600 379.400 311.200 ;
        RECT 378.800 310.400 379.400 310.600 ;
        RECT 381.200 310.400 382.000 310.800 ;
        RECT 378.800 309.600 379.600 310.400 ;
        RECT 381.200 309.800 382.800 310.400 ;
        RECT 382.000 309.600 382.800 309.800 ;
        RECT 377.400 308.800 378.200 309.600 ;
        RECT 377.400 308.400 378.000 308.800 ;
        RECT 373.000 308.200 374.600 308.400 ;
        RECT 372.800 307.800 374.600 308.200 ;
        RECT 372.800 302.200 373.600 307.800 ;
        RECT 377.200 307.600 378.000 308.400 ;
        RECT 378.800 306.200 379.400 309.600 ;
        RECT 380.400 307.600 381.200 309.200 ;
        RECT 383.600 306.800 384.400 308.400 ;
        RECT 385.200 306.200 386.000 319.800 ;
        RECT 386.800 311.600 387.600 313.200 ;
        RECT 388.400 312.400 389.200 319.800 ;
        RECT 391.600 319.200 395.600 319.800 ;
        RECT 391.600 312.400 392.400 319.200 ;
        RECT 388.400 311.800 392.400 312.400 ;
        RECT 393.200 311.800 394.000 318.600 ;
        RECT 394.800 311.800 395.600 319.200 ;
        RECT 399.000 312.400 399.800 319.800 ;
        RECT 400.400 313.600 401.200 314.400 ;
        RECT 400.600 312.400 401.200 313.600 ;
        RECT 405.400 312.400 406.200 319.800 ;
        RECT 406.800 313.600 407.600 314.400 ;
        RECT 407.000 312.400 407.600 313.600 ;
        RECT 399.000 311.800 400.000 312.400 ;
        RECT 400.600 311.800 402.000 312.400 ;
        RECT 405.400 311.800 406.400 312.400 ;
        RECT 407.000 311.800 408.400 312.400 ;
        RECT 393.200 311.200 393.800 311.800 ;
        RECT 389.200 310.400 390.000 310.800 ;
        RECT 391.800 310.600 393.800 311.200 ;
        RECT 391.800 310.400 392.400 310.600 ;
        RECT 388.400 309.800 390.000 310.400 ;
        RECT 388.400 309.600 389.200 309.800 ;
        RECT 391.600 309.600 392.400 310.400 ;
        RECT 394.800 309.600 395.600 311.200 ;
        RECT 390.000 307.600 390.800 309.200 ;
        RECT 391.800 306.200 392.400 309.600 ;
        RECT 393.000 308.800 393.800 309.600 ;
        RECT 398.000 308.800 398.800 310.400 ;
        RECT 399.400 310.300 400.000 311.800 ;
        RECT 401.200 311.600 402.000 311.800 ;
        RECT 402.800 310.300 403.600 310.400 ;
        RECT 399.400 309.700 403.600 310.300 ;
        RECT 393.200 308.400 393.800 308.800 ;
        RECT 399.400 308.400 400.000 309.700 ;
        RECT 402.800 309.600 403.600 309.700 ;
        RECT 404.400 308.800 405.200 310.400 ;
        RECT 405.800 310.300 406.400 311.800 ;
        RECT 407.600 311.600 408.400 311.800 ;
        RECT 407.600 310.300 408.400 310.400 ;
        RECT 405.800 309.700 408.400 310.300 ;
        RECT 405.800 308.400 406.400 309.700 ;
        RECT 407.600 309.600 408.400 309.700 ;
        RECT 393.200 307.600 394.000 308.400 ;
        RECT 396.400 308.200 397.200 308.400 ;
        RECT 396.400 307.600 398.000 308.200 ;
        RECT 399.400 307.600 402.000 308.400 ;
        RECT 402.800 308.200 403.600 308.400 ;
        RECT 402.800 307.600 404.400 308.200 ;
        RECT 405.800 307.600 408.400 308.400 ;
        RECT 397.200 307.200 398.000 307.600 ;
        RECT 396.600 306.200 400.200 306.600 ;
        RECT 401.200 306.200 401.800 307.600 ;
        RECT 403.600 307.200 404.400 307.600 ;
        RECT 403.000 306.200 406.600 306.600 ;
        RECT 407.600 306.200 408.200 307.600 ;
        RECT 378.200 302.200 379.800 306.200 ;
        RECT 385.200 305.600 387.000 306.200 ;
        RECT 386.200 302.200 387.000 305.600 ;
        RECT 391.400 304.400 393.000 306.200 ;
        RECT 396.400 306.000 400.400 306.200 ;
        RECT 391.400 303.600 394.000 304.400 ;
        RECT 391.400 302.200 393.000 303.600 ;
        RECT 396.400 302.200 397.200 306.000 ;
        RECT 399.600 302.200 400.400 306.000 ;
        RECT 401.200 302.200 402.000 306.200 ;
        RECT 402.800 306.000 406.800 306.200 ;
        RECT 402.800 302.200 403.600 306.000 ;
        RECT 406.000 302.200 406.800 306.000 ;
        RECT 407.600 302.200 408.400 306.200 ;
        RECT 409.200 302.200 410.000 319.800 ;
        RECT 413.200 313.600 414.000 314.400 ;
        RECT 413.200 312.400 413.800 313.600 ;
        RECT 414.600 312.400 415.400 319.800 ;
        RECT 412.400 311.800 413.800 312.400 ;
        RECT 414.400 311.800 415.400 312.400 ;
        RECT 421.400 312.400 422.200 319.800 ;
        RECT 426.800 316.400 427.600 319.800 ;
        RECT 426.600 315.800 427.600 316.400 ;
        RECT 426.600 315.200 427.200 315.800 ;
        RECT 430.000 315.200 430.800 319.800 ;
        RECT 433.200 317.000 434.000 319.800 ;
        RECT 434.800 317.000 435.600 319.800 ;
        RECT 425.200 314.600 427.200 315.200 ;
        RECT 422.800 313.600 423.600 314.400 ;
        RECT 423.000 312.400 423.600 313.600 ;
        RECT 421.400 311.800 422.400 312.400 ;
        RECT 423.000 311.800 424.400 312.400 ;
        RECT 412.400 311.600 413.200 311.800 ;
        RECT 414.400 308.400 415.000 311.800 ;
        RECT 415.600 308.800 416.400 310.400 ;
        RECT 420.400 308.800 421.200 310.400 ;
        RECT 421.800 310.300 422.400 311.800 ;
        RECT 423.600 311.600 424.400 311.800 ;
        RECT 423.600 310.300 424.400 310.400 ;
        RECT 421.800 309.700 424.400 310.300 ;
        RECT 421.800 308.400 422.400 309.700 ;
        RECT 423.600 309.600 424.400 309.700 ;
        RECT 425.200 309.000 426.000 314.600 ;
        RECT 427.800 314.400 432.000 315.200 ;
        RECT 436.400 315.000 437.200 319.800 ;
        RECT 439.600 315.000 440.400 319.800 ;
        RECT 427.800 314.000 428.400 314.400 ;
        RECT 426.800 313.200 428.400 314.000 ;
        RECT 431.400 313.800 437.200 314.400 ;
        RECT 429.400 313.200 430.800 313.800 ;
        RECT 429.400 313.000 435.600 313.200 ;
        RECT 430.200 312.600 435.600 313.000 ;
        RECT 434.800 312.400 435.600 312.600 ;
        RECT 436.600 313.000 437.200 313.800 ;
        RECT 437.800 313.600 440.400 314.400 ;
        RECT 442.800 313.600 443.600 319.800 ;
        RECT 444.400 317.000 445.200 319.800 ;
        RECT 446.000 317.000 446.800 319.800 ;
        RECT 447.600 317.000 448.400 319.800 ;
        RECT 446.000 314.400 450.200 315.200 ;
        RECT 450.800 314.400 451.600 319.800 ;
        RECT 454.000 315.200 454.800 319.800 ;
        RECT 454.000 314.600 456.600 315.200 ;
        RECT 450.800 313.600 453.400 314.400 ;
        RECT 444.400 313.000 445.200 313.200 ;
        RECT 436.600 312.400 445.200 313.000 ;
        RECT 447.600 313.000 448.400 313.200 ;
        RECT 456.000 313.000 456.600 314.600 ;
        RECT 447.600 312.400 456.600 313.000 ;
        RECT 456.000 310.600 456.600 312.400 ;
        RECT 457.200 312.000 458.000 319.800 ;
        RECT 467.800 312.400 468.600 319.800 ;
        RECT 469.200 313.600 470.000 314.400 ;
        RECT 469.400 312.400 470.000 313.600 ;
        RECT 457.200 311.200 458.200 312.000 ;
        RECT 467.800 311.800 468.800 312.400 ;
        RECT 469.400 312.300 470.800 312.400 ;
        RECT 471.600 312.300 472.400 312.400 ;
        RECT 469.400 311.800 472.400 312.300 ;
        RECT 426.600 310.000 450.000 310.600 ;
        RECT 456.000 310.000 456.800 310.600 ;
        RECT 426.600 309.800 427.400 310.000 ;
        RECT 428.400 309.600 429.200 310.000 ;
        RECT 431.600 309.600 432.400 310.000 ;
        RECT 449.200 309.400 450.000 310.000 ;
        RECT 412.400 307.600 415.000 308.400 ;
        RECT 417.200 308.200 418.000 308.400 ;
        RECT 416.400 307.600 418.000 308.200 ;
        RECT 418.800 308.200 419.600 308.400 ;
        RECT 418.800 307.600 420.400 308.200 ;
        RECT 421.800 307.600 424.400 308.400 ;
        RECT 425.200 308.200 434.000 309.000 ;
        RECT 434.600 308.600 436.600 309.400 ;
        RECT 440.400 308.600 443.600 309.400 ;
        RECT 410.800 304.800 411.600 306.400 ;
        RECT 412.600 306.200 413.200 307.600 ;
        RECT 416.400 307.200 417.200 307.600 ;
        RECT 419.600 307.200 420.400 307.600 ;
        RECT 414.200 306.200 417.800 306.600 ;
        RECT 419.000 306.200 422.600 306.600 ;
        RECT 423.600 306.200 424.200 307.600 ;
        RECT 412.400 302.200 413.200 306.200 ;
        RECT 414.000 306.000 418.000 306.200 ;
        RECT 414.000 302.200 414.800 306.000 ;
        RECT 417.200 302.200 418.000 306.000 ;
        RECT 418.800 306.000 422.800 306.200 ;
        RECT 418.800 302.200 419.600 306.000 ;
        RECT 422.000 302.200 422.800 306.000 ;
        RECT 423.600 302.200 424.400 306.200 ;
        RECT 425.200 302.200 426.000 308.200 ;
        RECT 427.600 306.800 430.600 307.600 ;
        RECT 429.800 306.200 430.600 306.800 ;
        RECT 435.800 306.200 436.600 308.600 ;
        RECT 438.000 306.800 438.800 308.400 ;
        RECT 443.200 307.800 444.000 308.000 ;
        RECT 439.600 307.200 444.000 307.800 ;
        RECT 439.600 307.000 440.400 307.200 ;
        RECT 446.000 306.400 446.800 309.200 ;
        RECT 451.800 308.600 455.600 309.400 ;
        RECT 451.800 307.400 452.600 308.600 ;
        RECT 456.200 308.000 456.800 310.000 ;
        RECT 439.600 306.200 440.400 306.400 ;
        RECT 429.800 305.400 432.400 306.200 ;
        RECT 435.800 305.600 440.400 306.200 ;
        RECT 441.200 305.600 442.800 306.400 ;
        RECT 445.800 305.600 446.800 306.400 ;
        RECT 450.800 306.800 452.600 307.400 ;
        RECT 455.600 307.400 456.800 308.000 ;
        RECT 450.800 306.200 451.600 306.800 ;
        RECT 431.600 302.200 432.400 305.400 ;
        RECT 449.200 305.400 451.600 306.200 ;
        RECT 433.200 302.200 434.000 305.000 ;
        RECT 434.800 302.200 435.600 305.000 ;
        RECT 436.400 302.200 437.200 305.000 ;
        RECT 439.600 302.200 440.400 305.000 ;
        RECT 442.800 302.200 443.600 305.000 ;
        RECT 444.400 302.200 445.200 305.000 ;
        RECT 446.000 302.200 446.800 305.000 ;
        RECT 447.600 302.200 448.400 305.000 ;
        RECT 449.200 302.200 450.000 305.400 ;
        RECT 455.600 302.200 456.400 307.400 ;
        RECT 457.400 306.800 458.200 311.200 ;
        RECT 466.800 308.800 467.600 310.400 ;
        RECT 468.200 310.300 468.800 311.800 ;
        RECT 470.000 311.700 472.400 311.800 ;
        RECT 470.000 311.600 470.800 311.700 ;
        RECT 471.600 311.600 472.400 311.700 ;
        RECT 471.600 310.300 472.400 310.400 ;
        RECT 468.200 309.700 472.400 310.300 ;
        RECT 468.200 308.400 468.800 309.700 ;
        RECT 471.600 309.600 472.400 309.700 ;
        RECT 465.200 308.200 466.000 308.400 ;
        RECT 465.200 307.600 466.800 308.200 ;
        RECT 468.200 307.600 470.800 308.400 ;
        RECT 473.200 308.300 474.000 319.800 ;
        RECT 477.400 312.400 478.200 319.800 ;
        RECT 478.800 313.600 479.600 314.400 ;
        RECT 479.000 312.400 479.600 313.600 ;
        RECT 482.000 313.600 482.800 314.400 ;
        RECT 482.000 312.400 482.600 313.600 ;
        RECT 483.400 312.400 484.200 319.800 ;
        RECT 488.400 313.600 489.200 314.400 ;
        RECT 488.400 312.400 489.000 313.600 ;
        RECT 489.800 312.400 490.600 319.800 ;
        RECT 477.400 311.800 478.400 312.400 ;
        RECT 479.000 311.800 480.400 312.400 ;
        RECT 476.400 308.800 477.200 310.400 ;
        RECT 477.800 308.400 478.400 311.800 ;
        RECT 479.600 311.600 480.400 311.800 ;
        RECT 481.200 311.800 482.600 312.400 ;
        RECT 483.200 311.800 484.200 312.400 ;
        RECT 487.600 311.800 489.000 312.400 ;
        RECT 489.600 311.800 490.600 312.400 ;
        RECT 494.000 311.800 494.800 319.800 ;
        RECT 495.600 312.400 496.400 319.800 ;
        RECT 498.800 312.400 499.600 319.800 ;
        RECT 503.000 314.400 503.800 319.800 ;
        RECT 509.400 314.400 510.200 319.800 ;
        RECT 502.000 313.600 503.800 314.400 ;
        RECT 504.400 313.600 505.200 314.400 ;
        RECT 508.400 313.600 510.200 314.400 ;
        RECT 510.800 313.600 511.600 314.400 ;
        RECT 495.600 311.800 499.600 312.400 ;
        RECT 503.000 312.400 503.800 313.600 ;
        RECT 504.600 312.400 505.200 313.600 ;
        RECT 509.400 312.400 510.200 313.600 ;
        RECT 511.000 312.400 511.600 313.600 ;
        RECT 503.000 311.800 504.000 312.400 ;
        RECT 504.600 311.800 506.000 312.400 ;
        RECT 509.400 311.800 510.400 312.400 ;
        RECT 511.000 311.800 512.400 312.400 ;
        RECT 481.200 311.600 482.000 311.800 ;
        RECT 483.200 308.400 483.800 311.800 ;
        RECT 487.600 311.600 488.400 311.800 ;
        RECT 484.400 308.800 485.200 310.400 ;
        RECT 489.600 308.400 490.200 311.800 ;
        RECT 494.200 310.400 494.800 311.800 ;
        RECT 498.000 310.400 498.800 310.800 ;
        RECT 490.800 310.300 491.600 310.400 ;
        RECT 494.000 310.300 496.400 310.400 ;
        RECT 490.800 309.800 496.400 310.300 ;
        RECT 498.000 310.300 499.600 310.400 ;
        RECT 500.400 310.300 501.200 310.400 ;
        RECT 498.000 309.800 501.200 310.300 ;
        RECT 490.800 309.700 494.800 309.800 ;
        RECT 490.800 308.800 491.600 309.700 ;
        RECT 494.000 309.600 494.800 309.700 ;
        RECT 474.800 308.300 475.600 308.400 ;
        RECT 473.200 308.200 475.600 308.300 ;
        RECT 473.200 307.700 476.400 308.200 ;
        RECT 466.000 307.200 466.800 307.600 ;
        RECT 457.200 306.000 458.200 306.800 ;
        RECT 465.400 306.200 469.000 306.600 ;
        RECT 470.000 306.200 470.600 307.600 ;
        RECT 465.200 306.000 469.200 306.200 ;
        RECT 457.200 302.200 458.000 306.000 ;
        RECT 465.200 302.200 466.000 306.000 ;
        RECT 468.400 302.200 469.200 306.000 ;
        RECT 470.000 302.200 470.800 306.200 ;
        RECT 471.600 304.800 472.400 306.400 ;
        RECT 473.200 302.200 474.000 307.700 ;
        RECT 474.800 307.600 476.400 307.700 ;
        RECT 477.800 307.600 480.400 308.400 ;
        RECT 481.200 307.600 483.800 308.400 ;
        RECT 486.000 308.200 486.800 308.400 ;
        RECT 485.200 307.600 486.800 308.200 ;
        RECT 487.600 307.600 490.200 308.400 ;
        RECT 492.400 308.200 493.200 308.400 ;
        RECT 491.600 307.600 493.200 308.200 ;
        RECT 475.600 307.200 476.400 307.600 ;
        RECT 475.000 306.200 478.600 306.600 ;
        RECT 479.600 306.400 480.200 307.600 ;
        RECT 474.800 306.000 478.800 306.200 ;
        RECT 474.800 302.200 475.600 306.000 ;
        RECT 478.000 302.200 478.800 306.000 ;
        RECT 479.600 302.200 480.400 306.400 ;
        RECT 481.400 306.200 482.000 307.600 ;
        RECT 485.200 307.200 486.000 307.600 ;
        RECT 483.000 306.200 486.600 306.600 ;
        RECT 487.800 306.200 488.400 307.600 ;
        RECT 491.600 307.200 492.400 307.600 ;
        RECT 489.400 306.200 493.000 306.600 ;
        RECT 481.200 302.200 482.000 306.200 ;
        RECT 482.800 306.000 486.800 306.200 ;
        RECT 482.800 302.200 483.600 306.000 ;
        RECT 486.000 302.200 486.800 306.000 ;
        RECT 487.600 302.200 488.400 306.200 ;
        RECT 489.200 306.000 493.200 306.200 ;
        RECT 489.200 302.200 490.000 306.000 ;
        RECT 492.400 302.200 493.200 306.000 ;
        RECT 494.000 305.600 494.800 306.400 ;
        RECT 495.800 306.200 496.400 309.800 ;
        RECT 498.800 309.700 501.200 309.800 ;
        RECT 498.800 309.600 499.600 309.700 ;
        RECT 500.400 309.600 501.200 309.700 ;
        RECT 497.200 307.600 498.000 309.200 ;
        RECT 502.000 308.800 502.800 310.400 ;
        RECT 503.400 308.400 504.000 311.800 ;
        RECT 505.200 311.600 506.000 311.800 ;
        RECT 508.400 308.800 509.200 310.400 ;
        RECT 509.800 308.400 510.400 311.800 ;
        RECT 511.600 311.600 512.400 311.800 ;
        RECT 513.200 311.600 514.000 313.200 ;
        RECT 511.600 310.300 512.400 310.400 ;
        RECT 514.800 310.300 515.600 319.800 ;
        RECT 518.000 311.600 518.800 313.200 ;
        RECT 511.600 309.700 515.600 310.300 ;
        RECT 511.600 309.600 512.400 309.700 ;
        RECT 500.400 308.200 501.200 308.400 ;
        RECT 500.400 307.600 502.000 308.200 ;
        RECT 503.400 307.600 506.000 308.400 ;
        RECT 506.800 308.200 507.600 308.400 ;
        RECT 506.800 307.600 508.400 308.200 ;
        RECT 509.800 307.600 512.400 308.400 ;
        RECT 501.200 307.200 502.000 307.600 ;
        RECT 500.600 306.200 504.200 306.600 ;
        RECT 505.200 306.200 505.800 307.600 ;
        RECT 507.600 307.200 508.400 307.600 ;
        RECT 507.000 306.200 510.600 306.600 ;
        RECT 511.600 306.200 512.200 307.600 ;
        RECT 514.800 306.200 515.600 309.700 ;
        RECT 516.400 306.800 517.200 308.400 ;
        RECT 519.600 306.200 520.400 319.800 ;
        RECT 525.000 318.400 525.800 319.800 ;
        RECT 525.000 317.600 526.800 318.400 ;
        RECT 521.200 314.300 522.000 314.400 ;
        RECT 523.600 314.300 524.400 314.400 ;
        RECT 521.200 313.700 524.400 314.300 ;
        RECT 521.200 313.600 522.000 313.700 ;
        RECT 523.600 313.600 524.400 313.700 ;
        RECT 523.600 312.400 524.200 313.600 ;
        RECT 525.000 312.400 525.800 317.600 ;
        RECT 522.800 311.800 524.200 312.400 ;
        RECT 524.800 311.800 525.800 312.400 ;
        RECT 529.200 312.400 530.000 319.800 ;
        RECT 529.200 311.800 531.400 312.400 ;
        RECT 532.400 311.800 533.200 319.800 ;
        RECT 522.800 311.600 523.600 311.800 ;
        RECT 524.800 308.400 525.400 311.800 ;
        RECT 530.800 311.200 531.400 311.800 ;
        RECT 530.800 310.400 532.000 311.200 ;
        RECT 526.000 308.800 526.800 310.400 ;
        RECT 529.200 308.800 530.000 310.400 ;
        RECT 521.200 306.800 522.000 308.400 ;
        RECT 522.800 307.600 525.400 308.400 ;
        RECT 527.600 308.200 528.400 308.400 ;
        RECT 526.800 307.600 528.400 308.200 ;
        RECT 523.000 306.200 523.600 307.600 ;
        RECT 526.800 307.200 527.600 307.600 ;
        RECT 530.800 307.400 531.400 310.400 ;
        RECT 532.600 309.600 533.200 311.800 ;
        RECT 529.200 306.800 531.400 307.400 ;
        RECT 524.600 306.200 528.200 306.600 ;
        RECT 494.200 304.800 495.000 305.600 ;
        RECT 495.600 302.200 496.400 306.200 ;
        RECT 500.400 306.000 504.400 306.200 ;
        RECT 500.400 302.200 501.200 306.000 ;
        RECT 503.600 302.200 504.400 306.000 ;
        RECT 505.200 302.200 506.000 306.200 ;
        RECT 506.800 306.000 510.800 306.200 ;
        RECT 506.800 302.200 507.600 306.000 ;
        RECT 510.000 302.200 510.800 306.000 ;
        RECT 511.600 302.200 512.400 306.200 ;
        RECT 513.800 305.600 515.600 306.200 ;
        RECT 518.600 305.600 520.400 306.200 ;
        RECT 513.800 302.200 514.600 305.600 ;
        RECT 518.600 304.400 519.400 305.600 ;
        RECT 518.000 303.600 519.400 304.400 ;
        RECT 518.600 302.200 519.400 303.600 ;
        RECT 522.800 302.200 523.600 306.200 ;
        RECT 524.400 306.000 528.400 306.200 ;
        RECT 524.400 302.200 525.200 306.000 ;
        RECT 527.600 302.200 528.400 306.000 ;
        RECT 529.200 302.200 530.000 306.800 ;
        RECT 532.400 302.200 533.200 309.600 ;
        RECT 534.000 306.800 534.800 308.400 ;
        RECT 535.600 306.200 536.400 319.800 ;
        RECT 537.200 311.600 538.000 313.200 ;
        RECT 538.800 312.400 539.600 319.800 ;
        RECT 542.000 312.800 542.800 319.800 ;
        RECT 538.800 311.800 541.400 312.400 ;
        RECT 542.000 311.800 543.000 312.800 ;
        RECT 538.800 309.600 539.800 310.400 ;
        RECT 539.000 308.800 539.800 309.600 ;
        RECT 540.800 309.800 541.400 311.800 ;
        RECT 540.800 309.000 541.800 309.800 ;
        RECT 540.800 307.400 541.400 309.000 ;
        RECT 542.400 308.400 543.000 311.800 ;
        RECT 542.000 307.600 543.000 308.400 ;
        RECT 538.800 306.800 541.400 307.400 ;
        RECT 535.600 305.600 537.400 306.200 ;
        RECT 536.600 304.400 537.400 305.600 ;
        RECT 536.600 303.600 538.000 304.400 ;
        RECT 536.600 302.200 537.400 303.600 ;
        RECT 538.800 302.200 539.600 306.800 ;
        RECT 542.400 306.200 543.000 307.600 ;
        RECT 542.000 305.600 543.000 306.200 ;
        RECT 542.000 302.200 542.800 305.600 ;
        RECT 546.800 302.200 547.600 319.800 ;
        RECT 551.600 316.400 552.400 319.800 ;
        RECT 551.400 315.800 552.400 316.400 ;
        RECT 551.400 315.200 552.000 315.800 ;
        RECT 554.800 315.200 555.600 319.800 ;
        RECT 558.000 317.000 558.800 319.800 ;
        RECT 559.600 317.000 560.400 319.800 ;
        RECT 550.000 314.600 552.000 315.200 ;
        RECT 550.000 309.000 550.800 314.600 ;
        RECT 552.600 314.400 556.800 315.200 ;
        RECT 561.200 315.000 562.000 319.800 ;
        RECT 564.400 315.000 565.200 319.800 ;
        RECT 552.600 314.000 553.200 314.400 ;
        RECT 551.600 313.200 553.200 314.000 ;
        RECT 556.200 313.800 562.000 314.400 ;
        RECT 554.200 313.200 555.600 313.800 ;
        RECT 554.200 313.000 560.400 313.200 ;
        RECT 555.000 312.600 560.400 313.000 ;
        RECT 559.600 312.400 560.400 312.600 ;
        RECT 561.400 313.000 562.000 313.800 ;
        RECT 562.600 313.600 565.200 314.400 ;
        RECT 567.600 313.600 568.400 319.800 ;
        RECT 569.200 317.000 570.000 319.800 ;
        RECT 570.800 317.000 571.600 319.800 ;
        RECT 572.400 317.000 573.200 319.800 ;
        RECT 570.800 314.400 575.000 315.200 ;
        RECT 575.600 314.400 576.400 319.800 ;
        RECT 578.800 315.200 579.600 319.800 ;
        RECT 578.800 314.600 581.400 315.200 ;
        RECT 575.600 313.600 578.200 314.400 ;
        RECT 569.200 313.000 570.000 313.200 ;
        RECT 561.400 312.400 570.000 313.000 ;
        RECT 572.400 313.000 573.200 313.200 ;
        RECT 580.800 313.000 581.400 314.600 ;
        RECT 572.400 312.400 581.400 313.000 ;
        RECT 580.800 310.600 581.400 312.400 ;
        RECT 582.000 312.000 582.800 319.800 ;
        RECT 586.000 313.600 586.800 314.400 ;
        RECT 586.000 312.400 586.600 313.600 ;
        RECT 587.400 312.400 588.200 319.800 ;
        RECT 582.000 311.200 583.000 312.000 ;
        RECT 585.200 311.800 586.600 312.400 ;
        RECT 587.200 311.800 588.200 312.400 ;
        RECT 585.200 311.600 586.000 311.800 ;
        RECT 551.400 310.000 574.800 310.600 ;
        RECT 580.800 310.000 581.600 310.600 ;
        RECT 551.400 309.800 552.200 310.000 ;
        RECT 556.400 309.600 557.200 310.000 ;
        RECT 574.000 309.400 574.800 310.000 ;
        RECT 550.000 308.200 558.800 309.000 ;
        RECT 559.400 308.600 561.400 309.400 ;
        RECT 565.200 308.600 568.400 309.400 ;
        RECT 550.000 302.200 550.800 308.200 ;
        RECT 552.400 306.800 555.400 307.600 ;
        RECT 554.600 306.200 555.400 306.800 ;
        RECT 560.600 306.200 561.400 308.600 ;
        RECT 562.800 306.800 563.600 308.400 ;
        RECT 568.000 307.800 568.800 308.000 ;
        RECT 564.400 307.200 568.800 307.800 ;
        RECT 564.400 307.000 565.200 307.200 ;
        RECT 570.800 306.400 571.600 309.200 ;
        RECT 576.600 308.600 580.400 309.400 ;
        RECT 576.600 307.400 577.400 308.600 ;
        RECT 581.000 308.000 581.600 310.000 ;
        RECT 564.400 306.200 565.200 306.400 ;
        RECT 554.600 305.400 557.200 306.200 ;
        RECT 560.600 305.600 565.200 306.200 ;
        RECT 566.000 305.600 567.600 306.400 ;
        RECT 570.600 305.600 571.600 306.400 ;
        RECT 575.600 306.800 577.400 307.400 ;
        RECT 580.400 307.400 581.600 308.000 ;
        RECT 575.600 306.200 576.400 306.800 ;
        RECT 556.400 302.200 557.200 305.400 ;
        RECT 574.000 305.400 576.400 306.200 ;
        RECT 558.000 302.200 558.800 305.000 ;
        RECT 559.600 302.200 560.400 305.000 ;
        RECT 561.200 302.200 562.000 305.000 ;
        RECT 564.400 302.200 565.200 305.000 ;
        RECT 567.600 302.200 568.400 305.000 ;
        RECT 569.200 302.200 570.000 305.000 ;
        RECT 570.800 302.200 571.600 305.000 ;
        RECT 572.400 302.200 573.200 305.000 ;
        RECT 574.000 302.200 574.800 305.400 ;
        RECT 580.400 302.200 581.200 307.400 ;
        RECT 582.200 306.800 583.000 311.200 ;
        RECT 587.200 308.400 587.800 311.800 ;
        RECT 588.400 310.300 589.200 310.400 ;
        RECT 591.600 310.300 592.400 319.800 ;
        RECT 595.600 313.600 596.400 314.400 ;
        RECT 595.600 312.400 596.200 313.600 ;
        RECT 597.000 312.400 597.800 319.800 ;
        RECT 593.200 312.300 594.000 312.400 ;
        RECT 594.800 312.300 596.200 312.400 ;
        RECT 593.200 311.800 596.200 312.300 ;
        RECT 596.800 311.800 597.800 312.400 ;
        RECT 593.200 311.700 595.600 311.800 ;
        RECT 593.200 311.600 594.000 311.700 ;
        RECT 594.800 311.600 595.600 311.700 ;
        RECT 588.400 309.700 592.400 310.300 ;
        RECT 588.400 308.800 589.200 309.700 ;
        RECT 585.200 307.600 587.800 308.400 ;
        RECT 590.000 308.200 590.800 308.400 ;
        RECT 589.200 307.600 590.800 308.200 ;
        RECT 582.000 306.000 583.000 306.800 ;
        RECT 585.400 306.200 586.000 307.600 ;
        RECT 589.200 307.200 590.000 307.600 ;
        RECT 587.000 306.200 590.600 306.600 ;
        RECT 582.000 302.200 582.800 306.000 ;
        RECT 585.200 302.200 586.000 306.200 ;
        RECT 586.800 306.000 590.800 306.200 ;
        RECT 586.800 302.200 587.600 306.000 ;
        RECT 590.000 302.200 590.800 306.000 ;
        RECT 591.600 302.200 592.400 309.700 ;
        RECT 596.800 308.400 597.400 311.800 ;
        RECT 598.000 310.300 598.800 310.400 ;
        RECT 601.200 310.300 602.000 319.800 ;
        RECT 604.400 312.400 605.200 319.800 ;
        RECT 604.400 311.800 606.600 312.400 ;
        RECT 606.000 311.200 606.600 311.800 ;
        RECT 606.000 310.400 607.200 311.200 ;
        RECT 598.000 309.700 602.000 310.300 ;
        RECT 598.000 308.800 598.800 309.700 ;
        RECT 594.800 307.600 597.400 308.400 ;
        RECT 599.600 308.200 600.400 308.400 ;
        RECT 598.800 307.600 600.400 308.200 ;
        RECT 593.200 304.800 594.000 306.400 ;
        RECT 595.000 306.200 595.600 307.600 ;
        RECT 598.800 307.200 599.600 307.600 ;
        RECT 596.600 306.200 600.200 306.600 ;
        RECT 594.800 302.200 595.600 306.200 ;
        RECT 596.400 306.000 600.400 306.200 ;
        RECT 596.400 302.200 597.200 306.000 ;
        RECT 599.600 302.200 600.400 306.000 ;
        RECT 601.200 302.200 602.000 309.700 ;
        RECT 604.400 308.800 605.200 310.400 ;
        RECT 606.000 307.400 606.600 310.400 ;
        RECT 604.400 306.800 606.600 307.400 ;
        RECT 602.800 304.800 603.600 306.400 ;
        RECT 604.400 302.200 605.200 306.800 ;
        RECT 2.800 295.200 3.600 299.800 ;
        RECT 6.000 295.200 6.800 299.800 ;
        RECT 9.200 295.200 10.000 299.800 ;
        RECT 12.400 295.200 13.200 299.800 ;
        RECT 2.800 294.400 4.600 295.200 ;
        RECT 6.000 294.400 8.200 295.200 ;
        RECT 9.200 294.400 11.400 295.200 ;
        RECT 12.400 294.400 14.800 295.200 ;
        RECT 1.200 293.800 2.000 294.400 ;
        RECT 3.800 293.800 4.600 294.400 ;
        RECT 7.400 293.800 8.200 294.400 ;
        RECT 10.600 293.800 11.400 294.400 ;
        RECT 1.200 293.000 3.000 293.800 ;
        RECT 3.800 293.000 6.400 293.800 ;
        RECT 7.400 293.000 9.800 293.800 ;
        RECT 10.600 293.000 13.200 293.800 ;
        RECT 3.800 291.600 4.600 293.000 ;
        RECT 7.400 291.600 8.200 293.000 ;
        RECT 10.600 291.600 11.400 293.000 ;
        RECT 14.000 291.600 14.800 294.400 ;
        RECT 2.800 290.800 4.600 291.600 ;
        RECT 6.000 290.800 8.200 291.600 ;
        RECT 9.200 290.800 11.400 291.600 ;
        RECT 12.400 290.800 14.800 291.600 ;
        RECT 15.600 293.800 16.400 299.800 ;
        RECT 22.000 296.600 22.800 299.800 ;
        RECT 23.600 297.000 24.400 299.800 ;
        RECT 25.200 297.000 26.000 299.800 ;
        RECT 26.800 297.000 27.600 299.800 ;
        RECT 30.000 297.000 30.800 299.800 ;
        RECT 33.200 297.000 34.000 299.800 ;
        RECT 34.800 297.000 35.600 299.800 ;
        RECT 36.400 297.000 37.200 299.800 ;
        RECT 38.000 297.000 38.800 299.800 ;
        RECT 20.200 295.800 22.800 296.600 ;
        RECT 39.600 296.600 40.400 299.800 ;
        RECT 26.200 295.800 30.800 296.400 ;
        RECT 20.200 295.200 21.000 295.800 ;
        RECT 18.000 294.400 21.000 295.200 ;
        RECT 15.600 293.000 24.400 293.800 ;
        RECT 26.200 293.400 27.000 295.800 ;
        RECT 30.000 295.600 30.800 295.800 ;
        RECT 31.600 295.600 33.200 296.400 ;
        RECT 36.200 295.600 37.200 296.400 ;
        RECT 39.600 295.800 42.000 296.600 ;
        RECT 28.400 293.600 29.200 295.200 ;
        RECT 30.000 294.800 30.800 295.000 ;
        RECT 30.000 294.200 34.400 294.800 ;
        RECT 33.600 294.000 34.400 294.200 ;
        RECT 2.800 282.200 3.600 290.800 ;
        RECT 6.000 282.200 6.800 290.800 ;
        RECT 9.200 282.200 10.000 290.800 ;
        RECT 12.400 282.200 13.200 290.800 ;
        RECT 15.600 287.400 16.400 293.000 ;
        RECT 25.000 292.600 27.000 293.400 ;
        RECT 30.800 292.600 34.000 293.400 ;
        RECT 36.400 292.800 37.200 295.600 ;
        RECT 41.200 295.200 42.000 295.800 ;
        RECT 41.200 294.600 43.000 295.200 ;
        RECT 42.200 293.400 43.000 294.600 ;
        RECT 46.000 294.600 46.800 299.800 ;
        RECT 47.600 296.300 48.400 299.800 ;
        RECT 52.400 297.800 53.200 299.800 ;
        RECT 50.800 296.300 51.600 297.200 ;
        RECT 52.600 296.300 53.200 297.800 ;
        RECT 55.800 296.400 56.600 297.200 ;
        RECT 55.600 296.300 56.400 296.400 ;
        RECT 47.600 295.700 51.600 296.300 ;
        RECT 52.500 295.700 56.400 296.300 ;
        RECT 47.600 295.200 48.600 295.700 ;
        RECT 50.800 295.600 51.600 295.700 ;
        RECT 46.000 294.000 47.200 294.600 ;
        RECT 42.200 292.600 46.000 293.400 ;
        RECT 17.000 292.000 17.800 292.200 ;
        RECT 18.800 292.000 19.600 292.400 ;
        RECT 22.000 292.000 22.800 292.400 ;
        RECT 28.400 292.000 29.200 292.400 ;
        RECT 39.600 292.000 40.400 292.600 ;
        RECT 46.600 292.000 47.200 294.000 ;
        RECT 17.000 291.400 40.400 292.000 ;
        RECT 46.400 291.400 47.200 292.000 ;
        RECT 46.400 289.600 47.000 291.400 ;
        RECT 47.800 290.800 48.600 295.200 ;
        RECT 52.600 294.400 53.200 295.700 ;
        RECT 55.600 295.600 56.400 295.700 ;
        RECT 57.200 295.600 58.000 299.800 ;
        RECT 52.400 293.600 53.200 294.400 ;
        RECT 25.200 289.400 26.000 289.600 ;
        RECT 20.600 289.000 26.000 289.400 ;
        RECT 19.800 288.800 26.000 289.000 ;
        RECT 27.000 289.000 35.600 289.600 ;
        RECT 17.200 288.000 18.800 288.800 ;
        RECT 19.800 288.200 21.200 288.800 ;
        RECT 27.000 288.200 27.600 289.000 ;
        RECT 34.800 288.800 35.600 289.000 ;
        RECT 38.000 289.000 47.000 289.600 ;
        RECT 38.000 288.800 38.800 289.000 ;
        RECT 18.200 287.600 18.800 288.000 ;
        RECT 21.800 287.600 27.600 288.200 ;
        RECT 28.200 287.600 30.800 288.400 ;
        RECT 15.600 286.800 17.600 287.400 ;
        RECT 18.200 286.800 22.400 287.600 ;
        RECT 17.000 286.200 17.600 286.800 ;
        RECT 17.000 285.600 18.000 286.200 ;
        RECT 17.200 282.200 18.000 285.600 ;
        RECT 20.400 282.200 21.200 286.800 ;
        RECT 23.600 282.200 24.400 285.000 ;
        RECT 25.200 282.200 26.000 285.000 ;
        RECT 26.800 282.200 27.600 287.000 ;
        RECT 30.000 282.200 30.800 287.000 ;
        RECT 33.200 282.200 34.000 288.400 ;
        RECT 41.200 287.600 43.800 288.400 ;
        RECT 36.400 286.800 40.600 287.600 ;
        RECT 34.800 282.200 35.600 285.000 ;
        RECT 36.400 282.200 37.200 285.000 ;
        RECT 38.000 282.200 38.800 285.000 ;
        RECT 41.200 282.200 42.000 287.600 ;
        RECT 46.400 287.400 47.000 289.000 ;
        RECT 44.400 286.800 47.000 287.400 ;
        RECT 47.600 290.000 48.600 290.800 ;
        RECT 52.600 290.200 53.200 293.600 ;
        RECT 54.000 290.800 54.800 292.400 ;
        RECT 55.600 292.200 56.400 292.400 ;
        RECT 57.400 292.200 58.000 295.600 ;
        RECT 58.800 292.800 59.600 294.400 ;
        RECT 62.000 293.800 62.800 299.800 ;
        RECT 68.400 296.600 69.200 299.800 ;
        RECT 70.000 297.000 70.800 299.800 ;
        RECT 71.600 297.000 72.400 299.800 ;
        RECT 73.200 297.000 74.000 299.800 ;
        RECT 76.400 297.000 77.200 299.800 ;
        RECT 79.600 297.000 80.400 299.800 ;
        RECT 81.200 297.000 82.000 299.800 ;
        RECT 82.800 297.000 83.600 299.800 ;
        RECT 84.400 297.000 85.200 299.800 ;
        RECT 66.600 295.800 69.200 296.600 ;
        RECT 86.000 296.600 86.800 299.800 ;
        RECT 72.600 295.800 77.200 296.400 ;
        RECT 66.600 295.200 67.400 295.800 ;
        RECT 64.400 294.400 67.400 295.200 ;
        RECT 62.000 293.000 70.800 293.800 ;
        RECT 72.600 293.400 73.400 295.800 ;
        RECT 76.400 295.600 77.200 295.800 ;
        RECT 78.000 295.600 79.600 296.400 ;
        RECT 82.600 295.600 83.600 296.400 ;
        RECT 86.000 295.800 88.400 296.600 ;
        RECT 74.800 293.600 75.600 295.200 ;
        RECT 76.400 294.800 77.200 295.000 ;
        RECT 76.400 294.200 80.800 294.800 ;
        RECT 80.000 294.000 80.800 294.200 ;
        RECT 60.400 292.200 61.200 292.400 ;
        RECT 55.600 291.600 58.000 292.200 ;
        RECT 59.600 291.600 61.200 292.200 ;
        RECT 55.800 290.200 56.400 291.600 ;
        RECT 59.600 291.200 60.400 291.600 ;
        RECT 44.400 282.200 45.200 286.800 ;
        RECT 47.600 282.200 48.400 290.000 ;
        RECT 52.400 289.400 54.200 290.200 ;
        RECT 53.400 282.200 54.200 289.400 ;
        RECT 55.600 282.200 56.400 290.200 ;
        RECT 57.200 289.600 61.200 290.200 ;
        RECT 57.200 282.200 58.000 289.600 ;
        RECT 60.400 282.200 61.200 289.600 ;
        RECT 62.000 287.400 62.800 293.000 ;
        RECT 71.400 292.600 73.400 293.400 ;
        RECT 77.200 292.600 80.400 293.400 ;
        RECT 82.800 292.800 83.600 295.600 ;
        RECT 87.600 295.200 88.400 295.800 ;
        RECT 87.600 294.600 89.400 295.200 ;
        RECT 88.600 293.400 89.400 294.600 ;
        RECT 92.400 294.600 93.200 299.800 ;
        RECT 94.000 296.300 94.800 299.800 ;
        RECT 98.800 297.800 99.600 299.800 ;
        RECT 97.200 296.300 98.000 297.200 ;
        RECT 99.000 296.300 99.600 297.800 ;
        RECT 102.200 296.400 103.000 297.200 ;
        RECT 102.000 296.300 102.800 296.400 ;
        RECT 94.000 295.700 98.000 296.300 ;
        RECT 98.900 295.700 102.800 296.300 ;
        RECT 103.600 295.800 104.400 299.800 ;
        RECT 94.000 295.200 95.000 295.700 ;
        RECT 97.200 295.600 98.000 295.700 ;
        RECT 92.400 294.000 93.600 294.600 ;
        RECT 88.600 292.600 92.400 293.400 ;
        RECT 63.400 292.000 64.200 292.200 ;
        RECT 68.400 292.000 69.200 292.400 ;
        RECT 86.000 292.000 86.800 292.600 ;
        RECT 93.000 292.000 93.600 294.000 ;
        RECT 63.400 291.400 86.800 292.000 ;
        RECT 92.800 291.400 93.600 292.000 ;
        RECT 92.800 289.600 93.400 291.400 ;
        RECT 94.200 290.800 95.000 295.200 ;
        RECT 99.000 294.400 99.600 295.700 ;
        RECT 102.000 295.600 102.800 295.700 ;
        RECT 98.800 293.600 99.600 294.400 ;
        RECT 71.600 289.400 72.400 289.600 ;
        RECT 67.000 289.000 72.400 289.400 ;
        RECT 66.200 288.800 72.400 289.000 ;
        RECT 73.400 289.000 82.000 289.600 ;
        RECT 63.600 288.000 65.200 288.800 ;
        RECT 66.200 288.200 67.600 288.800 ;
        RECT 73.400 288.200 74.000 289.000 ;
        RECT 81.200 288.800 82.000 289.000 ;
        RECT 84.400 289.000 93.400 289.600 ;
        RECT 84.400 288.800 85.200 289.000 ;
        RECT 64.600 287.600 65.200 288.000 ;
        RECT 68.200 287.600 74.000 288.200 ;
        RECT 74.600 287.600 77.200 288.400 ;
        RECT 62.000 286.800 64.000 287.400 ;
        RECT 64.600 286.800 68.800 287.600 ;
        RECT 63.400 286.200 64.000 286.800 ;
        RECT 63.400 285.600 64.400 286.200 ;
        RECT 63.600 282.200 64.400 285.600 ;
        RECT 66.800 282.200 67.600 286.800 ;
        RECT 70.000 282.200 70.800 285.000 ;
        RECT 71.600 282.200 72.400 285.000 ;
        RECT 73.200 282.200 74.000 287.000 ;
        RECT 76.400 282.200 77.200 287.000 ;
        RECT 79.600 282.200 80.400 288.400 ;
        RECT 87.600 287.600 90.200 288.400 ;
        RECT 82.800 286.800 87.000 287.600 ;
        RECT 81.200 282.200 82.000 285.000 ;
        RECT 82.800 282.200 83.600 285.000 ;
        RECT 84.400 282.200 85.200 285.000 ;
        RECT 87.600 282.200 88.400 287.600 ;
        RECT 92.800 287.400 93.400 289.000 ;
        RECT 90.800 286.800 93.400 287.400 ;
        RECT 94.000 290.000 95.000 290.800 ;
        RECT 99.000 290.200 99.600 293.600 ;
        RECT 100.400 290.800 101.200 292.400 ;
        RECT 102.000 292.200 102.800 292.400 ;
        RECT 103.800 292.200 104.400 295.800 ;
        RECT 108.400 295.600 109.200 297.200 ;
        RECT 105.200 292.800 106.000 294.400 ;
        RECT 106.800 292.200 107.600 292.400 ;
        RECT 102.000 291.600 104.400 292.200 ;
        RECT 106.000 291.600 107.600 292.200 ;
        RECT 102.200 290.200 102.800 291.600 ;
        RECT 106.000 291.200 106.800 291.600 ;
        RECT 90.800 282.200 91.600 286.800 ;
        RECT 94.000 282.200 94.800 290.000 ;
        RECT 98.800 289.400 100.600 290.200 ;
        RECT 99.800 282.200 100.600 289.400 ;
        RECT 102.000 282.200 102.800 290.200 ;
        RECT 103.600 289.600 107.600 290.200 ;
        RECT 103.600 282.200 104.400 289.600 ;
        RECT 106.800 282.200 107.600 289.600 ;
        RECT 110.000 282.200 110.800 299.800 ;
        RECT 111.600 297.000 112.400 299.000 ;
        RECT 111.600 294.800 112.200 297.000 ;
        RECT 115.800 296.000 116.600 299.000 ;
        RECT 122.800 296.000 123.600 299.800 ;
        RECT 115.800 295.400 117.400 296.000 ;
        RECT 116.600 295.000 117.400 295.400 ;
        RECT 111.600 294.200 115.800 294.800 ;
        RECT 114.800 293.800 115.800 294.200 ;
        RECT 116.800 294.400 117.400 295.000 ;
        RECT 122.600 295.200 123.600 296.000 ;
        RECT 111.600 291.600 112.400 293.200 ;
        RECT 113.200 291.600 114.000 293.200 ;
        RECT 114.800 293.000 116.200 293.800 ;
        RECT 116.800 293.600 118.800 294.400 ;
        RECT 114.800 291.000 115.400 293.000 ;
        RECT 111.600 290.400 115.400 291.000 ;
        RECT 111.600 287.000 112.200 290.400 ;
        RECT 116.800 289.800 117.400 293.600 ;
        RECT 118.000 290.800 118.800 292.400 ;
        RECT 122.600 290.800 123.400 295.200 ;
        RECT 124.400 294.600 125.200 299.800 ;
        RECT 130.800 296.600 131.600 299.800 ;
        RECT 132.400 297.000 133.200 299.800 ;
        RECT 134.000 297.000 134.800 299.800 ;
        RECT 135.600 297.000 136.400 299.800 ;
        RECT 137.200 297.000 138.000 299.800 ;
        RECT 140.400 297.000 141.200 299.800 ;
        RECT 143.600 297.000 144.400 299.800 ;
        RECT 145.200 297.000 146.000 299.800 ;
        RECT 146.800 297.000 147.600 299.800 ;
        RECT 129.200 295.800 131.600 296.600 ;
        RECT 148.400 296.600 149.200 299.800 ;
        RECT 129.200 295.200 130.000 295.800 ;
        RECT 124.000 294.000 125.200 294.600 ;
        RECT 128.200 294.600 130.000 295.200 ;
        RECT 134.000 295.600 135.000 296.400 ;
        RECT 138.000 295.600 139.600 296.400 ;
        RECT 140.400 295.800 145.000 296.400 ;
        RECT 148.400 295.800 151.000 296.600 ;
        RECT 140.400 295.600 141.200 295.800 ;
        RECT 124.000 292.000 124.600 294.000 ;
        RECT 128.200 293.400 129.000 294.600 ;
        RECT 125.200 292.600 129.000 293.400 ;
        RECT 134.000 292.800 134.800 295.600 ;
        RECT 140.400 294.800 141.200 295.000 ;
        RECT 136.800 294.200 141.200 294.800 ;
        RECT 136.800 294.000 137.600 294.200 ;
        RECT 142.000 293.600 142.800 295.200 ;
        RECT 144.200 293.400 145.000 295.800 ;
        RECT 150.200 295.200 151.000 295.800 ;
        RECT 150.200 294.400 153.200 295.200 ;
        RECT 154.800 293.800 155.600 299.800 ;
        RECT 161.200 295.600 162.000 297.200 ;
        RECT 137.200 292.600 140.400 293.400 ;
        RECT 144.200 292.600 146.200 293.400 ;
        RECT 146.800 293.000 155.600 293.800 ;
        RECT 130.800 292.000 131.600 292.600 ;
        RECT 148.400 292.000 149.200 292.400 ;
        RECT 151.600 292.000 152.400 292.400 ;
        RECT 153.400 292.000 154.200 292.200 ;
        RECT 124.000 291.400 124.800 292.000 ;
        RECT 130.800 291.400 154.200 292.000 ;
        RECT 122.600 290.000 123.600 290.800 ;
        RECT 115.800 289.200 117.400 289.800 ;
        RECT 111.600 283.000 112.400 287.000 ;
        RECT 115.800 284.400 116.600 289.200 ;
        RECT 114.800 283.600 116.600 284.400 ;
        RECT 115.800 282.200 116.600 283.600 ;
        RECT 122.800 282.200 123.600 290.000 ;
        RECT 124.200 289.600 124.800 291.400 ;
        RECT 124.200 289.000 133.200 289.600 ;
        RECT 124.200 287.400 124.800 289.000 ;
        RECT 132.400 288.800 133.200 289.000 ;
        RECT 135.600 289.000 144.200 289.600 ;
        RECT 135.600 288.800 136.400 289.000 ;
        RECT 127.400 287.600 130.000 288.400 ;
        RECT 124.200 286.800 126.800 287.400 ;
        RECT 126.000 282.200 126.800 286.800 ;
        RECT 129.200 282.200 130.000 287.600 ;
        RECT 130.600 286.800 134.800 287.600 ;
        RECT 132.400 282.200 133.200 285.000 ;
        RECT 134.000 282.200 134.800 285.000 ;
        RECT 135.600 282.200 136.400 285.000 ;
        RECT 137.200 282.200 138.000 288.400 ;
        RECT 140.400 287.600 143.000 288.400 ;
        RECT 143.600 288.200 144.200 289.000 ;
        RECT 145.200 289.400 146.000 289.600 ;
        RECT 145.200 289.000 150.600 289.400 ;
        RECT 145.200 288.800 151.400 289.000 ;
        RECT 150.000 288.200 151.400 288.800 ;
        RECT 143.600 287.600 149.400 288.200 ;
        RECT 152.400 288.000 154.000 288.800 ;
        RECT 152.400 287.600 153.000 288.000 ;
        RECT 140.400 282.200 141.200 287.000 ;
        RECT 143.600 282.200 144.400 287.000 ;
        RECT 148.800 286.800 153.000 287.600 ;
        RECT 154.800 287.400 155.600 293.000 ;
        RECT 153.600 286.800 155.600 287.400 ;
        RECT 162.800 294.300 163.600 299.800 ;
        RECT 164.400 296.000 165.200 299.800 ;
        RECT 167.600 296.000 168.400 299.800 ;
        RECT 164.400 295.800 168.400 296.000 ;
        RECT 169.200 295.800 170.000 299.800 ;
        RECT 164.600 295.400 168.200 295.800 ;
        RECT 165.200 294.400 166.000 294.800 ;
        RECT 169.200 294.400 169.800 295.800 ;
        RECT 164.400 294.300 166.000 294.400 ;
        RECT 162.800 293.800 166.000 294.300 ;
        RECT 162.800 293.700 165.200 293.800 ;
        RECT 145.200 282.200 146.000 285.000 ;
        RECT 146.800 282.200 147.600 285.000 ;
        RECT 150.000 282.200 150.800 286.800 ;
        RECT 153.600 286.200 154.200 286.800 ;
        RECT 153.200 285.600 154.200 286.200 ;
        RECT 153.200 282.200 154.000 285.600 ;
        RECT 162.800 282.200 163.600 293.700 ;
        RECT 164.400 293.600 165.200 293.700 ;
        RECT 167.400 293.600 170.000 294.400 ;
        RECT 170.800 293.800 171.600 299.800 ;
        RECT 177.200 296.600 178.000 299.800 ;
        RECT 178.800 297.000 179.600 299.800 ;
        RECT 180.400 297.000 181.200 299.800 ;
        RECT 182.000 297.000 182.800 299.800 ;
        RECT 185.200 297.000 186.000 299.800 ;
        RECT 188.400 297.000 189.200 299.800 ;
        RECT 190.000 297.000 190.800 299.800 ;
        RECT 191.600 297.000 192.400 299.800 ;
        RECT 193.200 297.000 194.000 299.800 ;
        RECT 175.400 295.800 178.000 296.600 ;
        RECT 194.800 296.600 195.600 299.800 ;
        RECT 181.400 295.800 186.000 296.400 ;
        RECT 175.400 295.200 176.200 295.800 ;
        RECT 173.200 294.400 176.200 295.200 ;
        RECT 166.000 291.600 166.800 293.200 ;
        RECT 167.400 290.200 168.000 293.600 ;
        RECT 170.800 293.000 179.600 293.800 ;
        RECT 181.400 293.400 182.200 295.800 ;
        RECT 185.200 295.600 186.000 295.800 ;
        RECT 186.800 295.600 188.400 296.400 ;
        RECT 191.400 295.600 192.400 296.400 ;
        RECT 194.800 295.800 197.200 296.600 ;
        RECT 183.600 293.600 184.400 295.200 ;
        RECT 185.200 294.800 186.000 295.000 ;
        RECT 185.200 294.200 189.600 294.800 ;
        RECT 188.800 294.000 189.600 294.200 ;
        RECT 169.200 290.200 170.000 290.400 ;
        RECT 167.000 289.600 168.000 290.200 ;
        RECT 168.600 289.600 170.000 290.200 ;
        RECT 167.000 282.200 167.800 289.600 ;
        RECT 168.600 288.400 169.200 289.600 ;
        RECT 168.400 287.600 169.200 288.400 ;
        RECT 170.800 287.400 171.600 293.000 ;
        RECT 180.200 292.600 182.200 293.400 ;
        RECT 186.000 292.600 189.200 293.400 ;
        RECT 191.600 292.800 192.400 295.600 ;
        RECT 196.400 295.200 197.200 295.800 ;
        RECT 196.400 294.600 198.200 295.200 ;
        RECT 197.400 293.400 198.200 294.600 ;
        RECT 201.200 294.600 202.000 299.800 ;
        RECT 202.800 296.000 203.600 299.800 ;
        RECT 202.800 295.200 203.800 296.000 ;
        RECT 201.200 294.000 202.400 294.600 ;
        RECT 197.400 292.600 201.200 293.400 ;
        RECT 172.200 292.000 173.000 292.200 ;
        RECT 175.600 292.000 176.400 292.400 ;
        RECT 177.200 292.000 178.000 292.400 ;
        RECT 194.800 292.000 195.600 292.600 ;
        RECT 201.800 292.000 202.400 294.000 ;
        RECT 172.200 291.400 195.600 292.000 ;
        RECT 201.600 291.400 202.400 292.000 ;
        RECT 203.000 294.300 203.800 295.200 ;
        RECT 206.000 294.300 206.800 295.200 ;
        RECT 203.000 293.700 206.800 294.300 ;
        RECT 201.600 289.600 202.200 291.400 ;
        RECT 203.000 290.800 203.800 293.700 ;
        RECT 206.000 293.600 206.800 293.700 ;
        RECT 180.400 289.400 181.200 289.600 ;
        RECT 175.800 289.000 181.200 289.400 ;
        RECT 175.000 288.800 181.200 289.000 ;
        RECT 182.200 289.000 190.800 289.600 ;
        RECT 172.400 288.000 174.000 288.800 ;
        RECT 175.000 288.200 176.400 288.800 ;
        RECT 182.200 288.200 182.800 289.000 ;
        RECT 190.000 288.800 190.800 289.000 ;
        RECT 193.200 289.000 202.200 289.600 ;
        RECT 193.200 288.800 194.000 289.000 ;
        RECT 173.400 287.600 174.000 288.000 ;
        RECT 177.000 287.600 182.800 288.200 ;
        RECT 183.400 287.600 186.000 288.400 ;
        RECT 170.800 286.800 172.800 287.400 ;
        RECT 173.400 286.800 177.600 287.600 ;
        RECT 172.200 286.200 172.800 286.800 ;
        RECT 172.200 285.600 173.200 286.200 ;
        RECT 172.400 282.200 173.200 285.600 ;
        RECT 175.600 282.200 176.400 286.800 ;
        RECT 178.800 282.200 179.600 285.000 ;
        RECT 180.400 282.200 181.200 285.000 ;
        RECT 182.000 282.200 182.800 287.000 ;
        RECT 185.200 282.200 186.000 287.000 ;
        RECT 188.400 282.200 189.200 288.400 ;
        RECT 196.400 287.600 199.000 288.400 ;
        RECT 191.600 286.800 195.800 287.600 ;
        RECT 190.000 282.200 190.800 285.000 ;
        RECT 191.600 282.200 192.400 285.000 ;
        RECT 193.200 282.200 194.000 285.000 ;
        RECT 196.400 282.200 197.200 287.600 ;
        RECT 201.600 287.400 202.200 289.000 ;
        RECT 199.600 286.800 202.200 287.400 ;
        RECT 202.800 290.000 203.800 290.800 ;
        RECT 199.600 282.200 200.400 286.800 ;
        RECT 202.800 282.200 203.600 290.000 ;
        RECT 207.600 282.200 208.400 299.800 ;
        RECT 211.800 296.400 212.600 299.800 ;
        RECT 216.600 296.400 217.400 299.800 ;
        RECT 210.800 295.800 212.600 296.400 ;
        RECT 215.600 295.800 217.400 296.400 ;
        RECT 209.200 293.600 210.000 295.200 ;
        RECT 210.800 294.300 211.600 295.800 ;
        RECT 214.000 294.300 214.800 295.200 ;
        RECT 210.800 293.700 214.800 294.300 ;
        RECT 210.800 282.200 211.600 293.700 ;
        RECT 214.000 293.600 214.800 293.700 ;
        RECT 212.400 292.300 213.200 292.400 ;
        RECT 215.600 292.300 216.400 295.800 ;
        RECT 212.400 291.700 216.400 292.300 ;
        RECT 212.400 291.600 213.200 291.700 ;
        RECT 212.400 290.300 213.200 290.400 ;
        RECT 214.000 290.300 214.800 290.400 ;
        RECT 212.400 289.700 214.800 290.300 ;
        RECT 212.400 288.800 213.200 289.700 ;
        RECT 214.000 289.600 214.800 289.700 ;
        RECT 215.600 282.200 216.400 291.700 ;
        RECT 218.800 293.800 219.600 299.800 ;
        RECT 225.200 296.600 226.000 299.800 ;
        RECT 226.800 297.000 227.600 299.800 ;
        RECT 228.400 297.000 229.200 299.800 ;
        RECT 230.000 297.000 230.800 299.800 ;
        RECT 233.200 297.000 234.000 299.800 ;
        RECT 236.400 297.000 237.200 299.800 ;
        RECT 238.000 297.000 238.800 299.800 ;
        RECT 239.600 297.000 240.400 299.800 ;
        RECT 241.200 297.000 242.000 299.800 ;
        RECT 223.400 295.800 226.000 296.600 ;
        RECT 242.800 296.600 243.600 299.800 ;
        RECT 229.400 295.800 234.000 296.400 ;
        RECT 223.400 295.200 224.200 295.800 ;
        RECT 221.200 294.400 224.200 295.200 ;
        RECT 218.800 293.000 227.600 293.800 ;
        RECT 229.400 293.400 230.200 295.800 ;
        RECT 233.200 295.600 234.000 295.800 ;
        RECT 234.800 295.600 236.400 296.400 ;
        RECT 239.400 295.600 240.400 296.400 ;
        RECT 242.800 295.800 245.200 296.600 ;
        RECT 231.600 293.600 232.400 295.200 ;
        RECT 233.200 294.800 234.000 295.000 ;
        RECT 233.200 294.200 237.600 294.800 ;
        RECT 236.800 294.000 237.600 294.200 ;
        RECT 217.200 288.800 218.000 290.400 ;
        RECT 218.800 287.400 219.600 293.000 ;
        RECT 228.200 292.600 230.200 293.400 ;
        RECT 234.000 292.600 237.200 293.400 ;
        RECT 239.600 292.800 240.400 295.600 ;
        RECT 244.400 295.200 245.200 295.800 ;
        RECT 244.400 294.600 246.200 295.200 ;
        RECT 245.400 293.400 246.200 294.600 ;
        RECT 249.200 294.600 250.000 299.800 ;
        RECT 250.800 296.300 251.600 299.800 ;
        RECT 254.000 296.300 254.800 297.200 ;
        RECT 250.800 295.700 254.800 296.300 ;
        RECT 250.800 295.200 251.800 295.700 ;
        RECT 254.000 295.600 254.800 295.700 ;
        RECT 249.200 294.000 250.400 294.600 ;
        RECT 245.400 292.600 249.200 293.400 ;
        RECT 220.200 292.000 221.000 292.200 ;
        RECT 222.000 292.000 222.800 292.400 ;
        RECT 225.200 292.000 226.000 292.400 ;
        RECT 242.800 292.000 243.600 292.600 ;
        RECT 249.800 292.000 250.400 294.000 ;
        RECT 220.200 291.400 243.600 292.000 ;
        RECT 249.600 291.400 250.400 292.000 ;
        RECT 249.600 289.600 250.200 291.400 ;
        RECT 251.000 290.800 251.800 295.200 ;
        RECT 228.400 289.400 229.200 289.600 ;
        RECT 223.800 289.000 229.200 289.400 ;
        RECT 223.000 288.800 229.200 289.000 ;
        RECT 230.200 289.000 238.800 289.600 ;
        RECT 220.400 288.000 222.000 288.800 ;
        RECT 223.000 288.200 224.400 288.800 ;
        RECT 230.200 288.200 230.800 289.000 ;
        RECT 238.000 288.800 238.800 289.000 ;
        RECT 241.200 289.000 250.200 289.600 ;
        RECT 241.200 288.800 242.000 289.000 ;
        RECT 221.400 287.600 222.000 288.000 ;
        RECT 225.000 287.600 230.800 288.200 ;
        RECT 231.400 287.600 234.000 288.400 ;
        RECT 218.800 286.800 220.800 287.400 ;
        RECT 221.400 286.800 225.600 287.600 ;
        RECT 220.200 286.200 220.800 286.800 ;
        RECT 220.200 285.600 221.200 286.200 ;
        RECT 220.400 282.200 221.200 285.600 ;
        RECT 223.600 282.200 224.400 286.800 ;
        RECT 226.800 282.200 227.600 285.000 ;
        RECT 228.400 282.200 229.200 285.000 ;
        RECT 230.000 282.200 230.800 287.000 ;
        RECT 233.200 282.200 234.000 287.000 ;
        RECT 236.400 282.200 237.200 288.400 ;
        RECT 244.400 287.600 247.000 288.400 ;
        RECT 239.600 286.800 243.800 287.600 ;
        RECT 238.000 282.200 238.800 285.000 ;
        RECT 239.600 282.200 240.400 285.000 ;
        RECT 241.200 282.200 242.000 285.000 ;
        RECT 244.400 282.200 245.200 287.600 ;
        RECT 249.600 287.400 250.200 289.000 ;
        RECT 247.600 286.800 250.200 287.400 ;
        RECT 250.800 290.000 251.800 290.800 ;
        RECT 255.600 292.300 256.400 299.800 ;
        RECT 261.000 296.000 261.800 299.000 ;
        RECT 265.200 297.000 266.000 299.000 ;
        RECT 260.200 295.400 261.800 296.000 ;
        RECT 260.200 295.000 261.000 295.400 ;
        RECT 260.200 294.400 260.800 295.000 ;
        RECT 265.400 294.800 266.000 297.000 ;
        RECT 257.200 294.300 258.000 294.400 ;
        RECT 258.800 294.300 260.800 294.400 ;
        RECT 257.200 293.700 260.800 294.300 ;
        RECT 261.800 294.200 266.000 294.800 ;
        RECT 261.800 293.800 262.800 294.200 ;
        RECT 257.200 293.600 258.000 293.700 ;
        RECT 258.800 293.600 260.800 293.700 ;
        RECT 258.800 292.300 259.600 292.400 ;
        RECT 255.600 291.700 259.600 292.300 ;
        RECT 247.600 282.200 248.400 286.800 ;
        RECT 250.800 282.200 251.600 290.000 ;
        RECT 255.600 282.200 256.400 291.700 ;
        RECT 258.800 290.800 259.600 291.700 ;
        RECT 260.200 289.800 260.800 293.600 ;
        RECT 261.400 293.000 262.800 293.800 ;
        RECT 266.800 293.800 267.600 299.800 ;
        RECT 273.200 296.600 274.000 299.800 ;
        RECT 274.800 297.000 275.600 299.800 ;
        RECT 276.400 297.000 277.200 299.800 ;
        RECT 278.000 297.000 278.800 299.800 ;
        RECT 281.200 297.000 282.000 299.800 ;
        RECT 284.400 297.000 285.200 299.800 ;
        RECT 286.000 297.000 286.800 299.800 ;
        RECT 287.600 297.000 288.400 299.800 ;
        RECT 289.200 297.000 290.000 299.800 ;
        RECT 271.400 295.800 274.000 296.600 ;
        RECT 290.800 296.600 291.600 299.800 ;
        RECT 277.400 295.800 282.000 296.400 ;
        RECT 271.400 295.200 272.200 295.800 ;
        RECT 269.200 294.400 272.200 295.200 ;
        RECT 262.200 291.000 262.800 293.000 ;
        RECT 263.600 291.600 264.400 293.200 ;
        RECT 265.200 291.600 266.000 293.200 ;
        RECT 266.800 293.000 275.600 293.800 ;
        RECT 277.400 293.400 278.200 295.800 ;
        RECT 281.200 295.600 282.000 295.800 ;
        RECT 282.800 295.600 284.400 296.400 ;
        RECT 287.400 295.600 288.400 296.400 ;
        RECT 290.800 295.800 293.200 296.600 ;
        RECT 279.600 293.600 280.400 295.200 ;
        RECT 281.200 294.800 282.000 295.000 ;
        RECT 281.200 294.200 285.600 294.800 ;
        RECT 284.800 294.000 285.600 294.200 ;
        RECT 262.200 290.400 266.000 291.000 ;
        RECT 260.200 289.200 261.800 289.800 ;
        RECT 261.000 282.200 261.800 289.200 ;
        RECT 265.400 287.000 266.000 290.400 ;
        RECT 265.200 283.000 266.000 287.000 ;
        RECT 266.800 287.400 267.600 293.000 ;
        RECT 276.200 292.600 278.200 293.400 ;
        RECT 282.000 292.600 285.200 293.400 ;
        RECT 287.600 292.800 288.400 295.600 ;
        RECT 292.400 295.200 293.200 295.800 ;
        RECT 292.400 294.600 294.200 295.200 ;
        RECT 293.400 293.400 294.200 294.600 ;
        RECT 297.200 294.600 298.000 299.800 ;
        RECT 298.800 296.000 299.600 299.800 ;
        RECT 304.600 296.400 305.400 299.800 ;
        RECT 314.200 296.400 315.000 299.800 ;
        RECT 319.000 296.400 319.800 299.800 ;
        RECT 298.800 295.200 299.800 296.000 ;
        RECT 303.600 295.800 305.400 296.400 ;
        RECT 313.200 295.800 315.000 296.400 ;
        RECT 318.000 295.800 319.800 296.400 ;
        RECT 321.200 296.000 322.000 299.800 ;
        RECT 324.400 296.000 325.200 299.800 ;
        RECT 321.200 295.800 325.200 296.000 ;
        RECT 326.000 295.800 326.800 299.800 ;
        RECT 327.600 296.000 328.400 299.800 ;
        RECT 330.800 296.000 331.600 299.800 ;
        RECT 327.600 295.800 331.600 296.000 ;
        RECT 332.400 295.800 333.200 299.800 ;
        RECT 336.600 298.400 337.400 299.800 ;
        RECT 335.600 297.600 337.400 298.400 ;
        RECT 340.400 297.800 341.200 299.800 ;
        RECT 336.600 296.400 337.400 297.600 ;
        RECT 335.600 295.800 337.400 296.400 ;
        RECT 297.200 294.000 298.400 294.600 ;
        RECT 293.400 292.600 297.200 293.400 ;
        RECT 268.200 292.000 269.000 292.200 ;
        RECT 270.000 292.000 270.800 292.400 ;
        RECT 273.200 292.000 274.000 292.400 ;
        RECT 290.800 292.000 291.600 292.600 ;
        RECT 297.800 292.000 298.400 294.000 ;
        RECT 268.200 291.400 291.600 292.000 ;
        RECT 297.600 291.400 298.400 292.000 ;
        RECT 299.000 294.300 299.800 295.200 ;
        RECT 302.000 294.300 302.800 295.200 ;
        RECT 299.000 293.700 302.800 294.300 ;
        RECT 297.600 289.600 298.200 291.400 ;
        RECT 299.000 290.800 299.800 293.700 ;
        RECT 302.000 293.600 302.800 293.700 ;
        RECT 303.600 294.300 304.400 295.800 ;
        RECT 311.600 294.300 312.400 295.200 ;
        RECT 303.600 293.700 312.400 294.300 ;
        RECT 276.400 289.400 277.200 289.600 ;
        RECT 271.800 289.000 277.200 289.400 ;
        RECT 271.000 288.800 277.200 289.000 ;
        RECT 278.200 289.000 286.800 289.600 ;
        RECT 268.400 288.000 270.000 288.800 ;
        RECT 271.000 288.200 272.400 288.800 ;
        RECT 278.200 288.200 278.800 289.000 ;
        RECT 286.000 288.800 286.800 289.000 ;
        RECT 289.200 289.000 298.200 289.600 ;
        RECT 289.200 288.800 290.000 289.000 ;
        RECT 269.400 287.600 270.000 288.000 ;
        RECT 273.000 287.600 278.800 288.200 ;
        RECT 279.400 287.600 282.000 288.400 ;
        RECT 266.800 286.800 268.800 287.400 ;
        RECT 269.400 286.800 273.600 287.600 ;
        RECT 268.200 286.200 268.800 286.800 ;
        RECT 268.200 285.600 269.200 286.200 ;
        RECT 268.400 282.200 269.200 285.600 ;
        RECT 271.600 282.200 272.400 286.800 ;
        RECT 274.800 282.200 275.600 285.000 ;
        RECT 276.400 282.200 277.200 285.000 ;
        RECT 278.000 282.200 278.800 287.000 ;
        RECT 281.200 282.200 282.000 287.000 ;
        RECT 284.400 282.200 285.200 288.400 ;
        RECT 292.400 287.600 295.000 288.400 ;
        RECT 287.600 286.800 291.800 287.600 ;
        RECT 286.000 282.200 286.800 285.000 ;
        RECT 287.600 282.200 288.400 285.000 ;
        RECT 289.200 282.200 290.000 285.000 ;
        RECT 292.400 282.200 293.200 287.600 ;
        RECT 297.600 287.400 298.200 289.000 ;
        RECT 295.600 286.800 298.200 287.400 ;
        RECT 298.800 290.000 299.800 290.800 ;
        RECT 295.600 282.200 296.400 286.800 ;
        RECT 298.800 282.200 299.600 290.000 ;
        RECT 303.600 282.200 304.400 293.700 ;
        RECT 311.600 293.600 312.400 293.700 ;
        RECT 305.200 292.300 306.000 292.400 ;
        RECT 313.200 292.300 314.000 295.800 ;
        RECT 316.400 293.600 317.200 295.200 ;
        RECT 318.000 294.300 318.800 295.800 ;
        RECT 321.400 295.400 325.000 295.800 ;
        RECT 322.000 294.400 322.800 294.800 ;
        RECT 326.000 294.400 326.600 295.800 ;
        RECT 327.800 295.400 331.400 295.800 ;
        RECT 328.400 294.400 329.200 294.800 ;
        RECT 332.400 294.400 333.000 295.800 ;
        RECT 321.200 294.300 322.800 294.400 ;
        RECT 318.000 293.800 322.800 294.300 ;
        RECT 318.000 293.700 322.000 293.800 ;
        RECT 305.200 291.700 314.000 292.300 ;
        RECT 305.200 291.600 306.000 291.700 ;
        RECT 305.200 288.800 306.000 290.400 ;
        RECT 313.200 282.200 314.000 291.700 ;
        RECT 314.800 288.800 315.600 290.400 ;
        RECT 318.000 282.200 318.800 293.700 ;
        RECT 321.200 293.600 322.000 293.700 ;
        RECT 324.200 293.600 326.800 294.400 ;
        RECT 327.600 293.800 329.200 294.400 ;
        RECT 327.600 293.600 328.400 293.800 ;
        RECT 330.600 293.600 333.200 294.400 ;
        RECT 334.000 293.600 334.800 295.200 ;
        RECT 322.800 291.600 323.600 293.200 ;
        RECT 324.200 290.400 324.800 293.600 ;
        RECT 329.200 291.600 330.000 293.200 ;
        RECT 330.600 292.400 331.200 293.600 ;
        RECT 330.600 291.600 331.600 292.400 ;
        RECT 319.600 288.800 320.400 290.400 ;
        RECT 322.800 289.600 324.800 290.400 ;
        RECT 326.000 290.200 326.800 290.400 ;
        RECT 330.600 290.200 331.200 291.600 ;
        RECT 332.400 290.200 333.200 290.400 ;
        RECT 325.400 289.600 326.800 290.200 ;
        RECT 330.200 289.600 331.200 290.200 ;
        RECT 331.800 289.600 333.200 290.200 ;
        RECT 323.800 282.200 324.600 289.600 ;
        RECT 325.400 288.400 326.000 289.600 ;
        RECT 325.200 287.600 326.000 288.400 ;
        RECT 330.200 282.200 331.000 289.600 ;
        RECT 331.800 288.400 332.400 289.600 ;
        RECT 331.600 287.600 332.400 288.400 ;
        RECT 335.600 282.200 336.400 295.800 ;
        RECT 338.800 295.600 339.600 297.200 ;
        RECT 340.600 294.400 341.200 297.800 ;
        RECT 340.400 293.600 341.200 294.400 ;
        RECT 340.600 292.300 341.200 293.600 ;
        RECT 337.300 291.700 341.200 292.300 ;
        RECT 337.300 290.400 337.900 291.700 ;
        RECT 337.200 288.800 338.000 290.400 ;
        RECT 340.600 290.200 341.200 291.700 ;
        RECT 342.000 292.300 342.800 292.400 ;
        RECT 343.600 292.300 344.400 299.800 ;
        RECT 350.400 294.200 351.200 299.800 ;
        RECT 356.800 294.200 357.600 299.800 ;
        RECT 359.600 297.000 360.400 299.000 ;
        RECT 359.600 294.800 360.200 297.000 ;
        RECT 363.800 296.000 364.600 299.000 ;
        RECT 369.800 298.400 370.600 299.800 ;
        RECT 369.200 297.600 370.600 298.400 ;
        RECT 369.800 296.400 370.600 297.600 ;
        RECT 363.800 295.400 365.400 296.000 ;
        RECT 369.800 295.800 371.600 296.400 ;
        RECT 364.600 295.000 365.400 295.400 ;
        RECT 359.600 294.200 363.800 294.800 ;
        RECT 350.400 293.800 352.200 294.200 ;
        RECT 356.800 293.800 358.600 294.200 ;
        RECT 350.600 293.600 352.200 293.800 ;
        RECT 357.000 293.600 358.600 293.800 ;
        RECT 342.000 291.700 344.400 292.300 ;
        RECT 342.000 290.800 342.800 291.700 ;
        RECT 340.400 289.400 342.200 290.200 ;
        RECT 341.400 282.200 342.200 289.400 ;
        RECT 343.600 288.300 344.400 291.700 ;
        RECT 348.400 291.600 350.000 292.400 ;
        RECT 346.800 289.600 347.600 291.200 ;
        RECT 351.600 290.400 352.200 293.600 ;
        RECT 354.800 291.600 356.400 292.400 ;
        RECT 358.000 290.400 358.600 293.600 ;
        RECT 362.800 293.800 363.800 294.200 ;
        RECT 364.800 294.400 365.400 295.000 ;
        RECT 359.600 291.600 360.400 293.200 ;
        RECT 361.200 291.600 362.000 293.200 ;
        RECT 362.800 293.000 364.200 293.800 ;
        RECT 364.800 293.600 366.800 294.400 ;
        RECT 362.800 291.000 363.400 293.000 ;
        RECT 359.600 290.400 363.400 291.000 ;
        RECT 351.600 289.600 352.400 290.400 ;
        RECT 358.000 289.600 358.800 290.400 ;
        RECT 350.000 288.300 350.800 289.200 ;
        RECT 343.600 287.700 350.800 288.300 ;
        RECT 343.600 282.200 344.400 287.700 ;
        RECT 350.000 287.600 350.800 287.700 ;
        RECT 351.600 287.000 352.200 289.600 ;
        RECT 356.400 287.600 357.200 289.200 ;
        RECT 358.000 287.000 358.600 289.600 ;
        RECT 348.600 286.400 352.200 287.000 ;
        RECT 355.000 286.400 358.600 287.000 ;
        RECT 348.600 286.200 349.200 286.400 ;
        RECT 348.400 282.200 349.200 286.200 ;
        RECT 351.600 286.200 352.200 286.400 ;
        RECT 351.600 282.200 352.400 286.200 ;
        RECT 354.800 282.200 355.600 286.400 ;
        RECT 358.000 286.200 358.600 286.400 ;
        RECT 359.600 287.000 360.200 290.400 ;
        RECT 364.800 289.800 365.400 293.600 ;
        RECT 366.000 290.800 366.800 292.400 ;
        RECT 363.800 289.200 365.400 289.800 ;
        RECT 358.000 282.200 358.800 286.200 ;
        RECT 359.600 283.000 360.400 287.000 ;
        RECT 363.800 284.400 364.600 289.200 ;
        RECT 369.200 288.800 370.000 290.400 ;
        RECT 362.800 283.600 364.600 284.400 ;
        RECT 363.800 282.200 364.600 283.600 ;
        RECT 370.800 282.200 371.600 295.800 ;
        RECT 372.400 293.600 373.200 295.200 ;
        RECT 377.600 294.200 378.400 299.800 ;
        RECT 377.600 293.800 379.400 294.200 ;
        RECT 377.800 293.600 379.400 293.800 ;
        RECT 380.400 293.600 381.200 295.200 ;
        RECT 374.000 289.600 374.800 291.200 ;
        RECT 378.800 290.400 379.400 293.600 ;
        RECT 378.800 289.600 379.600 290.400 ;
        RECT 372.400 288.300 373.200 288.400 ;
        RECT 372.400 287.700 376.300 288.300 ;
        RECT 372.400 287.600 373.200 287.700 ;
        RECT 375.700 287.000 376.300 287.700 ;
        RECT 377.200 287.600 378.000 289.200 ;
        RECT 378.800 287.000 379.400 289.600 ;
        RECT 375.700 286.400 379.400 287.000 ;
        RECT 375.700 286.200 376.400 286.400 ;
        RECT 375.600 282.200 376.400 286.200 ;
        RECT 378.800 286.200 379.400 286.400 ;
        RECT 378.800 282.200 379.600 286.200 ;
        RECT 382.000 282.200 382.800 299.800 ;
        RECT 387.800 298.400 389.400 299.800 ;
        RECT 386.800 297.600 389.400 298.400 ;
        RECT 387.800 295.800 389.400 297.600 ;
        RECT 395.800 298.400 396.600 299.800 ;
        RECT 395.800 297.600 397.200 298.400 ;
        RECT 395.800 296.400 396.600 297.600 ;
        RECT 394.800 295.800 396.600 296.400 ;
        RECT 399.600 296.000 400.400 299.800 ;
        RECT 386.800 293.600 387.600 294.400 ;
        RECT 387.000 293.200 387.600 293.600 ;
        RECT 387.000 292.400 387.800 293.200 ;
        RECT 388.400 292.400 389.000 295.800 ;
        RECT 390.000 292.800 390.800 294.400 ;
        RECT 393.200 293.600 394.000 295.200 ;
        RECT 385.200 290.800 386.000 292.400 ;
        RECT 388.400 291.600 389.200 292.400 ;
        RECT 391.600 292.200 392.400 292.400 ;
        RECT 390.800 291.600 392.400 292.200 ;
        RECT 388.400 291.400 389.000 291.600 ;
        RECT 387.000 290.800 389.000 291.400 ;
        RECT 390.800 291.200 391.600 291.600 ;
        RECT 387.000 290.200 387.600 290.800 ;
        RECT 385.200 282.800 386.000 290.200 ;
        RECT 386.800 283.400 387.600 290.200 ;
        RECT 388.400 289.600 392.400 290.200 ;
        RECT 388.400 282.800 389.200 289.600 ;
        RECT 385.200 282.200 389.200 282.800 ;
        RECT 391.600 282.200 392.400 289.600 ;
        RECT 394.800 282.200 395.600 295.800 ;
        RECT 399.400 295.200 400.400 296.000 ;
        RECT 399.400 290.800 400.200 295.200 ;
        RECT 401.200 294.600 402.000 299.800 ;
        RECT 407.600 296.600 408.400 299.800 ;
        RECT 409.200 297.000 410.000 299.800 ;
        RECT 410.800 297.000 411.600 299.800 ;
        RECT 412.400 297.000 413.200 299.800 ;
        RECT 414.000 297.000 414.800 299.800 ;
        RECT 417.200 297.000 418.000 299.800 ;
        RECT 420.400 297.000 421.200 299.800 ;
        RECT 422.000 297.000 422.800 299.800 ;
        RECT 423.600 297.000 424.400 299.800 ;
        RECT 406.000 295.800 408.400 296.600 ;
        RECT 425.200 296.600 426.000 299.800 ;
        RECT 406.000 295.200 406.800 295.800 ;
        RECT 400.800 294.000 402.000 294.600 ;
        RECT 405.000 294.600 406.800 295.200 ;
        RECT 410.800 295.600 411.800 296.400 ;
        RECT 414.800 295.600 416.400 296.400 ;
        RECT 417.200 295.800 421.800 296.400 ;
        RECT 425.200 295.800 427.800 296.600 ;
        RECT 417.200 295.600 418.000 295.800 ;
        RECT 400.800 292.000 401.400 294.000 ;
        RECT 405.000 293.400 405.800 294.600 ;
        RECT 402.000 292.600 405.800 293.400 ;
        RECT 410.800 292.800 411.600 295.600 ;
        RECT 417.200 294.800 418.000 295.000 ;
        RECT 413.600 294.200 418.000 294.800 ;
        RECT 413.600 294.000 414.400 294.200 ;
        RECT 418.800 293.600 419.600 295.200 ;
        RECT 421.000 293.400 421.800 295.800 ;
        RECT 427.000 295.200 427.800 295.800 ;
        RECT 427.000 294.400 430.000 295.200 ;
        RECT 431.600 293.800 432.400 299.800 ;
        RECT 435.800 298.400 437.400 299.800 ;
        RECT 443.800 298.400 445.400 299.800 ;
        RECT 434.800 297.600 437.400 298.400 ;
        RECT 442.800 297.600 445.400 298.400 ;
        RECT 435.800 295.800 437.400 297.600 ;
        RECT 443.800 295.800 445.400 297.600 ;
        RECT 414.000 292.600 417.200 293.400 ;
        RECT 421.000 292.600 423.000 293.400 ;
        RECT 423.600 293.000 432.400 293.800 ;
        RECT 434.800 293.600 435.600 294.400 ;
        RECT 407.600 292.000 408.400 292.600 ;
        RECT 425.200 292.000 426.000 292.400 ;
        RECT 428.400 292.000 429.200 292.400 ;
        RECT 430.200 292.000 431.000 292.200 ;
        RECT 400.800 291.400 401.600 292.000 ;
        RECT 407.600 291.400 431.000 292.000 ;
        RECT 396.400 290.300 397.200 290.400 ;
        RECT 398.000 290.300 398.800 290.400 ;
        RECT 396.400 289.700 398.800 290.300 ;
        RECT 399.400 290.000 400.400 290.800 ;
        RECT 396.400 288.800 397.200 289.700 ;
        RECT 398.000 289.600 398.800 289.700 ;
        RECT 399.600 282.200 400.400 290.000 ;
        RECT 401.000 289.600 401.600 291.400 ;
        RECT 401.000 289.000 410.000 289.600 ;
        RECT 401.000 287.400 401.600 289.000 ;
        RECT 409.200 288.800 410.000 289.000 ;
        RECT 412.400 289.000 421.000 289.600 ;
        RECT 412.400 288.800 413.200 289.000 ;
        RECT 404.200 287.600 406.800 288.400 ;
        RECT 401.000 286.800 403.600 287.400 ;
        RECT 402.800 282.200 403.600 286.800 ;
        RECT 406.000 282.200 406.800 287.600 ;
        RECT 407.400 286.800 411.600 287.600 ;
        RECT 409.200 282.200 410.000 285.000 ;
        RECT 410.800 282.200 411.600 285.000 ;
        RECT 412.400 282.200 413.200 285.000 ;
        RECT 414.000 282.200 414.800 288.400 ;
        RECT 417.200 287.600 419.800 288.400 ;
        RECT 420.400 288.200 421.000 289.000 ;
        RECT 422.000 289.400 422.800 289.600 ;
        RECT 422.000 289.000 427.400 289.400 ;
        RECT 422.000 288.800 428.200 289.000 ;
        RECT 426.800 288.200 428.200 288.800 ;
        RECT 420.400 287.600 426.200 288.200 ;
        RECT 429.200 288.000 430.800 288.800 ;
        RECT 429.200 287.600 429.800 288.000 ;
        RECT 417.200 282.200 418.000 287.000 ;
        RECT 420.400 282.200 421.200 287.000 ;
        RECT 425.600 286.800 429.800 287.600 ;
        RECT 431.600 287.400 432.400 293.000 ;
        RECT 435.000 293.200 435.600 293.600 ;
        RECT 435.000 292.400 435.800 293.200 ;
        RECT 436.400 292.400 437.000 295.800 ;
        RECT 438.000 292.800 438.800 294.400 ;
        RECT 442.800 293.600 443.600 294.400 ;
        RECT 443.000 293.200 443.600 293.600 ;
        RECT 443.000 292.400 443.800 293.200 ;
        RECT 444.400 292.400 445.000 295.800 ;
        RECT 446.000 294.300 446.800 294.400 ;
        RECT 447.600 294.300 448.400 294.400 ;
        RECT 446.000 293.700 448.400 294.300 ;
        RECT 446.000 292.800 446.800 293.700 ;
        RECT 447.600 293.600 448.400 293.700 ;
        RECT 433.200 290.800 434.000 292.400 ;
        RECT 436.400 291.600 437.200 292.400 ;
        RECT 439.600 292.200 440.400 292.400 ;
        RECT 438.800 291.600 440.400 292.200 ;
        RECT 436.400 291.400 437.000 291.600 ;
        RECT 435.000 290.800 437.000 291.400 ;
        RECT 438.800 291.200 439.600 291.600 ;
        RECT 441.200 290.800 442.000 292.400 ;
        RECT 444.400 291.600 445.200 292.400 ;
        RECT 447.600 292.300 448.400 292.400 ;
        RECT 449.200 292.300 450.000 299.800 ;
        RECT 450.800 295.600 451.600 297.200 ;
        RECT 450.800 294.300 451.600 294.400 ;
        RECT 452.400 294.300 453.200 299.800 ;
        RECT 454.000 296.300 454.800 297.200 ;
        RECT 458.800 296.300 459.600 296.400 ;
        RECT 454.000 295.700 459.600 296.300 ;
        RECT 454.000 295.600 454.800 295.700 ;
        RECT 458.800 295.600 459.600 295.700 ;
        RECT 464.000 294.400 464.800 299.800 ;
        RECT 450.800 293.700 453.200 294.300 ;
        RECT 450.800 293.600 451.600 293.700 ;
        RECT 447.600 292.200 450.000 292.300 ;
        RECT 446.800 291.700 450.000 292.200 ;
        RECT 446.800 291.600 448.400 291.700 ;
        RECT 444.400 291.400 445.000 291.600 ;
        RECT 443.000 290.800 445.000 291.400 ;
        RECT 446.800 291.200 447.600 291.600 ;
        RECT 435.000 290.200 435.600 290.800 ;
        RECT 443.000 290.200 443.600 290.800 ;
        RECT 430.400 286.800 432.400 287.400 ;
        RECT 422.000 282.200 422.800 285.000 ;
        RECT 423.600 282.200 424.400 285.000 ;
        RECT 426.800 282.200 427.600 286.800 ;
        RECT 430.400 286.200 431.000 286.800 ;
        RECT 430.000 285.600 431.000 286.200 ;
        RECT 430.000 282.200 430.800 285.600 ;
        RECT 433.200 282.800 434.000 290.200 ;
        RECT 434.800 283.400 435.600 290.200 ;
        RECT 436.400 289.600 440.400 290.200 ;
        RECT 436.400 282.800 437.200 289.600 ;
        RECT 433.200 282.200 437.200 282.800 ;
        RECT 439.600 282.200 440.400 289.600 ;
        RECT 441.200 282.800 442.000 290.200 ;
        RECT 442.800 283.400 443.600 290.200 ;
        RECT 444.400 289.600 448.400 290.200 ;
        RECT 444.400 282.800 445.200 289.600 ;
        RECT 441.200 282.200 445.200 282.800 ;
        RECT 447.600 282.200 448.400 289.600 ;
        RECT 449.200 282.200 450.000 291.700 ;
        RECT 452.400 282.200 453.200 293.700 ;
        RECT 463.600 294.200 464.800 294.400 ;
        RECT 470.400 294.200 471.200 299.800 ;
        RECT 476.400 295.800 477.200 299.800 ;
        RECT 477.800 296.400 478.600 297.200 ;
        RECT 480.200 296.400 481.000 299.800 ;
        RECT 463.600 293.600 465.800 294.200 ;
        RECT 470.400 293.800 472.200 294.200 ;
        RECT 470.600 293.600 472.200 293.800 ;
        RECT 462.000 291.600 463.600 292.400 ;
        RECT 460.400 289.600 461.200 291.200 ;
        RECT 465.200 290.400 465.800 293.600 ;
        RECT 468.400 291.600 470.000 292.400 ;
        RECT 465.200 289.600 466.000 290.400 ;
        RECT 466.800 289.600 467.600 291.200 ;
        RECT 471.600 290.400 472.200 293.600 ;
        RECT 474.800 292.800 475.600 294.400 ;
        RECT 473.200 292.200 474.000 292.400 ;
        RECT 476.400 292.200 477.000 295.800 ;
        RECT 478.000 295.600 478.800 296.400 ;
        RECT 480.200 295.800 482.000 296.400 ;
        RECT 479.600 294.300 480.400 294.400 ;
        RECT 481.200 294.300 482.000 295.800 ;
        RECT 487.600 295.800 488.400 299.800 ;
        RECT 492.400 297.800 493.200 299.800 ;
        RECT 498.200 298.400 499.000 299.800 ;
        RECT 489.000 296.400 489.800 297.200 ;
        RECT 479.600 293.700 482.000 294.300 ;
        RECT 479.600 293.600 480.400 293.700 ;
        RECT 478.000 292.200 478.800 292.400 ;
        RECT 473.200 291.600 474.800 292.200 ;
        RECT 476.400 291.600 478.800 292.200 ;
        RECT 474.000 291.200 474.800 291.600 ;
        RECT 471.600 289.600 472.400 290.400 ;
        RECT 478.000 290.200 478.600 291.600 ;
        RECT 473.200 289.600 477.200 290.200 ;
        RECT 463.600 287.600 464.400 289.200 ;
        RECT 465.200 287.000 465.800 289.600 ;
        RECT 466.800 288.300 467.600 288.400 ;
        RECT 470.000 288.300 470.800 289.200 ;
        RECT 466.800 287.700 470.800 288.300 ;
        RECT 466.800 287.600 467.600 287.700 ;
        RECT 470.000 287.600 470.800 287.700 ;
        RECT 471.600 287.000 472.200 289.600 ;
        RECT 462.200 286.400 465.800 287.000 ;
        RECT 462.200 286.200 462.800 286.400 ;
        RECT 462.000 282.200 462.800 286.200 ;
        RECT 465.200 286.200 465.800 286.400 ;
        RECT 468.600 286.400 472.200 287.000 ;
        RECT 468.600 286.200 469.200 286.400 ;
        RECT 465.200 282.200 466.000 286.200 ;
        RECT 468.400 282.200 469.200 286.200 ;
        RECT 471.600 286.200 472.200 286.400 ;
        RECT 471.600 282.200 472.400 286.200 ;
        RECT 473.200 282.200 474.000 289.600 ;
        RECT 476.400 282.200 477.200 289.600 ;
        RECT 478.000 282.200 478.800 290.200 ;
        RECT 479.600 288.800 480.400 290.400 ;
        RECT 481.200 282.200 482.000 293.700 ;
        RECT 482.800 293.600 483.600 295.200 ;
        RECT 486.000 292.800 486.800 294.400 ;
        RECT 484.400 292.200 485.200 292.400 ;
        RECT 487.600 292.200 488.200 295.800 ;
        RECT 489.200 295.600 490.000 296.400 ;
        RECT 490.800 295.600 491.600 297.200 ;
        RECT 489.300 294.300 489.900 295.600 ;
        RECT 492.600 294.400 493.200 297.800 ;
        RECT 497.200 297.600 499.000 298.400 ;
        RECT 498.200 296.400 499.000 297.600 ;
        RECT 497.200 295.800 499.000 296.400 ;
        RECT 500.400 295.800 501.200 299.800 ;
        RECT 502.000 296.000 502.800 299.800 ;
        RECT 505.200 296.000 506.000 299.800 ;
        RECT 502.000 295.800 506.000 296.000 ;
        RECT 506.800 296.000 507.600 299.800 ;
        RECT 510.000 296.000 510.800 299.800 ;
        RECT 506.800 295.800 510.800 296.000 ;
        RECT 511.600 295.800 512.400 299.800 ;
        RECT 515.800 296.400 516.600 299.800 ;
        RECT 514.800 295.800 516.600 296.400 ;
        RECT 519.600 297.800 520.400 299.800 ;
        RECT 524.400 297.800 525.200 299.800 ;
        RECT 490.800 294.300 491.600 294.400 ;
        RECT 489.300 293.700 491.600 294.300 ;
        RECT 490.800 293.600 491.600 293.700 ;
        RECT 492.400 293.600 493.200 294.400 ;
        RECT 495.600 293.600 496.400 295.200 ;
        RECT 489.200 292.200 490.000 292.400 ;
        RECT 484.400 291.600 486.000 292.200 ;
        RECT 487.600 291.600 490.000 292.200 ;
        RECT 485.200 291.200 486.000 291.600 ;
        RECT 489.200 290.200 489.800 291.600 ;
        RECT 492.600 290.200 493.200 293.600 ;
        RECT 494.000 290.800 494.800 292.400 ;
        RECT 484.400 289.600 488.400 290.200 ;
        RECT 484.400 282.200 485.200 289.600 ;
        RECT 487.600 282.200 488.400 289.600 ;
        RECT 489.200 282.200 490.000 290.200 ;
        RECT 492.400 289.400 494.200 290.200 ;
        RECT 493.400 288.300 494.200 289.400 ;
        RECT 495.600 288.300 496.400 288.400 ;
        RECT 493.400 287.700 496.400 288.300 ;
        RECT 493.400 282.200 494.200 287.700 ;
        RECT 495.600 287.600 496.400 287.700 ;
        RECT 497.200 282.200 498.000 295.800 ;
        RECT 500.600 294.400 501.200 295.800 ;
        RECT 502.200 295.400 505.800 295.800 ;
        RECT 507.000 295.400 510.600 295.800 ;
        RECT 504.400 294.400 505.200 294.800 ;
        RECT 507.600 294.400 508.400 294.800 ;
        RECT 511.600 294.400 512.200 295.800 ;
        RECT 500.400 293.600 503.000 294.400 ;
        RECT 504.400 294.300 506.000 294.400 ;
        RECT 506.800 294.300 508.400 294.400 ;
        RECT 504.400 293.800 508.400 294.300 ;
        RECT 505.200 293.700 507.600 293.800 ;
        RECT 505.200 293.600 506.000 293.700 ;
        RECT 506.800 293.600 507.600 293.700 ;
        RECT 509.800 293.600 512.400 294.400 ;
        RECT 513.200 293.600 514.000 295.200 ;
        RECT 498.800 292.300 499.600 292.400 ;
        RECT 502.400 292.300 503.000 293.600 ;
        RECT 498.800 291.700 503.000 292.300 ;
        RECT 498.800 291.600 499.600 291.700 ;
        RECT 498.800 288.800 499.600 290.400 ;
        RECT 500.400 290.200 501.200 290.400 ;
        RECT 502.400 290.200 503.000 291.700 ;
        RECT 503.600 292.300 504.400 293.200 ;
        RECT 508.400 292.300 509.200 293.200 ;
        RECT 503.600 291.700 509.200 292.300 ;
        RECT 503.600 291.600 504.400 291.700 ;
        RECT 508.400 291.600 509.200 291.700 ;
        RECT 509.800 290.200 510.400 293.600 ;
        RECT 511.600 290.300 512.400 290.400 ;
        RECT 514.800 290.300 515.600 295.800 ;
        RECT 519.600 294.400 520.200 297.800 ;
        RECT 521.200 295.600 522.000 297.200 ;
        RECT 522.800 295.600 523.600 297.200 ;
        RECT 524.600 294.400 525.200 297.800 ;
        RECT 519.600 293.600 520.400 294.400 ;
        RECT 524.400 293.600 525.200 294.400 ;
        RECT 526.000 294.300 526.800 294.400 ;
        RECT 527.600 294.300 528.400 295.200 ;
        RECT 526.000 293.700 528.400 294.300 ;
        RECT 526.000 293.600 526.800 293.700 ;
        RECT 527.600 293.600 528.400 293.700 ;
        RECT 518.000 290.800 518.800 292.400 ;
        RECT 511.600 290.200 515.600 290.300 ;
        RECT 500.400 289.600 501.800 290.200 ;
        RECT 502.400 289.600 503.400 290.200 ;
        RECT 501.200 288.400 501.800 289.600 ;
        RECT 501.200 287.600 502.000 288.400 ;
        RECT 502.600 282.200 503.400 289.600 ;
        RECT 509.400 289.600 510.400 290.200 ;
        RECT 511.000 289.700 515.600 290.200 ;
        RECT 511.000 289.600 512.400 289.700 ;
        RECT 509.400 282.200 510.200 289.600 ;
        RECT 511.000 288.400 511.600 289.600 ;
        RECT 510.800 287.600 511.600 288.400 ;
        RECT 514.800 282.200 515.600 289.700 ;
        RECT 516.400 288.800 517.200 290.400 ;
        RECT 519.600 290.200 520.200 293.600 ;
        RECT 524.600 290.200 525.200 293.600 ;
        RECT 526.000 290.800 526.800 292.400 ;
        RECT 518.600 289.400 520.400 290.200 ;
        RECT 524.400 289.400 526.200 290.200 ;
        RECT 518.600 284.400 519.400 289.400 ;
        RECT 525.400 284.400 526.200 289.400 ;
        RECT 518.600 283.600 520.400 284.400 ;
        RECT 525.400 283.600 526.800 284.400 ;
        RECT 518.600 282.200 519.400 283.600 ;
        RECT 525.400 282.200 526.200 283.600 ;
        RECT 529.200 282.200 530.000 299.800 ;
        RECT 530.800 295.800 531.600 299.800 ;
        RECT 532.400 296.000 533.200 299.800 ;
        RECT 535.600 296.000 536.400 299.800 ;
        RECT 538.800 296.000 539.600 299.800 ;
        RECT 532.400 295.800 536.400 296.000 ;
        RECT 531.000 294.400 531.600 295.800 ;
        RECT 532.600 295.400 536.200 295.800 ;
        RECT 538.600 295.200 539.600 296.000 ;
        RECT 534.800 294.400 535.600 294.800 ;
        RECT 530.800 293.600 533.400 294.400 ;
        RECT 534.800 293.800 536.400 294.400 ;
        RECT 535.600 293.600 536.400 293.800 ;
        RECT 530.800 290.200 531.600 290.400 ;
        RECT 532.800 290.200 533.400 293.600 ;
        RECT 534.000 291.600 534.800 293.200 ;
        RECT 538.600 290.800 539.400 295.200 ;
        RECT 540.400 294.600 541.200 299.800 ;
        RECT 546.800 296.600 547.600 299.800 ;
        RECT 548.400 297.000 549.200 299.800 ;
        RECT 550.000 297.000 550.800 299.800 ;
        RECT 551.600 297.000 552.400 299.800 ;
        RECT 553.200 297.000 554.000 299.800 ;
        RECT 556.400 297.000 557.200 299.800 ;
        RECT 559.600 297.000 560.400 299.800 ;
        RECT 561.200 297.000 562.000 299.800 ;
        RECT 562.800 297.000 563.600 299.800 ;
        RECT 545.200 295.800 547.600 296.600 ;
        RECT 564.400 296.600 565.200 299.800 ;
        RECT 545.200 295.200 546.000 295.800 ;
        RECT 540.000 294.000 541.200 294.600 ;
        RECT 544.200 294.600 546.000 295.200 ;
        RECT 550.000 295.600 551.000 296.400 ;
        RECT 554.000 295.600 555.600 296.400 ;
        RECT 556.400 295.800 561.000 296.400 ;
        RECT 564.400 295.800 567.000 296.600 ;
        RECT 556.400 295.600 557.200 295.800 ;
        RECT 540.000 292.000 540.600 294.000 ;
        RECT 544.200 293.400 545.000 294.600 ;
        RECT 541.200 292.600 545.000 293.400 ;
        RECT 550.000 292.800 550.800 295.600 ;
        RECT 556.400 294.800 557.200 295.000 ;
        RECT 552.800 294.200 557.200 294.800 ;
        RECT 552.800 294.000 553.600 294.200 ;
        RECT 558.000 293.600 558.800 295.200 ;
        RECT 560.200 293.400 561.000 295.800 ;
        RECT 566.200 295.200 567.000 295.800 ;
        RECT 566.200 294.400 569.200 295.200 ;
        RECT 570.800 293.800 571.600 299.800 ;
        RECT 575.000 298.400 575.800 299.800 ;
        RECT 575.000 297.600 576.400 298.400 ;
        RECT 575.000 296.400 575.800 297.600 ;
        RECT 574.000 295.800 575.800 296.400 ;
        RECT 553.200 292.600 556.400 293.400 ;
        RECT 560.200 292.600 562.200 293.400 ;
        RECT 562.800 293.000 571.600 293.800 ;
        RECT 572.400 293.600 573.200 295.200 ;
        RECT 546.800 292.000 547.600 292.600 ;
        RECT 558.000 292.000 558.800 292.400 ;
        RECT 564.400 292.000 565.200 292.400 ;
        RECT 569.200 292.200 570.000 292.400 ;
        RECT 569.200 292.000 570.200 292.200 ;
        RECT 540.000 291.400 540.800 292.000 ;
        RECT 546.800 291.400 570.200 292.000 ;
        RECT 530.800 289.600 532.200 290.200 ;
        RECT 532.800 289.600 533.800 290.200 ;
        RECT 538.600 290.000 539.600 290.800 ;
        RECT 531.600 288.400 532.200 289.600 ;
        RECT 531.600 287.600 532.400 288.400 ;
        RECT 533.000 282.200 533.800 289.600 ;
        RECT 538.800 282.200 539.600 290.000 ;
        RECT 540.200 289.600 540.800 291.400 ;
        RECT 540.200 289.000 549.200 289.600 ;
        RECT 540.200 287.400 540.800 289.000 ;
        RECT 548.400 288.800 549.200 289.000 ;
        RECT 551.600 289.000 560.200 289.600 ;
        RECT 551.600 288.800 552.400 289.000 ;
        RECT 543.400 287.600 546.000 288.400 ;
        RECT 540.200 286.800 542.800 287.400 ;
        RECT 542.000 282.200 542.800 286.800 ;
        RECT 545.200 282.200 546.000 287.600 ;
        RECT 546.600 286.800 550.800 287.600 ;
        RECT 548.400 282.200 549.200 285.000 ;
        RECT 550.000 282.200 550.800 285.000 ;
        RECT 551.600 282.200 552.400 285.000 ;
        RECT 553.200 282.200 554.000 288.400 ;
        RECT 556.400 287.600 559.000 288.400 ;
        RECT 559.600 288.200 560.200 289.000 ;
        RECT 561.200 289.400 562.000 289.600 ;
        RECT 561.200 289.000 566.600 289.400 ;
        RECT 561.200 288.800 567.400 289.000 ;
        RECT 566.000 288.200 567.400 288.800 ;
        RECT 559.600 287.600 565.400 288.200 ;
        RECT 568.400 288.000 570.000 288.800 ;
        RECT 568.400 287.600 569.000 288.000 ;
        RECT 556.400 282.200 557.200 287.000 ;
        RECT 559.600 282.200 560.400 287.000 ;
        RECT 564.800 286.800 569.000 287.600 ;
        RECT 570.800 287.400 571.600 293.000 ;
        RECT 569.600 286.800 571.600 287.400 ;
        RECT 561.200 282.200 562.000 285.000 ;
        RECT 562.800 282.200 563.600 285.000 ;
        RECT 566.000 282.200 566.800 286.800 ;
        RECT 569.600 286.200 570.200 286.800 ;
        RECT 569.200 285.600 570.200 286.200 ;
        RECT 569.200 282.200 570.000 285.600 ;
        RECT 574.000 282.200 574.800 295.800 ;
        RECT 577.200 293.800 578.000 299.800 ;
        RECT 583.600 296.600 584.400 299.800 ;
        RECT 585.200 297.000 586.000 299.800 ;
        RECT 586.800 297.000 587.600 299.800 ;
        RECT 588.400 297.000 589.200 299.800 ;
        RECT 591.600 297.000 592.400 299.800 ;
        RECT 594.800 297.000 595.600 299.800 ;
        RECT 596.400 297.000 597.200 299.800 ;
        RECT 598.000 297.000 598.800 299.800 ;
        RECT 599.600 297.000 600.400 299.800 ;
        RECT 581.800 295.800 584.400 296.600 ;
        RECT 601.200 296.600 602.000 299.800 ;
        RECT 587.800 295.800 592.400 296.400 ;
        RECT 581.800 295.200 582.600 295.800 ;
        RECT 579.600 294.400 582.600 295.200 ;
        RECT 577.200 293.000 586.000 293.800 ;
        RECT 587.800 293.400 588.600 295.800 ;
        RECT 591.600 295.600 592.400 295.800 ;
        RECT 593.200 295.600 594.800 296.400 ;
        RECT 597.800 295.600 598.800 296.400 ;
        RECT 601.200 295.800 603.600 296.600 ;
        RECT 590.000 293.600 590.800 295.200 ;
        RECT 591.600 294.800 592.400 295.000 ;
        RECT 591.600 294.200 596.000 294.800 ;
        RECT 595.200 294.000 596.000 294.200 ;
        RECT 575.600 288.800 576.400 290.400 ;
        RECT 577.200 287.400 578.000 293.000 ;
        RECT 586.600 292.600 588.600 293.400 ;
        RECT 592.400 292.600 595.600 293.400 ;
        RECT 598.000 292.800 598.800 295.600 ;
        RECT 602.800 295.200 603.600 295.800 ;
        RECT 602.800 294.600 604.600 295.200 ;
        RECT 603.800 293.400 604.600 294.600 ;
        RECT 607.600 294.600 608.400 299.800 ;
        RECT 609.200 296.000 610.000 299.800 ;
        RECT 609.200 295.200 610.200 296.000 ;
        RECT 607.600 294.000 608.800 294.600 ;
        RECT 603.800 292.600 607.600 293.400 ;
        RECT 578.800 292.200 579.600 292.400 ;
        RECT 578.600 292.000 579.600 292.200 ;
        RECT 583.600 292.000 584.400 292.400 ;
        RECT 601.200 292.000 602.000 292.600 ;
        RECT 608.200 292.000 608.800 294.000 ;
        RECT 578.600 291.400 602.000 292.000 ;
        RECT 608.000 291.400 608.800 292.000 ;
        RECT 608.000 289.600 608.600 291.400 ;
        RECT 609.400 290.800 610.200 295.200 ;
        RECT 586.800 289.400 587.600 289.600 ;
        RECT 582.200 289.000 587.600 289.400 ;
        RECT 581.400 288.800 587.600 289.000 ;
        RECT 588.600 289.000 597.200 289.600 ;
        RECT 578.800 288.000 580.400 288.800 ;
        RECT 581.400 288.200 582.800 288.800 ;
        RECT 588.600 288.200 589.200 289.000 ;
        RECT 596.400 288.800 597.200 289.000 ;
        RECT 599.600 289.000 608.600 289.600 ;
        RECT 599.600 288.800 600.400 289.000 ;
        RECT 579.800 287.600 580.400 288.000 ;
        RECT 583.400 287.600 589.200 288.200 ;
        RECT 589.800 287.600 592.400 288.400 ;
        RECT 577.200 286.800 579.200 287.400 ;
        RECT 579.800 286.800 584.000 287.600 ;
        RECT 578.600 286.200 579.200 286.800 ;
        RECT 578.600 285.600 579.600 286.200 ;
        RECT 578.800 282.200 579.600 285.600 ;
        RECT 582.000 282.200 582.800 286.800 ;
        RECT 585.200 282.200 586.000 285.000 ;
        RECT 586.800 282.200 587.600 285.000 ;
        RECT 588.400 282.200 589.200 287.000 ;
        RECT 591.600 282.200 592.400 287.000 ;
        RECT 594.800 282.200 595.600 288.400 ;
        RECT 602.800 287.600 605.400 288.400 ;
        RECT 598.000 286.800 602.200 287.600 ;
        RECT 596.400 282.200 597.200 285.000 ;
        RECT 598.000 282.200 598.800 285.000 ;
        RECT 599.600 282.200 600.400 285.000 ;
        RECT 602.800 282.200 603.600 287.600 ;
        RECT 608.000 287.400 608.600 289.000 ;
        RECT 606.000 286.800 608.600 287.400 ;
        RECT 609.200 290.000 610.200 290.800 ;
        RECT 606.000 282.200 606.800 286.800 ;
        RECT 609.200 282.200 610.000 290.000 ;
        RECT 2.800 276.400 3.600 279.800 ;
        RECT 2.600 275.800 3.600 276.400 ;
        RECT 2.600 275.200 3.200 275.800 ;
        RECT 6.000 275.200 6.800 279.800 ;
        RECT 9.200 277.000 10.000 279.800 ;
        RECT 10.800 277.000 11.600 279.800 ;
        RECT 1.200 274.600 3.200 275.200 ;
        RECT 1.200 269.000 2.000 274.600 ;
        RECT 3.800 274.400 8.000 275.200 ;
        RECT 12.400 275.000 13.200 279.800 ;
        RECT 15.600 275.000 16.400 279.800 ;
        RECT 3.800 274.000 4.400 274.400 ;
        RECT 2.800 273.200 4.400 274.000 ;
        RECT 7.400 273.800 13.200 274.400 ;
        RECT 5.400 273.200 6.800 273.800 ;
        RECT 5.400 273.000 11.600 273.200 ;
        RECT 6.200 272.600 11.600 273.000 ;
        RECT 10.800 272.400 11.600 272.600 ;
        RECT 12.600 273.000 13.200 273.800 ;
        RECT 13.800 273.600 16.400 274.400 ;
        RECT 18.800 273.600 19.600 279.800 ;
        RECT 20.400 277.000 21.200 279.800 ;
        RECT 22.000 277.000 22.800 279.800 ;
        RECT 23.600 277.000 24.400 279.800 ;
        RECT 22.000 274.400 26.200 275.200 ;
        RECT 26.800 274.400 27.600 279.800 ;
        RECT 30.000 275.200 30.800 279.800 ;
        RECT 30.000 274.600 32.600 275.200 ;
        RECT 26.800 273.600 29.400 274.400 ;
        RECT 20.400 273.000 21.200 273.200 ;
        RECT 12.600 272.400 21.200 273.000 ;
        RECT 23.600 273.000 24.400 273.200 ;
        RECT 32.000 273.000 32.600 274.600 ;
        RECT 23.600 272.400 32.600 273.000 ;
        RECT 32.000 270.600 32.600 272.400 ;
        RECT 33.200 272.000 34.000 279.800 ;
        RECT 38.000 272.000 38.800 279.800 ;
        RECT 41.200 275.200 42.000 279.800 ;
        RECT 33.200 271.200 34.200 272.000 ;
        RECT 2.600 270.000 26.000 270.600 ;
        RECT 32.000 270.000 32.800 270.600 ;
        RECT 2.600 269.800 3.400 270.000 ;
        RECT 7.600 269.600 8.400 270.000 ;
        RECT 25.200 269.400 26.000 270.000 ;
        RECT 1.200 268.200 10.000 269.000 ;
        RECT 10.600 268.600 12.600 269.400 ;
        RECT 16.400 268.600 19.600 269.400 ;
        RECT 1.200 262.200 2.000 268.200 ;
        RECT 3.600 266.800 6.600 267.600 ;
        RECT 5.800 266.200 6.600 266.800 ;
        RECT 11.800 266.200 12.600 268.600 ;
        RECT 14.000 266.800 14.800 268.400 ;
        RECT 19.200 267.800 20.000 268.000 ;
        RECT 15.600 267.200 20.000 267.800 ;
        RECT 15.600 267.000 16.400 267.200 ;
        RECT 22.000 266.400 22.800 269.200 ;
        RECT 27.800 268.600 31.600 269.400 ;
        RECT 27.800 267.400 28.600 268.600 ;
        RECT 32.200 268.000 32.800 270.000 ;
        RECT 15.600 266.200 16.400 266.400 ;
        RECT 5.800 265.400 8.400 266.200 ;
        RECT 11.800 265.600 16.400 266.200 ;
        RECT 17.200 265.600 18.800 266.400 ;
        RECT 21.800 265.600 22.800 266.400 ;
        RECT 26.800 266.800 28.600 267.400 ;
        RECT 31.600 267.400 32.800 268.000 ;
        RECT 26.800 266.200 27.600 266.800 ;
        RECT 7.600 262.200 8.400 265.400 ;
        RECT 25.200 265.400 27.600 266.200 ;
        RECT 9.200 262.200 10.000 265.000 ;
        RECT 10.800 262.200 11.600 265.000 ;
        RECT 12.400 262.200 13.200 265.000 ;
        RECT 15.600 262.200 16.400 265.000 ;
        RECT 18.800 262.200 19.600 265.000 ;
        RECT 20.400 262.200 21.200 265.000 ;
        RECT 22.000 262.200 22.800 265.000 ;
        RECT 23.600 262.200 24.400 265.000 ;
        RECT 25.200 262.200 26.000 265.400 ;
        RECT 31.600 262.200 32.400 267.400 ;
        RECT 33.400 266.800 34.200 271.200 ;
        RECT 33.200 266.000 34.200 266.800 ;
        RECT 37.800 271.200 38.800 272.000 ;
        RECT 39.400 274.600 42.000 275.200 ;
        RECT 39.400 273.000 40.000 274.600 ;
        RECT 44.400 274.400 45.200 279.800 ;
        RECT 47.600 277.000 48.400 279.800 ;
        RECT 49.200 277.000 50.000 279.800 ;
        RECT 50.800 277.000 51.600 279.800 ;
        RECT 45.800 274.400 50.000 275.200 ;
        RECT 42.600 273.600 45.200 274.400 ;
        RECT 52.400 273.600 53.200 279.800 ;
        RECT 55.600 275.000 56.400 279.800 ;
        RECT 58.800 275.000 59.600 279.800 ;
        RECT 60.400 277.000 61.200 279.800 ;
        RECT 62.000 277.000 62.800 279.800 ;
        RECT 65.200 275.200 66.000 279.800 ;
        RECT 68.400 276.400 69.200 279.800 ;
        RECT 68.400 275.800 69.400 276.400 ;
        RECT 68.800 275.200 69.400 275.800 ;
        RECT 64.000 274.400 68.200 275.200 ;
        RECT 68.800 274.600 70.800 275.200 ;
        RECT 55.600 273.600 58.200 274.400 ;
        RECT 58.800 273.800 64.600 274.400 ;
        RECT 67.600 274.000 68.200 274.400 ;
        RECT 47.600 273.000 48.400 273.200 ;
        RECT 39.400 272.400 48.400 273.000 ;
        RECT 50.800 273.000 51.600 273.200 ;
        RECT 58.800 273.000 59.400 273.800 ;
        RECT 65.200 273.200 66.600 273.800 ;
        RECT 67.600 273.200 69.200 274.000 ;
        RECT 50.800 272.400 59.400 273.000 ;
        RECT 60.400 273.000 66.600 273.200 ;
        RECT 60.400 272.600 65.800 273.000 ;
        RECT 60.400 272.400 61.200 272.600 ;
        RECT 37.800 266.800 38.600 271.200 ;
        RECT 39.400 270.600 40.000 272.400 ;
        RECT 39.200 270.000 40.000 270.600 ;
        RECT 46.000 270.000 69.400 270.600 ;
        RECT 39.200 268.000 39.800 270.000 ;
        RECT 46.000 269.400 46.800 270.000 ;
        RECT 63.600 269.600 64.400 270.000 ;
        RECT 65.200 269.600 66.000 270.000 ;
        RECT 68.600 269.800 69.400 270.000 ;
        RECT 40.400 268.600 44.200 269.400 ;
        RECT 39.200 267.400 40.400 268.000 ;
        RECT 37.800 266.000 38.800 266.800 ;
        RECT 33.200 262.200 34.000 266.000 ;
        RECT 38.000 262.200 38.800 266.000 ;
        RECT 39.600 262.200 40.400 267.400 ;
        RECT 43.400 267.400 44.200 268.600 ;
        RECT 43.400 266.800 45.200 267.400 ;
        RECT 44.400 266.200 45.200 266.800 ;
        RECT 49.200 266.400 50.000 269.200 ;
        RECT 52.400 268.600 55.600 269.400 ;
        RECT 59.400 268.600 61.400 269.400 ;
        RECT 70.000 269.000 70.800 274.600 ;
        RECT 74.200 272.600 75.000 279.800 ;
        RECT 73.200 271.800 75.000 272.600 ;
        RECT 76.400 271.800 77.200 279.800 ;
        RECT 78.000 272.400 78.800 279.800 ;
        RECT 81.200 272.400 82.000 279.800 ;
        RECT 78.000 271.800 82.000 272.400 ;
        RECT 84.400 272.000 85.200 279.800 ;
        RECT 87.600 275.200 88.400 279.800 ;
        RECT 52.000 267.800 52.800 268.000 ;
        RECT 52.000 267.200 56.400 267.800 ;
        RECT 55.600 267.000 56.400 267.200 ;
        RECT 57.200 266.800 58.000 268.400 ;
        RECT 44.400 265.400 46.800 266.200 ;
        RECT 49.200 265.600 50.200 266.400 ;
        RECT 53.200 265.600 54.800 266.400 ;
        RECT 55.600 266.200 56.400 266.400 ;
        RECT 59.400 266.200 60.200 268.600 ;
        RECT 62.000 268.200 70.800 269.000 ;
        RECT 73.400 268.400 74.000 271.800 ;
        RECT 74.800 269.600 75.600 271.200 ;
        RECT 76.600 270.400 77.200 271.800 ;
        RECT 84.200 271.200 85.200 272.000 ;
        RECT 85.800 274.600 88.400 275.200 ;
        RECT 85.800 273.000 86.400 274.600 ;
        RECT 90.800 274.400 91.600 279.800 ;
        RECT 94.000 277.000 94.800 279.800 ;
        RECT 95.600 277.000 96.400 279.800 ;
        RECT 97.200 277.000 98.000 279.800 ;
        RECT 92.200 274.400 96.400 275.200 ;
        RECT 89.000 273.600 91.600 274.400 ;
        RECT 98.800 273.600 99.600 279.800 ;
        RECT 102.000 275.000 102.800 279.800 ;
        RECT 105.200 275.000 106.000 279.800 ;
        RECT 106.800 277.000 107.600 279.800 ;
        RECT 108.400 277.000 109.200 279.800 ;
        RECT 111.600 275.200 112.400 279.800 ;
        RECT 114.800 276.400 115.600 279.800 ;
        RECT 114.800 275.800 115.800 276.400 ;
        RECT 115.200 275.200 115.800 275.800 ;
        RECT 110.400 274.400 114.600 275.200 ;
        RECT 115.200 274.600 117.200 275.200 ;
        RECT 102.000 273.600 104.600 274.400 ;
        RECT 105.200 273.800 111.000 274.400 ;
        RECT 114.000 274.000 114.600 274.400 ;
        RECT 94.000 273.000 94.800 273.200 ;
        RECT 85.800 272.400 94.800 273.000 ;
        RECT 97.200 273.000 98.000 273.200 ;
        RECT 105.200 273.000 105.800 273.800 ;
        RECT 111.600 273.200 113.000 273.800 ;
        RECT 114.000 273.200 115.600 274.000 ;
        RECT 97.200 272.400 105.800 273.000 ;
        RECT 106.800 273.000 113.000 273.200 ;
        RECT 106.800 272.600 112.200 273.000 ;
        RECT 106.800 272.400 107.600 272.600 ;
        RECT 80.400 270.400 81.200 270.800 ;
        RECT 76.400 269.800 78.800 270.400 ;
        RECT 80.400 269.800 82.000 270.400 ;
        RECT 76.400 269.600 77.200 269.800 ;
        RECT 65.400 266.800 68.400 267.600 ;
        RECT 65.400 266.200 66.200 266.800 ;
        RECT 55.600 265.600 60.200 266.200 ;
        RECT 46.000 262.200 46.800 265.400 ;
        RECT 63.600 265.400 66.200 266.200 ;
        RECT 47.600 262.200 48.400 265.000 ;
        RECT 49.200 262.200 50.000 265.000 ;
        RECT 50.800 262.200 51.600 265.000 ;
        RECT 52.400 262.200 53.200 265.000 ;
        RECT 55.600 262.200 56.400 265.000 ;
        RECT 58.800 262.200 59.600 265.000 ;
        RECT 60.400 262.200 61.200 265.000 ;
        RECT 62.000 262.200 62.800 265.000 ;
        RECT 63.600 262.200 64.400 265.400 ;
        RECT 70.000 262.200 70.800 268.200 ;
        RECT 73.200 267.600 74.000 268.400 ;
        RECT 74.800 268.300 75.600 268.400 ;
        RECT 78.200 268.300 78.800 269.800 ;
        RECT 81.200 269.600 82.000 269.800 ;
        RECT 74.800 267.700 78.800 268.300 ;
        RECT 74.800 267.600 75.600 267.700 ;
        RECT 71.600 264.800 72.400 266.400 ;
        RECT 73.400 266.300 74.000 267.600 ;
        RECT 76.400 266.300 77.200 266.400 ;
        RECT 73.300 265.700 77.200 266.300 ;
        RECT 78.200 266.200 78.800 267.700 ;
        RECT 79.600 267.600 80.400 269.200 ;
        RECT 73.400 264.200 74.000 265.700 ;
        RECT 76.400 265.600 77.200 265.700 ;
        RECT 76.600 264.800 77.400 265.600 ;
        RECT 73.200 262.200 74.000 264.200 ;
        RECT 78.000 262.200 78.800 266.200 ;
        RECT 84.200 266.800 85.000 271.200 ;
        RECT 85.800 270.600 86.400 272.400 ;
        RECT 85.600 270.000 86.400 270.600 ;
        RECT 92.400 270.000 115.800 270.600 ;
        RECT 85.600 268.000 86.200 270.000 ;
        RECT 92.400 269.400 93.200 270.000 ;
        RECT 110.000 269.600 110.800 270.000 ;
        RECT 113.200 269.600 114.000 270.000 ;
        RECT 115.000 269.800 115.800 270.000 ;
        RECT 86.800 268.600 90.600 269.400 ;
        RECT 85.600 267.400 86.800 268.000 ;
        RECT 84.200 266.000 85.200 266.800 ;
        RECT 84.400 262.200 85.200 266.000 ;
        RECT 86.000 262.200 86.800 267.400 ;
        RECT 89.800 267.400 90.600 268.600 ;
        RECT 89.800 266.800 91.600 267.400 ;
        RECT 90.800 266.200 91.600 266.800 ;
        RECT 95.600 266.400 96.400 269.200 ;
        RECT 98.800 268.600 102.000 269.400 ;
        RECT 105.800 268.600 107.800 269.400 ;
        RECT 116.400 269.000 117.200 274.600 ;
        RECT 118.000 271.800 118.800 279.800 ;
        RECT 119.600 272.400 120.400 279.800 ;
        RECT 122.800 272.400 123.600 279.800 ;
        RECT 119.600 271.800 123.600 272.400 ;
        RECT 118.200 270.400 118.800 271.800 ;
        RECT 126.000 271.200 126.800 279.800 ;
        RECT 129.200 271.200 130.000 279.800 ;
        RECT 132.400 271.200 133.200 279.800 ;
        RECT 135.600 271.200 136.400 279.800 ;
        RECT 122.000 270.400 122.800 270.800 ;
        RECT 124.400 270.400 126.800 271.200 ;
        RECT 127.800 270.400 130.000 271.200 ;
        RECT 131.000 270.400 133.200 271.200 ;
        RECT 134.600 270.400 136.400 271.200 ;
        RECT 140.400 271.200 141.200 279.800 ;
        RECT 143.600 271.200 144.400 279.800 ;
        RECT 146.800 271.200 147.600 279.800 ;
        RECT 150.000 271.200 150.800 279.800 ;
        RECT 158.000 272.400 158.800 279.800 ;
        RECT 161.200 272.800 162.000 279.800 ;
        RECT 165.000 278.400 165.800 279.800 ;
        RECT 164.400 277.600 165.800 278.400 ;
        RECT 158.000 271.800 160.600 272.400 ;
        RECT 161.200 271.800 162.200 272.800 ;
        RECT 165.000 272.600 165.800 277.600 ;
        RECT 165.000 271.800 166.800 272.600 ;
        RECT 169.800 272.400 170.600 279.800 ;
        RECT 169.200 271.800 170.600 272.400 ;
        RECT 140.400 270.400 142.200 271.200 ;
        RECT 143.600 270.400 145.800 271.200 ;
        RECT 146.800 270.400 149.000 271.200 ;
        RECT 150.000 270.400 152.400 271.200 ;
        RECT 118.000 269.800 120.400 270.400 ;
        RECT 122.000 269.800 123.600 270.400 ;
        RECT 118.000 269.600 118.800 269.800 ;
        RECT 98.400 267.800 99.200 268.000 ;
        RECT 98.400 267.200 102.800 267.800 ;
        RECT 102.000 267.000 102.800 267.200 ;
        RECT 103.600 266.800 104.400 268.400 ;
        RECT 90.800 265.400 93.200 266.200 ;
        RECT 95.600 265.600 96.600 266.400 ;
        RECT 99.600 265.600 101.200 266.400 ;
        RECT 102.000 266.200 102.800 266.400 ;
        RECT 105.800 266.200 106.600 268.600 ;
        RECT 108.400 268.200 117.200 269.000 ;
        RECT 111.800 266.800 114.800 267.600 ;
        RECT 111.800 266.200 112.600 266.800 ;
        RECT 102.000 265.600 106.600 266.200 ;
        RECT 92.400 262.200 93.200 265.400 ;
        RECT 110.000 265.400 112.600 266.200 ;
        RECT 94.000 262.200 94.800 265.000 ;
        RECT 95.600 262.200 96.400 265.000 ;
        RECT 97.200 262.200 98.000 265.000 ;
        RECT 98.800 262.200 99.600 265.000 ;
        RECT 102.000 262.200 102.800 265.000 ;
        RECT 105.200 262.200 106.000 265.000 ;
        RECT 106.800 262.200 107.600 265.000 ;
        RECT 108.400 262.200 109.200 265.000 ;
        RECT 110.000 262.200 110.800 265.400 ;
        RECT 116.400 262.200 117.200 268.200 ;
        RECT 118.000 265.600 118.800 266.400 ;
        RECT 119.800 266.200 120.400 269.800 ;
        RECT 122.800 269.600 123.600 269.800 ;
        RECT 121.200 267.600 122.000 269.200 ;
        RECT 124.400 267.600 125.200 270.400 ;
        RECT 127.800 269.000 128.600 270.400 ;
        RECT 131.000 269.000 131.800 270.400 ;
        RECT 134.600 269.000 135.400 270.400 ;
        RECT 141.400 269.000 142.200 270.400 ;
        RECT 145.000 269.000 145.800 270.400 ;
        RECT 148.200 269.000 149.000 270.400 ;
        RECT 126.000 268.200 128.600 269.000 ;
        RECT 129.400 268.200 131.800 269.000 ;
        RECT 132.800 268.200 135.400 269.000 ;
        RECT 136.200 268.300 138.000 269.000 ;
        RECT 138.800 268.300 140.600 269.000 ;
        RECT 136.200 268.200 140.600 268.300 ;
        RECT 141.400 268.200 144.000 269.000 ;
        RECT 145.000 268.200 147.400 269.000 ;
        RECT 148.200 268.200 150.800 269.000 ;
        RECT 127.800 267.600 128.600 268.200 ;
        RECT 131.000 267.600 131.800 268.200 ;
        RECT 134.600 267.600 135.400 268.200 ;
        RECT 137.200 267.700 139.600 268.200 ;
        RECT 137.200 267.600 138.000 267.700 ;
        RECT 138.800 267.600 139.600 267.700 ;
        RECT 141.400 267.600 142.200 268.200 ;
        RECT 145.000 267.600 145.800 268.200 ;
        RECT 148.200 267.600 149.000 268.200 ;
        RECT 151.600 267.600 152.400 270.400 ;
        RECT 153.200 270.300 154.000 270.400 ;
        RECT 158.000 270.300 159.000 270.400 ;
        RECT 153.200 269.700 159.000 270.300 ;
        RECT 153.200 269.600 154.000 269.700 ;
        RECT 158.000 269.600 159.000 269.700 ;
        RECT 158.200 268.800 159.000 269.600 ;
        RECT 160.000 269.800 160.600 271.800 ;
        RECT 160.000 269.000 161.000 269.800 ;
        RECT 124.400 266.800 126.800 267.600 ;
        RECT 127.800 266.800 130.000 267.600 ;
        RECT 131.000 266.800 133.200 267.600 ;
        RECT 134.600 266.800 136.400 267.600 ;
        RECT 118.200 264.800 119.000 265.600 ;
        RECT 119.600 262.200 120.400 266.200 ;
        RECT 126.000 262.200 126.800 266.800 ;
        RECT 129.200 262.200 130.000 266.800 ;
        RECT 132.400 262.200 133.200 266.800 ;
        RECT 135.600 262.200 136.400 266.800 ;
        RECT 140.400 266.800 142.200 267.600 ;
        RECT 143.600 266.800 145.800 267.600 ;
        RECT 146.800 266.800 149.000 267.600 ;
        RECT 150.000 266.800 152.400 267.600 ;
        RECT 160.000 267.400 160.600 269.000 ;
        RECT 161.600 268.400 162.200 271.800 ;
        RECT 164.400 269.600 165.200 271.200 ;
        RECT 166.000 268.400 166.600 271.800 ;
        RECT 169.200 271.600 170.000 271.800 ;
        RECT 169.200 270.400 169.800 271.600 ;
        RECT 174.000 271.200 174.800 279.800 ;
        RECT 177.200 276.400 178.000 279.800 ;
        RECT 177.000 275.800 178.000 276.400 ;
        RECT 177.000 275.200 177.600 275.800 ;
        RECT 180.400 275.200 181.200 279.800 ;
        RECT 183.600 277.000 184.400 279.800 ;
        RECT 185.200 277.000 186.000 279.800 ;
        RECT 170.800 270.800 174.800 271.200 ;
        RECT 170.600 270.600 174.800 270.800 ;
        RECT 175.600 274.600 177.600 275.200 ;
        RECT 169.200 269.600 170.000 270.400 ;
        RECT 170.600 270.000 171.400 270.600 ;
        RECT 161.200 268.300 162.200 268.400 ;
        RECT 162.800 268.300 163.600 268.400 ;
        RECT 161.200 267.700 163.600 268.300 ;
        RECT 161.200 267.600 162.200 267.700 ;
        RECT 162.800 267.600 163.600 267.700 ;
        RECT 166.000 267.600 166.800 268.400 ;
        RECT 158.000 266.800 160.600 267.400 ;
        RECT 140.400 262.200 141.200 266.800 ;
        RECT 143.600 262.200 144.400 266.800 ;
        RECT 146.800 262.200 147.600 266.800 ;
        RECT 150.000 262.200 150.800 266.800 ;
        RECT 158.000 262.200 158.800 266.800 ;
        RECT 161.600 266.200 162.200 267.600 ;
        RECT 161.200 265.600 162.200 266.200 ;
        RECT 161.200 262.200 162.000 265.600 ;
        RECT 166.000 264.200 166.600 267.600 ;
        RECT 167.600 264.800 168.400 266.400 ;
        RECT 169.200 266.200 169.800 269.600 ;
        RECT 170.600 267.000 171.200 270.000 ;
        RECT 175.600 269.000 176.400 274.600 ;
        RECT 178.200 274.400 182.400 275.200 ;
        RECT 186.800 275.000 187.600 279.800 ;
        RECT 190.000 275.000 190.800 279.800 ;
        RECT 178.200 274.000 178.800 274.400 ;
        RECT 177.200 273.200 178.800 274.000 ;
        RECT 181.800 273.800 187.600 274.400 ;
        RECT 179.800 273.200 181.200 273.800 ;
        RECT 179.800 273.000 186.000 273.200 ;
        RECT 180.600 272.600 186.000 273.000 ;
        RECT 185.200 272.400 186.000 272.600 ;
        RECT 187.000 273.000 187.600 273.800 ;
        RECT 188.200 273.600 190.800 274.400 ;
        RECT 193.200 273.600 194.000 279.800 ;
        RECT 194.800 277.000 195.600 279.800 ;
        RECT 196.400 277.000 197.200 279.800 ;
        RECT 198.000 277.000 198.800 279.800 ;
        RECT 196.400 274.400 200.600 275.200 ;
        RECT 201.200 274.400 202.000 279.800 ;
        RECT 204.400 275.200 205.200 279.800 ;
        RECT 204.400 274.600 207.000 275.200 ;
        RECT 201.200 273.600 203.800 274.400 ;
        RECT 194.800 273.000 195.600 273.200 ;
        RECT 187.000 272.400 195.600 273.000 ;
        RECT 198.000 273.000 198.800 273.200 ;
        RECT 206.400 273.000 207.000 274.600 ;
        RECT 198.000 272.400 207.000 273.000 ;
        RECT 206.400 270.600 207.000 272.400 ;
        RECT 207.600 272.000 208.400 279.800 ;
        RECT 207.600 271.200 208.600 272.000 ;
        RECT 177.000 270.000 200.400 270.600 ;
        RECT 206.400 270.000 207.200 270.600 ;
        RECT 177.000 269.800 177.800 270.000 ;
        RECT 178.800 269.600 179.600 270.000 ;
        RECT 182.000 269.600 182.800 270.000 ;
        RECT 199.600 269.400 200.400 270.000 ;
        RECT 175.600 268.200 184.400 269.000 ;
        RECT 185.000 268.600 187.000 269.400 ;
        RECT 190.800 268.600 194.000 269.400 ;
        RECT 170.600 266.400 173.000 267.000 ;
        RECT 166.000 262.200 166.800 264.200 ;
        RECT 169.200 262.200 170.000 266.200 ;
        RECT 172.400 264.200 173.000 266.400 ;
        RECT 174.000 264.800 174.800 266.400 ;
        RECT 172.400 262.200 173.200 264.200 ;
        RECT 175.600 262.200 176.400 268.200 ;
        RECT 178.000 266.800 181.000 267.600 ;
        RECT 180.200 266.200 181.000 266.800 ;
        RECT 186.200 266.200 187.000 268.600 ;
        RECT 188.400 266.800 189.200 268.400 ;
        RECT 193.600 267.800 194.400 268.000 ;
        RECT 190.000 267.200 194.400 267.800 ;
        RECT 190.000 267.000 190.800 267.200 ;
        RECT 196.400 266.400 197.200 269.200 ;
        RECT 202.200 268.600 206.000 269.400 ;
        RECT 202.200 267.400 203.000 268.600 ;
        RECT 206.600 268.000 207.200 270.000 ;
        RECT 190.000 266.200 190.800 266.400 ;
        RECT 180.200 265.400 182.800 266.200 ;
        RECT 186.200 265.600 190.800 266.200 ;
        RECT 191.600 265.600 193.200 266.400 ;
        RECT 196.200 265.600 197.200 266.400 ;
        RECT 201.200 266.800 203.000 267.400 ;
        RECT 206.000 267.400 207.200 268.000 ;
        RECT 201.200 266.200 202.000 266.800 ;
        RECT 182.000 262.200 182.800 265.400 ;
        RECT 199.600 265.400 202.000 266.200 ;
        RECT 183.600 262.200 184.400 265.000 ;
        RECT 185.200 262.200 186.000 265.000 ;
        RECT 186.800 262.200 187.600 265.000 ;
        RECT 190.000 262.200 190.800 265.000 ;
        RECT 193.200 262.200 194.000 265.000 ;
        RECT 194.800 262.200 195.600 265.000 ;
        RECT 196.400 262.200 197.200 265.000 ;
        RECT 198.000 262.200 198.800 265.000 ;
        RECT 199.600 262.200 200.400 265.400 ;
        RECT 206.000 262.200 206.800 267.400 ;
        RECT 207.800 266.800 208.600 271.200 ;
        RECT 207.600 266.000 208.600 266.800 ;
        RECT 210.800 270.300 211.600 279.800 ;
        RECT 212.400 270.300 213.200 270.400 ;
        RECT 210.800 269.700 213.200 270.300 ;
        RECT 207.600 262.200 208.400 266.000 ;
        RECT 210.800 262.200 211.600 269.700 ;
        RECT 212.400 269.600 213.200 269.700 ;
        RECT 212.400 268.300 213.200 268.400 ;
        RECT 214.000 268.300 214.800 268.400 ;
        RECT 212.400 267.700 214.800 268.300 ;
        RECT 212.400 266.800 213.200 267.700 ;
        RECT 214.000 266.800 214.800 267.700 ;
        RECT 215.600 268.300 216.400 279.800 ;
        RECT 217.200 271.600 218.000 273.200 ;
        RECT 218.800 268.300 219.600 268.400 ;
        RECT 215.600 267.700 219.600 268.300 ;
        RECT 215.600 266.200 216.400 267.700 ;
        RECT 218.800 266.800 219.600 267.700 ;
        RECT 220.400 266.200 221.200 279.800 ;
        RECT 222.000 271.600 222.800 273.200 ;
        RECT 225.200 271.200 226.000 279.800 ;
        RECT 228.400 271.200 229.200 279.800 ;
        RECT 233.200 276.400 234.000 279.800 ;
        RECT 233.000 275.800 234.000 276.400 ;
        RECT 233.000 275.200 233.600 275.800 ;
        RECT 236.400 275.200 237.200 279.800 ;
        RECT 239.600 277.000 240.400 279.800 ;
        RECT 241.200 277.000 242.000 279.800 ;
        RECT 225.200 270.400 229.200 271.200 ;
        RECT 231.600 274.600 233.600 275.200 ;
        RECT 225.200 267.600 226.000 270.400 ;
        RECT 231.600 269.000 232.400 274.600 ;
        RECT 234.200 274.400 238.400 275.200 ;
        RECT 242.800 275.000 243.600 279.800 ;
        RECT 246.000 275.000 246.800 279.800 ;
        RECT 234.200 274.000 234.800 274.400 ;
        RECT 233.200 273.200 234.800 274.000 ;
        RECT 237.800 273.800 243.600 274.400 ;
        RECT 235.800 273.200 237.200 273.800 ;
        RECT 235.800 273.000 242.000 273.200 ;
        RECT 236.600 272.600 242.000 273.000 ;
        RECT 241.200 272.400 242.000 272.600 ;
        RECT 243.000 273.000 243.600 273.800 ;
        RECT 244.200 273.600 246.800 274.400 ;
        RECT 249.200 273.600 250.000 279.800 ;
        RECT 250.800 277.000 251.600 279.800 ;
        RECT 252.400 277.000 253.200 279.800 ;
        RECT 254.000 277.000 254.800 279.800 ;
        RECT 252.400 274.400 256.600 275.200 ;
        RECT 257.200 274.400 258.000 279.800 ;
        RECT 260.400 275.200 261.200 279.800 ;
        RECT 260.400 274.600 263.000 275.200 ;
        RECT 257.200 273.600 259.800 274.400 ;
        RECT 250.800 273.000 251.600 273.200 ;
        RECT 243.000 272.400 251.600 273.000 ;
        RECT 254.000 273.000 254.800 273.200 ;
        RECT 262.400 273.000 263.000 274.600 ;
        RECT 254.000 272.400 263.000 273.000 ;
        RECT 262.400 270.600 263.000 272.400 ;
        RECT 263.600 272.000 264.400 279.800 ;
        RECT 266.800 275.000 267.600 279.000 ;
        RECT 263.600 271.200 264.600 272.000 ;
        RECT 233.000 270.000 256.400 270.600 ;
        RECT 262.400 270.000 263.200 270.600 ;
        RECT 233.000 269.800 233.800 270.000 ;
        RECT 238.000 269.600 238.800 270.000 ;
        RECT 255.600 269.400 256.400 270.000 ;
        RECT 231.600 268.200 240.400 269.000 ;
        RECT 241.000 268.600 243.000 269.400 ;
        RECT 246.800 268.600 250.000 269.400 ;
        RECT 225.200 266.800 229.200 267.600 ;
        RECT 215.600 265.600 217.400 266.200 ;
        RECT 220.400 265.600 222.200 266.200 ;
        RECT 216.600 262.200 217.400 265.600 ;
        RECT 221.400 262.200 222.200 265.600 ;
        RECT 225.200 262.200 226.000 266.800 ;
        RECT 228.400 262.200 229.200 266.800 ;
        RECT 231.600 262.200 232.400 268.200 ;
        RECT 234.000 266.800 237.000 267.600 ;
        RECT 236.200 266.200 237.000 266.800 ;
        RECT 242.200 266.200 243.000 268.600 ;
        RECT 244.400 266.800 245.200 268.400 ;
        RECT 249.600 267.800 250.400 268.000 ;
        RECT 246.000 267.200 250.400 267.800 ;
        RECT 246.000 267.000 246.800 267.200 ;
        RECT 252.400 266.400 253.200 269.200 ;
        RECT 258.200 268.600 262.000 269.400 ;
        RECT 258.200 267.400 259.000 268.600 ;
        RECT 262.600 268.000 263.200 270.000 ;
        RECT 246.000 266.200 246.800 266.400 ;
        RECT 236.200 265.400 238.800 266.200 ;
        RECT 242.200 265.600 246.800 266.200 ;
        RECT 247.600 265.600 249.200 266.400 ;
        RECT 252.200 265.600 253.200 266.400 ;
        RECT 257.200 266.800 259.000 267.400 ;
        RECT 262.000 267.400 263.200 268.000 ;
        RECT 257.200 266.200 258.000 266.800 ;
        RECT 238.000 262.200 238.800 265.400 ;
        RECT 255.600 265.400 258.000 266.200 ;
        RECT 239.600 262.200 240.400 265.000 ;
        RECT 241.200 262.200 242.000 265.000 ;
        RECT 242.800 262.200 243.600 265.000 ;
        RECT 246.000 262.200 246.800 265.000 ;
        RECT 249.200 262.200 250.000 265.000 ;
        RECT 250.800 262.200 251.600 265.000 ;
        RECT 252.400 262.200 253.200 265.000 ;
        RECT 254.000 262.200 254.800 265.000 ;
        RECT 255.600 262.200 256.400 265.400 ;
        RECT 262.000 262.200 262.800 267.400 ;
        RECT 263.800 266.800 264.600 271.200 ;
        RECT 266.800 271.600 267.400 275.000 ;
        RECT 271.000 272.800 271.800 279.800 ;
        RECT 271.000 272.200 272.600 272.800 ;
        RECT 266.800 271.000 270.600 271.600 ;
        RECT 266.800 268.800 267.600 270.400 ;
        RECT 268.400 268.800 269.200 270.400 ;
        RECT 270.000 269.000 270.600 271.000 ;
        RECT 270.000 268.200 271.400 269.000 ;
        RECT 272.000 268.400 272.600 272.200 ;
        RECT 273.200 270.300 274.000 271.200 ;
        RECT 276.400 270.300 277.200 279.800 ;
        RECT 280.400 273.600 281.200 274.400 ;
        RECT 280.400 272.400 281.000 273.600 ;
        RECT 281.800 272.400 282.600 279.800 ;
        RECT 288.600 272.400 289.400 279.800 ;
        RECT 290.000 273.600 290.800 274.400 ;
        RECT 290.200 272.400 290.800 273.600 ;
        RECT 279.600 271.800 281.000 272.400 ;
        RECT 281.600 271.800 282.600 272.400 ;
        RECT 279.600 271.600 280.400 271.800 ;
        RECT 273.200 269.700 277.200 270.300 ;
        RECT 273.200 269.600 274.000 269.700 ;
        RECT 270.000 267.800 271.000 268.200 ;
        RECT 263.600 266.000 264.600 266.800 ;
        RECT 266.800 267.200 271.000 267.800 ;
        RECT 272.000 267.600 274.000 268.400 ;
        RECT 263.600 262.200 264.400 266.000 ;
        RECT 266.800 265.000 267.400 267.200 ;
        RECT 272.000 267.000 272.600 267.600 ;
        RECT 271.800 266.600 272.600 267.000 ;
        RECT 271.000 266.400 272.600 266.600 ;
        RECT 270.000 266.000 272.600 266.400 ;
        RECT 270.000 265.600 271.800 266.000 ;
        RECT 266.800 263.000 267.600 265.000 ;
        RECT 271.000 263.000 271.800 265.600 ;
        RECT 276.400 262.200 277.200 269.700 ;
        RECT 278.000 270.300 278.800 270.400 ;
        RECT 281.600 270.300 282.200 271.800 ;
        RECT 287.600 271.600 289.600 272.400 ;
        RECT 290.200 271.800 291.600 272.400 ;
        RECT 290.800 271.600 291.600 271.800 ;
        RECT 278.000 269.700 282.200 270.300 ;
        RECT 278.000 269.600 278.800 269.700 ;
        RECT 281.600 268.400 282.200 269.700 ;
        RECT 282.800 270.300 283.600 270.400 ;
        RECT 286.000 270.300 286.800 270.400 ;
        RECT 282.800 269.700 286.800 270.300 ;
        RECT 282.800 268.800 283.600 269.700 ;
        RECT 286.000 269.600 286.800 269.700 ;
        RECT 287.600 268.800 288.400 270.400 ;
        RECT 289.000 268.400 289.600 271.600 ;
        RECT 279.600 267.600 282.200 268.400 ;
        RECT 284.400 268.200 285.200 268.400 ;
        RECT 283.600 267.600 285.200 268.200 ;
        RECT 286.000 268.200 286.800 268.400 ;
        RECT 286.000 267.600 287.600 268.200 ;
        RECT 289.000 267.600 291.600 268.400 ;
        RECT 278.000 264.800 278.800 266.400 ;
        RECT 279.800 266.200 280.400 267.600 ;
        RECT 283.600 267.200 284.400 267.600 ;
        RECT 286.800 267.200 287.600 267.600 ;
        RECT 281.400 266.200 285.000 266.600 ;
        RECT 286.200 266.200 289.800 266.600 ;
        RECT 290.800 266.200 291.400 267.600 ;
        RECT 279.600 262.200 280.400 266.200 ;
        RECT 281.200 266.000 285.200 266.200 ;
        RECT 281.200 262.200 282.000 266.000 ;
        RECT 284.400 262.200 285.200 266.000 ;
        RECT 286.000 266.000 290.000 266.200 ;
        RECT 286.000 262.200 286.800 266.000 ;
        RECT 289.200 262.200 290.000 266.000 ;
        RECT 290.800 262.200 291.600 266.200 ;
        RECT 292.400 264.800 293.200 266.400 ;
        RECT 294.000 262.200 294.800 279.800 ;
        RECT 295.600 275.000 296.400 279.000 ;
        RECT 295.600 271.600 296.200 275.000 ;
        RECT 299.800 272.800 300.600 279.800 ;
        RECT 311.600 276.400 312.400 279.800 ;
        RECT 311.400 275.800 312.400 276.400 ;
        RECT 311.400 275.200 312.000 275.800 ;
        RECT 314.800 275.200 315.600 279.800 ;
        RECT 318.000 277.000 318.800 279.800 ;
        RECT 319.600 277.000 320.400 279.800 ;
        RECT 310.000 274.600 312.000 275.200 ;
        RECT 299.800 272.200 301.400 272.800 ;
        RECT 295.600 271.000 299.400 271.600 ;
        RECT 295.600 268.800 296.400 270.400 ;
        RECT 297.200 268.800 298.000 270.400 ;
        RECT 298.800 269.000 299.400 271.000 ;
        RECT 298.800 268.200 300.200 269.000 ;
        RECT 300.800 268.400 301.400 272.200 ;
        RECT 302.000 269.600 302.800 271.200 ;
        RECT 310.000 269.000 310.800 274.600 ;
        RECT 312.600 274.400 316.800 275.200 ;
        RECT 321.200 275.000 322.000 279.800 ;
        RECT 324.400 275.000 325.200 279.800 ;
        RECT 312.600 274.000 313.200 274.400 ;
        RECT 311.600 273.200 313.200 274.000 ;
        RECT 316.200 273.800 322.000 274.400 ;
        RECT 314.200 273.200 315.600 273.800 ;
        RECT 314.200 273.000 320.400 273.200 ;
        RECT 315.000 272.600 320.400 273.000 ;
        RECT 319.600 272.400 320.400 272.600 ;
        RECT 321.400 273.000 322.000 273.800 ;
        RECT 322.600 273.600 325.200 274.400 ;
        RECT 327.600 273.600 328.400 279.800 ;
        RECT 329.200 277.000 330.000 279.800 ;
        RECT 330.800 277.000 331.600 279.800 ;
        RECT 332.400 277.000 333.200 279.800 ;
        RECT 330.800 274.400 335.000 275.200 ;
        RECT 335.600 274.400 336.400 279.800 ;
        RECT 338.800 275.200 339.600 279.800 ;
        RECT 338.800 274.600 341.400 275.200 ;
        RECT 335.600 273.600 338.200 274.400 ;
        RECT 329.200 273.000 330.000 273.200 ;
        RECT 321.400 272.400 330.000 273.000 ;
        RECT 332.400 273.000 333.200 273.200 ;
        RECT 340.800 273.000 341.400 274.600 ;
        RECT 332.400 272.400 341.400 273.000 ;
        RECT 340.800 270.600 341.400 272.400 ;
        RECT 342.000 272.000 342.800 279.800 ;
        RECT 343.600 274.300 344.400 274.400 ;
        RECT 345.200 274.300 346.000 279.800 ;
        RECT 343.600 273.700 346.000 274.300 ;
        RECT 343.600 273.600 344.400 273.700 ;
        RECT 342.000 271.200 343.000 272.000 ;
        RECT 311.400 270.000 334.800 270.600 ;
        RECT 340.800 270.000 341.600 270.600 ;
        RECT 311.400 269.800 312.200 270.000 ;
        RECT 316.400 269.600 317.200 270.000 ;
        RECT 322.800 269.600 323.600 270.000 ;
        RECT 334.000 269.400 334.800 270.000 ;
        RECT 300.800 268.300 302.800 268.400 ;
        RECT 308.400 268.300 309.200 268.400 ;
        RECT 298.800 267.800 299.800 268.200 ;
        RECT 295.600 267.200 299.800 267.800 ;
        RECT 300.800 267.700 309.200 268.300 ;
        RECT 300.800 267.600 302.800 267.700 ;
        RECT 308.400 267.600 309.200 267.700 ;
        RECT 310.000 268.200 318.800 269.000 ;
        RECT 319.400 268.600 321.400 269.400 ;
        RECT 325.200 268.600 328.400 269.400 ;
        RECT 295.600 265.000 296.200 267.200 ;
        RECT 300.800 267.000 301.400 267.600 ;
        RECT 300.600 266.600 301.400 267.000 ;
        RECT 299.800 266.000 301.400 266.600 ;
        RECT 295.600 263.000 296.400 265.000 ;
        RECT 299.800 263.000 300.600 266.000 ;
        RECT 310.000 262.200 310.800 268.200 ;
        RECT 312.400 266.800 315.400 267.600 ;
        RECT 314.600 266.200 315.400 266.800 ;
        RECT 320.600 266.200 321.400 268.600 ;
        RECT 322.800 266.800 323.600 268.400 ;
        RECT 328.000 267.800 328.800 268.000 ;
        RECT 324.400 267.200 328.800 267.800 ;
        RECT 324.400 267.000 325.200 267.200 ;
        RECT 330.800 266.400 331.600 269.200 ;
        RECT 336.600 268.600 340.400 269.400 ;
        RECT 336.600 267.400 337.400 268.600 ;
        RECT 341.000 268.000 341.600 270.000 ;
        RECT 324.400 266.200 325.200 266.400 ;
        RECT 314.600 265.400 317.200 266.200 ;
        RECT 320.600 265.600 325.200 266.200 ;
        RECT 326.000 265.600 327.600 266.400 ;
        RECT 330.600 265.600 331.600 266.400 ;
        RECT 335.600 266.800 337.400 267.400 ;
        RECT 340.400 267.400 341.600 268.000 ;
        RECT 335.600 266.200 336.400 266.800 ;
        RECT 316.400 262.200 317.200 265.400 ;
        RECT 334.000 265.400 336.400 266.200 ;
        RECT 318.000 262.200 318.800 265.000 ;
        RECT 319.600 262.200 320.400 265.000 ;
        RECT 321.200 262.200 322.000 265.000 ;
        RECT 324.400 262.200 325.200 265.000 ;
        RECT 327.600 262.200 328.400 265.000 ;
        RECT 329.200 262.200 330.000 265.000 ;
        RECT 330.800 262.200 331.600 265.000 ;
        RECT 332.400 262.200 333.200 265.000 ;
        RECT 334.000 262.200 334.800 265.400 ;
        RECT 340.400 262.200 341.200 267.400 ;
        RECT 342.200 266.800 343.000 271.200 ;
        RECT 342.000 266.000 343.000 266.800 ;
        RECT 342.000 262.200 342.800 266.000 ;
        RECT 345.200 262.200 346.000 273.700 ;
        RECT 349.200 273.600 350.000 274.400 ;
        RECT 349.200 272.400 349.800 273.600 ;
        RECT 350.600 272.400 351.400 279.800 ;
        RECT 357.400 272.400 358.200 279.800 ;
        RECT 358.800 273.600 359.600 274.400 ;
        RECT 359.000 272.400 359.600 273.600 ;
        RECT 346.800 272.300 347.600 272.400 ;
        RECT 348.400 272.300 349.800 272.400 ;
        RECT 346.800 271.800 349.800 272.300 ;
        RECT 350.400 271.800 351.400 272.400 ;
        RECT 346.800 271.700 349.200 271.800 ;
        RECT 346.800 271.600 347.600 271.700 ;
        RECT 348.400 271.600 349.200 271.700 ;
        RECT 348.400 270.300 349.200 270.400 ;
        RECT 350.400 270.300 351.000 271.800 ;
        RECT 356.400 271.600 358.400 272.400 ;
        RECT 359.000 271.800 360.400 272.400 ;
        RECT 359.600 271.600 360.400 271.800 ;
        RECT 348.400 269.700 351.000 270.300 ;
        RECT 348.400 269.600 349.200 269.700 ;
        RECT 350.400 268.400 351.000 269.700 ;
        RECT 351.600 268.800 352.400 270.400 ;
        RECT 353.200 270.300 354.000 270.400 ;
        RECT 356.400 270.300 357.200 270.400 ;
        RECT 353.200 269.700 357.200 270.300 ;
        RECT 353.200 269.600 354.000 269.700 ;
        RECT 356.400 268.800 357.200 269.700 ;
        RECT 357.800 268.400 358.400 271.600 ;
        RECT 359.600 270.300 360.400 270.400 ;
        RECT 361.200 270.300 362.000 279.800 ;
        RECT 364.400 271.600 365.200 273.200 ;
        RECT 359.600 269.700 362.000 270.300 ;
        RECT 359.600 269.600 360.400 269.700 ;
        RECT 348.400 267.600 351.000 268.400 ;
        RECT 353.200 268.200 354.000 268.400 ;
        RECT 352.400 267.600 354.000 268.200 ;
        RECT 354.800 268.200 355.600 268.400 ;
        RECT 354.800 267.600 356.400 268.200 ;
        RECT 357.800 267.600 360.400 268.400 ;
        RECT 346.800 264.800 347.600 266.400 ;
        RECT 348.600 266.200 349.200 267.600 ;
        RECT 352.400 267.200 353.200 267.600 ;
        RECT 355.600 267.200 356.400 267.600 ;
        RECT 350.200 266.200 353.800 266.600 ;
        RECT 355.000 266.200 358.600 266.600 ;
        RECT 359.600 266.200 360.200 267.600 ;
        RECT 348.400 262.200 349.200 266.200 ;
        RECT 350.000 266.000 354.000 266.200 ;
        RECT 350.000 262.200 350.800 266.000 ;
        RECT 353.200 262.200 354.000 266.000 ;
        RECT 354.800 266.000 358.800 266.200 ;
        RECT 354.800 262.200 355.600 266.000 ;
        RECT 358.000 262.200 358.800 266.000 ;
        RECT 359.600 262.200 360.400 266.200 ;
        RECT 361.200 262.200 362.000 269.700 ;
        RECT 362.800 264.800 363.600 266.400 ;
        RECT 366.000 266.200 366.800 279.800 ;
        RECT 370.800 275.800 371.600 279.800 ;
        RECT 371.000 275.600 371.600 275.800 ;
        RECT 374.000 275.800 374.800 279.800 ;
        RECT 377.200 275.800 378.000 279.800 ;
        RECT 374.000 275.600 374.600 275.800 ;
        RECT 371.000 275.000 374.600 275.600 ;
        RECT 377.400 275.600 378.000 275.800 ;
        RECT 380.400 275.800 381.200 279.800 ;
        RECT 383.600 275.800 384.400 279.800 ;
        RECT 380.400 275.600 381.000 275.800 ;
        RECT 377.400 275.000 381.000 275.600 ;
        RECT 383.800 275.600 384.400 275.800 ;
        RECT 386.800 275.800 387.600 279.800 ;
        RECT 390.000 275.800 390.800 279.800 ;
        RECT 386.800 275.600 387.400 275.800 ;
        RECT 383.800 275.000 387.400 275.600 ;
        RECT 390.200 275.600 390.800 275.800 ;
        RECT 393.200 275.800 394.000 279.800 ;
        RECT 393.200 275.600 393.800 275.800 ;
        RECT 390.200 275.000 393.800 275.600 ;
        RECT 372.400 272.800 373.200 274.400 ;
        RECT 374.000 272.400 374.600 275.000 ;
        RECT 378.800 272.800 379.600 274.400 ;
        RECT 380.400 272.400 381.000 275.000 ;
        RECT 385.200 272.800 386.000 274.400 ;
        RECT 386.800 272.400 387.400 275.000 ;
        RECT 391.600 272.800 392.400 274.400 ;
        RECT 393.200 272.400 393.800 275.000 ;
        RECT 394.800 272.400 395.600 279.800 ;
        RECT 398.000 279.200 402.000 279.800 ;
        RECT 398.000 272.400 398.800 279.200 ;
        RECT 369.200 270.800 370.000 272.400 ;
        RECT 374.000 271.600 374.800 272.400 ;
        RECT 374.000 268.400 374.600 271.600 ;
        RECT 375.600 270.800 376.400 272.400 ;
        RECT 380.400 271.600 381.200 272.400 ;
        RECT 377.200 269.600 378.800 270.400 ;
        RECT 380.400 268.400 381.000 271.600 ;
        RECT 382.000 270.800 382.800 272.400 ;
        RECT 386.800 271.600 387.600 272.400 ;
        RECT 393.200 271.600 394.000 272.400 ;
        RECT 394.800 271.800 398.800 272.400 ;
        RECT 399.600 271.800 400.400 278.600 ;
        RECT 401.200 271.800 402.000 279.200 ;
        RECT 402.800 272.400 403.600 279.800 ;
        RECT 406.000 279.200 410.000 279.800 ;
        RECT 406.000 272.400 406.800 279.200 ;
        RECT 402.800 271.800 406.800 272.400 ;
        RECT 407.600 271.800 408.400 278.600 ;
        RECT 409.200 271.800 410.000 279.200 ;
        RECT 383.600 269.600 385.200 270.400 ;
        RECT 386.800 268.400 387.400 271.600 ;
        RECT 390.000 269.600 391.600 270.400 ;
        RECT 393.200 268.400 393.800 271.600 ;
        RECT 399.600 271.200 400.200 271.800 ;
        RECT 407.600 271.200 408.200 271.800 ;
        RECT 395.600 270.400 396.400 270.800 ;
        RECT 398.200 270.600 400.200 271.200 ;
        RECT 398.200 270.400 398.800 270.600 ;
        RECT 394.800 269.800 396.400 270.400 ;
        RECT 394.800 269.600 395.600 269.800 ;
        RECT 398.000 269.600 398.800 270.400 ;
        RECT 401.200 270.300 402.000 271.200 ;
        RECT 403.600 270.400 404.400 270.800 ;
        RECT 406.200 270.600 408.200 271.200 ;
        RECT 406.200 270.400 406.800 270.600 ;
        RECT 402.800 270.300 404.400 270.400 ;
        RECT 401.200 269.800 404.400 270.300 ;
        RECT 401.200 269.700 403.600 269.800 ;
        RECT 401.200 269.600 402.000 269.700 ;
        RECT 402.800 269.600 403.600 269.700 ;
        RECT 406.000 269.600 406.800 270.400 ;
        RECT 409.200 269.600 410.000 271.200 ;
        RECT 367.600 266.800 368.400 268.400 ;
        RECT 372.400 267.800 374.600 268.400 ;
        RECT 379.400 268.200 381.000 268.400 ;
        RECT 385.800 268.200 387.400 268.400 ;
        RECT 392.200 268.200 393.800 268.400 ;
        RECT 379.200 267.800 381.000 268.200 ;
        RECT 385.600 267.800 387.400 268.200 ;
        RECT 392.000 267.800 393.800 268.200 ;
        RECT 372.400 267.600 373.600 267.800 ;
        RECT 365.000 265.600 366.800 266.200 ;
        RECT 365.000 264.400 365.800 265.600 ;
        RECT 365.000 263.600 366.800 264.400 ;
        RECT 365.000 262.200 365.800 263.600 ;
        RECT 372.800 262.200 373.600 267.600 ;
        RECT 379.200 262.200 380.000 267.800 ;
        RECT 385.600 262.200 386.400 267.800 ;
        RECT 392.000 262.200 392.800 267.800 ;
        RECT 396.400 267.600 397.200 269.200 ;
        RECT 398.200 266.200 398.800 269.600 ;
        RECT 399.400 268.800 400.200 269.600 ;
        RECT 399.600 268.400 400.200 268.800 ;
        RECT 399.600 268.300 400.400 268.400 ;
        RECT 401.200 268.300 402.000 268.400 ;
        RECT 399.600 267.700 402.000 268.300 ;
        RECT 399.600 267.600 400.400 267.700 ;
        RECT 401.200 267.600 402.000 267.700 ;
        RECT 404.400 267.600 405.200 269.200 ;
        RECT 406.200 266.200 406.800 269.600 ;
        RECT 407.400 268.800 408.200 269.600 ;
        RECT 407.600 268.400 408.200 268.800 ;
        RECT 407.600 267.600 408.400 268.400 ;
        RECT 410.800 266.800 411.600 268.400 ;
        RECT 412.400 268.300 413.200 279.800 ;
        RECT 415.600 279.200 419.600 279.800 ;
        RECT 414.000 271.600 414.800 273.200 ;
        RECT 415.600 271.800 416.400 279.200 ;
        RECT 417.200 271.800 418.000 278.600 ;
        RECT 418.800 272.400 419.600 279.200 ;
        RECT 422.000 272.400 422.800 279.800 ;
        RECT 418.800 271.800 422.800 272.400 ;
        RECT 423.600 279.200 427.600 279.800 ;
        RECT 423.600 271.800 424.400 279.200 ;
        RECT 425.200 271.800 426.000 278.600 ;
        RECT 426.800 272.400 427.600 279.200 ;
        RECT 430.000 272.400 430.800 279.800 ;
        RECT 433.200 275.800 434.000 279.800 ;
        RECT 433.400 275.600 434.000 275.800 ;
        RECT 436.400 275.800 437.200 279.800 ;
        RECT 438.000 275.800 438.800 279.800 ;
        RECT 436.400 275.600 437.000 275.800 ;
        RECT 433.400 275.000 437.000 275.600 ;
        RECT 434.800 272.800 435.600 274.400 ;
        RECT 436.400 272.400 437.000 275.000 ;
        RECT 438.200 275.600 438.800 275.800 ;
        RECT 441.200 275.800 442.000 279.800 ;
        RECT 444.400 279.200 448.400 279.800 ;
        RECT 441.200 275.600 441.800 275.800 ;
        RECT 438.200 275.000 441.800 275.600 ;
        RECT 438.200 272.400 438.800 275.000 ;
        RECT 439.600 272.800 440.400 274.400 ;
        RECT 426.800 271.800 430.800 272.400 ;
        RECT 417.400 271.200 418.000 271.800 ;
        RECT 425.400 271.200 426.000 271.800 ;
        RECT 414.000 270.300 414.800 270.400 ;
        RECT 415.600 270.300 416.400 271.200 ;
        RECT 417.400 270.600 419.400 271.200 ;
        RECT 414.000 269.700 416.400 270.300 ;
        RECT 414.000 269.600 414.800 269.700 ;
        RECT 415.600 269.600 416.400 269.700 ;
        RECT 418.800 270.400 419.400 270.600 ;
        RECT 421.200 270.400 422.000 270.800 ;
        RECT 418.800 269.600 419.600 270.400 ;
        RECT 421.200 270.300 422.800 270.400 ;
        RECT 423.600 270.300 424.400 271.200 ;
        RECT 425.400 270.600 427.400 271.200 ;
        RECT 431.600 270.800 432.400 272.400 ;
        RECT 436.400 271.600 437.200 272.400 ;
        RECT 438.000 271.600 438.800 272.400 ;
        RECT 421.200 269.800 424.400 270.300 ;
        RECT 422.000 269.700 424.400 269.800 ;
        RECT 422.000 269.600 422.800 269.700 ;
        RECT 423.600 269.600 424.400 269.700 ;
        RECT 426.800 270.400 427.400 270.600 ;
        RECT 429.200 270.400 430.000 270.800 ;
        RECT 426.800 269.600 427.600 270.400 ;
        RECT 429.200 269.800 430.800 270.400 ;
        RECT 430.000 269.600 430.800 269.800 ;
        RECT 433.200 269.600 434.800 270.400 ;
        RECT 417.400 268.800 418.200 269.600 ;
        RECT 417.400 268.400 418.000 268.800 ;
        RECT 415.600 268.300 416.400 268.400 ;
        RECT 412.400 267.700 416.400 268.300 ;
        RECT 412.400 266.200 413.200 267.700 ;
        RECT 415.600 267.600 416.400 267.700 ;
        RECT 417.200 267.600 418.000 268.400 ;
        RECT 418.800 266.200 419.400 269.600 ;
        RECT 420.400 267.600 421.200 269.200 ;
        RECT 425.400 268.800 426.200 269.600 ;
        RECT 425.400 268.400 426.000 268.800 ;
        RECT 425.200 267.600 426.000 268.400 ;
        RECT 426.800 266.200 427.400 269.600 ;
        RECT 428.400 267.600 429.200 269.200 ;
        RECT 436.400 268.400 437.000 271.600 ;
        RECT 435.400 268.200 437.000 268.400 ;
        RECT 435.200 267.800 437.000 268.200 ;
        RECT 438.200 268.400 438.800 271.600 ;
        RECT 442.800 270.800 443.600 272.400 ;
        RECT 444.400 271.800 445.200 279.200 ;
        RECT 446.000 271.600 446.800 278.600 ;
        RECT 447.600 272.400 448.400 279.200 ;
        RECT 450.800 272.400 451.600 279.800 ;
        RECT 452.400 275.800 453.200 279.800 ;
        RECT 452.600 275.600 453.200 275.800 ;
        RECT 455.600 275.800 456.400 279.800 ;
        RECT 465.200 275.800 466.000 279.800 ;
        RECT 455.600 275.600 456.200 275.800 ;
        RECT 452.600 275.000 456.200 275.600 ;
        RECT 465.300 275.600 466.000 275.800 ;
        RECT 468.400 275.800 469.200 279.800 ;
        RECT 471.600 275.800 472.400 279.800 ;
        RECT 468.400 275.600 469.000 275.800 ;
        RECT 465.300 275.000 469.000 275.600 ;
        RECT 471.800 275.600 472.400 275.800 ;
        RECT 474.800 275.800 475.600 279.800 ;
        RECT 474.800 275.600 475.400 275.800 ;
        RECT 478.000 275.600 478.800 279.800 ;
        RECT 481.200 275.800 482.000 279.800 ;
        RECT 481.200 275.600 481.800 275.800 ;
        RECT 471.800 275.000 475.400 275.600 ;
        RECT 478.200 275.000 481.800 275.600 ;
        RECT 452.600 272.400 453.200 275.000 ;
        RECT 454.000 274.300 454.800 274.400 ;
        RECT 455.600 274.300 456.400 274.400 ;
        RECT 465.300 274.300 465.900 275.000 ;
        RECT 454.000 273.700 456.400 274.300 ;
        RECT 454.000 272.800 454.800 273.700 ;
        RECT 455.600 273.600 456.400 273.700 ;
        RECT 457.300 273.700 465.900 274.300 ;
        RECT 457.300 272.400 457.900 273.700 ;
        RECT 466.800 272.800 467.600 274.400 ;
        RECT 468.400 272.400 469.000 275.000 ;
        RECT 470.000 274.300 470.800 274.400 ;
        RECT 473.200 274.300 474.000 274.400 ;
        RECT 470.000 273.700 474.000 274.300 ;
        RECT 470.000 273.600 470.800 273.700 ;
        RECT 473.200 272.800 474.000 273.700 ;
        RECT 474.800 272.400 475.400 275.000 ;
        RECT 479.600 272.800 480.400 274.400 ;
        RECT 481.200 272.400 481.800 275.000 ;
        RECT 483.400 274.400 484.200 279.800 ;
        RECT 482.800 273.600 484.200 274.400 ;
        RECT 483.400 272.600 484.200 273.600 ;
        RECT 490.200 278.400 492.200 279.800 ;
        RECT 490.200 277.600 493.200 278.400 ;
        RECT 447.600 271.800 451.600 272.400 ;
        RECT 452.400 271.600 453.200 272.400 ;
        RECT 446.200 271.200 446.800 271.600 ;
        RECT 440.400 269.600 442.000 270.400 ;
        RECT 444.400 269.600 445.200 271.200 ;
        RECT 446.200 270.600 448.200 271.200 ;
        RECT 447.600 270.400 448.200 270.600 ;
        RECT 450.000 270.400 450.800 270.800 ;
        RECT 447.600 269.600 448.400 270.400 ;
        RECT 450.000 269.800 451.600 270.400 ;
        RECT 450.800 269.600 451.600 269.800 ;
        RECT 446.200 268.800 447.000 269.600 ;
        RECT 446.200 268.400 446.800 268.800 ;
        RECT 438.200 268.200 439.800 268.400 ;
        RECT 438.200 267.800 440.000 268.200 ;
        RECT 397.800 262.200 399.400 266.200 ;
        RECT 405.800 262.200 407.400 266.200 ;
        RECT 412.400 265.600 414.200 266.200 ;
        RECT 413.400 262.200 414.200 265.600 ;
        RECT 418.200 262.200 419.800 266.200 ;
        RECT 426.200 262.200 427.800 266.200 ;
        RECT 435.200 262.200 436.000 267.800 ;
        RECT 439.200 262.200 440.000 267.800 ;
        RECT 446.000 267.600 446.800 268.400 ;
        RECT 447.600 266.200 448.200 269.600 ;
        RECT 449.200 267.600 450.000 269.200 ;
        RECT 452.600 268.400 453.200 271.600 ;
        RECT 457.200 270.800 458.000 272.400 ;
        RECT 463.600 270.800 464.400 272.400 ;
        RECT 468.400 271.600 469.200 272.400 ;
        RECT 470.000 272.300 470.800 272.400 ;
        RECT 471.600 272.300 472.400 272.400 ;
        RECT 470.000 271.700 472.400 272.300 ;
        RECT 454.000 269.600 456.400 270.400 ;
        RECT 465.200 269.600 466.800 270.400 ;
        RECT 468.400 268.400 469.000 271.600 ;
        RECT 470.000 270.800 470.800 271.700 ;
        RECT 471.600 271.600 472.400 271.700 ;
        RECT 474.800 271.600 475.600 272.400 ;
        RECT 471.600 269.600 473.200 270.400 ;
        RECT 474.800 268.400 475.400 271.600 ;
        RECT 476.400 270.800 477.200 272.400 ;
        RECT 481.200 271.600 482.000 272.400 ;
        RECT 483.400 271.800 485.200 272.600 ;
        RECT 490.200 271.800 492.200 277.600 ;
        RECT 495.600 272.400 496.400 279.800 ;
        RECT 498.800 272.400 499.600 279.800 ;
        RECT 495.600 271.800 499.600 272.400 ;
        RECT 500.400 271.800 501.200 279.800 ;
        RECT 504.600 278.400 505.400 279.800 ;
        RECT 504.600 277.600 506.000 278.400 ;
        RECT 504.600 272.600 505.400 277.600 ;
        RECT 509.000 274.400 509.800 279.800 ;
        RECT 503.600 271.800 505.400 272.600 ;
        RECT 507.600 273.600 508.400 274.400 ;
        RECT 509.000 273.600 510.800 274.400 ;
        RECT 507.600 272.400 508.200 273.600 ;
        RECT 509.000 272.400 509.800 273.600 ;
        RECT 515.800 272.600 516.600 279.800 ;
        RECT 506.800 271.800 508.200 272.400 ;
        RECT 508.800 271.800 509.800 272.400 ;
        RECT 514.800 271.800 516.600 272.600 ;
        RECT 518.600 272.600 519.400 279.800 ;
        RECT 525.400 278.400 526.200 279.800 ;
        RECT 531.800 278.400 533.800 279.800 ;
        RECT 524.400 277.600 526.200 278.400 ;
        RECT 530.800 277.600 533.800 278.400 ;
        RECT 518.600 271.800 520.400 272.600 ;
        RECT 525.400 272.400 526.200 277.600 ;
        RECT 526.800 273.600 527.600 274.400 ;
        RECT 527.000 272.400 527.600 273.600 ;
        RECT 525.400 271.800 526.400 272.400 ;
        RECT 527.000 271.800 528.400 272.400 ;
        RECT 531.800 271.800 533.800 277.600 ;
        RECT 478.000 269.600 479.600 270.400 ;
        RECT 481.200 268.400 481.800 271.600 ;
        RECT 482.800 269.600 483.600 271.200 ;
        RECT 452.600 268.200 454.200 268.400 ;
        RECT 467.400 268.200 469.000 268.400 ;
        RECT 473.800 268.200 475.400 268.400 ;
        RECT 480.200 268.200 481.800 268.400 ;
        RECT 452.600 267.800 454.400 268.200 ;
        RECT 447.000 262.200 448.600 266.200 ;
        RECT 453.600 262.200 454.400 267.800 ;
        RECT 467.200 267.800 469.000 268.200 ;
        RECT 473.600 267.800 475.400 268.200 ;
        RECT 480.000 267.800 481.800 268.200 ;
        RECT 484.400 268.400 485.000 271.800 ;
        RECT 467.200 262.200 468.000 267.800 ;
        RECT 473.600 262.200 474.400 267.800 ;
        RECT 480.000 262.200 480.800 267.800 ;
        RECT 484.400 267.600 485.200 268.400 ;
        RECT 487.600 267.600 488.400 269.200 ;
        RECT 489.200 268.800 490.000 270.400 ;
        RECT 491.000 268.400 491.600 271.800 ;
        RECT 496.400 270.400 497.200 270.800 ;
        RECT 500.400 270.400 501.000 271.800 ;
        RECT 492.400 268.800 493.200 270.400 ;
        RECT 495.600 269.800 497.200 270.400 ;
        RECT 498.800 269.800 501.200 270.400 ;
        RECT 495.600 269.600 496.400 269.800 ;
        RECT 490.800 268.200 491.600 268.400 ;
        RECT 494.000 268.200 494.800 268.400 ;
        RECT 489.200 267.600 491.600 268.200 ;
        RECT 493.200 267.600 494.800 268.200 ;
        RECT 497.200 267.600 498.000 269.200 ;
        RECT 484.400 264.400 485.000 267.600 ;
        RECT 486.000 264.800 486.800 266.400 ;
        RECT 489.200 266.200 489.800 267.600 ;
        RECT 493.200 267.200 494.000 267.600 ;
        RECT 491.000 266.200 494.600 266.600 ;
        RECT 498.800 266.200 499.400 269.800 ;
        RECT 500.400 269.600 501.200 269.800 ;
        RECT 503.800 268.400 504.400 271.800 ;
        RECT 506.800 271.600 507.600 271.800 ;
        RECT 505.200 269.600 506.000 271.200 ;
        RECT 508.800 268.400 509.400 271.800 ;
        RECT 510.000 270.300 510.800 270.400 ;
        RECT 511.600 270.300 512.400 270.400 ;
        RECT 510.000 269.700 512.400 270.300 ;
        RECT 510.000 268.800 510.800 269.700 ;
        RECT 511.600 269.600 512.400 269.700 ;
        RECT 515.000 268.400 515.600 271.800 ;
        RECT 516.400 269.600 517.200 271.200 ;
        RECT 518.000 269.600 518.800 271.200 ;
        RECT 519.600 270.300 520.200 271.800 ;
        RECT 524.400 270.300 525.200 270.400 ;
        RECT 519.600 269.700 525.200 270.300 ;
        RECT 503.600 267.600 504.400 268.400 ;
        RECT 506.800 267.600 509.400 268.400 ;
        RECT 511.600 268.200 512.400 268.400 ;
        RECT 510.800 267.600 512.400 268.200 ;
        RECT 514.800 268.300 515.600 268.400 ;
        RECT 518.100 268.300 518.700 269.600 ;
        RECT 514.800 267.700 518.700 268.300 ;
        RECT 519.600 268.400 520.200 269.700 ;
        RECT 524.400 268.800 525.200 269.700 ;
        RECT 525.800 268.400 526.400 271.800 ;
        RECT 527.600 271.600 528.400 271.800 ;
        RECT 530.800 268.800 531.600 270.400 ;
        RECT 532.400 268.400 533.000 271.800 ;
        RECT 537.200 271.600 538.000 273.200 ;
        RECT 534.000 268.800 534.800 270.400 ;
        RECT 514.800 267.600 515.600 267.700 ;
        RECT 484.400 262.200 485.200 264.400 ;
        RECT 487.600 262.800 488.400 266.200 ;
        RECT 489.200 263.400 490.000 266.200 ;
        RECT 490.800 266.000 494.800 266.200 ;
        RECT 490.800 262.800 491.600 266.000 ;
        RECT 487.600 262.200 491.600 262.800 ;
        RECT 494.000 262.200 494.800 266.000 ;
        RECT 498.800 262.200 499.600 266.200 ;
        RECT 500.400 265.600 501.200 266.400 ;
        RECT 500.200 264.800 501.000 265.600 ;
        RECT 502.000 264.800 502.800 266.400 ;
        RECT 503.800 264.200 504.400 267.600 ;
        RECT 507.000 266.200 507.600 267.600 ;
        RECT 510.800 267.200 511.600 267.600 ;
        RECT 508.600 266.200 512.200 266.600 ;
        RECT 515.000 266.400 515.600 267.600 ;
        RECT 503.600 262.200 504.400 264.200 ;
        RECT 506.800 262.200 507.600 266.200 ;
        RECT 508.400 266.000 512.400 266.200 ;
        RECT 508.400 262.200 509.200 266.000 ;
        RECT 511.600 262.200 512.400 266.000 ;
        RECT 513.200 264.800 514.000 266.400 ;
        RECT 514.800 265.600 515.600 266.400 ;
        RECT 515.000 264.200 515.600 265.600 ;
        RECT 514.800 262.200 515.600 264.200 ;
        RECT 519.600 267.600 520.400 268.400 ;
        RECT 522.800 268.200 523.600 268.400 ;
        RECT 522.800 267.600 524.400 268.200 ;
        RECT 525.800 267.600 528.400 268.400 ;
        RECT 529.200 268.200 530.000 268.400 ;
        RECT 532.400 268.200 533.200 268.400 ;
        RECT 529.200 267.600 530.800 268.200 ;
        RECT 532.400 267.600 534.800 268.200 ;
        RECT 535.600 267.600 536.400 269.200 ;
        RECT 519.600 264.200 520.200 267.600 ;
        RECT 523.600 267.200 524.400 267.600 ;
        RECT 521.200 264.800 522.000 266.400 ;
        RECT 523.000 266.200 526.600 266.600 ;
        RECT 527.600 266.200 528.200 267.600 ;
        RECT 530.000 267.200 530.800 267.600 ;
        RECT 529.400 266.200 533.000 266.600 ;
        RECT 534.200 266.200 534.800 267.600 ;
        RECT 538.800 266.200 539.600 279.800 ;
        RECT 540.400 266.800 541.200 268.400 ;
        RECT 522.800 266.000 526.800 266.200 ;
        RECT 519.600 262.200 520.400 264.200 ;
        RECT 522.800 262.200 523.600 266.000 ;
        RECT 526.000 262.200 526.800 266.000 ;
        RECT 527.600 262.200 528.400 266.200 ;
        RECT 529.200 266.000 533.200 266.200 ;
        RECT 529.200 262.200 530.000 266.000 ;
        RECT 532.400 262.800 533.200 266.000 ;
        RECT 534.000 263.400 534.800 266.200 ;
        RECT 535.600 262.800 536.400 266.200 ;
        RECT 532.400 262.200 536.400 262.800 ;
        RECT 537.800 265.600 539.600 266.200 ;
        RECT 537.800 264.400 538.600 265.600 ;
        RECT 537.800 263.600 539.600 264.400 ;
        RECT 537.800 262.200 538.600 263.600 ;
        RECT 542.000 262.200 542.800 279.800 ;
        RECT 545.200 271.600 546.000 273.200 ;
        RECT 543.600 264.800 544.400 266.400 ;
        RECT 546.800 266.200 547.600 279.800 ;
        RECT 550.000 271.600 550.800 273.200 ;
        RECT 548.400 266.800 549.200 268.400 ;
        RECT 551.600 266.200 552.400 279.800 ;
        RECT 557.400 272.400 558.200 279.800 ;
        RECT 558.800 273.600 559.600 274.400 ;
        RECT 559.000 272.400 559.600 273.600 ;
        RECT 557.400 271.800 558.400 272.400 ;
        RECT 559.000 272.300 560.400 272.400 ;
        RECT 561.200 272.300 562.000 272.400 ;
        RECT 559.000 271.800 562.000 272.300 ;
        RECT 556.400 268.800 557.200 270.400 ;
        RECT 557.800 268.400 558.400 271.800 ;
        RECT 559.600 271.700 562.000 271.800 ;
        RECT 559.600 271.600 560.400 271.700 ;
        RECT 561.200 271.600 562.000 271.700 ;
        RECT 553.200 268.300 554.000 268.400 ;
        RECT 554.800 268.300 555.600 268.400 ;
        RECT 553.200 268.200 555.600 268.300 ;
        RECT 557.800 268.300 560.400 268.400 ;
        RECT 561.200 268.300 562.000 268.400 ;
        RECT 553.200 267.700 556.400 268.200 ;
        RECT 553.200 266.800 554.000 267.700 ;
        RECT 554.800 267.600 556.400 267.700 ;
        RECT 557.800 267.700 562.000 268.300 ;
        RECT 557.800 267.600 560.400 267.700 ;
        RECT 555.600 267.200 556.400 267.600 ;
        RECT 555.000 266.200 558.600 266.600 ;
        RECT 559.600 266.200 560.200 267.600 ;
        RECT 561.200 266.800 562.000 267.700 ;
        RECT 562.800 266.200 563.600 279.800 ;
        RECT 564.400 271.600 565.200 273.200 ;
        RECT 568.600 272.400 569.400 279.800 ;
        RECT 570.000 274.300 570.800 274.400 ;
        RECT 572.400 274.300 573.200 274.400 ;
        RECT 570.000 273.700 573.200 274.300 ;
        RECT 570.000 273.600 570.800 273.700 ;
        RECT 572.400 273.600 573.200 273.700 ;
        RECT 570.200 272.400 570.800 273.600 ;
        RECT 568.600 271.800 569.600 272.400 ;
        RECT 570.200 271.800 571.600 272.400 ;
        RECT 567.600 268.800 568.400 270.400 ;
        RECT 569.000 268.400 569.600 271.800 ;
        RECT 570.800 271.600 571.600 271.800 ;
        RECT 564.400 268.300 565.200 268.400 ;
        RECT 566.000 268.300 566.800 268.400 ;
        RECT 564.400 268.200 566.800 268.300 ;
        RECT 569.000 268.300 571.600 268.400 ;
        RECT 572.400 268.300 573.200 268.400 ;
        RECT 564.400 267.700 567.600 268.200 ;
        RECT 564.400 267.600 565.200 267.700 ;
        RECT 566.000 267.600 567.600 267.700 ;
        RECT 569.000 267.700 573.200 268.300 ;
        RECT 569.000 267.600 571.600 267.700 ;
        RECT 566.800 267.200 567.600 267.600 ;
        RECT 566.200 266.200 569.800 266.600 ;
        RECT 570.800 266.200 571.400 267.600 ;
        RECT 572.400 266.800 573.200 267.700 ;
        RECT 574.000 268.300 574.800 279.800 ;
        RECT 575.600 271.600 576.400 273.200 ;
        RECT 578.800 272.000 579.600 279.800 ;
        RECT 582.000 275.200 582.800 279.800 ;
        RECT 578.600 271.200 579.600 272.000 ;
        RECT 580.200 274.600 582.800 275.200 ;
        RECT 580.200 273.000 580.800 274.600 ;
        RECT 585.200 274.400 586.000 279.800 ;
        RECT 588.400 277.000 589.200 279.800 ;
        RECT 590.000 277.000 590.800 279.800 ;
        RECT 591.600 277.000 592.400 279.800 ;
        RECT 586.600 274.400 590.800 275.200 ;
        RECT 583.400 273.600 586.000 274.400 ;
        RECT 593.200 273.600 594.000 279.800 ;
        RECT 596.400 275.000 597.200 279.800 ;
        RECT 599.600 275.000 600.400 279.800 ;
        RECT 601.200 277.000 602.000 279.800 ;
        RECT 602.800 277.000 603.600 279.800 ;
        RECT 606.000 275.200 606.800 279.800 ;
        RECT 609.200 276.400 610.000 279.800 ;
        RECT 609.200 275.800 610.200 276.400 ;
        RECT 609.600 275.200 610.200 275.800 ;
        RECT 604.800 274.400 609.000 275.200 ;
        RECT 609.600 274.600 611.600 275.200 ;
        RECT 596.400 273.600 599.000 274.400 ;
        RECT 599.600 273.800 605.400 274.400 ;
        RECT 608.400 274.000 609.000 274.400 ;
        RECT 588.400 273.000 589.200 273.200 ;
        RECT 580.200 272.400 589.200 273.000 ;
        RECT 591.600 273.000 592.400 273.200 ;
        RECT 599.600 273.000 600.200 273.800 ;
        RECT 606.000 273.200 607.400 273.800 ;
        RECT 608.400 273.200 610.000 274.000 ;
        RECT 591.600 272.400 600.200 273.000 ;
        RECT 601.200 273.000 607.400 273.200 ;
        RECT 601.200 272.600 606.600 273.000 ;
        RECT 601.200 272.400 602.000 272.600 ;
        RECT 577.200 268.300 578.000 268.400 ;
        RECT 574.000 267.700 578.000 268.300 ;
        RECT 574.000 266.200 574.800 267.700 ;
        RECT 577.200 267.600 578.000 267.700 ;
        RECT 578.600 266.800 579.400 271.200 ;
        RECT 580.200 270.600 580.800 272.400 ;
        RECT 580.000 270.000 580.800 270.600 ;
        RECT 586.800 270.000 610.200 270.600 ;
        RECT 580.000 268.000 580.600 270.000 ;
        RECT 586.800 269.400 587.600 270.000 ;
        RECT 604.400 269.600 605.200 270.000 ;
        RECT 609.400 269.800 610.200 270.000 ;
        RECT 581.200 268.600 585.000 269.400 ;
        RECT 580.000 267.400 581.200 268.000 ;
        RECT 545.800 265.600 547.600 266.200 ;
        RECT 550.600 265.600 552.400 266.200 ;
        RECT 554.800 266.000 558.800 266.200 ;
        RECT 545.800 264.400 546.600 265.600 ;
        RECT 545.200 263.600 546.600 264.400 ;
        RECT 545.800 262.200 546.600 263.600 ;
        RECT 550.600 264.400 551.400 265.600 ;
        RECT 550.600 263.600 552.400 264.400 ;
        RECT 550.600 262.200 551.400 263.600 ;
        RECT 554.800 262.200 555.600 266.000 ;
        RECT 558.000 262.200 558.800 266.000 ;
        RECT 559.600 262.200 560.400 266.200 ;
        RECT 562.800 265.600 564.600 266.200 ;
        RECT 563.800 264.400 564.600 265.600 ;
        RECT 566.000 266.000 570.000 266.200 ;
        RECT 563.800 263.600 565.200 264.400 ;
        RECT 563.800 262.200 564.600 263.600 ;
        RECT 566.000 262.200 566.800 266.000 ;
        RECT 569.200 262.200 570.000 266.000 ;
        RECT 570.800 262.200 571.600 266.200 ;
        RECT 574.000 265.600 575.800 266.200 ;
        RECT 578.600 266.000 579.600 266.800 ;
        RECT 575.000 262.200 575.800 265.600 ;
        RECT 578.800 262.200 579.600 266.000 ;
        RECT 580.400 262.200 581.200 267.400 ;
        RECT 584.200 267.400 585.000 268.600 ;
        RECT 584.200 266.800 586.000 267.400 ;
        RECT 585.200 266.200 586.000 266.800 ;
        RECT 590.000 266.400 590.800 269.200 ;
        RECT 593.200 268.600 596.400 269.400 ;
        RECT 600.200 268.600 602.200 269.400 ;
        RECT 610.800 269.000 611.600 274.600 ;
        RECT 592.800 267.800 593.600 268.000 ;
        RECT 592.800 267.200 597.200 267.800 ;
        RECT 596.400 267.000 597.200 267.200 ;
        RECT 598.000 266.800 598.800 268.400 ;
        RECT 585.200 265.400 587.600 266.200 ;
        RECT 590.000 265.600 591.000 266.400 ;
        RECT 594.000 265.600 595.600 266.400 ;
        RECT 596.400 266.200 597.200 266.400 ;
        RECT 600.200 266.200 601.000 268.600 ;
        RECT 602.800 268.200 611.600 269.000 ;
        RECT 606.200 266.800 609.200 267.600 ;
        RECT 606.200 266.200 607.000 266.800 ;
        RECT 596.400 265.600 601.000 266.200 ;
        RECT 586.800 262.200 587.600 265.400 ;
        RECT 604.400 265.400 607.000 266.200 ;
        RECT 588.400 262.200 589.200 265.000 ;
        RECT 590.000 262.200 590.800 265.000 ;
        RECT 591.600 262.200 592.400 265.000 ;
        RECT 593.200 262.200 594.000 265.000 ;
        RECT 596.400 262.200 597.200 265.000 ;
        RECT 599.600 262.200 600.400 265.000 ;
        RECT 601.200 262.200 602.000 265.000 ;
        RECT 602.800 262.200 603.600 265.000 ;
        RECT 604.400 262.200 605.200 265.400 ;
        RECT 610.800 262.200 611.600 268.200 ;
        RECT 1.200 253.800 2.000 259.800 ;
        RECT 7.600 256.600 8.400 259.800 ;
        RECT 9.200 257.000 10.000 259.800 ;
        RECT 10.800 257.000 11.600 259.800 ;
        RECT 12.400 257.000 13.200 259.800 ;
        RECT 15.600 257.000 16.400 259.800 ;
        RECT 18.800 257.000 19.600 259.800 ;
        RECT 20.400 257.000 21.200 259.800 ;
        RECT 22.000 257.000 22.800 259.800 ;
        RECT 23.600 257.000 24.400 259.800 ;
        RECT 5.800 255.800 8.400 256.600 ;
        RECT 25.200 256.600 26.000 259.800 ;
        RECT 11.800 255.800 16.400 256.400 ;
        RECT 5.800 255.200 6.600 255.800 ;
        RECT 3.600 254.400 6.600 255.200 ;
        RECT 1.200 253.000 10.000 253.800 ;
        RECT 11.800 253.400 12.600 255.800 ;
        RECT 15.600 255.600 16.400 255.800 ;
        RECT 17.200 255.600 18.800 256.400 ;
        RECT 21.800 255.600 22.800 256.400 ;
        RECT 25.200 255.800 27.600 256.600 ;
        RECT 14.000 253.600 14.800 255.200 ;
        RECT 15.600 254.800 16.400 255.000 ;
        RECT 15.600 254.200 20.000 254.800 ;
        RECT 19.200 254.000 20.000 254.200 ;
        RECT 1.200 247.400 2.000 253.000 ;
        RECT 10.600 252.600 12.600 253.400 ;
        RECT 16.400 252.600 19.600 253.400 ;
        RECT 22.000 252.800 22.800 255.600 ;
        RECT 26.800 255.200 27.600 255.800 ;
        RECT 26.800 254.600 28.600 255.200 ;
        RECT 27.800 253.400 28.600 254.600 ;
        RECT 31.600 254.600 32.400 259.800 ;
        RECT 33.200 256.000 34.000 259.800 ;
        RECT 33.200 255.200 34.200 256.000 ;
        RECT 31.600 254.000 32.800 254.600 ;
        RECT 27.800 252.600 31.600 253.400 ;
        RECT 2.600 252.000 3.400 252.200 ;
        RECT 7.600 252.000 8.400 252.400 ;
        RECT 25.200 252.000 26.000 252.600 ;
        RECT 32.200 252.000 32.800 254.000 ;
        RECT 2.600 251.400 26.000 252.000 ;
        RECT 32.000 251.400 32.800 252.000 ;
        RECT 32.000 249.600 32.600 251.400 ;
        RECT 33.400 250.800 34.200 255.200 ;
        RECT 10.800 249.400 11.600 249.600 ;
        RECT 6.200 249.000 11.600 249.400 ;
        RECT 5.400 248.800 11.600 249.000 ;
        RECT 12.600 249.000 21.200 249.600 ;
        RECT 2.800 248.000 4.400 248.800 ;
        RECT 5.400 248.200 6.800 248.800 ;
        RECT 12.600 248.200 13.200 249.000 ;
        RECT 20.400 248.800 21.200 249.000 ;
        RECT 23.600 249.000 32.600 249.600 ;
        RECT 23.600 248.800 24.400 249.000 ;
        RECT 3.800 247.600 4.400 248.000 ;
        RECT 7.400 247.600 13.200 248.200 ;
        RECT 13.800 247.600 16.400 248.400 ;
        RECT 1.200 246.800 3.200 247.400 ;
        RECT 3.800 246.800 8.000 247.600 ;
        RECT 2.600 246.200 3.200 246.800 ;
        RECT 2.600 245.600 3.600 246.200 ;
        RECT 2.800 242.200 3.600 245.600 ;
        RECT 6.000 242.200 6.800 246.800 ;
        RECT 9.200 242.200 10.000 245.000 ;
        RECT 10.800 242.200 11.600 245.000 ;
        RECT 12.400 242.200 13.200 247.000 ;
        RECT 15.600 242.200 16.400 247.000 ;
        RECT 18.800 242.200 19.600 248.400 ;
        RECT 26.800 247.600 29.400 248.400 ;
        RECT 22.000 246.800 26.200 247.600 ;
        RECT 20.400 242.200 21.200 245.000 ;
        RECT 22.000 242.200 22.800 245.000 ;
        RECT 23.600 242.200 24.400 245.000 ;
        RECT 26.800 242.200 27.600 247.600 ;
        RECT 32.000 247.400 32.600 249.000 ;
        RECT 30.000 246.800 32.600 247.400 ;
        RECT 33.200 250.000 34.200 250.800 ;
        RECT 30.000 242.200 30.800 246.800 ;
        RECT 33.200 242.200 34.000 250.000 ;
        RECT 34.800 248.300 35.600 248.400 ;
        RECT 36.400 248.300 37.200 259.800 ;
        RECT 38.000 255.600 38.800 257.200 ;
        RECT 34.800 247.700 37.200 248.300 ;
        RECT 34.800 247.600 35.600 247.700 ;
        RECT 36.400 242.200 37.200 247.700 ;
        RECT 39.600 253.800 40.400 259.800 ;
        RECT 46.000 256.600 46.800 259.800 ;
        RECT 47.600 257.000 48.400 259.800 ;
        RECT 49.200 257.000 50.000 259.800 ;
        RECT 50.800 257.000 51.600 259.800 ;
        RECT 54.000 257.000 54.800 259.800 ;
        RECT 57.200 257.000 58.000 259.800 ;
        RECT 58.800 257.000 59.600 259.800 ;
        RECT 60.400 257.000 61.200 259.800 ;
        RECT 62.000 257.000 62.800 259.800 ;
        RECT 44.200 255.800 46.800 256.600 ;
        RECT 63.600 256.600 64.400 259.800 ;
        RECT 50.200 255.800 54.800 256.400 ;
        RECT 44.200 255.200 45.000 255.800 ;
        RECT 42.000 254.400 45.000 255.200 ;
        RECT 39.600 253.000 48.400 253.800 ;
        RECT 50.200 253.400 51.000 255.800 ;
        RECT 54.000 255.600 54.800 255.800 ;
        RECT 55.600 255.600 57.200 256.400 ;
        RECT 60.200 255.600 61.200 256.400 ;
        RECT 63.600 255.800 66.000 256.600 ;
        RECT 52.400 253.600 53.200 255.200 ;
        RECT 54.000 254.800 54.800 255.000 ;
        RECT 54.000 254.200 58.400 254.800 ;
        RECT 57.600 254.000 58.400 254.200 ;
        RECT 39.600 247.400 40.400 253.000 ;
        RECT 49.000 252.600 51.000 253.400 ;
        RECT 54.800 252.600 58.000 253.400 ;
        RECT 60.400 252.800 61.200 255.600 ;
        RECT 65.200 255.200 66.000 255.800 ;
        RECT 65.200 254.600 67.000 255.200 ;
        RECT 66.200 253.400 67.000 254.600 ;
        RECT 70.000 254.600 70.800 259.800 ;
        RECT 71.600 256.000 72.400 259.800 ;
        RECT 76.400 257.800 77.200 259.800 ;
        RECT 71.600 255.200 72.600 256.000 ;
        RECT 74.800 255.600 75.600 257.200 ;
        RECT 76.600 256.300 77.200 257.800 ;
        RECT 79.800 256.400 80.600 257.200 ;
        RECT 79.600 256.300 80.400 256.400 ;
        RECT 76.500 255.700 80.400 256.300 ;
        RECT 81.200 255.800 82.000 259.800 ;
        RECT 70.000 254.000 71.200 254.600 ;
        RECT 66.200 252.600 70.000 253.400 ;
        RECT 41.200 252.200 42.000 252.400 ;
        RECT 41.000 252.000 42.000 252.200 ;
        RECT 46.000 252.000 46.800 252.400 ;
        RECT 63.600 252.000 64.400 252.600 ;
        RECT 70.600 252.000 71.200 254.000 ;
        RECT 41.000 251.400 64.400 252.000 ;
        RECT 70.400 251.400 71.200 252.000 ;
        RECT 70.400 249.600 71.000 251.400 ;
        RECT 71.800 250.800 72.600 255.200 ;
        RECT 76.600 254.400 77.200 255.700 ;
        RECT 79.600 255.600 80.400 255.700 ;
        RECT 76.400 253.600 77.200 254.400 ;
        RECT 49.200 249.400 50.000 249.600 ;
        RECT 44.600 249.000 50.000 249.400 ;
        RECT 43.800 248.800 50.000 249.000 ;
        RECT 51.000 249.000 59.600 249.600 ;
        RECT 41.200 248.000 42.800 248.800 ;
        RECT 43.800 248.200 45.200 248.800 ;
        RECT 51.000 248.200 51.600 249.000 ;
        RECT 58.800 248.800 59.600 249.000 ;
        RECT 62.000 249.000 71.000 249.600 ;
        RECT 62.000 248.800 62.800 249.000 ;
        RECT 42.200 247.600 42.800 248.000 ;
        RECT 45.800 247.600 51.600 248.200 ;
        RECT 52.200 247.600 54.800 248.400 ;
        RECT 39.600 246.800 41.600 247.400 ;
        RECT 42.200 246.800 46.400 247.600 ;
        RECT 41.000 246.200 41.600 246.800 ;
        RECT 41.000 245.600 42.000 246.200 ;
        RECT 41.200 242.200 42.000 245.600 ;
        RECT 44.400 242.200 45.200 246.800 ;
        RECT 47.600 242.200 48.400 245.000 ;
        RECT 49.200 242.200 50.000 245.000 ;
        RECT 50.800 242.200 51.600 247.000 ;
        RECT 54.000 242.200 54.800 247.000 ;
        RECT 57.200 242.200 58.000 248.400 ;
        RECT 65.200 247.600 67.800 248.400 ;
        RECT 60.400 246.800 64.600 247.600 ;
        RECT 58.800 242.200 59.600 245.000 ;
        RECT 60.400 242.200 61.200 245.000 ;
        RECT 62.000 242.200 62.800 245.000 ;
        RECT 65.200 242.200 66.000 247.600 ;
        RECT 70.400 247.400 71.000 249.000 ;
        RECT 68.400 246.800 71.000 247.400 ;
        RECT 71.600 250.000 72.600 250.800 ;
        RECT 76.600 250.200 77.200 253.600 ;
        RECT 78.000 250.800 78.800 252.400 ;
        RECT 79.600 252.200 80.400 252.400 ;
        RECT 81.400 252.200 82.000 255.800 ;
        RECT 82.800 252.800 83.600 254.400 ;
        RECT 84.400 252.200 85.200 252.400 ;
        RECT 79.600 251.600 82.000 252.200 ;
        RECT 83.600 251.600 85.200 252.200 ;
        RECT 79.800 250.200 80.400 251.600 ;
        RECT 83.600 251.200 84.400 251.600 ;
        RECT 68.400 242.200 69.200 246.800 ;
        RECT 71.600 242.200 72.400 250.000 ;
        RECT 76.400 249.400 78.200 250.200 ;
        RECT 77.400 242.200 78.200 249.400 ;
        RECT 79.600 242.200 80.400 250.200 ;
        RECT 81.200 249.600 85.200 250.200 ;
        RECT 81.200 242.200 82.000 249.600 ;
        RECT 84.400 242.200 85.200 249.600 ;
        RECT 86.000 242.200 86.800 259.800 ;
        RECT 90.800 257.600 91.600 259.800 ;
        RECT 87.600 256.300 88.400 257.200 ;
        RECT 89.200 256.300 90.000 256.400 ;
        RECT 87.600 255.700 90.000 256.300 ;
        RECT 87.600 255.600 88.400 255.700 ;
        RECT 89.200 255.600 90.000 255.700 ;
        RECT 90.800 254.400 91.400 257.600 ;
        RECT 92.400 256.300 93.200 257.200 ;
        RECT 95.600 256.300 96.400 259.800 ;
        RECT 92.400 255.700 96.400 256.300 ;
        RECT 92.400 255.600 93.200 255.700 ;
        RECT 95.400 255.200 96.400 255.700 ;
        RECT 90.800 253.600 91.600 254.400 ;
        RECT 87.600 252.300 88.400 252.400 ;
        RECT 89.200 252.300 90.000 252.400 ;
        RECT 87.600 251.700 90.000 252.300 ;
        RECT 87.600 251.600 88.400 251.700 ;
        RECT 89.200 250.800 90.000 251.700 ;
        RECT 90.800 250.200 91.400 253.600 ;
        RECT 95.400 250.800 96.200 255.200 ;
        RECT 97.200 254.600 98.000 259.800 ;
        RECT 103.600 256.600 104.400 259.800 ;
        RECT 105.200 257.000 106.000 259.800 ;
        RECT 106.800 257.000 107.600 259.800 ;
        RECT 108.400 257.000 109.200 259.800 ;
        RECT 110.000 257.000 110.800 259.800 ;
        RECT 113.200 257.000 114.000 259.800 ;
        RECT 116.400 257.000 117.200 259.800 ;
        RECT 118.000 257.000 118.800 259.800 ;
        RECT 119.600 257.000 120.400 259.800 ;
        RECT 102.000 255.800 104.400 256.600 ;
        RECT 121.200 256.600 122.000 259.800 ;
        RECT 102.000 255.200 102.800 255.800 ;
        RECT 96.800 254.000 98.000 254.600 ;
        RECT 101.000 254.600 102.800 255.200 ;
        RECT 106.800 255.600 107.800 256.400 ;
        RECT 110.800 255.600 112.400 256.400 ;
        RECT 113.200 255.800 117.800 256.400 ;
        RECT 121.200 255.800 123.800 256.600 ;
        RECT 113.200 255.600 114.000 255.800 ;
        RECT 96.800 252.000 97.400 254.000 ;
        RECT 101.000 253.400 101.800 254.600 ;
        RECT 98.000 252.600 101.800 253.400 ;
        RECT 106.800 252.800 107.600 255.600 ;
        RECT 113.200 254.800 114.000 255.000 ;
        RECT 109.600 254.200 114.000 254.800 ;
        RECT 109.600 254.000 110.400 254.200 ;
        RECT 114.800 253.600 115.600 255.200 ;
        RECT 117.000 253.400 117.800 255.800 ;
        RECT 123.000 255.200 123.800 255.800 ;
        RECT 123.000 254.400 126.000 255.200 ;
        RECT 127.600 253.800 128.400 259.800 ;
        RECT 110.000 252.600 113.200 253.400 ;
        RECT 117.000 252.600 119.000 253.400 ;
        RECT 119.600 253.000 128.400 253.800 ;
        RECT 103.600 252.000 104.400 252.600 ;
        RECT 121.200 252.000 122.000 252.400 ;
        RECT 124.400 252.000 125.200 252.400 ;
        RECT 126.200 252.000 127.000 252.200 ;
        RECT 96.800 251.400 97.600 252.000 ;
        RECT 103.600 251.400 127.000 252.000 ;
        RECT 89.800 249.400 91.600 250.200 ;
        RECT 95.400 250.000 96.400 250.800 ;
        RECT 89.800 242.200 90.600 249.400 ;
        RECT 95.600 242.200 96.400 250.000 ;
        RECT 97.000 249.600 97.600 251.400 ;
        RECT 97.000 249.000 106.000 249.600 ;
        RECT 97.000 247.400 97.600 249.000 ;
        RECT 105.200 248.800 106.000 249.000 ;
        RECT 108.400 249.000 117.000 249.600 ;
        RECT 108.400 248.800 109.200 249.000 ;
        RECT 100.200 247.600 102.800 248.400 ;
        RECT 97.000 246.800 99.600 247.400 ;
        RECT 98.800 242.200 99.600 246.800 ;
        RECT 102.000 242.200 102.800 247.600 ;
        RECT 103.400 246.800 107.600 247.600 ;
        RECT 105.200 242.200 106.000 245.000 ;
        RECT 106.800 242.200 107.600 245.000 ;
        RECT 108.400 242.200 109.200 245.000 ;
        RECT 110.000 242.200 110.800 248.400 ;
        RECT 113.200 247.600 115.800 248.400 ;
        RECT 116.400 248.200 117.000 249.000 ;
        RECT 118.000 249.400 118.800 249.600 ;
        RECT 118.000 249.000 123.400 249.400 ;
        RECT 118.000 248.800 124.200 249.000 ;
        RECT 122.800 248.200 124.200 248.800 ;
        RECT 116.400 247.600 122.200 248.200 ;
        RECT 125.200 248.000 126.800 248.800 ;
        RECT 125.200 247.600 125.800 248.000 ;
        RECT 113.200 242.200 114.000 247.000 ;
        RECT 116.400 242.200 117.200 247.000 ;
        RECT 121.600 246.800 125.800 247.600 ;
        RECT 127.600 247.400 128.400 253.000 ;
        RECT 126.400 246.800 128.400 247.400 ;
        RECT 118.000 242.200 118.800 245.000 ;
        RECT 119.600 242.200 120.400 245.000 ;
        RECT 122.800 242.200 123.600 246.800 ;
        RECT 126.400 246.200 127.000 246.800 ;
        RECT 126.000 245.600 127.000 246.200 ;
        RECT 126.000 242.200 126.800 245.600 ;
        RECT 129.200 242.200 130.000 259.800 ;
        RECT 130.800 255.600 131.600 257.200 ;
        RECT 134.000 256.400 134.800 259.800 ;
        RECT 133.800 255.800 134.800 256.400 ;
        RECT 133.800 254.400 134.400 255.800 ;
        RECT 137.200 255.200 138.000 259.800 ;
        RECT 145.200 256.000 146.000 259.800 ;
        RECT 135.400 254.600 138.000 255.200 ;
        RECT 145.000 255.200 146.000 256.000 ;
        RECT 130.800 254.300 131.600 254.400 ;
        RECT 133.800 254.300 134.800 254.400 ;
        RECT 130.800 253.700 134.800 254.300 ;
        RECT 130.800 253.600 131.600 253.700 ;
        RECT 133.800 253.600 134.800 253.700 ;
        RECT 133.800 250.200 134.400 253.600 ;
        RECT 135.400 253.000 136.000 254.600 ;
        RECT 135.000 252.200 136.000 253.000 ;
        RECT 135.400 250.200 136.000 252.200 ;
        RECT 137.000 252.400 137.800 253.200 ;
        RECT 137.000 251.600 138.000 252.400 ;
        RECT 145.000 250.800 145.800 255.200 ;
        RECT 146.800 254.600 147.600 259.800 ;
        RECT 153.200 256.600 154.000 259.800 ;
        RECT 154.800 257.000 155.600 259.800 ;
        RECT 156.400 257.000 157.200 259.800 ;
        RECT 158.000 257.000 158.800 259.800 ;
        RECT 159.600 257.000 160.400 259.800 ;
        RECT 162.800 257.000 163.600 259.800 ;
        RECT 166.000 257.000 166.800 259.800 ;
        RECT 167.600 257.000 168.400 259.800 ;
        RECT 169.200 257.000 170.000 259.800 ;
        RECT 151.600 255.800 154.000 256.600 ;
        RECT 170.800 256.600 171.600 259.800 ;
        RECT 151.600 255.200 152.400 255.800 ;
        RECT 146.400 254.000 147.600 254.600 ;
        RECT 150.600 254.600 152.400 255.200 ;
        RECT 156.400 255.600 157.400 256.400 ;
        RECT 160.400 255.600 162.000 256.400 ;
        RECT 162.800 255.800 167.400 256.400 ;
        RECT 170.800 255.800 173.400 256.600 ;
        RECT 162.800 255.600 163.600 255.800 ;
        RECT 146.400 252.000 147.000 254.000 ;
        RECT 150.600 253.400 151.400 254.600 ;
        RECT 147.600 252.600 151.400 253.400 ;
        RECT 156.400 252.800 157.200 255.600 ;
        RECT 162.800 254.800 163.600 255.000 ;
        RECT 159.200 254.200 163.600 254.800 ;
        RECT 159.200 254.000 160.000 254.200 ;
        RECT 164.400 253.600 165.200 255.200 ;
        RECT 166.600 253.400 167.400 255.800 ;
        RECT 172.600 255.200 173.400 255.800 ;
        RECT 172.600 254.400 175.600 255.200 ;
        RECT 177.200 253.800 178.000 259.800 ;
        RECT 181.400 256.400 182.200 259.800 ;
        RECT 180.400 255.800 182.200 256.400 ;
        RECT 183.600 255.800 184.400 259.800 ;
        RECT 185.200 256.000 186.000 259.800 ;
        RECT 188.400 256.000 189.200 259.800 ;
        RECT 185.200 255.800 189.200 256.000 ;
        RECT 159.600 252.600 162.800 253.400 ;
        RECT 166.600 252.600 168.600 253.400 ;
        RECT 169.200 253.000 178.000 253.800 ;
        RECT 178.800 253.600 179.600 255.200 ;
        RECT 153.200 252.000 154.000 252.600 ;
        RECT 170.800 252.000 171.600 252.400 ;
        RECT 174.000 252.000 174.800 252.400 ;
        RECT 175.800 252.000 176.600 252.200 ;
        RECT 146.400 251.400 147.200 252.000 ;
        RECT 153.200 251.400 176.600 252.000 ;
        RECT 133.800 249.200 134.800 250.200 ;
        RECT 135.400 249.600 138.000 250.200 ;
        RECT 145.000 250.000 146.000 250.800 ;
        RECT 134.000 242.200 134.800 249.200 ;
        RECT 137.200 242.200 138.000 249.600 ;
        RECT 145.200 242.200 146.000 250.000 ;
        RECT 146.600 249.600 147.200 251.400 ;
        RECT 146.600 249.000 155.600 249.600 ;
        RECT 146.600 247.400 147.200 249.000 ;
        RECT 154.800 248.800 155.600 249.000 ;
        RECT 158.000 249.000 166.600 249.600 ;
        RECT 158.000 248.800 158.800 249.000 ;
        RECT 149.800 247.600 152.400 248.400 ;
        RECT 146.600 246.800 149.200 247.400 ;
        RECT 148.400 242.200 149.200 246.800 ;
        RECT 151.600 242.200 152.400 247.600 ;
        RECT 153.000 246.800 157.200 247.600 ;
        RECT 154.800 242.200 155.600 245.000 ;
        RECT 156.400 242.200 157.200 245.000 ;
        RECT 158.000 242.200 158.800 245.000 ;
        RECT 159.600 242.200 160.400 248.400 ;
        RECT 162.800 247.600 165.400 248.400 ;
        RECT 166.000 248.200 166.600 249.000 ;
        RECT 167.600 249.400 168.400 249.600 ;
        RECT 167.600 249.000 173.000 249.400 ;
        RECT 167.600 248.800 173.800 249.000 ;
        RECT 172.400 248.200 173.800 248.800 ;
        RECT 166.000 247.600 171.800 248.200 ;
        RECT 174.800 248.000 176.400 248.800 ;
        RECT 174.800 247.600 175.400 248.000 ;
        RECT 162.800 242.200 163.600 247.000 ;
        RECT 166.000 242.200 166.800 247.000 ;
        RECT 171.200 246.800 175.400 247.600 ;
        RECT 177.200 247.400 178.000 253.000 ;
        RECT 176.000 246.800 178.000 247.400 ;
        RECT 180.400 252.300 181.200 255.800 ;
        RECT 183.800 254.400 184.400 255.800 ;
        RECT 185.400 255.400 189.000 255.800 ;
        RECT 187.600 254.400 188.400 254.800 ;
        RECT 182.000 254.300 182.800 254.400 ;
        RECT 183.600 254.300 186.200 254.400 ;
        RECT 182.000 253.700 186.200 254.300 ;
        RECT 187.600 254.300 189.200 254.400 ;
        RECT 191.600 254.300 192.400 259.800 ;
        RECT 187.600 253.800 192.400 254.300 ;
        RECT 182.000 253.600 182.800 253.700 ;
        RECT 183.600 253.600 186.200 253.700 ;
        RECT 188.400 253.700 192.400 253.800 ;
        RECT 188.400 253.600 189.200 253.700 ;
        RECT 180.400 251.700 184.300 252.300 ;
        RECT 167.600 242.200 168.400 245.000 ;
        RECT 169.200 242.200 170.000 245.000 ;
        RECT 172.400 242.200 173.200 246.800 ;
        RECT 176.000 246.200 176.600 246.800 ;
        RECT 175.600 245.600 176.600 246.200 ;
        RECT 175.600 242.200 176.400 245.600 ;
        RECT 180.400 242.200 181.200 251.700 ;
        RECT 183.700 250.400 184.300 251.700 ;
        RECT 182.000 248.800 182.800 250.400 ;
        RECT 183.600 250.200 184.400 250.400 ;
        RECT 185.600 250.200 186.200 253.600 ;
        RECT 186.800 251.600 187.600 253.200 ;
        RECT 183.600 249.600 185.000 250.200 ;
        RECT 185.600 249.600 186.600 250.200 ;
        RECT 184.400 248.400 185.000 249.600 ;
        RECT 184.400 247.600 185.200 248.400 ;
        RECT 185.800 242.200 186.600 249.600 ;
        RECT 191.600 242.200 192.400 253.700 ;
        RECT 193.200 253.600 194.000 255.200 ;
        RECT 194.800 253.800 195.600 259.800 ;
        RECT 201.200 256.600 202.000 259.800 ;
        RECT 202.800 257.000 203.600 259.800 ;
        RECT 204.400 257.000 205.200 259.800 ;
        RECT 206.000 257.000 206.800 259.800 ;
        RECT 209.200 257.000 210.000 259.800 ;
        RECT 212.400 257.000 213.200 259.800 ;
        RECT 214.000 257.000 214.800 259.800 ;
        RECT 215.600 257.000 216.400 259.800 ;
        RECT 217.200 257.000 218.000 259.800 ;
        RECT 199.400 255.800 202.000 256.600 ;
        RECT 218.800 256.600 219.600 259.800 ;
        RECT 205.400 255.800 210.000 256.400 ;
        RECT 199.400 255.200 200.200 255.800 ;
        RECT 197.200 254.400 200.200 255.200 ;
        RECT 194.800 253.000 203.600 253.800 ;
        RECT 205.400 253.400 206.200 255.800 ;
        RECT 209.200 255.600 210.000 255.800 ;
        RECT 210.800 255.600 212.400 256.400 ;
        RECT 215.400 255.600 216.400 256.400 ;
        RECT 218.800 255.800 221.200 256.600 ;
        RECT 207.600 253.600 208.400 255.200 ;
        RECT 209.200 254.800 210.000 255.000 ;
        RECT 209.200 254.200 213.600 254.800 ;
        RECT 212.800 254.000 213.600 254.200 ;
        RECT 194.800 247.400 195.600 253.000 ;
        RECT 204.200 252.600 206.200 253.400 ;
        RECT 210.000 252.600 213.200 253.400 ;
        RECT 215.600 252.800 216.400 255.600 ;
        RECT 220.400 255.200 221.200 255.800 ;
        RECT 220.400 254.600 222.200 255.200 ;
        RECT 221.400 253.400 222.200 254.600 ;
        RECT 225.200 254.600 226.000 259.800 ;
        RECT 226.800 256.300 227.600 259.800 ;
        RECT 230.000 256.300 230.800 257.200 ;
        RECT 226.800 255.700 230.800 256.300 ;
        RECT 226.800 255.200 227.800 255.700 ;
        RECT 230.000 255.600 230.800 255.700 ;
        RECT 225.200 254.000 226.400 254.600 ;
        RECT 221.400 252.600 225.200 253.400 ;
        RECT 196.200 252.000 197.000 252.200 ;
        RECT 199.600 252.000 200.400 252.400 ;
        RECT 201.200 252.000 202.000 252.400 ;
        RECT 218.800 252.000 219.600 252.600 ;
        RECT 225.800 252.000 226.400 254.000 ;
        RECT 196.200 251.400 219.600 252.000 ;
        RECT 225.600 251.400 226.400 252.000 ;
        RECT 225.600 249.600 226.200 251.400 ;
        RECT 227.000 250.800 227.800 255.200 ;
        RECT 204.400 249.400 205.200 249.600 ;
        RECT 199.800 249.000 205.200 249.400 ;
        RECT 199.000 248.800 205.200 249.000 ;
        RECT 206.200 249.000 214.800 249.600 ;
        RECT 196.400 248.000 198.000 248.800 ;
        RECT 199.000 248.200 200.400 248.800 ;
        RECT 206.200 248.200 206.800 249.000 ;
        RECT 214.000 248.800 214.800 249.000 ;
        RECT 217.200 249.000 226.200 249.600 ;
        RECT 217.200 248.800 218.000 249.000 ;
        RECT 197.400 247.600 198.000 248.000 ;
        RECT 201.000 247.600 206.800 248.200 ;
        RECT 207.400 247.600 210.000 248.400 ;
        RECT 194.800 246.800 196.800 247.400 ;
        RECT 197.400 246.800 201.600 247.600 ;
        RECT 196.200 246.200 196.800 246.800 ;
        RECT 196.200 245.600 197.200 246.200 ;
        RECT 196.400 242.200 197.200 245.600 ;
        RECT 199.600 242.200 200.400 246.800 ;
        RECT 202.800 242.200 203.600 245.000 ;
        RECT 204.400 242.200 205.200 245.000 ;
        RECT 206.000 242.200 206.800 247.000 ;
        RECT 209.200 242.200 210.000 247.000 ;
        RECT 212.400 242.200 213.200 248.400 ;
        RECT 220.400 247.600 223.000 248.400 ;
        RECT 215.600 246.800 219.800 247.600 ;
        RECT 214.000 242.200 214.800 245.000 ;
        RECT 215.600 242.200 216.400 245.000 ;
        RECT 217.200 242.200 218.000 245.000 ;
        RECT 220.400 242.200 221.200 247.600 ;
        RECT 225.600 247.400 226.200 249.000 ;
        RECT 223.600 246.800 226.200 247.400 ;
        RECT 226.800 250.000 227.800 250.800 ;
        RECT 231.600 252.300 232.400 259.800 ;
        RECT 237.000 256.000 237.800 259.000 ;
        RECT 241.200 257.000 242.000 259.000 ;
        RECT 236.200 255.400 237.800 256.000 ;
        RECT 236.200 255.000 237.000 255.400 ;
        RECT 236.200 254.400 236.800 255.000 ;
        RECT 241.400 254.800 242.000 257.000 ;
        RECT 244.400 256.400 245.200 259.800 ;
        RECT 233.200 254.300 234.000 254.400 ;
        RECT 234.800 254.300 236.800 254.400 ;
        RECT 233.200 253.700 236.800 254.300 ;
        RECT 237.800 254.200 242.000 254.800 ;
        RECT 244.200 255.800 245.200 256.400 ;
        RECT 244.200 254.400 244.800 255.800 ;
        RECT 247.600 255.200 248.400 259.800 ;
        RECT 250.800 256.000 251.600 259.800 ;
        RECT 245.800 254.600 248.400 255.200 ;
        RECT 250.600 255.200 251.600 256.000 ;
        RECT 237.800 253.800 238.800 254.200 ;
        RECT 233.200 253.600 234.000 253.700 ;
        RECT 234.800 253.600 236.800 253.700 ;
        RECT 234.800 252.300 235.600 252.400 ;
        RECT 231.600 251.700 235.600 252.300 ;
        RECT 223.600 242.200 224.400 246.800 ;
        RECT 226.800 242.200 227.600 250.000 ;
        RECT 231.600 242.200 232.400 251.700 ;
        RECT 234.800 250.800 235.600 251.700 ;
        RECT 236.200 249.800 236.800 253.600 ;
        RECT 237.400 253.000 238.800 253.800 ;
        RECT 244.200 253.600 245.200 254.400 ;
        RECT 238.200 251.000 238.800 253.000 ;
        RECT 239.600 251.600 240.400 253.200 ;
        RECT 241.200 252.300 242.000 253.200 ;
        RECT 242.800 252.300 243.600 252.400 ;
        RECT 241.200 251.700 243.600 252.300 ;
        RECT 241.200 251.600 242.000 251.700 ;
        RECT 242.800 251.600 243.600 251.700 ;
        RECT 238.200 250.400 242.000 251.000 ;
        RECT 236.200 249.200 237.800 249.800 ;
        RECT 237.000 242.200 237.800 249.200 ;
        RECT 241.400 247.000 242.000 250.400 ;
        RECT 244.200 250.200 244.800 253.600 ;
        RECT 245.800 253.000 246.400 254.600 ;
        RECT 245.400 252.200 246.400 253.000 ;
        RECT 245.800 250.200 246.400 252.200 ;
        RECT 247.400 252.400 248.200 253.200 ;
        RECT 247.400 251.600 248.400 252.400 ;
        RECT 250.600 250.800 251.400 255.200 ;
        RECT 252.400 254.600 253.200 259.800 ;
        RECT 258.800 256.600 259.600 259.800 ;
        RECT 260.400 257.000 261.200 259.800 ;
        RECT 262.000 257.000 262.800 259.800 ;
        RECT 263.600 257.000 264.400 259.800 ;
        RECT 265.200 257.000 266.000 259.800 ;
        RECT 268.400 257.000 269.200 259.800 ;
        RECT 271.600 257.000 272.400 259.800 ;
        RECT 273.200 257.000 274.000 259.800 ;
        RECT 274.800 257.000 275.600 259.800 ;
        RECT 257.200 255.800 259.600 256.600 ;
        RECT 276.400 256.600 277.200 259.800 ;
        RECT 257.200 255.200 258.000 255.800 ;
        RECT 252.000 254.000 253.200 254.600 ;
        RECT 256.200 254.600 258.000 255.200 ;
        RECT 262.000 255.600 263.000 256.400 ;
        RECT 266.000 255.600 267.600 256.400 ;
        RECT 268.400 255.800 273.000 256.400 ;
        RECT 276.400 255.800 279.000 256.600 ;
        RECT 268.400 255.600 269.200 255.800 ;
        RECT 252.000 252.000 252.600 254.000 ;
        RECT 256.200 253.400 257.000 254.600 ;
        RECT 253.200 252.600 257.000 253.400 ;
        RECT 262.000 252.800 262.800 255.600 ;
        RECT 268.400 254.800 269.200 255.000 ;
        RECT 264.800 254.200 269.200 254.800 ;
        RECT 264.800 254.000 265.600 254.200 ;
        RECT 270.000 253.600 270.800 255.200 ;
        RECT 272.200 253.400 273.000 255.800 ;
        RECT 278.200 255.200 279.000 255.800 ;
        RECT 278.200 254.400 281.200 255.200 ;
        RECT 282.800 253.800 283.600 259.800 ;
        RECT 284.400 259.200 288.400 259.800 ;
        RECT 284.400 255.800 285.200 259.200 ;
        RECT 286.000 255.800 286.800 258.600 ;
        RECT 287.600 256.000 288.400 259.200 ;
        RECT 290.800 256.000 291.600 259.800 ;
        RECT 287.600 255.800 291.600 256.000 ;
        RECT 292.400 255.800 293.200 259.800 ;
        RECT 294.000 256.000 294.800 259.800 ;
        RECT 297.200 256.000 298.000 259.800 ;
        RECT 301.400 258.400 302.200 259.800 ;
        RECT 300.400 257.600 302.200 258.400 ;
        RECT 310.000 257.800 310.800 259.800 ;
        RECT 301.400 256.400 302.200 257.600 ;
        RECT 294.000 255.800 298.000 256.000 ;
        RECT 300.400 255.800 302.200 256.400 ;
        RECT 286.000 254.400 286.600 255.800 ;
        RECT 287.800 255.400 291.400 255.800 ;
        RECT 290.000 254.400 290.800 254.800 ;
        RECT 292.600 254.400 293.200 255.800 ;
        RECT 294.200 255.400 297.800 255.800 ;
        RECT 296.400 254.400 297.200 254.800 ;
        RECT 265.200 252.600 268.400 253.400 ;
        RECT 272.200 252.600 274.200 253.400 ;
        RECT 274.800 253.000 283.600 253.800 ;
        RECT 258.800 252.000 259.600 252.600 ;
        RECT 276.400 252.000 277.200 252.400 ;
        RECT 281.400 252.000 282.200 252.200 ;
        RECT 252.000 251.400 252.800 252.000 ;
        RECT 258.800 251.400 282.200 252.000 ;
        RECT 244.200 249.200 245.200 250.200 ;
        RECT 245.800 249.600 248.400 250.200 ;
        RECT 250.600 250.000 251.600 250.800 ;
        RECT 241.200 243.000 242.000 247.000 ;
        RECT 244.400 242.200 245.200 249.200 ;
        RECT 247.600 242.200 248.400 249.600 ;
        RECT 250.800 242.200 251.600 250.000 ;
        RECT 252.200 249.600 252.800 251.400 ;
        RECT 252.200 249.000 261.200 249.600 ;
        RECT 252.200 247.400 252.800 249.000 ;
        RECT 260.400 248.800 261.200 249.000 ;
        RECT 263.600 249.000 272.200 249.600 ;
        RECT 263.600 248.800 264.400 249.000 ;
        RECT 255.400 247.600 258.000 248.400 ;
        RECT 252.200 246.800 254.800 247.400 ;
        RECT 254.000 242.200 254.800 246.800 ;
        RECT 257.200 242.200 258.000 247.600 ;
        RECT 258.600 246.800 262.800 247.600 ;
        RECT 260.400 242.200 261.200 245.000 ;
        RECT 262.000 242.200 262.800 245.000 ;
        RECT 263.600 242.200 264.400 245.000 ;
        RECT 265.200 242.200 266.000 248.400 ;
        RECT 268.400 247.600 271.000 248.400 ;
        RECT 271.600 248.200 272.200 249.000 ;
        RECT 273.200 249.400 274.000 249.600 ;
        RECT 273.200 249.000 278.600 249.400 ;
        RECT 273.200 248.800 279.400 249.000 ;
        RECT 278.000 248.200 279.400 248.800 ;
        RECT 271.600 247.600 277.400 248.200 ;
        RECT 280.400 248.000 282.000 248.800 ;
        RECT 280.400 247.600 281.000 248.000 ;
        RECT 268.400 242.200 269.200 247.000 ;
        RECT 271.600 242.200 272.400 247.000 ;
        RECT 276.800 246.800 281.000 247.600 ;
        RECT 282.800 247.400 283.600 253.000 ;
        RECT 284.400 252.800 285.200 254.400 ;
        RECT 286.000 253.800 288.400 254.400 ;
        RECT 290.000 253.800 291.600 254.400 ;
        RECT 287.600 253.600 288.400 253.800 ;
        RECT 290.800 253.600 291.600 253.800 ;
        RECT 292.400 253.600 295.000 254.400 ;
        RECT 296.400 253.800 298.000 254.400 ;
        RECT 297.200 253.600 298.000 253.800 ;
        RECT 298.800 253.600 299.600 255.200 ;
        RECT 286.000 251.600 286.800 253.200 ;
        RECT 287.800 250.200 288.400 253.600 ;
        RECT 289.200 252.300 290.000 253.200 ;
        RECT 294.400 252.300 295.000 253.600 ;
        RECT 289.200 251.700 295.000 252.300 ;
        RECT 289.200 251.600 290.000 251.700 ;
        RECT 292.400 250.200 293.200 250.400 ;
        RECT 294.400 250.200 295.000 251.700 ;
        RECT 281.600 246.800 283.600 247.400 ;
        RECT 273.200 242.200 274.000 245.000 ;
        RECT 274.800 242.200 275.600 245.000 ;
        RECT 278.000 242.200 278.800 246.800 ;
        RECT 281.600 246.200 282.200 246.800 ;
        RECT 281.200 245.600 282.200 246.200 ;
        RECT 281.200 242.200 282.000 245.600 ;
        RECT 287.000 242.200 289.000 250.200 ;
        RECT 292.400 249.600 293.800 250.200 ;
        RECT 294.400 249.600 295.400 250.200 ;
        RECT 293.200 248.400 293.800 249.600 ;
        RECT 293.200 247.600 294.000 248.400 ;
        RECT 294.600 242.200 295.400 249.600 ;
        RECT 300.400 242.200 301.200 255.800 ;
        RECT 308.400 255.600 309.200 257.200 ;
        RECT 310.200 255.600 310.800 257.800 ;
        RECT 313.200 255.600 314.000 259.800 ;
        RECT 316.400 256.400 317.200 259.800 ;
        RECT 310.200 255.000 312.600 255.600 ;
        RECT 312.000 252.000 312.600 255.000 ;
        RECT 313.400 252.400 314.000 255.600 ;
        RECT 316.200 255.800 317.200 256.400 ;
        RECT 316.200 254.400 316.800 255.800 ;
        RECT 319.600 255.200 320.400 259.800 ;
        RECT 321.200 255.800 322.000 259.800 ;
        RECT 322.800 256.000 323.600 259.800 ;
        RECT 326.000 256.000 326.800 259.800 ;
        RECT 322.800 255.800 326.800 256.000 ;
        RECT 327.600 259.200 331.600 259.800 ;
        RECT 327.600 255.800 328.400 259.200 ;
        RECT 329.200 255.800 330.000 258.600 ;
        RECT 330.800 256.000 331.600 259.200 ;
        RECT 334.000 256.000 334.800 259.800 ;
        RECT 330.800 255.800 334.800 256.000 ;
        RECT 336.200 256.400 337.000 259.800 ;
        RECT 336.200 255.800 338.000 256.400 ;
        RECT 317.800 254.600 320.400 255.200 ;
        RECT 314.800 254.300 315.600 254.400 ;
        RECT 316.200 254.300 317.200 254.400 ;
        RECT 314.800 253.700 317.200 254.300 ;
        RECT 314.800 253.600 315.600 253.700 ;
        RECT 316.200 253.600 317.200 253.700 ;
        RECT 311.800 251.400 312.600 252.000 ;
        RECT 313.200 251.600 314.000 252.400 ;
        RECT 308.400 251.200 312.600 251.400 ;
        RECT 308.400 250.800 312.400 251.200 ;
        RECT 302.000 248.800 302.800 250.400 ;
        RECT 308.400 242.200 309.200 250.800 ;
        RECT 313.400 250.200 314.000 251.600 ;
        RECT 312.600 249.600 314.000 250.200 ;
        RECT 316.200 250.200 316.800 253.600 ;
        RECT 317.800 253.000 318.400 254.600 ;
        RECT 321.400 254.400 322.000 255.800 ;
        RECT 323.000 255.400 326.600 255.800 ;
        RECT 329.200 254.400 329.800 255.800 ;
        RECT 331.000 255.400 334.600 255.800 ;
        RECT 333.200 254.400 334.000 254.800 ;
        RECT 321.200 253.600 323.800 254.400 ;
        RECT 317.400 252.200 318.400 253.000 ;
        RECT 317.800 250.200 318.400 252.200 ;
        RECT 319.400 252.400 320.200 253.200 ;
        RECT 319.400 251.600 320.400 252.400 ;
        RECT 321.200 250.200 322.000 250.400 ;
        RECT 323.200 250.200 323.800 253.600 ;
        RECT 324.400 251.600 325.200 253.200 ;
        RECT 327.600 252.800 328.400 254.400 ;
        RECT 329.200 253.800 331.600 254.400 ;
        RECT 333.200 253.800 334.800 254.400 ;
        RECT 330.800 253.600 331.600 253.800 ;
        RECT 334.000 253.600 334.800 253.800 ;
        RECT 329.200 251.600 330.000 253.200 ;
        RECT 331.000 250.200 331.600 253.600 ;
        RECT 332.400 252.300 333.200 253.200 ;
        RECT 337.200 252.300 338.000 255.800 ;
        RECT 338.800 253.600 339.600 255.200 ;
        RECT 344.000 254.200 344.800 259.800 ;
        RECT 346.800 255.200 347.600 259.800 ;
        RECT 346.800 254.600 349.000 255.200 ;
        RECT 344.000 253.800 345.800 254.200 ;
        RECT 344.200 253.600 345.800 253.800 ;
        RECT 332.400 251.700 338.000 252.300 ;
        RECT 332.400 251.600 333.200 251.700 ;
        RECT 312.600 244.400 313.400 249.600 ;
        RECT 316.200 249.200 317.200 250.200 ;
        RECT 317.800 249.600 320.400 250.200 ;
        RECT 321.200 249.600 322.600 250.200 ;
        RECT 323.200 249.600 324.200 250.200 ;
        RECT 312.600 243.600 314.000 244.400 ;
        RECT 312.600 242.200 313.400 243.600 ;
        RECT 316.400 242.200 317.200 249.200 ;
        RECT 319.600 242.200 320.400 249.600 ;
        RECT 322.000 248.400 322.600 249.600 ;
        RECT 323.400 248.400 324.200 249.600 ;
        RECT 322.000 247.600 322.800 248.400 ;
        RECT 323.400 247.600 325.200 248.400 ;
        RECT 323.400 242.200 324.200 247.600 ;
        RECT 330.200 244.400 332.200 250.200 ;
        RECT 335.600 248.800 336.400 250.400 ;
        RECT 329.200 243.600 332.200 244.400 ;
        RECT 330.200 242.200 332.200 243.600 ;
        RECT 337.200 242.200 338.000 251.700 ;
        RECT 342.000 251.600 343.600 252.400 ;
        RECT 345.200 250.400 345.800 253.600 ;
        RECT 346.800 251.600 347.600 253.200 ;
        RECT 348.400 251.600 349.000 254.600 ;
        RECT 350.000 252.400 350.800 259.800 ;
        RECT 348.400 250.800 349.600 251.600 ;
        RECT 345.200 249.600 346.000 250.400 ;
        RECT 348.400 250.200 349.000 250.800 ;
        RECT 350.200 250.200 350.800 252.400 ;
        RECT 346.800 249.600 349.000 250.200 ;
        RECT 343.600 247.600 344.400 249.200 ;
        RECT 345.200 247.000 345.800 249.600 ;
        RECT 342.200 246.400 345.800 247.000 ;
        RECT 342.200 246.200 342.800 246.400 ;
        RECT 342.000 242.200 342.800 246.200 ;
        RECT 345.200 246.200 345.800 246.400 ;
        RECT 345.200 242.200 346.000 246.200 ;
        RECT 346.800 242.200 347.600 249.600 ;
        RECT 350.000 242.200 350.800 250.200 ;
        RECT 351.600 253.800 352.400 259.800 ;
        RECT 358.000 256.600 358.800 259.800 ;
        RECT 359.600 257.000 360.400 259.800 ;
        RECT 361.200 257.000 362.000 259.800 ;
        RECT 362.800 257.000 363.600 259.800 ;
        RECT 366.000 257.000 366.800 259.800 ;
        RECT 369.200 257.000 370.000 259.800 ;
        RECT 370.800 257.000 371.600 259.800 ;
        RECT 372.400 257.000 373.200 259.800 ;
        RECT 374.000 257.000 374.800 259.800 ;
        RECT 356.200 255.800 358.800 256.600 ;
        RECT 375.600 256.600 376.400 259.800 ;
        RECT 362.200 255.800 366.800 256.400 ;
        RECT 356.200 255.200 357.000 255.800 ;
        RECT 354.000 254.400 357.000 255.200 ;
        RECT 351.600 253.000 360.400 253.800 ;
        RECT 362.200 253.400 363.000 255.800 ;
        RECT 366.000 255.600 366.800 255.800 ;
        RECT 367.600 255.600 369.200 256.400 ;
        RECT 372.200 255.600 373.200 256.400 ;
        RECT 375.600 255.800 378.000 256.600 ;
        RECT 364.400 253.600 365.200 255.200 ;
        RECT 366.000 254.800 366.800 255.000 ;
        RECT 366.000 254.200 370.400 254.800 ;
        RECT 369.600 254.000 370.400 254.200 ;
        RECT 351.600 247.400 352.400 253.000 ;
        RECT 361.000 252.600 363.000 253.400 ;
        RECT 366.800 252.600 370.000 253.400 ;
        RECT 372.400 252.800 373.200 255.600 ;
        RECT 377.200 255.200 378.000 255.800 ;
        RECT 377.200 254.600 379.000 255.200 ;
        RECT 378.200 253.400 379.000 254.600 ;
        RECT 382.000 254.600 382.800 259.800 ;
        RECT 383.600 256.000 384.400 259.800 ;
        RECT 383.600 255.200 384.600 256.000 ;
        RECT 382.000 254.000 383.200 254.600 ;
        RECT 378.200 252.600 382.000 253.400 ;
        RECT 353.000 252.000 353.800 252.200 ;
        RECT 356.400 252.000 357.200 252.400 ;
        RECT 358.000 252.000 358.800 252.400 ;
        RECT 375.600 252.000 376.400 252.600 ;
        RECT 382.600 252.000 383.200 254.000 ;
        RECT 353.000 251.400 376.400 252.000 ;
        RECT 382.400 251.400 383.200 252.000 ;
        RECT 382.400 249.600 383.000 251.400 ;
        RECT 383.800 250.800 384.600 255.200 ;
        RECT 361.200 249.400 362.000 249.600 ;
        RECT 356.600 249.000 362.000 249.400 ;
        RECT 355.800 248.800 362.000 249.000 ;
        RECT 363.000 249.000 371.600 249.600 ;
        RECT 353.200 248.000 354.800 248.800 ;
        RECT 355.800 248.200 357.200 248.800 ;
        RECT 363.000 248.200 363.600 249.000 ;
        RECT 370.800 248.800 371.600 249.000 ;
        RECT 374.000 249.000 383.000 249.600 ;
        RECT 374.000 248.800 374.800 249.000 ;
        RECT 354.200 247.600 354.800 248.000 ;
        RECT 357.800 247.600 363.600 248.200 ;
        RECT 364.200 247.600 366.800 248.400 ;
        RECT 351.600 246.800 353.600 247.400 ;
        RECT 354.200 246.800 358.400 247.600 ;
        RECT 353.000 246.200 353.600 246.800 ;
        RECT 353.000 245.600 354.000 246.200 ;
        RECT 353.200 242.200 354.000 245.600 ;
        RECT 356.400 242.200 357.200 246.800 ;
        RECT 359.600 242.200 360.400 245.000 ;
        RECT 361.200 242.200 362.000 245.000 ;
        RECT 362.800 242.200 363.600 247.000 ;
        RECT 366.000 242.200 366.800 247.000 ;
        RECT 369.200 242.200 370.000 248.400 ;
        RECT 377.200 247.600 379.800 248.400 ;
        RECT 372.400 246.800 376.600 247.600 ;
        RECT 370.800 242.200 371.600 245.000 ;
        RECT 372.400 242.200 373.200 245.000 ;
        RECT 374.000 242.200 374.800 245.000 ;
        RECT 377.200 242.200 378.000 247.600 ;
        RECT 382.400 247.400 383.000 249.000 ;
        RECT 380.400 246.800 383.000 247.400 ;
        RECT 383.600 250.000 384.600 250.800 ;
        RECT 380.400 242.200 381.200 246.800 ;
        RECT 383.600 242.200 384.400 250.000 ;
        RECT 386.800 242.200 387.600 259.800 ;
        RECT 388.400 255.600 389.200 257.200 ;
        RECT 393.600 254.200 394.400 259.800 ;
        RECT 399.000 258.400 400.600 259.800 ;
        RECT 398.000 257.600 400.600 258.400 ;
        RECT 399.000 255.800 400.600 257.600 ;
        RECT 407.000 255.800 408.600 259.800 ;
        RECT 415.000 256.400 415.800 259.800 ;
        RECT 414.000 255.800 415.800 256.400 ;
        RECT 393.600 253.800 395.400 254.200 ;
        RECT 393.800 253.600 395.400 253.800 ;
        RECT 398.000 253.600 398.800 254.400 ;
        RECT 391.600 251.600 393.200 252.400 ;
        RECT 394.800 250.400 395.400 253.600 ;
        RECT 398.200 253.200 398.800 253.600 ;
        RECT 398.200 252.400 399.000 253.200 ;
        RECT 399.600 252.400 400.200 255.800 ;
        RECT 401.200 254.300 402.000 254.400 ;
        RECT 404.400 254.300 405.200 254.400 ;
        RECT 401.200 253.700 405.200 254.300 ;
        RECT 401.200 252.800 402.000 253.700 ;
        RECT 404.400 253.600 405.200 253.700 ;
        RECT 406.000 253.600 406.800 254.400 ;
        RECT 406.200 253.200 406.800 253.600 ;
        RECT 406.200 252.400 407.000 253.200 ;
        RECT 407.600 252.400 408.200 255.800 ;
        RECT 409.200 252.800 410.000 254.400 ;
        RECT 412.400 253.600 413.200 255.200 ;
        RECT 396.400 250.800 397.200 252.400 ;
        RECT 399.600 251.600 400.400 252.400 ;
        RECT 402.800 252.200 403.600 252.400 ;
        RECT 402.000 251.600 403.600 252.200 ;
        RECT 399.600 251.400 400.200 251.600 ;
        RECT 398.200 250.800 400.200 251.400 ;
        RECT 402.000 251.200 402.800 251.600 ;
        RECT 404.400 250.800 405.200 252.400 ;
        RECT 407.600 251.600 408.400 252.400 ;
        RECT 410.800 252.200 411.600 252.400 ;
        RECT 410.000 251.600 411.600 252.200 ;
        RECT 407.600 251.400 408.200 251.600 ;
        RECT 406.200 250.800 408.200 251.400 ;
        RECT 410.000 251.200 410.800 251.600 ;
        RECT 394.800 249.600 395.600 250.400 ;
        RECT 398.200 250.200 398.800 250.800 ;
        RECT 406.200 250.200 406.800 250.800 ;
        RECT 393.200 247.600 394.000 249.200 ;
        RECT 394.800 247.000 395.400 249.600 ;
        RECT 391.800 246.400 395.400 247.000 ;
        RECT 391.600 242.200 392.400 246.400 ;
        RECT 394.800 246.200 395.400 246.400 ;
        RECT 394.800 242.200 395.600 246.200 ;
        RECT 396.400 242.800 397.200 250.200 ;
        RECT 398.000 243.400 398.800 250.200 ;
        RECT 399.600 249.600 403.600 250.200 ;
        RECT 399.600 242.800 400.400 249.600 ;
        RECT 396.400 242.200 400.400 242.800 ;
        RECT 402.800 242.200 403.600 249.600 ;
        RECT 404.400 242.800 405.200 250.200 ;
        RECT 406.000 243.400 406.800 250.200 ;
        RECT 407.600 249.600 411.600 250.200 ;
        RECT 407.600 242.800 408.400 249.600 ;
        RECT 404.400 242.200 408.400 242.800 ;
        RECT 410.800 242.200 411.600 249.600 ;
        RECT 414.000 242.200 414.800 255.800 ;
        RECT 420.800 254.200 421.600 259.800 ;
        RECT 424.200 256.400 425.000 259.800 ;
        RECT 431.400 258.400 433.000 259.800 ;
        RECT 431.400 257.600 434.000 258.400 ;
        RECT 423.600 255.600 426.000 256.400 ;
        RECT 431.400 255.800 433.000 257.600 ;
        RECT 439.000 256.400 439.800 259.800 ;
        RECT 438.000 255.800 439.800 256.400 ;
        RECT 441.800 256.400 442.600 259.800 ;
        RECT 441.800 255.800 443.600 256.400 ;
        RECT 420.800 253.800 422.600 254.200 ;
        RECT 421.000 253.600 422.600 253.800 ;
        RECT 418.800 251.600 420.400 252.400 ;
        RECT 422.000 252.300 422.600 253.600 ;
        RECT 423.600 252.300 424.400 252.400 ;
        RECT 422.000 251.700 424.400 252.300 ;
        RECT 415.600 248.800 416.400 250.400 ;
        RECT 417.200 249.600 418.000 251.200 ;
        RECT 422.000 250.400 422.600 251.700 ;
        RECT 423.600 251.600 424.400 251.700 ;
        RECT 422.000 249.600 422.800 250.400 ;
        RECT 420.400 247.600 421.200 249.200 ;
        RECT 422.000 247.000 422.600 249.600 ;
        RECT 423.600 248.800 424.400 250.400 ;
        RECT 419.000 246.400 422.600 247.000 ;
        RECT 419.000 246.200 419.600 246.400 ;
        RECT 418.800 242.200 419.600 246.200 ;
        RECT 422.000 246.200 422.600 246.400 ;
        RECT 422.000 242.200 422.800 246.200 ;
        RECT 425.200 242.200 426.000 255.600 ;
        RECT 426.800 253.600 427.600 255.200 ;
        RECT 430.000 252.800 430.800 254.400 ;
        RECT 431.800 252.400 432.400 255.800 ;
        RECT 433.200 253.600 434.000 254.400 ;
        RECT 436.400 253.600 437.200 255.200 ;
        RECT 438.000 254.300 438.800 255.800 ;
        RECT 439.600 254.300 440.400 254.400 ;
        RECT 438.000 253.700 440.400 254.300 ;
        RECT 433.200 253.200 433.800 253.600 ;
        RECT 433.000 252.400 433.800 253.200 ;
        RECT 428.400 252.200 429.200 252.400 ;
        RECT 428.400 251.600 430.000 252.200 ;
        RECT 431.600 251.600 432.400 252.400 ;
        RECT 429.200 251.200 430.000 251.600 ;
        RECT 431.800 251.400 432.400 251.600 ;
        RECT 431.800 250.800 433.800 251.400 ;
        RECT 434.800 250.800 435.600 252.400 ;
        RECT 433.200 250.200 433.800 250.800 ;
        RECT 428.400 249.600 432.400 250.200 ;
        RECT 428.400 242.200 429.200 249.600 ;
        RECT 431.600 242.800 432.400 249.600 ;
        RECT 433.200 243.400 434.000 250.200 ;
        RECT 434.800 242.800 435.600 250.200 ;
        RECT 431.600 242.200 435.600 242.800 ;
        RECT 438.000 242.200 438.800 253.700 ;
        RECT 439.600 253.600 440.400 253.700 ;
        RECT 439.600 248.800 440.400 250.400 ;
        RECT 441.200 248.800 442.000 250.400 ;
        RECT 442.800 250.300 443.600 255.800 ;
        RECT 444.400 253.600 445.200 255.200 ;
        RECT 449.600 254.300 450.400 259.800 ;
        RECT 455.000 255.800 456.600 259.800 ;
        RECT 467.800 255.800 469.400 259.800 ;
        RECT 476.800 258.400 477.600 259.800 ;
        RECT 476.800 257.600 478.800 258.400 ;
        RECT 481.200 257.600 482.000 259.800 ;
        RECT 452.400 254.300 453.200 254.400 ;
        RECT 449.600 253.800 453.200 254.300 ;
        RECT 449.800 253.700 453.200 253.800 ;
        RECT 449.800 253.600 451.400 253.700 ;
        RECT 452.400 253.600 453.200 253.700 ;
        RECT 454.000 253.600 454.800 254.400 ;
        RECT 447.600 251.600 449.200 252.400 ;
        RECT 446.000 250.300 446.800 251.200 ;
        RECT 442.800 249.700 446.800 250.300 ;
        RECT 442.800 242.200 443.600 249.700 ;
        RECT 446.000 249.600 446.800 249.700 ;
        RECT 450.800 250.400 451.400 253.600 ;
        RECT 454.200 253.200 454.800 253.600 ;
        RECT 454.200 252.400 455.000 253.200 ;
        RECT 455.600 252.400 456.200 255.800 ;
        RECT 457.200 252.800 458.000 254.400 ;
        RECT 465.200 254.300 466.000 254.400 ;
        RECT 466.800 254.300 467.600 254.400 ;
        RECT 465.200 253.700 467.600 254.300 ;
        RECT 465.200 253.600 466.000 253.700 ;
        RECT 466.800 253.600 467.600 253.700 ;
        RECT 467.000 253.200 467.600 253.600 ;
        RECT 467.000 252.400 467.800 253.200 ;
        RECT 468.400 252.400 469.000 255.800 ;
        RECT 470.000 252.800 470.800 254.400 ;
        RECT 476.800 254.200 477.600 257.600 ;
        RECT 479.600 255.600 480.400 257.200 ;
        RECT 481.400 254.400 482.000 257.600 ;
        RECT 476.800 253.800 478.600 254.200 ;
        RECT 477.000 253.600 478.600 253.800 ;
        RECT 481.200 253.600 482.000 254.400 ;
        RECT 452.400 250.800 453.200 252.400 ;
        RECT 455.600 251.600 456.400 252.400 ;
        RECT 458.800 252.200 459.600 252.400 ;
        RECT 458.000 251.600 459.600 252.200 ;
        RECT 455.600 251.400 456.200 251.600 ;
        RECT 454.200 250.800 456.200 251.400 ;
        RECT 458.000 251.200 458.800 251.600 ;
        RECT 465.200 250.800 466.000 252.400 ;
        RECT 468.400 251.600 469.200 252.400 ;
        RECT 471.600 252.200 472.400 252.400 ;
        RECT 470.800 251.600 472.400 252.200 ;
        RECT 474.800 251.600 476.400 252.400 ;
        RECT 468.400 251.400 469.000 251.600 ;
        RECT 467.000 250.800 469.000 251.400 ;
        RECT 470.800 251.200 471.600 251.600 ;
        RECT 450.800 249.600 451.600 250.400 ;
        RECT 454.200 250.200 454.800 250.800 ;
        RECT 467.000 250.200 467.600 250.800 ;
        RECT 449.200 247.600 450.000 249.200 ;
        RECT 450.800 247.000 451.400 249.600 ;
        RECT 447.800 246.400 451.400 247.000 ;
        RECT 447.800 246.200 448.400 246.400 ;
        RECT 447.600 242.200 448.400 246.200 ;
        RECT 450.800 246.200 451.400 246.400 ;
        RECT 450.800 242.200 451.600 246.200 ;
        RECT 452.400 242.800 453.200 250.200 ;
        RECT 454.000 243.400 454.800 250.200 ;
        RECT 455.600 249.600 459.600 250.200 ;
        RECT 455.600 242.800 456.400 249.600 ;
        RECT 452.400 242.200 456.400 242.800 ;
        RECT 458.800 242.200 459.600 249.600 ;
        RECT 465.200 242.800 466.000 250.200 ;
        RECT 466.800 243.400 467.600 250.200 ;
        RECT 468.400 249.600 472.400 250.200 ;
        RECT 473.200 249.600 474.000 251.200 ;
        RECT 478.000 250.400 478.600 253.600 ;
        RECT 478.000 249.600 478.800 250.400 ;
        RECT 481.400 250.200 482.000 253.600 ;
        RECT 486.000 257.800 486.800 259.800 ;
        RECT 486.000 254.400 486.600 257.800 ;
        RECT 487.600 255.600 488.400 257.200 ;
        RECT 486.000 253.600 486.800 254.400 ;
        RECT 482.800 250.800 483.600 252.400 ;
        RECT 484.400 250.800 485.200 252.400 ;
        RECT 486.000 250.200 486.600 253.600 ;
        RECT 468.400 242.800 469.200 249.600 ;
        RECT 465.200 242.200 469.200 242.800 ;
        RECT 471.600 242.200 472.400 249.600 ;
        RECT 476.400 247.600 477.200 249.200 ;
        RECT 478.000 247.000 478.600 249.600 ;
        RECT 481.200 249.400 483.000 250.200 ;
        RECT 475.000 246.400 478.600 247.000 ;
        RECT 475.000 246.200 475.600 246.400 ;
        RECT 474.800 242.200 475.600 246.200 ;
        RECT 478.000 246.200 478.600 246.400 ;
        RECT 478.000 242.200 478.800 246.200 ;
        RECT 482.200 244.400 483.000 249.400 ;
        RECT 485.000 249.400 486.800 250.200 ;
        RECT 485.000 244.400 485.800 249.400 ;
        RECT 481.200 243.600 483.000 244.400 ;
        RECT 484.400 243.600 485.800 244.400 ;
        RECT 482.200 242.200 483.000 243.600 ;
        RECT 485.000 242.200 485.800 243.600 ;
        RECT 489.200 242.200 490.000 259.800 ;
        RECT 490.800 255.600 491.600 257.200 ;
        RECT 492.400 242.200 493.200 259.800 ;
        RECT 494.000 255.600 494.800 257.200 ;
        RECT 498.800 255.800 499.600 259.800 ;
        RECT 500.200 256.400 501.000 257.200 ;
        RECT 502.600 256.400 503.400 259.800 ;
        RECT 497.200 252.800 498.000 254.400 ;
        RECT 498.800 254.300 499.400 255.800 ;
        RECT 500.400 255.600 501.200 256.400 ;
        RECT 502.600 255.800 504.400 256.400 ;
        RECT 502.000 254.300 502.800 254.400 ;
        RECT 498.800 253.700 502.800 254.300 ;
        RECT 495.600 252.200 496.400 252.400 ;
        RECT 498.800 252.200 499.400 253.700 ;
        RECT 502.000 253.600 502.800 253.700 ;
        RECT 500.400 252.200 501.200 252.400 ;
        RECT 495.600 251.600 497.200 252.200 ;
        RECT 498.800 251.600 501.200 252.200 ;
        RECT 496.400 251.200 497.200 251.600 ;
        RECT 500.400 250.200 501.000 251.600 ;
        RECT 495.600 249.600 499.600 250.200 ;
        RECT 495.600 242.200 496.400 249.600 ;
        RECT 498.800 242.200 499.600 249.600 ;
        RECT 500.400 242.200 501.200 250.200 ;
        RECT 502.000 248.800 502.800 250.400 ;
        RECT 503.600 242.200 504.400 255.800 ;
        RECT 505.200 253.600 506.000 255.200 ;
        RECT 508.000 254.200 508.800 259.800 ;
        RECT 507.000 253.800 508.800 254.200 ;
        RECT 514.800 257.600 515.600 259.800 ;
        RECT 518.000 259.200 522.000 259.800 ;
        RECT 514.800 254.400 515.400 257.600 ;
        RECT 516.400 255.600 517.200 257.200 ;
        RECT 518.000 255.800 518.800 259.200 ;
        RECT 519.600 255.800 520.400 258.600 ;
        RECT 521.200 256.000 522.000 259.200 ;
        RECT 524.400 256.000 525.200 259.800 ;
        RECT 521.200 255.800 525.200 256.000 ;
        RECT 526.000 259.200 530.000 259.800 ;
        RECT 526.000 255.800 526.800 259.200 ;
        RECT 527.600 255.800 528.400 258.600 ;
        RECT 529.200 256.000 530.000 259.200 ;
        RECT 532.400 256.000 533.200 259.800 ;
        RECT 529.200 255.800 533.200 256.000 ;
        RECT 519.600 254.400 520.200 255.800 ;
        RECT 521.400 255.400 525.000 255.800 ;
        RECT 523.600 254.400 524.400 254.800 ;
        RECT 527.600 254.400 528.200 255.800 ;
        RECT 529.400 255.400 533.000 255.800 ;
        RECT 534.000 255.600 534.800 257.200 ;
        RECT 531.600 254.400 532.400 254.800 ;
        RECT 507.000 253.600 508.600 253.800 ;
        RECT 514.800 253.600 515.600 254.400 ;
        RECT 507.000 250.400 507.600 253.600 ;
        RECT 509.200 251.600 510.800 252.400 ;
        RECT 506.800 249.600 507.600 250.400 ;
        RECT 511.600 249.600 512.400 251.200 ;
        RECT 513.200 250.800 514.000 252.400 ;
        RECT 514.800 250.200 515.400 253.600 ;
        RECT 518.000 252.800 518.800 254.400 ;
        RECT 519.600 253.800 522.000 254.400 ;
        RECT 523.600 254.300 525.200 254.400 ;
        RECT 526.000 254.300 526.800 254.400 ;
        RECT 523.600 253.800 526.800 254.300 ;
        RECT 527.600 253.800 530.000 254.400 ;
        RECT 531.600 254.300 533.200 254.400 ;
        RECT 535.600 254.300 536.400 259.800 ;
        RECT 537.200 259.200 541.200 259.800 ;
        RECT 537.200 255.800 538.000 259.200 ;
        RECT 538.800 255.800 539.600 258.600 ;
        RECT 540.400 256.000 541.200 259.200 ;
        RECT 543.600 256.000 544.400 259.800 ;
        RECT 540.400 255.800 544.400 256.000 ;
        RECT 538.800 254.400 539.400 255.800 ;
        RECT 540.600 255.400 544.200 255.800 ;
        RECT 542.800 254.400 543.600 254.800 ;
        RECT 537.200 254.300 538.000 254.400 ;
        RECT 531.600 253.800 538.000 254.300 ;
        RECT 538.800 253.800 541.200 254.400 ;
        RECT 542.800 253.800 544.400 254.400 ;
        RECT 521.200 253.600 522.000 253.800 ;
        RECT 524.400 253.700 526.800 253.800 ;
        RECT 524.400 253.600 525.200 253.700 ;
        RECT 519.600 251.600 520.400 253.200 ;
        RECT 521.400 250.200 522.000 253.600 ;
        RECT 522.800 251.600 523.600 253.200 ;
        RECT 526.000 252.800 526.800 253.700 ;
        RECT 529.200 253.600 530.000 253.800 ;
        RECT 532.400 253.700 538.000 253.800 ;
        RECT 532.400 253.600 533.200 253.700 ;
        RECT 527.600 251.600 528.400 253.200 ;
        RECT 529.400 250.200 530.000 253.600 ;
        RECT 530.800 252.300 531.600 253.200 ;
        RECT 534.000 252.300 534.800 252.400 ;
        RECT 530.800 251.700 534.800 252.300 ;
        RECT 530.800 251.600 531.600 251.700 ;
        RECT 534.000 251.600 534.800 251.700 ;
        RECT 507.000 247.000 507.600 249.600 ;
        RECT 513.800 249.400 515.600 250.200 ;
        RECT 508.400 247.600 509.200 249.200 ;
        RECT 507.000 246.400 510.600 247.000 ;
        RECT 507.000 246.200 507.600 246.400 ;
        RECT 506.800 242.200 507.600 246.200 ;
        RECT 510.000 246.200 510.600 246.400 ;
        RECT 510.000 242.200 510.800 246.200 ;
        RECT 513.800 242.200 514.600 249.400 ;
        RECT 520.600 242.200 522.600 250.200 ;
        RECT 528.600 242.200 530.600 250.200 ;
        RECT 535.600 242.200 536.400 253.700 ;
        RECT 537.200 252.800 538.000 253.700 ;
        RECT 540.400 253.600 541.200 253.800 ;
        RECT 543.600 253.600 544.400 253.800 ;
        RECT 545.200 253.600 546.000 255.200 ;
        RECT 538.800 251.600 539.600 253.200 ;
        RECT 540.600 250.400 541.200 253.600 ;
        RECT 542.000 251.600 542.800 253.200 ;
        RECT 546.800 252.300 547.600 259.800 ;
        RECT 548.400 256.000 549.200 259.800 ;
        RECT 551.600 256.000 552.400 259.800 ;
        RECT 548.400 255.800 552.400 256.000 ;
        RECT 553.200 255.800 554.000 259.800 ;
        RECT 548.600 255.400 552.200 255.800 ;
        RECT 549.200 254.400 550.000 254.800 ;
        RECT 553.200 254.400 553.800 255.800 ;
        RECT 556.400 255.200 557.200 259.800 ;
        RECT 559.600 255.200 560.400 259.800 ;
        RECT 562.800 255.200 563.600 259.800 ;
        RECT 566.000 255.200 566.800 259.800 ;
        RECT 570.800 256.000 571.600 259.800 ;
        RECT 570.600 255.200 571.600 256.000 ;
        RECT 556.400 254.400 558.200 255.200 ;
        RECT 559.600 254.400 561.800 255.200 ;
        RECT 562.800 254.400 565.000 255.200 ;
        RECT 566.000 254.400 568.400 255.200 ;
        RECT 548.400 253.800 550.000 254.400 ;
        RECT 548.400 253.600 549.200 253.800 ;
        RECT 551.400 253.600 554.000 254.400 ;
        RECT 554.800 253.800 555.600 254.400 ;
        RECT 557.400 253.800 558.200 254.400 ;
        RECT 561.000 253.800 561.800 254.400 ;
        RECT 564.200 253.800 565.000 254.400 ;
        RECT 550.000 252.300 550.800 253.200 ;
        RECT 546.800 251.700 550.800 252.300 ;
        RECT 538.800 250.200 541.200 250.400 ;
        RECT 538.800 249.600 541.800 250.200 ;
        RECT 539.800 242.200 541.800 249.600 ;
        RECT 546.800 242.200 547.600 251.700 ;
        RECT 550.000 251.600 550.800 251.700 ;
        RECT 551.400 250.200 552.000 253.600 ;
        RECT 554.800 253.000 556.600 253.800 ;
        RECT 557.400 253.000 560.000 253.800 ;
        RECT 561.000 253.000 563.400 253.800 ;
        RECT 564.200 253.000 566.800 253.800 ;
        RECT 557.400 251.600 558.200 253.000 ;
        RECT 561.000 251.600 561.800 253.000 ;
        RECT 564.200 251.600 565.000 253.000 ;
        RECT 567.600 251.600 568.400 254.400 ;
        RECT 556.400 250.800 558.200 251.600 ;
        RECT 559.600 250.800 561.800 251.600 ;
        RECT 562.800 250.800 565.000 251.600 ;
        RECT 566.000 250.800 568.400 251.600 ;
        RECT 570.600 250.800 571.400 255.200 ;
        RECT 572.400 254.600 573.200 259.800 ;
        RECT 578.800 256.600 579.600 259.800 ;
        RECT 580.400 257.000 581.200 259.800 ;
        RECT 582.000 257.000 582.800 259.800 ;
        RECT 583.600 257.000 584.400 259.800 ;
        RECT 585.200 257.000 586.000 259.800 ;
        RECT 588.400 257.000 589.200 259.800 ;
        RECT 591.600 257.000 592.400 259.800 ;
        RECT 593.200 257.000 594.000 259.800 ;
        RECT 594.800 257.000 595.600 259.800 ;
        RECT 577.200 255.800 579.600 256.600 ;
        RECT 596.400 256.600 597.200 259.800 ;
        RECT 577.200 255.200 578.000 255.800 ;
        RECT 572.000 254.000 573.200 254.600 ;
        RECT 576.200 254.600 578.000 255.200 ;
        RECT 582.000 255.600 583.000 256.400 ;
        RECT 586.000 255.600 587.600 256.400 ;
        RECT 588.400 255.800 593.000 256.400 ;
        RECT 596.400 255.800 599.000 256.600 ;
        RECT 588.400 255.600 589.200 255.800 ;
        RECT 572.000 252.000 572.600 254.000 ;
        RECT 576.200 253.400 577.000 254.600 ;
        RECT 573.200 252.600 577.000 253.400 ;
        RECT 582.000 252.800 582.800 255.600 ;
        RECT 588.400 254.800 589.200 255.000 ;
        RECT 584.800 254.200 589.200 254.800 ;
        RECT 584.800 254.000 585.600 254.200 ;
        RECT 590.000 253.600 590.800 255.200 ;
        RECT 592.200 253.400 593.000 255.800 ;
        RECT 598.200 255.200 599.000 255.800 ;
        RECT 598.200 254.400 601.200 255.200 ;
        RECT 602.800 253.800 603.600 259.800 ;
        RECT 604.400 255.200 605.200 259.800 ;
        RECT 604.400 254.600 606.600 255.200 ;
        RECT 585.200 252.600 588.400 253.400 ;
        RECT 592.200 252.600 594.200 253.400 ;
        RECT 594.800 253.000 603.600 253.800 ;
        RECT 578.800 252.000 579.600 252.600 ;
        RECT 596.400 252.000 597.200 252.400 ;
        RECT 601.400 252.000 602.200 252.200 ;
        RECT 572.000 251.400 572.800 252.000 ;
        RECT 578.800 251.400 602.200 252.000 ;
        RECT 553.200 250.200 554.000 250.400 ;
        RECT 551.000 249.600 552.000 250.200 ;
        RECT 552.600 249.600 554.000 250.200 ;
        RECT 551.000 244.400 551.800 249.600 ;
        RECT 552.600 248.400 553.200 249.600 ;
        RECT 552.400 247.600 553.200 248.400 ;
        RECT 550.000 243.600 551.800 244.400 ;
        RECT 551.000 242.200 551.800 243.600 ;
        RECT 556.400 242.200 557.200 250.800 ;
        RECT 559.600 242.200 560.400 250.800 ;
        RECT 562.800 242.200 563.600 250.800 ;
        RECT 566.000 242.200 566.800 250.800 ;
        RECT 570.600 250.000 571.600 250.800 ;
        RECT 570.800 242.200 571.600 250.000 ;
        RECT 572.200 249.600 572.800 251.400 ;
        RECT 572.200 249.000 581.200 249.600 ;
        RECT 572.200 247.400 572.800 249.000 ;
        RECT 580.400 248.800 581.200 249.000 ;
        RECT 583.600 249.000 592.200 249.600 ;
        RECT 583.600 248.800 584.400 249.000 ;
        RECT 575.400 247.600 578.000 248.400 ;
        RECT 572.200 246.800 574.800 247.400 ;
        RECT 574.000 242.200 574.800 246.800 ;
        RECT 577.200 242.200 578.000 247.600 ;
        RECT 578.600 246.800 582.800 247.600 ;
        RECT 580.400 242.200 581.200 245.000 ;
        RECT 582.000 242.200 582.800 245.000 ;
        RECT 583.600 242.200 584.400 245.000 ;
        RECT 585.200 242.200 586.000 248.400 ;
        RECT 588.400 247.600 591.000 248.400 ;
        RECT 591.600 248.200 592.200 249.000 ;
        RECT 593.200 249.400 594.000 249.600 ;
        RECT 593.200 249.000 598.600 249.400 ;
        RECT 593.200 248.800 599.400 249.000 ;
        RECT 598.000 248.200 599.400 248.800 ;
        RECT 591.600 247.600 597.400 248.200 ;
        RECT 600.400 248.000 602.000 248.800 ;
        RECT 600.400 247.600 601.000 248.000 ;
        RECT 588.400 242.200 589.200 247.000 ;
        RECT 591.600 242.200 592.400 247.000 ;
        RECT 596.800 246.800 601.000 247.600 ;
        RECT 602.800 247.400 603.600 253.000 ;
        RECT 604.400 251.600 605.200 253.200 ;
        RECT 606.000 251.600 606.600 254.600 ;
        RECT 606.000 250.800 607.200 251.600 ;
        RECT 606.000 250.200 606.600 250.800 ;
        RECT 601.600 246.800 603.600 247.400 ;
        RECT 604.400 249.600 606.600 250.200 ;
        RECT 593.200 242.200 594.000 245.000 ;
        RECT 594.800 242.200 595.600 245.000 ;
        RECT 598.000 242.200 598.800 246.800 ;
        RECT 601.600 246.200 602.200 246.800 ;
        RECT 601.200 245.600 602.200 246.200 ;
        RECT 601.200 242.200 602.000 245.600 ;
        RECT 604.400 242.200 605.200 249.600 ;
        RECT 2.800 222.200 3.600 239.800 ;
        RECT 6.000 222.200 6.800 239.800 ;
        RECT 10.200 232.400 11.000 239.800 ;
        RECT 16.600 234.400 17.400 239.800 ;
        RECT 23.000 238.400 23.800 239.800 ;
        RECT 22.000 237.600 23.800 238.400 ;
        RECT 11.600 233.600 12.400 234.400 ;
        RECT 15.600 233.600 17.400 234.400 ;
        RECT 18.000 233.600 18.800 234.400 ;
        RECT 11.800 232.400 12.400 233.600 ;
        RECT 16.600 232.400 17.400 233.600 ;
        RECT 18.200 232.400 18.800 233.600 ;
        RECT 23.000 232.400 23.800 237.600 ;
        RECT 24.400 233.600 25.200 234.400 ;
        RECT 24.600 232.400 25.200 233.600 ;
        RECT 10.200 231.800 11.200 232.400 ;
        RECT 11.800 231.800 13.200 232.400 ;
        RECT 16.600 231.800 17.600 232.400 ;
        RECT 18.200 231.800 19.600 232.400 ;
        RECT 23.000 231.800 24.000 232.400 ;
        RECT 24.600 231.800 26.000 232.400 ;
        RECT 9.200 228.800 10.000 230.400 ;
        RECT 10.600 230.300 11.200 231.800 ;
        RECT 12.400 231.600 13.200 231.800 ;
        RECT 14.000 230.300 14.800 230.400 ;
        RECT 10.600 229.700 14.800 230.300 ;
        RECT 10.600 228.400 11.200 229.700 ;
        RECT 14.000 229.600 14.800 229.700 ;
        RECT 15.600 228.800 16.400 230.400 ;
        RECT 17.000 228.400 17.600 231.800 ;
        RECT 18.800 231.600 19.600 231.800 ;
        RECT 22.000 228.800 22.800 230.400 ;
        RECT 23.400 228.400 24.000 231.800 ;
        RECT 25.200 231.600 26.000 231.800 ;
        RECT 7.600 228.200 8.400 228.400 ;
        RECT 7.600 227.600 9.200 228.200 ;
        RECT 10.600 227.600 13.200 228.400 ;
        RECT 14.000 228.200 14.800 228.400 ;
        RECT 14.000 227.600 15.600 228.200 ;
        RECT 17.000 227.600 19.600 228.400 ;
        RECT 20.400 228.200 21.200 228.400 ;
        RECT 20.400 227.600 22.000 228.200 ;
        RECT 23.400 227.600 26.000 228.400 ;
        RECT 8.400 227.200 9.200 227.600 ;
        RECT 7.800 226.200 11.400 226.600 ;
        RECT 12.400 226.200 13.000 227.600 ;
        RECT 14.800 227.200 15.600 227.600 ;
        RECT 14.200 226.200 17.800 226.600 ;
        RECT 18.800 226.200 19.400 227.600 ;
        RECT 21.200 227.200 22.000 227.600 ;
        RECT 20.600 226.200 24.200 226.600 ;
        RECT 25.200 226.200 25.800 227.600 ;
        RECT 26.800 226.800 27.600 228.400 ;
        RECT 28.400 226.200 29.200 239.800 ;
        RECT 30.000 231.600 30.800 234.400 ;
        RECT 34.200 232.400 35.000 239.800 ;
        RECT 35.600 233.600 36.400 234.400 ;
        RECT 35.800 232.400 36.400 233.600 ;
        RECT 33.200 231.600 35.200 232.400 ;
        RECT 35.800 231.800 37.200 232.400 ;
        RECT 36.400 231.600 37.200 231.800 ;
        RECT 33.200 228.800 34.000 230.400 ;
        RECT 34.600 228.400 35.200 231.600 ;
        RECT 31.600 228.200 32.400 228.400 ;
        RECT 31.600 227.600 33.200 228.200 ;
        RECT 34.600 227.600 37.200 228.400 ;
        RECT 32.400 227.200 33.200 227.600 ;
        RECT 31.800 226.200 35.400 226.600 ;
        RECT 36.400 226.200 37.000 227.600 ;
        RECT 7.600 226.000 11.600 226.200 ;
        RECT 7.600 222.200 8.400 226.000 ;
        RECT 10.800 222.200 11.600 226.000 ;
        RECT 12.400 222.200 13.200 226.200 ;
        RECT 14.000 226.000 18.000 226.200 ;
        RECT 14.000 222.200 14.800 226.000 ;
        RECT 17.200 222.200 18.000 226.000 ;
        RECT 18.800 222.200 19.600 226.200 ;
        RECT 20.400 226.000 24.400 226.200 ;
        RECT 20.400 222.200 21.200 226.000 ;
        RECT 23.600 222.200 24.400 226.000 ;
        RECT 25.200 222.200 26.000 226.200 ;
        RECT 28.400 225.600 30.200 226.200 ;
        RECT 29.400 224.400 30.200 225.600 ;
        RECT 28.400 223.600 30.200 224.400 ;
        RECT 29.400 222.200 30.200 223.600 ;
        RECT 31.600 226.000 35.600 226.200 ;
        RECT 31.600 222.200 32.400 226.000 ;
        RECT 34.800 222.200 35.600 226.000 ;
        RECT 36.400 222.200 37.200 226.200 ;
        RECT 38.000 222.200 38.800 239.800 ;
        RECT 39.600 224.800 40.400 226.400 ;
        RECT 41.200 224.800 42.000 226.400 ;
        RECT 42.800 222.200 43.600 239.800 ;
        RECT 46.000 236.400 46.800 239.800 ;
        RECT 45.800 235.800 46.800 236.400 ;
        RECT 45.800 235.200 46.400 235.800 ;
        RECT 49.200 235.200 50.000 239.800 ;
        RECT 52.400 237.000 53.200 239.800 ;
        RECT 54.000 237.000 54.800 239.800 ;
        RECT 44.400 234.600 46.400 235.200 ;
        RECT 44.400 229.000 45.200 234.600 ;
        RECT 47.000 234.400 51.200 235.200 ;
        RECT 55.600 235.000 56.400 239.800 ;
        RECT 58.800 235.000 59.600 239.800 ;
        RECT 47.000 234.000 47.600 234.400 ;
        RECT 46.000 233.200 47.600 234.000 ;
        RECT 50.600 233.800 56.400 234.400 ;
        RECT 48.600 233.200 50.000 233.800 ;
        RECT 48.600 233.000 54.800 233.200 ;
        RECT 49.400 232.600 54.800 233.000 ;
        RECT 54.000 232.400 54.800 232.600 ;
        RECT 55.800 233.000 56.400 233.800 ;
        RECT 57.000 233.600 59.600 234.400 ;
        RECT 62.000 233.600 62.800 239.800 ;
        RECT 63.600 237.000 64.400 239.800 ;
        RECT 65.200 237.000 66.000 239.800 ;
        RECT 66.800 237.000 67.600 239.800 ;
        RECT 65.200 234.400 69.400 235.200 ;
        RECT 70.000 234.400 70.800 239.800 ;
        RECT 73.200 235.200 74.000 239.800 ;
        RECT 73.200 234.600 75.800 235.200 ;
        RECT 70.000 233.600 72.600 234.400 ;
        RECT 63.600 233.000 64.400 233.200 ;
        RECT 55.800 232.400 64.400 233.000 ;
        RECT 66.800 233.000 67.600 233.200 ;
        RECT 75.200 233.000 75.800 234.600 ;
        RECT 66.800 232.400 75.800 233.000 ;
        RECT 75.200 230.600 75.800 232.400 ;
        RECT 76.400 232.000 77.200 239.800 ;
        RECT 78.000 234.300 78.800 234.400 ;
        RECT 81.200 234.300 82.000 239.800 ;
        RECT 82.800 234.300 83.600 234.400 ;
        RECT 78.000 233.700 80.400 234.300 ;
        RECT 78.000 233.600 78.800 233.700 ;
        RECT 76.400 231.200 77.400 232.000 ;
        RECT 79.600 231.600 80.400 233.700 ;
        RECT 81.200 233.700 83.600 234.300 ;
        RECT 45.800 230.000 69.200 230.600 ;
        RECT 75.200 230.000 76.000 230.600 ;
        RECT 45.800 229.800 46.600 230.000 ;
        RECT 47.600 229.600 48.400 230.000 ;
        RECT 50.800 229.600 51.600 230.000 ;
        RECT 68.400 229.400 69.200 230.000 ;
        RECT 44.400 228.200 53.200 229.000 ;
        RECT 53.800 228.600 55.800 229.400 ;
        RECT 59.600 228.600 62.800 229.400 ;
        RECT 44.400 222.200 45.200 228.200 ;
        RECT 46.800 226.800 49.800 227.600 ;
        RECT 49.000 226.200 49.800 226.800 ;
        RECT 55.000 226.200 55.800 228.600 ;
        RECT 57.200 226.800 58.000 228.400 ;
        RECT 62.400 227.800 63.200 228.000 ;
        RECT 58.800 227.200 63.200 227.800 ;
        RECT 58.800 227.000 59.600 227.200 ;
        RECT 65.200 226.400 66.000 229.200 ;
        RECT 71.000 228.600 74.800 229.400 ;
        RECT 71.000 227.400 71.800 228.600 ;
        RECT 75.400 228.000 76.000 230.000 ;
        RECT 58.800 226.200 59.600 226.400 ;
        RECT 49.000 225.400 51.600 226.200 ;
        RECT 55.000 225.600 59.600 226.200 ;
        RECT 60.400 225.600 62.000 226.400 ;
        RECT 65.000 225.600 66.000 226.400 ;
        RECT 70.000 226.800 71.800 227.400 ;
        RECT 74.800 227.400 76.000 228.000 ;
        RECT 70.000 226.200 70.800 226.800 ;
        RECT 50.800 222.200 51.600 225.400 ;
        RECT 68.400 225.400 70.800 226.200 ;
        RECT 52.400 222.200 53.200 225.000 ;
        RECT 54.000 222.200 54.800 225.000 ;
        RECT 55.600 222.200 56.400 225.000 ;
        RECT 58.800 222.200 59.600 225.000 ;
        RECT 62.000 222.200 62.800 225.000 ;
        RECT 63.600 222.200 64.400 225.000 ;
        RECT 65.200 222.200 66.000 225.000 ;
        RECT 66.800 222.200 67.600 225.000 ;
        RECT 68.400 222.200 69.200 225.400 ;
        RECT 74.800 222.200 75.600 227.400 ;
        RECT 76.600 226.800 77.400 231.200 ;
        RECT 76.400 226.000 77.400 226.800 ;
        RECT 81.200 226.200 82.000 233.700 ;
        RECT 82.800 233.600 83.600 233.700 ;
        RECT 86.000 231.200 86.800 239.800 ;
        RECT 89.200 231.200 90.000 239.800 ;
        RECT 92.400 231.200 93.200 239.800 ;
        RECT 95.600 231.200 96.400 239.800 ;
        RECT 98.800 232.400 99.600 239.800 ;
        RECT 102.000 232.800 102.800 239.800 ;
        RECT 98.800 231.800 101.400 232.400 ;
        RECT 102.000 231.800 103.000 232.800 ;
        RECT 86.000 230.400 87.800 231.200 ;
        RECT 89.200 230.400 91.400 231.200 ;
        RECT 92.400 230.400 94.600 231.200 ;
        RECT 95.600 230.400 98.000 231.200 ;
        RECT 87.000 229.000 87.800 230.400 ;
        RECT 90.600 229.000 91.400 230.400 ;
        RECT 93.800 229.000 94.600 230.400 ;
        RECT 82.800 226.800 83.600 228.400 ;
        RECT 84.400 228.200 86.200 229.000 ;
        RECT 87.000 228.200 89.600 229.000 ;
        RECT 90.600 228.200 93.000 229.000 ;
        RECT 93.800 228.200 96.400 229.000 ;
        RECT 84.400 227.600 85.200 228.200 ;
        RECT 87.000 227.600 87.800 228.200 ;
        RECT 90.600 227.600 91.400 228.200 ;
        RECT 93.800 227.600 94.600 228.200 ;
        RECT 97.200 227.600 98.000 230.400 ;
        RECT 86.000 226.800 87.800 227.600 ;
        RECT 89.200 226.800 91.400 227.600 ;
        RECT 92.400 226.800 94.600 227.600 ;
        RECT 95.600 226.800 98.000 227.600 ;
        RECT 100.800 229.800 101.400 231.800 ;
        RECT 100.800 229.000 101.800 229.800 ;
        RECT 100.800 227.400 101.400 229.000 ;
        RECT 102.400 228.400 103.000 231.800 ;
        RECT 105.200 231.400 106.000 239.800 ;
        RECT 109.600 236.400 110.400 239.800 ;
        RECT 108.400 235.800 110.400 236.400 ;
        RECT 114.000 235.800 114.800 239.800 ;
        RECT 118.200 235.800 119.400 239.800 ;
        RECT 108.400 235.000 109.200 235.800 ;
        RECT 114.000 235.200 114.600 235.800 ;
        RECT 111.800 234.600 115.400 235.200 ;
        RECT 118.000 235.000 118.800 235.800 ;
        RECT 111.800 234.400 112.600 234.600 ;
        RECT 114.600 234.400 115.400 234.600 ;
        RECT 108.400 233.000 109.200 233.200 ;
        RECT 113.000 233.000 113.800 233.200 ;
        RECT 108.400 232.400 113.800 233.000 ;
        RECT 114.400 233.000 116.600 233.600 ;
        RECT 114.400 231.800 115.000 233.000 ;
        RECT 115.800 232.800 116.600 233.000 ;
        RECT 118.200 233.200 119.600 234.000 ;
        RECT 118.200 232.200 118.800 233.200 ;
        RECT 110.200 231.400 115.000 231.800 ;
        RECT 105.200 231.200 115.000 231.400 ;
        RECT 116.400 231.600 118.800 232.200 ;
        RECT 105.200 231.000 111.000 231.200 ;
        RECT 105.200 230.800 110.800 231.000 ;
        RECT 111.600 230.300 112.400 230.400 ;
        RECT 114.800 230.300 115.600 230.400 ;
        RECT 111.600 230.200 115.600 230.300 ;
        RECT 107.400 229.700 115.600 230.200 ;
        RECT 107.400 229.600 112.400 229.700 ;
        RECT 114.800 229.600 115.600 229.700 ;
        RECT 107.400 229.400 108.200 229.600 ;
        RECT 109.000 228.400 109.800 228.600 ;
        RECT 116.400 228.400 117.000 231.600 ;
        RECT 122.800 231.200 123.600 239.800 ;
        RECT 125.200 233.600 126.000 234.400 ;
        RECT 125.200 232.400 125.800 233.600 ;
        RECT 126.600 232.400 127.400 239.800 ;
        RECT 131.400 232.600 132.200 239.800 ;
        RECT 124.400 231.800 125.800 232.400 ;
        RECT 124.400 231.600 125.200 231.800 ;
        RECT 126.400 231.600 128.400 232.400 ;
        RECT 131.400 231.800 133.200 232.600 ;
        RECT 138.200 232.400 139.000 239.800 ;
        RECT 139.600 233.600 140.400 234.400 ;
        RECT 139.800 232.400 140.400 233.600 ;
        RECT 138.200 231.800 139.200 232.400 ;
        RECT 139.800 232.300 141.200 232.400 ;
        RECT 142.000 232.300 142.800 239.800 ;
        RECT 151.600 236.400 152.400 239.800 ;
        RECT 151.400 235.800 152.400 236.400 ;
        RECT 151.400 235.200 152.000 235.800 ;
        RECT 154.800 235.200 155.600 239.800 ;
        RECT 158.000 237.000 158.800 239.800 ;
        RECT 159.600 237.000 160.400 239.800 ;
        RECT 139.800 231.800 142.800 232.300 ;
        RECT 119.400 230.600 123.600 231.200 ;
        RECT 119.400 230.400 120.200 230.600 ;
        RECT 121.000 229.800 121.800 230.000 ;
        RECT 118.000 229.200 121.800 229.800 ;
        RECT 118.000 229.000 118.800 229.200 ;
        RECT 102.000 227.600 103.000 228.400 ;
        RECT 106.000 227.800 117.000 228.400 ;
        RECT 106.000 227.600 107.600 227.800 ;
        RECT 98.800 226.800 101.400 227.400 ;
        RECT 76.400 222.200 77.200 226.000 ;
        RECT 80.200 225.600 82.000 226.200 ;
        RECT 80.200 222.200 81.000 225.600 ;
        RECT 86.000 222.200 86.800 226.800 ;
        RECT 89.200 222.200 90.000 226.800 ;
        RECT 92.400 222.200 93.200 226.800 ;
        RECT 95.600 222.200 96.400 226.800 ;
        RECT 98.800 222.200 99.600 226.800 ;
        RECT 102.400 226.200 103.000 227.600 ;
        RECT 102.000 225.600 103.000 226.200 ;
        RECT 102.000 222.200 102.800 225.600 ;
        RECT 105.200 222.200 106.000 227.000 ;
        RECT 110.200 225.600 110.800 227.800 ;
        RECT 115.800 227.600 116.600 227.800 ;
        RECT 122.800 227.200 123.600 230.600 ;
        RECT 126.400 228.400 127.000 231.600 ;
        RECT 127.600 230.300 128.400 230.400 ;
        RECT 129.200 230.300 130.000 230.400 ;
        RECT 127.600 229.700 130.000 230.300 ;
        RECT 127.600 228.800 128.400 229.700 ;
        RECT 129.200 229.600 130.000 229.700 ;
        RECT 130.800 229.600 131.600 231.200 ;
        RECT 124.400 227.600 127.000 228.400 ;
        RECT 129.200 228.300 130.000 228.400 ;
        RECT 130.900 228.300 131.500 229.600 ;
        RECT 129.200 228.200 131.500 228.300 ;
        RECT 128.400 227.700 131.500 228.200 ;
        RECT 132.400 228.400 133.000 231.800 ;
        RECT 134.000 230.300 134.800 230.400 ;
        RECT 137.200 230.300 138.000 230.400 ;
        RECT 134.000 229.700 138.000 230.300 ;
        RECT 134.000 229.600 134.800 229.700 ;
        RECT 137.200 228.800 138.000 229.700 ;
        RECT 138.600 228.400 139.200 231.800 ;
        RECT 140.400 231.700 142.800 231.800 ;
        RECT 140.400 231.600 141.200 231.700 ;
        RECT 128.400 227.600 130.000 227.700 ;
        RECT 132.400 227.600 133.200 228.400 ;
        RECT 135.600 228.300 136.400 228.400 ;
        RECT 134.100 228.200 136.400 228.300 ;
        RECT 134.100 227.700 137.200 228.200 ;
        RECT 119.800 226.600 123.600 227.200 ;
        RECT 119.800 226.400 120.600 226.600 ;
        RECT 108.400 224.200 109.200 225.000 ;
        RECT 110.000 224.800 110.800 225.600 ;
        RECT 111.800 225.400 112.600 225.600 ;
        RECT 111.800 224.800 114.600 225.400 ;
        RECT 114.000 224.200 114.600 224.800 ;
        RECT 118.000 224.200 118.800 225.000 ;
        RECT 108.400 223.600 110.400 224.200 ;
        RECT 109.600 222.200 110.400 223.600 ;
        RECT 114.000 222.200 114.800 224.200 ;
        RECT 118.000 223.600 119.400 224.200 ;
        RECT 118.200 222.200 119.400 223.600 ;
        RECT 122.800 222.200 123.600 226.600 ;
        RECT 124.600 226.200 125.200 227.600 ;
        RECT 128.400 227.200 129.200 227.600 ;
        RECT 126.200 226.200 129.800 226.600 ;
        RECT 124.400 222.200 125.200 226.200 ;
        RECT 126.000 226.000 130.000 226.200 ;
        RECT 126.000 222.200 126.800 226.000 ;
        RECT 129.200 222.200 130.000 226.000 ;
        RECT 132.400 224.400 133.000 227.600 ;
        RECT 134.100 226.400 134.700 227.700 ;
        RECT 135.600 227.600 137.200 227.700 ;
        RECT 138.600 227.600 141.200 228.400 ;
        RECT 136.400 227.200 137.200 227.600 ;
        RECT 134.000 224.800 134.800 226.400 ;
        RECT 135.800 226.200 139.400 226.600 ;
        RECT 140.400 226.200 141.000 227.600 ;
        RECT 135.600 226.000 139.600 226.200 ;
        RECT 132.400 222.200 133.200 224.400 ;
        RECT 135.600 222.200 136.400 226.000 ;
        RECT 138.800 222.200 139.600 226.000 ;
        RECT 140.400 222.200 141.200 226.200 ;
        RECT 142.000 222.200 142.800 231.700 ;
        RECT 150.000 234.600 152.000 235.200 ;
        RECT 150.000 229.000 150.800 234.600 ;
        RECT 152.600 234.400 156.800 235.200 ;
        RECT 161.200 235.000 162.000 239.800 ;
        RECT 164.400 235.000 165.200 239.800 ;
        RECT 152.600 234.000 153.200 234.400 ;
        RECT 151.600 233.200 153.200 234.000 ;
        RECT 156.200 233.800 162.000 234.400 ;
        RECT 154.200 233.200 155.600 233.800 ;
        RECT 154.200 233.000 160.400 233.200 ;
        RECT 155.000 232.600 160.400 233.000 ;
        RECT 159.600 232.400 160.400 232.600 ;
        RECT 161.400 233.000 162.000 233.800 ;
        RECT 162.600 233.600 165.200 234.400 ;
        RECT 167.600 233.600 168.400 239.800 ;
        RECT 169.200 237.000 170.000 239.800 ;
        RECT 170.800 237.000 171.600 239.800 ;
        RECT 172.400 237.000 173.200 239.800 ;
        RECT 170.800 234.400 175.000 235.200 ;
        RECT 175.600 234.400 176.400 239.800 ;
        RECT 178.800 235.200 179.600 239.800 ;
        RECT 178.800 234.600 181.400 235.200 ;
        RECT 175.600 233.600 178.200 234.400 ;
        RECT 169.200 233.000 170.000 233.200 ;
        RECT 161.400 232.400 170.000 233.000 ;
        RECT 172.400 233.000 173.200 233.200 ;
        RECT 180.800 233.000 181.400 234.600 ;
        RECT 172.400 232.400 181.400 233.000 ;
        RECT 180.800 230.600 181.400 232.400 ;
        RECT 182.000 232.000 182.800 239.800 ;
        RECT 182.000 231.200 183.000 232.000 ;
        RECT 151.400 230.000 174.800 230.600 ;
        RECT 180.800 230.000 181.600 230.600 ;
        RECT 151.400 229.800 152.200 230.000 ;
        RECT 156.400 229.600 157.200 230.000 ;
        RECT 174.000 229.400 174.800 230.000 ;
        RECT 150.000 228.200 158.800 229.000 ;
        RECT 159.400 228.600 161.400 229.400 ;
        RECT 165.200 228.600 168.400 229.400 ;
        RECT 143.600 224.800 144.400 226.400 ;
        RECT 150.000 222.200 150.800 228.200 ;
        RECT 152.400 226.800 155.400 227.600 ;
        RECT 154.600 226.200 155.400 226.800 ;
        RECT 160.600 226.200 161.400 228.600 ;
        RECT 162.800 226.800 163.600 228.400 ;
        RECT 168.000 227.800 168.800 228.000 ;
        RECT 164.400 227.200 168.800 227.800 ;
        RECT 164.400 227.000 165.200 227.200 ;
        RECT 170.800 226.400 171.600 229.200 ;
        RECT 176.600 228.600 180.400 229.400 ;
        RECT 176.600 227.400 177.400 228.600 ;
        RECT 181.000 228.000 181.600 230.000 ;
        RECT 164.400 226.200 165.200 226.400 ;
        RECT 154.600 225.400 157.200 226.200 ;
        RECT 160.600 225.600 165.200 226.200 ;
        RECT 166.000 225.600 167.600 226.400 ;
        RECT 170.600 225.600 171.600 226.400 ;
        RECT 175.600 226.800 177.400 227.400 ;
        RECT 180.400 227.400 181.600 228.000 ;
        RECT 175.600 226.200 176.400 226.800 ;
        RECT 156.400 222.200 157.200 225.400 ;
        RECT 174.000 225.400 176.400 226.200 ;
        RECT 158.000 222.200 158.800 225.000 ;
        RECT 159.600 222.200 160.400 225.000 ;
        RECT 161.200 222.200 162.000 225.000 ;
        RECT 164.400 222.200 165.200 225.000 ;
        RECT 167.600 222.200 168.400 225.000 ;
        RECT 169.200 222.200 170.000 225.000 ;
        RECT 170.800 222.200 171.600 225.000 ;
        RECT 172.400 222.200 173.200 225.000 ;
        RECT 174.000 222.200 174.800 225.400 ;
        RECT 180.400 222.200 181.200 227.400 ;
        RECT 182.200 226.800 183.000 231.200 ;
        RECT 182.000 226.000 183.000 226.800 ;
        RECT 182.000 222.200 182.800 226.000 ;
        RECT 185.200 224.800 186.000 226.400 ;
        RECT 186.800 222.200 187.600 239.800 ;
        RECT 190.000 236.400 190.800 239.800 ;
        RECT 189.800 235.800 190.800 236.400 ;
        RECT 189.800 235.200 190.400 235.800 ;
        RECT 193.200 235.200 194.000 239.800 ;
        RECT 196.400 237.000 197.200 239.800 ;
        RECT 198.000 237.000 198.800 239.800 ;
        RECT 188.400 234.600 190.400 235.200 ;
        RECT 188.400 229.000 189.200 234.600 ;
        RECT 191.000 234.400 195.200 235.200 ;
        RECT 199.600 235.000 200.400 239.800 ;
        RECT 202.800 235.000 203.600 239.800 ;
        RECT 191.000 234.000 191.600 234.400 ;
        RECT 190.000 233.200 191.600 234.000 ;
        RECT 194.600 233.800 200.400 234.400 ;
        RECT 192.600 233.200 194.000 233.800 ;
        RECT 192.600 233.000 198.800 233.200 ;
        RECT 193.400 232.600 198.800 233.000 ;
        RECT 198.000 232.400 198.800 232.600 ;
        RECT 199.800 233.000 200.400 233.800 ;
        RECT 201.000 233.600 203.600 234.400 ;
        RECT 206.000 233.600 206.800 239.800 ;
        RECT 207.600 237.000 208.400 239.800 ;
        RECT 209.200 237.000 210.000 239.800 ;
        RECT 210.800 237.000 211.600 239.800 ;
        RECT 209.200 234.400 213.400 235.200 ;
        RECT 214.000 234.400 214.800 239.800 ;
        RECT 217.200 235.200 218.000 239.800 ;
        RECT 217.200 234.600 219.800 235.200 ;
        RECT 214.000 233.600 216.600 234.400 ;
        RECT 207.600 233.000 208.400 233.200 ;
        RECT 199.800 232.400 208.400 233.000 ;
        RECT 210.800 233.000 211.600 233.200 ;
        RECT 219.200 233.000 219.800 234.600 ;
        RECT 210.800 232.400 219.800 233.000 ;
        RECT 219.200 230.600 219.800 232.400 ;
        RECT 220.400 232.000 221.200 239.800 ;
        RECT 220.400 231.200 221.400 232.000 ;
        RECT 189.800 230.000 213.200 230.600 ;
        RECT 219.200 230.000 220.000 230.600 ;
        RECT 189.800 229.800 190.600 230.000 ;
        RECT 194.800 229.600 195.600 230.000 ;
        RECT 212.400 229.400 213.200 230.000 ;
        RECT 188.400 228.200 197.200 229.000 ;
        RECT 197.800 228.600 199.800 229.400 ;
        RECT 203.600 228.600 206.800 229.400 ;
        RECT 188.400 222.200 189.200 228.200 ;
        RECT 190.800 226.800 193.800 227.600 ;
        RECT 193.000 226.200 193.800 226.800 ;
        RECT 199.000 226.200 199.800 228.600 ;
        RECT 201.200 226.800 202.000 228.400 ;
        RECT 206.400 227.800 207.200 228.000 ;
        RECT 202.800 227.200 207.200 227.800 ;
        RECT 202.800 227.000 203.600 227.200 ;
        RECT 209.200 226.400 210.000 229.200 ;
        RECT 215.000 228.600 218.800 229.400 ;
        RECT 215.000 227.400 215.800 228.600 ;
        RECT 219.400 228.000 220.000 230.000 ;
        RECT 202.800 226.200 203.600 226.400 ;
        RECT 193.000 225.400 195.600 226.200 ;
        RECT 199.000 225.600 203.600 226.200 ;
        RECT 204.400 225.600 206.000 226.400 ;
        RECT 209.000 225.600 210.000 226.400 ;
        RECT 214.000 226.800 215.800 227.400 ;
        RECT 218.800 227.400 220.000 228.000 ;
        RECT 214.000 226.200 214.800 226.800 ;
        RECT 194.800 222.200 195.600 225.400 ;
        RECT 212.400 225.400 214.800 226.200 ;
        RECT 196.400 222.200 197.200 225.000 ;
        RECT 198.000 222.200 198.800 225.000 ;
        RECT 199.600 222.200 200.400 225.000 ;
        RECT 202.800 222.200 203.600 225.000 ;
        RECT 206.000 222.200 206.800 225.000 ;
        RECT 207.600 222.200 208.400 225.000 ;
        RECT 209.200 222.200 210.000 225.000 ;
        RECT 210.800 222.200 211.600 225.000 ;
        RECT 212.400 222.200 213.200 225.400 ;
        RECT 218.800 222.200 219.600 227.400 ;
        RECT 220.600 226.800 221.400 231.200 ;
        RECT 220.400 226.000 221.400 226.800 ;
        RECT 225.200 231.200 226.000 239.800 ;
        RECT 228.400 231.200 229.200 239.800 ;
        RECT 233.200 236.400 234.000 239.800 ;
        RECT 233.000 235.800 234.000 236.400 ;
        RECT 233.000 235.200 233.600 235.800 ;
        RECT 236.400 235.200 237.200 239.800 ;
        RECT 239.600 237.000 240.400 239.800 ;
        RECT 241.200 237.000 242.000 239.800 ;
        RECT 225.200 230.400 229.200 231.200 ;
        RECT 231.600 234.600 233.600 235.200 ;
        RECT 225.200 227.600 226.000 230.400 ;
        RECT 231.600 229.000 232.400 234.600 ;
        RECT 234.200 234.400 238.400 235.200 ;
        RECT 242.800 235.000 243.600 239.800 ;
        RECT 246.000 235.000 246.800 239.800 ;
        RECT 234.200 234.000 234.800 234.400 ;
        RECT 233.200 233.200 234.800 234.000 ;
        RECT 237.800 233.800 243.600 234.400 ;
        RECT 235.800 233.200 237.200 233.800 ;
        RECT 235.800 233.000 242.000 233.200 ;
        RECT 236.600 232.600 242.000 233.000 ;
        RECT 241.200 232.400 242.000 232.600 ;
        RECT 243.000 233.000 243.600 233.800 ;
        RECT 244.200 233.600 246.800 234.400 ;
        RECT 249.200 233.600 250.000 239.800 ;
        RECT 250.800 237.000 251.600 239.800 ;
        RECT 252.400 237.000 253.200 239.800 ;
        RECT 254.000 237.000 254.800 239.800 ;
        RECT 252.400 234.400 256.600 235.200 ;
        RECT 257.200 234.400 258.000 239.800 ;
        RECT 260.400 235.200 261.200 239.800 ;
        RECT 260.400 234.600 263.000 235.200 ;
        RECT 257.200 233.600 259.800 234.400 ;
        RECT 250.800 233.000 251.600 233.200 ;
        RECT 243.000 232.400 251.600 233.000 ;
        RECT 254.000 233.000 254.800 233.200 ;
        RECT 262.400 233.000 263.000 234.600 ;
        RECT 254.000 232.400 263.000 233.000 ;
        RECT 262.400 230.600 263.000 232.400 ;
        RECT 263.600 232.000 264.400 239.800 ;
        RECT 263.600 231.200 264.600 232.000 ;
        RECT 266.800 231.600 267.600 233.200 ;
        RECT 233.000 230.000 256.400 230.600 ;
        RECT 262.400 230.000 263.200 230.600 ;
        RECT 233.000 229.800 233.800 230.000 ;
        RECT 238.000 229.600 238.800 230.000 ;
        RECT 244.400 229.600 245.200 230.000 ;
        RECT 255.600 229.400 256.400 230.000 ;
        RECT 231.600 228.200 240.400 229.000 ;
        RECT 241.000 228.600 243.000 229.400 ;
        RECT 246.800 228.600 250.000 229.400 ;
        RECT 225.200 226.800 229.200 227.600 ;
        RECT 220.400 222.200 221.200 226.000 ;
        RECT 225.200 222.200 226.000 226.800 ;
        RECT 228.400 222.200 229.200 226.800 ;
        RECT 231.600 222.200 232.400 228.200 ;
        RECT 234.000 226.800 237.000 227.600 ;
        RECT 236.200 226.200 237.000 226.800 ;
        RECT 242.200 226.200 243.000 228.600 ;
        RECT 244.400 226.800 245.200 228.400 ;
        RECT 249.600 227.800 250.400 228.000 ;
        RECT 246.000 227.200 250.400 227.800 ;
        RECT 246.000 227.000 246.800 227.200 ;
        RECT 252.400 226.400 253.200 229.200 ;
        RECT 258.200 228.600 262.000 229.400 ;
        RECT 258.200 227.400 259.000 228.600 ;
        RECT 262.600 228.000 263.200 230.000 ;
        RECT 246.000 226.200 246.800 226.400 ;
        RECT 236.200 225.400 238.800 226.200 ;
        RECT 242.200 225.600 246.800 226.200 ;
        RECT 247.600 225.600 249.200 226.400 ;
        RECT 252.200 225.600 253.200 226.400 ;
        RECT 257.200 226.800 259.000 227.400 ;
        RECT 262.000 227.400 263.200 228.000 ;
        RECT 257.200 226.200 258.000 226.800 ;
        RECT 238.000 222.200 238.800 225.400 ;
        RECT 255.600 225.400 258.000 226.200 ;
        RECT 239.600 222.200 240.400 225.000 ;
        RECT 241.200 222.200 242.000 225.000 ;
        RECT 242.800 222.200 243.600 225.000 ;
        RECT 246.000 222.200 246.800 225.000 ;
        RECT 249.200 222.200 250.000 225.000 ;
        RECT 250.800 222.200 251.600 225.000 ;
        RECT 252.400 222.200 253.200 225.000 ;
        RECT 254.000 222.200 254.800 225.000 ;
        RECT 255.600 222.200 256.400 225.400 ;
        RECT 262.000 222.200 262.800 227.400 ;
        RECT 263.800 226.800 264.600 231.200 ;
        RECT 265.200 230.300 266.000 230.400 ;
        RECT 268.400 230.300 269.200 239.800 ;
        RECT 271.600 231.600 272.400 233.200 ;
        RECT 265.200 229.700 269.200 230.300 ;
        RECT 265.200 229.600 266.000 229.700 ;
        RECT 263.600 226.000 264.600 226.800 ;
        RECT 268.400 226.200 269.200 229.700 ;
        RECT 270.000 228.300 270.800 228.400 ;
        RECT 273.200 228.300 274.000 239.800 ;
        RECT 276.400 230.300 277.200 230.400 ;
        RECT 278.000 230.300 278.800 239.800 ;
        RECT 280.400 233.600 281.200 234.400 ;
        RECT 280.400 232.400 281.000 233.600 ;
        RECT 281.800 232.400 282.600 239.800 ;
        RECT 279.600 231.800 281.000 232.400 ;
        RECT 281.600 231.800 282.600 232.400 ;
        RECT 279.600 231.600 280.400 231.800 ;
        RECT 276.400 229.700 278.800 230.300 ;
        RECT 276.400 229.600 277.200 229.700 ;
        RECT 270.000 227.700 274.000 228.300 ;
        RECT 270.000 226.800 270.800 227.700 ;
        RECT 273.200 226.200 274.000 227.700 ;
        RECT 274.800 228.300 275.600 228.400 ;
        RECT 276.400 228.300 277.200 228.400 ;
        RECT 274.800 227.700 277.200 228.300 ;
        RECT 274.800 226.800 275.600 227.700 ;
        RECT 276.400 226.800 277.200 227.700 ;
        RECT 263.600 222.200 264.400 226.000 ;
        RECT 267.400 225.600 269.200 226.200 ;
        RECT 272.200 225.600 274.000 226.200 ;
        RECT 267.400 222.200 268.200 225.600 ;
        RECT 272.200 222.200 273.000 225.600 ;
        RECT 278.000 222.200 278.800 229.700 ;
        RECT 281.600 228.400 282.200 231.800 ;
        RECT 282.800 228.800 283.600 230.400 ;
        RECT 279.600 227.600 282.200 228.400 ;
        RECT 284.400 228.200 285.200 228.400 ;
        RECT 283.600 227.600 285.200 228.200 ;
        RECT 279.800 226.200 280.400 227.600 ;
        RECT 283.600 227.200 284.400 227.600 ;
        RECT 281.400 226.200 285.000 226.600 ;
        RECT 279.600 222.200 280.400 226.200 ;
        RECT 281.200 226.000 285.200 226.200 ;
        RECT 281.200 222.200 282.000 226.000 ;
        RECT 284.400 222.200 285.200 226.000 ;
        RECT 286.000 222.200 286.800 239.800 ;
        RECT 290.000 233.600 290.800 234.400 ;
        RECT 290.000 232.400 290.600 233.600 ;
        RECT 291.400 232.400 292.200 239.800 ;
        RECT 298.200 232.400 299.000 239.800 ;
        RECT 299.600 233.600 300.400 234.400 ;
        RECT 299.800 232.400 300.400 233.600 ;
        RECT 289.200 231.800 290.600 232.400 ;
        RECT 291.200 231.800 292.200 232.400 ;
        RECT 289.200 231.600 290.000 231.800 ;
        RECT 287.600 230.300 288.400 230.400 ;
        RECT 291.200 230.300 291.800 231.800 ;
        RECT 297.200 231.600 299.200 232.400 ;
        RECT 299.800 231.800 301.200 232.400 ;
        RECT 300.400 231.600 301.200 231.800 ;
        RECT 287.600 229.700 291.800 230.300 ;
        RECT 287.600 229.600 288.400 229.700 ;
        RECT 291.200 228.400 291.800 229.700 ;
        RECT 292.400 230.300 293.200 230.400 ;
        RECT 295.600 230.300 296.400 230.400 ;
        RECT 292.400 229.700 296.400 230.300 ;
        RECT 292.400 228.800 293.200 229.700 ;
        RECT 295.600 229.600 296.400 229.700 ;
        RECT 297.200 228.800 298.000 230.400 ;
        RECT 298.600 228.400 299.200 231.600 ;
        RECT 289.200 227.600 291.800 228.400 ;
        RECT 294.000 228.200 294.800 228.400 ;
        RECT 293.200 227.600 294.800 228.200 ;
        RECT 295.600 228.200 296.400 228.400 ;
        RECT 295.600 227.600 297.200 228.200 ;
        RECT 298.600 227.600 301.200 228.400 ;
        RECT 287.600 224.800 288.400 226.400 ;
        RECT 289.400 226.200 290.000 227.600 ;
        RECT 293.200 227.200 294.000 227.600 ;
        RECT 296.400 227.200 297.200 227.600 ;
        RECT 291.000 226.200 294.600 226.600 ;
        RECT 295.800 226.200 299.400 226.600 ;
        RECT 300.400 226.200 301.000 227.600 ;
        RECT 302.000 226.800 302.800 228.400 ;
        RECT 303.600 226.200 304.400 239.800 ;
        RECT 305.200 231.600 306.000 233.200 ;
        RECT 314.200 232.400 315.000 239.800 ;
        RECT 319.600 235.800 320.400 239.800 ;
        RECT 319.800 235.600 320.400 235.800 ;
        RECT 322.800 235.800 323.600 239.800 ;
        RECT 322.800 235.600 323.400 235.800 ;
        RECT 319.800 235.000 323.400 235.600 ;
        RECT 315.600 233.600 316.400 234.400 ;
        RECT 315.800 232.400 316.400 233.600 ;
        RECT 321.200 232.800 322.000 234.400 ;
        RECT 322.800 232.400 323.400 235.000 ;
        RECT 313.200 231.600 315.200 232.400 ;
        RECT 315.800 231.800 317.200 232.400 ;
        RECT 316.400 231.600 317.200 231.800 ;
        RECT 311.600 230.300 312.400 230.400 ;
        RECT 313.200 230.300 314.000 230.400 ;
        RECT 311.600 229.700 314.000 230.300 ;
        RECT 311.600 229.600 312.400 229.700 ;
        RECT 313.200 228.800 314.000 229.700 ;
        RECT 314.600 228.400 315.200 231.600 ;
        RECT 318.000 230.800 318.800 232.400 ;
        RECT 322.800 231.600 323.600 232.400 ;
        RECT 319.600 229.600 321.200 230.400 ;
        RECT 322.800 228.400 323.400 231.600 ;
        RECT 326.000 231.200 326.800 239.800 ;
        RECT 329.200 231.200 330.000 239.800 ;
        RECT 332.400 231.200 333.200 239.800 ;
        RECT 335.600 231.200 336.400 239.800 ;
        RECT 340.400 235.800 341.200 239.800 ;
        RECT 340.600 235.600 341.200 235.800 ;
        RECT 343.600 235.800 344.400 239.800 ;
        RECT 346.800 235.800 347.600 239.800 ;
        RECT 343.600 235.600 344.200 235.800 ;
        RECT 340.600 235.000 344.200 235.600 ;
        RECT 347.000 235.600 347.600 235.800 ;
        RECT 350.000 235.800 350.800 239.800 ;
        RECT 350.000 235.600 350.600 235.800 ;
        RECT 353.200 235.600 354.000 239.800 ;
        RECT 356.400 235.800 357.200 239.800 ;
        RECT 356.400 235.600 357.000 235.800 ;
        RECT 347.000 235.000 350.600 235.600 ;
        RECT 353.400 235.000 357.000 235.600 ;
        RECT 342.000 232.800 342.800 234.400 ;
        RECT 343.600 232.400 344.200 235.000 ;
        RECT 348.400 232.800 349.200 234.400 ;
        RECT 350.000 232.400 350.600 235.000 ;
        RECT 351.600 234.300 352.400 234.400 ;
        RECT 354.800 234.300 355.600 234.400 ;
        RECT 351.600 233.700 355.600 234.300 ;
        RECT 351.600 233.600 352.400 233.700 ;
        RECT 354.800 232.800 355.600 233.700 ;
        RECT 356.400 232.400 357.000 235.000 ;
        RECT 358.000 235.000 358.800 239.000 ;
        RECT 311.600 228.200 312.400 228.400 ;
        RECT 311.600 227.600 313.200 228.200 ;
        RECT 314.600 227.600 317.200 228.400 ;
        RECT 321.800 228.200 323.400 228.400 ;
        RECT 321.600 227.800 323.400 228.200 ;
        RECT 324.400 230.400 326.800 231.200 ;
        RECT 327.800 230.400 330.000 231.200 ;
        RECT 331.000 230.400 333.200 231.200 ;
        RECT 334.600 230.400 336.400 231.200 ;
        RECT 338.800 230.800 339.600 232.400 ;
        RECT 343.600 231.600 344.400 232.400 ;
        RECT 345.200 232.300 346.000 232.400 ;
        RECT 346.800 232.300 347.600 232.400 ;
        RECT 345.200 231.700 347.600 232.300 ;
        RECT 312.400 227.200 313.200 227.600 ;
        RECT 311.800 226.200 315.400 226.600 ;
        RECT 316.400 226.200 317.000 227.600 ;
        RECT 289.200 222.200 290.000 226.200 ;
        RECT 290.800 226.000 294.800 226.200 ;
        RECT 290.800 222.200 291.600 226.000 ;
        RECT 294.000 222.200 294.800 226.000 ;
        RECT 295.600 226.000 299.600 226.200 ;
        RECT 295.600 222.200 296.400 226.000 ;
        RECT 298.800 222.200 299.600 226.000 ;
        RECT 300.400 222.200 301.200 226.200 ;
        RECT 303.600 225.600 305.400 226.200 ;
        RECT 304.600 222.200 305.400 225.600 ;
        RECT 311.600 226.000 315.600 226.200 ;
        RECT 311.600 222.200 312.400 226.000 ;
        RECT 314.800 222.200 315.600 226.000 ;
        RECT 316.400 222.200 317.200 226.200 ;
        RECT 321.600 222.200 322.400 227.800 ;
        RECT 324.400 227.600 325.200 230.400 ;
        RECT 327.800 229.000 328.600 230.400 ;
        RECT 331.000 229.000 331.800 230.400 ;
        RECT 334.600 229.000 335.400 230.400 ;
        RECT 340.400 229.600 342.000 230.400 ;
        RECT 326.000 228.200 328.600 229.000 ;
        RECT 329.400 228.200 331.800 229.000 ;
        RECT 332.800 228.200 335.400 229.000 ;
        RECT 336.200 228.200 338.000 229.000 ;
        RECT 343.600 228.400 344.200 231.600 ;
        RECT 345.200 230.800 346.000 231.700 ;
        RECT 346.800 231.600 347.600 231.700 ;
        RECT 350.000 231.600 350.800 232.400 ;
        RECT 346.800 229.600 348.400 230.400 ;
        RECT 350.000 228.400 350.600 231.600 ;
        RECT 351.600 230.800 352.400 232.400 ;
        RECT 356.400 231.600 357.200 232.400 ;
        RECT 358.000 231.600 358.600 235.000 ;
        RECT 362.200 232.800 363.000 239.800 ;
        RECT 369.200 236.400 370.000 239.800 ;
        RECT 369.000 235.800 370.000 236.400 ;
        RECT 369.000 235.200 369.600 235.800 ;
        RECT 372.400 235.200 373.200 239.800 ;
        RECT 375.600 237.000 376.400 239.800 ;
        RECT 377.200 237.000 378.000 239.800 ;
        RECT 367.600 234.600 369.600 235.200 ;
        RECT 362.200 232.200 363.800 232.800 ;
        RECT 353.200 229.600 354.800 230.400 ;
        RECT 356.400 228.400 357.000 231.600 ;
        RECT 358.000 231.000 361.800 231.600 ;
        RECT 358.000 228.800 358.800 230.400 ;
        RECT 359.600 228.800 360.400 230.400 ;
        RECT 361.200 229.000 361.800 231.000 ;
        RECT 342.600 228.200 344.200 228.400 ;
        RECT 327.800 227.600 328.600 228.200 ;
        RECT 331.000 227.600 331.800 228.200 ;
        RECT 334.600 227.600 335.400 228.200 ;
        RECT 337.200 227.600 338.000 228.200 ;
        RECT 342.400 227.800 344.200 228.200 ;
        RECT 348.400 227.800 350.600 228.400 ;
        RECT 355.400 228.200 357.000 228.400 ;
        RECT 355.200 227.800 357.000 228.200 ;
        RECT 361.200 228.200 362.600 229.000 ;
        RECT 363.200 228.400 363.800 232.200 ;
        RECT 364.400 229.600 365.200 231.200 ;
        RECT 367.600 229.000 368.400 234.600 ;
        RECT 370.200 234.400 374.400 235.200 ;
        RECT 378.800 235.000 379.600 239.800 ;
        RECT 382.000 235.000 382.800 239.800 ;
        RECT 370.200 234.000 370.800 234.400 ;
        RECT 369.200 233.200 370.800 234.000 ;
        RECT 373.800 233.800 379.600 234.400 ;
        RECT 371.800 233.200 373.200 233.800 ;
        RECT 371.800 233.000 378.000 233.200 ;
        RECT 372.600 232.600 378.000 233.000 ;
        RECT 377.200 232.400 378.000 232.600 ;
        RECT 379.000 233.000 379.600 233.800 ;
        RECT 380.200 233.600 382.800 234.400 ;
        RECT 385.200 233.600 386.000 239.800 ;
        RECT 386.800 237.000 387.600 239.800 ;
        RECT 388.400 237.000 389.200 239.800 ;
        RECT 390.000 237.000 390.800 239.800 ;
        RECT 388.400 234.400 392.600 235.200 ;
        RECT 393.200 234.400 394.000 239.800 ;
        RECT 396.400 235.200 397.200 239.800 ;
        RECT 396.400 234.600 399.000 235.200 ;
        RECT 393.200 233.600 395.800 234.400 ;
        RECT 386.800 233.000 387.600 233.200 ;
        RECT 379.000 232.400 387.600 233.000 ;
        RECT 390.000 233.000 390.800 233.200 ;
        RECT 398.400 233.000 399.000 234.600 ;
        RECT 390.000 232.400 399.000 233.000 ;
        RECT 398.400 230.600 399.000 232.400 ;
        RECT 399.600 232.000 400.400 239.800 ;
        RECT 399.600 231.200 400.600 232.000 ;
        RECT 369.000 230.000 392.400 230.600 ;
        RECT 398.400 230.000 399.200 230.600 ;
        RECT 369.000 229.800 369.800 230.000 ;
        RECT 370.800 229.600 371.600 230.000 ;
        RECT 374.000 229.600 374.800 230.000 ;
        RECT 391.600 229.400 392.400 230.000 ;
        RECT 363.200 228.300 365.200 228.400 ;
        RECT 366.000 228.300 366.800 228.400 ;
        RECT 361.200 227.800 362.200 228.200 ;
        RECT 324.400 226.800 326.800 227.600 ;
        RECT 327.800 226.800 330.000 227.600 ;
        RECT 331.000 226.800 333.200 227.600 ;
        RECT 334.600 226.800 336.400 227.600 ;
        RECT 326.000 222.200 326.800 226.800 ;
        RECT 329.200 222.200 330.000 226.800 ;
        RECT 332.400 222.200 333.200 226.800 ;
        RECT 335.600 222.200 336.400 226.800 ;
        RECT 342.400 222.200 343.200 227.800 ;
        RECT 348.400 227.600 349.600 227.800 ;
        RECT 348.800 222.200 349.600 227.600 ;
        RECT 355.200 222.200 356.000 227.800 ;
        RECT 358.000 227.200 362.200 227.800 ;
        RECT 363.200 227.700 366.800 228.300 ;
        RECT 363.200 227.600 365.200 227.700 ;
        RECT 366.000 227.600 366.800 227.700 ;
        RECT 367.600 228.200 376.400 229.000 ;
        RECT 377.000 228.600 379.000 229.400 ;
        RECT 382.800 228.600 386.000 229.400 ;
        RECT 358.000 225.000 358.600 227.200 ;
        RECT 363.200 227.000 363.800 227.600 ;
        RECT 363.000 226.600 363.800 227.000 ;
        RECT 362.200 226.000 363.800 226.600 ;
        RECT 358.000 223.000 358.800 225.000 ;
        RECT 362.200 223.000 363.000 226.000 ;
        RECT 367.600 222.200 368.400 228.200 ;
        RECT 370.000 226.800 373.000 227.600 ;
        RECT 372.200 226.200 373.000 226.800 ;
        RECT 378.200 226.200 379.000 228.600 ;
        RECT 380.400 226.800 381.200 228.400 ;
        RECT 385.600 227.800 386.400 228.000 ;
        RECT 382.000 227.200 386.400 227.800 ;
        RECT 382.000 227.000 382.800 227.200 ;
        RECT 388.400 226.400 389.200 229.200 ;
        RECT 394.200 228.600 398.000 229.400 ;
        RECT 394.200 227.400 395.000 228.600 ;
        RECT 398.600 228.000 399.200 230.000 ;
        RECT 382.000 226.200 382.800 226.400 ;
        RECT 372.200 225.400 374.800 226.200 ;
        RECT 378.200 225.600 382.800 226.200 ;
        RECT 383.600 225.600 385.200 226.400 ;
        RECT 388.200 225.600 389.200 226.400 ;
        RECT 393.200 226.800 395.000 227.400 ;
        RECT 398.000 227.400 399.200 228.000 ;
        RECT 393.200 226.200 394.000 226.800 ;
        RECT 374.000 222.200 374.800 225.400 ;
        RECT 391.600 225.400 394.000 226.200 ;
        RECT 375.600 222.200 376.400 225.000 ;
        RECT 377.200 222.200 378.000 225.000 ;
        RECT 378.800 222.200 379.600 225.000 ;
        RECT 382.000 222.200 382.800 225.000 ;
        RECT 385.200 222.200 386.000 225.000 ;
        RECT 386.800 222.200 387.600 225.000 ;
        RECT 388.400 222.200 389.200 225.000 ;
        RECT 390.000 222.200 390.800 225.000 ;
        RECT 391.600 222.200 392.400 225.400 ;
        RECT 398.000 222.200 398.800 227.400 ;
        RECT 399.800 226.800 400.600 231.200 ;
        RECT 401.200 230.300 402.000 230.400 ;
        RECT 402.800 230.300 403.600 239.800 ;
        RECT 406.000 231.600 406.800 233.200 ;
        RECT 401.200 229.700 403.600 230.300 ;
        RECT 401.200 229.600 402.000 229.700 ;
        RECT 399.600 226.000 400.600 226.800 ;
        RECT 399.600 222.200 400.400 226.000 ;
        RECT 402.800 222.200 403.600 229.700 ;
        RECT 404.400 224.800 405.200 226.400 ;
        RECT 407.600 226.200 408.400 239.800 ;
        RECT 410.800 232.400 411.600 239.800 ;
        RECT 414.000 232.800 414.800 239.800 ;
        RECT 410.800 231.800 413.400 232.400 ;
        RECT 414.000 231.800 415.000 232.800 ;
        RECT 412.800 229.800 413.400 231.800 ;
        RECT 412.800 229.000 413.800 229.800 ;
        RECT 409.200 226.800 410.000 228.400 ;
        RECT 412.800 227.400 413.400 229.000 ;
        RECT 414.400 228.400 415.000 231.800 ;
        RECT 418.800 231.200 419.600 239.800 ;
        RECT 422.000 231.200 422.800 239.800 ;
        RECT 425.200 231.200 426.000 239.800 ;
        RECT 428.400 231.200 429.200 239.800 ;
        RECT 417.200 230.400 419.600 231.200 ;
        RECT 420.600 230.400 422.800 231.200 ;
        RECT 423.800 230.400 426.000 231.200 ;
        RECT 427.400 230.400 429.200 231.200 ;
        RECT 433.200 231.200 434.000 239.800 ;
        RECT 436.400 231.200 437.200 239.800 ;
        RECT 439.600 231.200 440.400 239.800 ;
        RECT 442.800 231.200 443.600 239.800 ;
        RECT 446.000 232.400 446.800 239.800 ;
        RECT 449.200 239.200 453.200 239.800 ;
        RECT 449.200 232.400 450.000 239.200 ;
        RECT 446.000 231.800 450.000 232.400 ;
        RECT 450.800 231.800 451.600 238.600 ;
        RECT 452.400 231.800 453.200 239.200 ;
        RECT 454.000 239.200 458.000 239.800 ;
        RECT 454.000 231.800 454.800 239.200 ;
        RECT 455.600 231.800 456.400 238.600 ;
        RECT 457.200 232.400 458.000 239.200 ;
        RECT 460.400 232.400 461.200 239.800 ;
        RECT 462.000 234.300 462.800 234.400 ;
        RECT 466.800 234.300 467.600 234.400 ;
        RECT 462.000 233.700 467.600 234.300 ;
        RECT 462.000 233.600 462.800 233.700 ;
        RECT 466.800 233.600 467.600 233.700 ;
        RECT 457.200 231.800 461.200 232.400 ;
        RECT 450.800 231.200 451.400 231.800 ;
        RECT 455.800 231.200 456.400 231.800 ;
        RECT 433.200 230.400 435.000 231.200 ;
        RECT 436.400 230.400 438.600 231.200 ;
        RECT 439.600 230.400 441.800 231.200 ;
        RECT 442.800 230.400 445.200 231.200 ;
        RECT 446.800 230.400 447.600 230.800 ;
        RECT 449.400 230.600 451.400 231.200 ;
        RECT 449.400 230.400 450.000 230.600 ;
        RECT 414.000 228.300 415.000 228.400 ;
        RECT 415.600 228.300 416.400 228.400 ;
        RECT 414.000 227.700 416.400 228.300 ;
        RECT 414.000 227.600 415.000 227.700 ;
        RECT 415.600 227.600 416.400 227.700 ;
        RECT 417.200 227.600 418.000 230.400 ;
        RECT 420.600 229.000 421.400 230.400 ;
        RECT 423.800 229.000 424.600 230.400 ;
        RECT 427.400 229.000 428.200 230.400 ;
        RECT 434.200 229.000 435.000 230.400 ;
        RECT 437.800 229.000 438.600 230.400 ;
        RECT 441.000 229.000 441.800 230.400 ;
        RECT 418.800 228.200 421.400 229.000 ;
        RECT 422.200 228.200 424.600 229.000 ;
        RECT 425.600 228.200 428.200 229.000 ;
        RECT 429.000 228.300 430.800 229.000 ;
        RECT 431.600 228.300 433.400 229.000 ;
        RECT 429.000 228.200 433.400 228.300 ;
        RECT 434.200 228.200 436.800 229.000 ;
        RECT 437.800 228.200 440.200 229.000 ;
        RECT 441.000 228.200 443.600 229.000 ;
        RECT 420.600 227.600 421.400 228.200 ;
        RECT 423.800 227.600 424.600 228.200 ;
        RECT 427.400 227.600 428.200 228.200 ;
        RECT 430.000 227.700 432.400 228.200 ;
        RECT 430.000 227.600 430.800 227.700 ;
        RECT 431.600 227.600 432.400 227.700 ;
        RECT 434.200 227.600 435.000 228.200 ;
        RECT 437.800 227.600 438.600 228.200 ;
        RECT 441.000 227.600 441.800 228.200 ;
        RECT 444.400 227.600 445.200 230.400 ;
        RECT 446.000 229.800 447.600 230.400 ;
        RECT 446.000 229.600 446.800 229.800 ;
        RECT 449.200 229.600 450.000 230.400 ;
        RECT 452.400 229.600 453.200 231.200 ;
        RECT 454.000 229.600 454.800 231.200 ;
        RECT 455.800 230.600 457.800 231.200 ;
        RECT 457.200 230.400 457.800 230.600 ;
        RECT 459.600 230.400 460.400 230.800 ;
        RECT 457.200 229.600 458.000 230.400 ;
        RECT 459.600 229.800 461.200 230.400 ;
        RECT 460.400 229.600 461.200 229.800 ;
        RECT 468.400 230.300 469.200 239.800 ;
        RECT 473.200 235.800 474.000 239.800 ;
        RECT 473.400 235.600 474.000 235.800 ;
        RECT 476.400 235.800 477.200 239.800 ;
        RECT 476.400 235.600 477.000 235.800 ;
        RECT 473.400 235.000 477.000 235.600 ;
        RECT 470.000 231.600 470.800 233.200 ;
        RECT 474.800 232.800 475.600 234.400 ;
        RECT 476.400 232.400 477.000 235.000 ;
        RECT 471.600 230.800 472.400 232.400 ;
        RECT 476.400 231.600 477.200 232.400 ;
        RECT 478.000 232.300 478.800 232.400 ;
        RECT 479.600 232.300 480.400 239.800 ;
        RECT 478.000 231.700 480.400 232.300 ;
        RECT 478.000 231.600 478.800 231.700 ;
        RECT 470.000 230.300 470.800 230.400 ;
        RECT 468.400 229.700 470.800 230.300 ;
        RECT 447.600 227.600 448.400 229.200 ;
        RECT 410.800 226.800 413.400 227.400 ;
        RECT 406.600 225.600 408.400 226.200 ;
        RECT 406.600 222.200 407.400 225.600 ;
        RECT 410.800 222.200 411.600 226.800 ;
        RECT 414.400 226.200 415.000 227.600 ;
        RECT 417.200 226.800 419.600 227.600 ;
        RECT 420.600 226.800 422.800 227.600 ;
        RECT 423.800 226.800 426.000 227.600 ;
        RECT 427.400 226.800 429.200 227.600 ;
        RECT 414.000 225.600 415.000 226.200 ;
        RECT 414.000 222.200 414.800 225.600 ;
        RECT 418.800 222.200 419.600 226.800 ;
        RECT 422.000 222.200 422.800 226.800 ;
        RECT 425.200 222.200 426.000 226.800 ;
        RECT 428.400 222.200 429.200 226.800 ;
        RECT 433.200 226.800 435.000 227.600 ;
        RECT 436.400 226.800 438.600 227.600 ;
        RECT 439.600 226.800 441.800 227.600 ;
        RECT 442.800 226.800 445.200 227.600 ;
        RECT 433.200 222.200 434.000 226.800 ;
        RECT 436.400 222.200 437.200 226.800 ;
        RECT 439.600 222.200 440.400 226.800 ;
        RECT 442.800 222.200 443.600 226.800 ;
        RECT 449.400 226.200 450.000 229.600 ;
        RECT 450.600 228.800 451.400 229.600 ;
        RECT 450.800 228.400 451.400 228.800 ;
        RECT 455.800 228.800 456.600 229.600 ;
        RECT 455.800 228.400 456.400 228.800 ;
        RECT 450.800 227.600 451.600 228.400 ;
        RECT 455.600 227.600 456.400 228.400 ;
        RECT 457.200 226.200 457.800 229.600 ;
        RECT 458.800 227.600 459.600 229.200 ;
        RECT 466.800 226.800 467.600 228.400 ;
        RECT 468.400 226.200 469.200 229.700 ;
        RECT 470.000 229.600 470.800 229.700 ;
        RECT 473.200 229.600 474.800 230.400 ;
        RECT 476.400 228.400 477.000 231.600 ;
        RECT 475.400 228.200 477.000 228.400 ;
        RECT 475.200 227.800 477.000 228.200 ;
        RECT 449.000 222.200 450.600 226.200 ;
        RECT 456.600 222.200 458.200 226.200 ;
        RECT 468.400 225.600 470.200 226.200 ;
        RECT 469.400 222.200 470.200 225.600 ;
        RECT 475.200 222.200 476.000 227.800 ;
        RECT 478.000 226.800 478.800 228.400 ;
        RECT 479.600 226.200 480.400 231.700 ;
        RECT 481.200 231.600 482.000 233.200 ;
        RECT 482.800 232.400 483.600 239.800 ;
        RECT 486.000 239.200 490.000 239.800 ;
        RECT 486.000 232.400 486.800 239.200 ;
        RECT 482.800 231.800 486.800 232.400 ;
        RECT 487.600 231.800 488.400 238.600 ;
        RECT 489.200 231.800 490.000 239.200 ;
        RECT 490.800 235.800 491.600 239.800 ;
        RECT 491.000 235.600 491.600 235.800 ;
        RECT 494.000 235.800 494.800 239.800 ;
        RECT 494.000 235.600 494.600 235.800 ;
        RECT 491.000 235.000 494.600 235.600 ;
        RECT 491.000 232.400 491.600 235.000 ;
        RECT 492.400 232.800 493.200 234.400 ;
        RECT 487.600 231.200 488.200 231.800 ;
        RECT 490.800 231.600 491.600 232.400 ;
        RECT 483.600 230.400 484.400 230.800 ;
        RECT 486.200 230.600 488.200 231.200 ;
        RECT 486.200 230.400 486.800 230.600 ;
        RECT 482.800 229.800 484.400 230.400 ;
        RECT 482.800 229.600 483.600 229.800 ;
        RECT 486.000 229.600 486.800 230.400 ;
        RECT 489.200 229.600 490.000 231.200 ;
        RECT 481.200 228.300 482.000 228.400 ;
        RECT 484.400 228.300 485.200 229.200 ;
        RECT 481.200 227.700 485.200 228.300 ;
        RECT 481.200 227.600 482.000 227.700 ;
        RECT 484.400 227.600 485.200 227.700 ;
        RECT 486.200 226.200 486.800 229.600 ;
        RECT 487.400 228.800 488.200 229.600 ;
        RECT 487.600 228.400 488.200 228.800 ;
        RECT 491.000 228.400 491.600 231.600 ;
        RECT 495.600 230.800 496.400 232.400 ;
        RECT 497.200 231.800 498.000 239.800 ;
        RECT 498.800 232.400 499.600 239.800 ;
        RECT 502.000 232.400 502.800 239.800 ;
        RECT 503.600 235.800 504.400 239.800 ;
        RECT 503.800 235.600 504.400 235.800 ;
        RECT 506.800 235.600 507.600 239.800 ;
        RECT 510.000 235.800 510.800 239.800 ;
        RECT 510.200 235.600 510.800 235.800 ;
        RECT 513.200 235.800 514.000 239.800 ;
        RECT 518.000 235.800 518.800 239.800 ;
        RECT 513.200 235.600 513.800 235.800 ;
        RECT 503.800 235.000 507.400 235.600 ;
        RECT 510.200 235.000 513.800 235.600 ;
        RECT 518.200 235.600 518.800 235.800 ;
        RECT 521.200 235.800 522.000 239.800 ;
        RECT 524.400 235.800 525.200 239.800 ;
        RECT 521.200 235.600 521.800 235.800 ;
        RECT 518.200 235.000 521.800 235.600 ;
        RECT 524.600 235.600 525.200 235.800 ;
        RECT 527.600 235.800 528.400 239.800 ;
        RECT 527.600 235.600 528.200 235.800 ;
        RECT 530.800 235.600 531.600 239.800 ;
        RECT 534.000 235.800 534.800 239.800 ;
        RECT 535.600 235.800 536.400 239.800 ;
        RECT 534.000 235.600 534.600 235.800 ;
        RECT 524.600 235.000 528.200 235.600 ;
        RECT 531.000 235.000 534.600 235.600 ;
        RECT 503.800 232.400 504.400 235.000 ;
        RECT 505.200 234.300 506.000 234.400 ;
        RECT 508.400 234.300 509.200 234.400 ;
        RECT 505.200 233.700 509.200 234.300 ;
        RECT 505.200 232.800 506.000 233.700 ;
        RECT 508.400 233.600 509.200 233.700 ;
        RECT 510.200 232.400 510.800 235.000 ;
        RECT 511.600 232.800 512.400 234.400 ;
        RECT 519.600 232.800 520.400 234.400 ;
        RECT 521.200 232.400 521.800 235.000 ;
        RECT 526.000 232.800 526.800 234.400 ;
        RECT 527.600 232.400 528.200 235.000 ;
        RECT 530.800 234.300 531.600 234.400 ;
        RECT 532.400 234.300 533.200 234.400 ;
        RECT 530.800 233.700 533.200 234.300 ;
        RECT 530.800 233.600 531.600 233.700 ;
        RECT 532.400 232.800 533.200 233.700 ;
        RECT 534.000 232.400 534.600 235.000 ;
        RECT 535.800 235.600 536.400 235.800 ;
        RECT 538.800 235.800 539.600 239.800 ;
        RECT 542.000 235.800 542.800 239.800 ;
        RECT 538.800 235.600 539.400 235.800 ;
        RECT 535.800 235.000 539.400 235.600 ;
        RECT 542.200 235.600 542.800 235.800 ;
        RECT 545.200 235.800 546.000 239.800 ;
        RECT 545.200 235.600 545.800 235.800 ;
        RECT 542.200 235.000 545.800 235.600 ;
        RECT 535.800 232.400 536.400 235.000 ;
        RECT 537.200 232.800 538.000 234.400 ;
        RECT 542.200 232.400 542.800 235.000 ;
        RECT 543.600 232.800 544.400 234.400 ;
        RECT 498.800 231.800 502.800 232.400 ;
        RECT 497.400 230.400 498.000 231.800 ;
        RECT 503.600 231.600 504.400 232.400 ;
        RECT 501.200 230.400 502.000 230.800 ;
        RECT 493.200 229.600 494.800 230.400 ;
        RECT 497.200 229.800 499.600 230.400 ;
        RECT 501.200 229.800 502.800 230.400 ;
        RECT 497.200 229.600 498.000 229.800 ;
        RECT 487.600 227.600 488.400 228.400 ;
        RECT 491.000 228.200 492.600 228.400 ;
        RECT 491.000 227.800 492.800 228.200 ;
        RECT 479.600 225.600 481.400 226.200 ;
        RECT 480.600 222.200 481.400 225.600 ;
        RECT 485.800 222.200 487.400 226.200 ;
        RECT 492.000 222.200 492.800 227.800 ;
        RECT 497.200 225.600 498.000 226.400 ;
        RECT 499.000 226.200 499.600 229.800 ;
        RECT 502.000 229.600 502.800 229.800 ;
        RECT 500.400 227.600 501.200 229.200 ;
        RECT 503.800 228.400 504.400 231.600 ;
        RECT 508.400 230.800 509.200 232.400 ;
        RECT 510.000 231.600 510.800 232.400 ;
        RECT 506.000 229.600 507.600 230.400 ;
        RECT 510.200 228.400 510.800 231.600 ;
        RECT 514.800 230.800 515.600 232.400 ;
        RECT 516.400 232.300 517.200 232.400 ;
        RECT 518.000 232.300 518.800 232.400 ;
        RECT 516.400 231.700 518.800 232.300 ;
        RECT 512.400 229.600 514.000 230.400 ;
        RECT 516.400 229.600 517.200 231.700 ;
        RECT 518.000 231.600 518.800 231.700 ;
        RECT 521.200 231.600 522.000 232.400 ;
        RECT 518.000 229.600 519.600 230.400 ;
        RECT 521.200 228.400 521.800 231.600 ;
        RECT 522.800 230.800 523.600 232.400 ;
        RECT 527.600 231.600 528.400 232.400 ;
        RECT 524.400 229.600 526.000 230.400 ;
        RECT 527.600 228.400 528.200 231.600 ;
        RECT 529.200 230.800 530.000 232.400 ;
        RECT 534.000 231.600 534.800 232.400 ;
        RECT 535.600 231.600 536.400 232.400 ;
        RECT 530.800 229.600 532.400 230.400 ;
        RECT 534.000 228.400 534.600 231.600 ;
        RECT 503.800 228.200 505.400 228.400 ;
        RECT 510.200 228.200 511.800 228.400 ;
        RECT 503.800 227.800 505.600 228.200 ;
        RECT 510.200 227.800 512.000 228.200 ;
        RECT 497.400 224.800 498.200 225.600 ;
        RECT 498.800 222.200 499.600 226.200 ;
        RECT 504.800 222.200 505.600 227.800 ;
        RECT 511.200 222.200 512.000 227.800 ;
        RECT 519.600 227.800 521.800 228.400 ;
        RECT 526.600 228.200 528.200 228.400 ;
        RECT 533.000 228.200 534.600 228.400 ;
        RECT 526.400 227.800 528.200 228.200 ;
        RECT 532.800 227.800 534.600 228.200 ;
        RECT 535.800 228.400 536.400 231.600 ;
        RECT 540.400 230.800 541.200 232.400 ;
        RECT 542.000 231.600 542.800 232.400 ;
        RECT 542.200 230.400 542.800 231.600 ;
        RECT 546.800 230.800 547.600 232.400 ;
        RECT 548.400 231.600 549.200 233.200 ;
        RECT 538.000 229.600 539.600 230.400 ;
        RECT 542.000 229.600 542.800 230.400 ;
        RECT 544.400 229.600 546.000 230.400 ;
        RECT 542.200 228.400 542.800 229.600 ;
        RECT 535.800 228.200 537.400 228.400 ;
        RECT 542.200 228.200 543.800 228.400 ;
        RECT 535.800 227.800 537.600 228.200 ;
        RECT 542.200 227.800 544.000 228.200 ;
        RECT 519.600 227.600 520.800 227.800 ;
        RECT 520.000 222.200 520.800 227.600 ;
        RECT 526.400 222.200 527.200 227.800 ;
        RECT 532.800 222.200 533.600 227.800 ;
        RECT 536.800 222.200 537.600 227.800 ;
        RECT 543.200 222.200 544.000 227.800 ;
        RECT 550.000 226.200 550.800 239.800 ;
        RECT 554.800 232.300 555.600 239.800 ;
        RECT 558.000 235.800 558.800 239.800 ;
        RECT 558.200 235.600 558.800 235.800 ;
        RECT 561.200 235.800 562.000 239.800 ;
        RECT 561.200 235.600 561.800 235.800 ;
        RECT 558.200 235.000 561.800 235.600 ;
        RECT 559.600 232.800 560.400 234.400 ;
        RECT 561.200 232.400 561.800 235.000 ;
        RECT 556.400 232.300 557.200 232.400 ;
        RECT 554.800 231.700 557.200 232.300 ;
        RECT 551.600 226.800 552.400 228.400 ;
        RECT 553.200 226.800 554.000 228.400 ;
        RECT 549.000 225.600 550.800 226.200 ;
        RECT 549.000 224.400 549.800 225.600 ;
        RECT 548.400 223.600 549.800 224.400 ;
        RECT 549.000 222.200 549.800 223.600 ;
        RECT 554.800 222.200 555.600 231.700 ;
        RECT 556.400 230.800 557.200 231.700 ;
        RECT 561.200 231.600 562.000 232.400 ;
        RECT 562.800 231.600 563.600 233.200 ;
        RECT 558.000 229.600 559.600 230.400 ;
        RECT 561.200 228.400 561.800 231.600 ;
        RECT 562.800 230.300 563.600 230.400 ;
        RECT 564.400 230.300 565.200 239.800 ;
        RECT 569.200 232.000 570.000 239.800 ;
        RECT 572.400 235.200 573.200 239.800 ;
        RECT 562.800 229.700 565.200 230.300 ;
        RECT 562.800 229.600 563.600 229.700 ;
        RECT 560.200 228.200 561.800 228.400 ;
        RECT 560.000 227.800 561.800 228.200 ;
        RECT 560.000 222.200 560.800 227.800 ;
        RECT 564.400 226.200 565.200 229.700 ;
        RECT 569.000 231.200 570.000 232.000 ;
        RECT 570.600 234.600 573.200 235.200 ;
        RECT 570.600 233.000 571.200 234.600 ;
        RECT 575.600 234.400 576.400 239.800 ;
        RECT 578.800 237.000 579.600 239.800 ;
        RECT 580.400 237.000 581.200 239.800 ;
        RECT 582.000 237.000 582.800 239.800 ;
        RECT 577.000 234.400 581.200 235.200 ;
        RECT 573.800 233.600 576.400 234.400 ;
        RECT 583.600 233.600 584.400 239.800 ;
        RECT 586.800 235.000 587.600 239.800 ;
        RECT 590.000 235.000 590.800 239.800 ;
        RECT 591.600 237.000 592.400 239.800 ;
        RECT 593.200 237.000 594.000 239.800 ;
        RECT 596.400 235.200 597.200 239.800 ;
        RECT 599.600 236.400 600.400 239.800 ;
        RECT 599.600 235.800 600.600 236.400 ;
        RECT 600.000 235.200 600.600 235.800 ;
        RECT 595.200 234.400 599.400 235.200 ;
        RECT 600.000 234.600 602.000 235.200 ;
        RECT 586.800 233.600 589.400 234.400 ;
        RECT 590.000 233.800 595.800 234.400 ;
        RECT 598.800 234.000 599.400 234.400 ;
        RECT 578.800 233.000 579.600 233.200 ;
        RECT 570.600 232.400 579.600 233.000 ;
        RECT 582.000 233.000 582.800 233.200 ;
        RECT 590.000 233.000 590.600 233.800 ;
        RECT 596.400 233.200 597.800 233.800 ;
        RECT 598.800 233.200 600.400 234.000 ;
        RECT 582.000 232.400 590.600 233.000 ;
        RECT 591.600 233.000 597.800 233.200 ;
        RECT 591.600 232.600 597.000 233.000 ;
        RECT 591.600 232.400 592.400 232.600 ;
        RECT 566.000 226.800 566.800 228.400 ;
        RECT 569.000 226.800 569.800 231.200 ;
        RECT 570.600 230.600 571.200 232.400 ;
        RECT 570.400 230.000 571.200 230.600 ;
        RECT 577.200 230.000 600.600 230.600 ;
        RECT 570.400 228.000 571.000 230.000 ;
        RECT 577.200 229.400 578.000 230.000 ;
        RECT 594.800 229.600 595.600 230.000 ;
        RECT 599.800 229.800 600.600 230.000 ;
        RECT 571.600 228.600 575.400 229.400 ;
        RECT 570.400 227.400 571.600 228.000 ;
        RECT 563.400 225.600 565.200 226.200 ;
        RECT 569.000 226.000 570.000 226.800 ;
        RECT 563.400 222.200 564.200 225.600 ;
        RECT 569.200 222.200 570.000 226.000 ;
        RECT 570.800 222.200 571.600 227.400 ;
        RECT 574.600 227.400 575.400 228.600 ;
        RECT 574.600 226.800 576.400 227.400 ;
        RECT 575.600 226.200 576.400 226.800 ;
        RECT 580.400 226.400 581.200 229.200 ;
        RECT 583.600 228.600 586.800 229.400 ;
        RECT 590.600 228.600 592.600 229.400 ;
        RECT 601.200 229.000 602.000 234.600 ;
        RECT 605.400 232.400 606.200 239.800 ;
        RECT 606.800 233.600 607.600 234.400 ;
        RECT 607.000 232.400 607.600 233.600 ;
        RECT 604.400 231.600 606.400 232.400 ;
        RECT 607.000 231.800 608.400 232.400 ;
        RECT 607.600 231.600 608.400 231.800 ;
        RECT 583.200 227.800 584.000 228.000 ;
        RECT 583.200 227.200 587.600 227.800 ;
        RECT 586.800 227.000 587.600 227.200 ;
        RECT 588.400 226.800 589.200 228.400 ;
        RECT 575.600 225.400 578.000 226.200 ;
        RECT 580.400 225.600 581.400 226.400 ;
        RECT 584.400 225.600 586.000 226.400 ;
        RECT 586.800 226.200 587.600 226.400 ;
        RECT 590.600 226.200 591.400 228.600 ;
        RECT 593.200 228.200 602.000 229.000 ;
        RECT 604.400 228.800 605.200 230.400 ;
        RECT 605.800 228.400 606.400 231.600 ;
        RECT 596.600 226.800 599.600 227.600 ;
        RECT 596.600 226.200 597.400 226.800 ;
        RECT 586.800 225.600 591.400 226.200 ;
        RECT 577.200 222.200 578.000 225.400 ;
        RECT 594.800 225.400 597.400 226.200 ;
        RECT 578.800 222.200 579.600 225.000 ;
        RECT 580.400 222.200 581.200 225.000 ;
        RECT 582.000 222.200 582.800 225.000 ;
        RECT 583.600 222.200 584.400 225.000 ;
        RECT 586.800 222.200 587.600 225.000 ;
        RECT 590.000 222.200 590.800 225.000 ;
        RECT 591.600 222.200 592.400 225.000 ;
        RECT 593.200 222.200 594.000 225.000 ;
        RECT 594.800 222.200 595.600 225.400 ;
        RECT 601.200 222.200 602.000 228.200 ;
        RECT 602.800 228.200 603.600 228.400 ;
        RECT 602.800 227.600 604.400 228.200 ;
        RECT 605.800 227.600 608.400 228.400 ;
        RECT 603.600 227.200 604.400 227.600 ;
        RECT 603.000 226.200 606.600 226.600 ;
        RECT 607.600 226.200 608.200 227.600 ;
        RECT 602.800 226.000 606.800 226.200 ;
        RECT 602.800 222.200 603.600 226.000 ;
        RECT 606.000 222.200 606.800 226.000 ;
        RECT 607.600 222.200 608.400 226.200 ;
        RECT 2.800 214.300 3.600 219.800 ;
        RECT 4.400 216.000 5.200 219.800 ;
        RECT 7.600 216.000 8.400 219.800 ;
        RECT 4.400 215.800 8.400 216.000 ;
        RECT 9.200 215.800 10.000 219.800 ;
        RECT 10.800 215.800 11.600 219.800 ;
        RECT 14.000 217.800 14.800 219.800 ;
        RECT 4.600 215.400 8.200 215.800 ;
        RECT 5.200 214.400 6.000 214.800 ;
        RECT 9.200 214.400 9.800 215.800 ;
        RECT 4.400 214.300 6.000 214.400 ;
        RECT 2.800 213.800 6.000 214.300 ;
        RECT 2.800 213.700 5.200 213.800 ;
        RECT 2.800 202.200 3.600 213.700 ;
        RECT 4.400 213.600 5.200 213.700 ;
        RECT 7.400 213.600 10.000 214.400 ;
        RECT 6.000 211.600 6.800 213.200 ;
        RECT 7.400 210.200 8.000 213.600 ;
        RECT 10.800 212.400 11.400 215.800 ;
        RECT 14.000 215.600 14.600 217.800 ;
        RECT 15.600 215.600 16.400 217.200 ;
        RECT 17.200 216.000 18.000 219.800 ;
        RECT 20.400 216.000 21.200 219.800 ;
        RECT 17.200 215.800 21.200 216.000 ;
        RECT 22.000 215.800 22.800 219.800 ;
        RECT 26.200 216.400 27.000 219.800 ;
        RECT 25.200 215.800 27.000 216.400 ;
        RECT 28.400 215.800 29.200 219.800 ;
        RECT 30.000 216.000 30.800 219.800 ;
        RECT 33.200 216.000 34.000 219.800 ;
        RECT 30.000 215.800 34.000 216.000 ;
        RECT 34.800 215.800 35.600 219.800 ;
        RECT 36.400 216.000 37.200 219.800 ;
        RECT 39.600 216.000 40.400 219.800 ;
        RECT 36.400 215.800 40.400 216.000 ;
        RECT 12.200 215.000 14.600 215.600 ;
        RECT 9.200 212.300 10.000 212.400 ;
        RECT 10.800 212.300 11.600 212.400 ;
        RECT 9.200 211.700 11.600 212.300 ;
        RECT 9.200 211.600 10.000 211.700 ;
        RECT 10.800 211.600 11.600 211.700 ;
        RECT 12.200 212.000 12.800 215.000 ;
        RECT 13.800 213.600 14.800 214.400 ;
        RECT 15.700 214.300 16.300 215.600 ;
        RECT 17.400 215.400 21.000 215.800 ;
        RECT 18.000 214.400 18.800 214.800 ;
        RECT 22.000 214.400 22.600 215.800 ;
        RECT 17.200 214.300 18.800 214.400 ;
        RECT 15.700 213.800 18.800 214.300 ;
        RECT 15.700 213.700 18.000 213.800 ;
        RECT 17.200 213.600 18.000 213.700 ;
        RECT 20.200 213.600 22.800 214.400 ;
        RECT 23.600 213.600 24.400 215.200 ;
        RECT 13.600 212.800 14.400 213.600 ;
        RECT 9.200 210.200 10.000 210.400 ;
        RECT 7.000 209.600 8.000 210.200 ;
        RECT 8.600 209.600 10.000 210.200 ;
        RECT 10.800 210.200 11.400 211.600 ;
        RECT 12.200 211.400 13.000 212.000 ;
        RECT 18.800 211.600 19.600 213.200 ;
        RECT 12.200 211.200 16.400 211.400 ;
        RECT 12.400 210.800 16.400 211.200 ;
        RECT 10.800 209.600 12.200 210.200 ;
        RECT 7.000 204.400 7.800 209.600 ;
        RECT 8.600 208.400 9.200 209.600 ;
        RECT 8.400 207.600 9.200 208.400 ;
        RECT 6.000 203.600 7.800 204.400 ;
        RECT 7.000 202.200 7.800 203.600 ;
        RECT 11.400 202.200 12.200 209.600 ;
        RECT 15.600 202.200 16.400 210.800 ;
        RECT 20.200 210.400 20.800 213.600 ;
        RECT 18.800 209.600 20.800 210.400 ;
        RECT 22.000 210.200 22.800 210.400 ;
        RECT 21.400 209.600 22.800 210.200 ;
        RECT 19.800 202.200 20.600 209.600 ;
        RECT 21.400 208.400 22.000 209.600 ;
        RECT 21.200 207.600 22.000 208.400 ;
        RECT 25.200 202.200 26.000 215.800 ;
        RECT 28.600 214.400 29.200 215.800 ;
        RECT 30.200 215.400 33.800 215.800 ;
        RECT 32.400 214.400 33.200 214.800 ;
        RECT 35.000 214.400 35.600 215.800 ;
        RECT 36.600 215.400 40.200 215.800 ;
        RECT 42.800 215.200 43.600 219.800 ;
        RECT 46.000 215.200 46.800 219.800 ;
        RECT 49.200 215.200 50.000 219.800 ;
        RECT 52.400 215.200 53.200 219.800 ;
        RECT 38.800 214.400 39.600 214.800 ;
        RECT 41.200 214.400 43.600 215.200 ;
        RECT 44.600 214.400 46.800 215.200 ;
        RECT 47.800 214.400 50.000 215.200 ;
        RECT 51.400 214.400 53.200 215.200 ;
        RECT 57.200 215.200 58.000 219.800 ;
        RECT 60.400 215.200 61.200 219.800 ;
        RECT 63.600 215.200 64.400 219.800 ;
        RECT 66.800 215.200 67.600 219.800 ;
        RECT 73.800 216.400 74.600 219.000 ;
        RECT 78.000 217.000 78.800 219.000 ;
        RECT 73.800 216.000 75.600 216.400 ;
        RECT 73.000 215.600 75.600 216.000 ;
        RECT 73.000 215.400 74.600 215.600 ;
        RECT 57.200 214.400 59.000 215.200 ;
        RECT 60.400 214.400 62.600 215.200 ;
        RECT 63.600 214.400 65.800 215.200 ;
        RECT 66.800 214.400 69.200 215.200 ;
        RECT 73.000 215.000 73.800 215.400 ;
        RECT 73.000 214.400 73.600 215.000 ;
        RECT 78.200 214.800 78.800 217.000 ;
        RECT 28.400 213.600 31.000 214.400 ;
        RECT 32.400 213.800 34.000 214.400 ;
        RECT 33.200 213.600 34.000 213.800 ;
        RECT 34.800 213.600 37.400 214.400 ;
        RECT 38.800 213.800 40.400 214.400 ;
        RECT 39.600 213.600 40.400 213.800 ;
        RECT 30.400 212.400 31.000 213.600 ;
        RECT 30.000 211.600 31.000 212.400 ;
        RECT 31.600 212.300 32.400 213.200 ;
        RECT 34.800 212.300 35.600 212.400 ;
        RECT 31.600 211.700 35.600 212.300 ;
        RECT 31.600 211.600 32.400 211.700 ;
        RECT 34.800 211.600 35.600 211.700 ;
        RECT 26.800 208.800 27.600 210.400 ;
        RECT 28.400 210.200 29.200 210.400 ;
        RECT 30.400 210.200 31.000 211.600 ;
        RECT 34.800 210.200 35.600 210.400 ;
        RECT 36.800 210.200 37.400 213.600 ;
        RECT 38.000 211.600 38.800 213.200 ;
        RECT 41.200 211.600 42.000 214.400 ;
        RECT 44.600 213.800 45.400 214.400 ;
        RECT 47.800 213.800 48.600 214.400 ;
        RECT 51.400 213.800 52.200 214.400 ;
        RECT 54.000 214.300 54.800 214.400 ;
        RECT 55.600 214.300 56.400 214.400 ;
        RECT 54.000 213.800 56.400 214.300 ;
        RECT 58.200 213.800 59.000 214.400 ;
        RECT 61.800 213.800 62.600 214.400 ;
        RECT 65.000 213.800 65.800 214.400 ;
        RECT 42.800 213.000 45.400 213.800 ;
        RECT 46.200 213.000 48.600 213.800 ;
        RECT 49.600 213.000 52.200 213.800 ;
        RECT 53.000 213.700 57.400 213.800 ;
        RECT 53.000 213.000 54.800 213.700 ;
        RECT 55.600 213.000 57.400 213.700 ;
        RECT 58.200 213.000 60.800 213.800 ;
        RECT 61.800 213.000 64.200 213.800 ;
        RECT 65.000 213.000 67.600 213.800 ;
        RECT 44.600 211.600 45.400 213.000 ;
        RECT 47.800 211.600 48.600 213.000 ;
        RECT 51.400 211.600 52.200 213.000 ;
        RECT 58.200 211.600 59.000 213.000 ;
        RECT 61.800 211.600 62.600 213.000 ;
        RECT 65.000 211.600 65.800 213.000 ;
        RECT 68.400 211.600 69.200 214.400 ;
        RECT 71.600 213.600 73.600 214.400 ;
        RECT 74.600 214.200 78.800 214.800 ;
        RECT 79.600 215.400 80.400 219.800 ;
        RECT 83.800 218.400 85.000 219.800 ;
        RECT 83.800 217.800 85.200 218.400 ;
        RECT 88.400 217.800 89.200 219.800 ;
        RECT 92.800 218.400 93.600 219.800 ;
        RECT 92.800 217.800 94.800 218.400 ;
        RECT 84.400 217.000 85.200 217.800 ;
        RECT 88.600 217.200 89.200 217.800 ;
        RECT 88.600 216.600 91.400 217.200 ;
        RECT 90.600 216.400 91.400 216.600 ;
        RECT 92.400 215.600 93.200 217.200 ;
        RECT 94.000 217.000 94.800 217.800 ;
        RECT 82.600 215.400 83.400 215.600 ;
        RECT 79.600 214.800 83.400 215.400 ;
        RECT 74.600 213.800 75.600 214.200 ;
        RECT 41.200 210.800 43.600 211.600 ;
        RECT 44.600 210.800 46.800 211.600 ;
        RECT 47.800 210.800 50.000 211.600 ;
        RECT 51.400 210.800 53.200 211.600 ;
        RECT 28.400 209.600 29.800 210.200 ;
        RECT 30.400 209.600 31.400 210.200 ;
        RECT 34.800 209.600 36.200 210.200 ;
        RECT 36.800 209.600 37.800 210.200 ;
        RECT 29.200 208.400 29.800 209.600 ;
        RECT 29.200 207.600 30.000 208.400 ;
        RECT 30.600 202.200 31.400 209.600 ;
        RECT 35.600 208.400 36.200 209.600 ;
        RECT 35.600 207.600 36.400 208.400 ;
        RECT 37.000 204.400 37.800 209.600 ;
        RECT 37.000 203.600 38.800 204.400 ;
        RECT 37.000 202.200 37.800 203.600 ;
        RECT 42.800 202.200 43.600 210.800 ;
        RECT 46.000 202.200 46.800 210.800 ;
        RECT 49.200 202.200 50.000 210.800 ;
        RECT 52.400 202.200 53.200 210.800 ;
        RECT 57.200 210.800 59.000 211.600 ;
        RECT 60.400 210.800 62.600 211.600 ;
        RECT 63.600 210.800 65.800 211.600 ;
        RECT 66.800 210.800 69.200 211.600 ;
        RECT 71.600 210.800 72.400 212.400 ;
        RECT 57.200 202.200 58.000 210.800 ;
        RECT 60.400 202.200 61.200 210.800 ;
        RECT 63.600 202.200 64.400 210.800 ;
        RECT 66.800 202.200 67.600 210.800 ;
        RECT 73.000 209.800 73.600 213.600 ;
        RECT 74.200 213.000 75.600 213.800 ;
        RECT 75.000 211.000 75.600 213.000 ;
        RECT 76.400 211.600 77.200 213.200 ;
        RECT 78.000 211.600 78.800 213.200 ;
        RECT 79.600 211.400 80.400 214.800 ;
        RECT 86.600 214.200 87.400 214.400 ;
        RECT 92.400 214.200 93.000 215.600 ;
        RECT 97.200 215.000 98.000 219.800 ;
        RECT 98.800 216.000 99.600 219.800 ;
        RECT 102.000 216.000 102.800 219.800 ;
        RECT 98.800 215.800 102.800 216.000 ;
        RECT 103.600 215.800 104.400 219.800 ;
        RECT 105.200 215.800 106.000 219.800 ;
        RECT 106.800 216.000 107.600 219.800 ;
        RECT 110.000 216.000 110.800 219.800 ;
        RECT 106.800 215.800 110.800 216.000 ;
        RECT 111.600 216.000 112.400 219.800 ;
        RECT 114.800 216.000 115.600 219.800 ;
        RECT 111.600 215.800 115.600 216.000 ;
        RECT 116.400 215.800 117.200 219.800 ;
        RECT 118.000 215.800 118.800 219.800 ;
        RECT 119.600 216.000 120.400 219.800 ;
        RECT 122.800 216.000 123.600 219.800 ;
        RECT 119.600 215.800 123.600 216.000 ;
        RECT 124.400 216.000 125.200 219.800 ;
        RECT 127.600 216.000 128.400 219.800 ;
        RECT 124.400 215.800 128.400 216.000 ;
        RECT 129.200 215.800 130.000 219.800 ;
        RECT 130.800 215.800 131.600 219.800 ;
        RECT 132.400 216.000 133.200 219.800 ;
        RECT 135.600 216.000 136.400 219.800 ;
        RECT 132.400 215.800 136.400 216.000 ;
        RECT 99.000 215.400 102.600 215.800 ;
        RECT 99.600 214.400 100.400 214.800 ;
        RECT 103.600 214.400 104.200 215.800 ;
        RECT 105.400 214.400 106.000 215.800 ;
        RECT 107.000 215.400 110.600 215.800 ;
        RECT 111.800 215.400 115.400 215.800 ;
        RECT 109.200 214.400 110.000 214.800 ;
        RECT 112.400 214.400 113.200 214.800 ;
        RECT 116.400 214.400 117.000 215.800 ;
        RECT 118.200 214.400 118.800 215.800 ;
        RECT 119.800 215.400 123.400 215.800 ;
        RECT 124.600 215.400 128.200 215.800 ;
        RECT 122.000 214.400 122.800 214.800 ;
        RECT 125.200 214.400 126.000 214.800 ;
        RECT 129.200 214.400 129.800 215.800 ;
        RECT 131.000 214.400 131.600 215.800 ;
        RECT 132.600 215.400 136.200 215.800 ;
        RECT 137.200 215.400 138.000 219.800 ;
        RECT 141.400 218.400 142.600 219.800 ;
        RECT 141.400 217.800 142.800 218.400 ;
        RECT 146.000 217.800 146.800 219.800 ;
        RECT 150.400 218.400 151.200 219.800 ;
        RECT 150.400 217.800 152.400 218.400 ;
        RECT 142.000 217.000 142.800 217.800 ;
        RECT 146.200 217.200 146.800 217.800 ;
        RECT 146.200 216.600 149.000 217.200 ;
        RECT 148.200 216.400 149.000 216.600 ;
        RECT 150.000 215.600 150.800 217.200 ;
        RECT 151.600 217.000 152.400 217.800 ;
        RECT 140.200 215.400 141.000 215.600 ;
        RECT 137.200 214.800 141.000 215.400 ;
        RECT 134.800 214.400 135.600 214.800 ;
        RECT 95.600 214.200 97.200 214.400 ;
        RECT 86.200 213.600 97.200 214.200 ;
        RECT 98.800 213.800 100.400 214.400 ;
        RECT 98.800 213.600 99.600 213.800 ;
        RECT 101.800 213.600 104.400 214.400 ;
        RECT 105.200 213.600 107.800 214.400 ;
        RECT 109.200 213.800 110.800 214.400 ;
        RECT 110.000 213.600 110.800 213.800 ;
        RECT 111.600 213.800 113.200 214.400 ;
        RECT 111.600 213.600 112.400 213.800 ;
        RECT 114.600 213.600 117.200 214.400 ;
        RECT 118.000 213.600 120.600 214.400 ;
        RECT 122.000 214.300 123.600 214.400 ;
        RECT 124.400 214.300 126.000 214.400 ;
        RECT 122.000 213.800 126.000 214.300 ;
        RECT 122.800 213.700 125.200 213.800 ;
        RECT 122.800 213.600 123.600 213.700 ;
        RECT 124.400 213.600 125.200 213.700 ;
        RECT 127.400 213.600 130.000 214.400 ;
        RECT 130.800 213.600 133.400 214.400 ;
        RECT 134.800 213.800 136.400 214.400 ;
        RECT 135.600 213.600 136.400 213.800 ;
        RECT 84.400 212.800 85.200 213.000 ;
        RECT 81.400 212.200 85.200 212.800 ;
        RECT 81.400 212.000 82.200 212.200 ;
        RECT 83.000 211.400 83.800 211.600 ;
        RECT 75.000 210.400 78.800 211.000 ;
        RECT 73.000 209.200 74.600 209.800 ;
        RECT 73.800 202.200 74.600 209.200 ;
        RECT 78.200 207.000 78.800 210.400 ;
        RECT 78.000 203.000 78.800 207.000 ;
        RECT 79.600 210.800 83.800 211.400 ;
        RECT 79.600 202.200 80.400 210.800 ;
        RECT 86.200 210.400 86.800 213.600 ;
        RECT 93.400 213.400 94.200 213.600 ;
        RECT 92.400 212.400 93.200 212.600 ;
        RECT 95.000 212.400 95.800 212.600 ;
        RECT 90.800 211.800 95.800 212.400 ;
        RECT 90.800 211.600 91.600 211.800 ;
        RECT 100.400 211.600 101.200 213.200 ;
        RECT 92.400 211.000 98.000 211.200 ;
        RECT 92.200 210.800 98.000 211.000 ;
        RECT 84.400 209.800 86.800 210.400 ;
        RECT 88.200 210.600 98.000 210.800 ;
        RECT 88.200 210.200 93.000 210.600 ;
        RECT 84.400 208.800 85.000 209.800 ;
        RECT 83.600 208.000 85.000 208.800 ;
        RECT 86.600 209.000 87.400 209.200 ;
        RECT 88.200 209.000 88.800 210.200 ;
        RECT 86.600 208.400 88.800 209.000 ;
        RECT 89.400 209.000 94.800 209.600 ;
        RECT 89.400 208.800 90.200 209.000 ;
        RECT 94.000 208.800 94.800 209.000 ;
        RECT 87.800 207.400 88.600 207.600 ;
        RECT 90.600 207.400 91.400 207.600 ;
        RECT 84.400 206.200 85.200 207.000 ;
        RECT 87.800 206.800 91.400 207.400 ;
        RECT 88.600 206.200 89.200 206.800 ;
        RECT 94.000 206.200 94.800 207.000 ;
        RECT 83.800 202.200 85.000 206.200 ;
        RECT 88.400 202.200 89.200 206.200 ;
        RECT 92.800 205.600 94.800 206.200 ;
        RECT 92.800 202.200 93.600 205.600 ;
        RECT 97.200 202.200 98.000 210.600 ;
        RECT 101.800 210.200 102.400 213.600 ;
        RECT 107.200 212.300 107.800 213.600 ;
        RECT 103.700 211.700 107.800 212.300 ;
        RECT 103.700 210.400 104.300 211.700 ;
        RECT 103.600 210.200 104.400 210.400 ;
        RECT 101.400 209.600 102.400 210.200 ;
        RECT 103.000 209.600 104.400 210.200 ;
        RECT 105.200 210.200 106.000 210.400 ;
        RECT 107.200 210.200 107.800 211.700 ;
        RECT 108.400 211.600 109.200 213.200 ;
        RECT 113.200 211.600 114.000 213.200 ;
        RECT 114.600 210.200 115.200 213.600 ;
        RECT 120.000 212.300 120.600 213.600 ;
        RECT 116.500 211.700 120.600 212.300 ;
        RECT 116.500 210.400 117.100 211.700 ;
        RECT 116.400 210.200 117.200 210.400 ;
        RECT 105.200 209.600 106.600 210.200 ;
        RECT 107.200 209.600 108.200 210.200 ;
        RECT 101.400 202.200 102.200 209.600 ;
        RECT 103.000 208.400 103.600 209.600 ;
        RECT 102.800 207.600 103.600 208.400 ;
        RECT 106.000 208.400 106.600 209.600 ;
        RECT 106.000 207.600 106.800 208.400 ;
        RECT 107.400 202.200 108.200 209.600 ;
        RECT 114.200 209.600 115.200 210.200 ;
        RECT 115.800 209.600 117.200 210.200 ;
        RECT 118.000 210.200 118.800 210.400 ;
        RECT 120.000 210.200 120.600 211.700 ;
        RECT 121.200 212.300 122.000 213.200 ;
        RECT 126.000 212.300 126.800 213.200 ;
        RECT 121.200 211.700 126.800 212.300 ;
        RECT 121.200 211.600 122.000 211.700 ;
        RECT 126.000 211.600 126.800 211.700 ;
        RECT 127.400 212.300 128.000 213.600 ;
        RECT 127.400 211.700 131.500 212.300 ;
        RECT 127.400 210.200 128.000 211.700 ;
        RECT 130.900 210.400 131.500 211.700 ;
        RECT 132.800 210.400 133.400 213.600 ;
        RECT 134.000 211.600 134.800 213.200 ;
        RECT 137.200 211.400 138.000 214.800 ;
        RECT 144.200 214.200 145.000 214.400 ;
        RECT 150.000 214.200 150.600 215.600 ;
        RECT 154.800 215.000 155.600 219.800 ;
        RECT 162.800 217.800 163.600 219.800 ;
        RECT 158.000 216.300 158.800 216.400 ;
        RECT 161.200 216.300 162.000 217.200 ;
        RECT 158.000 215.700 162.000 216.300 ;
        RECT 158.000 215.600 158.800 215.700 ;
        RECT 161.200 215.600 162.000 215.700 ;
        RECT 163.000 214.400 163.600 217.800 ;
        RECT 166.000 215.800 166.800 219.800 ;
        RECT 170.400 218.400 172.000 219.800 ;
        RECT 170.400 217.600 173.200 218.400 ;
        RECT 170.400 216.200 172.000 217.600 ;
        RECT 166.000 215.200 168.400 215.800 ;
        RECT 167.600 215.000 168.400 215.200 ;
        RECT 169.000 214.800 169.800 215.600 ;
        RECT 169.000 214.400 169.600 214.800 ;
        RECT 153.200 214.200 154.800 214.400 ;
        RECT 143.800 213.600 154.800 214.200 ;
        RECT 162.800 214.300 163.600 214.400 ;
        RECT 164.400 214.300 165.200 214.400 ;
        RECT 162.800 213.700 165.200 214.300 ;
        RECT 162.800 213.600 163.600 213.700 ;
        RECT 164.400 213.600 165.200 213.700 ;
        RECT 166.000 213.600 167.600 214.400 ;
        RECT 168.800 213.600 169.600 214.400 ;
        RECT 142.000 212.800 142.800 213.000 ;
        RECT 139.000 212.200 142.800 212.800 ;
        RECT 139.000 212.000 139.800 212.200 ;
        RECT 140.600 211.400 141.400 211.600 ;
        RECT 137.200 210.800 141.400 211.400 ;
        RECT 129.200 210.200 130.000 210.400 ;
        RECT 118.000 209.600 119.400 210.200 ;
        RECT 120.000 209.600 121.000 210.200 ;
        RECT 114.200 202.200 115.000 209.600 ;
        RECT 115.800 208.400 116.400 209.600 ;
        RECT 115.600 207.600 116.400 208.400 ;
        RECT 118.800 208.400 119.400 209.600 ;
        RECT 118.800 207.600 119.600 208.400 ;
        RECT 120.200 202.200 121.000 209.600 ;
        RECT 127.000 209.600 128.000 210.200 ;
        RECT 128.600 209.600 130.000 210.200 ;
        RECT 130.800 210.200 131.600 210.400 ;
        RECT 130.800 209.600 132.200 210.200 ;
        RECT 132.800 209.600 134.800 210.400 ;
        RECT 127.000 202.200 127.800 209.600 ;
        RECT 128.600 208.400 129.200 209.600 ;
        RECT 128.400 207.600 129.200 208.400 ;
        RECT 131.600 208.400 132.200 209.600 ;
        RECT 131.600 207.600 132.400 208.400 ;
        RECT 133.000 202.200 133.800 209.600 ;
        RECT 137.200 202.200 138.000 210.800 ;
        RECT 143.800 210.400 144.400 213.600 ;
        RECT 151.000 213.400 151.800 213.600 ;
        RECT 152.600 212.400 153.400 212.600 ;
        RECT 148.400 211.800 153.400 212.400 ;
        RECT 148.400 211.600 149.200 211.800 ;
        RECT 150.000 211.000 155.600 211.200 ;
        RECT 149.800 210.800 155.600 211.000 ;
        RECT 142.000 209.800 144.400 210.400 ;
        RECT 145.800 210.600 155.600 210.800 ;
        RECT 145.800 210.200 150.600 210.600 ;
        RECT 142.000 208.800 142.600 209.800 ;
        RECT 141.200 208.000 142.600 208.800 ;
        RECT 144.200 209.000 145.000 209.200 ;
        RECT 145.800 209.000 146.400 210.200 ;
        RECT 144.200 208.400 146.400 209.000 ;
        RECT 147.000 209.000 152.400 209.600 ;
        RECT 147.000 208.800 147.800 209.000 ;
        RECT 151.600 208.800 152.400 209.000 ;
        RECT 145.400 207.400 146.200 207.600 ;
        RECT 148.200 207.400 149.000 207.600 ;
        RECT 142.000 206.200 142.800 207.000 ;
        RECT 145.400 206.800 149.000 207.400 ;
        RECT 146.200 206.200 146.800 206.800 ;
        RECT 151.600 206.200 152.400 207.000 ;
        RECT 141.400 202.200 142.600 206.200 ;
        RECT 146.000 202.200 146.800 206.200 ;
        RECT 150.400 205.600 152.400 206.200 ;
        RECT 150.400 202.200 151.200 205.600 ;
        RECT 154.800 202.200 155.600 210.600 ;
        RECT 163.000 210.200 163.600 213.600 ;
        RECT 170.400 212.800 171.000 216.200 ;
        RECT 175.600 215.800 176.400 219.800 ;
        RECT 178.800 216.000 179.600 219.800 ;
        RECT 171.600 215.400 173.200 215.600 ;
        RECT 171.600 214.800 173.600 215.400 ;
        RECT 174.200 215.200 176.400 215.800 ;
        RECT 178.600 215.200 179.600 216.000 ;
        RECT 174.200 215.000 175.000 215.200 ;
        RECT 173.000 214.400 173.600 214.800 ;
        RECT 171.600 213.400 172.400 214.200 ;
        RECT 173.000 213.800 176.400 214.400 ;
        RECT 174.800 213.600 176.400 213.800 ;
        RECT 170.000 212.400 171.000 212.800 ;
        RECT 164.400 210.800 165.200 212.400 ;
        RECT 169.200 212.200 171.000 212.400 ;
        RECT 171.800 212.800 172.400 213.400 ;
        RECT 171.800 212.200 174.400 212.800 ;
        RECT 169.200 211.600 170.600 212.200 ;
        RECT 173.600 212.000 174.400 212.200 ;
        RECT 170.000 210.200 170.600 211.600 ;
        RECT 171.400 211.400 172.200 211.600 ;
        RECT 171.400 210.800 174.800 211.400 ;
        RECT 174.200 210.200 174.800 210.800 ;
        RECT 178.600 210.800 179.400 215.200 ;
        RECT 180.400 214.600 181.200 219.800 ;
        RECT 186.800 216.600 187.600 219.800 ;
        RECT 188.400 217.000 189.200 219.800 ;
        RECT 190.000 217.000 190.800 219.800 ;
        RECT 191.600 217.000 192.400 219.800 ;
        RECT 193.200 217.000 194.000 219.800 ;
        RECT 196.400 217.000 197.200 219.800 ;
        RECT 199.600 217.000 200.400 219.800 ;
        RECT 201.200 217.000 202.000 219.800 ;
        RECT 202.800 217.000 203.600 219.800 ;
        RECT 185.200 215.800 187.600 216.600 ;
        RECT 204.400 216.600 205.200 219.800 ;
        RECT 185.200 215.200 186.000 215.800 ;
        RECT 180.000 214.000 181.200 214.600 ;
        RECT 184.200 214.600 186.000 215.200 ;
        RECT 190.000 215.600 191.000 216.400 ;
        RECT 194.000 215.600 195.600 216.400 ;
        RECT 196.400 215.800 201.000 216.400 ;
        RECT 204.400 215.800 207.000 216.600 ;
        RECT 196.400 215.600 197.200 215.800 ;
        RECT 180.000 212.000 180.600 214.000 ;
        RECT 184.200 213.400 185.000 214.600 ;
        RECT 181.200 212.600 185.000 213.400 ;
        RECT 190.000 212.800 190.800 215.600 ;
        RECT 196.400 214.800 197.200 215.000 ;
        RECT 192.800 214.200 197.200 214.800 ;
        RECT 192.800 214.000 193.600 214.200 ;
        RECT 198.000 213.600 198.800 215.200 ;
        RECT 200.200 213.400 201.000 215.800 ;
        RECT 206.200 215.200 207.000 215.800 ;
        RECT 206.200 214.400 209.200 215.200 ;
        RECT 210.800 213.800 211.600 219.800 ;
        RECT 193.200 212.600 196.400 213.400 ;
        RECT 200.200 212.600 202.200 213.400 ;
        RECT 202.800 213.000 211.600 213.800 ;
        RECT 186.800 212.000 187.600 212.600 ;
        RECT 204.400 212.000 205.200 212.400 ;
        RECT 209.400 212.000 210.200 212.200 ;
        RECT 180.000 211.400 180.800 212.000 ;
        RECT 186.800 211.400 210.200 212.000 ;
        RECT 162.800 209.400 164.600 210.200 ;
        RECT 163.800 202.200 164.600 209.400 ;
        RECT 166.000 209.600 168.400 210.200 ;
        RECT 170.000 209.600 172.000 210.200 ;
        RECT 166.000 202.200 166.800 209.600 ;
        RECT 167.600 209.400 168.400 209.600 ;
        RECT 170.400 202.200 172.000 209.600 ;
        RECT 174.200 209.600 176.400 210.200 ;
        RECT 178.600 210.000 179.600 210.800 ;
        RECT 174.200 209.400 175.000 209.600 ;
        RECT 175.600 202.200 176.400 209.600 ;
        RECT 178.800 202.200 179.600 210.000 ;
        RECT 180.200 209.600 180.800 211.400 ;
        RECT 180.200 209.000 189.200 209.600 ;
        RECT 180.200 207.400 180.800 209.000 ;
        RECT 188.400 208.800 189.200 209.000 ;
        RECT 191.600 209.000 200.200 209.600 ;
        RECT 191.600 208.800 192.400 209.000 ;
        RECT 183.400 207.600 186.000 208.400 ;
        RECT 180.200 206.800 182.800 207.400 ;
        RECT 182.000 202.200 182.800 206.800 ;
        RECT 185.200 202.200 186.000 207.600 ;
        RECT 186.600 206.800 190.800 207.600 ;
        RECT 188.400 202.200 189.200 205.000 ;
        RECT 190.000 202.200 190.800 205.000 ;
        RECT 191.600 202.200 192.400 205.000 ;
        RECT 193.200 202.200 194.000 208.400 ;
        RECT 196.400 207.600 199.000 208.400 ;
        RECT 199.600 208.200 200.200 209.000 ;
        RECT 201.200 209.400 202.000 209.600 ;
        RECT 201.200 209.000 206.600 209.400 ;
        RECT 201.200 208.800 207.400 209.000 ;
        RECT 206.000 208.200 207.400 208.800 ;
        RECT 199.600 207.600 205.400 208.200 ;
        RECT 208.400 208.000 210.000 208.800 ;
        RECT 208.400 207.600 209.000 208.000 ;
        RECT 196.400 202.200 197.200 207.000 ;
        RECT 199.600 202.200 200.400 207.000 ;
        RECT 204.800 206.800 209.000 207.600 ;
        RECT 210.800 207.400 211.600 213.000 ;
        RECT 209.600 206.800 211.600 207.400 ;
        RECT 212.400 213.800 213.200 219.800 ;
        RECT 218.800 216.600 219.600 219.800 ;
        RECT 220.400 217.000 221.200 219.800 ;
        RECT 222.000 217.000 222.800 219.800 ;
        RECT 223.600 217.000 224.400 219.800 ;
        RECT 226.800 217.000 227.600 219.800 ;
        RECT 230.000 217.000 230.800 219.800 ;
        RECT 231.600 217.000 232.400 219.800 ;
        RECT 233.200 217.000 234.000 219.800 ;
        RECT 234.800 217.000 235.600 219.800 ;
        RECT 217.000 215.800 219.600 216.600 ;
        RECT 236.400 216.600 237.200 219.800 ;
        RECT 223.000 215.800 227.600 216.400 ;
        RECT 217.000 215.200 217.800 215.800 ;
        RECT 214.800 214.400 217.800 215.200 ;
        RECT 212.400 213.000 221.200 213.800 ;
        RECT 223.000 213.400 223.800 215.800 ;
        RECT 226.800 215.600 227.600 215.800 ;
        RECT 228.400 215.600 230.000 216.400 ;
        RECT 233.000 215.600 234.000 216.400 ;
        RECT 236.400 215.800 238.800 216.600 ;
        RECT 225.200 213.600 226.000 215.200 ;
        RECT 226.800 214.800 227.600 215.000 ;
        RECT 226.800 214.200 231.200 214.800 ;
        RECT 230.400 214.000 231.200 214.200 ;
        RECT 212.400 207.400 213.200 213.000 ;
        RECT 221.800 212.600 223.800 213.400 ;
        RECT 227.600 212.600 230.800 213.400 ;
        RECT 233.200 212.800 234.000 215.600 ;
        RECT 238.000 215.200 238.800 215.800 ;
        RECT 238.000 214.600 239.800 215.200 ;
        RECT 239.000 213.400 239.800 214.600 ;
        RECT 242.800 214.600 243.600 219.800 ;
        RECT 244.400 216.000 245.200 219.800 ;
        RECT 246.000 216.300 246.800 216.400 ;
        RECT 247.600 216.300 248.400 217.200 ;
        RECT 244.400 215.200 245.400 216.000 ;
        RECT 246.000 215.700 248.400 216.300 ;
        RECT 246.000 215.600 246.800 215.700 ;
        RECT 247.600 215.600 248.400 215.700 ;
        RECT 242.800 214.000 244.000 214.600 ;
        RECT 239.000 212.600 242.800 213.400 ;
        RECT 213.800 212.000 214.600 212.200 ;
        RECT 215.600 212.000 216.400 212.400 ;
        RECT 218.800 212.000 219.600 212.400 ;
        RECT 236.400 212.000 237.200 212.600 ;
        RECT 243.400 212.000 244.000 214.000 ;
        RECT 213.800 211.400 237.200 212.000 ;
        RECT 243.200 211.400 244.000 212.000 ;
        RECT 243.200 209.600 243.800 211.400 ;
        RECT 244.600 210.800 245.400 215.200 ;
        RECT 222.000 209.400 222.800 209.600 ;
        RECT 217.400 209.000 222.800 209.400 ;
        RECT 216.600 208.800 222.800 209.000 ;
        RECT 223.800 209.000 232.400 209.600 ;
        RECT 214.000 208.000 215.600 208.800 ;
        RECT 216.600 208.200 218.000 208.800 ;
        RECT 223.800 208.200 224.400 209.000 ;
        RECT 231.600 208.800 232.400 209.000 ;
        RECT 234.800 209.000 243.800 209.600 ;
        RECT 234.800 208.800 235.600 209.000 ;
        RECT 215.000 207.600 215.600 208.000 ;
        RECT 218.600 207.600 224.400 208.200 ;
        RECT 225.000 207.600 227.600 208.400 ;
        RECT 212.400 206.800 214.400 207.400 ;
        RECT 215.000 206.800 219.200 207.600 ;
        RECT 201.200 202.200 202.000 205.000 ;
        RECT 202.800 202.200 203.600 205.000 ;
        RECT 206.000 202.200 206.800 206.800 ;
        RECT 209.600 206.200 210.200 206.800 ;
        RECT 209.200 205.600 210.200 206.200 ;
        RECT 213.800 206.200 214.400 206.800 ;
        RECT 213.800 205.600 214.800 206.200 ;
        RECT 209.200 202.200 210.000 205.600 ;
        RECT 214.000 202.200 214.800 205.600 ;
        RECT 217.200 202.200 218.000 206.800 ;
        RECT 220.400 202.200 221.200 205.000 ;
        RECT 222.000 202.200 222.800 205.000 ;
        RECT 223.600 202.200 224.400 207.000 ;
        RECT 226.800 202.200 227.600 207.000 ;
        RECT 230.000 202.200 230.800 208.400 ;
        RECT 238.000 207.600 240.600 208.400 ;
        RECT 233.200 206.800 237.400 207.600 ;
        RECT 231.600 202.200 232.400 205.000 ;
        RECT 233.200 202.200 234.000 205.000 ;
        RECT 234.800 202.200 235.600 205.000 ;
        RECT 238.000 202.200 238.800 207.600 ;
        RECT 243.200 207.400 243.800 209.000 ;
        RECT 241.200 206.800 243.800 207.400 ;
        RECT 244.400 210.000 245.400 210.800 ;
        RECT 241.200 202.200 242.000 206.800 ;
        RECT 244.400 202.200 245.200 210.000 ;
        RECT 249.200 202.200 250.000 219.800 ;
        RECT 250.800 213.800 251.600 219.800 ;
        RECT 257.200 216.600 258.000 219.800 ;
        RECT 258.800 217.000 259.600 219.800 ;
        RECT 260.400 217.000 261.200 219.800 ;
        RECT 262.000 217.000 262.800 219.800 ;
        RECT 265.200 217.000 266.000 219.800 ;
        RECT 268.400 217.000 269.200 219.800 ;
        RECT 270.000 217.000 270.800 219.800 ;
        RECT 271.600 217.000 272.400 219.800 ;
        RECT 273.200 217.000 274.000 219.800 ;
        RECT 255.400 215.800 258.000 216.600 ;
        RECT 274.800 216.600 275.600 219.800 ;
        RECT 261.400 215.800 266.000 216.400 ;
        RECT 255.400 215.200 256.200 215.800 ;
        RECT 253.200 214.400 256.200 215.200 ;
        RECT 250.800 213.000 259.600 213.800 ;
        RECT 261.400 213.400 262.200 215.800 ;
        RECT 265.200 215.600 266.000 215.800 ;
        RECT 266.800 215.600 268.400 216.400 ;
        RECT 271.400 215.600 272.400 216.400 ;
        RECT 274.800 215.800 277.200 216.600 ;
        RECT 263.600 213.600 264.400 215.200 ;
        RECT 265.200 214.800 266.000 215.000 ;
        RECT 265.200 214.200 269.600 214.800 ;
        RECT 268.800 214.000 269.600 214.200 ;
        RECT 250.800 207.400 251.600 213.000 ;
        RECT 260.200 212.600 262.200 213.400 ;
        RECT 266.000 212.600 269.200 213.400 ;
        RECT 271.600 212.800 272.400 215.600 ;
        RECT 276.400 215.200 277.200 215.800 ;
        RECT 276.400 214.600 278.200 215.200 ;
        RECT 277.400 213.400 278.200 214.600 ;
        RECT 281.200 214.600 282.000 219.800 ;
        RECT 282.800 216.000 283.600 219.800 ;
        RECT 284.400 216.300 285.200 216.400 ;
        RECT 286.000 216.300 286.800 219.800 ;
        RECT 282.800 215.200 283.800 216.000 ;
        RECT 284.400 215.700 286.800 216.300 ;
        RECT 284.400 215.600 285.200 215.700 ;
        RECT 281.200 214.000 282.400 214.600 ;
        RECT 277.400 212.600 281.200 213.400 ;
        RECT 252.200 212.000 253.000 212.200 ;
        RECT 255.600 212.000 256.400 212.400 ;
        RECT 257.200 212.000 258.000 212.400 ;
        RECT 274.800 212.000 275.600 212.600 ;
        RECT 281.800 212.000 282.400 214.000 ;
        RECT 252.200 211.400 275.600 212.000 ;
        RECT 281.600 211.400 282.400 212.000 ;
        RECT 281.600 209.600 282.200 211.400 ;
        RECT 283.000 210.800 283.800 215.200 ;
        RECT 260.400 209.400 261.200 209.600 ;
        RECT 255.800 209.000 261.200 209.400 ;
        RECT 255.000 208.800 261.200 209.000 ;
        RECT 262.200 209.000 270.800 209.600 ;
        RECT 252.400 208.000 254.000 208.800 ;
        RECT 255.000 208.200 256.400 208.800 ;
        RECT 262.200 208.200 262.800 209.000 ;
        RECT 270.000 208.800 270.800 209.000 ;
        RECT 273.200 209.000 282.200 209.600 ;
        RECT 273.200 208.800 274.000 209.000 ;
        RECT 253.400 207.600 254.000 208.000 ;
        RECT 257.000 207.600 262.800 208.200 ;
        RECT 263.400 207.600 266.000 208.400 ;
        RECT 250.800 206.800 252.800 207.400 ;
        RECT 253.400 206.800 257.600 207.600 ;
        RECT 252.200 206.200 252.800 206.800 ;
        RECT 252.200 205.600 253.200 206.200 ;
        RECT 252.400 202.200 253.200 205.600 ;
        RECT 255.600 202.200 256.400 206.800 ;
        RECT 258.800 202.200 259.600 205.000 ;
        RECT 260.400 202.200 261.200 205.000 ;
        RECT 262.000 202.200 262.800 207.000 ;
        RECT 265.200 202.200 266.000 207.000 ;
        RECT 268.400 202.200 269.200 208.400 ;
        RECT 276.400 207.600 279.000 208.400 ;
        RECT 271.600 206.800 275.800 207.600 ;
        RECT 270.000 202.200 270.800 205.000 ;
        RECT 271.600 202.200 272.400 205.000 ;
        RECT 273.200 202.200 274.000 205.000 ;
        RECT 276.400 202.200 277.200 207.600 ;
        RECT 281.600 207.400 282.200 209.000 ;
        RECT 279.600 206.800 282.200 207.400 ;
        RECT 282.800 210.000 283.800 210.800 ;
        RECT 279.600 202.200 280.400 206.800 ;
        RECT 282.800 202.200 283.600 210.000 ;
        RECT 286.000 202.200 286.800 215.700 ;
        RECT 287.600 215.600 288.400 217.200 ;
        RECT 290.800 215.200 291.600 219.800 ;
        RECT 294.000 215.200 294.800 219.800 ;
        RECT 297.200 215.200 298.000 219.800 ;
        RECT 300.400 215.200 301.200 219.800 ;
        RECT 310.000 216.000 310.800 219.800 ;
        RECT 289.200 214.400 291.600 215.200 ;
        RECT 292.600 214.400 294.800 215.200 ;
        RECT 295.800 214.400 298.000 215.200 ;
        RECT 299.400 214.400 301.200 215.200 ;
        RECT 309.800 215.200 310.800 216.000 ;
        RECT 289.200 211.600 290.000 214.400 ;
        RECT 292.600 213.800 293.400 214.400 ;
        RECT 295.800 213.800 296.600 214.400 ;
        RECT 299.400 213.800 300.200 214.400 ;
        RECT 302.000 213.800 302.800 214.400 ;
        RECT 290.800 213.000 293.400 213.800 ;
        RECT 294.200 213.000 296.600 213.800 ;
        RECT 297.600 213.000 300.200 213.800 ;
        RECT 301.000 213.000 302.800 213.800 ;
        RECT 292.600 211.600 293.400 213.000 ;
        RECT 295.800 211.600 296.600 213.000 ;
        RECT 299.400 211.600 300.200 213.000 ;
        RECT 289.200 210.800 291.600 211.600 ;
        RECT 292.600 210.800 294.800 211.600 ;
        RECT 295.800 210.800 298.000 211.600 ;
        RECT 299.400 210.800 301.200 211.600 ;
        RECT 290.800 202.200 291.600 210.800 ;
        RECT 294.000 202.200 294.800 210.800 ;
        RECT 297.200 202.200 298.000 210.800 ;
        RECT 300.400 202.200 301.200 210.800 ;
        RECT 309.800 210.800 310.600 215.200 ;
        RECT 311.600 214.600 312.400 219.800 ;
        RECT 318.000 216.600 318.800 219.800 ;
        RECT 319.600 217.000 320.400 219.800 ;
        RECT 321.200 217.000 322.000 219.800 ;
        RECT 322.800 217.000 323.600 219.800 ;
        RECT 324.400 217.000 325.200 219.800 ;
        RECT 327.600 217.000 328.400 219.800 ;
        RECT 330.800 217.000 331.600 219.800 ;
        RECT 332.400 217.000 333.200 219.800 ;
        RECT 334.000 217.000 334.800 219.800 ;
        RECT 316.400 215.800 318.800 216.600 ;
        RECT 335.600 216.600 336.400 219.800 ;
        RECT 316.400 215.200 317.200 215.800 ;
        RECT 311.200 214.000 312.400 214.600 ;
        RECT 315.400 214.600 317.200 215.200 ;
        RECT 321.200 215.600 322.200 216.400 ;
        RECT 325.200 215.600 326.800 216.400 ;
        RECT 327.600 215.800 332.200 216.400 ;
        RECT 335.600 215.800 338.200 216.600 ;
        RECT 327.600 215.600 328.400 215.800 ;
        RECT 311.200 212.000 311.800 214.000 ;
        RECT 315.400 213.400 316.200 214.600 ;
        RECT 312.400 212.600 316.200 213.400 ;
        RECT 321.200 212.800 322.000 215.600 ;
        RECT 327.600 214.800 328.400 215.000 ;
        RECT 324.000 214.200 328.400 214.800 ;
        RECT 324.000 214.000 324.800 214.200 ;
        RECT 329.200 213.600 330.000 215.200 ;
        RECT 331.400 213.400 332.200 215.800 ;
        RECT 337.400 215.200 338.200 215.800 ;
        RECT 337.400 214.400 340.400 215.200 ;
        RECT 342.000 213.800 342.800 219.800 ;
        RECT 343.600 216.000 344.400 219.800 ;
        RECT 346.800 216.000 347.600 219.800 ;
        RECT 343.600 215.800 347.600 216.000 ;
        RECT 348.400 215.800 349.200 219.800 ;
        RECT 351.600 216.000 352.400 219.800 ;
        RECT 343.800 215.400 347.400 215.800 ;
        RECT 344.400 214.400 345.200 214.800 ;
        RECT 348.400 214.400 349.000 215.800 ;
        RECT 351.400 215.200 352.400 216.000 ;
        RECT 324.400 212.600 327.600 213.400 ;
        RECT 331.400 212.600 333.400 213.400 ;
        RECT 334.000 213.000 342.800 213.800 ;
        RECT 343.600 213.800 345.200 214.400 ;
        RECT 346.600 214.300 349.200 214.400 ;
        RECT 350.000 214.300 350.800 214.400 ;
        RECT 343.600 213.600 344.400 213.800 ;
        RECT 346.600 213.700 350.800 214.300 ;
        RECT 346.600 213.600 349.200 213.700 ;
        RECT 350.000 213.600 350.800 213.700 ;
        RECT 318.000 212.000 318.800 212.600 ;
        RECT 335.600 212.000 336.400 212.400 ;
        RECT 340.400 212.200 341.200 212.400 ;
        RECT 340.400 212.000 341.400 212.200 ;
        RECT 311.200 211.400 312.000 212.000 ;
        RECT 318.000 211.400 341.400 212.000 ;
        RECT 309.800 210.000 310.800 210.800 ;
        RECT 310.000 202.200 310.800 210.000 ;
        RECT 311.400 209.600 312.000 211.400 ;
        RECT 311.400 209.000 320.400 209.600 ;
        RECT 311.400 207.400 312.000 209.000 ;
        RECT 319.600 208.800 320.400 209.000 ;
        RECT 322.800 209.000 331.400 209.600 ;
        RECT 322.800 208.800 323.600 209.000 ;
        RECT 314.600 207.600 317.200 208.400 ;
        RECT 311.400 206.800 314.000 207.400 ;
        RECT 313.200 202.200 314.000 206.800 ;
        RECT 316.400 202.200 317.200 207.600 ;
        RECT 317.800 206.800 322.000 207.600 ;
        RECT 319.600 202.200 320.400 205.000 ;
        RECT 321.200 202.200 322.000 205.000 ;
        RECT 322.800 202.200 323.600 205.000 ;
        RECT 324.400 202.200 325.200 208.400 ;
        RECT 327.600 207.600 330.200 208.400 ;
        RECT 330.800 208.200 331.400 209.000 ;
        RECT 332.400 209.400 333.200 209.600 ;
        RECT 332.400 209.000 337.800 209.400 ;
        RECT 332.400 208.800 338.600 209.000 ;
        RECT 337.200 208.200 338.600 208.800 ;
        RECT 330.800 207.600 336.600 208.200 ;
        RECT 339.600 208.000 341.200 208.800 ;
        RECT 339.600 207.600 340.200 208.000 ;
        RECT 327.600 202.200 328.400 207.000 ;
        RECT 330.800 202.200 331.600 207.000 ;
        RECT 336.000 206.800 340.200 207.600 ;
        RECT 342.000 207.400 342.800 213.000 ;
        RECT 345.200 211.600 346.000 213.200 ;
        RECT 346.600 210.200 347.200 213.600 ;
        RECT 351.400 210.800 352.200 215.200 ;
        RECT 353.200 214.600 354.000 219.800 ;
        RECT 359.600 216.600 360.400 219.800 ;
        RECT 361.200 217.000 362.000 219.800 ;
        RECT 362.800 217.000 363.600 219.800 ;
        RECT 364.400 217.000 365.200 219.800 ;
        RECT 366.000 217.000 366.800 219.800 ;
        RECT 369.200 217.000 370.000 219.800 ;
        RECT 372.400 217.000 373.200 219.800 ;
        RECT 374.000 217.000 374.800 219.800 ;
        RECT 375.600 217.000 376.400 219.800 ;
        RECT 358.000 215.800 360.400 216.600 ;
        RECT 377.200 216.600 378.000 219.800 ;
        RECT 358.000 215.200 358.800 215.800 ;
        RECT 352.800 214.000 354.000 214.600 ;
        RECT 357.000 214.600 358.800 215.200 ;
        RECT 362.800 215.600 363.800 216.400 ;
        RECT 366.800 215.600 368.400 216.400 ;
        RECT 369.200 215.800 373.800 216.400 ;
        RECT 377.200 215.800 379.800 216.600 ;
        RECT 369.200 215.600 370.000 215.800 ;
        RECT 352.800 212.000 353.400 214.000 ;
        RECT 357.000 213.400 357.800 214.600 ;
        RECT 354.000 212.600 357.800 213.400 ;
        RECT 362.800 212.800 363.600 215.600 ;
        RECT 369.200 214.800 370.000 215.000 ;
        RECT 365.600 214.200 370.000 214.800 ;
        RECT 365.600 214.000 366.400 214.200 ;
        RECT 370.800 213.600 371.600 215.200 ;
        RECT 373.000 213.400 373.800 215.800 ;
        RECT 379.000 215.200 379.800 215.800 ;
        RECT 379.000 214.400 382.000 215.200 ;
        RECT 383.600 213.800 384.400 219.800 ;
        RECT 387.800 216.400 388.600 219.800 ;
        RECT 386.800 215.800 388.600 216.400 ;
        RECT 366.000 212.600 369.200 213.400 ;
        RECT 373.000 212.600 375.000 213.400 ;
        RECT 375.600 213.000 384.400 213.800 ;
        RECT 385.200 213.600 386.000 215.200 ;
        RECT 359.600 212.000 360.400 212.600 ;
        RECT 377.200 212.000 378.000 212.400 ;
        RECT 378.800 212.000 379.600 212.400 ;
        RECT 382.200 212.000 383.000 212.200 ;
        RECT 352.800 211.400 353.600 212.000 ;
        RECT 359.600 211.400 383.000 212.000 ;
        RECT 348.400 210.300 349.200 210.400 ;
        RECT 351.400 210.300 352.400 210.800 ;
        RECT 348.400 210.200 352.400 210.300 ;
        RECT 340.800 206.800 342.800 207.400 ;
        RECT 346.200 209.600 347.200 210.200 ;
        RECT 347.800 209.700 352.400 210.200 ;
        RECT 347.800 209.600 349.200 209.700 ;
        RECT 332.400 202.200 333.200 205.000 ;
        RECT 334.000 202.200 334.800 205.000 ;
        RECT 337.200 202.200 338.000 206.800 ;
        RECT 340.800 206.200 341.400 206.800 ;
        RECT 340.400 205.600 341.400 206.200 ;
        RECT 340.400 202.200 341.200 205.600 ;
        RECT 346.200 202.200 347.000 209.600 ;
        RECT 347.800 208.400 348.400 209.600 ;
        RECT 347.600 207.600 348.400 208.400 ;
        RECT 351.600 202.200 352.400 209.700 ;
        RECT 353.000 209.600 353.600 211.400 ;
        RECT 353.000 209.000 362.000 209.600 ;
        RECT 353.000 207.400 353.600 209.000 ;
        RECT 361.200 208.800 362.000 209.000 ;
        RECT 364.400 209.000 373.000 209.600 ;
        RECT 364.400 208.800 365.200 209.000 ;
        RECT 356.200 207.600 358.800 208.400 ;
        RECT 353.000 206.800 355.600 207.400 ;
        RECT 354.800 202.200 355.600 206.800 ;
        RECT 358.000 202.200 358.800 207.600 ;
        RECT 359.400 206.800 363.600 207.600 ;
        RECT 361.200 202.200 362.000 205.000 ;
        RECT 362.800 202.200 363.600 205.000 ;
        RECT 364.400 202.200 365.200 205.000 ;
        RECT 366.000 202.200 366.800 208.400 ;
        RECT 369.200 207.600 371.800 208.400 ;
        RECT 372.400 208.200 373.000 209.000 ;
        RECT 374.000 209.400 374.800 209.600 ;
        RECT 374.000 209.000 379.400 209.400 ;
        RECT 374.000 208.800 380.200 209.000 ;
        RECT 378.800 208.200 380.200 208.800 ;
        RECT 372.400 207.600 378.200 208.200 ;
        RECT 381.200 208.000 382.800 208.800 ;
        RECT 381.200 207.600 381.800 208.000 ;
        RECT 369.200 202.200 370.000 207.000 ;
        RECT 372.400 202.200 373.200 207.000 ;
        RECT 377.600 206.800 381.800 207.600 ;
        RECT 383.600 207.400 384.400 213.000 ;
        RECT 382.400 206.800 384.400 207.400 ;
        RECT 374.000 202.200 374.800 205.000 ;
        RECT 375.600 202.200 376.400 205.000 ;
        RECT 378.800 202.200 379.600 206.800 ;
        RECT 382.400 206.200 383.000 206.800 ;
        RECT 382.000 205.600 383.000 206.200 ;
        RECT 382.000 202.200 382.800 205.600 ;
        RECT 386.800 202.200 387.600 215.800 ;
        RECT 391.600 215.200 392.400 219.800 ;
        RECT 394.800 215.200 395.600 219.800 ;
        RECT 391.600 214.400 395.600 215.200 ;
        RECT 398.000 215.200 398.800 219.800 ;
        RECT 401.200 216.400 402.000 219.800 ;
        RECT 401.200 215.800 402.200 216.400 ;
        RECT 404.400 216.000 405.200 219.800 ;
        RECT 407.600 216.000 408.400 219.800 ;
        RECT 404.400 215.800 408.400 216.000 ;
        RECT 409.200 215.800 410.000 219.800 ;
        RECT 398.000 214.600 400.600 215.200 ;
        RECT 394.800 211.600 395.600 214.400 ;
        RECT 398.200 212.400 399.000 213.200 ;
        RECT 398.000 211.600 399.000 212.400 ;
        RECT 400.000 213.000 400.600 214.600 ;
        RECT 401.600 214.400 402.200 215.800 ;
        RECT 404.600 215.400 408.200 215.800 ;
        RECT 405.200 214.400 406.000 214.800 ;
        RECT 409.200 214.400 409.800 215.800 ;
        RECT 410.800 215.600 411.600 217.200 ;
        RECT 401.200 214.300 402.200 214.400 ;
        RECT 404.400 214.300 406.000 214.400 ;
        RECT 401.200 213.800 406.000 214.300 ;
        RECT 407.400 214.300 410.000 214.400 ;
        RECT 410.800 214.300 411.600 214.400 ;
        RECT 401.200 213.700 405.200 213.800 ;
        RECT 401.200 213.600 402.200 213.700 ;
        RECT 404.400 213.600 405.200 213.700 ;
        RECT 407.400 213.700 411.600 214.300 ;
        RECT 407.400 213.600 410.000 213.700 ;
        RECT 410.800 213.600 411.600 213.700 ;
        RECT 400.000 212.200 401.000 213.000 ;
        RECT 391.600 210.800 395.600 211.600 ;
        RECT 388.400 208.800 389.200 210.400 ;
        RECT 391.600 202.200 392.400 210.800 ;
        RECT 394.800 202.200 395.600 210.800 ;
        RECT 400.000 210.200 400.600 212.200 ;
        RECT 401.600 210.200 402.200 213.600 ;
        RECT 402.800 212.300 403.600 212.400 ;
        RECT 406.000 212.300 406.800 213.200 ;
        RECT 402.800 211.700 406.800 212.300 ;
        RECT 402.800 211.600 403.600 211.700 ;
        RECT 406.000 211.600 406.800 211.700 ;
        RECT 407.400 210.200 408.000 213.600 ;
        RECT 409.200 210.300 410.000 210.400 ;
        RECT 410.800 210.300 411.600 210.400 ;
        RECT 409.200 210.200 411.600 210.300 ;
        RECT 398.000 209.600 400.600 210.200 ;
        RECT 398.000 202.200 398.800 209.600 ;
        RECT 401.200 209.200 402.200 210.200 ;
        RECT 407.000 209.600 408.000 210.200 ;
        RECT 408.600 209.700 411.600 210.200 ;
        RECT 408.600 209.600 410.000 209.700 ;
        RECT 410.800 209.600 411.600 209.700 ;
        RECT 401.200 202.200 402.000 209.200 ;
        RECT 407.000 202.200 407.800 209.600 ;
        RECT 408.600 208.400 409.200 209.600 ;
        RECT 408.400 207.600 409.200 208.400 ;
        RECT 412.400 202.200 413.200 219.800 ;
        RECT 414.000 215.200 414.800 219.800 ;
        RECT 417.200 216.400 418.000 219.800 ;
        RECT 423.000 216.400 423.800 219.800 ;
        RECT 417.200 215.800 418.200 216.400 ;
        RECT 414.000 214.600 416.600 215.200 ;
        RECT 416.000 213.000 416.600 214.600 ;
        RECT 417.600 214.400 418.200 215.800 ;
        RECT 422.000 215.800 423.800 216.400 ;
        RECT 426.800 216.000 427.600 219.800 ;
        RECT 417.200 213.600 418.200 214.400 ;
        RECT 420.400 213.600 421.200 215.200 ;
        RECT 422.000 214.300 422.800 215.800 ;
        RECT 426.600 215.200 427.600 216.000 ;
        RECT 425.200 214.300 426.000 214.400 ;
        RECT 422.000 213.700 426.000 214.300 ;
        RECT 416.000 212.200 417.000 213.000 ;
        RECT 416.000 210.200 416.600 212.200 ;
        RECT 417.600 210.200 418.200 213.600 ;
        RECT 414.000 209.600 416.600 210.200 ;
        RECT 414.000 202.200 414.800 209.600 ;
        RECT 417.200 209.200 418.200 210.200 ;
        RECT 417.200 202.200 418.000 209.200 ;
        RECT 422.000 202.200 422.800 213.700 ;
        RECT 425.200 213.600 426.000 213.700 ;
        RECT 426.600 210.800 427.400 215.200 ;
        RECT 428.400 214.600 429.200 219.800 ;
        RECT 434.800 216.600 435.600 219.800 ;
        RECT 436.400 217.000 437.200 219.800 ;
        RECT 438.000 217.000 438.800 219.800 ;
        RECT 439.600 217.000 440.400 219.800 ;
        RECT 441.200 217.000 442.000 219.800 ;
        RECT 444.400 217.000 445.200 219.800 ;
        RECT 447.600 217.000 448.400 219.800 ;
        RECT 449.200 217.000 450.000 219.800 ;
        RECT 450.800 217.000 451.600 219.800 ;
        RECT 433.200 215.800 435.600 216.600 ;
        RECT 452.400 216.600 453.200 219.800 ;
        RECT 433.200 215.200 434.000 215.800 ;
        RECT 428.000 214.000 429.200 214.600 ;
        RECT 432.200 214.600 434.000 215.200 ;
        RECT 438.000 215.600 439.000 216.400 ;
        RECT 442.000 215.600 443.600 216.400 ;
        RECT 444.400 215.800 449.000 216.400 ;
        RECT 452.400 215.800 455.000 216.600 ;
        RECT 444.400 215.600 445.200 215.800 ;
        RECT 428.000 212.000 428.600 214.000 ;
        RECT 432.200 213.400 433.000 214.600 ;
        RECT 429.200 212.600 433.000 213.400 ;
        RECT 438.000 212.800 438.800 215.600 ;
        RECT 444.400 214.800 445.200 215.000 ;
        RECT 440.800 214.200 445.200 214.800 ;
        RECT 440.800 214.000 441.600 214.200 ;
        RECT 446.000 213.600 446.800 215.200 ;
        RECT 448.200 213.400 449.000 215.800 ;
        RECT 454.200 215.200 455.000 215.800 ;
        RECT 454.200 214.400 457.200 215.200 ;
        RECT 458.800 213.800 459.600 219.800 ;
        RECT 465.200 215.600 466.000 217.200 ;
        RECT 441.200 212.600 444.400 213.400 ;
        RECT 448.200 212.600 450.200 213.400 ;
        RECT 450.800 213.000 459.600 213.800 ;
        RECT 434.800 212.000 435.600 212.600 ;
        RECT 452.400 212.000 453.200 212.400 ;
        RECT 457.400 212.000 458.200 212.200 ;
        RECT 428.000 211.400 428.800 212.000 ;
        RECT 434.800 211.400 458.200 212.000 ;
        RECT 423.600 208.800 424.400 210.400 ;
        RECT 426.600 210.000 427.600 210.800 ;
        RECT 426.800 202.200 427.600 210.000 ;
        RECT 428.200 209.600 428.800 211.400 ;
        RECT 428.200 209.000 437.200 209.600 ;
        RECT 428.200 207.400 428.800 209.000 ;
        RECT 436.400 208.800 437.200 209.000 ;
        RECT 439.600 209.000 448.200 209.600 ;
        RECT 439.600 208.800 440.400 209.000 ;
        RECT 431.400 207.600 434.000 208.400 ;
        RECT 428.200 206.800 430.800 207.400 ;
        RECT 430.000 202.200 430.800 206.800 ;
        RECT 433.200 202.200 434.000 207.600 ;
        RECT 434.600 206.800 438.800 207.600 ;
        RECT 436.400 202.200 437.200 205.000 ;
        RECT 438.000 202.200 438.800 205.000 ;
        RECT 439.600 202.200 440.400 205.000 ;
        RECT 441.200 202.200 442.000 208.400 ;
        RECT 444.400 207.600 447.000 208.400 ;
        RECT 447.600 208.200 448.200 209.000 ;
        RECT 449.200 209.400 450.000 209.600 ;
        RECT 449.200 209.000 454.600 209.400 ;
        RECT 449.200 208.800 455.400 209.000 ;
        RECT 454.000 208.200 455.400 208.800 ;
        RECT 447.600 207.600 453.400 208.200 ;
        RECT 456.400 208.000 458.000 208.800 ;
        RECT 456.400 207.600 457.000 208.000 ;
        RECT 444.400 202.200 445.200 207.000 ;
        RECT 447.600 202.200 448.400 207.000 ;
        RECT 452.800 206.800 457.000 207.600 ;
        RECT 458.800 207.400 459.600 213.000 ;
        RECT 457.600 206.800 459.600 207.400 ;
        RECT 449.200 202.200 450.000 205.000 ;
        RECT 450.800 202.200 451.600 205.000 ;
        RECT 454.000 202.200 454.800 206.800 ;
        RECT 457.600 206.200 458.200 206.800 ;
        RECT 457.200 205.600 458.200 206.200 ;
        RECT 457.200 202.200 458.000 205.600 ;
        RECT 466.800 202.200 467.600 219.800 ;
        RECT 468.400 215.600 469.200 217.200 ;
        RECT 470.000 202.200 470.800 219.800 ;
        RECT 471.600 215.600 472.400 217.200 ;
        RECT 473.200 202.200 474.000 219.800 ;
        RECT 474.800 215.600 475.600 217.200 ;
        RECT 476.400 202.200 477.200 219.800 ;
        RECT 478.000 215.600 478.800 217.200 ;
        RECT 479.600 202.200 480.400 219.800 ;
        RECT 481.800 218.400 482.600 219.800 ;
        RECT 481.200 217.600 482.600 218.400 ;
        RECT 481.800 216.800 482.600 217.600 ;
        RECT 481.200 215.800 482.600 216.800 ;
        RECT 486.000 215.800 486.800 219.800 ;
        RECT 481.200 212.400 481.800 215.800 ;
        RECT 486.000 215.600 486.600 215.800 ;
        RECT 484.800 215.200 486.600 215.600 ;
        RECT 482.400 215.000 486.600 215.200 ;
        RECT 482.400 214.600 485.400 215.000 ;
        RECT 482.400 214.400 483.200 214.600 ;
        RECT 481.200 211.600 482.000 212.400 ;
        RECT 481.200 210.200 481.800 211.600 ;
        RECT 482.600 211.000 483.200 214.400 ;
        RECT 484.000 213.800 484.800 214.000 ;
        RECT 484.000 213.200 485.000 213.800 ;
        RECT 484.400 212.400 485.000 213.200 ;
        RECT 486.000 212.800 486.800 214.400 ;
        RECT 487.600 213.800 488.400 219.800 ;
        RECT 494.000 216.600 494.800 219.800 ;
        RECT 495.600 217.000 496.400 219.800 ;
        RECT 497.200 217.000 498.000 219.800 ;
        RECT 498.800 217.000 499.600 219.800 ;
        RECT 502.000 217.000 502.800 219.800 ;
        RECT 505.200 217.000 506.000 219.800 ;
        RECT 506.800 217.000 507.600 219.800 ;
        RECT 508.400 217.000 509.200 219.800 ;
        RECT 510.000 217.000 510.800 219.800 ;
        RECT 492.200 215.800 494.800 216.600 ;
        RECT 511.600 216.600 512.400 219.800 ;
        RECT 498.200 215.800 502.800 216.400 ;
        RECT 492.200 215.200 493.000 215.800 ;
        RECT 490.000 214.400 493.000 215.200 ;
        RECT 487.600 213.000 496.400 213.800 ;
        RECT 498.200 213.400 499.000 215.800 ;
        RECT 502.000 215.600 502.800 215.800 ;
        RECT 503.600 215.600 505.200 216.400 ;
        RECT 508.200 215.600 509.200 216.400 ;
        RECT 511.600 215.800 514.000 216.600 ;
        RECT 500.400 213.600 501.200 215.200 ;
        RECT 502.000 214.800 502.800 215.000 ;
        RECT 502.000 214.200 506.400 214.800 ;
        RECT 505.600 214.000 506.400 214.200 ;
        RECT 484.400 211.600 485.200 212.400 ;
        RECT 482.600 210.400 485.000 211.000 ;
        RECT 481.200 202.200 482.000 210.200 ;
        RECT 484.400 206.200 485.000 210.400 ;
        RECT 487.600 207.400 488.400 213.000 ;
        RECT 497.000 212.600 499.000 213.400 ;
        RECT 502.800 212.600 506.000 213.400 ;
        RECT 508.400 212.800 509.200 215.600 ;
        RECT 513.200 215.200 514.000 215.800 ;
        RECT 513.200 214.600 515.000 215.200 ;
        RECT 514.200 213.400 515.000 214.600 ;
        RECT 518.000 214.600 518.800 219.800 ;
        RECT 519.600 216.000 520.400 219.800 ;
        RECT 519.600 215.200 520.600 216.000 ;
        RECT 522.800 215.600 523.600 217.200 ;
        RECT 518.000 214.000 519.200 214.600 ;
        RECT 514.200 212.600 518.000 213.400 ;
        RECT 489.000 212.000 489.800 212.200 ;
        RECT 494.000 212.000 494.800 212.400 ;
        RECT 511.600 212.000 512.400 212.600 ;
        RECT 518.600 212.000 519.200 214.000 ;
        RECT 489.000 211.400 512.400 212.000 ;
        RECT 518.400 211.400 519.200 212.000 ;
        RECT 518.400 209.600 519.000 211.400 ;
        RECT 519.800 210.800 520.600 215.200 ;
        RECT 497.200 209.400 498.000 209.600 ;
        RECT 492.600 209.000 498.000 209.400 ;
        RECT 491.800 208.800 498.000 209.000 ;
        RECT 499.000 209.000 507.600 209.600 ;
        RECT 489.200 208.000 490.800 208.800 ;
        RECT 491.800 208.200 493.200 208.800 ;
        RECT 499.000 208.200 499.600 209.000 ;
        RECT 506.800 208.800 507.600 209.000 ;
        RECT 510.000 209.000 519.000 209.600 ;
        RECT 510.000 208.800 510.800 209.000 ;
        RECT 490.200 207.600 490.800 208.000 ;
        RECT 493.800 207.600 499.600 208.200 ;
        RECT 500.200 207.600 502.800 208.400 ;
        RECT 487.600 206.800 489.600 207.400 ;
        RECT 490.200 206.800 494.400 207.600 ;
        RECT 489.000 206.200 489.600 206.800 ;
        RECT 484.400 202.200 485.200 206.200 ;
        RECT 489.000 205.600 490.000 206.200 ;
        RECT 489.200 202.200 490.000 205.600 ;
        RECT 492.400 202.200 493.200 206.800 ;
        RECT 495.600 202.200 496.400 205.000 ;
        RECT 497.200 202.200 498.000 205.000 ;
        RECT 498.800 202.200 499.600 207.000 ;
        RECT 502.000 202.200 502.800 207.000 ;
        RECT 505.200 202.200 506.000 208.400 ;
        RECT 513.200 207.600 515.800 208.400 ;
        RECT 508.400 206.800 512.600 207.600 ;
        RECT 506.800 202.200 507.600 205.000 ;
        RECT 508.400 202.200 509.200 205.000 ;
        RECT 510.000 202.200 510.800 205.000 ;
        RECT 513.200 202.200 514.000 207.600 ;
        RECT 518.400 207.400 519.000 209.000 ;
        RECT 516.400 206.800 519.000 207.400 ;
        RECT 519.600 210.000 520.600 210.800 ;
        RECT 524.400 212.300 525.200 219.800 ;
        RECT 526.000 216.000 526.800 219.800 ;
        RECT 529.200 216.000 530.000 219.800 ;
        RECT 526.000 215.800 530.000 216.000 ;
        RECT 530.800 215.800 531.600 219.800 ;
        RECT 533.000 218.400 533.800 219.800 ;
        RECT 533.000 217.600 534.800 218.400 ;
        RECT 533.000 216.400 533.800 217.600 ;
        RECT 533.000 215.800 534.800 216.400 ;
        RECT 538.800 216.000 539.600 219.800 ;
        RECT 526.200 215.400 529.800 215.800 ;
        RECT 526.800 214.400 527.600 214.800 ;
        RECT 530.800 214.400 531.400 215.800 ;
        RECT 526.000 213.800 527.600 214.400 ;
        RECT 526.000 213.600 526.800 213.800 ;
        RECT 529.000 213.600 531.600 214.400 ;
        RECT 527.600 212.300 528.400 213.200 ;
        RECT 524.400 211.700 528.400 212.300 ;
        RECT 516.400 202.200 517.200 206.800 ;
        RECT 519.600 202.200 520.400 210.000 ;
        RECT 524.400 202.200 525.200 211.700 ;
        RECT 527.600 211.600 528.400 211.700 ;
        RECT 529.000 212.300 529.600 213.600 ;
        RECT 529.000 211.700 533.100 212.300 ;
        RECT 529.000 210.200 529.600 211.700 ;
        RECT 532.500 210.400 533.100 211.700 ;
        RECT 530.800 210.200 531.600 210.400 ;
        RECT 528.600 209.600 529.600 210.200 ;
        RECT 530.200 209.600 531.600 210.200 ;
        RECT 528.600 202.200 529.400 209.600 ;
        RECT 530.200 208.400 530.800 209.600 ;
        RECT 532.400 208.800 533.200 210.400 ;
        RECT 530.000 207.600 530.800 208.400 ;
        RECT 534.000 202.200 534.800 215.800 ;
        RECT 538.600 215.200 539.600 216.000 ;
        RECT 535.600 213.600 536.400 215.200 ;
        RECT 538.600 210.800 539.400 215.200 ;
        RECT 540.400 214.600 541.200 219.800 ;
        RECT 546.800 216.600 547.600 219.800 ;
        RECT 548.400 217.000 549.200 219.800 ;
        RECT 550.000 217.000 550.800 219.800 ;
        RECT 551.600 217.000 552.400 219.800 ;
        RECT 553.200 217.000 554.000 219.800 ;
        RECT 556.400 217.000 557.200 219.800 ;
        RECT 559.600 217.000 560.400 219.800 ;
        RECT 561.200 217.000 562.000 219.800 ;
        RECT 562.800 217.000 563.600 219.800 ;
        RECT 545.200 215.800 547.600 216.600 ;
        RECT 564.400 216.600 565.200 219.800 ;
        RECT 545.200 215.200 546.000 215.800 ;
        RECT 540.000 214.000 541.200 214.600 ;
        RECT 544.200 214.600 546.000 215.200 ;
        RECT 550.000 215.600 551.000 216.400 ;
        RECT 554.000 215.600 555.600 216.400 ;
        RECT 556.400 215.800 561.000 216.400 ;
        RECT 564.400 215.800 567.000 216.600 ;
        RECT 556.400 215.600 557.200 215.800 ;
        RECT 540.000 212.000 540.600 214.000 ;
        RECT 544.200 213.400 545.000 214.600 ;
        RECT 541.200 212.600 545.000 213.400 ;
        RECT 550.000 212.800 550.800 215.600 ;
        RECT 556.400 214.800 557.200 215.000 ;
        RECT 552.800 214.200 557.200 214.800 ;
        RECT 552.800 214.000 553.600 214.200 ;
        RECT 558.000 213.600 558.800 215.200 ;
        RECT 560.200 213.400 561.000 215.800 ;
        RECT 566.200 215.200 567.000 215.800 ;
        RECT 566.200 214.400 569.200 215.200 ;
        RECT 570.800 213.800 571.600 219.800 ;
        RECT 572.400 216.000 573.200 219.800 ;
        RECT 575.600 216.000 576.400 219.800 ;
        RECT 572.400 215.800 576.400 216.000 ;
        RECT 577.200 215.800 578.000 219.800 ;
        RECT 572.600 215.400 576.200 215.800 ;
        RECT 573.200 214.400 574.000 214.800 ;
        RECT 577.200 214.400 577.800 215.800 ;
        RECT 580.400 215.200 581.200 219.800 ;
        RECT 583.600 215.200 584.400 219.800 ;
        RECT 586.800 215.200 587.600 219.800 ;
        RECT 590.000 215.200 590.800 219.800 ;
        RECT 578.800 214.400 581.200 215.200 ;
        RECT 582.200 214.400 584.400 215.200 ;
        RECT 585.400 214.400 587.600 215.200 ;
        RECT 589.000 214.400 590.800 215.200 ;
        RECT 594.800 215.200 595.600 219.800 ;
        RECT 598.000 215.200 598.800 219.800 ;
        RECT 601.200 215.200 602.000 219.800 ;
        RECT 604.400 215.200 605.200 219.800 ;
        RECT 594.800 214.400 596.600 215.200 ;
        RECT 598.000 214.400 600.200 215.200 ;
        RECT 601.200 214.400 603.400 215.200 ;
        RECT 604.400 214.400 606.800 215.200 ;
        RECT 553.200 212.600 556.400 213.400 ;
        RECT 560.200 212.600 562.200 213.400 ;
        RECT 562.800 213.000 571.600 213.800 ;
        RECT 572.400 213.800 574.000 214.400 ;
        RECT 572.400 213.600 573.200 213.800 ;
        RECT 575.400 213.600 578.000 214.400 ;
        RECT 546.800 212.000 547.600 212.600 ;
        RECT 564.400 212.000 565.200 212.400 ;
        RECT 567.600 212.000 568.400 212.400 ;
        RECT 569.400 212.000 570.200 212.200 ;
        RECT 540.000 211.400 540.800 212.000 ;
        RECT 546.800 211.400 570.200 212.000 ;
        RECT 538.600 210.000 539.600 210.800 ;
        RECT 538.800 202.200 539.600 210.000 ;
        RECT 540.200 209.600 540.800 211.400 ;
        RECT 540.200 209.000 549.200 209.600 ;
        RECT 540.200 207.400 540.800 209.000 ;
        RECT 548.400 208.800 549.200 209.000 ;
        RECT 551.600 209.000 560.200 209.600 ;
        RECT 551.600 208.800 552.400 209.000 ;
        RECT 543.400 207.600 546.000 208.400 ;
        RECT 540.200 206.800 542.800 207.400 ;
        RECT 542.000 202.200 542.800 206.800 ;
        RECT 545.200 202.200 546.000 207.600 ;
        RECT 546.600 206.800 550.800 207.600 ;
        RECT 548.400 202.200 549.200 205.000 ;
        RECT 550.000 202.200 550.800 205.000 ;
        RECT 551.600 202.200 552.400 205.000 ;
        RECT 553.200 202.200 554.000 208.400 ;
        RECT 556.400 207.600 559.000 208.400 ;
        RECT 559.600 208.200 560.200 209.000 ;
        RECT 561.200 209.400 562.000 209.600 ;
        RECT 561.200 209.000 566.600 209.400 ;
        RECT 561.200 208.800 567.400 209.000 ;
        RECT 566.000 208.200 567.400 208.800 ;
        RECT 559.600 207.600 565.400 208.200 ;
        RECT 568.400 208.000 570.000 208.800 ;
        RECT 568.400 207.600 569.000 208.000 ;
        RECT 556.400 202.200 557.200 207.000 ;
        RECT 559.600 202.200 560.400 207.000 ;
        RECT 564.800 206.800 569.000 207.600 ;
        RECT 570.800 207.400 571.600 213.000 ;
        RECT 574.000 211.600 574.800 213.200 ;
        RECT 575.400 212.400 576.000 213.600 ;
        RECT 575.400 211.600 576.400 212.400 ;
        RECT 578.800 211.600 579.600 214.400 ;
        RECT 582.200 213.800 583.000 214.400 ;
        RECT 585.400 213.800 586.200 214.400 ;
        RECT 589.000 213.800 589.800 214.400 ;
        RECT 591.600 214.300 592.400 214.400 ;
        RECT 593.200 214.300 594.000 214.400 ;
        RECT 591.600 213.800 594.000 214.300 ;
        RECT 595.800 213.800 596.600 214.400 ;
        RECT 599.400 213.800 600.200 214.400 ;
        RECT 602.600 213.800 603.400 214.400 ;
        RECT 580.400 213.000 583.000 213.800 ;
        RECT 583.800 213.000 586.200 213.800 ;
        RECT 587.200 213.000 589.800 213.800 ;
        RECT 590.600 213.700 595.000 213.800 ;
        RECT 590.600 213.000 592.400 213.700 ;
        RECT 593.200 213.000 595.000 213.700 ;
        RECT 595.800 213.000 598.400 213.800 ;
        RECT 599.400 213.000 601.800 213.800 ;
        RECT 602.600 213.000 605.200 213.800 ;
        RECT 582.200 211.600 583.000 213.000 ;
        RECT 585.400 211.600 586.200 213.000 ;
        RECT 589.000 211.600 589.800 213.000 ;
        RECT 595.800 211.600 596.600 213.000 ;
        RECT 599.400 211.600 600.200 213.000 ;
        RECT 602.600 211.600 603.400 213.000 ;
        RECT 606.000 211.600 606.800 214.400 ;
        RECT 575.400 210.200 576.000 211.600 ;
        RECT 578.800 210.800 581.200 211.600 ;
        RECT 582.200 210.800 584.400 211.600 ;
        RECT 585.400 210.800 587.600 211.600 ;
        RECT 589.000 210.800 590.800 211.600 ;
        RECT 577.200 210.200 578.000 210.400 ;
        RECT 569.600 206.800 571.600 207.400 ;
        RECT 575.000 209.600 576.000 210.200 ;
        RECT 576.600 209.600 578.000 210.200 ;
        RECT 561.200 202.200 562.000 205.000 ;
        RECT 562.800 202.200 563.600 205.000 ;
        RECT 566.000 202.200 566.800 206.800 ;
        RECT 569.600 206.200 570.200 206.800 ;
        RECT 569.200 205.600 570.200 206.200 ;
        RECT 569.200 202.200 570.000 205.600 ;
        RECT 575.000 202.200 575.800 209.600 ;
        RECT 576.600 208.400 577.200 209.600 ;
        RECT 576.400 207.600 577.200 208.400 ;
        RECT 580.400 202.200 581.200 210.800 ;
        RECT 583.600 202.200 584.400 210.800 ;
        RECT 586.800 202.200 587.600 210.800 ;
        RECT 590.000 202.200 590.800 210.800 ;
        RECT 594.800 210.800 596.600 211.600 ;
        RECT 598.000 210.800 600.200 211.600 ;
        RECT 601.200 210.800 603.400 211.600 ;
        RECT 604.400 210.800 606.800 211.600 ;
        RECT 594.800 202.200 595.600 210.800 ;
        RECT 598.000 202.200 598.800 210.800 ;
        RECT 601.200 202.200 602.000 210.800 ;
        RECT 604.400 202.200 605.200 210.800 ;
        RECT 2.800 196.400 3.600 199.800 ;
        RECT 2.600 195.800 3.600 196.400 ;
        RECT 2.600 195.200 3.200 195.800 ;
        RECT 6.000 195.200 6.800 199.800 ;
        RECT 9.200 197.000 10.000 199.800 ;
        RECT 10.800 197.000 11.600 199.800 ;
        RECT 1.200 194.600 3.200 195.200 ;
        RECT 1.200 189.000 2.000 194.600 ;
        RECT 3.800 194.400 8.000 195.200 ;
        RECT 12.400 195.000 13.200 199.800 ;
        RECT 15.600 195.000 16.400 199.800 ;
        RECT 3.800 194.000 4.400 194.400 ;
        RECT 2.800 193.200 4.400 194.000 ;
        RECT 7.400 193.800 13.200 194.400 ;
        RECT 5.400 193.200 6.800 193.800 ;
        RECT 5.400 193.000 11.600 193.200 ;
        RECT 6.200 192.600 11.600 193.000 ;
        RECT 10.800 192.400 11.600 192.600 ;
        RECT 12.600 193.000 13.200 193.800 ;
        RECT 13.800 193.600 16.400 194.400 ;
        RECT 18.800 193.600 19.600 199.800 ;
        RECT 20.400 197.000 21.200 199.800 ;
        RECT 22.000 197.000 22.800 199.800 ;
        RECT 23.600 197.000 24.400 199.800 ;
        RECT 22.000 194.400 26.200 195.200 ;
        RECT 26.800 194.400 27.600 199.800 ;
        RECT 30.000 195.200 30.800 199.800 ;
        RECT 30.000 194.600 32.600 195.200 ;
        RECT 26.800 193.600 29.400 194.400 ;
        RECT 20.400 193.000 21.200 193.200 ;
        RECT 12.600 192.400 21.200 193.000 ;
        RECT 23.600 193.000 24.400 193.200 ;
        RECT 32.000 193.000 32.600 194.600 ;
        RECT 23.600 192.400 32.600 193.000 ;
        RECT 32.000 190.600 32.600 192.400 ;
        RECT 33.200 192.000 34.000 199.800 ;
        RECT 33.200 191.200 34.200 192.000 ;
        RECT 2.600 190.000 26.000 190.600 ;
        RECT 32.000 190.000 32.800 190.600 ;
        RECT 2.600 189.800 3.400 190.000 ;
        RECT 7.600 189.600 8.400 190.000 ;
        RECT 25.200 189.400 26.000 190.000 ;
        RECT 1.200 188.200 10.000 189.000 ;
        RECT 10.600 188.600 12.600 189.400 ;
        RECT 16.400 188.600 19.600 189.400 ;
        RECT 1.200 182.200 2.000 188.200 ;
        RECT 3.600 186.800 6.600 187.600 ;
        RECT 5.800 186.200 6.600 186.800 ;
        RECT 11.800 186.200 12.600 188.600 ;
        RECT 14.000 186.800 14.800 188.400 ;
        RECT 19.200 187.800 20.000 188.000 ;
        RECT 15.600 187.200 20.000 187.800 ;
        RECT 15.600 187.000 16.400 187.200 ;
        RECT 22.000 186.400 22.800 189.200 ;
        RECT 27.800 188.600 31.600 189.400 ;
        RECT 27.800 187.400 28.600 188.600 ;
        RECT 32.200 188.000 32.800 190.000 ;
        RECT 15.600 186.200 16.400 186.400 ;
        RECT 5.800 185.400 8.400 186.200 ;
        RECT 11.800 185.600 16.400 186.200 ;
        RECT 17.200 185.600 18.800 186.400 ;
        RECT 21.800 185.600 22.800 186.400 ;
        RECT 26.800 186.800 28.600 187.400 ;
        RECT 31.600 187.400 32.800 188.000 ;
        RECT 26.800 186.200 27.600 186.800 ;
        RECT 7.600 182.200 8.400 185.400 ;
        RECT 25.200 185.400 27.600 186.200 ;
        RECT 9.200 182.200 10.000 185.000 ;
        RECT 10.800 182.200 11.600 185.000 ;
        RECT 12.400 182.200 13.200 185.000 ;
        RECT 15.600 182.200 16.400 185.000 ;
        RECT 18.800 182.200 19.600 185.000 ;
        RECT 20.400 182.200 21.200 185.000 ;
        RECT 22.000 182.200 22.800 185.000 ;
        RECT 23.600 182.200 24.400 185.000 ;
        RECT 25.200 182.200 26.000 185.400 ;
        RECT 31.600 182.200 32.400 187.400 ;
        RECT 33.400 186.800 34.200 191.200 ;
        RECT 33.200 186.000 34.200 186.800 ;
        RECT 33.200 182.200 34.000 186.000 ;
        RECT 36.400 182.200 37.200 199.800 ;
        RECT 39.600 191.400 40.400 199.800 ;
        RECT 44.000 196.400 44.800 199.800 ;
        RECT 42.800 195.800 44.800 196.400 ;
        RECT 48.400 195.800 49.200 199.800 ;
        RECT 52.600 195.800 53.800 199.800 ;
        RECT 42.800 195.000 43.600 195.800 ;
        RECT 48.400 195.200 49.000 195.800 ;
        RECT 46.200 194.600 49.800 195.200 ;
        RECT 52.400 195.000 53.200 195.800 ;
        RECT 46.200 194.400 47.000 194.600 ;
        RECT 49.000 194.400 49.800 194.600 ;
        RECT 42.800 193.000 43.600 193.200 ;
        RECT 47.400 193.000 48.200 193.200 ;
        RECT 42.800 192.400 48.200 193.000 ;
        RECT 48.800 193.000 51.000 193.600 ;
        RECT 48.800 191.800 49.400 193.000 ;
        RECT 50.200 192.800 51.000 193.000 ;
        RECT 52.600 193.200 54.000 194.000 ;
        RECT 52.600 192.200 53.200 193.200 ;
        RECT 44.600 191.400 49.400 191.800 ;
        RECT 39.600 191.200 49.400 191.400 ;
        RECT 50.800 191.600 53.200 192.200 ;
        RECT 39.600 191.000 45.400 191.200 ;
        RECT 39.600 190.800 45.200 191.000 ;
        RECT 46.000 190.300 46.800 190.400 ;
        RECT 47.600 190.300 48.400 190.400 ;
        RECT 46.000 190.200 48.400 190.300 ;
        RECT 41.800 189.700 48.400 190.200 ;
        RECT 41.800 189.600 46.800 189.700 ;
        RECT 47.600 189.600 48.400 189.700 ;
        RECT 41.800 189.400 42.600 189.600 ;
        RECT 43.400 188.400 44.200 188.600 ;
        RECT 50.800 188.400 51.400 191.600 ;
        RECT 57.200 191.200 58.000 199.800 ;
        RECT 59.600 193.600 60.400 194.400 ;
        RECT 59.600 192.400 60.200 193.600 ;
        RECT 61.000 192.400 61.800 199.800 ;
        RECT 67.800 192.400 68.600 199.800 ;
        RECT 69.200 193.600 70.000 194.400 ;
        RECT 69.400 192.400 70.000 193.600 ;
        RECT 75.400 192.800 76.200 199.800 ;
        RECT 79.600 195.000 80.400 199.000 ;
        RECT 58.800 191.800 60.200 192.400 ;
        RECT 60.800 191.800 61.800 192.400 ;
        RECT 58.800 191.600 59.600 191.800 ;
        RECT 53.800 190.600 58.000 191.200 ;
        RECT 53.800 190.400 54.600 190.600 ;
        RECT 55.400 189.800 56.200 190.000 ;
        RECT 52.400 189.200 56.200 189.800 ;
        RECT 52.400 189.000 53.200 189.200 ;
        RECT 40.400 187.800 51.400 188.400 ;
        RECT 40.400 187.600 42.000 187.800 ;
        RECT 38.000 184.800 38.800 186.400 ;
        RECT 39.600 182.200 40.400 187.000 ;
        RECT 44.600 185.600 45.200 187.800 ;
        RECT 50.200 187.600 51.000 187.800 ;
        RECT 57.200 187.200 58.000 190.600 ;
        RECT 58.800 190.300 59.600 190.400 ;
        RECT 60.800 190.300 61.400 191.800 ;
        RECT 66.800 191.600 68.800 192.400 ;
        RECT 69.400 191.800 70.800 192.400 ;
        RECT 70.000 191.600 70.800 191.800 ;
        RECT 74.600 192.200 76.200 192.800 ;
        RECT 58.800 189.700 61.400 190.300 ;
        RECT 58.800 189.600 59.600 189.700 ;
        RECT 60.800 188.400 61.400 189.700 ;
        RECT 62.000 188.800 62.800 190.400 ;
        RECT 66.800 188.800 67.600 190.400 ;
        RECT 68.200 188.400 68.800 191.600 ;
        RECT 73.200 189.600 74.000 191.200 ;
        RECT 74.600 188.400 75.200 192.200 ;
        RECT 79.800 191.600 80.400 195.000 ;
        RECT 82.800 192.800 83.600 199.800 ;
        RECT 76.600 191.000 80.400 191.600 ;
        RECT 82.600 191.800 83.600 192.800 ;
        RECT 86.000 192.400 86.800 199.800 ;
        RECT 84.200 191.800 86.800 192.400 ;
        RECT 76.600 189.000 77.200 191.000 ;
        RECT 58.800 187.600 61.400 188.400 ;
        RECT 63.600 188.200 64.400 188.400 ;
        RECT 62.800 187.600 64.400 188.200 ;
        RECT 65.200 188.200 66.000 188.400 ;
        RECT 65.200 187.600 66.800 188.200 ;
        RECT 68.200 187.600 70.800 188.400 ;
        RECT 71.600 188.300 72.400 188.400 ;
        RECT 73.200 188.300 75.200 188.400 ;
        RECT 71.600 187.700 75.200 188.300 ;
        RECT 75.800 188.200 77.200 189.000 ;
        RECT 78.000 188.800 78.800 190.400 ;
        RECT 79.600 188.800 80.400 190.400 ;
        RECT 71.600 187.600 72.400 187.700 ;
        RECT 73.200 187.600 75.200 187.700 ;
        RECT 54.200 186.600 58.000 187.200 ;
        RECT 54.200 186.400 55.000 186.600 ;
        RECT 42.800 184.200 43.600 185.000 ;
        RECT 44.400 184.800 45.200 185.600 ;
        RECT 46.200 185.400 47.000 185.600 ;
        RECT 46.200 184.800 49.000 185.400 ;
        RECT 48.400 184.200 49.000 184.800 ;
        RECT 52.400 184.200 53.200 185.000 ;
        RECT 42.800 183.600 44.800 184.200 ;
        RECT 44.000 182.200 44.800 183.600 ;
        RECT 48.400 182.200 49.200 184.200 ;
        RECT 52.400 183.600 53.800 184.200 ;
        RECT 52.600 182.200 53.800 183.600 ;
        RECT 57.200 182.200 58.000 186.600 ;
        RECT 59.000 186.200 59.600 187.600 ;
        RECT 62.800 187.200 63.600 187.600 ;
        RECT 66.000 187.200 66.800 187.600 ;
        RECT 60.600 186.200 64.200 186.600 ;
        RECT 65.400 186.200 69.000 186.600 ;
        RECT 70.000 186.200 70.600 187.600 ;
        RECT 74.600 187.000 75.200 187.600 ;
        RECT 76.200 187.800 77.200 188.200 ;
        RECT 82.600 188.400 83.200 191.800 ;
        RECT 84.200 189.800 84.800 191.800 ;
        RECT 87.600 191.400 88.400 199.800 ;
        RECT 92.000 196.400 92.800 199.800 ;
        RECT 90.800 195.800 92.800 196.400 ;
        RECT 96.400 195.800 97.200 199.800 ;
        RECT 100.600 195.800 101.800 199.800 ;
        RECT 90.800 195.000 91.600 195.800 ;
        RECT 96.400 195.200 97.000 195.800 ;
        RECT 94.200 194.600 97.800 195.200 ;
        RECT 100.400 195.000 101.200 195.800 ;
        RECT 94.200 194.400 95.000 194.600 ;
        RECT 97.000 194.400 97.800 194.600 ;
        RECT 90.800 193.000 91.600 193.200 ;
        RECT 95.400 193.000 96.200 193.200 ;
        RECT 90.800 192.400 96.200 193.000 ;
        RECT 96.800 193.000 99.000 193.600 ;
        RECT 96.800 191.800 97.400 193.000 ;
        RECT 98.200 192.800 99.000 193.000 ;
        RECT 100.600 193.200 102.000 194.000 ;
        RECT 100.600 192.200 101.200 193.200 ;
        RECT 92.600 191.400 97.400 191.800 ;
        RECT 87.600 191.200 97.400 191.400 ;
        RECT 98.800 191.600 101.200 192.200 ;
        RECT 87.600 191.000 93.400 191.200 ;
        RECT 87.600 190.800 93.200 191.000 ;
        RECT 83.800 189.000 84.800 189.800 ;
        RECT 76.200 187.200 80.400 187.800 ;
        RECT 74.600 186.600 75.400 187.000 ;
        RECT 58.800 182.200 59.600 186.200 ;
        RECT 60.400 186.000 64.400 186.200 ;
        RECT 60.400 182.200 61.200 186.000 ;
        RECT 63.600 182.200 64.400 186.000 ;
        RECT 65.200 186.000 69.200 186.200 ;
        RECT 65.200 182.200 66.000 186.000 ;
        RECT 68.400 182.200 69.200 186.000 ;
        RECT 70.000 182.200 70.800 186.200 ;
        RECT 74.600 186.000 76.200 186.600 ;
        RECT 75.400 183.000 76.200 186.000 ;
        RECT 79.800 185.000 80.400 187.200 ;
        RECT 82.600 187.600 83.600 188.400 ;
        RECT 82.600 186.200 83.200 187.600 ;
        RECT 84.200 187.400 84.800 189.000 ;
        RECT 85.800 189.600 86.800 190.400 ;
        RECT 94.000 190.200 94.800 190.400 ;
        RECT 89.800 189.600 94.800 190.200 ;
        RECT 85.800 188.800 86.600 189.600 ;
        RECT 89.800 189.400 90.600 189.600 ;
        RECT 91.400 188.400 92.200 188.600 ;
        RECT 98.800 188.400 99.400 191.600 ;
        RECT 105.200 191.200 106.000 199.800 ;
        RECT 109.400 192.400 110.200 199.800 ;
        RECT 113.200 195.000 114.000 199.000 ;
        RECT 117.400 198.400 118.200 199.800 ;
        RECT 116.400 197.600 118.200 198.400 ;
        RECT 110.800 193.600 111.600 194.400 ;
        RECT 111.000 192.400 111.600 193.600 ;
        RECT 108.400 191.600 110.400 192.400 ;
        RECT 111.000 191.800 112.400 192.400 ;
        RECT 111.600 191.600 112.400 191.800 ;
        RECT 113.200 191.600 113.800 195.000 ;
        RECT 117.400 192.800 118.200 197.600 ;
        RECT 123.600 193.600 124.400 194.400 ;
        RECT 117.400 192.200 119.000 192.800 ;
        RECT 123.600 192.400 124.200 193.600 ;
        RECT 125.000 192.400 125.800 199.800 ;
        RECT 101.800 190.600 106.000 191.200 ;
        RECT 101.800 190.400 102.600 190.600 ;
        RECT 103.400 189.800 104.200 190.000 ;
        RECT 100.400 189.200 104.200 189.800 ;
        RECT 100.400 189.000 101.200 189.200 ;
        RECT 88.400 187.800 99.400 188.400 ;
        RECT 88.400 187.600 90.000 187.800 ;
        RECT 84.200 186.800 86.800 187.400 ;
        RECT 82.600 185.600 83.600 186.200 ;
        RECT 79.600 183.000 80.400 185.000 ;
        RECT 82.800 182.200 83.600 185.600 ;
        RECT 86.000 182.200 86.800 186.800 ;
        RECT 87.600 182.200 88.400 187.000 ;
        RECT 92.600 185.600 93.200 187.800 ;
        RECT 98.200 187.600 99.000 187.800 ;
        RECT 105.200 187.200 106.000 190.600 ;
        RECT 108.400 188.800 109.200 190.400 ;
        RECT 109.800 188.400 110.400 191.600 ;
        RECT 113.200 191.000 117.000 191.600 ;
        RECT 113.200 188.800 114.000 190.400 ;
        RECT 114.800 188.800 115.600 190.400 ;
        RECT 116.400 189.000 117.000 191.000 ;
        RECT 106.800 188.200 107.600 188.400 ;
        RECT 106.800 187.600 108.400 188.200 ;
        RECT 109.800 187.600 112.400 188.400 ;
        RECT 116.400 188.200 117.800 189.000 ;
        RECT 118.400 188.400 119.000 192.200 ;
        RECT 122.800 191.800 124.200 192.400 ;
        RECT 124.800 191.800 125.800 192.400 ;
        RECT 129.200 195.000 130.000 199.000 ;
        RECT 133.400 198.400 134.200 199.800 ;
        RECT 132.400 197.600 134.200 198.400 ;
        RECT 122.800 191.600 123.600 191.800 ;
        RECT 119.600 189.600 120.400 191.200 ;
        RECT 121.200 190.300 122.000 190.400 ;
        RECT 124.800 190.300 125.400 191.800 ;
        RECT 129.200 191.600 129.800 195.000 ;
        RECT 133.400 192.800 134.200 197.600 ;
        RECT 133.400 192.200 135.000 192.800 ;
        RECT 129.200 191.000 133.000 191.600 ;
        RECT 121.200 189.700 125.400 190.300 ;
        RECT 121.200 189.600 122.000 189.700 ;
        RECT 124.800 188.400 125.400 189.700 ;
        RECT 126.000 188.800 126.800 190.400 ;
        RECT 129.200 188.800 130.000 190.400 ;
        RECT 130.800 188.800 131.600 190.400 ;
        RECT 132.400 189.000 133.000 191.000 ;
        RECT 116.400 187.800 117.400 188.200 ;
        RECT 107.600 187.200 108.400 187.600 ;
        RECT 102.200 186.600 106.000 187.200 ;
        RECT 102.200 186.400 103.000 186.600 ;
        RECT 90.800 184.200 91.600 185.000 ;
        RECT 92.400 184.800 93.200 185.600 ;
        RECT 94.200 185.400 95.000 185.600 ;
        RECT 94.200 184.800 97.000 185.400 ;
        RECT 96.400 184.200 97.000 184.800 ;
        RECT 100.400 184.200 101.200 185.000 ;
        RECT 90.800 183.600 92.800 184.200 ;
        RECT 92.000 182.200 92.800 183.600 ;
        RECT 96.400 182.200 97.200 184.200 ;
        RECT 100.400 183.600 101.800 184.200 ;
        RECT 100.600 182.200 101.800 183.600 ;
        RECT 105.200 182.200 106.000 186.600 ;
        RECT 107.000 186.200 110.600 186.600 ;
        RECT 111.600 186.200 112.200 187.600 ;
        RECT 113.200 187.200 117.400 187.800 ;
        RECT 118.400 187.600 120.400 188.400 ;
        RECT 122.800 187.600 125.400 188.400 ;
        RECT 127.600 188.200 128.400 188.400 ;
        RECT 126.800 187.600 128.400 188.200 ;
        RECT 132.400 188.200 133.800 189.000 ;
        RECT 134.400 188.400 135.000 192.200 ;
        RECT 138.800 192.400 139.600 199.800 ;
        RECT 142.000 192.800 142.800 199.800 ;
        RECT 138.800 191.800 141.400 192.400 ;
        RECT 142.000 191.800 143.000 192.800 ;
        RECT 135.600 189.600 136.400 191.200 ;
        RECT 138.800 189.600 139.800 190.400 ;
        RECT 139.000 188.800 139.800 189.600 ;
        RECT 140.800 189.800 141.400 191.800 ;
        RECT 140.800 189.000 141.800 189.800 ;
        RECT 132.400 187.800 133.400 188.200 ;
        RECT 106.800 186.000 110.800 186.200 ;
        RECT 106.800 182.200 107.600 186.000 ;
        RECT 110.000 182.200 110.800 186.000 ;
        RECT 111.600 182.200 112.400 186.200 ;
        RECT 113.200 185.000 113.800 187.200 ;
        RECT 118.400 187.000 119.000 187.600 ;
        RECT 118.200 186.600 119.000 187.000 ;
        RECT 117.400 186.000 119.000 186.600 ;
        RECT 123.000 186.200 123.600 187.600 ;
        RECT 126.800 187.200 127.600 187.600 ;
        RECT 129.200 187.200 133.400 187.800 ;
        RECT 134.400 187.600 136.400 188.400 ;
        RECT 124.600 186.200 128.200 186.600 ;
        RECT 113.200 183.000 114.000 185.000 ;
        RECT 117.400 183.000 118.200 186.000 ;
        RECT 122.800 182.200 123.600 186.200 ;
        RECT 124.400 186.000 128.400 186.200 ;
        RECT 124.400 182.200 125.200 186.000 ;
        RECT 127.600 182.200 128.400 186.000 ;
        RECT 129.200 185.000 129.800 187.200 ;
        RECT 134.400 187.000 135.000 187.600 ;
        RECT 140.800 187.400 141.400 189.000 ;
        RECT 142.400 188.400 143.000 191.800 ;
        RECT 142.000 187.600 143.000 188.400 ;
        RECT 134.200 186.600 135.000 187.000 ;
        RECT 133.400 186.000 135.000 186.600 ;
        RECT 138.800 186.800 141.400 187.400 ;
        RECT 129.200 183.000 130.000 185.000 ;
        RECT 133.400 183.000 134.200 186.000 ;
        RECT 138.800 182.200 139.600 186.800 ;
        RECT 142.400 186.200 143.000 187.600 ;
        RECT 142.000 185.600 143.000 186.200 ;
        RECT 142.000 182.200 142.800 185.600 ;
        RECT 145.200 182.200 146.000 199.800 ;
        RECT 151.000 192.600 151.800 199.800 ;
        RECT 150.000 191.800 151.800 192.600 ;
        RECT 150.200 188.400 150.800 191.800 ;
        RECT 151.600 189.600 152.400 191.200 ;
        RECT 150.000 187.600 150.800 188.400 ;
        RECT 150.200 186.400 150.800 187.600 ;
        RECT 146.800 186.300 147.600 186.400 ;
        RECT 148.400 186.300 149.200 186.400 ;
        RECT 146.800 185.700 149.200 186.300 ;
        RECT 146.800 184.800 147.600 185.700 ;
        RECT 148.400 184.800 149.200 185.700 ;
        RECT 150.000 185.600 150.800 186.400 ;
        RECT 150.200 184.200 150.800 185.600 ;
        RECT 150.000 182.200 150.800 184.200 ;
        RECT 156.400 184.300 157.200 184.400 ;
        RECT 158.000 184.300 158.800 199.800 ;
        RECT 161.200 192.400 162.000 199.800 ;
        RECT 162.600 192.400 163.400 192.600 ;
        RECT 161.200 191.800 163.400 192.400 ;
        RECT 165.600 192.400 167.200 199.800 ;
        RECT 169.200 192.400 170.000 192.600 ;
        RECT 170.800 192.400 171.600 199.800 ;
        RECT 165.600 191.800 167.600 192.400 ;
        RECT 169.200 191.800 171.600 192.400 ;
        RECT 174.000 192.000 174.800 199.800 ;
        RECT 177.200 195.200 178.000 199.800 ;
        RECT 162.800 191.200 163.400 191.800 ;
        RECT 162.800 190.600 166.200 191.200 ;
        RECT 165.400 190.400 166.200 190.600 ;
        RECT 167.000 190.400 167.600 191.800 ;
        RECT 173.800 191.200 174.800 192.000 ;
        RECT 175.400 194.600 178.000 195.200 ;
        RECT 175.400 193.000 176.000 194.600 ;
        RECT 180.400 194.400 181.200 199.800 ;
        RECT 183.600 197.000 184.400 199.800 ;
        RECT 185.200 197.000 186.000 199.800 ;
        RECT 186.800 197.000 187.600 199.800 ;
        RECT 181.800 194.400 186.000 195.200 ;
        RECT 178.600 193.600 181.200 194.400 ;
        RECT 188.400 193.600 189.200 199.800 ;
        RECT 191.600 195.000 192.400 199.800 ;
        RECT 194.800 195.000 195.600 199.800 ;
        RECT 196.400 197.000 197.200 199.800 ;
        RECT 198.000 197.000 198.800 199.800 ;
        RECT 201.200 195.200 202.000 199.800 ;
        RECT 204.400 196.400 205.200 199.800 ;
        RECT 204.400 195.800 205.400 196.400 ;
        RECT 204.800 195.200 205.400 195.800 ;
        RECT 200.000 194.400 204.200 195.200 ;
        RECT 204.800 194.600 206.800 195.200 ;
        RECT 191.600 193.600 194.200 194.400 ;
        RECT 194.800 193.800 200.600 194.400 ;
        RECT 203.600 194.000 204.200 194.400 ;
        RECT 183.600 193.000 184.400 193.200 ;
        RECT 175.400 192.400 184.400 193.000 ;
        RECT 186.800 193.000 187.600 193.200 ;
        RECT 194.800 193.000 195.400 193.800 ;
        RECT 201.200 193.200 202.600 193.800 ;
        RECT 203.600 193.200 205.200 194.000 ;
        RECT 186.800 192.400 195.400 193.000 ;
        RECT 196.400 193.000 202.600 193.200 ;
        RECT 196.400 192.600 201.800 193.000 ;
        RECT 196.400 192.400 197.200 192.600 ;
        RECT 167.000 190.300 168.400 190.400 ;
        RECT 172.400 190.300 173.200 190.400 ;
        RECT 163.200 189.800 164.000 190.000 ;
        RECT 167.000 189.800 173.200 190.300 ;
        RECT 163.200 189.200 165.800 189.800 ;
        RECT 165.200 188.600 165.800 189.200 ;
        RECT 166.600 189.700 173.200 189.800 ;
        RECT 166.600 189.600 168.400 189.700 ;
        RECT 172.400 189.600 173.200 189.700 ;
        RECT 166.600 189.200 167.600 189.600 ;
        RECT 161.200 188.200 162.800 188.400 ;
        RECT 161.200 187.600 164.600 188.200 ;
        RECT 165.200 187.800 166.000 188.600 ;
        RECT 164.000 187.200 164.600 187.600 ;
        RECT 162.600 186.800 163.400 187.000 ;
        RECT 159.600 184.800 160.400 186.400 ;
        RECT 161.200 186.200 163.400 186.800 ;
        RECT 164.000 186.600 166.000 187.200 ;
        RECT 164.400 186.400 166.000 186.600 ;
        RECT 156.400 183.700 158.800 184.300 ;
        RECT 156.400 183.600 157.200 183.700 ;
        RECT 158.000 182.200 158.800 183.700 ;
        RECT 161.200 182.200 162.000 186.200 ;
        RECT 166.600 185.800 167.200 189.200 ;
        RECT 168.000 187.600 168.800 188.400 ;
        RECT 170.000 188.300 171.600 188.400 ;
        RECT 173.800 188.300 174.600 191.200 ;
        RECT 175.400 190.600 176.000 192.400 ;
        RECT 170.000 187.700 174.600 188.300 ;
        RECT 170.000 187.600 171.600 187.700 ;
        RECT 168.000 187.200 168.600 187.600 ;
        RECT 167.800 186.400 168.600 187.200 ;
        RECT 169.200 186.800 170.000 187.000 ;
        RECT 173.800 186.800 174.600 187.700 ;
        RECT 175.200 190.000 176.000 190.600 ;
        RECT 182.000 190.000 205.400 190.600 ;
        RECT 175.200 188.000 175.800 190.000 ;
        RECT 182.000 189.400 182.800 190.000 ;
        RECT 199.600 189.600 200.400 190.000 ;
        RECT 204.400 189.800 205.400 190.000 ;
        RECT 204.400 189.600 205.200 189.800 ;
        RECT 176.400 188.600 180.200 189.400 ;
        RECT 175.200 187.400 176.400 188.000 ;
        RECT 169.200 186.200 171.600 186.800 ;
        RECT 165.600 182.200 167.200 185.800 ;
        RECT 170.800 182.200 171.600 186.200 ;
        RECT 173.800 186.000 174.800 186.800 ;
        RECT 174.000 182.200 174.800 186.000 ;
        RECT 175.600 182.200 176.400 187.400 ;
        RECT 179.400 187.400 180.200 188.600 ;
        RECT 179.400 186.800 181.200 187.400 ;
        RECT 180.400 186.200 181.200 186.800 ;
        RECT 185.200 186.400 186.000 189.200 ;
        RECT 188.400 188.600 191.600 189.400 ;
        RECT 195.400 188.600 197.400 189.400 ;
        RECT 206.000 189.000 206.800 194.600 ;
        RECT 207.600 191.600 208.400 193.200 ;
        RECT 188.000 187.800 188.800 188.000 ;
        RECT 188.000 187.200 192.400 187.800 ;
        RECT 191.600 187.000 192.400 187.200 ;
        RECT 193.200 186.800 194.000 188.400 ;
        RECT 180.400 185.400 182.800 186.200 ;
        RECT 185.200 185.600 186.200 186.400 ;
        RECT 189.200 185.600 190.800 186.400 ;
        RECT 191.600 186.200 192.400 186.400 ;
        RECT 195.400 186.200 196.200 188.600 ;
        RECT 198.000 188.200 206.800 189.000 ;
        RECT 201.400 186.800 204.400 187.600 ;
        RECT 201.400 186.200 202.200 186.800 ;
        RECT 191.600 185.600 196.200 186.200 ;
        RECT 182.000 182.200 182.800 185.400 ;
        RECT 199.600 185.400 202.200 186.200 ;
        RECT 183.600 182.200 184.400 185.000 ;
        RECT 185.200 182.200 186.000 185.000 ;
        RECT 186.800 182.200 187.600 185.000 ;
        RECT 188.400 182.200 189.200 185.000 ;
        RECT 191.600 182.200 192.400 185.000 ;
        RECT 194.800 182.200 195.600 185.000 ;
        RECT 196.400 182.200 197.200 185.000 ;
        RECT 198.000 182.200 198.800 185.000 ;
        RECT 199.600 182.200 200.400 185.400 ;
        RECT 206.000 182.200 206.800 188.200 ;
        RECT 209.200 186.200 210.000 199.800 ;
        RECT 215.000 192.400 215.800 199.800 ;
        RECT 216.400 193.600 218.000 194.400 ;
        RECT 216.600 192.400 217.200 193.600 ;
        RECT 218.800 192.400 219.600 199.800 ;
        RECT 215.000 191.800 216.000 192.400 ;
        RECT 216.600 191.800 218.000 192.400 ;
        RECT 218.800 191.800 221.000 192.400 ;
        RECT 222.000 191.800 222.800 199.800 ;
        RECT 214.000 188.800 214.800 190.400 ;
        RECT 215.400 188.400 216.000 191.800 ;
        RECT 217.200 191.600 218.000 191.800 ;
        RECT 220.400 191.200 221.000 191.800 ;
        RECT 220.400 190.400 221.600 191.200 ;
        RECT 218.800 188.800 219.600 190.400 ;
        RECT 210.800 186.800 211.600 188.400 ;
        RECT 212.400 188.200 213.200 188.400 ;
        RECT 212.400 187.600 214.000 188.200 ;
        RECT 215.400 187.600 218.000 188.400 ;
        RECT 213.200 187.200 214.000 187.600 ;
        RECT 212.600 186.200 216.200 186.600 ;
        RECT 217.200 186.200 217.800 187.600 ;
        RECT 220.400 187.400 221.000 190.400 ;
        RECT 222.200 189.600 222.800 191.800 ;
        RECT 218.800 186.800 221.000 187.400 ;
        RECT 222.000 188.300 222.800 189.600 ;
        RECT 225.200 191.200 226.000 199.800 ;
        RECT 228.400 191.200 229.200 199.800 ;
        RECT 234.200 192.400 235.000 199.800 ;
        RECT 235.600 193.600 237.200 194.400 ;
        RECT 235.800 192.400 236.400 193.600 ;
        RECT 240.600 192.400 241.400 199.800 ;
        RECT 242.000 194.300 242.800 194.400 ;
        RECT 244.400 194.300 245.200 194.400 ;
        RECT 242.000 193.700 245.200 194.300 ;
        RECT 242.000 193.600 242.800 193.700 ;
        RECT 244.400 193.600 245.200 193.700 ;
        RECT 242.200 192.400 242.800 193.600 ;
        RECT 234.200 191.800 235.200 192.400 ;
        RECT 235.800 191.800 237.200 192.400 ;
        RECT 240.600 191.800 241.600 192.400 ;
        RECT 242.200 191.800 243.600 192.400 ;
        RECT 225.200 190.400 229.200 191.200 ;
        RECT 234.600 190.400 235.200 191.800 ;
        RECT 236.400 191.600 237.200 191.800 ;
        RECT 223.600 188.300 224.400 188.400 ;
        RECT 222.000 187.700 224.400 188.300 ;
        RECT 208.200 185.600 210.000 186.200 ;
        RECT 212.400 186.000 216.400 186.200 ;
        RECT 208.200 182.200 209.000 185.600 ;
        RECT 212.400 182.200 213.200 186.000 ;
        RECT 215.600 182.200 216.400 186.000 ;
        RECT 217.200 182.200 218.000 186.200 ;
        RECT 218.800 182.200 219.600 186.800 ;
        RECT 222.000 182.200 222.800 187.700 ;
        RECT 223.600 187.600 224.400 187.700 ;
        RECT 225.200 187.600 226.000 190.400 ;
        RECT 233.200 188.800 234.000 190.400 ;
        RECT 234.600 189.600 235.600 190.400 ;
        RECT 234.600 188.400 235.200 189.600 ;
        RECT 239.600 188.800 240.400 190.400 ;
        RECT 241.000 188.400 241.600 191.800 ;
        RECT 242.800 191.600 243.600 191.800 ;
        RECT 231.600 188.200 232.400 188.400 ;
        RECT 231.600 187.600 233.200 188.200 ;
        RECT 234.600 187.600 237.200 188.400 ;
        RECT 238.000 188.200 238.800 188.400 ;
        RECT 241.000 188.300 243.600 188.400 ;
        RECT 244.400 188.300 245.200 188.400 ;
        RECT 238.000 187.600 239.600 188.200 ;
        RECT 241.000 187.700 245.200 188.300 ;
        RECT 241.000 187.600 243.600 187.700 ;
        RECT 225.200 186.800 229.200 187.600 ;
        RECT 232.400 187.200 233.200 187.600 ;
        RECT 225.200 182.200 226.000 186.800 ;
        RECT 228.400 182.200 229.200 186.800 ;
        RECT 231.800 186.200 235.400 186.600 ;
        RECT 236.400 186.200 237.000 187.600 ;
        RECT 238.800 187.200 239.600 187.600 ;
        RECT 238.200 186.200 241.800 186.600 ;
        RECT 242.800 186.200 243.400 187.600 ;
        RECT 244.400 186.800 245.200 187.700 ;
        RECT 246.000 188.300 246.800 199.800 ;
        RECT 247.600 191.600 248.400 193.200 ;
        RECT 250.800 192.800 251.600 199.800 ;
        RECT 250.600 191.800 251.600 192.800 ;
        RECT 254.000 192.400 254.800 199.800 ;
        RECT 257.200 196.400 258.000 199.800 ;
        RECT 257.000 195.800 258.000 196.400 ;
        RECT 257.000 195.200 257.600 195.800 ;
        RECT 260.400 195.200 261.200 199.800 ;
        RECT 263.600 197.000 264.400 199.800 ;
        RECT 265.200 197.000 266.000 199.800 ;
        RECT 252.200 191.800 254.800 192.400 ;
        RECT 255.600 194.600 257.600 195.200 ;
        RECT 250.600 188.400 251.200 191.800 ;
        RECT 252.200 189.800 252.800 191.800 ;
        RECT 251.800 189.000 252.800 189.800 ;
        RECT 247.600 188.300 248.400 188.400 ;
        RECT 246.000 187.700 248.400 188.300 ;
        RECT 246.000 186.200 246.800 187.700 ;
        RECT 247.600 187.600 248.400 187.700 ;
        RECT 249.200 188.300 250.000 188.400 ;
        RECT 250.600 188.300 251.600 188.400 ;
        RECT 249.200 187.700 251.600 188.300 ;
        RECT 249.200 187.600 250.000 187.700 ;
        RECT 250.600 187.600 251.600 187.700 ;
        RECT 250.600 186.200 251.200 187.600 ;
        RECT 252.200 187.400 252.800 189.000 ;
        RECT 253.800 189.600 254.800 190.400 ;
        RECT 253.800 188.800 254.600 189.600 ;
        RECT 255.600 189.000 256.400 194.600 ;
        RECT 258.200 194.400 262.400 195.200 ;
        RECT 266.800 195.000 267.600 199.800 ;
        RECT 270.000 195.000 270.800 199.800 ;
        RECT 258.200 194.000 258.800 194.400 ;
        RECT 257.200 193.200 258.800 194.000 ;
        RECT 261.800 193.800 267.600 194.400 ;
        RECT 259.800 193.200 261.200 193.800 ;
        RECT 259.800 193.000 266.000 193.200 ;
        RECT 260.600 192.600 266.000 193.000 ;
        RECT 265.200 192.400 266.000 192.600 ;
        RECT 267.000 193.000 267.600 193.800 ;
        RECT 268.200 193.600 270.800 194.400 ;
        RECT 273.200 193.600 274.000 199.800 ;
        RECT 274.800 197.000 275.600 199.800 ;
        RECT 276.400 197.000 277.200 199.800 ;
        RECT 278.000 197.000 278.800 199.800 ;
        RECT 276.400 194.400 280.600 195.200 ;
        RECT 281.200 194.400 282.000 199.800 ;
        RECT 284.400 195.200 285.200 199.800 ;
        RECT 284.400 194.600 287.000 195.200 ;
        RECT 281.200 193.600 283.800 194.400 ;
        RECT 274.800 193.000 275.600 193.200 ;
        RECT 267.000 192.400 275.600 193.000 ;
        RECT 278.000 193.000 278.800 193.200 ;
        RECT 286.400 193.000 287.000 194.600 ;
        RECT 278.000 192.400 287.000 193.000 ;
        RECT 286.400 190.600 287.000 192.400 ;
        RECT 287.600 192.000 288.400 199.800 ;
        RECT 291.600 193.600 292.400 194.400 ;
        RECT 291.600 192.400 292.200 193.600 ;
        RECT 293.000 192.400 293.800 199.800 ;
        RECT 289.200 192.300 290.000 192.400 ;
        RECT 290.800 192.300 292.200 192.400 ;
        RECT 287.600 191.200 288.600 192.000 ;
        RECT 289.200 191.800 292.200 192.300 ;
        RECT 292.800 191.800 293.800 192.400 ;
        RECT 297.200 192.400 298.000 199.800 ;
        RECT 300.400 192.800 301.200 199.800 ;
        RECT 297.200 191.800 299.800 192.400 ;
        RECT 300.400 191.800 301.400 192.800 ;
        RECT 289.200 191.700 291.600 191.800 ;
        RECT 289.200 191.600 290.000 191.700 ;
        RECT 290.800 191.600 291.600 191.700 ;
        RECT 257.000 190.000 280.400 190.600 ;
        RECT 286.400 190.000 287.200 190.600 ;
        RECT 257.000 189.800 257.800 190.000 ;
        RECT 258.800 189.600 259.600 190.000 ;
        RECT 262.000 189.600 262.800 190.000 ;
        RECT 279.600 189.400 280.400 190.000 ;
        RECT 255.600 188.200 264.400 189.000 ;
        RECT 265.000 188.600 267.000 189.400 ;
        RECT 270.800 188.600 274.000 189.400 ;
        RECT 252.200 186.800 254.800 187.400 ;
        RECT 231.600 186.000 235.600 186.200 ;
        RECT 231.600 182.200 232.400 186.000 ;
        RECT 234.800 182.200 235.600 186.000 ;
        RECT 236.400 182.200 237.200 186.200 ;
        RECT 238.000 186.000 242.000 186.200 ;
        RECT 238.000 182.200 238.800 186.000 ;
        RECT 241.200 182.200 242.000 186.000 ;
        RECT 242.800 182.200 243.600 186.200 ;
        RECT 246.000 185.600 247.800 186.200 ;
        RECT 250.600 185.600 251.600 186.200 ;
        RECT 247.000 182.200 247.800 185.600 ;
        RECT 250.800 182.200 251.600 185.600 ;
        RECT 254.000 182.200 254.800 186.800 ;
        RECT 255.600 182.200 256.400 188.200 ;
        RECT 258.000 186.800 261.000 187.600 ;
        RECT 260.200 186.200 261.000 186.800 ;
        RECT 266.200 186.200 267.000 188.600 ;
        RECT 268.400 186.800 269.200 188.400 ;
        RECT 273.600 187.800 274.400 188.000 ;
        RECT 270.000 187.200 274.400 187.800 ;
        RECT 270.000 187.000 270.800 187.200 ;
        RECT 276.400 186.400 277.200 189.200 ;
        RECT 282.200 188.600 286.000 189.400 ;
        RECT 282.200 187.400 283.000 188.600 ;
        RECT 286.600 188.000 287.200 190.000 ;
        RECT 270.000 186.200 270.800 186.400 ;
        RECT 260.200 185.400 262.800 186.200 ;
        RECT 266.200 185.600 270.800 186.200 ;
        RECT 271.600 185.600 273.200 186.400 ;
        RECT 276.200 185.600 277.200 186.400 ;
        RECT 281.200 186.800 283.000 187.400 ;
        RECT 286.000 187.400 287.200 188.000 ;
        RECT 281.200 186.200 282.000 186.800 ;
        RECT 262.000 182.200 262.800 185.400 ;
        RECT 279.600 185.400 282.000 186.200 ;
        RECT 263.600 182.200 264.400 185.000 ;
        RECT 265.200 182.200 266.000 185.000 ;
        RECT 266.800 182.200 267.600 185.000 ;
        RECT 270.000 182.200 270.800 185.000 ;
        RECT 273.200 182.200 274.000 185.000 ;
        RECT 274.800 182.200 275.600 185.000 ;
        RECT 276.400 182.200 277.200 185.000 ;
        RECT 278.000 182.200 278.800 185.000 ;
        RECT 279.600 182.200 280.400 185.400 ;
        RECT 286.000 182.200 286.800 187.400 ;
        RECT 287.800 186.800 288.600 191.200 ;
        RECT 292.800 188.400 293.400 191.800 ;
        RECT 294.000 188.800 294.800 190.400 ;
        RECT 295.600 190.300 296.400 190.400 ;
        RECT 297.200 190.300 298.200 190.400 ;
        RECT 295.600 189.700 298.200 190.300 ;
        RECT 295.600 189.600 296.400 189.700 ;
        RECT 297.200 189.600 298.200 189.700 ;
        RECT 297.400 188.800 298.200 189.600 ;
        RECT 299.200 189.800 299.800 191.800 ;
        RECT 299.200 189.000 300.200 189.800 ;
        RECT 290.800 187.600 293.400 188.400 ;
        RECT 295.600 188.200 296.400 188.400 ;
        RECT 294.800 187.600 296.400 188.200 ;
        RECT 287.600 186.000 288.600 186.800 ;
        RECT 291.000 186.200 291.600 187.600 ;
        RECT 294.800 187.200 295.600 187.600 ;
        RECT 299.200 187.400 299.800 189.000 ;
        RECT 300.800 188.400 301.400 191.800 ;
        RECT 300.400 187.600 301.400 188.400 ;
        RECT 297.200 186.800 299.800 187.400 ;
        RECT 292.600 186.200 296.200 186.600 ;
        RECT 287.600 182.200 288.400 186.000 ;
        RECT 290.800 182.200 291.600 186.200 ;
        RECT 292.400 186.000 296.400 186.200 ;
        RECT 292.400 182.200 293.200 186.000 ;
        RECT 295.600 182.200 296.400 186.000 ;
        RECT 297.200 182.200 298.000 186.800 ;
        RECT 300.800 186.200 301.400 187.600 ;
        RECT 300.400 185.600 301.400 186.200 ;
        RECT 300.400 182.200 301.200 185.600 ;
        RECT 308.400 184.800 309.200 186.400 ;
        RECT 310.000 182.200 310.800 199.800 ;
        RECT 314.200 192.600 315.000 199.800 ;
        RECT 313.200 191.800 315.000 192.600 ;
        RECT 319.000 192.400 319.800 199.800 ;
        RECT 320.400 194.300 321.200 194.400 ;
        RECT 324.400 194.300 325.200 199.800 ;
        RECT 327.600 195.200 328.400 199.800 ;
        RECT 320.400 193.700 325.200 194.300 ;
        RECT 320.400 193.600 321.200 193.700 ;
        RECT 320.600 192.400 321.200 193.600 ;
        RECT 319.000 191.800 320.000 192.400 ;
        RECT 320.600 191.800 322.000 192.400 ;
        RECT 324.400 192.000 325.200 193.700 ;
        RECT 313.400 190.400 314.000 191.800 ;
        RECT 313.200 189.600 314.000 190.400 ;
        RECT 314.800 189.600 315.600 191.200 ;
        RECT 313.400 188.400 314.000 189.600 ;
        RECT 318.000 188.800 318.800 190.400 ;
        RECT 319.400 188.400 320.000 191.800 ;
        RECT 321.200 191.600 322.000 191.800 ;
        RECT 324.200 191.200 325.200 192.000 ;
        RECT 325.800 194.600 328.400 195.200 ;
        RECT 325.800 193.000 326.400 194.600 ;
        RECT 330.800 194.400 331.600 199.800 ;
        RECT 334.000 197.000 334.800 199.800 ;
        RECT 335.600 197.000 336.400 199.800 ;
        RECT 337.200 197.000 338.000 199.800 ;
        RECT 332.200 194.400 336.400 195.200 ;
        RECT 329.000 193.600 331.600 194.400 ;
        RECT 338.800 193.600 339.600 199.800 ;
        RECT 342.000 195.000 342.800 199.800 ;
        RECT 345.200 195.000 346.000 199.800 ;
        RECT 346.800 197.000 347.600 199.800 ;
        RECT 348.400 197.000 349.200 199.800 ;
        RECT 351.600 195.200 352.400 199.800 ;
        RECT 354.800 196.400 355.600 199.800 ;
        RECT 354.800 195.800 355.800 196.400 ;
        RECT 355.200 195.200 355.800 195.800 ;
        RECT 350.400 194.400 354.600 195.200 ;
        RECT 355.200 194.600 357.200 195.200 ;
        RECT 342.000 193.600 344.600 194.400 ;
        RECT 345.200 193.800 351.000 194.400 ;
        RECT 354.000 194.000 354.600 194.400 ;
        RECT 334.000 193.000 334.800 193.200 ;
        RECT 325.800 192.400 334.800 193.000 ;
        RECT 337.200 193.000 338.000 193.200 ;
        RECT 345.200 193.000 345.800 193.800 ;
        RECT 351.600 193.200 353.000 193.800 ;
        RECT 354.000 193.200 355.600 194.000 ;
        RECT 337.200 192.400 345.800 193.000 ;
        RECT 346.800 193.000 353.000 193.200 ;
        RECT 346.800 192.600 352.200 193.000 ;
        RECT 346.800 192.400 347.600 192.600 ;
        RECT 313.200 187.600 314.000 188.400 ;
        RECT 316.400 188.200 317.200 188.400 ;
        RECT 316.400 187.600 318.000 188.200 ;
        RECT 319.400 187.600 322.000 188.400 ;
        RECT 311.600 184.800 312.400 186.400 ;
        RECT 313.400 184.200 314.000 187.600 ;
        RECT 317.200 187.200 318.000 187.600 ;
        RECT 316.600 186.200 320.200 186.600 ;
        RECT 321.200 186.200 321.800 187.600 ;
        RECT 324.200 186.800 325.000 191.200 ;
        RECT 325.800 190.600 326.400 192.400 ;
        RECT 325.600 190.000 326.400 190.600 ;
        RECT 332.400 190.000 355.800 190.600 ;
        RECT 325.600 188.000 326.200 190.000 ;
        RECT 332.400 189.400 333.200 190.000 ;
        RECT 350.000 189.600 350.800 190.000 ;
        RECT 355.000 189.800 355.800 190.000 ;
        RECT 326.800 188.600 330.600 189.400 ;
        RECT 325.600 187.400 326.800 188.000 ;
        RECT 313.200 182.200 314.000 184.200 ;
        RECT 316.400 186.000 320.400 186.200 ;
        RECT 316.400 182.200 317.200 186.000 ;
        RECT 319.600 182.200 320.400 186.000 ;
        RECT 321.200 182.200 322.000 186.200 ;
        RECT 324.200 186.000 325.200 186.800 ;
        RECT 324.400 182.200 325.200 186.000 ;
        RECT 326.000 182.200 326.800 187.400 ;
        RECT 329.800 187.400 330.600 188.600 ;
        RECT 329.800 186.800 331.600 187.400 ;
        RECT 330.800 186.200 331.600 186.800 ;
        RECT 335.600 186.400 336.400 189.200 ;
        RECT 338.800 188.600 342.000 189.400 ;
        RECT 345.800 188.600 347.800 189.400 ;
        RECT 356.400 189.000 357.200 194.600 ;
        RECT 358.000 193.600 359.600 194.400 ;
        RECT 358.800 192.400 359.400 193.600 ;
        RECT 360.200 192.400 361.000 199.800 ;
        RECT 358.000 191.800 359.400 192.400 ;
        RECT 360.000 191.800 361.000 192.400 ;
        RECT 366.000 192.000 366.800 199.800 ;
        RECT 369.200 195.200 370.000 199.800 ;
        RECT 358.000 191.600 358.800 191.800 ;
        RECT 338.400 187.800 339.200 188.000 ;
        RECT 338.400 187.200 342.800 187.800 ;
        RECT 342.000 187.000 342.800 187.200 ;
        RECT 343.600 186.800 344.400 188.400 ;
        RECT 330.800 185.400 333.200 186.200 ;
        RECT 335.600 185.600 336.600 186.400 ;
        RECT 339.600 185.600 341.200 186.400 ;
        RECT 342.000 186.200 342.800 186.400 ;
        RECT 345.800 186.200 346.600 188.600 ;
        RECT 348.400 188.200 357.200 189.000 ;
        RECT 360.000 188.400 360.600 191.800 ;
        RECT 365.800 191.200 366.800 192.000 ;
        RECT 367.400 194.600 370.000 195.200 ;
        RECT 367.400 193.000 368.000 194.600 ;
        RECT 372.400 194.400 373.200 199.800 ;
        RECT 375.600 197.000 376.400 199.800 ;
        RECT 377.200 197.000 378.000 199.800 ;
        RECT 378.800 197.000 379.600 199.800 ;
        RECT 373.800 194.400 378.000 195.200 ;
        RECT 370.600 193.600 373.200 194.400 ;
        RECT 380.400 193.600 381.200 199.800 ;
        RECT 383.600 195.000 384.400 199.800 ;
        RECT 386.800 195.000 387.600 199.800 ;
        RECT 388.400 197.000 389.200 199.800 ;
        RECT 390.000 197.000 390.800 199.800 ;
        RECT 393.200 195.200 394.000 199.800 ;
        RECT 396.400 196.400 397.200 199.800 ;
        RECT 401.200 196.400 402.000 199.800 ;
        RECT 396.400 195.800 397.400 196.400 ;
        RECT 396.800 195.200 397.400 195.800 ;
        RECT 401.000 195.800 402.000 196.400 ;
        RECT 401.000 195.200 401.600 195.800 ;
        RECT 404.400 195.200 405.200 199.800 ;
        RECT 407.600 197.000 408.400 199.800 ;
        RECT 409.200 197.000 410.000 199.800 ;
        RECT 392.000 194.400 396.200 195.200 ;
        RECT 396.800 194.600 398.800 195.200 ;
        RECT 383.600 193.600 386.200 194.400 ;
        RECT 386.800 193.800 392.600 194.400 ;
        RECT 395.600 194.000 396.200 194.400 ;
        RECT 375.600 193.000 376.400 193.200 ;
        RECT 367.400 192.400 376.400 193.000 ;
        RECT 378.800 193.000 379.600 193.200 ;
        RECT 386.800 193.000 387.400 193.800 ;
        RECT 393.200 193.200 394.600 193.800 ;
        RECT 395.600 193.200 397.200 194.000 ;
        RECT 378.800 192.400 387.400 193.000 ;
        RECT 388.400 193.000 394.600 193.200 ;
        RECT 388.400 192.600 393.800 193.000 ;
        RECT 388.400 192.400 389.200 192.600 ;
        RECT 361.200 188.800 362.000 190.400 ;
        RECT 351.800 186.800 354.800 187.600 ;
        RECT 351.800 186.200 352.600 186.800 ;
        RECT 342.000 185.600 346.600 186.200 ;
        RECT 332.400 182.200 333.200 185.400 ;
        RECT 350.000 185.400 352.600 186.200 ;
        RECT 334.000 182.200 334.800 185.000 ;
        RECT 335.600 182.200 336.400 185.000 ;
        RECT 337.200 182.200 338.000 185.000 ;
        RECT 338.800 182.200 339.600 185.000 ;
        RECT 342.000 182.200 342.800 185.000 ;
        RECT 345.200 182.200 346.000 185.000 ;
        RECT 346.800 182.200 347.600 185.000 ;
        RECT 348.400 182.200 349.200 185.000 ;
        RECT 350.000 182.200 350.800 185.400 ;
        RECT 356.400 182.200 357.200 188.200 ;
        RECT 358.000 187.600 360.600 188.400 ;
        RECT 362.800 188.300 363.600 188.400 ;
        RECT 364.400 188.300 365.200 188.400 ;
        RECT 362.800 188.200 365.200 188.300 ;
        RECT 362.000 187.700 365.200 188.200 ;
        RECT 362.000 187.600 363.600 187.700 ;
        RECT 364.400 187.600 365.200 187.700 ;
        RECT 358.200 186.200 358.800 187.600 ;
        RECT 362.000 187.200 362.800 187.600 ;
        RECT 365.800 186.800 366.600 191.200 ;
        RECT 367.400 190.600 368.000 192.400 ;
        RECT 367.200 190.000 368.000 190.600 ;
        RECT 374.000 190.000 397.400 190.600 ;
        RECT 367.200 188.000 367.800 190.000 ;
        RECT 374.000 189.400 374.800 190.000 ;
        RECT 391.600 189.600 392.400 190.000 ;
        RECT 396.400 189.800 397.400 190.000 ;
        RECT 396.400 189.600 397.200 189.800 ;
        RECT 368.400 188.600 372.200 189.400 ;
        RECT 367.200 187.400 368.400 188.000 ;
        RECT 359.800 186.200 363.400 186.600 ;
        RECT 358.000 182.200 358.800 186.200 ;
        RECT 359.600 186.000 363.600 186.200 ;
        RECT 365.800 186.000 366.800 186.800 ;
        RECT 359.600 182.200 360.400 186.000 ;
        RECT 362.800 182.200 363.600 186.000 ;
        RECT 366.000 182.200 366.800 186.000 ;
        RECT 367.600 182.200 368.400 187.400 ;
        RECT 371.400 187.400 372.200 188.600 ;
        RECT 371.400 186.800 373.200 187.400 ;
        RECT 372.400 186.200 373.200 186.800 ;
        RECT 377.200 186.400 378.000 189.200 ;
        RECT 380.400 188.600 383.600 189.400 ;
        RECT 387.400 188.600 389.400 189.400 ;
        RECT 398.000 189.000 398.800 194.600 ;
        RECT 380.000 187.800 380.800 188.000 ;
        RECT 380.000 187.200 384.400 187.800 ;
        RECT 383.600 187.000 384.400 187.200 ;
        RECT 385.200 186.800 386.000 188.400 ;
        RECT 372.400 185.400 374.800 186.200 ;
        RECT 377.200 185.600 378.200 186.400 ;
        RECT 381.200 185.600 382.800 186.400 ;
        RECT 383.600 186.200 384.400 186.400 ;
        RECT 387.400 186.200 388.200 188.600 ;
        RECT 390.000 188.200 398.800 189.000 ;
        RECT 393.400 186.800 396.400 187.600 ;
        RECT 393.400 186.200 394.200 186.800 ;
        RECT 383.600 185.600 388.200 186.200 ;
        RECT 374.000 182.200 374.800 185.400 ;
        RECT 391.600 185.400 394.200 186.200 ;
        RECT 375.600 182.200 376.400 185.000 ;
        RECT 377.200 182.200 378.000 185.000 ;
        RECT 378.800 182.200 379.600 185.000 ;
        RECT 380.400 182.200 381.200 185.000 ;
        RECT 383.600 182.200 384.400 185.000 ;
        RECT 386.800 182.200 387.600 185.000 ;
        RECT 388.400 182.200 389.200 185.000 ;
        RECT 390.000 182.200 390.800 185.000 ;
        RECT 391.600 182.200 392.400 185.400 ;
        RECT 398.000 182.200 398.800 188.200 ;
        RECT 399.600 194.600 401.600 195.200 ;
        RECT 399.600 189.000 400.400 194.600 ;
        RECT 402.200 194.400 406.400 195.200 ;
        RECT 410.800 195.000 411.600 199.800 ;
        RECT 414.000 195.000 414.800 199.800 ;
        RECT 402.200 194.000 402.800 194.400 ;
        RECT 401.200 193.200 402.800 194.000 ;
        RECT 405.800 193.800 411.600 194.400 ;
        RECT 403.800 193.200 405.200 193.800 ;
        RECT 403.800 193.000 410.000 193.200 ;
        RECT 404.600 192.600 410.000 193.000 ;
        RECT 409.200 192.400 410.000 192.600 ;
        RECT 411.000 193.000 411.600 193.800 ;
        RECT 412.200 193.600 414.800 194.400 ;
        RECT 417.200 193.600 418.000 199.800 ;
        RECT 418.800 197.000 419.600 199.800 ;
        RECT 420.400 197.000 421.200 199.800 ;
        RECT 422.000 197.000 422.800 199.800 ;
        RECT 420.400 194.400 424.600 195.200 ;
        RECT 425.200 194.400 426.000 199.800 ;
        RECT 428.400 195.200 429.200 199.800 ;
        RECT 428.400 194.600 431.000 195.200 ;
        RECT 425.200 193.600 427.800 194.400 ;
        RECT 418.800 193.000 419.600 193.200 ;
        RECT 411.000 192.400 419.600 193.000 ;
        RECT 422.000 193.000 422.800 193.200 ;
        RECT 430.400 193.000 431.000 194.600 ;
        RECT 422.000 192.400 431.000 193.000 ;
        RECT 430.400 190.600 431.000 192.400 ;
        RECT 431.600 192.000 432.400 199.800 ;
        RECT 436.400 196.400 437.200 199.800 ;
        RECT 436.200 195.800 437.200 196.400 ;
        RECT 436.200 195.200 436.800 195.800 ;
        RECT 439.600 195.200 440.400 199.800 ;
        RECT 442.800 197.000 443.600 199.800 ;
        RECT 444.400 197.000 445.200 199.800 ;
        RECT 434.800 194.600 436.800 195.200 ;
        RECT 431.600 191.200 432.600 192.000 ;
        RECT 401.000 190.000 424.400 190.600 ;
        RECT 430.400 190.000 431.200 190.600 ;
        RECT 401.000 189.800 401.800 190.000 ;
        RECT 404.400 189.600 405.200 190.000 ;
        RECT 406.000 189.600 406.800 190.000 ;
        RECT 423.600 189.400 424.400 190.000 ;
        RECT 399.600 188.200 408.400 189.000 ;
        RECT 409.000 188.600 411.000 189.400 ;
        RECT 414.800 188.600 418.000 189.400 ;
        RECT 399.600 182.200 400.400 188.200 ;
        RECT 402.000 186.800 405.000 187.600 ;
        RECT 404.200 186.200 405.000 186.800 ;
        RECT 410.200 186.200 411.000 188.600 ;
        RECT 412.400 186.800 413.200 188.400 ;
        RECT 417.600 187.800 418.400 188.000 ;
        RECT 414.000 187.200 418.400 187.800 ;
        RECT 414.000 187.000 414.800 187.200 ;
        RECT 420.400 186.400 421.200 189.200 ;
        RECT 426.200 188.600 430.000 189.400 ;
        RECT 426.200 187.400 427.000 188.600 ;
        RECT 430.600 188.000 431.200 190.000 ;
        RECT 414.000 186.200 414.800 186.400 ;
        RECT 404.200 185.400 406.800 186.200 ;
        RECT 410.200 185.600 414.800 186.200 ;
        RECT 415.600 185.600 417.200 186.400 ;
        RECT 420.200 185.600 421.200 186.400 ;
        RECT 425.200 186.800 427.000 187.400 ;
        RECT 430.000 187.400 431.200 188.000 ;
        RECT 425.200 186.200 426.000 186.800 ;
        RECT 406.000 182.200 406.800 185.400 ;
        RECT 423.600 185.400 426.000 186.200 ;
        RECT 407.600 182.200 408.400 185.000 ;
        RECT 409.200 182.200 410.000 185.000 ;
        RECT 410.800 182.200 411.600 185.000 ;
        RECT 414.000 182.200 414.800 185.000 ;
        RECT 417.200 182.200 418.000 185.000 ;
        RECT 418.800 182.200 419.600 185.000 ;
        RECT 420.400 182.200 421.200 185.000 ;
        RECT 422.000 182.200 422.800 185.000 ;
        RECT 423.600 182.200 424.400 185.400 ;
        RECT 430.000 182.200 430.800 187.400 ;
        RECT 431.800 186.800 432.600 191.200 ;
        RECT 431.600 186.000 432.600 186.800 ;
        RECT 434.800 189.000 435.600 194.600 ;
        RECT 437.400 194.400 441.600 195.200 ;
        RECT 446.000 195.000 446.800 199.800 ;
        RECT 449.200 195.000 450.000 199.800 ;
        RECT 437.400 194.000 438.000 194.400 ;
        RECT 436.400 193.200 438.000 194.000 ;
        RECT 441.000 193.800 446.800 194.400 ;
        RECT 439.000 193.200 440.400 193.800 ;
        RECT 439.000 193.000 445.200 193.200 ;
        RECT 439.800 192.600 445.200 193.000 ;
        RECT 444.400 192.400 445.200 192.600 ;
        RECT 446.200 193.000 446.800 193.800 ;
        RECT 447.400 193.600 450.000 194.400 ;
        RECT 452.400 193.600 453.200 199.800 ;
        RECT 454.000 197.000 454.800 199.800 ;
        RECT 455.600 197.000 456.400 199.800 ;
        RECT 457.200 197.000 458.000 199.800 ;
        RECT 455.600 194.400 459.800 195.200 ;
        RECT 460.400 194.400 461.200 199.800 ;
        RECT 463.600 195.200 464.400 199.800 ;
        RECT 463.600 194.600 466.200 195.200 ;
        RECT 460.400 193.600 463.000 194.400 ;
        RECT 454.000 193.000 454.800 193.200 ;
        RECT 446.200 192.400 454.800 193.000 ;
        RECT 457.200 193.000 458.000 193.200 ;
        RECT 465.600 193.000 466.200 194.600 ;
        RECT 457.200 192.400 466.200 193.000 ;
        RECT 465.600 190.600 466.200 192.400 ;
        RECT 466.800 192.000 467.600 199.800 ;
        RECT 466.800 191.200 467.800 192.000 ;
        RECT 436.200 190.000 459.600 190.600 ;
        RECT 465.600 190.000 466.400 190.600 ;
        RECT 436.200 189.800 437.000 190.000 ;
        RECT 438.000 189.600 438.800 190.000 ;
        RECT 441.200 189.600 442.000 190.000 ;
        RECT 458.800 189.400 459.600 190.000 ;
        RECT 434.800 188.200 443.600 189.000 ;
        RECT 444.200 188.600 446.200 189.400 ;
        RECT 450.000 188.600 453.200 189.400 ;
        RECT 431.600 182.200 432.400 186.000 ;
        RECT 434.800 182.200 435.600 188.200 ;
        RECT 437.200 186.800 440.200 187.600 ;
        RECT 439.400 186.200 440.200 186.800 ;
        RECT 445.400 186.200 446.200 188.600 ;
        RECT 447.600 186.800 448.400 188.400 ;
        RECT 452.800 187.800 453.600 188.000 ;
        RECT 449.200 187.200 453.600 187.800 ;
        RECT 449.200 187.000 450.000 187.200 ;
        RECT 455.600 186.400 456.400 189.200 ;
        RECT 461.400 188.600 465.200 189.400 ;
        RECT 461.400 187.400 462.200 188.600 ;
        RECT 465.800 188.000 466.400 190.000 ;
        RECT 449.200 186.200 450.000 186.400 ;
        RECT 439.400 185.400 442.000 186.200 ;
        RECT 445.400 185.600 450.000 186.200 ;
        RECT 450.800 185.600 452.400 186.400 ;
        RECT 455.400 185.600 456.400 186.400 ;
        RECT 460.400 186.800 462.200 187.400 ;
        RECT 465.200 187.400 466.400 188.000 ;
        RECT 460.400 186.200 461.200 186.800 ;
        RECT 441.200 182.200 442.000 185.400 ;
        RECT 458.800 185.400 461.200 186.200 ;
        RECT 442.800 182.200 443.600 185.000 ;
        RECT 444.400 182.200 445.200 185.000 ;
        RECT 446.000 182.200 446.800 185.000 ;
        RECT 449.200 182.200 450.000 185.000 ;
        RECT 452.400 182.200 453.200 185.000 ;
        RECT 454.000 182.200 454.800 185.000 ;
        RECT 455.600 182.200 456.400 185.000 ;
        RECT 457.200 182.200 458.000 185.000 ;
        RECT 458.800 182.200 459.600 185.400 ;
        RECT 465.200 182.200 466.000 187.400 ;
        RECT 467.000 186.800 467.800 191.200 ;
        RECT 474.800 191.400 475.600 199.800 ;
        RECT 479.200 196.400 480.000 199.800 ;
        RECT 478.000 195.800 480.000 196.400 ;
        RECT 483.600 195.800 484.400 199.800 ;
        RECT 487.800 195.800 489.000 199.800 ;
        RECT 478.000 195.000 478.800 195.800 ;
        RECT 483.600 195.200 484.200 195.800 ;
        RECT 481.400 194.600 485.000 195.200 ;
        RECT 487.600 195.000 488.400 195.800 ;
        RECT 481.400 194.400 482.200 194.600 ;
        RECT 484.200 194.400 485.000 194.600 ;
        RECT 488.600 194.000 490.000 194.400 ;
        RECT 487.800 193.600 490.000 194.000 ;
        RECT 478.000 193.000 478.800 193.200 ;
        RECT 482.600 193.000 483.400 193.200 ;
        RECT 478.000 192.400 483.400 193.000 ;
        RECT 484.000 193.000 486.200 193.600 ;
        RECT 484.000 191.800 484.600 193.000 ;
        RECT 485.400 192.800 486.200 193.000 ;
        RECT 487.800 193.200 489.200 193.600 ;
        RECT 487.800 192.200 488.400 193.200 ;
        RECT 479.800 191.400 484.600 191.800 ;
        RECT 474.800 191.200 484.600 191.400 ;
        RECT 486.000 191.600 488.400 192.200 ;
        RECT 474.800 191.000 480.600 191.200 ;
        RECT 474.800 190.800 480.400 191.000 ;
        RECT 481.200 190.200 482.000 190.400 ;
        RECT 477.000 189.600 482.000 190.200 ;
        RECT 477.000 189.400 477.800 189.600 ;
        RECT 479.600 189.400 480.400 189.600 ;
        RECT 478.600 188.400 479.400 188.600 ;
        RECT 486.000 188.400 486.600 191.600 ;
        RECT 492.400 191.200 493.200 199.800 ;
        RECT 496.600 192.400 497.400 199.800 ;
        RECT 498.000 193.600 498.800 194.400 ;
        RECT 498.200 192.400 498.800 193.600 ;
        RECT 502.000 194.300 502.800 199.800 ;
        RECT 503.600 194.300 504.400 194.400 ;
        RECT 502.000 193.700 504.400 194.300 ;
        RECT 496.600 191.800 497.600 192.400 ;
        RECT 498.200 191.800 499.600 192.400 ;
        RECT 489.000 190.600 493.200 191.200 ;
        RECT 489.000 190.400 489.800 190.600 ;
        RECT 490.600 189.800 491.400 190.000 ;
        RECT 487.600 189.200 491.400 189.800 ;
        RECT 487.600 189.000 488.400 189.200 ;
        RECT 475.600 187.800 486.600 188.400 ;
        RECT 475.600 187.600 477.200 187.800 ;
        RECT 466.800 186.000 467.800 186.800 ;
        RECT 466.800 182.200 467.600 186.000 ;
        RECT 474.800 182.200 475.600 187.000 ;
        RECT 479.800 185.600 480.400 187.800 ;
        RECT 481.200 187.600 482.000 187.800 ;
        RECT 485.400 187.600 486.200 187.800 ;
        RECT 492.400 187.200 493.200 190.600 ;
        RECT 495.600 188.800 496.400 190.400 ;
        RECT 497.000 188.400 497.600 191.800 ;
        RECT 498.800 191.600 499.600 191.800 ;
        RECT 500.400 191.600 501.200 193.200 ;
        RECT 494.000 188.200 494.800 188.400 ;
        RECT 494.000 187.600 495.600 188.200 ;
        RECT 497.000 187.600 499.600 188.400 ;
        RECT 494.800 187.200 495.600 187.600 ;
        RECT 489.400 186.600 493.200 187.200 ;
        RECT 489.400 186.400 490.200 186.600 ;
        RECT 478.000 184.200 478.800 185.000 ;
        RECT 479.600 184.800 480.400 185.600 ;
        RECT 481.400 185.400 482.200 185.600 ;
        RECT 481.400 184.800 484.200 185.400 ;
        RECT 483.600 184.200 484.200 184.800 ;
        RECT 487.600 184.200 488.400 185.000 ;
        RECT 478.000 183.600 480.000 184.200 ;
        RECT 479.200 182.200 480.000 183.600 ;
        RECT 483.600 182.200 484.400 184.200 ;
        RECT 487.600 183.600 489.000 184.200 ;
        RECT 487.800 182.200 489.000 183.600 ;
        RECT 492.400 182.200 493.200 186.600 ;
        RECT 494.200 186.200 497.800 186.600 ;
        RECT 498.800 186.200 499.400 187.600 ;
        RECT 502.000 186.200 502.800 193.700 ;
        RECT 503.600 193.600 504.400 193.700 ;
        RECT 506.800 191.200 507.600 199.800 ;
        RECT 510.000 191.200 510.800 199.800 ;
        RECT 513.800 192.600 514.600 199.800 ;
        RECT 518.800 193.600 519.600 194.400 ;
        RECT 513.800 191.800 515.600 192.600 ;
        RECT 518.800 192.400 519.400 193.600 ;
        RECT 520.200 192.400 521.000 199.800 ;
        RECT 518.000 191.800 519.400 192.400 ;
        RECT 520.000 191.800 521.000 192.400 ;
        RECT 506.800 190.400 510.800 191.200 ;
        RECT 503.600 186.800 504.400 188.400 ;
        RECT 506.800 187.600 507.600 190.400 ;
        RECT 513.200 189.600 514.000 191.200 ;
        RECT 514.800 188.400 515.400 191.800 ;
        RECT 518.000 191.600 518.800 191.800 ;
        RECT 520.000 188.400 520.600 191.800 ;
        RECT 521.200 190.300 522.000 190.400 ;
        RECT 524.400 190.300 525.200 199.800 ;
        RECT 529.200 192.000 530.000 199.800 ;
        RECT 532.400 195.200 533.200 199.800 ;
        RECT 521.200 189.700 525.200 190.300 ;
        RECT 521.200 188.800 522.000 189.700 ;
        RECT 514.800 187.600 515.600 188.400 ;
        RECT 518.000 187.600 520.600 188.400 ;
        RECT 522.800 188.200 523.600 188.400 ;
        RECT 522.000 187.600 523.600 188.200 ;
        RECT 506.800 186.800 510.800 187.600 ;
        RECT 494.000 186.000 498.000 186.200 ;
        RECT 494.000 182.200 494.800 186.000 ;
        RECT 497.200 182.200 498.000 186.000 ;
        RECT 498.800 182.200 499.600 186.200 ;
        RECT 501.000 185.600 502.800 186.200 ;
        RECT 501.000 182.200 501.800 185.600 ;
        RECT 506.800 182.200 507.600 186.800 ;
        RECT 510.000 182.200 510.800 186.800 ;
        RECT 514.800 184.400 515.400 187.600 ;
        RECT 516.400 184.800 517.200 186.400 ;
        RECT 518.200 186.200 518.800 187.600 ;
        RECT 522.000 187.200 522.800 187.600 ;
        RECT 519.800 186.200 523.400 186.600 ;
        RECT 514.800 182.200 515.600 184.400 ;
        RECT 518.000 182.200 518.800 186.200 ;
        RECT 519.600 186.000 523.600 186.200 ;
        RECT 519.600 182.200 520.400 186.000 ;
        RECT 522.800 182.200 523.600 186.000 ;
        RECT 524.400 182.200 525.200 189.700 ;
        RECT 529.000 191.200 530.000 192.000 ;
        RECT 530.600 194.600 533.200 195.200 ;
        RECT 530.600 193.000 531.200 194.600 ;
        RECT 535.600 194.400 536.400 199.800 ;
        RECT 538.800 197.000 539.600 199.800 ;
        RECT 540.400 197.000 541.200 199.800 ;
        RECT 542.000 197.000 542.800 199.800 ;
        RECT 537.000 194.400 541.200 195.200 ;
        RECT 533.800 193.600 536.400 194.400 ;
        RECT 543.600 193.600 544.400 199.800 ;
        RECT 546.800 195.000 547.600 199.800 ;
        RECT 550.000 195.000 550.800 199.800 ;
        RECT 551.600 197.000 552.400 199.800 ;
        RECT 553.200 197.000 554.000 199.800 ;
        RECT 556.400 195.200 557.200 199.800 ;
        RECT 559.600 196.400 560.400 199.800 ;
        RECT 564.400 196.400 565.200 199.800 ;
        RECT 559.600 195.800 560.600 196.400 ;
        RECT 560.000 195.200 560.600 195.800 ;
        RECT 564.200 195.800 565.200 196.400 ;
        RECT 564.200 195.200 564.800 195.800 ;
        RECT 567.600 195.200 568.400 199.800 ;
        RECT 570.800 197.000 571.600 199.800 ;
        RECT 572.400 197.000 573.200 199.800 ;
        RECT 555.200 194.400 559.400 195.200 ;
        RECT 560.000 194.600 562.000 195.200 ;
        RECT 546.800 193.600 549.400 194.400 ;
        RECT 550.000 193.800 555.800 194.400 ;
        RECT 558.800 194.000 559.400 194.400 ;
        RECT 538.800 193.000 539.600 193.200 ;
        RECT 530.600 192.400 539.600 193.000 ;
        RECT 542.000 193.000 542.800 193.200 ;
        RECT 550.000 193.000 550.600 193.800 ;
        RECT 556.400 193.200 557.800 193.800 ;
        RECT 558.800 193.200 560.400 194.000 ;
        RECT 542.000 192.400 550.600 193.000 ;
        RECT 551.600 193.000 557.800 193.200 ;
        RECT 551.600 192.600 557.000 193.000 ;
        RECT 551.600 192.400 552.400 192.600 ;
        RECT 529.000 186.800 529.800 191.200 ;
        RECT 530.600 190.600 531.200 192.400 ;
        RECT 530.400 190.000 531.200 190.600 ;
        RECT 537.200 190.000 560.600 190.600 ;
        RECT 530.400 188.000 531.000 190.000 ;
        RECT 537.200 189.400 538.000 190.000 ;
        RECT 554.800 189.600 555.600 190.000 ;
        RECT 559.600 189.800 560.600 190.000 ;
        RECT 559.600 189.600 560.400 189.800 ;
        RECT 531.600 188.600 535.400 189.400 ;
        RECT 530.400 187.400 531.600 188.000 ;
        RECT 526.000 184.800 526.800 186.400 ;
        RECT 529.000 186.000 530.000 186.800 ;
        RECT 529.200 182.200 530.000 186.000 ;
        RECT 530.800 182.200 531.600 187.400 ;
        RECT 534.600 187.400 535.400 188.600 ;
        RECT 534.600 186.800 536.400 187.400 ;
        RECT 535.600 186.200 536.400 186.800 ;
        RECT 540.400 186.400 541.200 189.200 ;
        RECT 543.600 188.600 546.800 189.400 ;
        RECT 550.600 188.600 552.600 189.400 ;
        RECT 561.200 189.000 562.000 194.600 ;
        RECT 543.200 187.800 544.000 188.000 ;
        RECT 543.200 187.200 547.600 187.800 ;
        RECT 546.800 187.000 547.600 187.200 ;
        RECT 548.400 186.800 549.200 188.400 ;
        RECT 535.600 185.400 538.000 186.200 ;
        RECT 540.400 185.600 541.400 186.400 ;
        RECT 544.400 185.600 546.000 186.400 ;
        RECT 546.800 186.200 547.600 186.400 ;
        RECT 550.600 186.200 551.400 188.600 ;
        RECT 553.200 188.200 562.000 189.000 ;
        RECT 556.600 186.800 559.600 187.600 ;
        RECT 556.600 186.200 557.400 186.800 ;
        RECT 546.800 185.600 551.400 186.200 ;
        RECT 537.200 182.200 538.000 185.400 ;
        RECT 554.800 185.400 557.400 186.200 ;
        RECT 538.800 182.200 539.600 185.000 ;
        RECT 540.400 182.200 541.200 185.000 ;
        RECT 542.000 182.200 542.800 185.000 ;
        RECT 543.600 182.200 544.400 185.000 ;
        RECT 546.800 182.200 547.600 185.000 ;
        RECT 550.000 182.200 550.800 185.000 ;
        RECT 551.600 182.200 552.400 185.000 ;
        RECT 553.200 182.200 554.000 185.000 ;
        RECT 554.800 182.200 555.600 185.400 ;
        RECT 561.200 182.200 562.000 188.200 ;
        RECT 562.800 194.600 564.800 195.200 ;
        RECT 562.800 189.000 563.600 194.600 ;
        RECT 565.400 194.400 569.600 195.200 ;
        RECT 574.000 195.000 574.800 199.800 ;
        RECT 577.200 195.000 578.000 199.800 ;
        RECT 565.400 194.000 566.000 194.400 ;
        RECT 564.400 193.200 566.000 194.000 ;
        RECT 569.000 193.800 574.800 194.400 ;
        RECT 567.000 193.200 568.400 193.800 ;
        RECT 567.000 193.000 573.200 193.200 ;
        RECT 567.800 192.600 573.200 193.000 ;
        RECT 572.400 192.400 573.200 192.600 ;
        RECT 574.200 193.000 574.800 193.800 ;
        RECT 575.400 193.600 578.000 194.400 ;
        RECT 580.400 193.600 581.200 199.800 ;
        RECT 582.000 197.000 582.800 199.800 ;
        RECT 583.600 197.000 584.400 199.800 ;
        RECT 585.200 197.000 586.000 199.800 ;
        RECT 583.600 194.400 587.800 195.200 ;
        RECT 588.400 194.400 589.200 199.800 ;
        RECT 591.600 195.200 592.400 199.800 ;
        RECT 591.600 194.600 594.200 195.200 ;
        RECT 588.400 193.600 591.000 194.400 ;
        RECT 582.000 193.000 582.800 193.200 ;
        RECT 574.200 192.400 582.800 193.000 ;
        RECT 585.200 193.000 586.000 193.200 ;
        RECT 593.600 193.000 594.200 194.600 ;
        RECT 585.200 192.400 594.200 193.000 ;
        RECT 593.600 190.600 594.200 192.400 ;
        RECT 594.800 192.000 595.600 199.800 ;
        RECT 598.800 193.600 599.600 194.400 ;
        RECT 598.800 192.400 599.400 193.600 ;
        RECT 600.200 192.400 601.000 199.800 ;
        RECT 594.800 191.200 595.800 192.000 ;
        RECT 598.000 191.800 599.400 192.400 ;
        RECT 600.000 191.800 601.000 192.400 ;
        RECT 604.400 192.400 605.200 199.800 ;
        RECT 604.400 191.800 606.600 192.400 ;
        RECT 598.000 191.600 598.800 191.800 ;
        RECT 564.200 190.000 587.600 190.600 ;
        RECT 593.600 190.000 594.400 190.600 ;
        RECT 564.200 189.800 565.000 190.000 ;
        RECT 566.000 189.600 566.800 190.000 ;
        RECT 569.200 189.600 570.000 190.000 ;
        RECT 586.800 189.400 587.600 190.000 ;
        RECT 562.800 188.200 571.600 189.000 ;
        RECT 572.200 188.600 574.200 189.400 ;
        RECT 578.000 188.600 581.200 189.400 ;
        RECT 562.800 182.200 563.600 188.200 ;
        RECT 565.200 186.800 568.200 187.600 ;
        RECT 567.400 186.200 568.200 186.800 ;
        RECT 573.400 186.200 574.200 188.600 ;
        RECT 575.600 186.800 576.400 188.400 ;
        RECT 580.800 187.800 581.600 188.000 ;
        RECT 577.200 187.200 581.600 187.800 ;
        RECT 577.200 187.000 578.000 187.200 ;
        RECT 583.600 186.400 584.400 189.200 ;
        RECT 589.400 188.600 593.200 189.400 ;
        RECT 589.400 187.400 590.200 188.600 ;
        RECT 593.800 188.000 594.400 190.000 ;
        RECT 577.200 186.200 578.000 186.400 ;
        RECT 567.400 185.400 570.000 186.200 ;
        RECT 573.400 185.600 578.000 186.200 ;
        RECT 578.800 185.600 580.400 186.400 ;
        RECT 583.400 185.600 584.400 186.400 ;
        RECT 588.400 186.800 590.200 187.400 ;
        RECT 593.200 187.400 594.400 188.000 ;
        RECT 588.400 186.200 589.200 186.800 ;
        RECT 569.200 182.200 570.000 185.400 ;
        RECT 586.800 185.400 589.200 186.200 ;
        RECT 570.800 182.200 571.600 185.000 ;
        RECT 572.400 182.200 573.200 185.000 ;
        RECT 574.000 182.200 574.800 185.000 ;
        RECT 577.200 182.200 578.000 185.000 ;
        RECT 580.400 182.200 581.200 185.000 ;
        RECT 582.000 182.200 582.800 185.000 ;
        RECT 583.600 182.200 584.400 185.000 ;
        RECT 585.200 182.200 586.000 185.000 ;
        RECT 586.800 182.200 587.600 185.400 ;
        RECT 593.200 182.200 594.000 187.400 ;
        RECT 595.000 186.800 595.800 191.200 ;
        RECT 600.000 188.400 600.600 191.800 ;
        RECT 606.000 191.200 606.600 191.800 ;
        RECT 606.000 190.400 607.200 191.200 ;
        RECT 601.200 188.800 602.000 190.400 ;
        RECT 602.800 190.300 603.600 190.400 ;
        RECT 604.400 190.300 605.200 190.400 ;
        RECT 602.800 189.700 605.200 190.300 ;
        RECT 602.800 189.600 603.600 189.700 ;
        RECT 604.400 188.800 605.200 189.700 ;
        RECT 598.000 187.600 600.600 188.400 ;
        RECT 602.800 188.200 603.600 188.400 ;
        RECT 602.000 187.600 603.600 188.200 ;
        RECT 594.800 186.000 595.800 186.800 ;
        RECT 598.200 186.200 598.800 187.600 ;
        RECT 602.000 187.200 602.800 187.600 ;
        RECT 606.000 187.400 606.600 190.400 ;
        RECT 604.400 186.800 606.600 187.400 ;
        RECT 599.800 186.200 603.400 186.600 ;
        RECT 594.800 182.200 595.600 186.000 ;
        RECT 598.000 182.200 598.800 186.200 ;
        RECT 599.600 186.000 603.600 186.200 ;
        RECT 599.600 182.200 600.400 186.000 ;
        RECT 602.800 182.200 603.600 186.000 ;
        RECT 604.400 182.200 605.200 186.800 ;
        RECT 1.200 175.000 2.000 179.800 ;
        RECT 5.600 178.400 6.400 179.800 ;
        RECT 4.400 177.800 6.400 178.400 ;
        RECT 10.000 177.800 10.800 179.800 ;
        RECT 14.200 178.400 15.400 179.800 ;
        RECT 14.000 177.800 15.400 178.400 ;
        RECT 4.400 177.000 5.200 177.800 ;
        RECT 10.000 177.200 10.600 177.800 ;
        RECT 6.000 175.600 6.800 177.200 ;
        RECT 7.800 176.600 10.600 177.200 ;
        RECT 14.000 177.000 14.800 177.800 ;
        RECT 7.800 176.400 8.600 176.600 ;
        RECT 2.000 174.200 3.600 174.400 ;
        RECT 6.200 174.200 6.800 175.600 ;
        RECT 15.800 175.400 16.600 175.600 ;
        RECT 18.800 175.400 19.600 179.800 ;
        RECT 20.400 175.800 21.200 179.800 ;
        RECT 22.000 176.000 22.800 179.800 ;
        RECT 25.200 176.000 26.000 179.800 ;
        RECT 22.000 175.800 26.000 176.000 ;
        RECT 26.800 177.000 27.600 179.000 ;
        RECT 15.800 174.800 19.600 175.400 ;
        RECT 11.800 174.200 12.600 174.400 ;
        RECT 2.000 173.600 13.000 174.200 ;
        RECT 5.000 173.400 5.800 173.600 ;
        RECT 3.400 172.400 4.200 172.600 ;
        RECT 3.400 172.300 8.400 172.400 ;
        RECT 9.200 172.300 10.000 172.400 ;
        RECT 3.400 171.800 10.000 172.300 ;
        RECT 7.600 171.700 10.000 171.800 ;
        RECT 7.600 171.600 8.400 171.700 ;
        RECT 9.200 171.600 10.000 171.700 ;
        RECT 1.200 171.000 6.800 171.200 ;
        RECT 1.200 170.800 7.000 171.000 ;
        RECT 1.200 170.600 11.000 170.800 ;
        RECT 1.200 162.200 2.000 170.600 ;
        RECT 6.200 170.200 11.000 170.600 ;
        RECT 4.400 169.000 9.800 169.600 ;
        RECT 4.400 168.800 5.200 169.000 ;
        RECT 9.000 168.800 9.800 169.000 ;
        RECT 10.400 169.000 11.000 170.200 ;
        RECT 12.400 170.400 13.000 173.600 ;
        RECT 14.000 172.800 14.800 173.000 ;
        RECT 14.000 172.200 17.800 172.800 ;
        RECT 17.000 172.000 17.800 172.200 ;
        RECT 15.400 171.400 16.200 171.600 ;
        RECT 18.800 171.400 19.600 174.800 ;
        RECT 20.600 174.400 21.200 175.800 ;
        RECT 22.200 175.400 25.800 175.800 ;
        RECT 26.800 174.800 27.400 177.000 ;
        RECT 31.000 176.000 31.800 179.000 ;
        RECT 38.000 176.400 38.800 179.800 ;
        RECT 31.000 175.400 32.600 176.000 ;
        RECT 31.800 175.000 32.600 175.400 ;
        RECT 24.400 174.400 25.200 174.800 ;
        RECT 20.400 173.600 23.000 174.400 ;
        RECT 24.400 173.800 26.000 174.400 ;
        RECT 26.800 174.200 31.000 174.800 ;
        RECT 25.200 173.600 26.000 173.800 ;
        RECT 30.000 173.800 31.000 174.200 ;
        RECT 32.000 174.400 32.600 175.000 ;
        RECT 37.800 175.800 38.800 176.400 ;
        RECT 37.800 174.400 38.400 175.800 ;
        RECT 41.200 175.200 42.000 179.800 ;
        RECT 42.800 175.800 43.600 179.800 ;
        RECT 44.400 176.000 45.200 179.800 ;
        RECT 47.600 176.000 48.400 179.800 ;
        RECT 44.400 175.800 48.400 176.000 ;
        RECT 39.400 174.600 42.000 175.200 ;
        RECT 20.400 172.300 21.200 172.400 ;
        RECT 22.400 172.300 23.000 173.600 ;
        RECT 20.400 171.700 23.000 172.300 ;
        RECT 20.400 171.600 21.200 171.700 ;
        RECT 15.400 170.800 19.600 171.400 ;
        RECT 12.400 169.800 14.800 170.400 ;
        RECT 11.800 169.000 12.600 169.200 ;
        RECT 10.400 168.400 12.600 169.000 ;
        RECT 14.200 168.800 14.800 169.800 ;
        RECT 14.200 168.000 15.600 168.800 ;
        RECT 7.800 167.400 8.600 167.600 ;
        RECT 10.600 167.400 11.400 167.600 ;
        RECT 4.400 166.200 5.200 167.000 ;
        RECT 7.800 166.800 11.400 167.400 ;
        RECT 10.000 166.200 10.600 166.800 ;
        RECT 14.000 166.200 14.800 167.000 ;
        RECT 4.400 165.600 6.400 166.200 ;
        RECT 5.600 162.200 6.400 165.600 ;
        RECT 10.000 162.200 10.800 166.200 ;
        RECT 14.200 162.200 15.400 166.200 ;
        RECT 18.800 162.200 19.600 170.800 ;
        RECT 20.400 170.200 21.200 170.400 ;
        RECT 22.400 170.200 23.000 171.700 ;
        RECT 23.600 171.600 24.400 173.200 ;
        RECT 26.800 171.600 27.600 173.200 ;
        RECT 28.400 171.600 29.200 173.200 ;
        RECT 30.000 173.000 31.400 173.800 ;
        RECT 32.000 173.600 34.000 174.400 ;
        RECT 37.800 173.600 38.800 174.400 ;
        RECT 30.000 171.000 30.600 173.000 ;
        RECT 32.000 172.400 32.600 173.600 ;
        RECT 31.600 171.600 32.600 172.400 ;
        RECT 26.800 170.400 30.600 171.000 ;
        RECT 20.400 169.600 21.800 170.200 ;
        RECT 22.400 169.600 23.400 170.200 ;
        RECT 21.200 168.400 21.800 169.600 ;
        RECT 21.200 167.600 22.000 168.400 ;
        RECT 22.600 162.200 23.400 169.600 ;
        RECT 26.800 167.000 27.400 170.400 ;
        RECT 32.000 169.800 32.600 171.600 ;
        RECT 33.200 170.800 34.000 172.400 ;
        RECT 31.000 169.200 32.600 169.800 ;
        RECT 37.800 170.200 38.400 173.600 ;
        RECT 39.400 173.000 40.000 174.600 ;
        RECT 43.000 174.400 43.600 175.800 ;
        RECT 44.600 175.400 48.200 175.800 ;
        RECT 46.800 174.400 47.600 174.800 ;
        RECT 42.800 173.600 45.400 174.400 ;
        RECT 46.800 173.800 48.400 174.400 ;
        RECT 47.600 173.600 48.400 173.800 ;
        RECT 39.000 172.200 40.000 173.000 ;
        RECT 39.400 170.200 40.000 172.200 ;
        RECT 41.000 172.400 41.800 173.200 ;
        RECT 41.000 171.600 42.000 172.400 ;
        RECT 42.800 170.200 43.600 170.400 ;
        RECT 44.800 170.200 45.400 173.600 ;
        RECT 46.000 172.300 46.800 173.200 ;
        RECT 49.200 172.300 50.000 179.800 ;
        RECT 50.800 175.600 51.600 177.200 ;
        RECT 46.000 171.700 50.000 172.300 ;
        RECT 46.000 171.600 46.800 171.700 ;
        RECT 37.800 169.200 38.800 170.200 ;
        RECT 39.400 169.600 42.000 170.200 ;
        RECT 42.800 169.600 44.200 170.200 ;
        RECT 44.800 169.600 45.800 170.200 ;
        RECT 26.800 163.000 27.600 167.000 ;
        RECT 31.000 162.200 31.800 169.200 ;
        RECT 38.000 162.200 38.800 169.200 ;
        RECT 41.200 162.200 42.000 169.600 ;
        RECT 43.600 168.400 44.200 169.600 ;
        RECT 43.600 167.600 44.400 168.400 ;
        RECT 45.000 164.400 45.800 169.600 ;
        RECT 45.000 163.600 46.800 164.400 ;
        RECT 45.000 162.200 45.800 163.600 ;
        RECT 49.200 162.200 50.000 171.700 ;
        RECT 52.400 175.400 53.200 179.800 ;
        RECT 56.600 178.400 57.800 179.800 ;
        RECT 56.600 177.800 58.000 178.400 ;
        RECT 61.200 177.800 62.000 179.800 ;
        RECT 65.600 178.400 66.400 179.800 ;
        RECT 65.600 177.800 67.600 178.400 ;
        RECT 57.200 177.000 58.000 177.800 ;
        RECT 61.400 177.200 62.000 177.800 ;
        RECT 61.400 176.600 64.200 177.200 ;
        RECT 63.400 176.400 64.200 176.600 ;
        RECT 65.200 176.400 66.000 177.200 ;
        RECT 66.800 177.000 67.600 177.800 ;
        RECT 55.400 175.400 56.200 175.600 ;
        RECT 52.400 174.800 56.200 175.400 ;
        RECT 52.400 171.400 53.200 174.800 ;
        RECT 59.400 174.200 60.200 174.400 ;
        RECT 65.200 174.200 65.800 176.400 ;
        RECT 70.000 175.000 70.800 179.800 ;
        RECT 75.400 176.400 76.200 179.000 ;
        RECT 79.600 177.000 80.400 179.000 ;
        RECT 75.400 176.000 77.200 176.400 ;
        RECT 74.600 175.600 77.200 176.000 ;
        RECT 74.600 175.400 76.200 175.600 ;
        RECT 74.600 175.000 75.400 175.400 ;
        RECT 74.600 174.400 75.200 175.000 ;
        RECT 79.800 174.800 80.400 177.000 ;
        RECT 81.200 176.000 82.000 179.800 ;
        RECT 84.400 176.000 85.200 179.800 ;
        RECT 81.200 175.800 85.200 176.000 ;
        RECT 86.000 175.800 86.800 179.800 ;
        RECT 87.600 175.800 88.400 179.800 ;
        RECT 89.200 176.000 90.000 179.800 ;
        RECT 92.400 176.000 93.200 179.800 ;
        RECT 89.200 175.800 93.200 176.000 ;
        RECT 81.400 175.400 85.000 175.800 ;
        RECT 68.400 174.200 70.000 174.400 ;
        RECT 59.000 173.600 70.000 174.200 ;
        RECT 73.200 173.600 75.200 174.400 ;
        RECT 76.200 174.200 80.400 174.800 ;
        RECT 82.000 174.400 82.800 174.800 ;
        RECT 86.000 174.400 86.600 175.800 ;
        RECT 87.800 174.400 88.400 175.800 ;
        RECT 89.400 175.400 93.000 175.800 ;
        RECT 94.000 175.600 94.800 177.200 ;
        RECT 91.600 174.400 92.400 174.800 ;
        RECT 76.200 173.800 77.200 174.200 ;
        RECT 57.200 172.800 58.000 173.000 ;
        RECT 54.200 172.200 58.000 172.800 ;
        RECT 54.200 172.000 55.000 172.200 ;
        RECT 55.800 171.400 56.600 171.600 ;
        RECT 52.400 170.800 56.600 171.400 ;
        RECT 52.400 162.200 53.200 170.800 ;
        RECT 59.000 170.400 59.600 173.600 ;
        RECT 66.200 173.400 67.000 173.600 ;
        RECT 65.200 172.400 66.000 172.600 ;
        RECT 67.800 172.400 68.600 172.600 ;
        RECT 63.600 171.800 68.600 172.400 ;
        RECT 63.600 171.600 64.400 171.800 ;
        RECT 65.200 171.000 70.800 171.200 ;
        RECT 65.000 170.800 70.800 171.000 ;
        RECT 73.200 170.800 74.000 172.400 ;
        RECT 57.200 169.800 59.600 170.400 ;
        RECT 61.000 170.600 70.800 170.800 ;
        RECT 61.000 170.200 65.800 170.600 ;
        RECT 57.200 168.800 57.800 169.800 ;
        RECT 56.400 168.000 57.800 168.800 ;
        RECT 59.400 169.000 60.200 169.200 ;
        RECT 61.000 169.000 61.600 170.200 ;
        RECT 59.400 168.400 61.600 169.000 ;
        RECT 62.200 169.000 67.600 169.600 ;
        RECT 62.200 168.800 63.000 169.000 ;
        RECT 66.800 168.800 67.600 169.000 ;
        RECT 60.600 167.400 61.400 167.600 ;
        RECT 63.400 167.400 64.200 167.600 ;
        RECT 57.200 166.200 58.000 167.000 ;
        RECT 60.600 166.800 64.200 167.400 ;
        RECT 61.400 166.200 62.000 166.800 ;
        RECT 66.800 166.200 67.600 167.000 ;
        RECT 56.600 162.200 57.800 166.200 ;
        RECT 61.200 162.200 62.000 166.200 ;
        RECT 65.600 165.600 67.600 166.200 ;
        RECT 65.600 162.200 66.400 165.600 ;
        RECT 70.000 162.200 70.800 170.600 ;
        RECT 74.600 169.800 75.200 173.600 ;
        RECT 75.800 173.000 77.200 173.800 ;
        RECT 81.200 173.800 82.800 174.400 ;
        RECT 81.200 173.600 82.000 173.800 ;
        RECT 84.200 173.600 86.800 174.400 ;
        RECT 87.600 173.600 90.200 174.400 ;
        RECT 91.600 173.800 93.200 174.400 ;
        RECT 92.400 173.600 93.200 173.800 ;
        RECT 76.600 171.000 77.200 173.000 ;
        RECT 78.000 171.600 78.800 173.200 ;
        RECT 79.600 171.600 80.400 173.200 ;
        RECT 82.800 171.600 83.600 173.200 ;
        RECT 76.600 170.400 80.400 171.000 ;
        RECT 84.200 170.400 84.800 173.600 ;
        RECT 89.600 172.300 90.200 173.600 ;
        RECT 86.100 171.700 90.200 172.300 ;
        RECT 86.100 170.400 86.700 171.700 ;
        RECT 74.600 169.200 76.200 169.800 ;
        RECT 75.400 162.200 76.200 169.200 ;
        RECT 79.800 167.000 80.400 170.400 ;
        RECT 82.800 169.600 84.800 170.400 ;
        RECT 86.000 170.200 86.800 170.400 ;
        RECT 85.400 169.600 86.800 170.200 ;
        RECT 87.600 170.200 88.400 170.400 ;
        RECT 89.600 170.200 90.200 171.700 ;
        RECT 90.800 171.600 91.600 173.200 ;
        RECT 95.600 172.300 96.400 179.800 ;
        RECT 101.000 178.400 101.800 179.000 ;
        RECT 101.000 177.600 102.800 178.400 ;
        RECT 101.000 176.000 101.800 177.600 ;
        RECT 105.200 177.000 106.000 179.000 ;
        RECT 100.200 175.400 101.800 176.000 ;
        RECT 100.200 175.000 101.000 175.400 ;
        RECT 100.200 174.400 100.800 175.000 ;
        RECT 105.400 174.800 106.000 177.000 ;
        RECT 106.800 175.600 107.600 177.200 ;
        RECT 98.800 173.600 100.800 174.400 ;
        RECT 101.800 174.200 106.000 174.800 ;
        RECT 101.800 173.800 102.800 174.200 ;
        RECT 97.200 172.300 98.000 172.400 ;
        RECT 95.600 171.700 98.000 172.300 ;
        RECT 87.600 169.600 89.000 170.200 ;
        RECT 89.600 169.600 90.600 170.200 ;
        RECT 79.600 163.000 80.400 167.000 ;
        RECT 83.800 162.200 84.600 169.600 ;
        RECT 85.400 168.400 86.000 169.600 ;
        RECT 85.200 167.600 86.000 168.400 ;
        RECT 88.400 168.400 89.000 169.600 ;
        RECT 88.400 167.600 89.200 168.400 ;
        RECT 89.800 162.200 90.600 169.600 ;
        RECT 95.600 162.200 96.400 171.700 ;
        RECT 97.200 171.600 98.000 171.700 ;
        RECT 98.800 170.800 99.600 172.400 ;
        RECT 100.200 169.800 100.800 173.600 ;
        RECT 101.400 173.000 102.800 173.800 ;
        RECT 102.200 171.000 102.800 173.000 ;
        RECT 103.600 171.600 104.400 173.200 ;
        RECT 105.200 171.600 106.000 173.200 ;
        RECT 102.200 170.400 106.000 171.000 ;
        RECT 100.200 169.200 101.800 169.800 ;
        RECT 101.000 162.200 101.800 169.200 ;
        RECT 105.400 167.000 106.000 170.400 ;
        RECT 105.200 163.000 106.000 167.000 ;
        RECT 108.400 168.300 109.200 179.800 ;
        RECT 112.600 176.400 113.400 179.800 ;
        RECT 111.600 175.800 113.400 176.400 ;
        RECT 110.000 173.600 110.800 175.200 ;
        RECT 110.000 168.300 110.800 168.400 ;
        RECT 108.400 167.700 110.800 168.300 ;
        RECT 108.400 162.200 109.200 167.700 ;
        RECT 110.000 167.600 110.800 167.700 ;
        RECT 111.600 162.200 112.400 175.800 ;
        RECT 114.800 175.600 115.600 177.200 ;
        RECT 113.200 168.800 114.000 170.400 ;
        RECT 116.400 162.200 117.200 179.800 ;
        RECT 118.000 175.600 118.800 177.200 ;
        RECT 119.600 162.200 120.400 179.800 ;
        RECT 121.800 178.400 122.600 179.800 ;
        RECT 121.200 177.600 122.600 178.400 ;
        RECT 127.600 177.800 128.400 179.800 ;
        RECT 121.800 176.400 122.600 177.600 ;
        RECT 121.800 175.800 123.600 176.400 ;
        RECT 121.200 168.800 122.000 170.400 ;
        RECT 122.800 162.200 123.600 175.800 ;
        RECT 126.000 175.600 126.800 177.200 ;
        RECT 127.800 176.300 128.400 177.800 ;
        RECT 132.400 176.400 133.200 179.800 ;
        RECT 129.200 176.300 130.000 176.400 ;
        RECT 127.700 175.700 130.000 176.300 ;
        RECT 124.400 174.300 125.200 175.200 ;
        RECT 126.100 174.300 126.700 175.600 ;
        RECT 127.800 174.400 128.400 175.700 ;
        RECT 129.200 175.600 130.000 175.700 ;
        RECT 132.200 175.800 133.200 176.400 ;
        RECT 124.400 173.700 126.700 174.300 ;
        RECT 124.400 173.600 125.200 173.700 ;
        RECT 127.600 173.600 128.400 174.400 ;
        RECT 127.800 170.200 128.400 173.600 ;
        RECT 132.200 174.400 132.800 175.800 ;
        RECT 135.600 175.200 136.400 179.800 ;
        RECT 137.200 175.600 138.000 177.200 ;
        RECT 133.800 174.600 136.400 175.200 ;
        RECT 132.200 173.600 133.200 174.400 ;
        RECT 129.200 170.800 130.000 172.400 ;
        RECT 132.200 170.200 132.800 173.600 ;
        RECT 133.800 173.000 134.400 174.600 ;
        RECT 133.400 172.200 134.400 173.000 ;
        RECT 133.800 170.200 134.400 172.200 ;
        RECT 135.400 172.400 136.200 173.200 ;
        RECT 135.400 171.600 136.400 172.400 ;
        RECT 127.600 169.400 129.400 170.200 ;
        RECT 128.600 162.200 129.400 169.400 ;
        RECT 132.200 169.200 133.200 170.200 ;
        RECT 133.800 169.600 136.400 170.200 ;
        RECT 132.400 162.200 133.200 169.200 ;
        RECT 135.600 162.200 136.400 169.600 ;
        RECT 138.800 162.200 139.600 179.800 ;
        RECT 142.000 177.800 142.800 179.800 ;
        RECT 142.000 174.400 142.600 177.800 ;
        RECT 143.600 176.300 144.400 177.200 ;
        RECT 145.200 176.300 146.000 176.400 ;
        RECT 143.600 175.700 146.000 176.300 ;
        RECT 151.600 176.000 152.400 179.800 ;
        RECT 143.600 175.600 144.400 175.700 ;
        RECT 145.200 175.600 146.000 175.700 ;
        RECT 151.400 175.200 152.400 176.000 ;
        RECT 142.000 173.600 142.800 174.400 ;
        RECT 140.400 170.800 141.200 172.400 ;
        RECT 142.000 170.200 142.600 173.600 ;
        RECT 151.400 170.800 152.200 175.200 ;
        RECT 153.200 174.600 154.000 179.800 ;
        RECT 159.600 176.600 160.400 179.800 ;
        RECT 161.200 177.000 162.000 179.800 ;
        RECT 162.800 177.000 163.600 179.800 ;
        RECT 164.400 177.000 165.200 179.800 ;
        RECT 166.000 177.000 166.800 179.800 ;
        RECT 169.200 177.000 170.000 179.800 ;
        RECT 172.400 177.000 173.200 179.800 ;
        RECT 174.000 177.000 174.800 179.800 ;
        RECT 175.600 177.000 176.400 179.800 ;
        RECT 158.000 175.800 160.400 176.600 ;
        RECT 177.200 176.600 178.000 179.800 ;
        RECT 158.000 175.200 158.800 175.800 ;
        RECT 152.800 174.000 154.000 174.600 ;
        RECT 157.000 174.600 158.800 175.200 ;
        RECT 162.800 175.600 163.800 176.400 ;
        RECT 166.800 175.600 168.400 176.400 ;
        RECT 169.200 175.800 173.800 176.400 ;
        RECT 177.200 175.800 179.800 176.600 ;
        RECT 169.200 175.600 170.000 175.800 ;
        RECT 152.800 172.000 153.400 174.000 ;
        RECT 157.000 173.400 157.800 174.600 ;
        RECT 154.000 172.600 157.800 173.400 ;
        RECT 162.800 172.800 163.600 175.600 ;
        RECT 169.200 174.800 170.000 175.000 ;
        RECT 165.600 174.200 170.000 174.800 ;
        RECT 165.600 174.000 166.400 174.200 ;
        RECT 170.800 173.600 171.600 175.200 ;
        RECT 173.000 173.400 173.800 175.800 ;
        RECT 179.000 175.200 179.800 175.800 ;
        RECT 179.000 174.400 182.000 175.200 ;
        RECT 183.600 173.800 184.400 179.800 ;
        RECT 186.800 176.400 187.600 179.800 ;
        RECT 186.600 175.800 187.600 176.400 ;
        RECT 186.600 174.400 187.200 175.800 ;
        RECT 190.000 175.200 190.800 179.800 ;
        RECT 192.200 178.400 193.000 179.800 ;
        RECT 192.200 177.600 194.000 178.400 ;
        RECT 192.200 176.400 193.000 177.600 ;
        RECT 197.000 176.400 197.800 179.800 ;
        RECT 192.200 175.800 194.000 176.400 ;
        RECT 197.000 175.800 198.800 176.400 ;
        RECT 201.200 175.800 202.000 179.800 ;
        RECT 202.800 176.000 203.600 179.800 ;
        RECT 206.000 176.000 206.800 179.800 ;
        RECT 209.200 176.000 210.000 179.800 ;
        RECT 202.800 175.800 206.800 176.000 ;
        RECT 188.200 174.600 190.800 175.200 ;
        RECT 166.000 172.600 169.200 173.400 ;
        RECT 173.000 172.600 175.000 173.400 ;
        RECT 175.600 173.000 184.400 173.800 ;
        RECT 185.200 174.300 186.000 174.400 ;
        RECT 186.600 174.300 187.600 174.400 ;
        RECT 185.200 173.700 187.600 174.300 ;
        RECT 185.200 173.600 186.000 173.700 ;
        RECT 186.600 173.600 187.600 173.700 ;
        RECT 159.600 172.000 160.400 172.600 ;
        RECT 177.200 172.000 178.000 172.400 ;
        RECT 180.400 172.000 181.200 172.400 ;
        RECT 182.200 172.000 183.000 172.200 ;
        RECT 152.800 171.400 153.600 172.000 ;
        RECT 159.600 171.400 183.000 172.000 ;
        RECT 141.000 169.400 142.800 170.200 ;
        RECT 151.400 170.000 152.400 170.800 ;
        RECT 141.000 164.400 141.800 169.400 ;
        RECT 140.400 163.600 141.800 164.400 ;
        RECT 141.000 162.200 141.800 163.600 ;
        RECT 151.600 162.200 152.400 170.000 ;
        RECT 153.000 169.600 153.600 171.400 ;
        RECT 153.000 169.000 162.000 169.600 ;
        RECT 153.000 167.400 153.600 169.000 ;
        RECT 161.200 168.800 162.000 169.000 ;
        RECT 164.400 169.000 173.000 169.600 ;
        RECT 164.400 168.800 165.200 169.000 ;
        RECT 156.200 167.600 158.800 168.400 ;
        RECT 153.000 166.800 155.600 167.400 ;
        RECT 154.800 162.200 155.600 166.800 ;
        RECT 158.000 162.200 158.800 167.600 ;
        RECT 159.400 166.800 163.600 167.600 ;
        RECT 161.200 162.200 162.000 165.000 ;
        RECT 162.800 162.200 163.600 165.000 ;
        RECT 164.400 162.200 165.200 165.000 ;
        RECT 166.000 162.200 166.800 168.400 ;
        RECT 169.200 167.600 171.800 168.400 ;
        RECT 172.400 168.200 173.000 169.000 ;
        RECT 174.000 169.400 174.800 169.600 ;
        RECT 174.000 169.000 179.400 169.400 ;
        RECT 174.000 168.800 180.200 169.000 ;
        RECT 178.800 168.200 180.200 168.800 ;
        RECT 172.400 167.600 178.200 168.200 ;
        RECT 181.200 168.000 182.800 168.800 ;
        RECT 181.200 167.600 181.800 168.000 ;
        RECT 169.200 162.200 170.000 167.000 ;
        RECT 172.400 162.200 173.200 167.000 ;
        RECT 177.600 166.800 181.800 167.600 ;
        RECT 183.600 167.400 184.400 173.000 ;
        RECT 186.600 170.200 187.200 173.600 ;
        RECT 188.200 173.000 188.800 174.600 ;
        RECT 187.800 172.200 188.800 173.000 ;
        RECT 188.200 170.200 188.800 172.200 ;
        RECT 189.800 172.400 190.600 173.200 ;
        RECT 189.800 171.600 190.800 172.400 ;
        RECT 186.600 169.200 187.600 170.200 ;
        RECT 188.200 169.600 190.800 170.200 ;
        RECT 182.400 166.800 184.400 167.400 ;
        RECT 174.000 162.200 174.800 165.000 ;
        RECT 175.600 162.200 176.400 165.000 ;
        RECT 178.800 162.200 179.600 166.800 ;
        RECT 182.400 166.200 183.000 166.800 ;
        RECT 182.000 165.600 183.000 166.200 ;
        RECT 182.000 162.200 182.800 165.600 ;
        RECT 186.800 162.200 187.600 169.200 ;
        RECT 190.000 162.200 190.800 169.600 ;
        RECT 191.600 168.800 192.400 170.400 ;
        RECT 193.200 162.200 194.000 175.800 ;
        RECT 194.800 173.600 195.600 175.200 ;
        RECT 198.000 172.300 198.800 175.800 ;
        RECT 199.600 174.300 200.400 175.200 ;
        RECT 201.400 174.400 202.000 175.800 ;
        RECT 203.000 175.400 206.600 175.800 ;
        RECT 209.000 175.200 210.000 176.000 ;
        RECT 205.200 174.400 206.000 174.800 ;
        RECT 201.200 174.300 203.800 174.400 ;
        RECT 199.600 173.700 203.800 174.300 ;
        RECT 205.200 173.800 206.800 174.400 ;
        RECT 199.600 173.600 200.400 173.700 ;
        RECT 201.200 173.600 203.800 173.700 ;
        RECT 206.000 173.600 206.800 173.800 ;
        RECT 201.200 172.300 202.000 172.400 ;
        RECT 198.000 171.700 202.000 172.300 ;
        RECT 196.400 168.800 197.200 170.400 ;
        RECT 198.000 162.200 198.800 171.700 ;
        RECT 201.200 171.600 202.000 171.700 ;
        RECT 201.200 170.200 202.000 170.400 ;
        RECT 203.200 170.200 203.800 173.600 ;
        RECT 204.400 171.600 205.200 173.200 ;
        RECT 209.000 170.800 209.800 175.200 ;
        RECT 210.800 174.600 211.600 179.800 ;
        RECT 217.200 176.600 218.000 179.800 ;
        RECT 218.800 177.000 219.600 179.800 ;
        RECT 220.400 177.000 221.200 179.800 ;
        RECT 222.000 177.000 222.800 179.800 ;
        RECT 223.600 177.000 224.400 179.800 ;
        RECT 226.800 177.000 227.600 179.800 ;
        RECT 230.000 177.000 230.800 179.800 ;
        RECT 231.600 177.000 232.400 179.800 ;
        RECT 233.200 177.000 234.000 179.800 ;
        RECT 215.600 175.800 218.000 176.600 ;
        RECT 234.800 176.600 235.600 179.800 ;
        RECT 215.600 175.200 216.400 175.800 ;
        RECT 210.400 174.000 211.600 174.600 ;
        RECT 214.600 174.600 216.400 175.200 ;
        RECT 220.400 175.600 221.400 176.400 ;
        RECT 224.400 175.600 226.000 176.400 ;
        RECT 226.800 175.800 231.400 176.400 ;
        RECT 234.800 175.800 237.400 176.600 ;
        RECT 226.800 175.600 227.600 175.800 ;
        RECT 210.400 172.000 211.000 174.000 ;
        RECT 214.600 173.400 215.400 174.600 ;
        RECT 211.600 172.600 215.400 173.400 ;
        RECT 220.400 172.800 221.200 175.600 ;
        RECT 226.800 174.800 227.600 175.000 ;
        RECT 223.200 174.200 227.600 174.800 ;
        RECT 223.200 174.000 224.000 174.200 ;
        RECT 228.400 173.600 229.200 175.200 ;
        RECT 230.600 173.400 231.400 175.800 ;
        RECT 236.600 175.200 237.400 175.800 ;
        RECT 236.600 174.400 239.600 175.200 ;
        RECT 241.200 173.800 242.000 179.800 ;
        RECT 223.600 172.600 226.800 173.400 ;
        RECT 230.600 172.600 232.600 173.400 ;
        RECT 233.200 173.000 242.000 173.800 ;
        RECT 217.200 172.000 218.000 172.600 ;
        RECT 234.800 172.000 235.600 172.400 ;
        RECT 238.000 172.000 238.800 172.400 ;
        RECT 239.800 172.000 240.600 172.200 ;
        RECT 210.400 171.400 211.200 172.000 ;
        RECT 217.200 171.400 240.600 172.000 ;
        RECT 201.200 169.600 202.600 170.200 ;
        RECT 203.200 169.600 204.200 170.200 ;
        RECT 209.000 170.000 210.000 170.800 ;
        RECT 202.000 168.400 202.600 169.600 ;
        RECT 202.000 167.600 202.800 168.400 ;
        RECT 203.400 162.200 204.200 169.600 ;
        RECT 209.200 162.200 210.000 170.000 ;
        RECT 210.600 169.600 211.200 171.400 ;
        RECT 210.600 169.000 219.600 169.600 ;
        RECT 210.600 167.400 211.200 169.000 ;
        RECT 218.800 168.800 219.600 169.000 ;
        RECT 222.000 169.000 230.600 169.600 ;
        RECT 222.000 168.800 222.800 169.000 ;
        RECT 213.800 167.600 216.400 168.400 ;
        RECT 210.600 166.800 213.200 167.400 ;
        RECT 212.400 162.200 213.200 166.800 ;
        RECT 215.600 162.200 216.400 167.600 ;
        RECT 217.000 166.800 221.200 167.600 ;
        RECT 218.800 162.200 219.600 165.000 ;
        RECT 220.400 162.200 221.200 165.000 ;
        RECT 222.000 162.200 222.800 165.000 ;
        RECT 223.600 162.200 224.400 168.400 ;
        RECT 226.800 167.600 229.400 168.400 ;
        RECT 230.000 168.200 230.600 169.000 ;
        RECT 231.600 169.400 232.400 169.600 ;
        RECT 231.600 169.000 237.000 169.400 ;
        RECT 231.600 168.800 237.800 169.000 ;
        RECT 236.400 168.200 237.800 168.800 ;
        RECT 230.000 167.600 235.800 168.200 ;
        RECT 238.800 168.000 240.400 168.800 ;
        RECT 238.800 167.600 239.400 168.000 ;
        RECT 226.800 162.200 227.600 167.000 ;
        RECT 230.000 162.200 230.800 167.000 ;
        RECT 235.200 166.800 239.400 167.600 ;
        RECT 241.200 167.400 242.000 173.000 ;
        RECT 240.000 166.800 242.000 167.400 ;
        RECT 242.800 173.800 243.600 179.800 ;
        RECT 249.200 176.600 250.000 179.800 ;
        RECT 250.800 177.000 251.600 179.800 ;
        RECT 252.400 177.000 253.200 179.800 ;
        RECT 254.000 177.000 254.800 179.800 ;
        RECT 257.200 177.000 258.000 179.800 ;
        RECT 260.400 177.000 261.200 179.800 ;
        RECT 262.000 177.000 262.800 179.800 ;
        RECT 263.600 177.000 264.400 179.800 ;
        RECT 265.200 177.000 266.000 179.800 ;
        RECT 247.400 175.800 250.000 176.600 ;
        RECT 266.800 176.600 267.600 179.800 ;
        RECT 253.400 175.800 258.000 176.400 ;
        RECT 247.400 175.200 248.200 175.800 ;
        RECT 245.200 174.400 248.200 175.200 ;
        RECT 242.800 173.000 251.600 173.800 ;
        RECT 253.400 173.400 254.200 175.800 ;
        RECT 257.200 175.600 258.000 175.800 ;
        RECT 258.800 175.600 260.400 176.400 ;
        RECT 263.400 175.600 264.400 176.400 ;
        RECT 266.800 175.800 269.200 176.600 ;
        RECT 255.600 173.600 256.400 175.200 ;
        RECT 257.200 174.800 258.000 175.000 ;
        RECT 257.200 174.200 261.600 174.800 ;
        RECT 260.800 174.000 261.600 174.200 ;
        RECT 242.800 167.400 243.600 173.000 ;
        RECT 252.200 172.600 254.200 173.400 ;
        RECT 258.000 172.600 261.200 173.400 ;
        RECT 263.600 172.800 264.400 175.600 ;
        RECT 268.400 175.200 269.200 175.800 ;
        RECT 268.400 174.600 270.200 175.200 ;
        RECT 269.400 173.400 270.200 174.600 ;
        RECT 273.200 174.600 274.000 179.800 ;
        RECT 274.800 176.000 275.600 179.800 ;
        RECT 278.600 176.400 279.400 179.800 ;
        RECT 274.800 175.200 275.800 176.000 ;
        RECT 278.600 175.800 280.400 176.400 ;
        RECT 273.200 174.000 274.400 174.600 ;
        RECT 269.400 172.600 273.200 173.400 ;
        RECT 244.200 172.000 245.000 172.200 ;
        RECT 249.200 172.000 250.000 172.400 ;
        RECT 266.800 172.000 267.600 172.600 ;
        RECT 273.800 172.000 274.400 174.000 ;
        RECT 244.200 171.400 267.600 172.000 ;
        RECT 273.600 171.400 274.400 172.000 ;
        RECT 273.600 169.600 274.200 171.400 ;
        RECT 275.000 170.800 275.800 175.200 ;
        RECT 276.400 174.300 277.200 174.400 ;
        RECT 279.600 174.300 280.400 175.800 ;
        RECT 284.400 175.200 285.200 179.800 ;
        RECT 287.600 175.200 288.400 179.800 ;
        RECT 290.800 175.200 291.600 179.800 ;
        RECT 294.000 175.200 294.800 179.800 ;
        RECT 276.400 173.700 280.400 174.300 ;
        RECT 276.400 173.600 277.200 173.700 ;
        RECT 252.400 169.400 253.200 169.600 ;
        RECT 247.800 169.000 253.200 169.400 ;
        RECT 247.000 168.800 253.200 169.000 ;
        RECT 254.200 169.000 262.800 169.600 ;
        RECT 244.400 168.000 246.000 168.800 ;
        RECT 247.000 168.200 248.400 168.800 ;
        RECT 254.200 168.200 254.800 169.000 ;
        RECT 262.000 168.800 262.800 169.000 ;
        RECT 265.200 169.000 274.200 169.600 ;
        RECT 265.200 168.800 266.000 169.000 ;
        RECT 245.400 167.600 246.000 168.000 ;
        RECT 249.000 167.600 254.800 168.200 ;
        RECT 255.400 167.600 258.000 168.400 ;
        RECT 242.800 166.800 244.800 167.400 ;
        RECT 245.400 166.800 249.600 167.600 ;
        RECT 231.600 162.200 232.400 165.000 ;
        RECT 233.200 162.200 234.000 165.000 ;
        RECT 236.400 162.200 237.200 166.800 ;
        RECT 240.000 166.200 240.600 166.800 ;
        RECT 239.600 165.600 240.600 166.200 ;
        RECT 244.200 166.200 244.800 166.800 ;
        RECT 244.200 165.600 245.200 166.200 ;
        RECT 239.600 162.200 240.400 165.600 ;
        RECT 244.400 162.200 245.200 165.600 ;
        RECT 247.600 162.200 248.400 166.800 ;
        RECT 250.800 162.200 251.600 165.000 ;
        RECT 252.400 162.200 253.200 165.000 ;
        RECT 254.000 162.200 254.800 167.000 ;
        RECT 257.200 162.200 258.000 167.000 ;
        RECT 260.400 162.200 261.200 168.400 ;
        RECT 268.400 167.600 271.000 168.400 ;
        RECT 263.600 166.800 267.800 167.600 ;
        RECT 262.000 162.200 262.800 165.000 ;
        RECT 263.600 162.200 264.400 165.000 ;
        RECT 265.200 162.200 266.000 165.000 ;
        RECT 268.400 162.200 269.200 167.600 ;
        RECT 273.600 167.400 274.200 169.000 ;
        RECT 271.600 166.800 274.200 167.400 ;
        RECT 274.800 170.000 275.800 170.800 ;
        RECT 271.600 162.200 272.400 166.800 ;
        RECT 274.800 162.200 275.600 170.000 ;
        RECT 278.000 168.800 278.800 170.400 ;
        RECT 279.600 162.200 280.400 173.700 ;
        RECT 281.200 173.600 282.000 175.200 ;
        RECT 282.800 174.400 285.200 175.200 ;
        RECT 286.200 174.400 288.400 175.200 ;
        RECT 289.400 174.400 291.600 175.200 ;
        RECT 293.000 174.400 294.800 175.200 ;
        RECT 282.800 171.600 283.600 174.400 ;
        RECT 286.200 173.800 287.000 174.400 ;
        RECT 289.400 173.800 290.200 174.400 ;
        RECT 293.000 173.800 293.800 174.400 ;
        RECT 295.600 174.300 296.400 174.400 ;
        RECT 297.200 174.300 298.000 174.400 ;
        RECT 295.600 173.800 298.000 174.300 ;
        RECT 284.400 173.000 287.000 173.800 ;
        RECT 287.800 173.000 290.200 173.800 ;
        RECT 291.200 173.000 293.800 173.800 ;
        RECT 294.600 173.700 298.000 173.800 ;
        RECT 294.600 173.000 296.400 173.700 ;
        RECT 297.200 173.600 298.000 173.700 ;
        RECT 302.000 173.800 302.800 179.800 ;
        RECT 308.400 176.600 309.200 179.800 ;
        RECT 310.000 177.000 310.800 179.800 ;
        RECT 311.600 177.000 312.400 179.800 ;
        RECT 313.200 177.000 314.000 179.800 ;
        RECT 316.400 177.000 317.200 179.800 ;
        RECT 319.600 177.000 320.400 179.800 ;
        RECT 321.200 177.000 322.000 179.800 ;
        RECT 322.800 177.000 323.600 179.800 ;
        RECT 324.400 177.000 325.200 179.800 ;
        RECT 306.600 175.800 309.200 176.600 ;
        RECT 326.000 176.600 326.800 179.800 ;
        RECT 312.600 175.800 317.200 176.400 ;
        RECT 306.600 175.200 307.400 175.800 ;
        RECT 304.400 174.400 307.400 175.200 ;
        RECT 302.000 173.000 310.800 173.800 ;
        RECT 312.600 173.400 313.400 175.800 ;
        RECT 316.400 175.600 317.200 175.800 ;
        RECT 318.000 175.600 319.600 176.400 ;
        RECT 322.600 175.600 323.600 176.400 ;
        RECT 326.000 175.800 328.400 176.600 ;
        RECT 314.800 173.600 315.600 175.200 ;
        RECT 316.400 174.800 317.200 175.000 ;
        RECT 316.400 174.200 320.800 174.800 ;
        RECT 320.000 174.000 320.800 174.200 ;
        RECT 286.200 171.600 287.000 173.000 ;
        RECT 289.400 171.600 290.200 173.000 ;
        RECT 293.000 171.600 293.800 173.000 ;
        RECT 282.800 170.800 285.200 171.600 ;
        RECT 286.200 170.800 288.400 171.600 ;
        RECT 289.400 170.800 291.600 171.600 ;
        RECT 293.000 170.800 294.800 171.600 ;
        RECT 284.400 162.200 285.200 170.800 ;
        RECT 287.600 162.200 288.400 170.800 ;
        RECT 290.800 162.200 291.600 170.800 ;
        RECT 294.000 162.200 294.800 170.800 ;
        RECT 302.000 167.400 302.800 173.000 ;
        RECT 311.400 172.600 313.400 173.400 ;
        RECT 317.200 172.600 320.400 173.400 ;
        RECT 322.800 172.800 323.600 175.600 ;
        RECT 327.600 175.200 328.400 175.800 ;
        RECT 327.600 174.600 329.400 175.200 ;
        RECT 328.600 173.400 329.400 174.600 ;
        RECT 332.400 174.600 333.200 179.800 ;
        RECT 334.000 176.000 334.800 179.800 ;
        RECT 339.800 178.400 340.600 179.800 ;
        RECT 339.800 177.600 341.200 178.400 ;
        RECT 339.800 176.400 340.600 177.600 ;
        RECT 334.000 175.200 335.000 176.000 ;
        RECT 338.800 175.800 340.600 176.400 ;
        RECT 342.000 175.800 342.800 179.800 ;
        RECT 343.600 176.000 344.400 179.800 ;
        RECT 346.800 176.000 347.600 179.800 ;
        RECT 351.000 176.400 351.800 179.800 ;
        RECT 343.600 175.800 347.600 176.000 ;
        RECT 350.000 175.800 351.800 176.400 ;
        RECT 332.400 174.000 333.600 174.600 ;
        RECT 328.600 172.600 332.400 173.400 ;
        RECT 303.400 172.000 304.200 172.200 ;
        RECT 308.400 172.000 309.200 172.400 ;
        RECT 326.000 172.000 326.800 172.600 ;
        RECT 333.000 172.000 333.600 174.000 ;
        RECT 303.400 171.400 326.800 172.000 ;
        RECT 332.800 171.400 333.600 172.000 ;
        RECT 332.800 169.600 333.400 171.400 ;
        RECT 334.200 170.800 335.000 175.200 ;
        RECT 337.200 173.600 338.000 175.200 ;
        RECT 311.600 169.400 312.400 169.600 ;
        RECT 307.000 169.000 312.400 169.400 ;
        RECT 306.200 168.800 312.400 169.000 ;
        RECT 313.400 169.000 322.000 169.600 ;
        RECT 303.600 168.000 305.200 168.800 ;
        RECT 306.200 168.200 307.600 168.800 ;
        RECT 313.400 168.200 314.000 169.000 ;
        RECT 321.200 168.800 322.000 169.000 ;
        RECT 324.400 169.000 333.400 169.600 ;
        RECT 324.400 168.800 325.200 169.000 ;
        RECT 304.600 167.600 305.200 168.000 ;
        RECT 308.200 167.600 314.000 168.200 ;
        RECT 314.600 167.600 317.200 168.400 ;
        RECT 302.000 166.800 304.000 167.400 ;
        RECT 304.600 166.800 308.800 167.600 ;
        RECT 303.400 166.200 304.000 166.800 ;
        RECT 303.400 165.600 304.400 166.200 ;
        RECT 303.600 162.200 304.400 165.600 ;
        RECT 306.800 162.200 307.600 166.800 ;
        RECT 310.000 162.200 310.800 165.000 ;
        RECT 311.600 162.200 312.400 165.000 ;
        RECT 313.200 162.200 314.000 167.000 ;
        RECT 316.400 162.200 317.200 167.000 ;
        RECT 319.600 162.200 320.400 168.400 ;
        RECT 327.600 167.600 330.200 168.400 ;
        RECT 322.800 166.800 327.000 167.600 ;
        RECT 321.200 162.200 322.000 165.000 ;
        RECT 322.800 162.200 323.600 165.000 ;
        RECT 324.400 162.200 325.200 165.000 ;
        RECT 327.600 162.200 328.400 167.600 ;
        RECT 332.800 167.400 333.400 169.000 ;
        RECT 330.800 166.800 333.400 167.400 ;
        RECT 334.000 170.000 335.000 170.800 ;
        RECT 330.800 162.200 331.600 166.800 ;
        RECT 334.000 162.200 334.800 170.000 ;
        RECT 338.800 162.200 339.600 175.800 ;
        RECT 342.200 174.400 342.800 175.800 ;
        RECT 343.800 175.400 347.400 175.800 ;
        RECT 346.000 174.400 346.800 174.800 ;
        RECT 342.000 173.600 344.600 174.400 ;
        RECT 346.000 173.800 347.600 174.400 ;
        RECT 346.800 173.600 347.600 173.800 ;
        RECT 348.400 173.600 349.200 175.200 ;
        RECT 340.400 168.800 341.200 170.400 ;
        RECT 342.000 170.200 342.800 170.400 ;
        RECT 344.000 170.200 344.600 173.600 ;
        RECT 345.200 171.600 346.000 173.200 ;
        RECT 342.000 169.600 343.400 170.200 ;
        RECT 344.000 169.600 345.000 170.200 ;
        RECT 342.800 168.400 343.400 169.600 ;
        RECT 342.800 167.600 343.600 168.400 ;
        RECT 344.200 162.200 345.000 169.600 ;
        RECT 350.000 162.200 350.800 175.800 ;
        RECT 353.200 175.200 354.000 179.800 ;
        RECT 356.400 176.400 357.200 179.800 ;
        RECT 362.200 178.400 363.000 179.800 ;
        RECT 362.200 177.600 363.600 178.400 ;
        RECT 362.200 176.400 363.000 177.600 ;
        RECT 356.400 175.800 357.400 176.400 ;
        RECT 353.200 174.600 355.800 175.200 ;
        RECT 353.400 172.400 354.200 173.200 ;
        RECT 353.200 171.600 354.200 172.400 ;
        RECT 355.200 173.000 355.800 174.600 ;
        RECT 356.800 174.400 357.400 175.800 ;
        RECT 361.200 175.800 363.000 176.400 ;
        RECT 364.400 176.000 365.200 179.800 ;
        RECT 367.600 176.000 368.400 179.800 ;
        RECT 364.400 175.800 368.400 176.000 ;
        RECT 369.200 175.800 370.000 179.800 ;
        RECT 356.400 173.600 357.400 174.400 ;
        RECT 358.000 174.300 358.800 174.400 ;
        RECT 359.600 174.300 360.400 175.200 ;
        RECT 358.000 173.700 360.400 174.300 ;
        RECT 358.000 173.600 358.800 173.700 ;
        RECT 359.600 173.600 360.400 173.700 ;
        RECT 355.200 172.200 356.200 173.000 ;
        RECT 351.600 168.800 352.400 170.400 ;
        RECT 355.200 170.200 355.800 172.200 ;
        RECT 356.800 170.200 357.400 173.600 ;
        RECT 353.200 169.600 355.800 170.200 ;
        RECT 353.200 162.200 354.000 169.600 ;
        RECT 356.400 169.200 357.400 170.200 ;
        RECT 356.400 162.200 357.200 169.200 ;
        RECT 361.200 162.200 362.000 175.800 ;
        RECT 364.600 175.400 368.200 175.800 ;
        RECT 365.200 174.400 366.000 174.800 ;
        RECT 369.200 174.400 369.800 175.800 ;
        RECT 370.800 175.200 371.600 179.800 ;
        RECT 374.000 176.400 374.800 179.800 ;
        RECT 379.800 178.400 380.600 179.800 ;
        RECT 379.800 177.600 381.200 178.400 ;
        RECT 379.800 176.400 380.600 177.600 ;
        RECT 374.000 175.800 375.000 176.400 ;
        RECT 370.800 174.600 373.400 175.200 ;
        RECT 364.400 173.800 366.000 174.400 ;
        RECT 364.400 173.600 365.200 173.800 ;
        RECT 367.400 173.600 370.000 174.400 ;
        RECT 366.000 172.300 366.800 173.200 ;
        RECT 364.500 171.700 366.800 172.300 ;
        RECT 366.000 171.600 366.800 171.700 ;
        RECT 362.800 168.800 363.600 170.400 ;
        RECT 367.400 170.200 368.000 173.600 ;
        RECT 371.000 172.400 371.800 173.200 ;
        RECT 370.800 171.600 371.800 172.400 ;
        RECT 372.800 173.000 373.400 174.600 ;
        RECT 374.400 174.400 375.000 175.800 ;
        RECT 378.800 175.800 380.600 176.400 ;
        RECT 374.000 173.600 375.000 174.400 ;
        RECT 377.200 173.600 378.000 175.200 ;
        RECT 372.800 172.200 373.800 173.000 ;
        RECT 369.200 170.200 370.000 170.400 ;
        RECT 372.800 170.200 373.400 172.200 ;
        RECT 374.400 170.200 375.000 173.600 ;
        RECT 367.000 169.600 368.000 170.200 ;
        RECT 368.600 169.600 370.000 170.200 ;
        RECT 370.800 169.600 373.400 170.200 ;
        RECT 367.000 162.200 367.800 169.600 ;
        RECT 368.600 168.400 369.200 169.600 ;
        RECT 368.400 167.600 369.200 168.400 ;
        RECT 370.800 162.200 371.600 169.600 ;
        RECT 374.000 169.200 375.000 170.200 ;
        RECT 374.000 162.200 374.800 169.200 ;
        RECT 378.800 162.200 379.600 175.800 ;
        RECT 380.400 168.800 381.200 170.400 ;
        RECT 382.000 168.300 382.800 179.800 ;
        RECT 383.600 176.300 384.400 177.200 ;
        RECT 385.200 176.300 386.000 179.800 ;
        RECT 389.400 178.400 390.600 179.800 ;
        RECT 389.400 177.800 390.800 178.400 ;
        RECT 394.000 177.800 394.800 179.800 ;
        RECT 398.400 178.400 399.200 179.800 ;
        RECT 398.400 177.800 400.400 178.400 ;
        RECT 390.000 177.000 390.800 177.800 ;
        RECT 394.200 177.200 394.800 177.800 ;
        RECT 394.200 176.600 397.000 177.200 ;
        RECT 396.200 176.400 397.000 176.600 ;
        RECT 398.000 176.400 398.800 177.200 ;
        RECT 399.600 177.000 400.400 177.800 ;
        RECT 383.600 175.700 386.000 176.300 ;
        RECT 383.600 175.600 384.400 175.700 ;
        RECT 385.200 175.400 386.000 175.700 ;
        RECT 388.200 175.400 389.000 175.600 ;
        RECT 385.200 174.800 389.000 175.400 ;
        RECT 385.200 171.400 386.000 174.800 ;
        RECT 392.200 174.200 393.000 174.400 ;
        RECT 398.000 174.200 398.600 176.400 ;
        RECT 402.800 175.000 403.600 179.800 ;
        RECT 404.400 176.000 405.200 179.800 ;
        RECT 407.600 176.000 408.400 179.800 ;
        RECT 404.400 175.800 408.400 176.000 ;
        RECT 409.200 175.800 410.000 179.800 ;
        RECT 404.600 175.400 408.200 175.800 ;
        RECT 405.200 174.400 406.000 174.800 ;
        RECT 409.200 174.400 409.800 175.800 ;
        RECT 410.800 175.600 411.600 179.800 ;
        RECT 412.400 176.000 413.200 179.800 ;
        RECT 415.600 176.000 416.400 179.800 ;
        RECT 421.000 176.000 421.800 179.000 ;
        RECT 425.200 177.000 426.000 179.000 ;
        RECT 412.400 175.800 416.400 176.000 ;
        RECT 411.000 174.400 411.600 175.600 ;
        RECT 412.600 175.400 416.200 175.800 ;
        RECT 420.200 175.400 421.800 176.000 ;
        RECT 420.200 175.000 421.000 175.400 ;
        RECT 414.800 174.400 415.600 174.800 ;
        RECT 420.200 174.400 420.800 175.000 ;
        RECT 425.400 174.800 426.000 177.000 ;
        RECT 426.800 175.000 427.600 179.800 ;
        RECT 431.200 178.400 432.000 179.800 ;
        RECT 430.000 177.800 432.000 178.400 ;
        RECT 435.600 177.800 436.400 179.800 ;
        RECT 439.800 178.400 441.000 179.800 ;
        RECT 439.600 177.800 441.000 178.400 ;
        RECT 430.000 177.000 430.800 177.800 ;
        RECT 435.600 177.200 436.200 177.800 ;
        RECT 431.600 176.400 432.400 177.200 ;
        RECT 433.400 176.600 436.200 177.200 ;
        RECT 439.600 177.000 440.400 177.800 ;
        RECT 433.400 176.400 434.200 176.600 ;
        RECT 401.200 174.200 402.800 174.400 ;
        RECT 391.800 173.600 402.800 174.200 ;
        RECT 404.400 173.800 406.000 174.400 ;
        RECT 404.400 173.600 405.200 173.800 ;
        RECT 407.400 173.600 410.000 174.400 ;
        RECT 410.800 173.600 413.400 174.400 ;
        RECT 414.800 173.800 416.400 174.400 ;
        RECT 415.600 173.600 416.400 173.800 ;
        RECT 417.200 174.300 418.000 174.400 ;
        RECT 418.800 174.300 420.800 174.400 ;
        RECT 417.200 173.700 420.800 174.300 ;
        RECT 421.800 174.200 426.000 174.800 ;
        RECT 427.600 174.200 429.200 174.400 ;
        RECT 431.800 174.200 432.400 176.400 ;
        RECT 441.400 175.400 442.200 175.600 ;
        RECT 444.400 175.400 445.200 179.800 ;
        RECT 446.000 176.000 446.800 179.800 ;
        RECT 449.200 176.000 450.000 179.800 ;
        RECT 446.000 175.800 450.000 176.000 ;
        RECT 450.800 175.800 451.600 179.800 ;
        RECT 452.400 175.800 453.200 179.800 ;
        RECT 454.000 176.000 454.800 179.800 ;
        RECT 457.200 176.000 458.000 179.800 ;
        RECT 454.000 175.800 458.000 176.000 ;
        RECT 463.600 176.000 464.400 179.800 ;
        RECT 466.800 176.000 467.600 179.800 ;
        RECT 463.600 175.800 467.600 176.000 ;
        RECT 468.400 175.800 469.200 179.800 ;
        RECT 470.000 176.000 470.800 179.800 ;
        RECT 473.200 176.000 474.000 179.800 ;
        RECT 470.000 175.800 474.000 176.000 ;
        RECT 474.800 175.800 475.600 179.800 ;
        RECT 480.200 176.000 481.000 179.000 ;
        RECT 484.400 177.000 485.200 179.000 ;
        RECT 446.200 175.400 449.800 175.800 ;
        RECT 441.400 174.800 445.200 175.400 ;
        RECT 433.200 174.200 434.000 174.400 ;
        RECT 437.400 174.200 438.200 174.400 ;
        RECT 421.800 173.800 422.800 174.200 ;
        RECT 417.200 173.600 418.000 173.700 ;
        RECT 418.800 173.600 420.800 173.700 ;
        RECT 390.000 172.800 390.800 173.000 ;
        RECT 387.000 172.200 390.800 172.800 ;
        RECT 387.000 172.000 387.800 172.200 ;
        RECT 388.600 171.400 389.400 171.600 ;
        RECT 385.200 170.800 389.400 171.400 ;
        RECT 383.600 168.300 384.400 168.400 ;
        RECT 382.000 167.700 384.400 168.300 ;
        RECT 382.000 162.200 382.800 167.700 ;
        RECT 383.600 167.600 384.400 167.700 ;
        RECT 385.200 162.200 386.000 170.800 ;
        RECT 391.800 170.400 392.400 173.600 ;
        RECT 399.000 173.400 399.800 173.600 ;
        RECT 398.000 172.400 398.800 172.600 ;
        RECT 400.600 172.400 401.400 172.600 ;
        RECT 396.400 171.800 401.400 172.400 ;
        RECT 396.400 171.600 397.200 171.800 ;
        RECT 406.000 171.600 406.800 173.200 ;
        RECT 407.400 172.300 408.000 173.600 ;
        RECT 407.400 171.700 411.500 172.300 ;
        RECT 398.000 171.000 403.600 171.200 ;
        RECT 397.800 170.800 403.600 171.000 ;
        RECT 390.000 169.800 392.400 170.400 ;
        RECT 393.800 170.600 403.600 170.800 ;
        RECT 393.800 170.200 398.600 170.600 ;
        RECT 390.000 168.800 390.600 169.800 ;
        RECT 389.200 168.000 390.600 168.800 ;
        RECT 392.200 169.000 393.000 169.200 ;
        RECT 393.800 169.000 394.400 170.200 ;
        RECT 392.200 168.400 394.400 169.000 ;
        RECT 395.000 169.000 400.400 169.600 ;
        RECT 395.000 168.800 395.800 169.000 ;
        RECT 399.600 168.800 400.400 169.000 ;
        RECT 393.400 167.400 394.200 167.600 ;
        RECT 396.200 167.400 397.000 167.600 ;
        RECT 390.000 166.200 390.800 167.000 ;
        RECT 393.400 166.800 397.000 167.400 ;
        RECT 394.200 166.200 394.800 166.800 ;
        RECT 399.600 166.200 400.400 167.000 ;
        RECT 389.400 162.200 390.600 166.200 ;
        RECT 394.000 162.200 394.800 166.200 ;
        RECT 398.400 165.600 400.400 166.200 ;
        RECT 398.400 162.200 399.200 165.600 ;
        RECT 402.800 162.200 403.600 170.600 ;
        RECT 407.400 170.200 408.000 171.700 ;
        RECT 410.900 170.400 411.500 171.700 ;
        RECT 409.200 170.200 410.000 170.400 ;
        RECT 407.000 169.600 408.000 170.200 ;
        RECT 408.600 169.600 410.000 170.200 ;
        RECT 410.800 170.200 411.600 170.400 ;
        RECT 412.800 170.200 413.400 173.600 ;
        RECT 414.000 171.600 414.800 173.200 ;
        RECT 417.200 172.300 418.000 172.400 ;
        RECT 418.800 172.300 419.600 172.400 ;
        RECT 417.200 171.700 419.600 172.300 ;
        RECT 417.200 171.600 418.000 171.700 ;
        RECT 418.800 170.800 419.600 171.700 ;
        RECT 410.800 169.600 412.200 170.200 ;
        RECT 412.800 169.600 413.800 170.200 ;
        RECT 407.000 162.200 407.800 169.600 ;
        RECT 408.600 168.400 409.200 169.600 ;
        RECT 408.400 167.600 409.200 168.400 ;
        RECT 411.600 168.400 412.200 169.600 ;
        RECT 411.600 167.600 412.400 168.400 ;
        RECT 413.000 162.200 413.800 169.600 ;
        RECT 420.200 169.800 420.800 173.600 ;
        RECT 421.400 173.000 422.800 173.800 ;
        RECT 427.600 173.600 438.600 174.200 ;
        RECT 430.600 173.400 431.400 173.600 ;
        RECT 422.200 171.000 422.800 173.000 ;
        RECT 423.600 171.600 424.400 173.200 ;
        RECT 425.200 171.600 426.000 173.200 ;
        RECT 429.000 172.400 429.800 172.600 ;
        RECT 429.000 171.800 434.000 172.400 ;
        RECT 433.200 171.600 434.000 171.800 ;
        RECT 426.800 171.000 432.400 171.200 ;
        RECT 422.200 170.400 426.000 171.000 ;
        RECT 420.200 169.200 421.800 169.800 ;
        RECT 421.000 162.200 421.800 169.200 ;
        RECT 425.400 167.000 426.000 170.400 ;
        RECT 425.200 163.000 426.000 167.000 ;
        RECT 426.800 170.800 432.600 171.000 ;
        RECT 426.800 170.600 436.600 170.800 ;
        RECT 426.800 162.200 427.600 170.600 ;
        RECT 431.800 170.200 436.600 170.600 ;
        RECT 430.000 169.000 435.400 169.600 ;
        RECT 430.000 168.800 430.800 169.000 ;
        RECT 434.600 168.800 435.400 169.000 ;
        RECT 436.000 169.000 436.600 170.200 ;
        RECT 438.000 170.400 438.600 173.600 ;
        RECT 439.600 172.800 440.400 173.000 ;
        RECT 439.600 172.200 443.400 172.800 ;
        RECT 442.600 172.000 443.400 172.200 ;
        RECT 441.000 171.400 441.800 171.600 ;
        RECT 444.400 171.400 445.200 174.800 ;
        RECT 446.800 174.400 447.600 174.800 ;
        RECT 450.800 174.400 451.400 175.800 ;
        RECT 452.600 174.400 453.200 175.800 ;
        RECT 454.200 175.400 457.800 175.800 ;
        RECT 463.800 175.400 467.400 175.800 ;
        RECT 456.400 174.400 457.200 174.800 ;
        RECT 464.400 174.400 465.200 174.800 ;
        RECT 468.400 174.400 469.000 175.800 ;
        RECT 470.200 175.400 473.800 175.800 ;
        RECT 470.800 174.400 471.600 174.800 ;
        RECT 474.800 174.400 475.400 175.800 ;
        RECT 479.400 175.400 481.000 176.000 ;
        RECT 479.400 175.000 480.200 175.400 ;
        RECT 479.400 174.400 480.000 175.000 ;
        RECT 484.600 174.800 485.200 177.000 ;
        RECT 446.000 173.800 447.600 174.400 ;
        RECT 446.000 173.600 446.800 173.800 ;
        RECT 449.000 173.600 451.600 174.400 ;
        RECT 452.400 173.600 455.000 174.400 ;
        RECT 456.400 174.300 458.000 174.400 ;
        RECT 463.600 174.300 465.200 174.400 ;
        RECT 456.400 173.800 465.200 174.300 ;
        RECT 457.200 173.700 464.400 173.800 ;
        RECT 457.200 173.600 458.000 173.700 ;
        RECT 463.600 173.600 464.400 173.700 ;
        RECT 466.600 173.600 469.200 174.400 ;
        RECT 470.000 173.800 471.600 174.400 ;
        RECT 473.000 174.300 475.600 174.400 ;
        RECT 476.400 174.300 477.200 174.400 ;
        RECT 470.000 173.600 470.800 173.800 ;
        RECT 473.000 173.700 477.200 174.300 ;
        RECT 473.000 173.600 475.600 173.700 ;
        RECT 476.400 173.600 477.200 173.700 ;
        RECT 478.000 173.600 480.000 174.400 ;
        RECT 481.000 174.200 485.200 174.800 ;
        RECT 486.000 175.400 486.800 179.800 ;
        RECT 490.200 178.400 491.400 179.800 ;
        RECT 490.200 177.800 491.600 178.400 ;
        RECT 494.800 177.800 495.600 179.800 ;
        RECT 499.200 178.400 500.000 179.800 ;
        RECT 499.200 177.800 501.200 178.400 ;
        RECT 490.800 177.000 491.600 177.800 ;
        RECT 495.000 177.200 495.600 177.800 ;
        RECT 495.000 176.600 497.800 177.200 ;
        RECT 497.000 176.400 497.800 176.600 ;
        RECT 498.800 176.400 499.600 177.200 ;
        RECT 500.400 177.000 501.200 177.800 ;
        RECT 489.000 175.400 489.800 175.600 ;
        RECT 486.000 174.800 489.800 175.400 ;
        RECT 481.000 173.800 482.000 174.200 ;
        RECT 447.600 171.600 448.400 173.200 ;
        RECT 449.000 172.400 449.600 173.600 ;
        RECT 449.000 171.600 450.000 172.400 ;
        RECT 454.400 172.300 455.000 173.600 ;
        RECT 450.900 171.700 455.000 172.300 ;
        RECT 441.000 170.800 445.200 171.400 ;
        RECT 438.000 169.800 440.400 170.400 ;
        RECT 437.400 169.000 438.200 169.200 ;
        RECT 436.000 168.400 438.200 169.000 ;
        RECT 439.800 168.800 440.400 169.800 ;
        RECT 439.800 168.000 441.200 168.800 ;
        RECT 433.400 167.400 434.200 167.600 ;
        RECT 436.200 167.400 437.000 167.600 ;
        RECT 430.000 166.200 430.800 167.000 ;
        RECT 433.400 166.800 437.000 167.400 ;
        RECT 435.600 166.200 436.200 166.800 ;
        RECT 439.600 166.200 440.400 167.000 ;
        RECT 430.000 165.600 432.000 166.200 ;
        RECT 431.200 162.200 432.000 165.600 ;
        RECT 435.600 162.200 436.400 166.200 ;
        RECT 439.800 162.200 441.000 166.200 ;
        RECT 444.400 162.200 445.200 170.800 ;
        RECT 449.000 170.200 449.600 171.600 ;
        RECT 450.900 170.400 451.500 171.700 ;
        RECT 450.800 170.200 451.600 170.400 ;
        RECT 448.600 169.600 449.600 170.200 ;
        RECT 450.200 169.600 451.600 170.200 ;
        RECT 452.400 170.200 453.200 170.400 ;
        RECT 454.400 170.200 455.000 171.700 ;
        RECT 455.600 172.300 456.400 173.200 ;
        RECT 463.600 172.300 464.400 172.400 ;
        RECT 465.200 172.300 466.000 173.200 ;
        RECT 455.600 171.700 466.000 172.300 ;
        RECT 455.600 171.600 456.400 171.700 ;
        RECT 463.600 171.600 464.400 171.700 ;
        RECT 465.200 171.600 466.000 171.700 ;
        RECT 466.600 170.400 467.200 173.600 ;
        RECT 471.600 171.600 472.400 173.200 ;
        RECT 452.400 169.600 453.800 170.200 ;
        RECT 454.400 169.600 455.400 170.200 ;
        RECT 465.200 169.600 467.200 170.400 ;
        RECT 468.400 170.200 469.200 170.400 ;
        RECT 473.000 170.200 473.600 173.600 ;
        RECT 474.800 172.300 475.600 172.400 ;
        RECT 478.000 172.300 478.800 172.400 ;
        RECT 474.800 171.700 478.800 172.300 ;
        RECT 474.800 171.600 475.600 171.700 ;
        RECT 478.000 170.800 478.800 171.700 ;
        RECT 474.800 170.200 475.600 170.400 ;
        RECT 467.800 169.600 469.200 170.200 ;
        RECT 472.600 169.600 473.600 170.200 ;
        RECT 474.200 169.600 475.600 170.200 ;
        RECT 479.400 169.800 480.000 173.600 ;
        RECT 480.600 173.000 482.000 173.800 ;
        RECT 481.400 171.000 482.000 173.000 ;
        RECT 482.800 171.600 483.600 173.200 ;
        RECT 484.400 171.600 485.200 173.200 ;
        RECT 486.000 171.400 486.800 174.800 ;
        RECT 493.000 174.200 493.800 174.400 ;
        RECT 498.800 174.200 499.400 176.400 ;
        RECT 503.600 175.000 504.400 179.800 ;
        RECT 505.200 176.000 506.000 179.800 ;
        RECT 508.400 176.000 509.200 179.800 ;
        RECT 505.200 175.800 509.200 176.000 ;
        RECT 510.000 175.800 510.800 179.800 ;
        RECT 511.600 175.800 512.400 179.800 ;
        RECT 513.200 176.000 514.000 179.800 ;
        RECT 516.400 176.000 517.200 179.800 ;
        RECT 513.200 175.800 517.200 176.000 ;
        RECT 518.000 177.000 518.800 179.000 ;
        RECT 505.400 175.400 509.000 175.800 ;
        RECT 506.000 174.400 506.800 174.800 ;
        RECT 510.000 174.400 510.600 175.800 ;
        RECT 511.800 174.400 512.400 175.800 ;
        RECT 513.400 175.400 517.000 175.800 ;
        RECT 518.000 174.800 518.600 177.000 ;
        RECT 522.200 176.400 523.000 179.000 ;
        RECT 521.200 176.000 523.000 176.400 ;
        RECT 527.600 177.000 528.400 179.000 ;
        RECT 521.200 175.600 523.800 176.000 ;
        RECT 522.200 175.400 523.800 175.600 ;
        RECT 523.000 175.000 523.800 175.400 ;
        RECT 515.600 174.400 516.400 174.800 ;
        RECT 502.000 174.200 503.600 174.400 ;
        RECT 492.600 173.600 503.600 174.200 ;
        RECT 505.200 173.800 506.800 174.400 ;
        RECT 505.200 173.600 506.000 173.800 ;
        RECT 508.200 173.600 510.800 174.400 ;
        RECT 511.600 173.600 514.200 174.400 ;
        RECT 515.600 173.800 517.200 174.400 ;
        RECT 518.000 174.200 522.200 174.800 ;
        RECT 516.400 173.600 517.200 173.800 ;
        RECT 521.200 173.800 522.200 174.200 ;
        RECT 523.200 174.400 523.800 175.000 ;
        RECT 527.600 174.800 528.200 177.000 ;
        RECT 531.800 176.000 532.600 179.000 ;
        RECT 537.200 176.000 538.000 179.800 ;
        RECT 540.400 176.000 541.200 179.800 ;
        RECT 531.800 175.400 533.400 176.000 ;
        RECT 537.200 175.800 541.200 176.000 ;
        RECT 542.000 175.800 542.800 179.800 ;
        RECT 543.600 176.000 544.400 179.800 ;
        RECT 546.800 176.000 547.600 179.800 ;
        RECT 543.600 175.800 547.600 176.000 ;
        RECT 548.400 175.800 549.200 179.800 ;
        RECT 537.400 175.400 541.000 175.800 ;
        RECT 532.600 175.000 533.400 175.400 ;
        RECT 490.800 172.800 491.600 173.000 ;
        RECT 487.800 172.200 491.600 172.800 ;
        RECT 487.800 172.000 488.600 172.200 ;
        RECT 489.400 171.400 490.200 171.600 ;
        RECT 481.400 170.400 485.200 171.000 ;
        RECT 448.600 162.200 449.400 169.600 ;
        RECT 450.200 168.400 450.800 169.600 ;
        RECT 450.000 167.600 450.800 168.400 ;
        RECT 453.200 168.400 453.800 169.600 ;
        RECT 453.200 167.600 454.000 168.400 ;
        RECT 454.600 162.200 455.400 169.600 ;
        RECT 466.200 162.200 467.000 169.600 ;
        RECT 467.800 168.400 468.400 169.600 ;
        RECT 467.600 167.600 468.400 168.400 ;
        RECT 472.600 162.200 473.400 169.600 ;
        RECT 474.200 168.400 474.800 169.600 ;
        RECT 479.400 169.200 481.000 169.800 ;
        RECT 474.000 167.600 474.800 168.400 ;
        RECT 480.200 162.200 481.000 169.200 ;
        RECT 484.600 167.000 485.200 170.400 ;
        RECT 484.400 163.000 485.200 167.000 ;
        RECT 486.000 170.800 490.200 171.400 ;
        RECT 486.000 162.200 486.800 170.800 ;
        RECT 492.600 170.400 493.200 173.600 ;
        RECT 499.800 173.400 500.600 173.600 ;
        RECT 501.400 172.400 502.200 172.600 ;
        RECT 497.200 171.800 502.200 172.400 ;
        RECT 497.200 171.600 498.000 171.800 ;
        RECT 506.800 171.600 507.600 173.200 ;
        RECT 498.800 171.000 504.400 171.200 ;
        RECT 498.600 170.800 504.400 171.000 ;
        RECT 490.800 169.800 493.200 170.400 ;
        RECT 494.600 170.600 504.400 170.800 ;
        RECT 494.600 170.200 499.400 170.600 ;
        RECT 490.800 168.800 491.400 169.800 ;
        RECT 490.000 168.400 491.400 168.800 ;
        RECT 493.000 169.000 493.800 169.200 ;
        RECT 494.600 169.000 495.200 170.200 ;
        RECT 493.000 168.400 495.200 169.000 ;
        RECT 495.800 169.000 501.200 169.600 ;
        RECT 495.800 168.800 496.600 169.000 ;
        RECT 500.400 168.800 501.200 169.000 ;
        RECT 489.200 168.000 491.400 168.400 ;
        RECT 489.200 167.600 490.600 168.000 ;
        RECT 494.200 167.400 495.000 167.600 ;
        RECT 497.000 167.400 497.800 167.600 ;
        RECT 490.800 166.200 491.600 167.000 ;
        RECT 494.200 166.800 497.800 167.400 ;
        RECT 495.000 166.200 495.600 166.800 ;
        RECT 500.400 166.200 501.200 167.000 ;
        RECT 490.200 162.200 491.400 166.200 ;
        RECT 494.800 162.200 495.600 166.200 ;
        RECT 499.200 165.600 501.200 166.200 ;
        RECT 499.200 162.200 500.000 165.600 ;
        RECT 503.600 162.200 504.400 170.600 ;
        RECT 508.200 170.200 508.800 173.600 ;
        RECT 513.600 172.300 514.200 173.600 ;
        RECT 510.100 171.700 514.200 172.300 ;
        RECT 510.100 170.400 510.700 171.700 ;
        RECT 510.000 170.200 510.800 170.400 ;
        RECT 507.800 169.600 508.800 170.200 ;
        RECT 509.400 169.600 510.800 170.200 ;
        RECT 511.600 170.200 512.400 170.400 ;
        RECT 513.600 170.200 514.200 171.700 ;
        RECT 514.800 171.600 515.600 173.200 ;
        RECT 518.000 171.600 518.800 173.200 ;
        RECT 519.600 171.600 520.400 173.200 ;
        RECT 521.200 173.000 522.600 173.800 ;
        RECT 523.200 173.600 525.200 174.400 ;
        RECT 527.600 174.200 531.800 174.800 ;
        RECT 530.800 173.800 531.800 174.200 ;
        RECT 532.800 174.400 533.400 175.000 ;
        RECT 538.000 174.400 538.800 174.800 ;
        RECT 542.000 174.400 542.600 175.800 ;
        RECT 543.800 175.400 547.400 175.800 ;
        RECT 544.400 174.400 545.200 174.800 ;
        RECT 548.400 174.400 549.000 175.800 ;
        RECT 521.200 171.000 521.800 173.000 ;
        RECT 518.000 170.400 521.800 171.000 ;
        RECT 511.600 169.600 513.000 170.200 ;
        RECT 513.600 169.600 514.600 170.200 ;
        RECT 507.800 162.200 508.600 169.600 ;
        RECT 509.400 168.400 510.000 169.600 ;
        RECT 509.200 167.600 510.000 168.400 ;
        RECT 512.400 168.400 513.000 169.600 ;
        RECT 512.400 167.600 513.200 168.400 ;
        RECT 513.800 162.200 514.600 169.600 ;
        RECT 518.000 167.000 518.600 170.400 ;
        RECT 523.200 169.800 523.800 173.600 ;
        RECT 524.400 170.800 525.200 172.400 ;
        RECT 527.600 171.600 528.400 173.200 ;
        RECT 529.200 171.600 530.000 173.200 ;
        RECT 530.800 173.000 532.200 173.800 ;
        RECT 532.800 173.600 534.800 174.400 ;
        RECT 537.200 173.800 538.800 174.400 ;
        RECT 537.200 173.600 538.000 173.800 ;
        RECT 540.200 173.600 542.800 174.400 ;
        RECT 543.600 173.800 545.200 174.400 ;
        RECT 543.600 173.600 544.400 173.800 ;
        RECT 546.600 173.600 549.200 174.400 ;
        RECT 530.800 171.000 531.400 173.000 ;
        RECT 522.200 169.200 523.800 169.800 ;
        RECT 527.600 170.400 531.400 171.000 ;
        RECT 518.000 163.000 518.800 167.000 ;
        RECT 522.200 162.200 523.000 169.200 ;
        RECT 527.600 167.000 528.200 170.400 ;
        RECT 532.800 169.800 533.400 173.600 ;
        RECT 534.000 170.800 534.800 172.400 ;
        RECT 538.800 171.600 539.600 173.200 ;
        RECT 540.200 172.400 540.800 173.600 ;
        RECT 540.200 171.600 541.200 172.400 ;
        RECT 545.200 171.600 546.000 173.200 ;
        RECT 540.200 170.200 540.800 171.600 ;
        RECT 546.600 170.400 547.200 173.600 ;
        RECT 542.000 170.200 542.800 170.400 ;
        RECT 531.800 169.200 533.400 169.800 ;
        RECT 539.800 169.600 540.800 170.200 ;
        RECT 541.400 169.600 542.800 170.200 ;
        RECT 545.200 169.600 547.200 170.400 ;
        RECT 548.400 170.200 549.200 170.400 ;
        RECT 547.800 169.600 549.200 170.200 ;
        RECT 527.600 163.000 528.400 167.000 ;
        RECT 531.800 164.400 532.600 169.200 ;
        RECT 531.800 163.600 533.200 164.400 ;
        RECT 531.800 162.200 532.600 163.600 ;
        RECT 539.800 162.200 540.600 169.600 ;
        RECT 541.400 168.400 542.000 169.600 ;
        RECT 541.200 167.600 542.000 168.400 ;
        RECT 546.200 162.200 547.000 169.600 ;
        RECT 547.800 168.400 548.400 169.600 ;
        RECT 547.600 167.600 548.400 168.400 ;
        RECT 550.000 162.200 550.800 179.800 ;
        RECT 555.800 178.400 556.600 179.800 ;
        RECT 554.800 177.600 556.600 178.400 ;
        RECT 551.600 175.600 552.400 177.200 ;
        RECT 555.800 176.400 556.600 177.600 ;
        RECT 554.800 175.800 556.600 176.400 ;
        RECT 558.000 176.000 558.800 179.800 ;
        RECT 561.200 176.000 562.000 179.800 ;
        RECT 558.000 175.800 562.000 176.000 ;
        RECT 562.800 175.800 563.600 179.800 ;
        RECT 566.000 176.000 566.800 179.800 ;
        RECT 551.600 174.300 552.400 174.400 ;
        RECT 553.200 174.300 554.000 175.200 ;
        RECT 551.600 173.700 554.000 174.300 ;
        RECT 551.600 173.600 552.400 173.700 ;
        RECT 553.200 173.600 554.000 173.700 ;
        RECT 554.800 162.200 555.600 175.800 ;
        RECT 558.200 175.400 561.800 175.800 ;
        RECT 558.800 174.400 559.600 174.800 ;
        RECT 562.800 174.400 563.400 175.800 ;
        RECT 565.800 175.200 566.800 176.000 ;
        RECT 558.000 173.800 559.600 174.400 ;
        RECT 558.000 173.600 558.800 173.800 ;
        RECT 561.000 173.600 563.600 174.400 ;
        RECT 559.600 171.600 560.400 173.200 ;
        RECT 561.000 172.300 561.600 173.600 ;
        RECT 564.400 172.300 565.200 172.400 ;
        RECT 561.000 171.700 565.200 172.300 ;
        RECT 556.400 168.800 557.200 170.400 ;
        RECT 561.000 170.200 561.600 171.700 ;
        RECT 564.400 171.600 565.200 171.700 ;
        RECT 565.800 170.800 566.600 175.200 ;
        RECT 567.600 174.600 568.400 179.800 ;
        RECT 574.000 176.600 574.800 179.800 ;
        RECT 575.600 177.000 576.400 179.800 ;
        RECT 577.200 177.000 578.000 179.800 ;
        RECT 578.800 177.000 579.600 179.800 ;
        RECT 580.400 177.000 581.200 179.800 ;
        RECT 583.600 177.000 584.400 179.800 ;
        RECT 586.800 177.000 587.600 179.800 ;
        RECT 588.400 177.000 589.200 179.800 ;
        RECT 590.000 177.000 590.800 179.800 ;
        RECT 572.400 175.800 574.800 176.600 ;
        RECT 591.600 176.600 592.400 179.800 ;
        RECT 572.400 175.200 573.200 175.800 ;
        RECT 567.200 174.000 568.400 174.600 ;
        RECT 571.400 174.600 573.200 175.200 ;
        RECT 577.200 175.600 578.200 176.400 ;
        RECT 581.200 175.600 582.800 176.400 ;
        RECT 583.600 175.800 588.200 176.400 ;
        RECT 591.600 175.800 594.200 176.600 ;
        RECT 583.600 175.600 584.400 175.800 ;
        RECT 567.200 172.000 567.800 174.000 ;
        RECT 571.400 173.400 572.200 174.600 ;
        RECT 568.400 172.600 572.200 173.400 ;
        RECT 577.200 172.800 578.000 175.600 ;
        RECT 583.600 174.800 584.400 175.000 ;
        RECT 580.000 174.200 584.400 174.800 ;
        RECT 580.000 174.000 580.800 174.200 ;
        RECT 585.200 173.600 586.000 175.200 ;
        RECT 587.400 173.400 588.200 175.800 ;
        RECT 593.400 175.200 594.200 175.800 ;
        RECT 593.400 174.400 596.400 175.200 ;
        RECT 598.000 173.800 598.800 179.800 ;
        RECT 599.600 175.800 600.400 179.800 ;
        RECT 601.200 176.000 602.000 179.800 ;
        RECT 604.400 176.000 605.200 179.800 ;
        RECT 601.200 175.800 605.200 176.000 ;
        RECT 599.800 174.400 600.400 175.800 ;
        RECT 601.400 175.400 605.000 175.800 ;
        RECT 603.600 174.400 604.400 174.800 ;
        RECT 580.400 172.600 583.600 173.400 ;
        RECT 587.400 172.600 589.400 173.400 ;
        RECT 590.000 173.000 598.800 173.800 ;
        RECT 599.600 173.600 602.200 174.400 ;
        RECT 603.600 174.300 605.200 174.400 ;
        RECT 606.000 174.300 606.800 179.800 ;
        RECT 603.600 173.800 606.800 174.300 ;
        RECT 604.400 173.700 606.800 173.800 ;
        RECT 604.400 173.600 605.200 173.700 ;
        RECT 574.000 172.000 574.800 172.600 ;
        RECT 591.600 172.000 592.400 172.400 ;
        RECT 594.800 172.000 595.600 172.400 ;
        RECT 596.600 172.000 597.400 172.200 ;
        RECT 567.200 171.400 568.000 172.000 ;
        RECT 574.000 171.400 597.400 172.000 ;
        RECT 562.800 170.300 563.600 170.400 ;
        RECT 565.800 170.300 566.800 170.800 ;
        RECT 562.800 170.200 566.800 170.300 ;
        RECT 560.600 169.600 561.600 170.200 ;
        RECT 562.200 169.700 566.800 170.200 ;
        RECT 562.200 169.600 563.600 169.700 ;
        RECT 560.600 162.200 561.400 169.600 ;
        RECT 562.200 168.400 562.800 169.600 ;
        RECT 562.000 167.600 562.800 168.400 ;
        RECT 566.000 162.200 566.800 169.700 ;
        RECT 567.400 169.600 568.000 171.400 ;
        RECT 567.400 169.000 576.400 169.600 ;
        RECT 567.400 167.400 568.000 169.000 ;
        RECT 575.600 168.800 576.400 169.000 ;
        RECT 578.800 169.000 587.400 169.600 ;
        RECT 578.800 168.800 579.600 169.000 ;
        RECT 570.600 167.600 573.200 168.400 ;
        RECT 567.400 166.800 570.000 167.400 ;
        RECT 569.200 162.200 570.000 166.800 ;
        RECT 572.400 162.200 573.200 167.600 ;
        RECT 573.800 166.800 578.000 167.600 ;
        RECT 575.600 162.200 576.400 165.000 ;
        RECT 577.200 162.200 578.000 165.000 ;
        RECT 578.800 162.200 579.600 165.000 ;
        RECT 580.400 162.200 581.200 168.400 ;
        RECT 583.600 167.600 586.200 168.400 ;
        RECT 586.800 168.200 587.400 169.000 ;
        RECT 588.400 169.400 589.200 169.600 ;
        RECT 588.400 169.000 593.800 169.400 ;
        RECT 588.400 168.800 594.600 169.000 ;
        RECT 593.200 168.200 594.600 168.800 ;
        RECT 586.800 167.600 592.600 168.200 ;
        RECT 595.600 168.000 597.200 168.800 ;
        RECT 595.600 167.600 596.200 168.000 ;
        RECT 583.600 162.200 584.400 167.000 ;
        RECT 586.800 162.200 587.600 167.000 ;
        RECT 592.000 166.800 596.200 167.600 ;
        RECT 598.000 167.400 598.800 173.000 ;
        RECT 599.600 170.200 600.400 170.400 ;
        RECT 601.600 170.200 602.200 173.600 ;
        RECT 602.800 171.600 603.600 173.200 ;
        RECT 599.600 169.600 601.000 170.200 ;
        RECT 601.600 169.600 602.600 170.200 ;
        RECT 600.400 168.400 601.000 169.600 ;
        RECT 600.400 167.600 601.200 168.400 ;
        RECT 596.800 166.800 598.800 167.400 ;
        RECT 588.400 162.200 589.200 165.000 ;
        RECT 590.000 162.200 590.800 165.000 ;
        RECT 593.200 162.200 594.000 166.800 ;
        RECT 596.800 166.200 597.400 166.800 ;
        RECT 596.400 165.600 597.400 166.200 ;
        RECT 596.400 162.200 597.200 165.600 ;
        RECT 601.800 162.200 602.600 169.600 ;
        RECT 606.000 162.200 606.800 173.700 ;
        RECT 1.200 151.400 2.000 159.800 ;
        RECT 5.600 156.400 6.400 159.800 ;
        RECT 4.400 155.800 6.400 156.400 ;
        RECT 10.000 155.800 10.800 159.800 ;
        RECT 14.200 155.800 15.400 159.800 ;
        RECT 4.400 155.000 5.200 155.800 ;
        RECT 10.000 155.200 10.600 155.800 ;
        RECT 7.800 154.600 11.400 155.200 ;
        RECT 14.000 155.000 14.800 155.800 ;
        RECT 7.800 154.400 8.600 154.600 ;
        RECT 10.600 154.400 11.400 154.600 ;
        RECT 4.400 153.000 5.200 153.200 ;
        RECT 9.000 153.000 9.800 153.200 ;
        RECT 4.400 152.400 9.800 153.000 ;
        RECT 10.400 153.000 12.600 153.600 ;
        RECT 10.400 151.800 11.000 153.000 ;
        RECT 11.800 152.800 12.600 153.000 ;
        RECT 14.200 153.200 15.600 154.000 ;
        RECT 14.200 152.200 14.800 153.200 ;
        RECT 6.200 151.400 11.000 151.800 ;
        RECT 1.200 151.200 11.000 151.400 ;
        RECT 12.400 151.600 14.800 152.200 ;
        RECT 1.200 151.000 7.000 151.200 ;
        RECT 1.200 150.800 6.800 151.000 ;
        RECT 7.600 150.200 8.400 150.400 ;
        RECT 3.400 149.600 8.400 150.200 ;
        RECT 3.400 149.400 4.200 149.600 ;
        RECT 5.000 148.400 5.800 148.600 ;
        RECT 12.400 148.400 13.000 151.600 ;
        RECT 18.800 151.200 19.600 159.800 ;
        RECT 22.600 158.400 23.400 159.800 ;
        RECT 22.600 157.600 24.400 158.400 ;
        RECT 21.200 153.600 22.000 154.400 ;
        RECT 21.200 152.400 21.800 153.600 ;
        RECT 22.600 152.400 23.400 157.600 ;
        RECT 20.400 151.800 21.800 152.400 ;
        RECT 22.400 151.800 23.400 152.400 ;
        RECT 29.400 152.400 30.200 159.800 ;
        RECT 30.800 153.600 31.600 154.400 ;
        RECT 31.000 152.400 31.600 153.600 ;
        RECT 34.000 153.600 34.800 154.400 ;
        RECT 34.000 152.400 34.600 153.600 ;
        RECT 35.400 152.400 36.200 159.800 ;
        RECT 43.400 152.800 44.200 159.800 ;
        RECT 47.600 155.000 48.400 159.000 ;
        RECT 29.400 151.800 30.400 152.400 ;
        RECT 31.000 151.800 32.400 152.400 ;
        RECT 20.400 151.600 21.200 151.800 ;
        RECT 15.400 150.600 19.600 151.200 ;
        RECT 15.400 150.400 16.200 150.600 ;
        RECT 17.000 149.800 17.800 150.000 ;
        RECT 14.000 149.200 17.800 149.800 ;
        RECT 14.000 149.000 14.800 149.200 ;
        RECT 2.000 147.800 13.000 148.400 ;
        RECT 2.000 147.600 3.600 147.800 ;
        RECT 6.000 147.600 6.800 147.800 ;
        RECT 11.800 147.600 12.600 147.800 ;
        RECT 1.200 142.200 2.000 147.000 ;
        RECT 6.200 145.600 6.800 147.600 ;
        RECT 18.800 147.200 19.600 150.600 ;
        RECT 22.400 148.400 23.000 151.800 ;
        RECT 23.600 150.300 24.400 150.400 ;
        RECT 28.400 150.300 29.200 150.400 ;
        RECT 23.600 149.700 29.200 150.300 ;
        RECT 23.600 148.800 24.400 149.700 ;
        RECT 28.400 148.800 29.200 149.700 ;
        RECT 29.800 150.300 30.400 151.800 ;
        RECT 31.600 151.600 32.400 151.800 ;
        RECT 33.200 151.800 34.600 152.400 ;
        RECT 35.200 151.800 36.200 152.400 ;
        RECT 42.600 152.200 44.200 152.800 ;
        RECT 33.200 151.600 34.000 151.800 ;
        RECT 33.300 150.300 33.900 151.600 ;
        RECT 29.800 149.700 33.900 150.300 ;
        RECT 29.800 148.400 30.400 149.700 ;
        RECT 35.200 148.400 35.800 151.800 ;
        RECT 36.400 148.800 37.200 150.400 ;
        RECT 39.600 150.300 40.400 150.400 ;
        RECT 41.200 150.300 42.000 151.200 ;
        RECT 39.600 149.700 42.000 150.300 ;
        RECT 39.600 149.600 40.400 149.700 ;
        RECT 41.200 149.600 42.000 149.700 ;
        RECT 42.600 148.400 43.200 152.200 ;
        RECT 47.800 151.600 48.400 155.000 ;
        RECT 53.000 152.800 53.800 159.800 ;
        RECT 57.200 155.000 58.000 159.000 ;
        RECT 44.600 151.000 48.400 151.600 ;
        RECT 52.200 152.200 53.800 152.800 ;
        RECT 44.600 149.000 45.200 151.000 ;
        RECT 20.400 147.600 23.000 148.400 ;
        RECT 25.200 148.300 26.000 148.400 ;
        RECT 26.800 148.300 27.600 148.400 ;
        RECT 25.200 148.200 27.600 148.300 ;
        RECT 24.400 147.700 28.400 148.200 ;
        RECT 24.400 147.600 26.000 147.700 ;
        RECT 26.800 147.600 28.400 147.700 ;
        RECT 29.800 147.600 32.400 148.400 ;
        RECT 33.200 147.600 35.800 148.400 ;
        RECT 38.000 148.200 38.800 148.400 ;
        RECT 37.200 147.600 38.800 148.200 ;
        RECT 39.600 148.300 40.400 148.400 ;
        RECT 41.200 148.300 43.200 148.400 ;
        RECT 39.600 147.700 43.200 148.300 ;
        RECT 43.800 148.200 45.200 149.000 ;
        RECT 46.000 148.800 46.800 150.400 ;
        RECT 47.600 148.800 48.400 150.400 ;
        RECT 50.800 149.600 51.600 151.200 ;
        RECT 52.200 148.400 52.800 152.200 ;
        RECT 57.400 151.600 58.000 155.000 ;
        RECT 61.400 152.400 62.200 159.800 ;
        RECT 62.800 153.600 63.600 154.400 ;
        RECT 63.000 152.400 63.600 153.600 ;
        RECT 66.000 153.600 66.800 154.400 ;
        RECT 66.000 152.400 66.600 153.600 ;
        RECT 67.400 152.400 68.200 159.800 ;
        RECT 61.400 151.800 62.400 152.400 ;
        RECT 63.000 151.800 64.400 152.400 ;
        RECT 54.200 151.000 58.000 151.600 ;
        RECT 54.200 149.000 54.800 151.000 ;
        RECT 39.600 147.600 40.400 147.700 ;
        RECT 41.200 147.600 43.200 147.700 ;
        RECT 15.800 146.600 19.600 147.200 ;
        RECT 15.800 146.400 16.600 146.600 ;
        RECT 4.400 144.200 5.200 145.000 ;
        RECT 6.000 144.800 6.800 145.600 ;
        RECT 7.800 145.400 8.600 145.600 ;
        RECT 7.800 144.800 10.600 145.400 ;
        RECT 10.000 144.200 10.600 144.800 ;
        RECT 14.000 144.200 14.800 145.000 ;
        RECT 4.400 143.600 6.400 144.200 ;
        RECT 5.600 142.200 6.400 143.600 ;
        RECT 10.000 142.200 10.800 144.200 ;
        RECT 14.000 143.600 15.400 144.200 ;
        RECT 14.200 142.200 15.400 143.600 ;
        RECT 18.800 142.200 19.600 146.600 ;
        RECT 20.600 146.200 21.200 147.600 ;
        RECT 24.400 147.200 25.200 147.600 ;
        RECT 27.600 147.200 28.400 147.600 ;
        RECT 22.200 146.200 25.800 146.600 ;
        RECT 27.000 146.200 30.600 146.600 ;
        RECT 31.600 146.200 32.200 147.600 ;
        RECT 33.400 146.200 34.000 147.600 ;
        RECT 37.200 147.200 38.000 147.600 ;
        RECT 42.600 147.000 43.200 147.600 ;
        RECT 44.200 147.800 45.200 148.200 ;
        RECT 44.200 147.200 48.400 147.800 ;
        RECT 50.800 147.600 52.800 148.400 ;
        RECT 53.400 148.200 54.800 149.000 ;
        RECT 55.600 148.800 56.400 150.400 ;
        RECT 57.200 148.800 58.000 150.400 ;
        RECT 60.400 148.800 61.200 150.400 ;
        RECT 61.800 150.300 62.400 151.800 ;
        RECT 63.600 151.600 64.400 151.800 ;
        RECT 65.200 151.800 66.600 152.400 ;
        RECT 67.200 151.800 68.200 152.400 ;
        RECT 65.200 151.600 66.000 151.800 ;
        RECT 65.300 150.300 65.900 151.600 ;
        RECT 67.200 150.400 67.800 151.800 ;
        RECT 71.600 151.400 72.400 159.800 ;
        RECT 76.000 156.400 76.800 159.800 ;
        RECT 74.800 155.800 76.800 156.400 ;
        RECT 80.400 155.800 81.200 159.800 ;
        RECT 84.600 155.800 85.800 159.800 ;
        RECT 74.800 155.000 75.600 155.800 ;
        RECT 80.400 155.200 81.000 155.800 ;
        RECT 78.200 154.600 81.800 155.200 ;
        RECT 84.400 155.000 85.200 155.800 ;
        RECT 78.200 154.400 79.000 154.600 ;
        RECT 81.000 154.400 81.800 154.600 ;
        RECT 74.800 153.000 75.600 153.200 ;
        RECT 79.400 153.000 80.200 153.200 ;
        RECT 74.800 152.400 80.200 153.000 ;
        RECT 80.800 153.000 83.000 153.600 ;
        RECT 80.800 151.800 81.400 153.000 ;
        RECT 82.200 152.800 83.000 153.000 ;
        RECT 84.600 153.200 86.000 154.000 ;
        RECT 84.600 152.200 85.200 153.200 ;
        RECT 76.600 151.400 81.400 151.800 ;
        RECT 71.600 151.200 81.400 151.400 ;
        RECT 82.800 151.600 85.200 152.200 ;
        RECT 89.200 152.300 90.000 159.800 ;
        RECT 92.400 155.800 93.200 159.800 ;
        RECT 92.600 155.600 93.200 155.800 ;
        RECT 95.600 155.800 96.400 159.800 ;
        RECT 95.600 155.600 96.200 155.800 ;
        RECT 92.600 155.000 96.200 155.600 ;
        RECT 94.000 152.800 94.800 154.400 ;
        RECT 95.600 152.400 96.200 155.000 ;
        RECT 99.800 152.400 100.600 159.800 ;
        RECT 105.200 155.800 106.000 159.800 ;
        RECT 105.400 155.600 106.000 155.800 ;
        RECT 108.400 155.800 109.200 159.800 ;
        RECT 108.400 155.600 109.000 155.800 ;
        RECT 105.400 155.000 109.000 155.600 ;
        RECT 101.200 153.600 102.000 154.400 ;
        RECT 101.400 152.400 102.000 153.600 ;
        RECT 106.800 152.800 107.600 154.400 ;
        RECT 108.400 152.400 109.000 155.000 ;
        RECT 112.600 154.400 113.400 159.800 ;
        RECT 111.600 153.600 113.400 154.400 ;
        RECT 114.000 153.600 114.800 154.400 ;
        RECT 112.600 152.400 113.400 153.600 ;
        RECT 114.200 152.400 114.800 153.600 ;
        RECT 117.200 153.600 118.000 154.400 ;
        RECT 117.200 152.400 117.800 153.600 ;
        RECT 118.600 152.400 119.400 159.800 ;
        RECT 90.800 152.300 91.600 152.400 ;
        RECT 89.200 151.700 91.600 152.300 ;
        RECT 71.600 151.000 77.400 151.200 ;
        RECT 71.600 150.800 77.200 151.000 ;
        RECT 61.800 149.700 65.900 150.300 ;
        RECT 61.800 148.400 62.400 149.700 ;
        RECT 66.800 149.600 67.800 150.400 ;
        RECT 67.200 148.400 67.800 149.600 ;
        RECT 68.400 148.800 69.200 150.400 ;
        RECT 78.000 150.200 78.800 150.400 ;
        RECT 73.800 149.600 78.800 150.200 ;
        RECT 73.800 149.400 74.600 149.600 ;
        RECT 76.400 149.400 77.200 149.600 ;
        RECT 75.400 148.400 76.200 148.600 ;
        RECT 82.800 148.400 83.400 151.600 ;
        RECT 89.200 151.200 90.000 151.700 ;
        RECT 85.800 150.600 90.000 151.200 ;
        RECT 90.800 150.800 91.600 151.700 ;
        RECT 95.600 151.600 96.400 152.400 ;
        RECT 99.800 151.800 100.800 152.400 ;
        RECT 101.400 151.800 102.800 152.400 ;
        RECT 85.800 150.400 86.600 150.600 ;
        RECT 87.400 149.800 88.200 150.000 ;
        RECT 84.400 149.200 88.200 149.800 ;
        RECT 84.400 149.000 85.200 149.200 ;
        RECT 42.600 146.600 43.400 147.000 ;
        RECT 35.000 146.200 38.600 146.600 ;
        RECT 20.400 142.200 21.200 146.200 ;
        RECT 22.000 146.000 26.000 146.200 ;
        RECT 22.000 142.200 22.800 146.000 ;
        RECT 25.200 142.200 26.000 146.000 ;
        RECT 26.800 146.000 30.800 146.200 ;
        RECT 26.800 142.200 27.600 146.000 ;
        RECT 30.000 142.200 30.800 146.000 ;
        RECT 31.600 142.200 32.400 146.200 ;
        RECT 33.200 142.200 34.000 146.200 ;
        RECT 34.800 146.000 38.800 146.200 ;
        RECT 42.600 146.000 44.200 146.600 ;
        RECT 34.800 142.200 35.600 146.000 ;
        RECT 38.000 142.200 38.800 146.000 ;
        RECT 43.400 143.000 44.200 146.000 ;
        RECT 47.800 145.000 48.400 147.200 ;
        RECT 52.200 147.000 52.800 147.600 ;
        RECT 53.800 147.800 54.800 148.200 ;
        RECT 58.800 148.200 59.600 148.400 ;
        RECT 53.800 147.200 58.000 147.800 ;
        RECT 58.800 147.600 60.400 148.200 ;
        RECT 61.800 147.600 64.400 148.400 ;
        RECT 65.200 147.600 67.800 148.400 ;
        RECT 70.000 148.200 70.800 148.400 ;
        RECT 69.200 147.600 70.800 148.200 ;
        RECT 72.400 147.800 83.400 148.400 ;
        RECT 72.400 147.600 74.000 147.800 ;
        RECT 59.600 147.200 60.400 147.600 ;
        RECT 52.200 146.600 53.000 147.000 ;
        RECT 52.200 146.400 53.800 146.600 ;
        RECT 52.200 146.000 54.800 146.400 ;
        RECT 47.600 143.000 48.400 145.000 ;
        RECT 53.000 145.600 54.800 146.000 ;
        RECT 53.000 143.000 53.800 145.600 ;
        RECT 57.400 145.000 58.000 147.200 ;
        RECT 59.000 146.200 62.600 146.600 ;
        RECT 63.600 146.200 64.200 147.600 ;
        RECT 65.400 146.200 66.000 147.600 ;
        RECT 69.200 147.200 70.000 147.600 ;
        RECT 67.000 146.200 70.600 146.600 ;
        RECT 57.200 143.000 58.000 145.000 ;
        RECT 58.800 146.000 62.800 146.200 ;
        RECT 58.800 142.200 59.600 146.000 ;
        RECT 62.000 142.200 62.800 146.000 ;
        RECT 63.600 142.200 64.400 146.200 ;
        RECT 65.200 142.200 66.000 146.200 ;
        RECT 66.800 146.000 70.800 146.200 ;
        RECT 66.800 142.200 67.600 146.000 ;
        RECT 70.000 142.200 70.800 146.000 ;
        RECT 71.600 142.200 72.400 147.000 ;
        RECT 76.600 146.400 77.200 147.800 ;
        RECT 82.200 147.600 83.000 147.800 ;
        RECT 89.200 147.200 90.000 150.600 ;
        RECT 92.400 149.600 94.000 150.400 ;
        RECT 95.600 148.400 96.200 151.600 ;
        RECT 98.800 148.800 99.600 150.400 ;
        RECT 100.200 148.400 100.800 151.800 ;
        RECT 102.000 151.600 102.800 151.800 ;
        RECT 103.600 150.800 104.400 152.400 ;
        RECT 108.400 151.600 109.200 152.400 ;
        RECT 112.600 151.800 113.600 152.400 ;
        RECT 114.200 151.800 115.600 152.400 ;
        RECT 105.200 149.600 106.800 150.400 ;
        RECT 108.400 148.400 109.000 151.600 ;
        RECT 111.600 148.800 112.400 150.400 ;
        RECT 113.000 148.400 113.600 151.800 ;
        RECT 114.800 151.600 115.600 151.800 ;
        RECT 116.400 151.800 117.800 152.400 ;
        RECT 118.400 151.800 119.400 152.400 ;
        RECT 125.400 152.400 126.200 159.800 ;
        RECT 126.800 153.600 127.600 154.400 ;
        RECT 127.000 152.400 127.600 153.600 ;
        RECT 131.800 152.400 132.600 159.800 ;
        RECT 138.200 158.400 139.000 159.800 ;
        RECT 137.200 157.600 139.000 158.400 ;
        RECT 133.200 153.600 134.000 154.400 ;
        RECT 133.400 152.400 134.000 153.600 ;
        RECT 138.200 152.400 139.000 157.600 ;
        RECT 139.600 153.600 140.400 154.400 ;
        RECT 139.800 152.400 140.400 153.600 ;
        RECT 125.400 151.800 126.400 152.400 ;
        RECT 127.000 151.800 128.400 152.400 ;
        RECT 116.400 151.600 117.200 151.800 ;
        RECT 118.400 150.400 119.000 151.800 ;
        RECT 118.000 149.600 119.000 150.400 ;
        RECT 118.400 148.400 119.000 149.600 ;
        RECT 119.600 148.800 120.400 150.400 ;
        RECT 124.400 148.800 125.200 150.400 ;
        RECT 125.800 148.400 126.400 151.800 ;
        RECT 127.600 151.600 128.400 151.800 ;
        RECT 130.800 151.600 132.800 152.400 ;
        RECT 133.400 151.800 134.800 152.400 ;
        RECT 138.200 151.800 139.200 152.400 ;
        RECT 139.800 151.800 141.200 152.400 ;
        RECT 134.000 151.600 134.800 151.800 ;
        RECT 127.600 150.300 128.400 150.400 ;
        RECT 127.600 149.700 129.900 150.300 ;
        RECT 127.600 149.600 128.400 149.700 ;
        RECT 129.300 148.400 129.900 149.700 ;
        RECT 130.800 148.800 131.600 150.400 ;
        RECT 132.200 148.400 132.800 151.600 ;
        RECT 137.200 148.800 138.000 150.400 ;
        RECT 138.600 148.400 139.200 151.800 ;
        RECT 140.400 151.600 141.200 151.800 ;
        RECT 94.600 148.200 96.200 148.400 ;
        RECT 86.200 146.600 90.000 147.200 ;
        RECT 86.200 146.400 87.000 146.600 ;
        RECT 74.800 144.200 75.600 145.000 ;
        RECT 76.400 144.800 77.200 146.400 ;
        RECT 78.200 145.400 79.000 145.600 ;
        RECT 78.200 144.800 81.000 145.400 ;
        RECT 80.400 144.200 81.000 144.800 ;
        RECT 84.400 144.200 85.200 145.000 ;
        RECT 74.800 143.600 76.800 144.200 ;
        RECT 76.000 142.200 76.800 143.600 ;
        RECT 80.400 142.200 81.200 144.200 ;
        RECT 84.400 143.600 85.800 144.200 ;
        RECT 84.600 142.200 85.800 143.600 ;
        RECT 89.200 142.200 90.000 146.600 ;
        RECT 94.400 147.800 96.200 148.200 ;
        RECT 97.200 148.200 98.000 148.400 ;
        RECT 94.400 142.200 95.200 147.800 ;
        RECT 97.200 147.600 98.800 148.200 ;
        RECT 100.200 147.600 102.800 148.400 ;
        RECT 107.400 148.200 109.000 148.400 ;
        RECT 107.200 147.800 109.000 148.200 ;
        RECT 110.000 148.200 110.800 148.400 ;
        RECT 98.000 147.200 98.800 147.600 ;
        RECT 97.400 146.200 101.000 146.600 ;
        RECT 102.000 146.200 102.600 147.600 ;
        RECT 97.200 146.000 101.200 146.200 ;
        RECT 97.200 142.200 98.000 146.000 ;
        RECT 100.400 142.200 101.200 146.000 ;
        RECT 102.000 142.200 102.800 146.200 ;
        RECT 107.200 142.200 108.000 147.800 ;
        RECT 110.000 147.600 111.600 148.200 ;
        RECT 113.000 147.600 115.600 148.400 ;
        RECT 116.400 147.600 119.000 148.400 ;
        RECT 121.200 148.200 122.000 148.400 ;
        RECT 120.400 147.600 122.000 148.200 ;
        RECT 122.800 148.200 123.600 148.400 ;
        RECT 122.800 147.600 124.400 148.200 ;
        RECT 125.800 147.600 128.400 148.400 ;
        RECT 129.200 148.200 130.000 148.400 ;
        RECT 129.200 147.600 130.800 148.200 ;
        RECT 132.200 147.600 134.800 148.400 ;
        RECT 135.600 148.200 136.400 148.400 ;
        RECT 135.600 147.600 137.200 148.200 ;
        RECT 138.600 147.600 141.200 148.400 ;
        RECT 110.800 147.200 111.600 147.600 ;
        RECT 110.200 146.200 113.800 146.600 ;
        RECT 114.800 146.200 115.400 147.600 ;
        RECT 116.600 146.200 117.200 147.600 ;
        RECT 120.400 147.200 121.200 147.600 ;
        RECT 123.600 147.200 124.400 147.600 ;
        RECT 118.200 146.200 121.800 146.600 ;
        RECT 123.000 146.200 126.600 146.600 ;
        RECT 127.600 146.200 128.200 147.600 ;
        RECT 130.000 147.200 130.800 147.600 ;
        RECT 129.400 146.200 133.000 146.600 ;
        RECT 134.000 146.200 134.600 147.600 ;
        RECT 136.400 147.200 137.200 147.600 ;
        RECT 135.800 146.200 139.400 146.600 ;
        RECT 140.400 146.200 141.000 147.600 ;
        RECT 142.000 146.800 142.800 148.400 ;
        RECT 143.600 148.300 144.400 159.800 ;
        RECT 145.200 152.400 146.000 159.800 ;
        RECT 149.600 158.400 151.200 159.800 ;
        RECT 149.600 157.600 152.400 158.400 ;
        RECT 146.800 152.400 147.600 152.600 ;
        RECT 149.600 152.400 151.200 157.600 ;
        RECT 145.200 151.800 147.600 152.400 ;
        RECT 149.200 151.800 151.200 152.400 ;
        RECT 153.400 152.400 154.200 152.600 ;
        RECT 154.800 152.400 155.600 159.800 ;
        RECT 162.800 156.400 163.600 159.800 ;
        RECT 162.600 155.800 163.600 156.400 ;
        RECT 162.600 155.200 163.200 155.800 ;
        RECT 166.000 155.200 166.800 159.800 ;
        RECT 169.200 157.000 170.000 159.800 ;
        RECT 170.800 157.000 171.600 159.800 ;
        RECT 153.400 151.800 155.600 152.400 ;
        RECT 161.200 154.600 163.200 155.200 ;
        RECT 149.200 150.400 149.800 151.800 ;
        RECT 153.400 151.200 154.000 151.800 ;
        RECT 150.600 150.600 154.000 151.200 ;
        RECT 150.600 150.400 151.400 150.600 ;
        RECT 148.400 149.800 149.800 150.400 ;
        RECT 152.800 149.800 153.600 150.000 ;
        RECT 148.400 149.600 150.200 149.800 ;
        RECT 149.200 149.200 150.200 149.600 ;
        RECT 145.200 148.300 146.800 148.400 ;
        RECT 143.600 147.700 146.800 148.300 ;
        RECT 110.000 146.000 114.000 146.200 ;
        RECT 110.000 142.200 110.800 146.000 ;
        RECT 113.200 142.200 114.000 146.000 ;
        RECT 114.800 142.200 115.600 146.200 ;
        RECT 116.400 142.200 117.200 146.200 ;
        RECT 118.000 146.000 122.000 146.200 ;
        RECT 118.000 142.200 118.800 146.000 ;
        RECT 121.200 142.200 122.000 146.000 ;
        RECT 122.800 146.000 126.800 146.200 ;
        RECT 122.800 142.200 123.600 146.000 ;
        RECT 126.000 142.200 126.800 146.000 ;
        RECT 127.600 142.200 128.400 146.200 ;
        RECT 129.200 146.000 133.200 146.200 ;
        RECT 129.200 142.200 130.000 146.000 ;
        RECT 132.400 142.200 133.200 146.000 ;
        RECT 134.000 142.200 134.800 146.200 ;
        RECT 135.600 146.000 139.600 146.200 ;
        RECT 135.600 142.200 136.400 146.000 ;
        RECT 138.800 142.200 139.600 146.000 ;
        RECT 140.400 142.200 141.200 146.200 ;
        RECT 143.600 142.200 144.400 147.700 ;
        RECT 145.200 147.600 146.800 147.700 ;
        RECT 148.000 147.600 148.800 148.400 ;
        RECT 148.200 147.200 148.800 147.600 ;
        RECT 146.800 146.800 147.600 147.000 ;
        RECT 145.200 146.200 147.600 146.800 ;
        RECT 148.200 146.400 149.000 147.200 ;
        RECT 145.200 142.200 146.000 146.200 ;
        RECT 149.600 145.800 150.200 149.200 ;
        RECT 151.000 149.200 153.600 149.800 ;
        RECT 151.000 148.600 151.600 149.200 ;
        RECT 150.800 147.800 151.600 148.600 ;
        RECT 161.200 149.000 162.000 154.600 ;
        RECT 163.800 154.400 168.000 155.200 ;
        RECT 172.400 155.000 173.200 159.800 ;
        RECT 175.600 155.000 176.400 159.800 ;
        RECT 163.800 154.000 164.400 154.400 ;
        RECT 162.800 153.200 164.400 154.000 ;
        RECT 167.400 153.800 173.200 154.400 ;
        RECT 165.400 153.200 166.800 153.800 ;
        RECT 165.400 153.000 171.600 153.200 ;
        RECT 166.200 152.600 171.600 153.000 ;
        RECT 170.800 152.400 171.600 152.600 ;
        RECT 172.600 153.000 173.200 153.800 ;
        RECT 173.800 153.600 176.400 154.400 ;
        RECT 178.800 153.600 179.600 159.800 ;
        RECT 180.400 157.000 181.200 159.800 ;
        RECT 182.000 157.000 182.800 159.800 ;
        RECT 183.600 157.000 184.400 159.800 ;
        RECT 182.000 154.400 186.200 155.200 ;
        RECT 186.800 154.400 187.600 159.800 ;
        RECT 190.000 155.200 190.800 159.800 ;
        RECT 190.000 154.600 192.600 155.200 ;
        RECT 186.800 153.600 189.400 154.400 ;
        RECT 180.400 153.000 181.200 153.200 ;
        RECT 172.600 152.400 181.200 153.000 ;
        RECT 183.600 153.000 184.400 153.200 ;
        RECT 192.000 153.000 192.600 154.600 ;
        RECT 183.600 152.400 192.600 153.000 ;
        RECT 192.000 150.600 192.600 152.400 ;
        RECT 193.200 154.300 194.000 159.800 ;
        RECT 197.200 154.300 198.000 154.400 ;
        RECT 193.200 153.700 198.000 154.300 ;
        RECT 193.200 152.000 194.000 153.700 ;
        RECT 197.200 153.600 198.000 153.700 ;
        RECT 197.200 152.400 197.800 153.600 ;
        RECT 198.600 152.400 199.400 159.800 ;
        RECT 204.400 152.800 205.200 159.800 ;
        RECT 193.200 151.200 194.200 152.000 ;
        RECT 196.400 151.800 197.800 152.400 ;
        RECT 198.400 151.800 199.400 152.400 ;
        RECT 204.200 151.800 205.200 152.800 ;
        RECT 207.600 152.400 208.400 159.800 ;
        RECT 205.800 151.800 208.400 152.400 ;
        RECT 209.800 152.600 210.600 159.800 ;
        RECT 209.800 151.800 211.600 152.600 ;
        RECT 196.400 151.600 197.200 151.800 ;
        RECT 162.600 150.000 186.000 150.600 ;
        RECT 192.000 150.000 192.800 150.600 ;
        RECT 162.600 149.800 163.400 150.000 ;
        RECT 167.600 149.600 168.400 150.000 ;
        RECT 185.200 149.400 186.000 150.000 ;
        RECT 154.000 148.200 155.600 148.400 ;
        RECT 152.200 147.600 155.600 148.200 ;
        RECT 161.200 148.200 170.000 149.000 ;
        RECT 170.600 148.600 172.600 149.400 ;
        RECT 176.400 148.600 179.600 149.400 ;
        RECT 152.200 147.200 152.800 147.600 ;
        RECT 150.800 146.600 152.800 147.200 ;
        RECT 153.400 146.800 154.200 147.000 ;
        RECT 150.800 146.400 152.400 146.600 ;
        RECT 153.400 146.200 155.600 146.800 ;
        RECT 149.600 142.200 151.200 145.800 ;
        RECT 154.800 142.200 155.600 146.200 ;
        RECT 161.200 142.200 162.000 148.200 ;
        RECT 163.600 146.800 166.600 147.600 ;
        RECT 165.800 146.200 166.600 146.800 ;
        RECT 171.800 146.200 172.600 148.600 ;
        RECT 174.000 146.800 174.800 148.400 ;
        RECT 179.200 147.800 180.000 148.000 ;
        RECT 175.600 147.200 180.000 147.800 ;
        RECT 175.600 147.000 176.400 147.200 ;
        RECT 182.000 146.400 182.800 149.200 ;
        RECT 187.800 148.600 191.600 149.400 ;
        RECT 187.800 147.400 188.600 148.600 ;
        RECT 192.200 148.000 192.800 150.000 ;
        RECT 175.600 146.200 176.400 146.400 ;
        RECT 165.800 145.400 168.400 146.200 ;
        RECT 171.800 145.600 176.400 146.200 ;
        RECT 177.200 145.600 178.800 146.400 ;
        RECT 181.800 145.600 182.800 146.400 ;
        RECT 186.800 146.800 188.600 147.400 ;
        RECT 191.600 147.400 192.800 148.000 ;
        RECT 186.800 146.200 187.600 146.800 ;
        RECT 167.600 142.200 168.400 145.400 ;
        RECT 185.200 145.400 187.600 146.200 ;
        RECT 169.200 142.200 170.000 145.000 ;
        RECT 170.800 142.200 171.600 145.000 ;
        RECT 172.400 142.200 173.200 145.000 ;
        RECT 175.600 142.200 176.400 145.000 ;
        RECT 178.800 142.200 179.600 145.000 ;
        RECT 180.400 142.200 181.200 145.000 ;
        RECT 182.000 142.200 182.800 145.000 ;
        RECT 183.600 142.200 184.400 145.000 ;
        RECT 185.200 142.200 186.000 145.400 ;
        RECT 191.600 142.200 192.400 147.400 ;
        RECT 193.400 146.800 194.200 151.200 ;
        RECT 198.400 148.400 199.000 151.800 ;
        RECT 199.600 150.300 200.400 150.400 ;
        RECT 201.200 150.300 202.000 150.400 ;
        RECT 199.600 149.700 202.000 150.300 ;
        RECT 199.600 148.800 200.400 149.700 ;
        RECT 201.200 149.600 202.000 149.700 ;
        RECT 204.200 148.400 204.800 151.800 ;
        RECT 205.800 149.800 206.400 151.800 ;
        RECT 205.400 149.000 206.400 149.800 ;
        RECT 196.400 147.600 199.000 148.400 ;
        RECT 201.200 148.300 202.000 148.400 ;
        RECT 204.200 148.300 205.200 148.400 ;
        RECT 201.200 148.200 205.200 148.300 ;
        RECT 200.400 147.700 205.200 148.200 ;
        RECT 200.400 147.600 202.000 147.700 ;
        RECT 204.200 147.600 205.200 147.700 ;
        RECT 193.200 146.000 194.200 146.800 ;
        RECT 196.600 146.200 197.200 147.600 ;
        RECT 200.400 147.200 201.200 147.600 ;
        RECT 198.200 146.200 201.800 146.600 ;
        RECT 204.200 146.400 204.800 147.600 ;
        RECT 205.800 147.400 206.400 149.000 ;
        RECT 207.400 149.600 208.400 150.400 ;
        RECT 209.200 149.600 210.000 151.200 ;
        RECT 210.800 150.300 211.400 151.800 ;
        RECT 214.000 151.600 214.800 153.200 ;
        RECT 214.000 150.300 214.800 150.400 ;
        RECT 210.800 149.700 214.800 150.300 ;
        RECT 207.400 148.800 208.200 149.600 ;
        RECT 210.800 148.400 211.400 149.700 ;
        RECT 214.000 149.600 214.800 149.700 ;
        RECT 210.800 147.600 211.600 148.400 ;
        RECT 205.800 146.800 208.400 147.400 ;
        RECT 193.200 142.200 194.000 146.000 ;
        RECT 196.400 142.200 197.200 146.200 ;
        RECT 198.000 146.000 202.000 146.200 ;
        RECT 198.000 142.200 198.800 146.000 ;
        RECT 201.200 142.200 202.000 146.000 ;
        RECT 204.200 145.600 205.200 146.400 ;
        RECT 204.400 142.200 205.200 145.600 ;
        RECT 207.600 142.200 208.400 146.800 ;
        RECT 210.800 144.400 211.400 147.600 ;
        RECT 212.400 144.800 213.200 146.400 ;
        RECT 215.600 146.200 216.400 159.800 ;
        RECT 221.400 152.400 222.200 159.800 ;
        RECT 226.800 156.400 227.600 159.800 ;
        RECT 226.600 155.800 227.600 156.400 ;
        RECT 226.600 155.200 227.200 155.800 ;
        RECT 230.000 155.200 230.800 159.800 ;
        RECT 233.200 157.000 234.000 159.800 ;
        RECT 234.800 157.000 235.600 159.800 ;
        RECT 225.200 154.600 227.200 155.200 ;
        RECT 222.800 153.600 224.400 154.400 ;
        RECT 223.000 152.400 223.600 153.600 ;
        RECT 221.400 151.800 222.400 152.400 ;
        RECT 223.000 151.800 224.400 152.400 ;
        RECT 220.400 148.800 221.200 150.400 ;
        RECT 221.800 148.400 222.400 151.800 ;
        RECT 223.600 151.600 224.400 151.800 ;
        RECT 225.200 149.000 226.000 154.600 ;
        RECT 227.800 154.400 232.000 155.200 ;
        RECT 236.400 155.000 237.200 159.800 ;
        RECT 239.600 155.000 240.400 159.800 ;
        RECT 227.800 154.000 228.400 154.400 ;
        RECT 226.800 153.200 228.400 154.000 ;
        RECT 231.400 153.800 237.200 154.400 ;
        RECT 229.400 153.200 230.800 153.800 ;
        RECT 229.400 153.000 235.600 153.200 ;
        RECT 230.200 152.600 235.600 153.000 ;
        RECT 234.800 152.400 235.600 152.600 ;
        RECT 236.600 153.000 237.200 153.800 ;
        RECT 237.800 153.600 240.400 154.400 ;
        RECT 242.800 153.600 243.600 159.800 ;
        RECT 244.400 157.000 245.200 159.800 ;
        RECT 246.000 157.000 246.800 159.800 ;
        RECT 247.600 157.000 248.400 159.800 ;
        RECT 246.000 154.400 250.200 155.200 ;
        RECT 250.800 154.400 251.600 159.800 ;
        RECT 254.000 155.200 254.800 159.800 ;
        RECT 254.000 154.600 256.600 155.200 ;
        RECT 250.800 153.600 253.400 154.400 ;
        RECT 244.400 153.000 245.200 153.200 ;
        RECT 236.600 152.400 245.200 153.000 ;
        RECT 247.600 153.000 248.400 153.200 ;
        RECT 256.000 153.000 256.600 154.600 ;
        RECT 247.600 152.400 256.600 153.000 ;
        RECT 256.000 150.600 256.600 152.400 ;
        RECT 257.200 152.000 258.000 159.800 ;
        RECT 257.200 151.200 258.200 152.000 ;
        RECT 260.400 151.600 261.200 153.200 ;
        RECT 226.600 150.000 250.000 150.600 ;
        RECT 256.000 150.000 256.800 150.600 ;
        RECT 226.600 149.800 227.400 150.000 ;
        RECT 231.600 149.600 232.400 150.000 ;
        RECT 238.000 149.600 238.800 150.000 ;
        RECT 249.200 149.400 250.000 150.000 ;
        RECT 217.200 146.800 218.000 148.400 ;
        RECT 218.800 148.200 219.600 148.400 ;
        RECT 218.800 147.600 220.400 148.200 ;
        RECT 221.800 147.600 224.400 148.400 ;
        RECT 225.200 148.200 234.000 149.000 ;
        RECT 234.600 148.600 236.600 149.400 ;
        RECT 240.400 148.600 243.600 149.400 ;
        RECT 219.600 147.200 220.400 147.600 ;
        RECT 219.000 146.200 222.600 146.600 ;
        RECT 223.600 146.200 224.200 147.600 ;
        RECT 214.600 145.600 216.400 146.200 ;
        RECT 218.800 146.000 222.800 146.200 ;
        RECT 214.600 144.400 215.400 145.600 ;
        RECT 210.800 142.200 211.600 144.400 ;
        RECT 214.600 143.600 216.400 144.400 ;
        RECT 214.600 142.200 215.400 143.600 ;
        RECT 218.800 142.200 219.600 146.000 ;
        RECT 222.000 142.200 222.800 146.000 ;
        RECT 223.600 142.200 224.400 146.200 ;
        RECT 225.200 142.200 226.000 148.200 ;
        RECT 227.600 146.800 230.600 147.600 ;
        RECT 229.800 146.200 230.600 146.800 ;
        RECT 235.800 146.200 236.600 148.600 ;
        RECT 238.000 146.800 238.800 148.400 ;
        RECT 243.200 147.800 244.000 148.000 ;
        RECT 239.600 147.200 244.000 147.800 ;
        RECT 239.600 147.000 240.400 147.200 ;
        RECT 246.000 146.400 246.800 149.200 ;
        RECT 251.800 148.600 255.600 149.400 ;
        RECT 251.800 147.400 252.600 148.600 ;
        RECT 256.200 148.000 256.800 150.000 ;
        RECT 239.600 146.200 240.400 146.400 ;
        RECT 229.800 145.400 232.400 146.200 ;
        RECT 235.800 145.600 240.400 146.200 ;
        RECT 241.200 145.600 242.800 146.400 ;
        RECT 245.800 145.600 246.800 146.400 ;
        RECT 250.800 146.800 252.600 147.400 ;
        RECT 255.600 147.400 256.800 148.000 ;
        RECT 250.800 146.200 251.600 146.800 ;
        RECT 231.600 142.200 232.400 145.400 ;
        RECT 249.200 145.400 251.600 146.200 ;
        RECT 233.200 142.200 234.000 145.000 ;
        RECT 234.800 142.200 235.600 145.000 ;
        RECT 236.400 142.200 237.200 145.000 ;
        RECT 239.600 142.200 240.400 145.000 ;
        RECT 242.800 142.200 243.600 145.000 ;
        RECT 244.400 142.200 245.200 145.000 ;
        RECT 246.000 142.200 246.800 145.000 ;
        RECT 247.600 142.200 248.400 145.000 ;
        RECT 249.200 142.200 250.000 145.400 ;
        RECT 255.600 142.200 256.400 147.400 ;
        RECT 257.400 146.800 258.200 151.200 ;
        RECT 257.200 146.000 258.200 146.800 ;
        RECT 262.000 146.200 262.800 159.800 ;
        RECT 266.800 156.400 267.600 159.800 ;
        RECT 266.600 155.800 267.600 156.400 ;
        RECT 266.600 155.200 267.200 155.800 ;
        RECT 270.000 155.200 270.800 159.800 ;
        RECT 273.200 157.000 274.000 159.800 ;
        RECT 274.800 157.000 275.600 159.800 ;
        RECT 265.200 154.600 267.200 155.200 ;
        RECT 265.200 149.000 266.000 154.600 ;
        RECT 267.800 154.400 272.000 155.200 ;
        RECT 276.400 155.000 277.200 159.800 ;
        RECT 279.600 155.000 280.400 159.800 ;
        RECT 267.800 154.000 268.400 154.400 ;
        RECT 266.800 153.200 268.400 154.000 ;
        RECT 271.400 153.800 277.200 154.400 ;
        RECT 269.400 153.200 270.800 153.800 ;
        RECT 269.400 153.000 275.600 153.200 ;
        RECT 270.200 152.600 275.600 153.000 ;
        RECT 274.800 152.400 275.600 152.600 ;
        RECT 276.600 153.000 277.200 153.800 ;
        RECT 277.800 153.600 280.400 154.400 ;
        RECT 282.800 153.600 283.600 159.800 ;
        RECT 284.400 157.000 285.200 159.800 ;
        RECT 286.000 157.000 286.800 159.800 ;
        RECT 287.600 157.000 288.400 159.800 ;
        RECT 286.000 154.400 290.200 155.200 ;
        RECT 290.800 154.400 291.600 159.800 ;
        RECT 294.000 155.200 294.800 159.800 ;
        RECT 294.000 154.600 296.600 155.200 ;
        RECT 290.800 153.600 293.400 154.400 ;
        RECT 284.400 153.000 285.200 153.200 ;
        RECT 276.600 152.400 285.200 153.000 ;
        RECT 287.600 153.000 288.400 153.200 ;
        RECT 296.000 153.000 296.600 154.600 ;
        RECT 287.600 152.400 296.600 153.000 ;
        RECT 296.000 150.600 296.600 152.400 ;
        RECT 297.200 154.300 298.000 159.800 ;
        RECT 298.800 154.300 299.600 154.400 ;
        RECT 297.200 153.700 299.600 154.300 ;
        RECT 297.200 152.000 298.000 153.700 ;
        RECT 298.800 153.600 299.600 153.700 ;
        RECT 297.200 151.200 298.200 152.000 ;
        RECT 266.600 150.000 290.000 150.600 ;
        RECT 296.000 150.000 296.800 150.600 ;
        RECT 266.600 149.800 267.600 150.000 ;
        RECT 266.800 149.600 267.600 149.800 ;
        RECT 271.600 149.600 272.400 150.000 ;
        RECT 289.200 149.400 290.000 150.000 ;
        RECT 263.600 146.800 264.400 148.400 ;
        RECT 265.200 148.200 274.000 149.000 ;
        RECT 274.600 148.600 276.600 149.400 ;
        RECT 280.400 148.600 283.600 149.400 ;
        RECT 257.200 142.200 258.000 146.000 ;
        RECT 261.000 145.600 262.800 146.200 ;
        RECT 261.000 144.400 261.800 145.600 ;
        RECT 261.000 143.600 262.800 144.400 ;
        RECT 261.000 142.200 261.800 143.600 ;
        RECT 265.200 142.200 266.000 148.200 ;
        RECT 267.600 146.800 270.600 147.600 ;
        RECT 269.800 146.200 270.600 146.800 ;
        RECT 275.800 146.200 276.600 148.600 ;
        RECT 278.000 146.800 278.800 148.400 ;
        RECT 283.200 147.800 284.000 148.000 ;
        RECT 279.600 147.200 284.000 147.800 ;
        RECT 279.600 147.000 280.400 147.200 ;
        RECT 286.000 146.400 286.800 149.200 ;
        RECT 291.800 148.600 295.600 149.400 ;
        RECT 291.800 147.400 292.600 148.600 ;
        RECT 296.200 148.000 296.800 150.000 ;
        RECT 279.600 146.200 280.400 146.400 ;
        RECT 269.800 145.400 272.400 146.200 ;
        RECT 275.800 145.600 280.400 146.200 ;
        RECT 281.200 145.600 282.800 146.400 ;
        RECT 285.800 145.600 286.800 146.400 ;
        RECT 290.800 146.800 292.600 147.400 ;
        RECT 295.600 147.400 296.800 148.000 ;
        RECT 290.800 146.200 291.600 146.800 ;
        RECT 271.600 142.200 272.400 145.400 ;
        RECT 289.200 145.400 291.600 146.200 ;
        RECT 273.200 142.200 274.000 145.000 ;
        RECT 274.800 142.200 275.600 145.000 ;
        RECT 276.400 142.200 277.200 145.000 ;
        RECT 279.600 142.200 280.400 145.000 ;
        RECT 282.800 142.200 283.600 145.000 ;
        RECT 284.400 142.200 285.200 145.000 ;
        RECT 286.000 142.200 286.800 145.000 ;
        RECT 287.600 142.200 288.400 145.000 ;
        RECT 289.200 142.200 290.000 145.400 ;
        RECT 295.600 142.200 296.400 147.400 ;
        RECT 297.400 146.800 298.200 151.200 ;
        RECT 298.800 148.300 299.600 148.400 ;
        RECT 300.400 148.300 301.200 159.800 ;
        RECT 311.000 152.400 311.800 159.800 ;
        RECT 312.400 153.600 313.200 154.400 ;
        RECT 312.600 152.400 313.200 153.600 ;
        RECT 311.000 151.800 312.000 152.400 ;
        RECT 312.600 152.300 314.000 152.400 ;
        RECT 314.800 152.300 315.600 152.400 ;
        RECT 312.600 151.800 315.600 152.300 ;
        RECT 310.000 148.800 310.800 150.400 ;
        RECT 311.400 148.400 312.000 151.800 ;
        RECT 313.200 151.700 315.600 151.800 ;
        RECT 313.200 151.600 314.000 151.700 ;
        RECT 314.800 151.600 315.600 151.700 ;
        RECT 308.400 148.300 309.200 148.400 ;
        RECT 298.800 147.700 301.200 148.300 ;
        RECT 298.800 147.600 299.600 147.700 ;
        RECT 297.200 146.000 298.200 146.800 ;
        RECT 297.200 142.200 298.000 146.000 ;
        RECT 300.400 142.200 301.200 147.700 ;
        RECT 302.100 148.200 309.200 148.300 ;
        RECT 311.400 148.300 314.000 148.400 ;
        RECT 314.800 148.300 315.600 148.400 ;
        RECT 302.100 147.700 310.000 148.200 ;
        RECT 302.100 146.400 302.700 147.700 ;
        RECT 308.400 147.600 310.000 147.700 ;
        RECT 311.400 147.700 315.600 148.300 ;
        RECT 311.400 147.600 314.000 147.700 ;
        RECT 309.200 147.200 310.000 147.600 ;
        RECT 302.000 144.800 302.800 146.400 ;
        RECT 308.600 146.200 312.200 146.600 ;
        RECT 313.200 146.200 313.800 147.600 ;
        RECT 314.800 146.800 315.600 147.700 ;
        RECT 316.400 146.200 317.200 159.800 ;
        RECT 321.200 156.400 322.000 159.800 ;
        RECT 321.000 155.800 322.000 156.400 ;
        RECT 321.000 155.200 321.600 155.800 ;
        RECT 324.400 155.200 325.200 159.800 ;
        RECT 327.600 157.000 328.400 159.800 ;
        RECT 329.200 157.000 330.000 159.800 ;
        RECT 319.600 154.600 321.600 155.200 ;
        RECT 318.000 151.600 318.800 153.200 ;
        RECT 319.600 149.000 320.400 154.600 ;
        RECT 322.200 154.400 326.400 155.200 ;
        RECT 330.800 155.000 331.600 159.800 ;
        RECT 334.000 155.000 334.800 159.800 ;
        RECT 322.200 154.000 322.800 154.400 ;
        RECT 321.200 153.200 322.800 154.000 ;
        RECT 325.800 153.800 331.600 154.400 ;
        RECT 323.800 153.200 325.200 153.800 ;
        RECT 323.800 153.000 330.000 153.200 ;
        RECT 324.600 152.600 330.000 153.000 ;
        RECT 329.200 152.400 330.000 152.600 ;
        RECT 331.000 153.000 331.600 153.800 ;
        RECT 332.200 153.600 334.800 154.400 ;
        RECT 337.200 153.600 338.000 159.800 ;
        RECT 338.800 157.000 339.600 159.800 ;
        RECT 340.400 157.000 341.200 159.800 ;
        RECT 342.000 157.000 342.800 159.800 ;
        RECT 340.400 154.400 344.600 155.200 ;
        RECT 345.200 154.400 346.000 159.800 ;
        RECT 348.400 155.200 349.200 159.800 ;
        RECT 348.400 154.600 351.000 155.200 ;
        RECT 345.200 153.600 347.800 154.400 ;
        RECT 338.800 153.000 339.600 153.200 ;
        RECT 331.000 152.400 339.600 153.000 ;
        RECT 342.000 153.000 342.800 153.200 ;
        RECT 350.400 153.000 351.000 154.600 ;
        RECT 342.000 152.400 351.000 153.000 ;
        RECT 350.400 150.600 351.000 152.400 ;
        RECT 351.600 152.000 352.400 159.800 ;
        RECT 351.600 151.200 352.600 152.000 ;
        RECT 354.800 151.600 355.600 153.200 ;
        RECT 321.000 150.000 344.400 150.600 ;
        RECT 350.400 150.000 351.200 150.600 ;
        RECT 321.000 149.800 321.800 150.000 ;
        RECT 326.000 149.600 326.800 150.000 ;
        RECT 332.400 149.600 333.200 150.000 ;
        RECT 343.600 149.400 344.400 150.000 ;
        RECT 319.600 148.200 328.400 149.000 ;
        RECT 329.000 148.600 331.000 149.400 ;
        RECT 334.800 148.600 338.000 149.400 ;
        RECT 308.400 146.000 312.400 146.200 ;
        RECT 308.400 142.200 309.200 146.000 ;
        RECT 311.600 142.200 312.400 146.000 ;
        RECT 313.200 142.200 314.000 146.200 ;
        RECT 316.400 145.600 318.200 146.200 ;
        RECT 317.400 144.400 318.200 145.600 ;
        RECT 317.400 143.600 318.800 144.400 ;
        RECT 317.400 142.200 318.200 143.600 ;
        RECT 319.600 142.200 320.400 148.200 ;
        RECT 322.000 146.800 325.000 147.600 ;
        RECT 324.200 146.200 325.000 146.800 ;
        RECT 330.200 146.200 331.000 148.600 ;
        RECT 332.400 146.800 333.200 148.400 ;
        RECT 337.600 147.800 338.400 148.000 ;
        RECT 334.000 147.200 338.400 147.800 ;
        RECT 334.000 147.000 334.800 147.200 ;
        RECT 340.400 146.400 341.200 149.200 ;
        RECT 346.200 148.600 350.000 149.400 ;
        RECT 346.200 147.400 347.000 148.600 ;
        RECT 350.600 148.000 351.200 150.000 ;
        RECT 334.000 146.200 334.800 146.400 ;
        RECT 324.200 145.400 326.800 146.200 ;
        RECT 330.200 145.600 334.800 146.200 ;
        RECT 335.600 145.600 337.200 146.400 ;
        RECT 340.200 145.600 341.200 146.400 ;
        RECT 345.200 146.800 347.000 147.400 ;
        RECT 350.000 147.400 351.200 148.000 ;
        RECT 345.200 146.200 346.000 146.800 ;
        RECT 326.000 142.200 326.800 145.400 ;
        RECT 343.600 145.400 346.000 146.200 ;
        RECT 327.600 142.200 328.400 145.000 ;
        RECT 329.200 142.200 330.000 145.000 ;
        RECT 330.800 142.200 331.600 145.000 ;
        RECT 334.000 142.200 334.800 145.000 ;
        RECT 337.200 142.200 338.000 145.000 ;
        RECT 338.800 142.200 339.600 145.000 ;
        RECT 340.400 142.200 341.200 145.000 ;
        RECT 342.000 142.200 342.800 145.000 ;
        RECT 343.600 142.200 344.400 145.400 ;
        RECT 350.000 142.200 350.800 147.400 ;
        RECT 351.800 146.800 352.600 151.200 ;
        RECT 354.800 148.300 355.600 148.400 ;
        RECT 356.400 148.300 357.200 159.800 ;
        RECT 358.000 154.300 358.800 154.400 ;
        RECT 360.400 154.300 361.200 154.400 ;
        RECT 358.000 153.700 361.200 154.300 ;
        RECT 358.000 153.600 358.800 153.700 ;
        RECT 360.400 153.600 361.200 153.700 ;
        RECT 360.400 152.400 361.000 153.600 ;
        RECT 361.800 152.400 362.600 159.800 ;
        RECT 359.600 151.800 361.000 152.400 ;
        RECT 361.600 151.800 362.600 152.400 ;
        RECT 359.600 151.600 360.400 151.800 ;
        RECT 361.600 148.400 362.200 151.800 ;
        RECT 362.800 148.800 363.600 150.400 ;
        RECT 354.800 147.700 357.200 148.300 ;
        RECT 354.800 147.600 355.600 147.700 ;
        RECT 351.600 146.000 352.600 146.800 ;
        RECT 356.400 146.200 357.200 147.700 ;
        RECT 358.000 148.300 358.800 148.400 ;
        RECT 359.600 148.300 362.200 148.400 ;
        RECT 358.000 147.700 362.200 148.300 ;
        RECT 364.400 148.200 365.200 148.400 ;
        RECT 358.000 146.800 358.800 147.700 ;
        RECT 359.600 147.600 362.200 147.700 ;
        RECT 363.600 147.600 365.200 148.200 ;
        RECT 359.800 146.200 360.400 147.600 ;
        RECT 363.600 147.200 364.400 147.600 ;
        RECT 366.000 146.800 366.800 148.400 ;
        RECT 361.400 146.200 365.000 146.600 ;
        RECT 367.600 146.200 368.400 159.800 ;
        RECT 373.000 158.400 373.800 159.800 ;
        RECT 379.400 158.400 380.200 159.800 ;
        RECT 373.000 157.600 374.800 158.400 ;
        RECT 379.400 157.600 381.200 158.400 ;
        RECT 371.600 153.600 372.400 154.400 ;
        RECT 369.200 151.600 370.000 153.200 ;
        RECT 371.600 152.400 372.200 153.600 ;
        RECT 373.000 152.400 373.800 157.600 ;
        RECT 378.000 153.600 378.800 154.400 ;
        RECT 378.000 152.400 378.600 153.600 ;
        RECT 379.400 152.400 380.200 157.600 ;
        RECT 386.200 152.400 387.000 159.800 ;
        RECT 387.600 153.600 388.400 154.400 ;
        RECT 387.800 152.400 388.400 153.600 ;
        RECT 390.800 153.600 391.600 154.400 ;
        RECT 390.800 152.400 391.400 153.600 ;
        RECT 392.200 152.400 393.000 159.800 ;
        RECT 396.400 155.800 397.200 159.800 ;
        RECT 396.600 155.600 397.200 155.800 ;
        RECT 399.600 155.800 400.400 159.800 ;
        RECT 399.600 155.600 400.200 155.800 ;
        RECT 402.800 155.600 403.600 159.800 ;
        RECT 406.000 155.800 406.800 159.800 ;
        RECT 406.000 155.600 406.600 155.800 ;
        RECT 396.600 155.000 400.200 155.600 ;
        RECT 403.000 155.000 406.600 155.600 ;
        RECT 396.600 152.400 397.200 155.000 ;
        RECT 398.000 152.800 398.800 154.400 ;
        RECT 403.000 152.400 403.600 155.000 ;
        RECT 404.400 152.800 405.200 154.400 ;
        RECT 411.800 152.400 412.600 159.800 ;
        RECT 413.200 153.600 414.000 154.400 ;
        RECT 413.400 152.400 414.000 153.600 ;
        RECT 416.400 153.600 417.200 154.400 ;
        RECT 416.400 152.400 417.000 153.600 ;
        RECT 417.800 152.400 418.600 159.800 ;
        RECT 425.800 152.800 426.600 159.800 ;
        RECT 430.000 155.000 430.800 159.000 ;
        RECT 370.800 151.800 372.200 152.400 ;
        RECT 372.800 151.800 373.800 152.400 ;
        RECT 377.200 151.800 378.600 152.400 ;
        RECT 379.200 151.800 380.200 152.400 ;
        RECT 370.800 151.600 371.600 151.800 ;
        RECT 372.800 148.400 373.400 151.800 ;
        RECT 377.200 151.600 378.000 151.800 ;
        RECT 374.000 148.800 374.800 150.400 ;
        RECT 379.200 148.400 379.800 151.800 ;
        RECT 385.200 151.600 387.200 152.400 ;
        RECT 387.800 151.800 389.200 152.400 ;
        RECT 388.400 151.600 389.200 151.800 ;
        RECT 390.000 151.800 391.400 152.400 ;
        RECT 392.000 151.800 393.000 152.400 ;
        RECT 390.000 151.600 390.800 151.800 ;
        RECT 380.400 148.800 381.200 150.400 ;
        RECT 385.200 148.800 386.000 150.400 ;
        RECT 386.600 148.400 387.200 151.600 ;
        RECT 392.000 148.400 392.600 151.800 ;
        RECT 396.400 151.600 397.200 152.400 ;
        RECT 393.200 148.800 394.000 150.400 ;
        RECT 396.600 148.400 397.200 151.600 ;
        RECT 401.200 150.800 402.000 152.400 ;
        RECT 402.800 151.600 403.600 152.400 ;
        RECT 398.800 149.600 400.400 150.400 ;
        RECT 403.000 148.400 403.600 151.600 ;
        RECT 407.600 150.800 408.400 152.400 ;
        RECT 411.800 151.800 412.800 152.400 ;
        RECT 413.400 151.800 414.800 152.400 ;
        RECT 405.200 149.600 406.800 150.400 ;
        RECT 410.800 148.800 411.600 150.400 ;
        RECT 412.200 150.300 412.800 151.800 ;
        RECT 414.000 151.600 414.800 151.800 ;
        RECT 415.600 151.800 417.000 152.400 ;
        RECT 417.600 151.800 418.600 152.400 ;
        RECT 425.000 152.200 426.600 152.800 ;
        RECT 415.600 151.600 416.400 151.800 ;
        RECT 415.700 150.300 416.300 151.600 ;
        RECT 412.200 149.700 416.300 150.300 ;
        RECT 412.200 148.400 412.800 149.700 ;
        RECT 417.600 148.400 418.200 151.800 ;
        RECT 418.800 150.300 419.600 150.400 ;
        RECT 418.800 149.700 422.700 150.300 ;
        RECT 418.800 148.800 419.600 149.700 ;
        RECT 370.800 147.600 373.400 148.400 ;
        RECT 375.600 148.200 376.400 148.400 ;
        RECT 374.800 147.600 376.400 148.200 ;
        RECT 377.200 147.600 379.800 148.400 ;
        RECT 382.000 148.200 382.800 148.400 ;
        RECT 381.200 147.600 382.800 148.200 ;
        RECT 383.600 148.200 384.400 148.400 ;
        RECT 383.600 147.600 385.200 148.200 ;
        RECT 386.600 147.600 389.200 148.400 ;
        RECT 390.000 147.600 392.600 148.400 ;
        RECT 394.800 148.200 395.600 148.400 ;
        RECT 394.000 147.600 395.600 148.200 ;
        RECT 396.600 148.200 398.200 148.400 ;
        RECT 403.000 148.200 404.600 148.400 ;
        RECT 409.200 148.200 410.000 148.400 ;
        RECT 396.600 147.800 398.400 148.200 ;
        RECT 403.000 147.800 404.800 148.200 ;
        RECT 371.000 146.200 371.600 147.600 ;
        RECT 374.800 147.200 375.600 147.600 ;
        RECT 372.600 146.200 376.200 146.600 ;
        RECT 377.400 146.200 378.000 147.600 ;
        RECT 381.200 147.200 382.000 147.600 ;
        RECT 384.400 147.200 385.200 147.600 ;
        RECT 379.000 146.200 382.600 146.600 ;
        RECT 383.800 146.200 387.400 146.600 ;
        RECT 388.400 146.200 389.000 147.600 ;
        RECT 390.200 146.200 390.800 147.600 ;
        RECT 394.000 147.200 394.800 147.600 ;
        RECT 391.800 146.200 395.400 146.600 ;
        RECT 351.600 142.200 352.400 146.000 ;
        RECT 355.400 145.600 357.200 146.200 ;
        RECT 355.400 142.200 356.200 145.600 ;
        RECT 359.600 142.200 360.400 146.200 ;
        RECT 361.200 146.000 365.200 146.200 ;
        RECT 361.200 142.200 362.000 146.000 ;
        RECT 364.400 142.200 365.200 146.000 ;
        RECT 367.600 145.600 369.400 146.200 ;
        RECT 368.600 144.400 369.400 145.600 ;
        RECT 368.600 143.600 370.000 144.400 ;
        RECT 368.600 142.200 369.400 143.600 ;
        RECT 370.800 142.200 371.600 146.200 ;
        RECT 372.400 146.000 376.400 146.200 ;
        RECT 372.400 142.200 373.200 146.000 ;
        RECT 375.600 142.200 376.400 146.000 ;
        RECT 377.200 142.200 378.000 146.200 ;
        RECT 378.800 146.000 382.800 146.200 ;
        RECT 378.800 142.200 379.600 146.000 ;
        RECT 382.000 142.200 382.800 146.000 ;
        RECT 383.600 146.000 387.600 146.200 ;
        RECT 383.600 142.200 384.400 146.000 ;
        RECT 386.800 142.200 387.600 146.000 ;
        RECT 388.400 142.200 389.200 146.200 ;
        RECT 390.000 142.200 390.800 146.200 ;
        RECT 391.600 146.000 395.600 146.200 ;
        RECT 391.600 142.200 392.400 146.000 ;
        RECT 394.800 142.200 395.600 146.000 ;
        RECT 397.600 142.200 398.400 147.800 ;
        RECT 404.000 142.200 404.800 147.800 ;
        RECT 409.200 147.600 410.800 148.200 ;
        RECT 412.200 147.600 414.800 148.400 ;
        RECT 415.600 147.600 418.200 148.400 ;
        RECT 420.400 148.200 421.200 148.400 ;
        RECT 419.600 147.600 421.200 148.200 ;
        RECT 422.100 148.300 422.700 149.700 ;
        RECT 423.600 149.600 424.400 151.200 ;
        RECT 425.000 148.400 425.600 152.200 ;
        RECT 430.200 151.600 430.800 155.000 ;
        RECT 432.400 153.600 433.200 154.400 ;
        RECT 432.400 152.400 433.000 153.600 ;
        RECT 433.800 152.400 434.600 159.800 ;
        RECT 431.600 151.800 433.000 152.400 ;
        RECT 433.600 151.800 434.600 152.400 ;
        RECT 431.600 151.600 432.400 151.800 ;
        RECT 427.000 151.000 430.800 151.600 ;
        RECT 427.000 149.000 427.600 151.000 ;
        RECT 423.600 148.300 425.600 148.400 ;
        RECT 422.100 147.700 425.600 148.300 ;
        RECT 426.200 148.200 427.600 149.000 ;
        RECT 428.400 148.800 429.200 150.400 ;
        RECT 430.000 148.800 430.800 150.400 ;
        RECT 433.600 148.400 434.200 151.800 ;
        RECT 434.800 148.800 435.600 150.400 ;
        RECT 423.600 147.600 425.600 147.700 ;
        RECT 410.000 147.200 410.800 147.600 ;
        RECT 409.400 146.200 413.000 146.600 ;
        RECT 414.000 146.200 414.600 147.600 ;
        RECT 415.800 146.200 416.400 147.600 ;
        RECT 419.600 147.200 420.400 147.600 ;
        RECT 425.000 147.000 425.600 147.600 ;
        RECT 426.600 147.800 427.600 148.200 ;
        RECT 426.600 147.200 430.800 147.800 ;
        RECT 431.600 147.600 434.200 148.400 ;
        RECT 436.400 148.300 437.200 148.400 ;
        RECT 438.000 148.300 438.800 159.800 ;
        RECT 441.200 155.000 442.000 159.000 ;
        RECT 445.400 158.400 446.200 159.800 ;
        RECT 445.400 157.600 446.800 158.400 ;
        RECT 441.200 151.600 441.800 155.000 ;
        RECT 445.400 152.800 446.200 157.600 ;
        RECT 445.400 152.200 447.000 152.800 ;
        RECT 441.200 151.000 445.000 151.600 ;
        RECT 441.200 148.800 442.000 150.400 ;
        RECT 442.800 148.800 443.600 150.400 ;
        RECT 444.400 149.000 445.000 151.000 ;
        RECT 436.400 148.200 438.800 148.300 ;
        RECT 435.600 147.700 438.800 148.200 ;
        RECT 444.400 148.200 445.800 149.000 ;
        RECT 446.400 148.400 447.000 152.200 ;
        RECT 450.800 151.600 451.600 153.200 ;
        RECT 447.600 149.600 448.400 151.200 ;
        RECT 449.200 150.300 450.000 150.400 ;
        RECT 452.400 150.300 453.200 159.800 ;
        RECT 449.200 149.700 453.200 150.300 ;
        RECT 449.200 149.600 450.000 149.700 ;
        RECT 444.400 147.800 445.400 148.200 ;
        RECT 435.600 147.600 437.200 147.700 ;
        RECT 425.000 146.600 425.800 147.000 ;
        RECT 417.400 146.200 421.000 146.600 ;
        RECT 409.200 146.000 413.200 146.200 ;
        RECT 409.200 142.200 410.000 146.000 ;
        RECT 412.400 142.200 413.200 146.000 ;
        RECT 414.000 142.200 414.800 146.200 ;
        RECT 415.600 142.200 416.400 146.200 ;
        RECT 417.200 146.000 421.200 146.200 ;
        RECT 425.000 146.000 426.600 146.600 ;
        RECT 417.200 142.200 418.000 146.000 ;
        RECT 420.400 142.200 421.200 146.000 ;
        RECT 425.800 143.000 426.600 146.000 ;
        RECT 430.200 145.000 430.800 147.200 ;
        RECT 431.800 146.200 432.400 147.600 ;
        RECT 435.600 147.200 436.400 147.600 ;
        RECT 433.400 146.200 437.000 146.600 ;
        RECT 430.000 143.000 430.800 145.000 ;
        RECT 431.600 142.200 432.400 146.200 ;
        RECT 433.200 146.000 437.200 146.200 ;
        RECT 433.200 142.200 434.000 146.000 ;
        RECT 436.400 142.200 437.200 146.000 ;
        RECT 438.000 142.200 438.800 147.700 ;
        RECT 441.200 147.200 445.400 147.800 ;
        RECT 446.400 147.600 448.400 148.400 ;
        RECT 439.600 144.800 440.400 146.400 ;
        RECT 441.200 145.000 441.800 147.200 ;
        RECT 446.400 147.000 447.000 147.600 ;
        RECT 446.200 146.600 447.000 147.000 ;
        RECT 445.400 146.000 447.000 146.600 ;
        RECT 452.400 146.200 453.200 149.700 ;
        RECT 460.400 151.200 461.200 159.800 ;
        RECT 464.600 155.800 465.800 159.800 ;
        RECT 469.200 155.800 470.000 159.800 ;
        RECT 473.600 156.400 474.400 159.800 ;
        RECT 473.600 155.800 475.600 156.400 ;
        RECT 465.200 155.000 466.000 155.800 ;
        RECT 469.400 155.200 470.000 155.800 ;
        RECT 468.600 154.600 472.200 155.200 ;
        RECT 474.800 155.000 475.600 155.800 ;
        RECT 468.600 154.400 469.400 154.600 ;
        RECT 471.400 154.400 472.200 154.600 ;
        RECT 464.400 153.200 465.800 154.000 ;
        RECT 465.200 152.200 465.800 153.200 ;
        RECT 467.400 153.000 469.600 153.600 ;
        RECT 467.400 152.800 468.200 153.000 ;
        RECT 465.200 151.600 467.600 152.200 ;
        RECT 460.400 150.600 464.600 151.200 ;
        RECT 454.000 146.800 454.800 148.400 ;
        RECT 460.400 147.200 461.200 150.600 ;
        RECT 463.800 150.400 464.600 150.600 ;
        RECT 462.200 149.800 463.000 150.000 ;
        RECT 462.200 149.200 466.000 149.800 ;
        RECT 465.200 149.000 466.000 149.200 ;
        RECT 467.000 148.400 467.600 151.600 ;
        RECT 469.000 151.800 469.600 153.000 ;
        RECT 470.200 153.000 471.000 153.200 ;
        RECT 474.800 153.000 475.600 153.200 ;
        RECT 470.200 152.400 475.600 153.000 ;
        RECT 469.000 151.400 473.800 151.800 ;
        RECT 478.000 151.400 478.800 159.800 ;
        RECT 469.000 151.200 478.800 151.400 ;
        RECT 473.000 151.000 478.800 151.200 ;
        RECT 473.200 150.800 478.800 151.000 ;
        RECT 471.600 150.200 472.400 150.400 ;
        RECT 471.600 149.600 476.600 150.200 ;
        RECT 475.800 149.400 476.600 149.600 ;
        RECT 474.200 148.400 475.000 148.600 ;
        RECT 467.000 147.800 478.000 148.400 ;
        RECT 467.400 147.600 468.200 147.800 ;
        RECT 441.200 143.000 442.000 145.000 ;
        RECT 445.400 143.000 446.200 146.000 ;
        RECT 451.400 145.600 453.200 146.200 ;
        RECT 460.400 146.600 464.200 147.200 ;
        RECT 451.400 142.200 452.200 145.600 ;
        RECT 460.400 142.200 461.200 146.600 ;
        RECT 463.400 146.400 464.200 146.600 ;
        RECT 473.200 145.600 473.800 147.800 ;
        RECT 476.400 147.600 478.000 147.800 ;
        RECT 471.400 145.400 472.200 145.600 ;
        RECT 465.200 144.200 466.000 145.000 ;
        RECT 469.400 144.800 472.200 145.400 ;
        RECT 473.200 144.800 474.000 145.600 ;
        RECT 469.400 144.200 470.000 144.800 ;
        RECT 474.800 144.200 475.600 145.000 ;
        RECT 464.600 143.600 466.000 144.200 ;
        RECT 464.600 142.200 465.800 143.600 ;
        RECT 469.200 142.200 470.000 144.200 ;
        RECT 473.600 143.600 475.600 144.200 ;
        RECT 473.600 142.200 474.400 143.600 ;
        RECT 478.000 142.200 478.800 147.000 ;
        RECT 479.600 142.200 480.400 159.800 ;
        RECT 482.800 155.000 483.600 159.000 ;
        RECT 482.800 151.600 483.400 155.000 ;
        RECT 487.000 154.400 487.800 159.800 ;
        RECT 487.000 153.600 488.400 154.400 ;
        RECT 487.000 152.800 487.800 153.600 ;
        RECT 487.000 152.200 488.600 152.800 ;
        RECT 482.800 151.000 486.600 151.600 ;
        RECT 482.800 148.800 483.600 150.400 ;
        RECT 484.400 148.800 485.200 150.400 ;
        RECT 486.000 149.000 486.600 151.000 ;
        RECT 486.000 148.200 487.400 149.000 ;
        RECT 488.000 148.400 488.600 152.200 ;
        RECT 489.200 149.600 490.000 151.200 ;
        RECT 494.000 150.300 494.800 159.800 ;
        RECT 498.000 153.600 498.800 154.400 ;
        RECT 495.600 151.600 496.400 153.200 ;
        RECT 498.000 152.400 498.600 153.600 ;
        RECT 499.400 152.400 500.200 159.800 ;
        RECT 497.200 151.800 498.600 152.400 ;
        RECT 499.200 151.800 500.200 152.400 ;
        RECT 506.200 152.400 507.000 159.800 ;
        RECT 507.600 153.600 508.400 154.400 ;
        RECT 507.800 152.400 508.400 153.600 ;
        RECT 510.800 153.600 511.600 154.400 ;
        RECT 510.800 152.400 511.400 153.600 ;
        RECT 512.200 152.400 513.000 159.800 ;
        RECT 506.200 151.800 507.200 152.400 ;
        RECT 507.800 151.800 509.200 152.400 ;
        RECT 497.200 151.600 498.000 151.800 ;
        RECT 497.300 150.300 497.900 151.600 ;
        RECT 494.000 149.700 497.900 150.300 ;
        RECT 486.000 147.800 487.000 148.200 ;
        RECT 482.800 147.200 487.000 147.800 ;
        RECT 488.000 147.600 490.000 148.400 ;
        RECT 481.200 144.800 482.000 146.400 ;
        RECT 482.800 145.000 483.400 147.200 ;
        RECT 488.000 147.000 488.600 147.600 ;
        RECT 487.800 146.600 488.600 147.000 ;
        RECT 492.400 146.800 493.200 148.400 ;
        RECT 487.000 146.000 488.600 146.600 ;
        RECT 494.000 146.200 494.800 149.700 ;
        RECT 499.200 148.400 499.800 151.800 ;
        RECT 500.400 148.800 501.200 150.400 ;
        RECT 505.200 148.800 506.000 150.400 ;
        RECT 506.600 148.400 507.200 151.800 ;
        RECT 508.400 151.600 509.200 151.800 ;
        RECT 510.000 151.800 511.400 152.400 ;
        RECT 512.000 151.800 513.000 152.400 ;
        RECT 510.000 151.600 510.800 151.800 ;
        RECT 508.500 150.300 509.100 151.600 ;
        RECT 512.000 150.300 512.600 151.800 ;
        RECT 516.400 151.200 517.200 159.800 ;
        RECT 520.600 155.800 521.800 159.800 ;
        RECT 525.200 155.800 526.000 159.800 ;
        RECT 529.600 156.400 530.400 159.800 ;
        RECT 529.600 155.800 531.600 156.400 ;
        RECT 521.200 155.000 522.000 155.800 ;
        RECT 525.400 155.200 526.000 155.800 ;
        RECT 524.600 154.600 528.200 155.200 ;
        RECT 530.800 155.000 531.600 155.800 ;
        RECT 524.600 154.400 525.400 154.600 ;
        RECT 527.400 154.400 528.200 154.600 ;
        RECT 519.600 154.000 521.000 154.400 ;
        RECT 519.600 153.600 521.800 154.000 ;
        RECT 520.400 153.200 521.800 153.600 ;
        RECT 521.200 152.200 521.800 153.200 ;
        RECT 523.400 153.000 525.600 153.600 ;
        RECT 523.400 152.800 524.200 153.000 ;
        RECT 521.200 151.600 523.600 152.200 ;
        RECT 516.400 150.600 520.600 151.200 ;
        RECT 508.500 149.700 512.600 150.300 ;
        RECT 512.000 148.400 512.600 149.700 ;
        RECT 513.200 148.800 514.000 150.400 ;
        RECT 497.200 147.600 499.800 148.400 ;
        RECT 502.000 148.200 502.800 148.400 ;
        RECT 501.200 147.600 502.800 148.200 ;
        RECT 503.600 148.200 504.400 148.400 ;
        RECT 503.600 147.600 505.200 148.200 ;
        RECT 506.600 147.600 509.200 148.400 ;
        RECT 510.000 147.600 512.600 148.400 ;
        RECT 514.800 148.200 515.600 148.400 ;
        RECT 514.000 147.600 515.600 148.200 ;
        RECT 497.400 146.200 498.000 147.600 ;
        RECT 501.200 147.200 502.000 147.600 ;
        RECT 504.400 147.200 505.200 147.600 ;
        RECT 499.000 146.200 502.600 146.600 ;
        RECT 503.800 146.200 507.400 146.600 ;
        RECT 508.400 146.200 509.000 147.600 ;
        RECT 510.200 146.200 510.800 147.600 ;
        RECT 514.000 147.200 514.800 147.600 ;
        RECT 516.400 147.200 517.200 150.600 ;
        RECT 519.800 150.400 520.600 150.600 ;
        RECT 518.200 149.800 519.000 150.000 ;
        RECT 518.200 149.200 522.000 149.800 ;
        RECT 521.200 149.000 522.000 149.200 ;
        RECT 523.000 148.400 523.600 151.600 ;
        RECT 525.000 151.800 525.600 153.000 ;
        RECT 526.200 153.000 527.000 153.200 ;
        RECT 530.800 153.000 531.600 153.200 ;
        RECT 526.200 152.400 531.600 153.000 ;
        RECT 525.000 151.400 529.800 151.800 ;
        RECT 534.000 151.400 534.800 159.800 ;
        RECT 538.200 152.400 539.000 159.800 ;
        RECT 539.600 153.600 540.400 154.400 ;
        RECT 539.800 152.400 540.400 153.600 ;
        RECT 538.200 151.800 539.200 152.400 ;
        RECT 539.800 151.800 541.200 152.400 ;
        RECT 525.000 151.200 534.800 151.400 ;
        RECT 529.000 151.000 534.800 151.200 ;
        RECT 529.200 150.800 534.800 151.000 ;
        RECT 527.600 150.200 528.400 150.400 ;
        RECT 527.600 149.600 532.600 150.200 ;
        RECT 531.800 149.400 532.600 149.600 ;
        RECT 537.200 148.800 538.000 150.400 ;
        RECT 538.600 150.300 539.200 151.800 ;
        RECT 540.400 151.600 541.200 151.800 ;
        RECT 542.000 151.200 542.800 159.800 ;
        RECT 546.200 155.800 547.400 159.800 ;
        RECT 550.800 155.800 551.600 159.800 ;
        RECT 555.200 156.400 556.000 159.800 ;
        RECT 555.200 155.800 557.200 156.400 ;
        RECT 546.800 155.000 547.600 155.800 ;
        RECT 551.000 155.200 551.600 155.800 ;
        RECT 550.200 154.600 553.800 155.200 ;
        RECT 556.400 155.000 557.200 155.800 ;
        RECT 550.200 154.400 551.000 154.600 ;
        RECT 553.000 154.400 553.800 154.600 ;
        RECT 545.200 154.000 546.600 154.400 ;
        RECT 545.200 153.600 547.400 154.000 ;
        RECT 546.000 153.200 547.400 153.600 ;
        RECT 546.800 152.200 547.400 153.200 ;
        RECT 549.000 153.000 551.200 153.600 ;
        RECT 549.000 152.800 549.800 153.000 ;
        RECT 546.800 151.600 549.200 152.200 ;
        RECT 542.000 150.600 546.200 151.200 ;
        RECT 540.400 150.300 541.200 150.400 ;
        RECT 538.600 149.700 541.200 150.300 ;
        RECT 530.200 148.400 531.000 148.600 ;
        RECT 538.600 148.400 539.200 149.700 ;
        RECT 540.400 149.600 541.200 149.700 ;
        RECT 523.000 147.800 534.000 148.400 ;
        RECT 523.400 147.600 524.200 147.800 ;
        RECT 516.400 146.600 520.200 147.200 ;
        RECT 511.800 146.200 515.400 146.600 ;
        RECT 482.800 143.000 483.600 145.000 ;
        RECT 487.000 143.000 487.800 146.000 ;
        RECT 494.000 145.600 495.800 146.200 ;
        RECT 495.000 142.200 495.800 145.600 ;
        RECT 497.200 142.200 498.000 146.200 ;
        RECT 498.800 146.000 502.800 146.200 ;
        RECT 498.800 142.200 499.600 146.000 ;
        RECT 502.000 142.200 502.800 146.000 ;
        RECT 503.600 146.000 507.600 146.200 ;
        RECT 503.600 142.200 504.400 146.000 ;
        RECT 506.800 142.200 507.600 146.000 ;
        RECT 508.400 142.200 509.200 146.200 ;
        RECT 510.000 142.200 510.800 146.200 ;
        RECT 511.600 146.000 515.600 146.200 ;
        RECT 511.600 142.200 512.400 146.000 ;
        RECT 514.800 142.200 515.600 146.000 ;
        RECT 516.400 142.200 517.200 146.600 ;
        RECT 519.400 146.400 520.200 146.600 ;
        RECT 529.200 146.400 529.800 147.800 ;
        RECT 532.400 147.600 534.000 147.800 ;
        RECT 535.600 148.200 536.400 148.400 ;
        RECT 535.600 147.600 537.200 148.200 ;
        RECT 538.600 147.600 541.200 148.400 ;
        RECT 536.400 147.200 537.200 147.600 ;
        RECT 527.400 145.400 528.200 145.600 ;
        RECT 521.200 144.200 522.000 145.000 ;
        RECT 525.400 144.800 528.200 145.400 ;
        RECT 529.200 144.800 530.000 146.400 ;
        RECT 525.400 144.200 526.000 144.800 ;
        RECT 530.800 144.200 531.600 145.000 ;
        RECT 520.600 143.600 522.000 144.200 ;
        RECT 520.600 142.200 521.800 143.600 ;
        RECT 525.200 142.200 526.000 144.200 ;
        RECT 529.600 143.600 531.600 144.200 ;
        RECT 529.600 142.200 530.400 143.600 ;
        RECT 534.000 142.200 534.800 147.000 ;
        RECT 535.800 146.200 539.400 146.600 ;
        RECT 540.400 146.200 541.000 147.600 ;
        RECT 542.000 147.200 542.800 150.600 ;
        RECT 545.400 150.400 546.200 150.600 ;
        RECT 543.800 149.800 544.600 150.000 ;
        RECT 543.800 149.200 547.600 149.800 ;
        RECT 546.800 149.000 547.600 149.200 ;
        RECT 548.600 148.400 549.200 151.600 ;
        RECT 550.600 151.800 551.200 153.000 ;
        RECT 551.800 153.000 552.600 153.200 ;
        RECT 556.400 153.000 557.200 153.200 ;
        RECT 551.800 152.400 557.200 153.000 ;
        RECT 550.600 151.400 555.400 151.800 ;
        RECT 559.600 151.400 560.400 159.800 ;
        RECT 550.600 151.200 560.400 151.400 ;
        RECT 554.600 151.000 560.400 151.200 ;
        RECT 554.800 150.800 560.400 151.000 ;
        RECT 561.200 151.200 562.000 159.800 ;
        RECT 565.400 154.300 566.200 159.800 ;
        RECT 567.600 154.300 568.400 154.400 ;
        RECT 565.400 153.700 568.400 154.300 ;
        RECT 565.400 152.400 566.200 153.700 ;
        RECT 567.600 153.600 568.400 153.700 ;
        RECT 565.400 151.800 566.800 152.400 ;
        RECT 569.200 152.000 570.000 159.800 ;
        RECT 572.400 155.200 573.200 159.800 ;
        RECT 561.200 150.800 565.200 151.200 ;
        RECT 561.200 150.600 565.400 150.800 ;
        RECT 550.000 150.300 550.800 150.400 ;
        RECT 553.200 150.300 554.000 150.400 ;
        RECT 550.000 150.200 554.000 150.300 ;
        RECT 550.000 149.700 558.200 150.200 ;
        RECT 564.600 150.000 565.400 150.600 ;
        RECT 566.200 150.400 566.800 151.800 ;
        RECT 550.000 149.600 550.800 149.700 ;
        RECT 553.200 149.600 558.200 149.700 ;
        RECT 557.400 149.400 558.200 149.600 ;
        RECT 555.800 148.400 556.600 148.600 ;
        RECT 563.200 148.400 564.000 149.200 ;
        RECT 548.600 147.800 559.600 148.400 ;
        RECT 549.000 147.600 549.800 147.800 ;
        RECT 553.200 147.600 554.000 147.800 ;
        RECT 542.000 146.600 545.800 147.200 ;
        RECT 535.600 146.000 539.600 146.200 ;
        RECT 535.600 142.200 536.400 146.000 ;
        RECT 538.800 142.200 539.600 146.000 ;
        RECT 540.400 142.200 541.200 146.200 ;
        RECT 542.000 142.200 542.800 146.600 ;
        RECT 545.000 146.400 545.800 146.600 ;
        RECT 554.800 145.600 555.400 147.800 ;
        RECT 558.000 147.600 559.600 147.800 ;
        RECT 562.800 147.600 563.800 148.400 ;
        RECT 564.800 147.000 565.400 150.000 ;
        RECT 566.000 149.600 566.800 150.400 ;
        RECT 553.000 145.400 553.800 145.600 ;
        RECT 546.800 144.200 547.600 145.000 ;
        RECT 551.000 144.800 553.800 145.400 ;
        RECT 554.800 144.800 555.600 145.600 ;
        RECT 551.000 144.200 551.600 144.800 ;
        RECT 556.400 144.200 557.200 145.000 ;
        RECT 546.200 143.600 547.600 144.200 ;
        RECT 546.200 142.200 547.400 143.600 ;
        RECT 550.800 142.200 551.600 144.200 ;
        RECT 555.200 143.600 557.200 144.200 ;
        RECT 555.200 142.200 556.000 143.600 ;
        RECT 559.600 142.200 560.400 147.000 ;
        RECT 563.000 146.400 565.400 147.000 ;
        RECT 561.200 144.800 562.000 146.400 ;
        RECT 563.000 144.200 563.600 146.400 ;
        RECT 566.200 146.200 566.800 149.600 ;
        RECT 562.800 142.200 563.600 144.200 ;
        RECT 566.000 142.200 566.800 146.200 ;
        RECT 569.000 151.200 570.000 152.000 ;
        RECT 570.600 154.600 573.200 155.200 ;
        RECT 570.600 153.000 571.200 154.600 ;
        RECT 575.600 154.400 576.400 159.800 ;
        RECT 578.800 157.000 579.600 159.800 ;
        RECT 580.400 157.000 581.200 159.800 ;
        RECT 582.000 157.000 582.800 159.800 ;
        RECT 577.000 154.400 581.200 155.200 ;
        RECT 573.800 153.600 576.400 154.400 ;
        RECT 583.600 153.600 584.400 159.800 ;
        RECT 586.800 155.000 587.600 159.800 ;
        RECT 590.000 155.000 590.800 159.800 ;
        RECT 591.600 157.000 592.400 159.800 ;
        RECT 593.200 157.000 594.000 159.800 ;
        RECT 596.400 155.200 597.200 159.800 ;
        RECT 599.600 156.400 600.400 159.800 ;
        RECT 599.600 155.800 600.600 156.400 ;
        RECT 600.000 155.200 600.600 155.800 ;
        RECT 595.200 154.400 599.400 155.200 ;
        RECT 600.000 154.600 602.000 155.200 ;
        RECT 586.800 153.600 589.400 154.400 ;
        RECT 590.000 153.800 595.800 154.400 ;
        RECT 598.800 154.000 599.400 154.400 ;
        RECT 578.800 153.000 579.600 153.200 ;
        RECT 570.600 152.400 579.600 153.000 ;
        RECT 582.000 153.000 582.800 153.200 ;
        RECT 590.000 153.000 590.600 153.800 ;
        RECT 596.400 153.200 597.800 153.800 ;
        RECT 598.800 153.200 600.400 154.000 ;
        RECT 582.000 152.400 590.600 153.000 ;
        RECT 591.600 153.000 597.800 153.200 ;
        RECT 591.600 152.600 597.000 153.000 ;
        RECT 591.600 152.400 592.400 152.600 ;
        RECT 569.000 146.800 569.800 151.200 ;
        RECT 570.600 150.600 571.200 152.400 ;
        RECT 570.400 150.000 571.200 150.600 ;
        RECT 577.200 150.000 600.600 150.600 ;
        RECT 570.400 148.000 571.000 150.000 ;
        RECT 577.200 149.400 578.000 150.000 ;
        RECT 594.800 149.600 595.600 150.000 ;
        RECT 598.000 149.600 598.800 150.000 ;
        RECT 599.800 149.800 600.600 150.000 ;
        RECT 571.600 148.600 575.400 149.400 ;
        RECT 570.400 147.400 571.600 148.000 ;
        RECT 569.000 146.000 570.000 146.800 ;
        RECT 569.200 142.200 570.000 146.000 ;
        RECT 570.800 142.200 571.600 147.400 ;
        RECT 574.600 147.400 575.400 148.600 ;
        RECT 574.600 146.800 576.400 147.400 ;
        RECT 575.600 146.200 576.400 146.800 ;
        RECT 580.400 146.400 581.200 149.200 ;
        RECT 583.600 148.600 586.800 149.400 ;
        RECT 590.600 148.600 592.600 149.400 ;
        RECT 601.200 149.000 602.000 154.600 ;
        RECT 583.200 147.800 584.000 148.000 ;
        RECT 583.200 147.200 587.600 147.800 ;
        RECT 586.800 147.000 587.600 147.200 ;
        RECT 588.400 146.800 589.200 148.400 ;
        RECT 575.600 145.400 578.000 146.200 ;
        RECT 580.400 145.600 581.400 146.400 ;
        RECT 584.400 145.600 586.000 146.400 ;
        RECT 586.800 146.200 587.600 146.400 ;
        RECT 590.600 146.200 591.400 148.600 ;
        RECT 593.200 148.200 602.000 149.000 ;
        RECT 596.600 146.800 599.600 147.600 ;
        RECT 596.600 146.200 597.400 146.800 ;
        RECT 586.800 145.600 591.400 146.200 ;
        RECT 577.200 142.200 578.000 145.400 ;
        RECT 594.800 145.400 597.400 146.200 ;
        RECT 578.800 142.200 579.600 145.000 ;
        RECT 580.400 142.200 581.200 145.000 ;
        RECT 582.000 142.200 582.800 145.000 ;
        RECT 583.600 142.200 584.400 145.000 ;
        RECT 586.800 142.200 587.600 145.000 ;
        RECT 590.000 142.200 590.800 145.000 ;
        RECT 591.600 142.200 592.400 145.000 ;
        RECT 593.200 142.200 594.000 145.000 ;
        RECT 594.800 142.200 595.600 145.400 ;
        RECT 601.200 142.200 602.000 148.200 ;
        RECT 602.800 142.200 603.600 159.800 ;
        RECT 606.000 152.400 606.800 159.800 ;
        RECT 606.000 151.800 608.200 152.400 ;
        RECT 607.600 151.200 608.200 151.800 ;
        RECT 607.600 150.400 608.800 151.200 ;
        RECT 606.000 148.800 606.800 150.400 ;
        RECT 607.600 147.400 608.200 150.400 ;
        RECT 606.000 146.800 608.200 147.400 ;
        RECT 606.000 142.200 606.800 146.800 ;
        RECT 2.800 136.000 3.600 139.800 ;
        RECT 2.600 135.200 3.600 136.000 ;
        RECT 2.600 130.800 3.400 135.200 ;
        RECT 4.400 134.600 5.200 139.800 ;
        RECT 10.800 136.600 11.600 139.800 ;
        RECT 12.400 137.000 13.200 139.800 ;
        RECT 14.000 137.000 14.800 139.800 ;
        RECT 15.600 137.000 16.400 139.800 ;
        RECT 17.200 137.000 18.000 139.800 ;
        RECT 20.400 137.000 21.200 139.800 ;
        RECT 23.600 137.000 24.400 139.800 ;
        RECT 25.200 137.000 26.000 139.800 ;
        RECT 26.800 137.000 27.600 139.800 ;
        RECT 9.200 135.800 11.600 136.600 ;
        RECT 28.400 136.600 29.200 139.800 ;
        RECT 9.200 135.200 10.000 135.800 ;
        RECT 4.000 134.000 5.200 134.600 ;
        RECT 8.200 134.600 10.000 135.200 ;
        RECT 14.000 135.600 15.000 136.400 ;
        RECT 18.000 135.600 19.600 136.400 ;
        RECT 20.400 135.800 25.000 136.400 ;
        RECT 28.400 135.800 31.000 136.600 ;
        RECT 20.400 135.600 21.200 135.800 ;
        RECT 4.000 132.000 4.600 134.000 ;
        RECT 8.200 133.400 9.000 134.600 ;
        RECT 5.200 132.600 9.000 133.400 ;
        RECT 14.000 132.800 14.800 135.600 ;
        RECT 20.400 134.800 21.200 135.000 ;
        RECT 16.800 134.200 21.200 134.800 ;
        RECT 16.800 134.000 17.600 134.200 ;
        RECT 22.000 133.600 22.800 135.200 ;
        RECT 24.200 133.400 25.000 135.800 ;
        RECT 30.200 135.200 31.000 135.800 ;
        RECT 30.200 134.400 33.200 135.200 ;
        RECT 34.800 133.800 35.600 139.800 ;
        RECT 39.000 136.400 39.800 139.800 ;
        RECT 38.000 135.800 39.800 136.400 ;
        RECT 17.200 132.600 20.400 133.400 ;
        RECT 24.200 132.600 26.200 133.400 ;
        RECT 26.800 133.000 35.600 133.800 ;
        RECT 36.400 133.600 37.200 135.200 ;
        RECT 10.800 132.000 11.600 132.600 ;
        RECT 28.400 132.000 29.200 132.400 ;
        RECT 30.000 132.000 30.800 132.400 ;
        RECT 33.400 132.000 34.200 132.200 ;
        RECT 4.000 131.400 4.800 132.000 ;
        RECT 10.800 131.400 34.200 132.000 ;
        RECT 2.600 130.000 3.600 130.800 ;
        RECT 2.800 122.200 3.600 130.000 ;
        RECT 4.200 129.600 4.800 131.400 ;
        RECT 4.200 129.000 13.200 129.600 ;
        RECT 4.200 127.400 4.800 129.000 ;
        RECT 12.400 128.800 13.200 129.000 ;
        RECT 15.600 129.000 24.200 129.600 ;
        RECT 15.600 128.800 16.400 129.000 ;
        RECT 7.400 127.600 10.000 128.400 ;
        RECT 4.200 126.800 6.800 127.400 ;
        RECT 6.000 122.200 6.800 126.800 ;
        RECT 9.200 122.200 10.000 127.600 ;
        RECT 10.600 126.800 14.800 127.600 ;
        RECT 12.400 122.200 13.200 125.000 ;
        RECT 14.000 122.200 14.800 125.000 ;
        RECT 15.600 122.200 16.400 125.000 ;
        RECT 17.200 122.200 18.000 128.400 ;
        RECT 20.400 127.600 23.000 128.400 ;
        RECT 23.600 128.200 24.200 129.000 ;
        RECT 25.200 129.400 26.000 129.600 ;
        RECT 25.200 129.000 30.600 129.400 ;
        RECT 25.200 128.800 31.400 129.000 ;
        RECT 30.000 128.200 31.400 128.800 ;
        RECT 23.600 127.600 29.400 128.200 ;
        RECT 32.400 128.000 34.000 128.800 ;
        RECT 32.400 127.600 33.000 128.000 ;
        RECT 20.400 122.200 21.200 127.000 ;
        RECT 23.600 122.200 24.400 127.000 ;
        RECT 28.800 126.800 33.000 127.600 ;
        RECT 34.800 127.400 35.600 133.000 ;
        RECT 33.600 126.800 35.600 127.400 ;
        RECT 38.000 132.300 38.800 135.800 ;
        RECT 41.200 135.600 42.000 139.800 ;
        RECT 42.800 136.000 43.600 139.800 ;
        RECT 46.000 136.000 46.800 139.800 ;
        RECT 51.400 136.000 52.200 139.000 ;
        RECT 55.600 137.000 56.400 139.000 ;
        RECT 42.800 135.800 46.800 136.000 ;
        RECT 41.400 134.400 42.000 135.600 ;
        RECT 43.000 135.400 46.600 135.800 ;
        RECT 50.600 135.400 52.200 136.000 ;
        RECT 50.600 135.000 51.400 135.400 ;
        RECT 45.200 134.400 46.000 134.800 ;
        RECT 50.600 134.400 51.200 135.000 ;
        RECT 55.800 134.800 56.400 137.000 ;
        RECT 57.200 136.000 58.000 139.800 ;
        RECT 60.400 136.000 61.200 139.800 ;
        RECT 57.200 135.800 61.200 136.000 ;
        RECT 62.000 135.800 62.800 139.800 ;
        RECT 63.600 135.800 64.400 139.800 ;
        RECT 65.200 136.000 66.000 139.800 ;
        RECT 68.400 136.000 69.200 139.800 ;
        RECT 65.200 135.800 69.200 136.000 ;
        RECT 57.400 135.400 61.000 135.800 ;
        RECT 41.200 133.600 43.800 134.400 ;
        RECT 45.200 133.800 46.800 134.400 ;
        RECT 46.000 133.600 46.800 133.800 ;
        RECT 49.200 133.600 51.200 134.400 ;
        RECT 52.200 134.200 56.400 134.800 ;
        RECT 58.000 134.400 58.800 134.800 ;
        RECT 62.000 134.400 62.600 135.800 ;
        RECT 63.800 134.400 64.400 135.800 ;
        RECT 65.400 135.400 69.000 135.800 ;
        RECT 70.000 135.000 70.800 139.800 ;
        RECT 74.400 138.400 75.200 139.800 ;
        RECT 73.200 137.800 75.200 138.400 ;
        RECT 78.800 137.800 79.600 139.800 ;
        RECT 83.000 138.400 84.200 139.800 ;
        RECT 82.800 137.800 84.200 138.400 ;
        RECT 73.200 137.000 74.000 137.800 ;
        RECT 78.800 137.200 79.400 137.800 ;
        RECT 74.800 136.400 75.600 137.200 ;
        RECT 76.600 136.600 79.400 137.200 ;
        RECT 82.800 137.000 83.600 137.800 ;
        RECT 76.600 136.400 77.400 136.600 ;
        RECT 67.600 134.400 68.400 134.800 ;
        RECT 52.200 133.800 53.200 134.200 ;
        RECT 38.000 131.700 41.900 132.300 ;
        RECT 25.200 122.200 26.000 125.000 ;
        RECT 26.800 122.200 27.600 125.000 ;
        RECT 30.000 122.200 30.800 126.800 ;
        RECT 33.600 126.200 34.200 126.800 ;
        RECT 33.200 125.600 34.200 126.200 ;
        RECT 33.200 122.200 34.000 125.600 ;
        RECT 38.000 122.200 38.800 131.700 ;
        RECT 41.300 130.400 41.900 131.700 ;
        RECT 39.600 128.800 40.400 130.400 ;
        RECT 41.200 130.200 42.000 130.400 ;
        RECT 43.200 130.200 43.800 133.600 ;
        RECT 44.400 131.600 45.200 133.200 ;
        RECT 49.200 130.800 50.000 132.400 ;
        RECT 41.200 129.600 42.600 130.200 ;
        RECT 43.200 129.600 44.200 130.200 ;
        RECT 42.000 128.400 42.600 129.600 ;
        RECT 42.000 127.600 42.800 128.400 ;
        RECT 43.400 122.200 44.200 129.600 ;
        RECT 50.600 129.800 51.200 133.600 ;
        RECT 51.800 133.000 53.200 133.800 ;
        RECT 57.200 133.800 58.800 134.400 ;
        RECT 57.200 133.600 58.000 133.800 ;
        RECT 60.200 133.600 62.800 134.400 ;
        RECT 63.600 133.600 66.200 134.400 ;
        RECT 67.600 133.800 69.200 134.400 ;
        RECT 68.400 133.600 69.200 133.800 ;
        RECT 70.800 134.200 72.400 134.400 ;
        RECT 75.000 134.200 75.600 136.400 ;
        RECT 84.600 135.400 85.400 135.600 ;
        RECT 87.600 135.400 88.400 139.800 ;
        RECT 90.800 136.400 91.600 139.800 ;
        RECT 84.600 134.800 88.400 135.400 ;
        RECT 76.400 134.200 77.200 134.400 ;
        RECT 80.600 134.200 81.400 134.400 ;
        RECT 70.800 133.600 81.800 134.200 ;
        RECT 52.600 131.000 53.200 133.000 ;
        RECT 54.000 131.600 54.800 133.200 ;
        RECT 55.600 131.600 56.400 133.200 ;
        RECT 58.800 131.600 59.600 133.200 ;
        RECT 60.200 132.300 60.800 133.600 ;
        RECT 65.600 132.400 66.200 133.600 ;
        RECT 73.800 133.400 74.600 133.600 ;
        RECT 60.200 131.700 64.300 132.300 ;
        RECT 52.600 130.400 56.400 131.000 ;
        RECT 50.600 129.200 52.200 129.800 ;
        RECT 51.400 124.400 52.200 129.200 ;
        RECT 55.800 127.000 56.400 130.400 ;
        RECT 60.200 130.200 60.800 131.700 ;
        RECT 63.700 130.400 64.300 131.700 ;
        RECT 65.200 131.600 66.200 132.400 ;
        RECT 66.800 131.600 67.600 133.200 ;
        RECT 72.200 132.400 73.000 132.600 ;
        RECT 74.800 132.400 75.600 132.600 ;
        RECT 72.200 131.800 77.200 132.400 ;
        RECT 76.400 131.600 77.200 131.800 ;
        RECT 62.000 130.200 62.800 130.400 ;
        RECT 50.800 123.600 52.200 124.400 ;
        RECT 51.400 122.200 52.200 123.600 ;
        RECT 55.600 123.000 56.400 127.000 ;
        RECT 59.800 129.600 60.800 130.200 ;
        RECT 61.400 129.600 62.800 130.200 ;
        RECT 63.600 130.200 64.400 130.400 ;
        RECT 65.600 130.200 66.200 131.600 ;
        RECT 70.000 131.000 75.600 131.200 ;
        RECT 70.000 130.800 75.800 131.000 ;
        RECT 70.000 130.600 79.800 130.800 ;
        RECT 63.600 129.600 65.000 130.200 ;
        RECT 65.600 129.600 66.600 130.200 ;
        RECT 59.800 122.200 60.600 129.600 ;
        RECT 61.400 128.400 62.000 129.600 ;
        RECT 61.200 127.600 62.000 128.400 ;
        RECT 64.400 128.400 65.000 129.600 ;
        RECT 64.400 127.600 65.200 128.400 ;
        RECT 65.800 122.200 66.600 129.600 ;
        RECT 70.000 122.200 70.800 130.600 ;
        RECT 75.000 130.200 79.800 130.600 ;
        RECT 73.200 129.000 78.600 129.600 ;
        RECT 73.200 128.800 74.000 129.000 ;
        RECT 77.800 128.800 78.600 129.000 ;
        RECT 79.200 129.000 79.800 130.200 ;
        RECT 81.200 130.400 81.800 133.600 ;
        RECT 82.800 132.800 83.600 133.000 ;
        RECT 82.800 132.200 86.600 132.800 ;
        RECT 85.800 132.000 86.600 132.200 ;
        RECT 84.200 131.400 85.000 131.600 ;
        RECT 87.600 131.400 88.400 134.800 ;
        RECT 90.600 135.800 91.600 136.400 ;
        RECT 90.600 134.400 91.200 135.800 ;
        RECT 94.000 135.200 94.800 139.800 ;
        RECT 95.600 135.800 96.400 139.800 ;
        RECT 97.200 136.000 98.000 139.800 ;
        RECT 100.400 136.000 101.200 139.800 ;
        RECT 97.200 135.800 101.200 136.000 ;
        RECT 92.200 134.600 94.800 135.200 ;
        RECT 89.200 134.300 90.000 134.400 ;
        RECT 90.600 134.300 91.600 134.400 ;
        RECT 89.200 133.700 91.600 134.300 ;
        RECT 89.200 133.600 90.000 133.700 ;
        RECT 90.600 133.600 91.600 133.700 ;
        RECT 84.200 130.800 88.400 131.400 ;
        RECT 81.200 129.800 83.600 130.400 ;
        RECT 80.600 129.000 81.400 129.200 ;
        RECT 79.200 128.400 81.400 129.000 ;
        RECT 83.000 128.800 83.600 129.800 ;
        RECT 83.000 128.000 84.400 128.800 ;
        RECT 76.600 127.400 77.400 127.600 ;
        RECT 79.400 127.400 80.200 127.600 ;
        RECT 73.200 126.200 74.000 127.000 ;
        RECT 76.600 126.800 80.200 127.400 ;
        RECT 78.800 126.200 79.400 126.800 ;
        RECT 82.800 126.200 83.600 127.000 ;
        RECT 73.200 125.600 75.200 126.200 ;
        RECT 74.400 122.200 75.200 125.600 ;
        RECT 78.800 122.200 79.600 126.200 ;
        RECT 83.000 122.200 84.200 126.200 ;
        RECT 87.600 122.200 88.400 130.800 ;
        RECT 90.600 130.200 91.200 133.600 ;
        RECT 92.200 133.000 92.800 134.600 ;
        RECT 95.800 134.400 96.400 135.800 ;
        RECT 97.400 135.400 101.000 135.800 ;
        RECT 102.000 135.000 102.800 139.800 ;
        RECT 106.400 138.400 107.200 139.800 ;
        RECT 105.200 137.800 107.200 138.400 ;
        RECT 110.800 137.800 111.600 139.800 ;
        RECT 115.000 138.400 116.200 139.800 ;
        RECT 114.800 137.800 116.200 138.400 ;
        RECT 105.200 137.000 106.000 137.800 ;
        RECT 110.800 137.200 111.400 137.800 ;
        RECT 106.800 136.400 107.600 137.200 ;
        RECT 108.600 136.600 111.400 137.200 ;
        RECT 114.800 137.000 115.600 137.800 ;
        RECT 108.600 136.400 109.400 136.600 ;
        RECT 99.600 134.400 100.400 134.800 ;
        RECT 95.600 133.600 98.200 134.400 ;
        RECT 99.600 133.800 101.200 134.400 ;
        RECT 100.400 133.600 101.200 133.800 ;
        RECT 102.800 134.200 104.400 134.400 ;
        RECT 107.000 134.200 107.600 136.400 ;
        RECT 116.600 135.400 117.400 135.600 ;
        RECT 119.600 135.400 120.400 139.800 ;
        RECT 123.800 138.400 124.600 139.800 ;
        RECT 122.800 137.600 124.600 138.400 ;
        RECT 123.800 136.400 124.600 137.600 ;
        RECT 116.600 134.800 120.400 135.400 ;
        RECT 122.800 135.800 124.600 136.400 ;
        RECT 112.600 134.200 113.400 134.400 ;
        RECT 102.800 133.600 113.800 134.200 ;
        RECT 91.800 132.200 92.800 133.000 ;
        RECT 92.200 130.200 92.800 132.200 ;
        RECT 93.800 132.400 94.600 133.200 ;
        RECT 93.800 131.600 94.800 132.400 ;
        RECT 95.600 130.200 96.400 130.400 ;
        RECT 97.600 130.200 98.200 133.600 ;
        RECT 105.800 133.400 106.600 133.600 ;
        RECT 98.800 131.600 99.600 133.200 ;
        RECT 104.200 132.400 105.000 132.600 ;
        RECT 106.800 132.400 107.600 132.600 ;
        RECT 104.200 131.800 109.200 132.400 ;
        RECT 108.400 131.600 109.200 131.800 ;
        RECT 102.000 131.000 107.600 131.200 ;
        RECT 102.000 130.800 107.800 131.000 ;
        RECT 102.000 130.600 111.800 130.800 ;
        RECT 90.600 129.200 91.600 130.200 ;
        RECT 92.200 129.600 94.800 130.200 ;
        RECT 95.600 129.600 97.000 130.200 ;
        RECT 97.600 129.600 98.600 130.200 ;
        RECT 90.800 122.200 91.600 129.200 ;
        RECT 94.000 122.200 94.800 129.600 ;
        RECT 96.400 128.400 97.000 129.600 ;
        RECT 96.400 127.600 97.200 128.400 ;
        RECT 97.800 122.200 98.600 129.600 ;
        RECT 102.000 122.200 102.800 130.600 ;
        RECT 107.000 130.200 111.800 130.600 ;
        RECT 105.200 129.000 110.600 129.600 ;
        RECT 105.200 128.800 106.000 129.000 ;
        RECT 109.800 128.800 110.600 129.000 ;
        RECT 111.200 129.000 111.800 130.200 ;
        RECT 113.200 130.400 113.800 133.600 ;
        RECT 114.800 132.800 115.600 133.000 ;
        RECT 114.800 132.200 118.600 132.800 ;
        RECT 117.800 132.000 118.600 132.200 ;
        RECT 116.200 131.400 117.000 131.600 ;
        RECT 119.600 131.400 120.400 134.800 ;
        RECT 121.200 133.600 122.000 135.200 ;
        RECT 116.200 130.800 120.400 131.400 ;
        RECT 113.200 129.800 115.600 130.400 ;
        RECT 112.600 129.000 113.400 129.200 ;
        RECT 111.200 128.400 113.400 129.000 ;
        RECT 115.000 128.800 115.600 129.800 ;
        RECT 115.000 128.000 116.400 128.800 ;
        RECT 108.600 127.400 109.400 127.600 ;
        RECT 111.400 127.400 112.200 127.600 ;
        RECT 105.200 126.200 106.000 127.000 ;
        RECT 108.600 126.800 112.200 127.400 ;
        RECT 110.800 126.200 111.400 126.800 ;
        RECT 114.800 126.200 115.600 127.000 ;
        RECT 105.200 125.600 107.200 126.200 ;
        RECT 106.400 122.200 107.200 125.600 ;
        RECT 110.800 122.200 111.600 126.200 ;
        RECT 115.000 122.200 116.200 126.200 ;
        RECT 119.600 122.200 120.400 130.800 ;
        RECT 122.800 122.200 123.600 135.800 ;
        RECT 126.000 135.600 126.800 137.200 ;
        RECT 124.400 128.800 125.200 130.400 ;
        RECT 127.600 122.200 128.400 139.800 ;
        RECT 131.800 136.400 132.600 139.800 ;
        RECT 130.800 135.800 132.600 136.400 ;
        RECT 134.000 136.000 134.800 139.800 ;
        RECT 137.200 136.000 138.000 139.800 ;
        RECT 134.000 135.800 138.000 136.000 ;
        RECT 129.200 133.600 130.000 135.200 ;
        RECT 130.800 122.200 131.600 135.800 ;
        RECT 134.200 135.400 137.800 135.800 ;
        RECT 138.800 135.600 139.600 139.800 ;
        RECT 140.400 136.000 141.200 139.800 ;
        RECT 143.600 136.000 144.400 139.800 ;
        RECT 140.400 135.800 144.400 136.000 ;
        RECT 145.200 135.800 146.000 139.800 ;
        RECT 147.400 136.400 148.200 139.800 ;
        RECT 147.400 135.800 149.200 136.400 ;
        RECT 156.400 136.000 157.200 139.800 ;
        RECT 159.600 136.000 160.400 139.800 ;
        RECT 156.400 135.800 160.400 136.000 ;
        RECT 161.200 135.800 162.000 139.800 ;
        RECT 164.400 136.000 165.200 139.800 ;
        RECT 134.800 134.400 135.600 134.800 ;
        RECT 138.800 134.400 139.400 135.600 ;
        RECT 140.600 135.400 144.200 135.800 ;
        RECT 141.200 134.400 142.000 134.800 ;
        RECT 145.200 134.400 145.800 135.800 ;
        RECT 134.000 133.800 135.600 134.400 ;
        RECT 134.000 133.600 134.800 133.800 ;
        RECT 137.000 133.600 139.600 134.400 ;
        RECT 140.400 133.800 142.000 134.400 ;
        RECT 140.400 133.600 141.200 133.800 ;
        RECT 143.400 133.600 146.000 134.400 ;
        RECT 135.600 131.600 136.400 133.200 ;
        RECT 132.400 128.800 133.200 130.400 ;
        RECT 137.000 130.200 137.600 133.600 ;
        RECT 142.000 131.600 142.800 133.200 ;
        RECT 138.800 130.200 139.600 130.400 ;
        RECT 143.400 130.200 144.000 133.600 ;
        RECT 145.200 132.300 146.000 132.400 ;
        RECT 148.400 132.300 149.200 135.800 ;
        RECT 156.600 135.400 160.200 135.800 ;
        RECT 150.000 133.600 150.800 135.200 ;
        RECT 157.200 134.400 158.000 134.800 ;
        RECT 161.200 134.400 161.800 135.800 ;
        RECT 164.200 135.200 165.200 136.000 ;
        RECT 156.400 133.800 158.000 134.400 ;
        RECT 156.400 133.600 157.200 133.800 ;
        RECT 159.400 133.600 162.000 134.400 ;
        RECT 145.200 131.700 149.200 132.300 ;
        RECT 145.200 131.600 146.000 131.700 ;
        RECT 145.200 130.200 146.000 130.400 ;
        RECT 136.600 129.600 137.600 130.200 ;
        RECT 138.200 129.600 139.600 130.200 ;
        RECT 143.000 129.600 144.000 130.200 ;
        RECT 144.600 129.600 146.000 130.200 ;
        RECT 136.600 122.200 137.400 129.600 ;
        RECT 138.200 128.400 138.800 129.600 ;
        RECT 138.000 127.600 138.800 128.400 ;
        RECT 143.000 124.400 143.800 129.600 ;
        RECT 144.600 128.400 145.200 129.600 ;
        RECT 146.800 128.800 147.600 130.400 ;
        RECT 144.400 127.600 145.200 128.400 ;
        RECT 148.400 128.300 149.200 131.700 ;
        RECT 158.000 131.600 158.800 133.200 ;
        RECT 159.400 130.200 160.000 133.600 ;
        RECT 164.200 130.800 165.000 135.200 ;
        RECT 166.000 134.600 166.800 139.800 ;
        RECT 172.400 136.600 173.200 139.800 ;
        RECT 174.000 137.000 174.800 139.800 ;
        RECT 175.600 137.000 176.400 139.800 ;
        RECT 177.200 137.000 178.000 139.800 ;
        RECT 178.800 137.000 179.600 139.800 ;
        RECT 182.000 137.000 182.800 139.800 ;
        RECT 185.200 137.000 186.000 139.800 ;
        RECT 186.800 137.000 187.600 139.800 ;
        RECT 188.400 137.000 189.200 139.800 ;
        RECT 170.800 135.800 173.200 136.600 ;
        RECT 190.000 136.600 190.800 139.800 ;
        RECT 170.800 135.200 171.600 135.800 ;
        RECT 165.600 134.000 166.800 134.600 ;
        RECT 169.800 134.600 171.600 135.200 ;
        RECT 175.600 135.600 176.600 136.400 ;
        RECT 179.600 135.600 181.200 136.400 ;
        RECT 182.000 135.800 186.600 136.400 ;
        RECT 190.000 135.800 192.600 136.600 ;
        RECT 182.000 135.600 182.800 135.800 ;
        RECT 165.600 132.000 166.200 134.000 ;
        RECT 169.800 133.400 170.600 134.600 ;
        RECT 166.800 132.600 170.600 133.400 ;
        RECT 175.600 132.800 176.400 135.600 ;
        RECT 182.000 134.800 182.800 135.000 ;
        RECT 178.400 134.200 182.800 134.800 ;
        RECT 178.400 134.000 179.200 134.200 ;
        RECT 183.600 133.600 184.400 135.200 ;
        RECT 185.800 133.400 186.600 135.800 ;
        RECT 191.800 135.200 192.600 135.800 ;
        RECT 191.800 134.400 194.800 135.200 ;
        RECT 196.400 133.800 197.200 139.800 ;
        RECT 198.600 138.400 199.400 139.800 ;
        RECT 198.000 137.600 199.400 138.400 ;
        RECT 198.600 136.400 199.400 137.600 ;
        RECT 204.400 136.400 205.200 139.800 ;
        RECT 198.600 135.800 200.400 136.400 ;
        RECT 178.800 132.600 182.000 133.400 ;
        RECT 185.800 132.600 187.800 133.400 ;
        RECT 188.400 133.000 197.200 133.800 ;
        RECT 172.400 132.000 173.200 132.600 ;
        RECT 183.600 132.000 184.400 132.400 ;
        RECT 190.000 132.000 190.800 132.400 ;
        RECT 193.200 132.000 194.000 132.400 ;
        RECT 195.000 132.000 195.800 132.200 ;
        RECT 165.600 131.400 166.400 132.000 ;
        RECT 172.400 131.400 195.800 132.000 ;
        RECT 161.200 130.200 162.000 130.400 ;
        RECT 159.000 129.600 160.000 130.200 ;
        RECT 160.600 129.600 162.000 130.200 ;
        RECT 164.200 130.000 165.200 130.800 ;
        RECT 153.200 128.300 154.000 128.400 ;
        RECT 148.400 127.700 154.000 128.300 ;
        RECT 142.000 123.600 143.800 124.400 ;
        RECT 143.000 122.200 143.800 123.600 ;
        RECT 148.400 122.200 149.200 127.700 ;
        RECT 153.200 127.600 154.000 127.700 ;
        RECT 159.000 122.200 159.800 129.600 ;
        RECT 160.600 128.400 161.200 129.600 ;
        RECT 160.400 127.600 161.200 128.400 ;
        RECT 164.400 122.200 165.200 130.000 ;
        RECT 165.800 129.600 166.400 131.400 ;
        RECT 165.800 129.000 174.800 129.600 ;
        RECT 165.800 127.400 166.400 129.000 ;
        RECT 174.000 128.800 174.800 129.000 ;
        RECT 177.200 129.000 185.800 129.600 ;
        RECT 177.200 128.800 178.000 129.000 ;
        RECT 169.000 127.600 171.600 128.400 ;
        RECT 165.800 126.800 168.400 127.400 ;
        RECT 167.600 122.200 168.400 126.800 ;
        RECT 170.800 122.200 171.600 127.600 ;
        RECT 172.200 126.800 176.400 127.600 ;
        RECT 174.000 122.200 174.800 125.000 ;
        RECT 175.600 122.200 176.400 125.000 ;
        RECT 177.200 122.200 178.000 125.000 ;
        RECT 178.800 122.200 179.600 128.400 ;
        RECT 182.000 127.600 184.600 128.400 ;
        RECT 185.200 128.200 185.800 129.000 ;
        RECT 186.800 129.400 187.600 129.600 ;
        RECT 186.800 129.000 192.200 129.400 ;
        RECT 186.800 128.800 193.000 129.000 ;
        RECT 191.600 128.200 193.000 128.800 ;
        RECT 185.200 127.600 191.000 128.200 ;
        RECT 194.000 128.000 195.600 128.800 ;
        RECT 194.000 127.600 194.600 128.000 ;
        RECT 182.000 122.200 182.800 127.000 ;
        RECT 185.200 122.200 186.000 127.000 ;
        RECT 190.400 126.800 194.600 127.600 ;
        RECT 196.400 127.400 197.200 133.000 ;
        RECT 198.000 128.800 198.800 130.400 ;
        RECT 195.200 126.800 197.200 127.400 ;
        RECT 186.800 122.200 187.600 125.000 ;
        RECT 188.400 122.200 189.200 125.000 ;
        RECT 191.600 122.200 192.400 126.800 ;
        RECT 195.200 126.200 195.800 126.800 ;
        RECT 194.800 125.600 195.800 126.200 ;
        RECT 194.800 122.200 195.600 125.600 ;
        RECT 199.600 122.200 200.400 135.800 ;
        RECT 204.200 135.800 205.200 136.400 ;
        RECT 201.200 133.600 202.000 135.200 ;
        RECT 204.200 134.400 204.800 135.800 ;
        RECT 207.600 135.200 208.400 139.800 ;
        RECT 210.800 136.000 211.600 139.800 ;
        RECT 205.800 134.600 208.400 135.200 ;
        RECT 210.600 135.200 211.600 136.000 ;
        RECT 202.800 134.300 203.600 134.400 ;
        RECT 204.200 134.300 205.200 134.400 ;
        RECT 202.800 133.700 205.200 134.300 ;
        RECT 202.800 133.600 203.600 133.700 ;
        RECT 204.200 133.600 205.200 133.700 ;
        RECT 204.200 130.200 204.800 133.600 ;
        RECT 205.800 133.000 206.400 134.600 ;
        RECT 205.400 132.200 206.400 133.000 ;
        RECT 205.800 130.200 206.400 132.200 ;
        RECT 207.400 132.400 208.200 133.200 ;
        RECT 207.400 131.600 208.400 132.400 ;
        RECT 210.600 130.800 211.400 135.200 ;
        RECT 212.400 134.600 213.200 139.800 ;
        RECT 218.800 136.600 219.600 139.800 ;
        RECT 220.400 137.000 221.200 139.800 ;
        RECT 222.000 137.000 222.800 139.800 ;
        RECT 223.600 137.000 224.400 139.800 ;
        RECT 225.200 137.000 226.000 139.800 ;
        RECT 228.400 137.000 229.200 139.800 ;
        RECT 231.600 137.000 232.400 139.800 ;
        RECT 233.200 137.000 234.000 139.800 ;
        RECT 234.800 137.000 235.600 139.800 ;
        RECT 217.200 135.800 219.600 136.600 ;
        RECT 236.400 136.600 237.200 139.800 ;
        RECT 217.200 135.200 218.000 135.800 ;
        RECT 212.000 134.000 213.200 134.600 ;
        RECT 216.200 134.600 218.000 135.200 ;
        RECT 222.000 135.600 223.000 136.400 ;
        RECT 226.000 135.600 227.600 136.400 ;
        RECT 228.400 135.800 233.000 136.400 ;
        RECT 236.400 135.800 239.000 136.600 ;
        RECT 228.400 135.600 229.200 135.800 ;
        RECT 212.000 132.000 212.600 134.000 ;
        RECT 216.200 133.400 217.000 134.600 ;
        RECT 213.200 132.600 217.000 133.400 ;
        RECT 222.000 132.800 222.800 135.600 ;
        RECT 228.400 134.800 229.200 135.000 ;
        RECT 224.800 134.200 229.200 134.800 ;
        RECT 224.800 134.000 225.600 134.200 ;
        RECT 230.000 133.600 230.800 135.200 ;
        RECT 232.200 133.400 233.000 135.800 ;
        RECT 238.200 135.200 239.000 135.800 ;
        RECT 238.200 134.400 241.200 135.200 ;
        RECT 242.800 133.800 243.600 139.800 ;
        RECT 246.000 137.800 246.800 139.800 ;
        RECT 250.800 137.800 251.600 139.800 ;
        RECT 246.000 134.400 246.600 137.800 ;
        RECT 247.600 135.600 248.400 137.200 ;
        RECT 249.200 135.600 250.000 137.200 ;
        RECT 251.000 134.400 251.600 137.800 ;
        RECT 254.000 135.200 254.800 139.800 ;
        RECT 257.200 136.400 258.000 139.800 ;
        RECT 257.200 135.800 258.200 136.400 ;
        RECT 260.400 136.000 261.200 139.800 ;
        RECT 263.600 136.000 264.400 139.800 ;
        RECT 260.400 135.800 264.400 136.000 ;
        RECT 265.200 135.800 266.000 139.800 ;
        RECT 268.400 136.000 269.200 139.800 ;
        RECT 254.000 134.600 256.600 135.200 ;
        RECT 225.200 132.600 228.400 133.400 ;
        RECT 232.200 132.600 234.200 133.400 ;
        RECT 234.800 133.000 243.600 133.800 ;
        RECT 244.400 134.300 245.200 134.400 ;
        RECT 246.000 134.300 246.800 134.400 ;
        RECT 244.400 133.700 246.800 134.300 ;
        RECT 244.400 133.600 245.200 133.700 ;
        RECT 246.000 133.600 246.800 133.700 ;
        RECT 250.800 133.600 251.600 134.400 ;
        RECT 218.800 132.000 219.600 132.600 ;
        RECT 236.400 132.000 237.200 132.400 ;
        RECT 241.400 132.000 242.200 132.200 ;
        RECT 212.000 131.400 212.800 132.000 ;
        RECT 218.800 131.400 242.200 132.000 ;
        RECT 209.200 130.300 210.000 130.400 ;
        RECT 210.600 130.300 211.600 130.800 ;
        RECT 204.200 129.200 205.200 130.200 ;
        RECT 205.800 129.600 208.400 130.200 ;
        RECT 209.200 129.700 211.600 130.300 ;
        RECT 209.200 129.600 210.000 129.700 ;
        RECT 204.400 122.200 205.200 129.200 ;
        RECT 207.600 122.200 208.400 129.600 ;
        RECT 210.800 122.200 211.600 129.700 ;
        RECT 212.200 129.600 212.800 131.400 ;
        RECT 212.200 129.000 221.200 129.600 ;
        RECT 212.200 127.400 212.800 129.000 ;
        RECT 220.400 128.800 221.200 129.000 ;
        RECT 223.600 129.000 232.200 129.600 ;
        RECT 223.600 128.800 224.400 129.000 ;
        RECT 215.400 127.600 218.000 128.400 ;
        RECT 212.200 126.800 214.800 127.400 ;
        RECT 214.000 122.200 214.800 126.800 ;
        RECT 217.200 122.200 218.000 127.600 ;
        RECT 218.600 126.800 222.800 127.600 ;
        RECT 220.400 122.200 221.200 125.000 ;
        RECT 222.000 122.200 222.800 125.000 ;
        RECT 223.600 122.200 224.400 125.000 ;
        RECT 225.200 122.200 226.000 128.400 ;
        RECT 228.400 127.600 231.000 128.400 ;
        RECT 231.600 128.200 232.200 129.000 ;
        RECT 233.200 129.400 234.000 129.600 ;
        RECT 233.200 129.000 238.600 129.400 ;
        RECT 233.200 128.800 239.400 129.000 ;
        RECT 238.000 128.200 239.400 128.800 ;
        RECT 231.600 127.600 237.400 128.200 ;
        RECT 240.400 128.000 242.000 128.800 ;
        RECT 240.400 127.600 241.000 128.000 ;
        RECT 228.400 122.200 229.200 127.000 ;
        RECT 231.600 122.200 232.400 127.000 ;
        RECT 236.800 126.800 241.000 127.600 ;
        RECT 242.800 127.400 243.600 133.000 ;
        RECT 244.400 130.800 245.200 132.400 ;
        RECT 246.000 130.200 246.600 133.600 ;
        RECT 251.000 130.200 251.600 133.600 ;
        RECT 254.200 132.400 255.000 133.200 ;
        RECT 252.400 130.800 253.200 132.400 ;
        RECT 254.000 131.600 255.000 132.400 ;
        RECT 256.000 133.000 256.600 134.600 ;
        RECT 257.600 134.400 258.200 135.800 ;
        RECT 260.600 135.400 264.200 135.800 ;
        RECT 261.200 134.400 262.000 134.800 ;
        RECT 265.200 134.400 265.800 135.800 ;
        RECT 268.200 135.200 269.200 136.000 ;
        RECT 257.200 133.600 258.200 134.400 ;
        RECT 260.400 133.800 262.000 134.400 ;
        RECT 260.400 133.600 261.200 133.800 ;
        RECT 263.400 133.600 266.000 134.400 ;
        RECT 256.000 132.200 257.000 133.000 ;
        RECT 256.000 130.200 256.600 132.200 ;
        RECT 257.600 130.200 258.200 133.600 ;
        RECT 262.000 131.600 262.800 133.200 ;
        RECT 263.400 130.200 264.000 133.600 ;
        RECT 268.200 130.800 269.000 135.200 ;
        RECT 270.000 134.600 270.800 139.800 ;
        RECT 276.400 136.600 277.200 139.800 ;
        RECT 278.000 137.000 278.800 139.800 ;
        RECT 279.600 137.000 280.400 139.800 ;
        RECT 281.200 137.000 282.000 139.800 ;
        RECT 282.800 137.000 283.600 139.800 ;
        RECT 286.000 137.000 286.800 139.800 ;
        RECT 289.200 137.000 290.000 139.800 ;
        RECT 290.800 137.000 291.600 139.800 ;
        RECT 292.400 137.000 293.200 139.800 ;
        RECT 274.800 135.800 277.200 136.600 ;
        RECT 294.000 136.600 294.800 139.800 ;
        RECT 274.800 135.200 275.600 135.800 ;
        RECT 269.600 134.000 270.800 134.600 ;
        RECT 273.800 134.600 275.600 135.200 ;
        RECT 279.600 135.600 280.600 136.400 ;
        RECT 283.600 135.600 285.200 136.400 ;
        RECT 286.000 135.800 290.600 136.400 ;
        RECT 294.000 135.800 296.600 136.600 ;
        RECT 286.000 135.600 286.800 135.800 ;
        RECT 269.600 132.000 270.200 134.000 ;
        RECT 273.800 133.400 274.600 134.600 ;
        RECT 270.800 132.600 274.600 133.400 ;
        RECT 279.600 132.800 280.400 135.600 ;
        RECT 286.000 134.800 286.800 135.000 ;
        RECT 282.400 134.200 286.800 134.800 ;
        RECT 282.400 134.000 283.200 134.200 ;
        RECT 287.600 133.600 288.400 135.200 ;
        RECT 289.800 133.400 290.600 135.800 ;
        RECT 295.800 135.200 296.600 135.800 ;
        RECT 295.800 134.400 298.800 135.200 ;
        RECT 300.400 133.800 301.200 139.800 ;
        RECT 308.400 135.200 309.200 139.800 ;
        RECT 311.600 135.200 312.400 139.800 ;
        RECT 314.800 135.200 315.600 139.800 ;
        RECT 318.000 135.200 318.800 139.800 ;
        RECT 282.800 132.600 286.000 133.400 ;
        RECT 289.800 132.600 291.800 133.400 ;
        RECT 292.400 133.000 301.200 133.800 ;
        RECT 276.400 132.000 277.200 132.600 ;
        RECT 287.600 132.000 288.400 132.400 ;
        RECT 294.000 132.000 294.800 132.400 ;
        RECT 299.000 132.000 299.800 132.200 ;
        RECT 269.600 131.400 270.400 132.000 ;
        RECT 276.400 131.400 299.800 132.000 ;
        RECT 265.200 130.300 266.000 130.400 ;
        RECT 268.200 130.300 269.200 130.800 ;
        RECT 265.200 130.200 269.200 130.300 ;
        RECT 241.600 126.800 243.600 127.400 ;
        RECT 245.000 129.400 246.800 130.200 ;
        RECT 250.800 129.400 252.600 130.200 ;
        RECT 233.200 122.200 234.000 125.000 ;
        RECT 234.800 122.200 235.600 125.000 ;
        RECT 238.000 122.200 238.800 126.800 ;
        RECT 241.600 126.200 242.200 126.800 ;
        RECT 241.200 125.600 242.200 126.200 ;
        RECT 241.200 122.200 242.000 125.600 ;
        RECT 245.000 122.200 245.800 129.400 ;
        RECT 251.800 124.400 252.600 129.400 ;
        RECT 250.800 123.600 252.600 124.400 ;
        RECT 251.800 122.200 252.600 123.600 ;
        RECT 254.000 129.600 256.600 130.200 ;
        RECT 254.000 122.200 254.800 129.600 ;
        RECT 257.200 129.200 258.200 130.200 ;
        RECT 263.000 129.600 264.000 130.200 ;
        RECT 264.600 129.700 269.200 130.200 ;
        RECT 264.600 129.600 266.000 129.700 ;
        RECT 257.200 122.200 258.000 129.200 ;
        RECT 263.000 122.200 263.800 129.600 ;
        RECT 264.600 128.400 265.200 129.600 ;
        RECT 264.400 127.600 266.000 128.400 ;
        RECT 268.400 122.200 269.200 129.700 ;
        RECT 269.800 129.600 270.400 131.400 ;
        RECT 269.800 129.000 278.800 129.600 ;
        RECT 269.800 127.400 270.400 129.000 ;
        RECT 278.000 128.800 278.800 129.000 ;
        RECT 281.200 129.000 289.800 129.600 ;
        RECT 281.200 128.800 282.000 129.000 ;
        RECT 273.000 127.600 275.600 128.400 ;
        RECT 269.800 126.800 272.400 127.400 ;
        RECT 271.600 122.200 272.400 126.800 ;
        RECT 274.800 122.200 275.600 127.600 ;
        RECT 276.200 126.800 280.400 127.600 ;
        RECT 278.000 122.200 278.800 125.000 ;
        RECT 279.600 122.200 280.400 125.000 ;
        RECT 281.200 122.200 282.000 125.000 ;
        RECT 282.800 122.200 283.600 128.400 ;
        RECT 286.000 127.600 288.600 128.400 ;
        RECT 289.200 128.200 289.800 129.000 ;
        RECT 290.800 129.400 291.600 129.600 ;
        RECT 290.800 129.000 296.200 129.400 ;
        RECT 290.800 128.800 297.000 129.000 ;
        RECT 295.600 128.200 297.000 128.800 ;
        RECT 289.200 127.600 295.000 128.200 ;
        RECT 298.000 128.000 299.600 128.800 ;
        RECT 298.000 127.600 298.600 128.000 ;
        RECT 286.000 122.200 286.800 127.000 ;
        RECT 289.200 122.200 290.000 127.000 ;
        RECT 294.400 126.800 298.600 127.600 ;
        RECT 300.400 127.400 301.200 133.000 ;
        RECT 306.800 134.400 309.200 135.200 ;
        RECT 310.200 134.400 312.400 135.200 ;
        RECT 313.400 134.400 315.600 135.200 ;
        RECT 317.000 134.400 318.800 135.200 ;
        RECT 306.800 131.600 307.600 134.400 ;
        RECT 310.200 133.800 311.000 134.400 ;
        RECT 313.400 133.800 314.200 134.400 ;
        RECT 317.000 133.800 317.800 134.400 ;
        RECT 319.600 133.800 320.400 134.400 ;
        RECT 308.400 133.000 311.000 133.800 ;
        RECT 311.800 133.000 314.200 133.800 ;
        RECT 315.200 133.000 317.800 133.800 ;
        RECT 318.600 133.000 320.400 133.800 ;
        RECT 321.200 133.800 322.000 139.800 ;
        RECT 327.600 136.600 328.400 139.800 ;
        RECT 329.200 137.000 330.000 139.800 ;
        RECT 330.800 137.000 331.600 139.800 ;
        RECT 332.400 137.000 333.200 139.800 ;
        RECT 335.600 137.000 336.400 139.800 ;
        RECT 338.800 137.000 339.600 139.800 ;
        RECT 340.400 137.000 341.200 139.800 ;
        RECT 342.000 137.000 342.800 139.800 ;
        RECT 343.600 137.000 344.400 139.800 ;
        RECT 325.800 135.800 328.400 136.600 ;
        RECT 345.200 136.600 346.000 139.800 ;
        RECT 331.800 135.800 336.400 136.400 ;
        RECT 325.800 135.200 326.600 135.800 ;
        RECT 323.600 134.400 326.600 135.200 ;
        RECT 321.200 133.000 330.000 133.800 ;
        RECT 331.800 133.400 332.600 135.800 ;
        RECT 335.600 135.600 336.400 135.800 ;
        RECT 337.200 135.600 338.800 136.400 ;
        RECT 341.800 135.600 342.800 136.400 ;
        RECT 345.200 135.800 347.600 136.600 ;
        RECT 334.000 133.600 334.800 135.200 ;
        RECT 335.600 134.800 336.400 135.000 ;
        RECT 335.600 134.200 340.000 134.800 ;
        RECT 339.200 134.000 340.000 134.200 ;
        RECT 310.200 131.600 311.000 133.000 ;
        RECT 313.400 131.600 314.200 133.000 ;
        RECT 317.000 131.600 317.800 133.000 ;
        RECT 306.800 130.800 309.200 131.600 ;
        RECT 310.200 130.800 312.400 131.600 ;
        RECT 313.400 130.800 315.600 131.600 ;
        RECT 317.000 130.800 318.800 131.600 ;
        RECT 299.200 126.800 301.200 127.400 ;
        RECT 290.800 122.200 291.600 125.000 ;
        RECT 292.400 122.200 293.200 125.000 ;
        RECT 295.600 122.200 296.400 126.800 ;
        RECT 299.200 126.200 299.800 126.800 ;
        RECT 298.800 125.600 299.800 126.200 ;
        RECT 298.800 122.200 299.600 125.600 ;
        RECT 308.400 122.200 309.200 130.800 ;
        RECT 311.600 122.200 312.400 130.800 ;
        RECT 314.800 122.200 315.600 130.800 ;
        RECT 318.000 122.200 318.800 130.800 ;
        RECT 321.200 127.400 322.000 133.000 ;
        RECT 330.600 132.600 332.600 133.400 ;
        RECT 336.400 132.600 339.600 133.400 ;
        RECT 342.000 132.800 342.800 135.600 ;
        RECT 346.800 135.200 347.600 135.800 ;
        RECT 346.800 134.600 348.600 135.200 ;
        RECT 347.800 133.400 348.600 134.600 ;
        RECT 351.600 134.600 352.400 139.800 ;
        RECT 353.200 136.300 354.000 139.800 ;
        RECT 354.800 136.300 355.600 136.400 ;
        RECT 353.200 135.700 355.600 136.300 ;
        RECT 353.200 135.200 354.200 135.700 ;
        RECT 354.800 135.600 355.600 135.700 ;
        RECT 351.600 134.000 352.800 134.600 ;
        RECT 347.800 132.600 351.600 133.400 ;
        RECT 322.800 132.200 323.600 132.400 ;
        RECT 322.600 132.000 323.600 132.200 ;
        RECT 327.600 132.000 328.400 132.400 ;
        RECT 345.200 132.000 346.000 132.600 ;
        RECT 352.200 132.000 352.800 134.000 ;
        RECT 322.600 131.400 346.000 132.000 ;
        RECT 352.000 131.400 352.800 132.000 ;
        RECT 352.000 129.600 352.600 131.400 ;
        RECT 353.400 130.800 354.200 135.200 ;
        RECT 356.400 135.200 357.200 139.800 ;
        RECT 359.600 136.400 360.400 139.800 ;
        RECT 359.600 135.600 360.600 136.400 ;
        RECT 356.400 134.600 359.000 135.200 ;
        RECT 356.600 132.400 357.400 133.200 ;
        RECT 356.400 131.600 357.400 132.400 ;
        RECT 358.400 133.000 359.000 134.600 ;
        RECT 360.000 134.400 360.600 135.600 ;
        RECT 359.600 133.600 360.600 134.400 ;
        RECT 358.400 132.200 359.400 133.000 ;
        RECT 330.800 129.400 331.600 129.600 ;
        RECT 326.200 129.000 331.600 129.400 ;
        RECT 325.400 128.800 331.600 129.000 ;
        RECT 332.600 129.000 341.200 129.600 ;
        RECT 322.800 128.000 324.400 128.800 ;
        RECT 325.400 128.200 326.800 128.800 ;
        RECT 332.600 128.200 333.200 129.000 ;
        RECT 340.400 128.800 341.200 129.000 ;
        RECT 343.600 129.000 352.600 129.600 ;
        RECT 343.600 128.800 344.400 129.000 ;
        RECT 323.800 127.600 324.400 128.000 ;
        RECT 327.400 127.600 333.200 128.200 ;
        RECT 333.800 127.600 336.400 128.400 ;
        RECT 321.200 126.800 323.200 127.400 ;
        RECT 323.800 126.800 328.000 127.600 ;
        RECT 322.600 126.200 323.200 126.800 ;
        RECT 322.600 125.600 323.600 126.200 ;
        RECT 322.800 122.200 323.600 125.600 ;
        RECT 326.000 122.200 326.800 126.800 ;
        RECT 329.200 122.200 330.000 125.000 ;
        RECT 330.800 122.200 331.600 125.000 ;
        RECT 332.400 122.200 333.200 127.000 ;
        RECT 335.600 122.200 336.400 127.000 ;
        RECT 338.800 122.200 339.600 128.400 ;
        RECT 346.800 127.600 349.400 128.400 ;
        RECT 342.000 126.800 346.200 127.600 ;
        RECT 340.400 122.200 341.200 125.000 ;
        RECT 342.000 122.200 342.800 125.000 ;
        RECT 343.600 122.200 344.400 125.000 ;
        RECT 346.800 122.200 347.600 127.600 ;
        RECT 352.000 127.400 352.600 129.000 ;
        RECT 350.000 126.800 352.600 127.400 ;
        RECT 353.200 130.000 354.200 130.800 ;
        RECT 358.400 130.200 359.000 132.200 ;
        RECT 360.000 130.200 360.600 133.600 ;
        RECT 350.000 122.200 350.800 126.800 ;
        RECT 353.200 122.200 354.000 130.000 ;
        RECT 356.400 129.600 359.000 130.200 ;
        RECT 356.400 122.200 357.200 129.600 ;
        RECT 359.600 129.200 360.600 130.200 ;
        RECT 362.800 132.400 363.600 139.800 ;
        RECT 366.000 135.200 366.800 139.800 ;
        RECT 367.600 136.000 368.400 139.800 ;
        RECT 370.800 136.000 371.600 139.800 ;
        RECT 367.600 135.800 371.600 136.000 ;
        RECT 372.400 135.800 373.200 139.800 ;
        RECT 376.600 136.400 377.400 139.800 ;
        RECT 375.600 135.800 377.400 136.400 ;
        RECT 367.800 135.400 371.400 135.800 ;
        RECT 364.600 134.600 366.800 135.200 ;
        RECT 362.800 130.200 363.400 132.400 ;
        RECT 364.600 131.600 365.200 134.600 ;
        RECT 368.400 134.400 369.200 134.800 ;
        RECT 372.400 134.400 373.000 135.800 ;
        RECT 367.600 133.800 369.200 134.400 ;
        RECT 370.600 134.300 373.200 134.400 ;
        RECT 374.000 134.300 374.800 135.200 ;
        RECT 367.600 133.600 368.400 133.800 ;
        RECT 370.600 133.700 374.800 134.300 ;
        RECT 370.600 133.600 373.200 133.700 ;
        RECT 374.000 133.600 374.800 133.700 ;
        RECT 375.600 134.300 376.400 135.800 ;
        RECT 377.200 134.300 378.000 134.400 ;
        RECT 375.600 133.700 378.000 134.300 ;
        RECT 366.000 131.600 366.800 133.200 ;
        RECT 369.200 131.600 370.000 133.200 ;
        RECT 364.000 130.800 365.200 131.600 ;
        RECT 364.600 130.200 365.200 130.800 ;
        RECT 370.600 130.200 371.200 133.600 ;
        RECT 372.400 130.200 373.200 130.400 ;
        RECT 359.600 122.200 360.400 129.200 ;
        RECT 362.800 122.200 363.600 130.200 ;
        RECT 364.600 129.600 366.800 130.200 ;
        RECT 366.000 122.200 366.800 129.600 ;
        RECT 370.200 129.600 371.200 130.200 ;
        RECT 371.800 129.600 373.200 130.200 ;
        RECT 370.200 122.200 371.000 129.600 ;
        RECT 371.800 128.400 372.400 129.600 ;
        RECT 371.600 128.300 372.400 128.400 ;
        RECT 374.000 128.300 374.800 128.400 ;
        RECT 371.600 127.700 374.800 128.300 ;
        RECT 371.600 127.600 372.400 127.700 ;
        RECT 374.000 127.600 374.800 127.700 ;
        RECT 375.600 122.200 376.400 133.700 ;
        RECT 377.200 133.600 378.000 133.700 ;
        RECT 378.800 133.800 379.600 139.800 ;
        RECT 385.200 136.600 386.000 139.800 ;
        RECT 386.800 137.000 387.600 139.800 ;
        RECT 388.400 137.000 389.200 139.800 ;
        RECT 390.000 137.000 390.800 139.800 ;
        RECT 393.200 137.000 394.000 139.800 ;
        RECT 396.400 137.000 397.200 139.800 ;
        RECT 398.000 137.000 398.800 139.800 ;
        RECT 399.600 137.000 400.400 139.800 ;
        RECT 401.200 137.000 402.000 139.800 ;
        RECT 383.400 135.800 386.000 136.600 ;
        RECT 402.800 136.600 403.600 139.800 ;
        RECT 389.400 135.800 394.000 136.400 ;
        RECT 383.400 135.200 384.200 135.800 ;
        RECT 381.200 134.400 384.200 135.200 ;
        RECT 378.800 133.000 387.600 133.800 ;
        RECT 389.400 133.400 390.200 135.800 ;
        RECT 393.200 135.600 394.000 135.800 ;
        RECT 394.800 135.600 396.400 136.400 ;
        RECT 399.400 135.600 400.400 136.400 ;
        RECT 402.800 135.800 405.200 136.600 ;
        RECT 391.600 133.600 392.400 135.200 ;
        RECT 393.200 134.800 394.000 135.000 ;
        RECT 393.200 134.200 397.600 134.800 ;
        RECT 396.800 134.000 397.600 134.200 ;
        RECT 377.200 128.800 378.000 130.400 ;
        RECT 378.800 127.400 379.600 133.000 ;
        RECT 388.200 132.600 390.200 133.400 ;
        RECT 394.000 132.600 397.200 133.400 ;
        RECT 399.600 132.800 400.400 135.600 ;
        RECT 404.400 135.200 405.200 135.800 ;
        RECT 404.400 134.600 406.200 135.200 ;
        RECT 405.400 133.400 406.200 134.600 ;
        RECT 409.200 134.600 410.000 139.800 ;
        RECT 410.800 136.000 411.600 139.800 ;
        RECT 410.800 135.200 411.800 136.000 ;
        RECT 415.600 135.200 416.400 139.800 ;
        RECT 418.800 135.200 419.600 139.800 ;
        RECT 422.000 135.200 422.800 139.800 ;
        RECT 425.200 135.200 426.000 139.800 ;
        RECT 428.400 135.800 429.200 139.800 ;
        RECT 430.000 136.000 430.800 139.800 ;
        RECT 433.200 136.000 434.000 139.800 ;
        RECT 430.000 135.800 434.000 136.000 ;
        RECT 409.200 134.000 410.400 134.600 ;
        RECT 405.400 132.600 409.200 133.400 ;
        RECT 380.200 132.000 381.000 132.200 ;
        RECT 382.000 132.000 382.800 132.400 ;
        RECT 385.200 132.000 386.000 132.400 ;
        RECT 402.800 132.000 403.600 132.600 ;
        RECT 409.800 132.000 410.400 134.000 ;
        RECT 380.200 131.400 403.600 132.000 ;
        RECT 409.600 131.400 410.400 132.000 ;
        RECT 409.600 129.600 410.200 131.400 ;
        RECT 411.000 130.800 411.800 135.200 ;
        RECT 414.000 134.400 416.400 135.200 ;
        RECT 417.400 134.400 419.600 135.200 ;
        RECT 420.600 134.400 422.800 135.200 ;
        RECT 424.200 134.400 426.000 135.200 ;
        RECT 428.600 134.400 429.200 135.800 ;
        RECT 430.200 135.400 433.800 135.800 ;
        RECT 434.800 135.200 435.600 139.800 ;
        RECT 438.000 136.400 438.800 139.800 ;
        RECT 438.000 135.800 439.000 136.400 ;
        RECT 432.400 134.400 433.200 134.800 ;
        RECT 434.800 134.600 437.400 135.200 ;
        RECT 414.000 131.600 414.800 134.400 ;
        RECT 417.400 133.800 418.200 134.400 ;
        RECT 420.600 133.800 421.400 134.400 ;
        RECT 424.200 133.800 425.000 134.400 ;
        RECT 426.800 133.800 427.600 134.400 ;
        RECT 415.600 133.000 418.200 133.800 ;
        RECT 419.000 133.000 421.400 133.800 ;
        RECT 422.400 133.000 425.000 133.800 ;
        RECT 425.800 133.000 427.600 133.800 ;
        RECT 428.400 133.600 431.000 134.400 ;
        RECT 432.400 133.800 434.000 134.400 ;
        RECT 433.200 133.600 434.000 133.800 ;
        RECT 417.400 131.600 418.200 133.000 ;
        RECT 420.600 131.600 421.400 133.000 ;
        RECT 424.200 131.600 425.000 133.000 ;
        RECT 414.000 130.800 416.400 131.600 ;
        RECT 417.400 130.800 419.600 131.600 ;
        RECT 420.600 130.800 422.800 131.600 ;
        RECT 424.200 130.800 426.000 131.600 ;
        RECT 388.400 129.400 389.200 129.600 ;
        RECT 383.800 129.000 389.200 129.400 ;
        RECT 383.000 128.800 389.200 129.000 ;
        RECT 390.200 129.000 398.800 129.600 ;
        RECT 380.400 128.000 382.000 128.800 ;
        RECT 383.000 128.200 384.400 128.800 ;
        RECT 390.200 128.200 390.800 129.000 ;
        RECT 398.000 128.800 398.800 129.000 ;
        RECT 401.200 129.000 410.200 129.600 ;
        RECT 401.200 128.800 402.000 129.000 ;
        RECT 381.400 127.600 382.000 128.000 ;
        RECT 385.000 127.600 390.800 128.200 ;
        RECT 391.400 127.600 394.000 128.400 ;
        RECT 378.800 126.800 380.800 127.400 ;
        RECT 381.400 126.800 385.600 127.600 ;
        RECT 380.200 126.200 380.800 126.800 ;
        RECT 380.200 125.600 381.200 126.200 ;
        RECT 380.400 122.200 381.200 125.600 ;
        RECT 383.600 122.200 384.400 126.800 ;
        RECT 386.800 122.200 387.600 125.000 ;
        RECT 388.400 122.200 389.200 125.000 ;
        RECT 390.000 122.200 390.800 127.000 ;
        RECT 393.200 122.200 394.000 127.000 ;
        RECT 396.400 122.200 397.200 128.400 ;
        RECT 404.400 127.600 407.000 128.400 ;
        RECT 399.600 126.800 403.800 127.600 ;
        RECT 398.000 122.200 398.800 125.000 ;
        RECT 399.600 122.200 400.400 125.000 ;
        RECT 401.200 122.200 402.000 125.000 ;
        RECT 404.400 122.200 405.200 127.600 ;
        RECT 409.600 127.400 410.200 129.000 ;
        RECT 407.600 126.800 410.200 127.400 ;
        RECT 410.800 130.000 411.800 130.800 ;
        RECT 407.600 122.200 408.400 126.800 ;
        RECT 410.800 122.200 411.600 130.000 ;
        RECT 415.600 122.200 416.400 130.800 ;
        RECT 418.800 122.200 419.600 130.800 ;
        RECT 422.000 122.200 422.800 130.800 ;
        RECT 425.200 122.200 426.000 130.800 ;
        RECT 428.400 130.200 429.200 130.400 ;
        RECT 430.400 130.200 431.000 133.600 ;
        RECT 431.600 131.600 432.400 133.200 ;
        RECT 435.000 132.400 435.800 133.200 ;
        RECT 433.200 132.300 434.000 132.400 ;
        RECT 434.800 132.300 435.800 132.400 ;
        RECT 433.200 131.700 435.800 132.300 ;
        RECT 433.200 131.600 434.000 131.700 ;
        RECT 434.800 131.600 435.800 131.700 ;
        RECT 436.800 133.000 437.400 134.600 ;
        RECT 438.400 134.400 439.000 135.800 ;
        RECT 438.000 133.600 439.000 134.400 ;
        RECT 442.400 134.200 443.200 139.800 ;
        RECT 449.200 137.800 450.000 139.800 ;
        RECT 447.600 135.600 448.400 137.200 ;
        RECT 449.400 134.400 450.000 137.800 ;
        RECT 452.400 135.800 453.200 139.800 ;
        RECT 456.800 138.400 458.400 139.800 ;
        RECT 455.600 137.600 458.400 138.400 ;
        RECT 456.800 136.200 458.400 137.600 ;
        RECT 452.400 135.200 454.600 135.800 ;
        RECT 455.600 135.400 457.200 135.600 ;
        RECT 453.800 135.000 454.600 135.200 ;
        RECT 455.200 134.800 457.200 135.400 ;
        RECT 455.200 134.400 455.800 134.800 ;
        RECT 436.800 132.200 437.800 133.000 ;
        RECT 436.800 130.200 437.400 132.200 ;
        RECT 438.400 130.200 439.000 133.600 ;
        RECT 441.400 133.800 443.200 134.200 ;
        RECT 449.200 134.300 450.000 134.400 ;
        RECT 452.400 134.300 455.800 134.400 ;
        RECT 449.200 133.800 455.800 134.300 ;
        RECT 441.400 133.600 443.000 133.800 ;
        RECT 449.200 133.700 454.000 133.800 ;
        RECT 449.200 133.600 450.000 133.700 ;
        RECT 452.400 133.600 454.000 133.700 ;
        RECT 441.400 130.400 442.000 133.600 ;
        RECT 443.600 131.600 445.200 132.400 ;
        RECT 428.400 129.600 429.800 130.200 ;
        RECT 430.400 129.600 431.400 130.200 ;
        RECT 429.200 128.400 429.800 129.600 ;
        RECT 429.200 127.600 430.000 128.400 ;
        RECT 430.600 124.400 431.400 129.600 ;
        RECT 434.800 129.600 437.400 130.200 ;
        RECT 430.600 123.600 432.400 124.400 ;
        RECT 430.600 122.200 431.400 123.600 ;
        RECT 434.800 122.200 435.600 129.600 ;
        RECT 438.000 129.200 439.000 130.200 ;
        RECT 441.200 129.600 442.000 130.400 ;
        RECT 444.400 130.300 445.200 130.400 ;
        RECT 446.000 130.300 446.800 131.200 ;
        RECT 444.400 129.700 446.800 130.300 ;
        RECT 449.400 130.200 450.000 133.600 ;
        RECT 456.400 133.400 457.200 134.200 ;
        RECT 456.400 132.800 457.000 133.400 ;
        RECT 450.800 130.800 451.600 132.400 ;
        RECT 454.400 132.200 457.000 132.800 ;
        RECT 457.800 132.800 458.400 136.200 ;
        RECT 462.000 135.800 462.800 139.800 ;
        RECT 459.000 134.800 459.800 135.600 ;
        RECT 460.400 135.200 462.800 135.800 ;
        RECT 460.400 135.000 461.200 135.200 ;
        RECT 459.200 134.400 459.800 134.800 ;
        RECT 459.200 133.600 460.000 134.400 ;
        RECT 461.200 134.300 462.800 134.400 ;
        RECT 468.400 134.300 469.200 139.800 ;
        RECT 473.200 137.800 474.000 139.800 ;
        RECT 470.000 135.600 470.800 137.200 ;
        RECT 471.600 135.600 472.400 137.200 ;
        RECT 473.400 136.400 474.000 137.800 ;
        RECT 473.200 135.600 474.000 136.400 ;
        RECT 476.400 136.000 477.200 139.800 ;
        RECT 479.600 136.000 480.400 139.800 ;
        RECT 476.400 135.800 480.400 136.000 ;
        RECT 481.200 135.800 482.000 139.800 ;
        RECT 484.400 136.400 485.200 139.800 ;
        RECT 484.200 135.800 485.200 136.400 ;
        RECT 471.700 134.300 472.300 135.600 ;
        RECT 473.400 134.400 474.000 135.600 ;
        RECT 476.600 135.400 480.200 135.800 ;
        RECT 477.200 134.400 478.000 134.800 ;
        RECT 481.200 134.400 481.800 135.800 ;
        RECT 484.200 134.400 484.800 135.800 ;
        RECT 487.600 135.200 488.400 139.800 ;
        RECT 489.200 135.800 490.000 139.800 ;
        RECT 490.800 136.000 491.600 139.800 ;
        RECT 494.000 136.000 494.800 139.800 ;
        RECT 499.400 136.000 500.200 139.000 ;
        RECT 503.600 137.000 504.400 139.000 ;
        RECT 490.800 135.800 494.800 136.000 ;
        RECT 485.800 134.600 488.400 135.200 ;
        RECT 461.200 133.700 472.300 134.300 ;
        RECT 461.200 133.600 462.800 133.700 ;
        RECT 457.800 132.400 458.800 132.800 ;
        RECT 457.800 132.200 459.600 132.400 ;
        RECT 454.400 132.000 455.200 132.200 ;
        RECT 458.200 131.600 459.600 132.200 ;
        RECT 456.600 131.400 457.400 131.600 ;
        RECT 454.000 130.800 457.400 131.400 ;
        RECT 454.000 130.200 454.600 130.800 ;
        RECT 458.200 130.200 458.800 131.600 ;
        RECT 444.400 129.600 445.200 129.700 ;
        RECT 446.000 129.600 446.800 129.700 ;
        RECT 438.000 122.200 438.800 129.200 ;
        RECT 441.400 127.000 442.000 129.600 ;
        RECT 449.200 129.400 451.000 130.200 ;
        RECT 442.800 127.600 443.600 129.200 ;
        RECT 441.400 126.400 445.000 127.000 ;
        RECT 441.400 126.200 442.000 126.400 ;
        RECT 441.200 122.200 442.000 126.200 ;
        RECT 444.400 126.200 445.000 126.400 ;
        RECT 444.400 122.200 445.200 126.200 ;
        RECT 450.200 122.200 451.000 129.400 ;
        RECT 452.400 129.600 454.600 130.200 ;
        RECT 452.400 122.200 453.200 129.600 ;
        RECT 453.800 129.400 454.600 129.600 ;
        RECT 456.800 129.600 458.800 130.200 ;
        RECT 460.400 129.600 462.800 130.200 ;
        RECT 456.800 122.200 458.400 129.600 ;
        RECT 460.400 129.400 461.200 129.600 ;
        RECT 462.000 122.200 462.800 129.600 ;
        RECT 468.400 122.200 469.200 133.700 ;
        RECT 473.200 133.600 474.000 134.400 ;
        RECT 476.400 133.800 478.000 134.400 ;
        RECT 476.400 133.600 477.200 133.800 ;
        RECT 479.400 133.600 482.000 134.400 ;
        RECT 482.800 134.300 483.600 134.400 ;
        RECT 484.200 134.300 485.200 134.400 ;
        RECT 482.800 133.700 485.200 134.300 ;
        RECT 482.800 133.600 483.600 133.700 ;
        RECT 484.200 133.600 485.200 133.700 ;
        RECT 473.400 130.200 474.000 133.600 ;
        RECT 474.800 130.800 475.600 132.400 ;
        RECT 478.000 131.600 478.800 133.200 ;
        RECT 479.400 132.300 480.000 133.600 ;
        RECT 482.800 132.300 483.600 132.400 ;
        RECT 479.400 131.700 483.600 132.300 ;
        RECT 479.400 130.200 480.000 131.700 ;
        RECT 482.800 131.600 483.600 131.700 ;
        RECT 481.200 130.200 482.000 130.400 ;
        RECT 473.200 129.400 475.000 130.200 ;
        RECT 474.200 122.200 475.000 129.400 ;
        RECT 479.000 129.600 480.000 130.200 ;
        RECT 480.600 129.600 482.000 130.200 ;
        RECT 484.200 130.200 484.800 133.600 ;
        RECT 485.800 133.000 486.400 134.600 ;
        RECT 489.400 134.400 490.000 135.800 ;
        RECT 491.000 135.400 494.600 135.800 ;
        RECT 498.600 135.400 500.200 136.000 ;
        RECT 498.600 135.000 499.400 135.400 ;
        RECT 493.200 134.400 494.000 134.800 ;
        RECT 498.600 134.400 499.200 135.000 ;
        RECT 503.800 134.800 504.400 137.000 ;
        RECT 506.800 136.400 507.600 139.800 ;
        RECT 489.200 133.600 491.800 134.400 ;
        RECT 493.200 133.800 494.800 134.400 ;
        RECT 497.200 134.300 499.200 134.400 ;
        RECT 494.000 133.600 494.800 133.800 ;
        RECT 495.700 133.700 499.200 134.300 ;
        RECT 500.200 134.200 504.400 134.800 ;
        RECT 506.600 135.800 507.600 136.400 ;
        RECT 506.600 134.400 507.200 135.800 ;
        RECT 510.000 135.200 510.800 139.800 ;
        RECT 511.600 136.000 512.400 139.800 ;
        RECT 514.800 136.000 515.600 139.800 ;
        RECT 511.600 135.800 515.600 136.000 ;
        RECT 516.400 135.800 517.200 139.800 ;
        RECT 511.800 135.400 515.400 135.800 ;
        RECT 508.200 134.600 510.800 135.200 ;
        RECT 500.200 133.800 501.200 134.200 ;
        RECT 485.400 132.200 486.400 133.000 ;
        RECT 485.800 130.200 486.400 132.200 ;
        RECT 487.400 132.400 488.200 133.200 ;
        RECT 487.400 131.600 488.400 132.400 ;
        RECT 491.200 130.400 491.800 133.600 ;
        RECT 492.400 132.300 493.200 133.200 ;
        RECT 495.700 132.300 496.300 133.700 ;
        RECT 497.200 133.600 499.200 133.700 ;
        RECT 492.400 131.700 496.300 132.300 ;
        RECT 492.400 131.600 493.200 131.700 ;
        RECT 497.200 130.800 498.000 132.400 ;
        RECT 489.200 130.200 490.000 130.400 ;
        RECT 479.000 122.200 479.800 129.600 ;
        RECT 480.600 128.400 481.200 129.600 ;
        RECT 484.200 129.200 485.200 130.200 ;
        RECT 485.800 129.600 488.400 130.200 ;
        RECT 489.200 129.600 490.600 130.200 ;
        RECT 491.200 129.600 493.200 130.400 ;
        RECT 498.600 129.800 499.200 133.600 ;
        RECT 499.800 133.000 501.200 133.800 ;
        RECT 506.600 133.600 507.600 134.400 ;
        RECT 500.600 131.000 501.200 133.000 ;
        RECT 502.000 131.600 502.800 133.200 ;
        RECT 503.600 131.600 504.400 133.200 ;
        RECT 500.600 130.400 504.400 131.000 ;
        RECT 480.400 127.600 481.200 128.400 ;
        RECT 484.400 122.200 485.200 129.200 ;
        RECT 487.600 122.200 488.400 129.600 ;
        RECT 490.000 128.400 490.600 129.600 ;
        RECT 490.000 127.600 490.800 128.400 ;
        RECT 491.400 122.200 492.200 129.600 ;
        RECT 498.600 129.200 500.200 129.800 ;
        RECT 499.400 122.200 500.200 129.200 ;
        RECT 503.800 127.000 504.400 130.400 ;
        RECT 506.600 130.200 507.200 133.600 ;
        RECT 508.200 133.000 508.800 134.600 ;
        RECT 512.400 134.400 513.200 134.800 ;
        RECT 516.400 134.400 517.000 135.800 ;
        RECT 518.000 135.400 518.800 139.800 ;
        RECT 522.200 138.400 523.400 139.800 ;
        RECT 522.200 137.800 523.600 138.400 ;
        RECT 526.800 137.800 527.600 139.800 ;
        RECT 531.200 138.400 532.000 139.800 ;
        RECT 531.200 137.800 533.200 138.400 ;
        RECT 522.800 137.000 523.600 137.800 ;
        RECT 527.000 137.200 527.600 137.800 ;
        RECT 527.000 136.600 529.800 137.200 ;
        RECT 529.000 136.400 529.800 136.600 ;
        RECT 530.800 136.400 531.600 137.200 ;
        RECT 532.400 137.000 533.200 137.800 ;
        RECT 521.000 135.400 521.800 135.600 ;
        RECT 518.000 134.800 521.800 135.400 ;
        RECT 511.600 133.800 513.200 134.400 ;
        RECT 511.600 133.600 512.400 133.800 ;
        RECT 514.600 133.600 517.200 134.400 ;
        RECT 507.800 132.200 508.800 133.000 ;
        RECT 508.200 130.200 508.800 132.200 ;
        RECT 509.800 132.400 510.600 133.200 ;
        RECT 509.800 131.600 510.800 132.400 ;
        RECT 513.200 131.600 514.000 133.200 ;
        RECT 514.600 132.400 515.200 133.600 ;
        RECT 514.600 131.600 515.600 132.400 ;
        RECT 514.600 130.200 515.200 131.600 ;
        RECT 518.000 131.400 518.800 134.800 ;
        RECT 525.000 134.200 525.800 134.400 ;
        RECT 529.200 134.200 530.000 134.400 ;
        RECT 530.800 134.200 531.400 136.400 ;
        RECT 535.600 135.000 536.400 139.800 ;
        RECT 537.200 136.000 538.000 139.800 ;
        RECT 540.400 136.000 541.200 139.800 ;
        RECT 537.200 135.800 541.200 136.000 ;
        RECT 542.000 135.800 542.800 139.800 ;
        RECT 537.400 135.400 541.000 135.800 ;
        RECT 538.000 134.400 538.800 134.800 ;
        RECT 542.000 134.400 542.600 135.800 ;
        RECT 534.000 134.200 535.600 134.400 ;
        RECT 524.600 133.600 535.600 134.200 ;
        RECT 537.200 133.800 538.800 134.400 ;
        RECT 537.200 133.600 538.000 133.800 ;
        RECT 540.200 133.600 542.800 134.400 ;
        RECT 522.800 132.800 523.600 133.000 ;
        RECT 519.800 132.200 523.600 132.800 ;
        RECT 519.800 132.000 520.600 132.200 ;
        RECT 521.400 131.400 522.200 131.600 ;
        RECT 518.000 130.800 522.200 131.400 ;
        RECT 516.400 130.200 517.200 130.400 ;
        RECT 506.600 129.200 507.600 130.200 ;
        RECT 508.200 129.600 510.800 130.200 ;
        RECT 503.600 123.000 504.400 127.000 ;
        RECT 506.800 122.200 507.600 129.200 ;
        RECT 510.000 122.200 510.800 129.600 ;
        RECT 514.200 129.600 515.200 130.200 ;
        RECT 515.800 129.600 517.200 130.200 ;
        RECT 514.200 122.200 515.000 129.600 ;
        RECT 515.800 128.400 516.400 129.600 ;
        RECT 515.600 127.600 516.400 128.400 ;
        RECT 518.000 122.200 518.800 130.800 ;
        RECT 524.600 130.400 525.200 133.600 ;
        RECT 531.800 133.400 532.600 133.600 ;
        RECT 533.400 132.400 534.200 132.600 ;
        RECT 529.200 131.800 534.200 132.400 ;
        RECT 529.200 131.600 530.000 131.800 ;
        RECT 538.800 131.600 539.600 133.200 ;
        RECT 540.200 132.400 540.800 133.600 ;
        RECT 540.200 131.600 541.200 132.400 ;
        RECT 530.800 131.000 536.400 131.200 ;
        RECT 530.600 130.800 536.400 131.000 ;
        RECT 522.800 129.800 525.200 130.400 ;
        RECT 526.600 130.600 536.400 130.800 ;
        RECT 526.600 130.200 531.400 130.600 ;
        RECT 522.800 128.800 523.400 129.800 ;
        RECT 522.000 128.000 523.400 128.800 ;
        RECT 525.000 129.000 525.800 129.200 ;
        RECT 526.600 129.000 527.200 130.200 ;
        RECT 525.000 128.400 527.200 129.000 ;
        RECT 527.800 129.000 533.200 129.600 ;
        RECT 527.800 128.800 528.600 129.000 ;
        RECT 532.400 128.800 533.200 129.000 ;
        RECT 526.200 127.400 527.000 127.600 ;
        RECT 529.000 127.400 529.800 127.600 ;
        RECT 522.800 126.200 523.600 127.000 ;
        RECT 526.200 126.800 529.800 127.400 ;
        RECT 527.000 126.200 527.600 126.800 ;
        RECT 532.400 126.200 533.200 127.000 ;
        RECT 522.200 122.200 523.400 126.200 ;
        RECT 526.800 122.200 527.600 126.200 ;
        RECT 531.200 125.600 533.200 126.200 ;
        RECT 531.200 122.200 532.000 125.600 ;
        RECT 535.600 122.200 536.400 130.600 ;
        RECT 540.200 130.200 540.800 131.600 ;
        RECT 542.000 130.300 542.800 130.400 ;
        RECT 543.600 130.300 544.400 139.800 ;
        RECT 545.200 135.600 546.000 137.200 ;
        RECT 546.800 135.200 547.600 139.800 ;
        RECT 550.000 136.400 550.800 139.800 ;
        RECT 550.000 135.800 551.000 136.400 ;
        RECT 546.800 134.600 549.400 135.200 ;
        RECT 547.000 132.400 547.800 133.200 ;
        RECT 546.800 131.600 547.800 132.400 ;
        RECT 548.800 133.000 549.400 134.600 ;
        RECT 550.400 134.400 551.000 135.800 ;
        RECT 553.200 135.200 554.000 139.800 ;
        RECT 556.400 136.400 557.200 139.800 ;
        RECT 556.400 135.600 557.400 136.400 ;
        RECT 553.200 134.600 555.800 135.200 ;
        RECT 550.000 134.300 551.000 134.400 ;
        RECT 551.600 134.300 552.400 134.400 ;
        RECT 550.000 133.700 552.400 134.300 ;
        RECT 550.000 133.600 551.000 133.700 ;
        RECT 551.600 133.600 552.400 133.700 ;
        RECT 548.800 132.200 549.800 133.000 ;
        RECT 542.000 130.200 544.400 130.300 ;
        RECT 548.800 130.200 549.400 132.200 ;
        RECT 550.400 130.200 551.000 133.600 ;
        RECT 553.400 132.400 554.200 133.200 ;
        RECT 553.200 131.600 554.200 132.400 ;
        RECT 555.200 133.000 555.800 134.600 ;
        RECT 556.800 134.400 557.400 135.600 ;
        RECT 556.400 133.600 557.400 134.400 ;
        RECT 555.200 132.200 556.200 133.000 ;
        RECT 555.200 130.200 555.800 132.200 ;
        RECT 556.800 130.200 557.400 133.600 ;
        RECT 539.800 129.600 540.800 130.200 ;
        RECT 541.400 129.700 544.400 130.200 ;
        RECT 541.400 129.600 542.800 129.700 ;
        RECT 539.800 122.200 540.600 129.600 ;
        RECT 541.400 128.400 542.000 129.600 ;
        RECT 541.200 127.600 542.000 128.400 ;
        RECT 543.600 122.200 544.400 129.700 ;
        RECT 546.800 129.600 549.400 130.200 ;
        RECT 546.800 122.200 547.600 129.600 ;
        RECT 550.000 129.200 551.000 130.200 ;
        RECT 553.200 129.600 555.800 130.200 ;
        RECT 550.000 122.200 550.800 129.200 ;
        RECT 553.200 122.200 554.000 129.600 ;
        RECT 556.400 129.200 557.400 130.200 ;
        RECT 556.400 122.200 557.200 129.200 ;
        RECT 559.600 122.200 560.400 139.800 ;
        RECT 561.200 135.600 562.000 137.200 ;
        RECT 562.800 136.000 563.600 139.800 ;
        RECT 566.000 136.000 566.800 139.800 ;
        RECT 562.800 135.800 566.800 136.000 ;
        RECT 567.600 135.800 568.400 139.800 ;
        RECT 569.200 137.000 570.000 139.000 ;
        RECT 563.000 135.400 566.600 135.800 ;
        RECT 563.600 134.400 564.400 134.800 ;
        RECT 567.600 134.400 568.200 135.800 ;
        RECT 569.200 134.800 569.800 137.000 ;
        RECT 573.400 136.000 574.200 139.000 ;
        RECT 578.800 136.000 579.600 139.800 ;
        RECT 582.000 136.000 582.800 139.800 ;
        RECT 573.400 135.400 575.000 136.000 ;
        RECT 578.800 135.800 582.800 136.000 ;
        RECT 583.600 135.800 584.400 139.800 ;
        RECT 585.800 138.400 586.600 139.800 ;
        RECT 585.200 137.600 586.600 138.400 ;
        RECT 585.800 136.400 586.600 137.600 ;
        RECT 585.800 135.800 587.600 136.400 ;
        RECT 579.000 135.400 582.600 135.800 ;
        RECT 574.200 135.000 575.000 135.400 ;
        RECT 562.800 133.800 564.400 134.400 ;
        RECT 562.800 133.600 563.600 133.800 ;
        RECT 565.800 133.600 568.400 134.400 ;
        RECT 569.200 134.200 573.400 134.800 ;
        RECT 572.400 133.800 573.400 134.200 ;
        RECT 574.400 134.400 575.000 135.000 ;
        RECT 579.600 134.400 580.400 134.800 ;
        RECT 583.600 134.400 584.200 135.800 ;
        RECT 574.400 134.300 576.400 134.400 ;
        RECT 564.400 131.600 565.200 133.200 ;
        RECT 565.800 132.300 566.400 133.600 ;
        RECT 567.600 132.300 568.400 132.400 ;
        RECT 565.800 131.700 568.400 132.300 ;
        RECT 565.800 130.200 566.400 131.700 ;
        RECT 567.600 131.600 568.400 131.700 ;
        RECT 569.200 131.600 570.000 133.200 ;
        RECT 570.800 131.600 571.600 133.200 ;
        RECT 572.400 133.000 573.800 133.800 ;
        RECT 574.400 133.700 577.900 134.300 ;
        RECT 574.400 133.600 576.400 133.700 ;
        RECT 572.400 131.000 573.000 133.000 ;
        RECT 569.200 130.400 573.000 131.000 ;
        RECT 567.600 130.200 568.400 130.400 ;
        RECT 565.400 129.600 566.400 130.200 ;
        RECT 567.000 129.600 568.400 130.200 ;
        RECT 565.400 122.200 566.200 129.600 ;
        RECT 567.000 128.400 567.600 129.600 ;
        RECT 566.800 127.600 567.600 128.400 ;
        RECT 569.200 127.000 569.800 130.400 ;
        RECT 574.400 129.800 575.000 133.600 ;
        RECT 575.600 130.800 576.400 132.400 ;
        RECT 577.300 132.300 577.900 133.700 ;
        RECT 578.800 133.800 580.400 134.400 ;
        RECT 578.800 133.600 579.600 133.800 ;
        RECT 581.800 133.600 584.400 134.400 ;
        RECT 580.400 132.300 581.200 133.200 ;
        RECT 577.300 131.700 581.200 132.300 ;
        RECT 580.400 131.600 581.200 131.700 ;
        RECT 581.800 132.300 582.400 133.600 ;
        RECT 585.200 132.300 586.000 132.400 ;
        RECT 581.800 131.700 586.000 132.300 ;
        RECT 581.800 130.200 582.400 131.700 ;
        RECT 585.200 131.600 586.000 131.700 ;
        RECT 583.600 130.200 584.400 130.400 ;
        RECT 573.400 129.200 575.000 129.800 ;
        RECT 581.400 129.600 582.400 130.200 ;
        RECT 583.000 129.600 584.400 130.200 ;
        RECT 569.200 123.000 570.000 127.000 ;
        RECT 573.400 122.200 574.200 129.200 ;
        RECT 581.400 122.200 582.200 129.600 ;
        RECT 583.000 128.400 583.600 129.600 ;
        RECT 582.800 127.600 583.600 128.400 ;
        RECT 585.200 127.600 586.000 130.400 ;
        RECT 586.800 122.200 587.600 135.800 ;
        RECT 588.400 133.600 589.200 135.200 ;
        RECT 590.000 135.000 590.800 139.800 ;
        RECT 594.400 138.400 595.200 139.800 ;
        RECT 593.200 137.800 595.200 138.400 ;
        RECT 598.800 137.800 599.600 139.800 ;
        RECT 603.000 138.400 604.200 139.800 ;
        RECT 602.800 137.800 604.200 138.400 ;
        RECT 593.200 137.000 594.000 137.800 ;
        RECT 598.800 137.200 599.400 137.800 ;
        RECT 594.800 136.400 595.600 137.200 ;
        RECT 596.600 136.600 599.400 137.200 ;
        RECT 602.800 137.000 603.600 137.800 ;
        RECT 596.600 136.400 597.400 136.600 ;
        RECT 590.800 134.200 592.400 134.400 ;
        RECT 595.000 134.200 595.600 136.400 ;
        RECT 604.600 135.400 605.400 135.600 ;
        RECT 607.600 135.400 608.400 139.800 ;
        RECT 604.600 134.800 608.400 135.400 ;
        RECT 600.600 134.200 601.400 134.400 ;
        RECT 590.800 133.600 601.800 134.200 ;
        RECT 593.800 133.400 594.600 133.600 ;
        RECT 592.200 132.400 593.000 132.600 ;
        RECT 594.800 132.400 595.600 132.600 ;
        RECT 592.200 131.800 597.200 132.400 ;
        RECT 596.400 131.600 597.200 131.800 ;
        RECT 590.000 131.000 595.600 131.200 ;
        RECT 590.000 130.800 595.800 131.000 ;
        RECT 590.000 130.600 599.800 130.800 ;
        RECT 590.000 122.200 590.800 130.600 ;
        RECT 595.000 130.200 599.800 130.600 ;
        RECT 593.200 129.000 598.600 129.600 ;
        RECT 593.200 128.800 594.000 129.000 ;
        RECT 597.800 128.800 598.600 129.000 ;
        RECT 599.200 129.000 599.800 130.200 ;
        RECT 601.200 130.400 601.800 133.600 ;
        RECT 602.800 132.800 603.600 133.000 ;
        RECT 602.800 132.200 606.600 132.800 ;
        RECT 605.800 132.000 606.600 132.200 ;
        RECT 604.200 131.400 605.000 131.600 ;
        RECT 607.600 131.400 608.400 134.800 ;
        RECT 604.200 130.800 608.400 131.400 ;
        RECT 601.200 129.800 603.600 130.400 ;
        RECT 600.600 129.000 601.400 129.200 ;
        RECT 599.200 128.400 601.400 129.000 ;
        RECT 603.000 128.800 603.600 129.800 ;
        RECT 603.000 128.000 604.400 128.800 ;
        RECT 596.600 127.400 597.400 127.600 ;
        RECT 599.400 127.400 600.200 127.600 ;
        RECT 593.200 126.200 594.000 127.000 ;
        RECT 596.600 126.800 600.200 127.400 ;
        RECT 598.800 126.200 599.400 126.800 ;
        RECT 602.800 126.200 603.600 127.000 ;
        RECT 593.200 125.600 595.200 126.200 ;
        RECT 594.400 122.200 595.200 125.600 ;
        RECT 598.800 122.200 599.600 126.200 ;
        RECT 603.000 122.200 604.200 126.200 ;
        RECT 607.600 122.200 608.400 130.800 ;
        RECT 1.200 111.400 2.000 119.800 ;
        RECT 5.600 116.400 6.400 119.800 ;
        RECT 4.400 115.800 6.400 116.400 ;
        RECT 10.000 115.800 10.800 119.800 ;
        RECT 14.200 115.800 15.400 119.800 ;
        RECT 4.400 115.000 5.200 115.800 ;
        RECT 10.000 115.200 10.600 115.800 ;
        RECT 7.800 114.600 11.400 115.200 ;
        RECT 14.000 115.000 14.800 115.800 ;
        RECT 7.800 114.400 8.600 114.600 ;
        RECT 10.600 114.400 11.400 114.600 ;
        RECT 4.400 113.000 5.200 113.200 ;
        RECT 9.000 113.000 9.800 113.200 ;
        RECT 4.400 112.400 9.800 113.000 ;
        RECT 10.400 113.000 12.600 113.600 ;
        RECT 10.400 111.800 11.000 113.000 ;
        RECT 11.800 112.800 12.600 113.000 ;
        RECT 14.200 113.200 15.600 114.000 ;
        RECT 14.200 112.200 14.800 113.200 ;
        RECT 6.200 111.400 11.000 111.800 ;
        RECT 1.200 111.200 11.000 111.400 ;
        RECT 12.400 111.600 14.800 112.200 ;
        RECT 1.200 111.000 7.000 111.200 ;
        RECT 1.200 110.800 6.800 111.000 ;
        RECT 7.600 110.300 8.400 110.400 ;
        RECT 9.200 110.300 10.000 110.400 ;
        RECT 7.600 110.200 10.000 110.300 ;
        RECT 3.400 109.700 10.000 110.200 ;
        RECT 3.400 109.600 8.400 109.700 ;
        RECT 9.200 109.600 10.000 109.700 ;
        RECT 3.400 109.400 4.200 109.600 ;
        RECT 5.000 108.400 5.800 108.600 ;
        RECT 12.400 108.400 13.000 111.600 ;
        RECT 18.800 111.200 19.600 119.800 ;
        RECT 21.200 113.600 22.000 114.400 ;
        RECT 21.200 112.400 21.800 113.600 ;
        RECT 22.600 112.400 23.400 119.800 ;
        RECT 27.600 113.600 28.400 114.400 ;
        RECT 27.600 112.400 28.200 113.600 ;
        RECT 29.000 112.400 29.800 119.800 ;
        RECT 34.800 112.800 35.600 119.800 ;
        RECT 20.400 111.800 21.800 112.400 ;
        RECT 22.400 111.800 23.400 112.400 ;
        RECT 26.800 111.800 28.200 112.400 ;
        RECT 28.800 111.800 29.800 112.400 ;
        RECT 34.600 111.800 35.600 112.800 ;
        RECT 38.000 112.400 38.800 119.800 ;
        RECT 43.400 118.400 44.200 119.800 ;
        RECT 42.800 117.600 44.200 118.400 ;
        RECT 43.400 112.800 44.200 117.600 ;
        RECT 47.600 115.000 48.400 119.000 ;
        RECT 36.200 111.800 38.800 112.400 ;
        RECT 42.600 112.200 44.200 112.800 ;
        RECT 20.400 111.600 21.200 111.800 ;
        RECT 15.400 110.600 19.600 111.200 ;
        RECT 15.400 110.400 16.200 110.600 ;
        RECT 17.000 109.800 17.800 110.000 ;
        RECT 14.000 109.200 17.800 109.800 ;
        RECT 14.000 109.000 14.800 109.200 ;
        RECT 2.000 107.800 13.000 108.400 ;
        RECT 2.000 107.600 3.600 107.800 ;
        RECT 6.000 107.600 6.800 107.800 ;
        RECT 11.800 107.600 12.600 107.800 ;
        RECT 1.200 102.200 2.000 107.000 ;
        RECT 6.200 105.600 6.800 107.600 ;
        RECT 18.800 107.200 19.600 110.600 ;
        RECT 22.400 110.400 23.000 111.800 ;
        RECT 26.800 111.600 27.600 111.800 ;
        RECT 22.000 109.600 23.000 110.400 ;
        RECT 22.400 108.400 23.000 109.600 ;
        RECT 23.600 108.800 24.400 110.400 ;
        RECT 28.800 108.400 29.400 111.800 ;
        RECT 30.000 108.800 30.800 110.400 ;
        RECT 34.600 108.400 35.200 111.800 ;
        RECT 36.200 109.800 36.800 111.800 ;
        RECT 35.800 109.000 36.800 109.800 ;
        RECT 20.400 107.600 23.000 108.400 ;
        RECT 25.200 108.200 26.000 108.400 ;
        RECT 24.400 107.600 26.000 108.200 ;
        RECT 26.800 107.600 29.400 108.400 ;
        RECT 31.600 108.300 32.400 108.400 ;
        RECT 34.600 108.300 35.600 108.400 ;
        RECT 31.600 108.200 35.600 108.300 ;
        RECT 30.800 107.700 35.600 108.200 ;
        RECT 30.800 107.600 32.400 107.700 ;
        RECT 34.600 107.600 35.600 107.700 ;
        RECT 15.800 106.600 19.600 107.200 ;
        RECT 15.800 106.400 16.600 106.600 ;
        RECT 4.400 104.200 5.200 105.000 ;
        RECT 6.000 104.800 6.800 105.600 ;
        RECT 7.800 105.400 8.600 105.600 ;
        RECT 7.800 104.800 10.600 105.400 ;
        RECT 10.000 104.200 10.600 104.800 ;
        RECT 14.000 104.200 14.800 105.000 ;
        RECT 4.400 103.600 6.400 104.200 ;
        RECT 5.600 102.200 6.400 103.600 ;
        RECT 10.000 102.200 10.800 104.200 ;
        RECT 14.000 103.600 15.400 104.200 ;
        RECT 14.200 102.200 15.400 103.600 ;
        RECT 18.800 102.200 19.600 106.600 ;
        RECT 20.600 106.200 21.200 107.600 ;
        RECT 24.400 107.200 25.200 107.600 ;
        RECT 22.200 106.200 25.800 106.600 ;
        RECT 27.000 106.200 27.600 107.600 ;
        RECT 30.800 107.200 31.600 107.600 ;
        RECT 28.600 106.200 32.200 106.600 ;
        RECT 34.600 106.200 35.200 107.600 ;
        RECT 36.200 107.400 36.800 109.000 ;
        RECT 37.800 109.600 38.800 110.400 ;
        RECT 39.600 110.300 40.400 110.400 ;
        RECT 41.200 110.300 42.000 111.200 ;
        RECT 39.600 109.700 42.000 110.300 ;
        RECT 39.600 109.600 40.400 109.700 ;
        RECT 41.200 109.600 42.000 109.700 ;
        RECT 37.800 108.800 38.600 109.600 ;
        RECT 42.600 108.400 43.200 112.200 ;
        RECT 47.800 111.600 48.400 115.000 ;
        RECT 51.800 112.400 52.600 119.800 ;
        RECT 53.200 113.600 54.000 114.400 ;
        RECT 53.400 112.400 54.000 113.600 ;
        RECT 56.400 113.600 57.200 114.400 ;
        RECT 56.400 112.400 57.000 113.600 ;
        RECT 57.800 112.400 58.600 119.800 ;
        RECT 65.800 112.800 66.600 119.800 ;
        RECT 70.000 115.000 70.800 119.000 ;
        RECT 51.800 111.800 52.800 112.400 ;
        RECT 53.400 111.800 54.800 112.400 ;
        RECT 44.600 111.000 48.400 111.600 ;
        RECT 44.600 109.000 45.200 111.000 ;
        RECT 41.200 107.600 43.200 108.400 ;
        RECT 43.800 108.200 45.200 109.000 ;
        RECT 46.000 108.800 46.800 110.400 ;
        RECT 47.600 108.800 48.400 110.400 ;
        RECT 50.800 108.800 51.600 110.400 ;
        RECT 52.200 110.300 52.800 111.800 ;
        RECT 54.000 111.600 54.800 111.800 ;
        RECT 55.600 111.800 57.000 112.400 ;
        RECT 57.600 111.800 58.600 112.400 ;
        RECT 65.000 112.200 66.600 112.800 ;
        RECT 55.600 111.600 56.400 111.800 ;
        RECT 55.700 110.300 56.300 111.600 ;
        RECT 57.600 110.400 58.200 111.800 ;
        RECT 52.200 109.700 56.300 110.300 ;
        RECT 52.200 108.400 52.800 109.700 ;
        RECT 57.200 109.600 58.200 110.400 ;
        RECT 57.600 108.400 58.200 109.600 ;
        RECT 58.800 110.300 59.600 110.400 ;
        RECT 58.800 109.700 62.700 110.300 ;
        RECT 58.800 108.800 59.600 109.700 ;
        RECT 36.200 106.800 38.800 107.400 ;
        RECT 20.400 102.200 21.200 106.200 ;
        RECT 22.000 106.000 26.000 106.200 ;
        RECT 22.000 102.200 22.800 106.000 ;
        RECT 25.200 102.200 26.000 106.000 ;
        RECT 26.800 102.200 27.600 106.200 ;
        RECT 28.400 106.000 32.400 106.200 ;
        RECT 28.400 102.200 29.200 106.000 ;
        RECT 31.600 102.200 32.400 106.000 ;
        RECT 34.600 105.600 35.600 106.200 ;
        RECT 34.800 102.200 35.600 105.600 ;
        RECT 38.000 102.200 38.800 106.800 ;
        RECT 42.600 107.000 43.200 107.600 ;
        RECT 44.200 107.800 45.200 108.200 ;
        RECT 49.200 108.200 50.000 108.400 ;
        RECT 44.200 107.200 48.400 107.800 ;
        RECT 49.200 107.600 50.800 108.200 ;
        RECT 52.200 107.600 54.800 108.400 ;
        RECT 55.600 107.600 58.200 108.400 ;
        RECT 60.400 108.200 61.200 108.400 ;
        RECT 59.600 107.600 61.200 108.200 ;
        RECT 62.100 108.300 62.700 109.700 ;
        RECT 63.600 109.600 64.400 111.200 ;
        RECT 65.000 108.400 65.600 112.200 ;
        RECT 70.200 111.600 70.800 115.000 ;
        RECT 73.200 112.800 74.000 119.800 ;
        RECT 67.000 111.000 70.800 111.600 ;
        RECT 73.000 111.600 74.000 112.800 ;
        RECT 76.400 112.400 77.200 119.800 ;
        RECT 79.600 112.800 80.400 119.800 ;
        RECT 74.600 111.800 77.200 112.400 ;
        RECT 79.400 111.800 80.400 112.800 ;
        RECT 82.800 112.400 83.600 119.800 ;
        RECT 81.000 111.800 83.600 112.400 ;
        RECT 67.000 109.000 67.600 111.000 ;
        RECT 63.600 108.300 65.600 108.400 ;
        RECT 62.100 107.700 65.600 108.300 ;
        RECT 66.200 108.200 67.600 109.000 ;
        RECT 68.400 108.800 69.200 110.400 ;
        RECT 70.000 108.800 70.800 110.400 ;
        RECT 63.600 107.600 65.600 107.700 ;
        RECT 50.000 107.200 50.800 107.600 ;
        RECT 42.600 106.600 43.400 107.000 ;
        RECT 42.600 106.000 44.200 106.600 ;
        RECT 43.400 103.000 44.200 106.000 ;
        RECT 47.800 105.000 48.400 107.200 ;
        RECT 49.400 106.200 53.000 106.600 ;
        RECT 54.000 106.200 54.600 107.600 ;
        RECT 55.800 106.200 56.400 107.600 ;
        RECT 59.600 107.200 60.400 107.600 ;
        RECT 65.000 107.000 65.600 107.600 ;
        RECT 66.600 107.800 67.600 108.200 ;
        RECT 73.000 108.400 73.600 111.600 ;
        RECT 74.600 109.800 75.200 111.800 ;
        RECT 74.200 109.000 75.200 109.800 ;
        RECT 66.600 107.200 70.800 107.800 ;
        RECT 65.000 106.600 65.800 107.000 ;
        RECT 57.400 106.200 61.000 106.600 ;
        RECT 47.600 103.000 48.400 105.000 ;
        RECT 49.200 106.000 53.200 106.200 ;
        RECT 49.200 102.200 50.000 106.000 ;
        RECT 52.400 102.200 53.200 106.000 ;
        RECT 54.000 102.200 54.800 106.200 ;
        RECT 55.600 102.200 56.400 106.200 ;
        RECT 57.200 106.000 61.200 106.200 ;
        RECT 65.000 106.000 66.600 106.600 ;
        RECT 57.200 102.200 58.000 106.000 ;
        RECT 60.400 102.200 61.200 106.000 ;
        RECT 65.800 103.000 66.600 106.000 ;
        RECT 70.200 105.000 70.800 107.200 ;
        RECT 73.000 107.600 74.000 108.400 ;
        RECT 73.000 106.200 73.600 107.600 ;
        RECT 74.600 107.400 75.200 109.000 ;
        RECT 76.200 110.300 77.200 110.400 ;
        RECT 78.000 110.300 78.800 110.400 ;
        RECT 76.200 109.700 78.800 110.300 ;
        RECT 76.200 109.600 77.200 109.700 ;
        RECT 78.000 109.600 78.800 109.700 ;
        RECT 76.200 108.800 77.000 109.600 ;
        RECT 79.400 108.400 80.000 111.800 ;
        RECT 81.000 109.800 81.600 111.800 ;
        RECT 80.600 109.000 81.600 109.800 ;
        RECT 79.400 107.600 80.400 108.400 ;
        RECT 74.600 106.800 77.200 107.400 ;
        RECT 73.000 105.600 74.000 106.200 ;
        RECT 70.000 103.000 70.800 105.000 ;
        RECT 73.200 102.200 74.000 105.600 ;
        RECT 76.400 102.200 77.200 106.800 ;
        RECT 79.400 106.200 80.000 107.600 ;
        RECT 81.000 107.400 81.600 109.000 ;
        RECT 82.600 109.600 83.600 110.400 ;
        RECT 82.600 108.800 83.400 109.600 ;
        RECT 81.000 106.800 83.600 107.400 ;
        RECT 84.400 106.800 85.200 108.400 ;
        RECT 79.400 105.600 80.400 106.200 ;
        RECT 79.600 102.200 80.400 105.600 ;
        RECT 82.800 102.200 83.600 106.800 ;
        RECT 86.000 106.200 86.800 119.800 ;
        RECT 90.800 115.800 91.600 119.800 ;
        RECT 91.000 115.600 91.600 115.800 ;
        RECT 94.000 115.800 94.800 119.800 ;
        RECT 94.000 115.600 94.600 115.800 ;
        RECT 91.000 115.000 94.600 115.600 ;
        RECT 87.600 111.600 88.400 113.200 ;
        RECT 92.400 112.800 93.200 114.400 ;
        RECT 94.000 112.400 94.600 115.000 ;
        RECT 96.400 113.600 97.200 114.400 ;
        RECT 96.400 112.400 97.000 113.600 ;
        RECT 97.800 112.400 98.600 119.800 ;
        RECT 104.600 118.400 105.400 119.800 ;
        RECT 103.600 117.600 105.400 118.400 ;
        RECT 104.600 112.400 105.400 117.600 ;
        RECT 106.000 113.600 106.800 114.400 ;
        RECT 106.200 112.400 106.800 113.600 ;
        RECT 111.000 112.400 111.800 119.800 ;
        RECT 112.400 113.600 113.200 114.400 ;
        RECT 112.600 112.400 113.200 113.600 ;
        RECT 117.400 112.400 118.200 119.800 ;
        RECT 118.800 113.600 119.600 114.400 ;
        RECT 119.000 112.400 119.600 113.600 ;
        RECT 121.200 112.400 122.000 119.800 ;
        RECT 124.400 112.800 125.200 119.800 ;
        RECT 89.200 110.800 90.000 112.400 ;
        RECT 94.000 111.600 94.800 112.400 ;
        RECT 95.600 111.800 97.000 112.400 ;
        RECT 95.600 111.600 96.400 111.800 ;
        RECT 97.600 111.600 99.600 112.400 ;
        RECT 104.600 111.800 105.600 112.400 ;
        RECT 106.200 111.800 107.600 112.400 ;
        RECT 111.000 111.800 112.000 112.400 ;
        RECT 112.600 111.800 114.000 112.400 ;
        RECT 117.400 111.800 118.400 112.400 ;
        RECT 119.000 111.800 120.400 112.400 ;
        RECT 121.200 111.800 123.800 112.400 ;
        RECT 124.400 111.800 125.400 112.800 ;
        RECT 90.800 109.600 92.400 110.400 ;
        RECT 94.000 108.400 94.600 111.600 ;
        RECT 97.600 108.400 98.200 111.600 ;
        RECT 98.800 108.800 99.600 110.400 ;
        RECT 100.400 110.300 101.200 110.400 ;
        RECT 103.600 110.300 104.400 110.400 ;
        RECT 100.400 109.700 104.400 110.300 ;
        RECT 100.400 109.600 101.200 109.700 ;
        RECT 103.600 108.800 104.400 109.700 ;
        RECT 105.000 108.400 105.600 111.800 ;
        RECT 106.800 111.600 107.600 111.800 ;
        RECT 110.000 108.800 110.800 110.400 ;
        RECT 111.400 110.300 112.000 111.800 ;
        RECT 113.200 111.600 114.000 111.800 ;
        RECT 117.800 110.400 118.400 111.800 ;
        RECT 119.600 111.600 120.400 111.800 ;
        RECT 116.400 110.300 117.200 110.400 ;
        RECT 111.400 109.700 117.200 110.300 ;
        RECT 111.400 108.400 112.000 109.700 ;
        RECT 116.400 108.800 117.200 109.700 ;
        RECT 117.800 109.600 118.800 110.400 ;
        RECT 121.200 109.600 122.200 110.400 ;
        RECT 117.800 108.400 118.400 109.600 ;
        RECT 121.400 108.800 122.200 109.600 ;
        RECT 123.200 109.800 123.800 111.800 ;
        RECT 123.200 109.000 124.200 109.800 ;
        RECT 93.000 108.200 94.600 108.400 ;
        RECT 92.800 107.800 94.600 108.200 ;
        RECT 86.000 105.600 87.800 106.200 ;
        RECT 87.000 102.200 87.800 105.600 ;
        RECT 92.800 102.200 93.600 107.800 ;
        RECT 95.600 107.600 98.200 108.400 ;
        RECT 100.400 108.200 101.200 108.400 ;
        RECT 99.600 107.600 101.200 108.200 ;
        RECT 102.000 108.200 102.800 108.400 ;
        RECT 102.000 107.600 103.600 108.200 ;
        RECT 105.000 107.600 107.600 108.400 ;
        RECT 108.400 108.200 109.200 108.400 ;
        RECT 108.400 107.600 110.000 108.200 ;
        RECT 111.400 107.600 114.000 108.400 ;
        RECT 114.800 108.200 115.600 108.400 ;
        RECT 114.800 107.600 116.400 108.200 ;
        RECT 117.800 107.600 120.400 108.400 ;
        RECT 95.800 106.200 96.400 107.600 ;
        RECT 99.600 107.200 100.400 107.600 ;
        RECT 102.800 107.200 103.600 107.600 ;
        RECT 97.400 106.200 101.000 106.600 ;
        RECT 102.200 106.200 105.800 106.600 ;
        RECT 106.800 106.200 107.400 107.600 ;
        RECT 109.200 107.200 110.000 107.600 ;
        RECT 108.600 106.200 112.200 106.600 ;
        RECT 113.200 106.200 113.800 107.600 ;
        RECT 115.600 107.200 116.400 107.600 ;
        RECT 115.000 106.200 118.600 106.600 ;
        RECT 119.600 106.200 120.200 107.600 ;
        RECT 123.200 107.400 123.800 109.000 ;
        RECT 124.800 108.400 125.400 111.800 ;
        RECT 127.600 111.600 128.400 113.200 ;
        RECT 124.400 107.600 125.400 108.400 ;
        RECT 121.200 106.800 123.800 107.400 ;
        RECT 95.600 102.200 96.400 106.200 ;
        RECT 97.200 106.000 101.200 106.200 ;
        RECT 97.200 102.200 98.000 106.000 ;
        RECT 100.400 102.200 101.200 106.000 ;
        RECT 102.000 106.000 106.000 106.200 ;
        RECT 102.000 102.200 102.800 106.000 ;
        RECT 105.200 102.200 106.000 106.000 ;
        RECT 106.800 102.200 107.600 106.200 ;
        RECT 108.400 106.000 112.400 106.200 ;
        RECT 108.400 102.200 109.200 106.000 ;
        RECT 111.600 102.200 112.400 106.000 ;
        RECT 113.200 102.200 114.000 106.200 ;
        RECT 114.800 106.000 118.800 106.200 ;
        RECT 114.800 102.200 115.600 106.000 ;
        RECT 118.000 102.200 118.800 106.000 ;
        RECT 119.600 102.200 120.400 106.200 ;
        RECT 121.200 102.200 122.000 106.800 ;
        RECT 124.800 106.400 125.400 107.600 ;
        RECT 124.400 105.600 125.400 106.400 ;
        RECT 129.200 106.200 130.000 119.800 ;
        RECT 130.800 108.300 131.600 108.400 ;
        RECT 132.400 108.300 133.200 108.400 ;
        RECT 130.800 107.700 133.200 108.300 ;
        RECT 130.800 106.800 131.600 107.700 ;
        RECT 132.400 107.600 133.200 107.700 ;
        RECT 132.500 106.400 133.100 107.600 ;
        RECT 128.200 105.600 130.000 106.200 ;
        RECT 124.400 102.200 125.200 105.600 ;
        RECT 128.200 104.400 129.000 105.600 ;
        RECT 132.400 104.800 133.200 106.400 ;
        RECT 128.200 103.600 130.000 104.400 ;
        RECT 128.200 102.200 129.000 103.600 ;
        RECT 134.000 102.200 134.800 119.800 ;
        RECT 136.400 113.600 137.200 114.400 ;
        RECT 136.400 112.400 137.000 113.600 ;
        RECT 137.800 112.400 138.600 119.800 ;
        RECT 142.800 113.600 143.600 114.400 ;
        RECT 142.800 112.400 143.400 113.600 ;
        RECT 144.200 112.400 145.000 119.800 ;
        RECT 155.400 118.400 156.200 119.800 ;
        RECT 155.400 117.600 157.200 118.400 ;
        RECT 154.000 113.600 154.800 114.400 ;
        RECT 154.000 112.400 154.600 113.600 ;
        RECT 155.400 112.400 156.200 117.600 ;
        RECT 135.600 111.800 137.000 112.400 ;
        RECT 137.600 111.800 138.600 112.400 ;
        RECT 142.000 111.800 143.400 112.400 ;
        RECT 144.000 111.800 145.000 112.400 ;
        RECT 153.200 111.800 154.600 112.400 ;
        RECT 155.200 111.800 156.200 112.400 ;
        RECT 135.600 111.600 136.400 111.800 ;
        RECT 137.600 108.400 138.200 111.800 ;
        RECT 142.000 111.600 142.800 111.800 ;
        RECT 138.800 110.300 139.600 110.400 ;
        RECT 140.400 110.300 141.200 110.400 ;
        RECT 138.800 109.700 141.200 110.300 ;
        RECT 138.800 108.800 139.600 109.700 ;
        RECT 140.400 109.600 141.200 109.700 ;
        RECT 142.000 110.300 142.800 110.400 ;
        RECT 144.000 110.300 144.600 111.800 ;
        RECT 153.200 111.600 154.000 111.800 ;
        RECT 142.000 109.700 144.600 110.300 ;
        RECT 142.000 109.600 142.800 109.700 ;
        RECT 144.000 108.400 144.600 109.700 ;
        RECT 145.200 108.800 146.000 110.400 ;
        RECT 155.200 108.400 155.800 111.800 ;
        RECT 161.200 111.200 162.000 119.800 ;
        RECT 164.400 111.200 165.200 119.800 ;
        RECT 167.600 111.200 168.400 119.800 ;
        RECT 170.800 111.200 171.600 119.800 ;
        RECT 174.000 115.000 174.800 119.000 ;
        RECT 174.000 111.600 174.600 115.000 ;
        RECT 178.200 112.800 179.000 119.800 ;
        RECT 183.600 115.000 184.400 119.000 ;
        RECT 178.200 112.200 179.800 112.800 ;
        RECT 161.200 110.400 163.000 111.200 ;
        RECT 164.400 110.400 166.600 111.200 ;
        RECT 167.600 110.400 169.800 111.200 ;
        RECT 170.800 110.400 173.200 111.200 ;
        RECT 174.000 111.000 177.800 111.600 ;
        RECT 156.400 110.300 157.200 110.400 ;
        RECT 158.000 110.300 158.800 110.400 ;
        RECT 156.400 109.700 158.800 110.300 ;
        RECT 156.400 108.800 157.200 109.700 ;
        RECT 158.000 109.600 158.800 109.700 ;
        RECT 162.200 109.000 163.000 110.400 ;
        RECT 165.800 109.000 166.600 110.400 ;
        RECT 169.000 109.000 169.800 110.400 ;
        RECT 135.600 107.600 138.200 108.400 ;
        RECT 140.400 108.200 141.200 108.400 ;
        RECT 139.600 107.600 141.200 108.200 ;
        RECT 142.000 107.600 144.600 108.400 ;
        RECT 146.800 108.200 147.600 108.400 ;
        RECT 146.000 107.600 147.600 108.200 ;
        RECT 153.200 107.600 155.800 108.400 ;
        RECT 158.000 108.200 158.800 108.400 ;
        RECT 157.200 107.600 158.800 108.200 ;
        RECT 159.600 108.200 161.400 109.000 ;
        RECT 162.200 108.200 164.800 109.000 ;
        RECT 165.800 108.200 168.200 109.000 ;
        RECT 169.000 108.200 171.600 109.000 ;
        RECT 159.600 107.600 160.400 108.200 ;
        RECT 162.200 107.600 163.000 108.200 ;
        RECT 165.800 107.600 166.600 108.200 ;
        RECT 169.000 107.600 169.800 108.200 ;
        RECT 172.400 107.600 173.200 110.400 ;
        RECT 174.000 108.800 174.800 110.400 ;
        RECT 175.600 108.800 176.400 110.400 ;
        RECT 177.200 109.000 177.800 111.000 ;
        RECT 177.200 108.200 178.600 109.000 ;
        RECT 179.200 108.400 179.800 112.200 ;
        RECT 183.600 111.600 184.200 115.000 ;
        RECT 187.800 112.800 188.600 119.800 ;
        RECT 187.800 112.200 189.400 112.800 ;
        RECT 180.400 109.600 181.200 111.200 ;
        RECT 183.600 111.000 187.400 111.600 ;
        RECT 183.600 108.800 184.400 110.400 ;
        RECT 185.200 108.800 186.000 110.400 ;
        RECT 186.800 109.000 187.400 111.000 ;
        RECT 177.200 107.800 178.200 108.200 ;
        RECT 135.800 106.200 136.400 107.600 ;
        RECT 139.600 107.200 140.400 107.600 ;
        RECT 137.400 106.200 141.000 106.600 ;
        RECT 142.200 106.200 142.800 107.600 ;
        RECT 146.000 107.200 146.800 107.600 ;
        RECT 143.800 106.200 147.400 106.600 ;
        RECT 153.400 106.200 154.000 107.600 ;
        RECT 157.200 107.200 158.000 107.600 ;
        RECT 161.200 106.800 163.000 107.600 ;
        RECT 164.400 106.800 166.600 107.600 ;
        RECT 167.600 106.800 169.800 107.600 ;
        RECT 170.800 106.800 173.200 107.600 ;
        RECT 174.000 107.200 178.200 107.800 ;
        RECT 179.200 107.600 181.200 108.400 ;
        RECT 186.800 108.200 188.200 109.000 ;
        RECT 188.800 108.400 189.400 112.200 ;
        RECT 193.200 112.400 194.000 119.800 ;
        RECT 195.000 112.400 195.800 112.600 ;
        RECT 193.200 111.800 195.800 112.400 ;
        RECT 197.600 111.800 199.200 119.800 ;
        RECT 201.200 112.400 202.000 112.600 ;
        RECT 202.800 112.400 203.600 119.800 ;
        RECT 205.000 112.400 205.800 119.800 ;
        RECT 201.200 111.800 203.600 112.400 ;
        RECT 204.400 111.800 205.800 112.400 ;
        RECT 190.000 110.300 190.800 111.200 ;
        RECT 196.200 110.400 197.000 110.600 ;
        RECT 198.200 110.400 198.800 111.800 ;
        RECT 190.000 109.700 192.300 110.300 ;
        RECT 190.000 109.600 190.800 109.700 ;
        RECT 191.700 108.400 192.300 109.700 ;
        RECT 195.400 109.800 197.000 110.400 ;
        RECT 195.400 109.600 196.200 109.800 ;
        RECT 198.000 109.600 198.800 110.400 ;
        RECT 196.800 108.600 197.600 108.800 ;
        RECT 194.800 108.400 197.600 108.600 ;
        RECT 186.800 107.800 187.800 108.200 ;
        RECT 155.000 106.200 158.600 106.600 ;
        RECT 135.600 102.200 136.400 106.200 ;
        RECT 137.200 106.000 141.200 106.200 ;
        RECT 137.200 102.200 138.000 106.000 ;
        RECT 140.400 102.200 141.200 106.000 ;
        RECT 142.000 102.200 142.800 106.200 ;
        RECT 143.600 106.000 147.600 106.200 ;
        RECT 143.600 102.200 144.400 106.000 ;
        RECT 146.800 102.200 147.600 106.000 ;
        RECT 153.200 102.200 154.000 106.200 ;
        RECT 154.800 106.000 158.800 106.200 ;
        RECT 154.800 102.200 155.600 106.000 ;
        RECT 158.000 102.200 158.800 106.000 ;
        RECT 161.200 102.200 162.000 106.800 ;
        RECT 164.400 102.200 165.200 106.800 ;
        RECT 167.600 102.200 168.400 106.800 ;
        RECT 170.800 102.200 171.600 106.800 ;
        RECT 174.000 105.000 174.600 107.200 ;
        RECT 179.200 107.000 179.800 107.600 ;
        RECT 179.000 106.600 179.800 107.000 ;
        RECT 178.200 106.000 179.800 106.600 ;
        RECT 183.600 107.200 187.800 107.800 ;
        RECT 188.800 107.600 190.800 108.400 ;
        RECT 191.600 108.300 192.400 108.400 ;
        RECT 193.200 108.300 197.600 108.400 ;
        RECT 191.600 108.000 197.600 108.300 ;
        RECT 198.200 108.400 198.800 109.600 ;
        RECT 204.400 110.400 205.000 111.800 ;
        RECT 209.200 111.200 210.000 119.800 ;
        RECT 210.800 111.800 211.600 119.800 ;
        RECT 212.400 112.400 213.200 119.800 ;
        RECT 215.600 112.400 216.400 119.800 ;
        RECT 218.800 115.600 219.600 119.800 ;
        RECT 222.000 115.800 222.800 119.800 ;
        RECT 222.000 115.600 222.600 115.800 ;
        RECT 219.000 115.000 222.600 115.600 ;
        RECT 220.400 112.800 221.200 114.400 ;
        RECT 222.000 112.400 222.600 115.000 ;
        RECT 212.400 111.800 216.400 112.400 ;
        RECT 206.000 110.800 210.000 111.200 ;
        RECT 205.800 110.600 210.000 110.800 ;
        RECT 204.400 109.600 205.200 110.400 ;
        RECT 205.800 110.000 206.600 110.600 ;
        RECT 211.000 110.400 211.600 111.800 ;
        RECT 217.200 110.800 218.000 112.400 ;
        RECT 222.000 111.600 222.800 112.400 ;
        RECT 214.800 110.400 215.600 110.800 ;
        RECT 191.600 107.800 195.400 108.000 ;
        RECT 198.200 107.800 199.200 108.400 ;
        RECT 191.600 107.700 194.800 107.800 ;
        RECT 191.600 107.600 192.400 107.700 ;
        RECT 193.200 107.600 194.800 107.700 ;
        RECT 174.000 103.000 174.800 105.000 ;
        RECT 178.200 104.400 179.000 106.000 ;
        RECT 183.600 105.000 184.200 107.200 ;
        RECT 188.800 107.000 189.400 107.600 ;
        RECT 188.600 106.600 189.400 107.000 ;
        RECT 195.000 106.800 195.800 107.000 ;
        RECT 187.800 106.400 189.400 106.600 ;
        RECT 186.800 106.000 189.400 106.400 ;
        RECT 193.200 106.200 195.800 106.800 ;
        RECT 196.400 106.400 198.000 107.200 ;
        RECT 186.800 105.600 188.600 106.000 ;
        RECT 178.200 103.600 179.600 104.400 ;
        RECT 178.200 103.000 179.000 103.600 ;
        RECT 183.600 103.000 184.400 105.000 ;
        RECT 187.800 103.000 188.600 105.600 ;
        RECT 193.200 102.200 194.000 106.200 ;
        RECT 198.600 105.800 199.200 107.800 ;
        RECT 200.000 107.600 200.800 108.400 ;
        RECT 202.000 107.600 203.600 108.400 ;
        RECT 200.000 107.200 200.600 107.600 ;
        RECT 199.800 106.400 200.600 107.200 ;
        RECT 201.200 106.800 202.000 107.000 ;
        RECT 201.200 106.200 203.600 106.800 ;
        RECT 197.600 102.200 199.200 105.800 ;
        RECT 202.800 102.200 203.600 106.200 ;
        RECT 204.400 106.200 205.000 109.600 ;
        RECT 205.800 107.000 206.400 110.000 ;
        RECT 210.800 109.800 213.200 110.400 ;
        RECT 214.800 109.800 216.400 110.400 ;
        RECT 210.800 109.600 211.600 109.800 ;
        RECT 207.200 108.400 208.000 109.200 ;
        RECT 207.400 107.600 208.400 108.400 ;
        RECT 210.800 108.300 211.600 108.400 ;
        RECT 209.300 107.700 211.600 108.300 ;
        RECT 205.800 106.400 208.200 107.000 ;
        RECT 209.300 106.400 209.900 107.700 ;
        RECT 210.800 107.600 211.600 107.700 ;
        RECT 204.400 102.200 205.200 106.200 ;
        RECT 207.600 104.200 208.200 106.400 ;
        RECT 209.200 104.800 210.000 106.400 ;
        RECT 210.800 105.600 211.600 106.400 ;
        RECT 212.600 106.200 213.200 109.800 ;
        RECT 215.600 109.600 216.400 109.800 ;
        RECT 218.800 109.600 220.400 110.400 ;
        RECT 214.000 107.600 214.800 109.200 ;
        RECT 222.000 108.400 222.600 111.600 ;
        RECT 221.000 108.200 222.600 108.400 ;
        RECT 220.800 107.800 222.600 108.200 ;
        RECT 211.000 104.800 211.800 105.600 ;
        RECT 207.600 102.200 208.400 104.200 ;
        RECT 212.400 102.200 213.200 106.200 ;
        RECT 220.800 102.200 221.600 107.800 ;
        RECT 223.600 102.200 224.400 119.800 ;
        RECT 226.800 111.200 227.600 119.800 ;
        RECT 231.000 112.400 231.800 119.800 ;
        RECT 235.800 112.600 236.600 119.800 ;
        RECT 231.000 111.800 232.400 112.400 ;
        RECT 234.800 111.800 236.600 112.600 ;
        RECT 238.800 113.600 239.600 114.400 ;
        RECT 238.800 112.400 239.400 113.600 ;
        RECT 240.200 112.400 241.000 119.800 ;
        RECT 246.000 116.400 246.800 119.800 ;
        RECT 245.800 115.800 246.800 116.400 ;
        RECT 245.800 115.200 246.400 115.800 ;
        RECT 249.200 115.200 250.000 119.800 ;
        RECT 252.400 117.000 253.200 119.800 ;
        RECT 254.000 117.000 254.800 119.800 ;
        RECT 238.000 111.800 239.400 112.400 ;
        RECT 240.000 111.800 241.000 112.400 ;
        RECT 244.400 114.600 246.400 115.200 ;
        RECT 226.800 110.800 230.800 111.200 ;
        RECT 226.800 110.600 231.000 110.800 ;
        RECT 230.200 110.000 231.000 110.600 ;
        RECT 231.800 110.400 232.400 111.800 ;
        RECT 228.800 108.400 229.600 109.200 ;
        RECT 225.200 108.300 226.000 108.400 ;
        RECT 228.400 108.300 229.400 108.400 ;
        RECT 225.200 107.700 229.400 108.300 ;
        RECT 225.200 107.600 226.000 107.700 ;
        RECT 228.400 107.600 229.400 107.700 ;
        RECT 230.400 107.000 231.000 110.000 ;
        RECT 231.600 110.300 232.400 110.400 ;
        RECT 233.200 110.300 234.000 110.400 ;
        RECT 231.600 109.700 234.000 110.300 ;
        RECT 231.600 109.600 232.400 109.700 ;
        RECT 233.200 109.600 234.000 109.700 ;
        RECT 228.600 106.400 231.000 107.000 ;
        RECT 225.200 104.800 226.000 106.400 ;
        RECT 226.800 104.800 227.600 106.400 ;
        RECT 228.600 104.200 229.200 106.400 ;
        RECT 231.800 106.200 232.400 109.600 ;
        RECT 235.000 108.400 235.600 111.800 ;
        RECT 238.000 111.600 238.800 111.800 ;
        RECT 236.400 109.600 237.200 111.200 ;
        RECT 240.000 108.400 240.600 111.800 ;
        RECT 241.200 108.800 242.000 110.400 ;
        RECT 244.400 109.000 245.200 114.600 ;
        RECT 247.000 114.400 251.200 115.200 ;
        RECT 255.600 115.000 256.400 119.800 ;
        RECT 258.800 115.000 259.600 119.800 ;
        RECT 247.000 114.000 247.600 114.400 ;
        RECT 246.000 113.200 247.600 114.000 ;
        RECT 250.600 113.800 256.400 114.400 ;
        RECT 248.600 113.200 250.000 113.800 ;
        RECT 248.600 113.000 254.800 113.200 ;
        RECT 249.400 112.600 254.800 113.000 ;
        RECT 254.000 112.400 254.800 112.600 ;
        RECT 255.800 113.000 256.400 113.800 ;
        RECT 257.000 113.600 259.600 114.400 ;
        RECT 262.000 113.600 262.800 119.800 ;
        RECT 263.600 117.000 264.400 119.800 ;
        RECT 265.200 117.000 266.000 119.800 ;
        RECT 266.800 117.000 267.600 119.800 ;
        RECT 265.200 114.400 269.400 115.200 ;
        RECT 270.000 114.400 270.800 119.800 ;
        RECT 273.200 115.200 274.000 119.800 ;
        RECT 273.200 114.600 275.800 115.200 ;
        RECT 270.000 113.600 272.600 114.400 ;
        RECT 263.600 113.000 264.400 113.200 ;
        RECT 255.800 112.400 264.400 113.000 ;
        RECT 266.800 113.000 267.600 113.200 ;
        RECT 275.200 113.000 275.800 114.600 ;
        RECT 266.800 112.400 275.800 113.000 ;
        RECT 247.600 111.800 248.400 112.400 ;
        RECT 250.800 111.800 251.800 112.000 ;
        RECT 247.600 111.200 274.600 111.800 ;
        RECT 273.800 111.000 274.600 111.200 ;
        RECT 275.200 110.600 275.800 112.400 ;
        RECT 276.400 112.000 277.200 119.800 ;
        RECT 280.400 113.600 281.200 114.400 ;
        RECT 280.400 112.400 281.000 113.600 ;
        RECT 281.800 112.400 282.600 119.800 ;
        RECT 287.600 112.800 288.400 119.800 ;
        RECT 276.400 111.200 277.400 112.000 ;
        RECT 279.600 111.800 281.000 112.400 ;
        RECT 281.600 111.800 282.600 112.400 ;
        RECT 287.400 111.800 288.400 112.800 ;
        RECT 290.800 112.400 291.600 119.800 ;
        RECT 289.000 111.800 291.600 112.400 ;
        RECT 292.400 112.400 293.200 119.800 ;
        RECT 294.200 112.400 295.000 112.600 ;
        RECT 292.400 111.800 295.000 112.400 ;
        RECT 296.800 111.800 298.400 119.800 ;
        RECT 300.400 112.400 301.200 112.600 ;
        RECT 302.000 112.400 302.800 119.800 ;
        RECT 300.400 111.800 302.800 112.400 ;
        RECT 279.600 111.600 280.400 111.800 ;
        RECT 275.200 110.000 276.000 110.600 ;
        RECT 234.800 107.600 235.600 108.400 ;
        RECT 238.000 107.600 240.600 108.400 ;
        RECT 242.800 108.200 243.600 108.400 ;
        RECT 242.000 107.600 243.600 108.200 ;
        RECT 244.400 108.200 253.200 109.000 ;
        RECT 253.800 108.600 255.800 109.400 ;
        RECT 259.600 108.600 262.800 109.400 ;
        RECT 228.400 102.200 229.200 104.200 ;
        RECT 231.600 102.200 232.400 106.200 ;
        RECT 233.200 104.800 234.000 106.400 ;
        RECT 235.000 106.300 235.600 107.600 ;
        RECT 236.400 106.300 237.200 106.400 ;
        RECT 234.900 105.700 237.200 106.300 ;
        RECT 238.200 106.200 238.800 107.600 ;
        RECT 242.000 107.200 242.800 107.600 ;
        RECT 239.800 106.200 243.400 106.600 ;
        RECT 235.000 104.200 235.600 105.700 ;
        RECT 236.400 105.600 237.200 105.700 ;
        RECT 234.800 102.200 235.600 104.200 ;
        RECT 238.000 102.200 238.800 106.200 ;
        RECT 239.600 106.000 243.600 106.200 ;
        RECT 239.600 102.200 240.400 106.000 ;
        RECT 242.800 102.200 243.600 106.000 ;
        RECT 244.400 102.200 245.200 108.200 ;
        RECT 246.800 106.800 249.800 107.600 ;
        RECT 249.000 106.200 249.800 106.800 ;
        RECT 255.000 106.200 255.800 108.600 ;
        RECT 257.200 106.800 258.000 108.400 ;
        RECT 262.400 107.800 263.200 108.000 ;
        RECT 258.800 107.200 263.200 107.800 ;
        RECT 258.800 107.000 259.600 107.200 ;
        RECT 265.200 106.400 266.000 109.200 ;
        RECT 271.000 108.600 274.800 109.400 ;
        RECT 271.000 107.400 271.800 108.600 ;
        RECT 275.400 108.000 276.000 110.000 ;
        RECT 258.800 106.200 259.600 106.400 ;
        RECT 249.000 105.400 251.600 106.200 ;
        RECT 255.000 105.600 259.600 106.200 ;
        RECT 260.400 105.600 262.000 106.400 ;
        RECT 265.000 105.600 266.000 106.400 ;
        RECT 270.000 106.800 271.800 107.400 ;
        RECT 274.800 107.400 276.000 108.000 ;
        RECT 270.000 106.200 270.800 106.800 ;
        RECT 250.800 102.200 251.600 105.400 ;
        RECT 268.400 105.400 270.800 106.200 ;
        RECT 252.400 102.200 253.200 105.000 ;
        RECT 254.000 102.200 254.800 105.000 ;
        RECT 255.600 102.200 256.400 105.000 ;
        RECT 258.800 102.200 259.600 105.000 ;
        RECT 262.000 102.200 262.800 105.000 ;
        RECT 263.600 102.200 264.400 105.000 ;
        RECT 265.200 102.200 266.000 105.000 ;
        RECT 266.800 102.200 267.600 105.000 ;
        RECT 268.400 102.200 269.200 105.400 ;
        RECT 274.800 102.200 275.600 107.400 ;
        RECT 276.600 106.800 277.400 111.200 ;
        RECT 281.600 108.400 282.200 111.800 ;
        RECT 282.800 108.800 283.600 110.400 ;
        RECT 287.400 108.400 288.000 111.800 ;
        RECT 289.000 109.800 289.600 111.800 ;
        RECT 295.400 110.400 296.200 110.600 ;
        RECT 297.400 110.400 298.000 111.800 ;
        RECT 288.600 109.000 289.600 109.800 ;
        RECT 279.600 107.600 282.200 108.400 ;
        RECT 284.400 108.300 285.200 108.400 ;
        RECT 287.400 108.300 288.400 108.400 ;
        RECT 284.400 108.200 288.400 108.300 ;
        RECT 283.600 107.700 288.400 108.200 ;
        RECT 283.600 107.600 285.200 107.700 ;
        RECT 287.400 107.600 288.400 107.700 ;
        RECT 276.400 106.000 277.400 106.800 ;
        RECT 279.800 106.200 280.400 107.600 ;
        RECT 283.600 107.200 284.400 107.600 ;
        RECT 281.400 106.200 285.000 106.600 ;
        RECT 287.400 106.200 288.000 107.600 ;
        RECT 289.000 107.400 289.600 109.000 ;
        RECT 290.600 109.600 291.600 110.400 ;
        RECT 294.600 109.800 296.200 110.400 ;
        RECT 294.600 109.600 295.400 109.800 ;
        RECT 297.200 109.600 298.000 110.400 ;
        RECT 290.600 108.800 291.400 109.600 ;
        RECT 296.000 108.600 296.800 108.800 ;
        RECT 294.000 108.400 296.800 108.600 ;
        RECT 292.400 108.000 296.800 108.400 ;
        RECT 297.400 108.400 298.000 109.600 ;
        RECT 292.400 107.800 294.600 108.000 ;
        RECT 297.400 107.800 298.400 108.400 ;
        RECT 292.400 107.600 294.000 107.800 ;
        RECT 289.000 106.800 291.600 107.400 ;
        RECT 294.200 106.800 295.000 107.000 ;
        RECT 276.400 102.200 277.200 106.000 ;
        RECT 279.600 102.200 280.400 106.200 ;
        RECT 281.200 106.000 285.200 106.200 ;
        RECT 281.200 102.200 282.000 106.000 ;
        RECT 284.400 102.200 285.200 106.000 ;
        RECT 287.400 105.600 288.400 106.200 ;
        RECT 287.600 102.200 288.400 105.600 ;
        RECT 290.800 102.200 291.600 106.800 ;
        RECT 292.400 106.200 295.000 106.800 ;
        RECT 295.600 106.400 297.200 107.200 ;
        RECT 292.400 102.200 293.200 106.200 ;
        RECT 297.800 105.800 298.400 107.800 ;
        RECT 299.200 107.600 300.000 108.400 ;
        RECT 301.200 107.600 302.800 108.400 ;
        RECT 299.200 107.200 299.800 107.600 ;
        RECT 299.000 106.400 299.800 107.200 ;
        RECT 300.400 106.800 301.200 107.000 ;
        RECT 308.400 106.800 309.200 108.400 ;
        RECT 300.400 106.200 302.800 106.800 ;
        RECT 296.800 102.200 298.400 105.800 ;
        RECT 302.000 102.200 302.800 106.200 ;
        RECT 310.000 106.200 310.800 119.800 ;
        RECT 311.600 112.300 312.400 113.200 ;
        RECT 314.800 112.300 315.600 119.800 ;
        RECT 318.000 115.200 318.800 119.800 ;
        RECT 311.600 111.700 315.600 112.300 ;
        RECT 311.600 111.600 312.400 111.700 ;
        RECT 314.600 111.200 315.600 111.700 ;
        RECT 316.200 114.600 318.800 115.200 ;
        RECT 316.200 113.000 316.800 114.600 ;
        RECT 321.200 114.400 322.000 119.800 ;
        RECT 324.400 117.000 325.200 119.800 ;
        RECT 326.000 117.000 326.800 119.800 ;
        RECT 327.600 117.000 328.400 119.800 ;
        RECT 322.600 114.400 326.800 115.200 ;
        RECT 319.400 113.600 322.000 114.400 ;
        RECT 329.200 113.600 330.000 119.800 ;
        RECT 332.400 115.000 333.200 119.800 ;
        RECT 335.600 115.000 336.400 119.800 ;
        RECT 337.200 117.000 338.000 119.800 ;
        RECT 338.800 117.000 339.600 119.800 ;
        RECT 342.000 115.200 342.800 119.800 ;
        RECT 345.200 116.400 346.000 119.800 ;
        RECT 345.200 115.800 346.200 116.400 ;
        RECT 345.600 115.200 346.200 115.800 ;
        RECT 340.800 114.400 345.000 115.200 ;
        RECT 345.600 114.600 347.600 115.200 ;
        RECT 332.400 113.600 335.000 114.400 ;
        RECT 335.600 113.800 341.400 114.400 ;
        RECT 344.400 114.000 345.000 114.400 ;
        RECT 324.400 113.000 325.200 113.200 ;
        RECT 316.200 112.400 325.200 113.000 ;
        RECT 327.600 113.000 328.400 113.200 ;
        RECT 335.600 113.000 336.200 113.800 ;
        RECT 342.000 113.200 343.400 113.800 ;
        RECT 344.400 113.200 346.000 114.000 ;
        RECT 327.600 112.400 336.200 113.000 ;
        RECT 337.200 113.000 343.400 113.200 ;
        RECT 337.200 112.600 342.600 113.000 ;
        RECT 337.200 112.400 338.000 112.600 ;
        RECT 314.600 106.800 315.400 111.200 ;
        RECT 316.200 110.600 316.800 112.400 ;
        RECT 316.000 110.000 316.800 110.600 ;
        RECT 322.800 110.000 346.200 110.600 ;
        RECT 316.000 108.000 316.600 110.000 ;
        RECT 322.800 109.400 323.600 110.000 ;
        RECT 340.400 109.600 341.200 110.000 ;
        RECT 343.600 109.600 344.400 110.000 ;
        RECT 345.400 109.800 346.200 110.000 ;
        RECT 317.200 108.600 321.000 109.400 ;
        RECT 316.000 107.400 317.200 108.000 ;
        RECT 310.000 105.600 311.800 106.200 ;
        RECT 314.600 106.000 315.600 106.800 ;
        RECT 311.000 104.400 311.800 105.600 ;
        RECT 310.000 103.600 311.800 104.400 ;
        RECT 311.000 102.200 311.800 103.600 ;
        RECT 314.800 102.200 315.600 106.000 ;
        RECT 316.400 102.200 317.200 107.400 ;
        RECT 320.200 107.400 321.000 108.600 ;
        RECT 320.200 106.800 322.000 107.400 ;
        RECT 321.200 106.200 322.000 106.800 ;
        RECT 326.000 106.400 326.800 109.200 ;
        RECT 329.200 108.600 332.400 109.400 ;
        RECT 336.200 108.600 338.200 109.400 ;
        RECT 346.800 109.000 347.600 114.600 ;
        RECT 350.000 112.800 350.800 119.800 ;
        RECT 328.800 107.800 329.600 108.000 ;
        RECT 328.800 107.200 333.200 107.800 ;
        RECT 332.400 107.000 333.200 107.200 ;
        RECT 334.000 106.800 334.800 108.400 ;
        RECT 321.200 105.400 323.600 106.200 ;
        RECT 326.000 105.600 327.000 106.400 ;
        RECT 330.000 105.600 331.600 106.400 ;
        RECT 332.400 106.200 333.200 106.400 ;
        RECT 336.200 106.200 337.000 108.600 ;
        RECT 338.800 108.200 347.600 109.000 ;
        RECT 342.200 106.800 345.200 107.600 ;
        RECT 342.200 106.200 343.000 106.800 ;
        RECT 332.400 105.600 337.000 106.200 ;
        RECT 322.800 102.200 323.600 105.400 ;
        RECT 340.400 105.400 343.000 106.200 ;
        RECT 324.400 102.200 325.200 105.000 ;
        RECT 326.000 102.200 326.800 105.000 ;
        RECT 327.600 102.200 328.400 105.000 ;
        RECT 329.200 102.200 330.000 105.000 ;
        RECT 332.400 102.200 333.200 105.000 ;
        RECT 335.600 102.200 336.400 105.000 ;
        RECT 337.200 102.200 338.000 105.000 ;
        RECT 338.800 102.200 339.600 105.000 ;
        RECT 340.400 102.200 341.200 105.400 ;
        RECT 346.800 102.200 347.600 108.200 ;
        RECT 349.800 111.800 350.800 112.800 ;
        RECT 353.200 112.400 354.000 119.800 ;
        RECT 351.400 111.800 354.000 112.400 ;
        RECT 354.800 112.400 355.600 119.800 ;
        RECT 358.000 112.800 358.800 119.800 ;
        RECT 354.800 111.800 357.400 112.400 ;
        RECT 358.000 111.800 359.000 112.800 ;
        RECT 349.800 108.400 350.400 111.800 ;
        RECT 351.400 109.800 352.000 111.800 ;
        RECT 351.000 109.000 352.000 109.800 ;
        RECT 349.800 107.600 350.800 108.400 ;
        RECT 349.800 106.200 350.400 107.600 ;
        RECT 351.400 107.400 352.000 109.000 ;
        RECT 353.000 110.300 354.000 110.400 ;
        RECT 354.800 110.300 355.800 110.400 ;
        RECT 353.000 109.700 355.800 110.300 ;
        RECT 353.000 109.600 354.000 109.700 ;
        RECT 354.800 109.600 355.800 109.700 ;
        RECT 353.000 108.800 353.800 109.600 ;
        RECT 355.000 108.800 355.800 109.600 ;
        RECT 356.800 109.800 357.400 111.800 ;
        RECT 356.800 109.000 357.800 109.800 ;
        RECT 356.800 107.400 357.400 109.000 ;
        RECT 358.400 108.400 359.000 111.800 ;
        RECT 358.000 107.600 359.000 108.400 ;
        RECT 351.400 106.800 354.000 107.400 ;
        RECT 349.800 105.600 350.800 106.200 ;
        RECT 350.000 102.200 350.800 105.600 ;
        RECT 353.200 102.200 354.000 106.800 ;
        RECT 354.800 106.800 357.400 107.400 ;
        RECT 354.800 102.200 355.600 106.800 ;
        RECT 358.400 106.200 359.000 107.600 ;
        RECT 358.000 105.600 359.000 106.200 ;
        RECT 361.200 110.300 362.000 119.800 ;
        RECT 367.000 112.400 367.800 119.800 ;
        RECT 372.400 116.400 373.200 119.800 ;
        RECT 372.200 115.800 373.200 116.400 ;
        RECT 372.200 115.200 372.800 115.800 ;
        RECT 375.600 115.200 376.400 119.800 ;
        RECT 378.800 117.000 379.600 119.800 ;
        RECT 380.400 117.000 381.200 119.800 ;
        RECT 370.800 114.600 372.800 115.200 ;
        RECT 368.400 113.600 369.200 114.400 ;
        RECT 368.600 112.400 369.200 113.600 ;
        RECT 367.000 111.800 368.000 112.400 ;
        RECT 368.600 111.800 370.000 112.400 ;
        RECT 366.000 110.300 366.800 110.400 ;
        RECT 361.200 109.700 366.800 110.300 ;
        RECT 358.000 102.200 358.800 105.600 ;
        RECT 361.200 102.200 362.000 109.700 ;
        RECT 366.000 108.800 366.800 109.700 ;
        RECT 367.400 108.400 368.000 111.800 ;
        RECT 369.200 111.600 370.000 111.800 ;
        RECT 370.800 109.000 371.600 114.600 ;
        RECT 373.400 114.400 377.600 115.200 ;
        RECT 382.000 115.000 382.800 119.800 ;
        RECT 385.200 115.000 386.000 119.800 ;
        RECT 373.400 114.000 374.000 114.400 ;
        RECT 372.400 113.200 374.000 114.000 ;
        RECT 377.000 113.800 382.800 114.400 ;
        RECT 375.000 113.200 376.400 113.800 ;
        RECT 375.000 113.000 381.200 113.200 ;
        RECT 375.800 112.600 381.200 113.000 ;
        RECT 380.400 112.400 381.200 112.600 ;
        RECT 382.200 113.000 382.800 113.800 ;
        RECT 383.400 113.600 386.000 114.400 ;
        RECT 388.400 113.600 389.200 119.800 ;
        RECT 390.000 117.000 390.800 119.800 ;
        RECT 391.600 117.000 392.400 119.800 ;
        RECT 393.200 117.000 394.000 119.800 ;
        RECT 391.600 114.400 395.800 115.200 ;
        RECT 396.400 114.400 397.200 119.800 ;
        RECT 399.600 115.200 400.400 119.800 ;
        RECT 399.600 114.600 402.200 115.200 ;
        RECT 396.400 113.600 399.000 114.400 ;
        RECT 390.000 113.000 390.800 113.200 ;
        RECT 382.200 112.400 390.800 113.000 ;
        RECT 393.200 113.000 394.000 113.200 ;
        RECT 401.600 113.000 402.200 114.600 ;
        RECT 393.200 112.400 402.200 113.000 ;
        RECT 401.600 110.600 402.200 112.400 ;
        RECT 402.800 112.000 403.600 119.800 ;
        RECT 402.800 111.200 403.800 112.000 ;
        RECT 372.200 110.000 395.600 110.600 ;
        RECT 401.600 110.000 402.400 110.600 ;
        RECT 372.200 109.800 373.000 110.000 ;
        RECT 377.200 109.600 378.000 110.000 ;
        RECT 394.800 109.400 395.600 110.000 ;
        RECT 364.400 108.200 365.200 108.400 ;
        RECT 364.400 107.600 366.000 108.200 ;
        RECT 367.400 107.600 370.000 108.400 ;
        RECT 370.800 108.200 379.600 109.000 ;
        RECT 380.200 108.600 382.200 109.400 ;
        RECT 386.000 108.600 389.200 109.400 ;
        RECT 365.200 107.200 366.000 107.600 ;
        RECT 362.800 104.800 363.600 106.400 ;
        RECT 364.600 106.200 368.200 106.600 ;
        RECT 369.200 106.200 369.800 107.600 ;
        RECT 364.400 106.000 368.400 106.200 ;
        RECT 364.400 102.200 365.200 106.000 ;
        RECT 367.600 102.200 368.400 106.000 ;
        RECT 369.200 102.200 370.000 106.200 ;
        RECT 370.800 102.200 371.600 108.200 ;
        RECT 373.200 106.800 376.200 107.600 ;
        RECT 375.400 106.200 376.200 106.800 ;
        RECT 381.400 106.200 382.200 108.600 ;
        RECT 383.600 106.800 384.400 108.400 ;
        RECT 388.800 107.800 389.600 108.000 ;
        RECT 385.200 107.200 389.600 107.800 ;
        RECT 385.200 107.000 386.000 107.200 ;
        RECT 391.600 106.400 392.400 109.200 ;
        RECT 397.400 108.600 401.200 109.400 ;
        RECT 397.400 107.400 398.200 108.600 ;
        RECT 401.800 108.000 402.400 110.000 ;
        RECT 385.200 106.200 386.000 106.400 ;
        RECT 375.400 105.400 378.000 106.200 ;
        RECT 381.400 105.600 386.000 106.200 ;
        RECT 386.800 105.600 388.400 106.400 ;
        RECT 391.400 105.600 392.400 106.400 ;
        RECT 396.400 106.800 398.200 107.400 ;
        RECT 401.200 107.400 402.400 108.000 ;
        RECT 396.400 106.200 397.200 106.800 ;
        RECT 377.200 102.200 378.000 105.400 ;
        RECT 394.800 105.400 397.200 106.200 ;
        RECT 378.800 102.200 379.600 105.000 ;
        RECT 380.400 102.200 381.200 105.000 ;
        RECT 382.000 102.200 382.800 105.000 ;
        RECT 385.200 102.200 386.000 105.000 ;
        RECT 388.400 102.200 389.200 105.000 ;
        RECT 390.000 102.200 390.800 105.000 ;
        RECT 391.600 102.200 392.400 105.000 ;
        RECT 393.200 102.200 394.000 105.000 ;
        RECT 394.800 102.200 395.600 105.400 ;
        RECT 401.200 102.200 402.000 107.400 ;
        RECT 403.000 106.800 403.800 111.200 ;
        RECT 402.800 106.000 403.800 106.800 ;
        RECT 406.000 111.200 406.800 119.800 ;
        RECT 410.200 115.800 411.400 119.800 ;
        RECT 414.800 115.800 415.600 119.800 ;
        RECT 419.200 116.400 420.000 119.800 ;
        RECT 419.200 115.800 421.200 116.400 ;
        RECT 410.800 115.000 411.600 115.800 ;
        RECT 415.000 115.200 415.600 115.800 ;
        RECT 414.200 114.600 417.800 115.200 ;
        RECT 420.400 115.000 421.200 115.800 ;
        RECT 414.200 114.400 415.000 114.600 ;
        RECT 417.000 114.400 417.800 114.600 ;
        RECT 410.000 113.200 411.400 114.000 ;
        RECT 410.800 112.200 411.400 113.200 ;
        RECT 413.000 113.000 415.200 113.600 ;
        RECT 413.000 112.800 413.800 113.000 ;
        RECT 410.800 111.600 413.200 112.200 ;
        RECT 406.000 110.600 410.200 111.200 ;
        RECT 406.000 107.200 406.800 110.600 ;
        RECT 409.400 110.400 410.200 110.600 ;
        RECT 407.800 109.800 408.600 110.000 ;
        RECT 407.800 109.200 411.600 109.800 ;
        RECT 410.800 109.000 411.600 109.200 ;
        RECT 412.600 108.400 413.200 111.600 ;
        RECT 414.600 111.800 415.200 113.000 ;
        RECT 415.800 113.000 416.600 113.200 ;
        RECT 420.400 113.000 421.200 113.200 ;
        RECT 415.800 112.400 421.200 113.000 ;
        RECT 414.600 111.400 419.400 111.800 ;
        RECT 423.600 111.400 424.400 119.800 ;
        RECT 414.600 111.200 424.400 111.400 ;
        RECT 418.600 111.000 424.400 111.200 ;
        RECT 418.800 110.800 424.400 111.000 ;
        RECT 417.200 110.200 418.000 110.400 ;
        RECT 417.200 109.600 422.200 110.200 ;
        RECT 418.800 109.400 419.600 109.600 ;
        RECT 421.400 109.400 422.200 109.600 ;
        RECT 419.800 108.400 420.600 108.600 ;
        RECT 407.600 107.200 408.400 108.400 ;
        RECT 412.600 107.800 423.600 108.400 ;
        RECT 413.000 107.600 413.800 107.800 ;
        RECT 415.600 107.600 416.400 107.800 ;
        RECT 406.000 106.600 409.800 107.200 ;
        RECT 402.800 102.200 403.600 106.000 ;
        RECT 406.000 102.200 406.800 106.600 ;
        RECT 409.000 106.400 409.800 106.600 ;
        RECT 418.800 105.600 419.400 107.800 ;
        RECT 422.000 107.600 423.600 107.800 ;
        RECT 417.000 105.400 417.800 105.600 ;
        RECT 410.800 104.200 411.600 105.000 ;
        RECT 415.000 104.800 417.800 105.400 ;
        RECT 418.800 104.800 419.600 105.600 ;
        RECT 415.000 104.200 415.600 104.800 ;
        RECT 420.400 104.200 421.200 105.000 ;
        RECT 410.200 103.600 411.600 104.200 ;
        RECT 410.200 102.200 411.400 103.600 ;
        RECT 414.800 102.200 415.600 104.200 ;
        RECT 419.200 103.600 421.200 104.200 ;
        RECT 419.200 102.200 420.000 103.600 ;
        RECT 423.600 102.200 424.400 107.000 ;
        RECT 425.200 104.800 426.000 106.400 ;
        RECT 426.800 102.200 427.600 119.800 ;
        RECT 429.200 113.600 430.000 114.400 ;
        RECT 429.200 112.400 429.800 113.600 ;
        RECT 430.600 112.400 431.400 119.800 ;
        RECT 438.600 112.800 439.400 119.800 ;
        RECT 442.800 115.000 443.600 119.000 ;
        RECT 428.400 111.800 429.800 112.400 ;
        RECT 430.400 111.800 431.400 112.400 ;
        RECT 437.800 112.200 439.400 112.800 ;
        RECT 428.400 111.600 429.200 111.800 ;
        RECT 430.400 108.400 431.000 111.800 ;
        RECT 431.600 110.300 432.400 110.400 ;
        RECT 431.600 109.700 435.500 110.300 ;
        RECT 431.600 108.800 432.400 109.700 ;
        RECT 428.400 107.600 431.000 108.400 ;
        RECT 433.200 108.200 434.000 108.400 ;
        RECT 432.400 107.600 434.000 108.200 ;
        RECT 434.900 108.300 435.500 109.700 ;
        RECT 436.400 109.600 437.200 111.200 ;
        RECT 437.800 108.400 438.400 112.200 ;
        RECT 443.000 111.600 443.600 115.000 ;
        RECT 445.200 113.600 446.000 114.400 ;
        RECT 445.200 112.400 445.800 113.600 ;
        RECT 446.600 112.400 447.400 119.800 ;
        RECT 451.600 113.600 452.400 114.400 ;
        RECT 451.600 112.400 452.200 113.600 ;
        RECT 453.000 112.400 453.800 119.800 ;
        RECT 444.400 111.800 445.800 112.400 ;
        RECT 446.400 111.800 447.400 112.400 ;
        RECT 450.800 111.800 452.200 112.400 ;
        RECT 452.800 111.800 453.800 112.400 ;
        RECT 444.400 111.600 445.200 111.800 ;
        RECT 439.800 111.000 443.600 111.600 ;
        RECT 439.800 109.000 440.400 111.000 ;
        RECT 436.400 108.300 438.400 108.400 ;
        RECT 434.900 107.700 438.400 108.300 ;
        RECT 439.000 108.200 440.400 109.000 ;
        RECT 441.200 108.800 442.000 110.400 ;
        RECT 442.800 110.300 443.600 110.400 ;
        RECT 444.400 110.300 445.200 110.400 ;
        RECT 442.800 109.700 445.200 110.300 ;
        RECT 442.800 108.800 443.600 109.700 ;
        RECT 444.400 109.600 445.200 109.700 ;
        RECT 446.400 108.400 447.000 111.800 ;
        RECT 450.800 111.600 451.600 111.800 ;
        RECT 447.600 110.300 448.400 110.400 ;
        RECT 450.800 110.300 451.600 110.400 ;
        RECT 447.600 109.700 451.600 110.300 ;
        RECT 447.600 108.800 448.400 109.700 ;
        RECT 450.800 109.600 451.600 109.700 ;
        RECT 452.800 108.400 453.400 111.800 ;
        RECT 454.000 108.800 454.800 110.400 ;
        RECT 436.400 107.600 438.400 107.700 ;
        RECT 428.600 106.200 429.200 107.600 ;
        RECT 432.400 107.200 433.200 107.600 ;
        RECT 437.800 107.000 438.400 107.600 ;
        RECT 439.400 107.800 440.400 108.200 ;
        RECT 439.400 107.200 443.600 107.800 ;
        RECT 444.400 107.600 447.000 108.400 ;
        RECT 449.200 108.300 450.000 108.400 ;
        RECT 450.800 108.300 453.400 108.400 ;
        RECT 449.200 108.200 453.400 108.300 ;
        RECT 455.600 108.200 456.400 108.400 ;
        RECT 448.400 107.700 453.400 108.200 ;
        RECT 448.400 107.600 450.000 107.700 ;
        RECT 450.800 107.600 453.400 107.700 ;
        RECT 454.800 107.600 456.400 108.200 ;
        RECT 437.800 106.600 438.600 107.000 ;
        RECT 430.200 106.200 433.800 106.600 ;
        RECT 428.400 102.200 429.200 106.200 ;
        RECT 430.000 106.000 434.000 106.200 ;
        RECT 437.800 106.000 439.400 106.600 ;
        RECT 430.000 102.200 430.800 106.000 ;
        RECT 433.200 102.200 434.000 106.000 ;
        RECT 438.600 103.000 439.400 106.000 ;
        RECT 443.000 105.000 443.600 107.200 ;
        RECT 444.600 106.400 445.200 107.600 ;
        RECT 448.400 107.200 449.200 107.600 ;
        RECT 442.800 103.000 443.600 105.000 ;
        RECT 444.400 102.200 445.200 106.400 ;
        RECT 446.200 106.200 449.800 106.600 ;
        RECT 451.000 106.200 451.600 107.600 ;
        RECT 454.800 107.200 455.600 107.600 ;
        RECT 462.000 106.800 462.800 108.400 ;
        RECT 452.600 106.200 456.200 106.600 ;
        RECT 463.600 106.200 464.400 119.800 ;
        RECT 465.200 112.300 466.000 113.200 ;
        RECT 466.800 112.300 467.600 119.800 ;
        RECT 465.200 111.700 467.600 112.300 ;
        RECT 465.200 111.600 466.000 111.700 ;
        RECT 446.000 106.000 450.000 106.200 ;
        RECT 446.000 102.200 446.800 106.000 ;
        RECT 449.200 102.200 450.000 106.000 ;
        RECT 450.800 102.200 451.600 106.200 ;
        RECT 452.400 106.000 456.400 106.200 ;
        RECT 452.400 102.200 453.200 106.000 ;
        RECT 455.600 102.200 456.400 106.000 ;
        RECT 463.600 105.600 465.400 106.200 ;
        RECT 464.600 104.400 465.400 105.600 ;
        RECT 463.600 103.600 465.400 104.400 ;
        RECT 464.600 102.200 465.400 103.600 ;
        RECT 466.800 102.200 467.600 111.700 ;
        RECT 468.400 110.300 469.200 110.400 ;
        RECT 470.000 110.300 470.800 119.800 ;
        RECT 471.600 114.300 472.400 114.400 ;
        RECT 474.800 114.300 475.600 119.800 ;
        RECT 471.600 113.700 475.600 114.300 ;
        RECT 471.600 113.600 472.400 113.700 ;
        RECT 468.400 109.700 470.800 110.300 ;
        RECT 468.400 109.600 469.200 109.700 ;
        RECT 468.400 104.800 469.200 106.400 ;
        RECT 470.000 102.200 470.800 109.700 ;
        RECT 471.600 108.300 472.400 108.400 ;
        RECT 473.200 108.300 474.000 108.400 ;
        RECT 471.600 107.700 474.000 108.300 ;
        RECT 471.600 107.600 472.400 107.700 ;
        RECT 473.200 106.800 474.000 107.700 ;
        RECT 471.600 104.800 472.400 106.400 ;
        RECT 474.800 106.200 475.600 113.700 ;
        RECT 480.600 118.400 481.400 119.800 ;
        RECT 480.600 117.600 482.000 118.400 ;
        RECT 476.400 111.600 477.200 113.200 ;
        RECT 480.600 112.600 481.400 117.600 ;
        RECT 479.600 111.800 481.400 112.600 ;
        RECT 483.600 113.600 484.400 114.400 ;
        RECT 483.600 112.400 484.200 113.600 ;
        RECT 485.000 112.400 485.800 119.800 ;
        RECT 482.800 111.800 484.200 112.400 ;
        RECT 484.800 111.800 485.800 112.400 ;
        RECT 479.800 108.400 480.400 111.800 ;
        RECT 482.800 111.600 483.600 111.800 ;
        RECT 481.200 109.600 482.000 111.200 ;
        RECT 484.800 108.400 485.400 111.800 ;
        RECT 489.200 111.600 490.000 113.200 ;
        RECT 486.000 108.800 486.800 110.400 ;
        RECT 489.200 110.300 490.000 110.400 ;
        RECT 490.800 110.300 491.600 119.800 ;
        RECT 496.600 112.400 497.400 119.800 ;
        RECT 498.000 113.600 498.800 114.400 ;
        RECT 498.200 112.400 498.800 113.600 ;
        RECT 496.600 111.800 497.600 112.400 ;
        RECT 498.200 112.300 499.600 112.400 ;
        RECT 502.000 112.300 502.800 119.800 ;
        RECT 498.200 111.800 502.800 112.300 ;
        RECT 489.200 109.700 491.600 110.300 ;
        RECT 489.200 109.600 490.000 109.700 ;
        RECT 479.600 107.600 480.400 108.400 ;
        RECT 482.800 107.600 485.400 108.400 ;
        RECT 487.600 108.200 488.400 108.400 ;
        RECT 486.800 107.600 488.400 108.200 ;
        RECT 474.800 105.600 476.600 106.200 ;
        RECT 475.800 104.400 476.600 105.600 ;
        RECT 478.000 104.800 478.800 106.400 ;
        RECT 474.800 103.600 476.600 104.400 ;
        RECT 479.800 104.200 480.400 107.600 ;
        RECT 483.000 106.200 483.600 107.600 ;
        RECT 486.800 107.200 487.600 107.600 ;
        RECT 484.600 106.200 488.200 106.600 ;
        RECT 490.800 106.200 491.600 109.700 ;
        RECT 492.400 110.300 493.200 110.400 ;
        RECT 495.600 110.300 496.400 110.400 ;
        RECT 492.400 109.700 496.400 110.300 ;
        RECT 492.400 109.600 493.200 109.700 ;
        RECT 495.600 108.800 496.400 109.700 ;
        RECT 497.000 108.400 497.600 111.800 ;
        RECT 498.800 111.700 502.800 111.800 ;
        RECT 498.800 111.600 499.600 111.700 ;
        RECT 492.400 106.800 493.200 108.400 ;
        RECT 494.000 108.200 494.800 108.400 ;
        RECT 494.000 107.600 495.600 108.200 ;
        RECT 497.000 107.600 499.600 108.400 ;
        RECT 494.800 107.200 495.600 107.600 ;
        RECT 494.200 106.200 497.800 106.600 ;
        RECT 498.800 106.200 499.400 107.600 ;
        RECT 500.400 106.800 501.200 108.400 ;
        RECT 502.000 106.200 502.800 111.700 ;
        RECT 503.600 111.600 504.400 114.400 ;
        RECT 475.800 102.200 476.600 103.600 ;
        RECT 479.600 102.200 480.400 104.200 ;
        RECT 482.800 102.200 483.600 106.200 ;
        RECT 484.400 106.000 488.400 106.200 ;
        RECT 484.400 102.200 485.200 106.000 ;
        RECT 487.600 102.200 488.400 106.000 ;
        RECT 489.800 105.600 491.600 106.200 ;
        RECT 494.000 106.000 498.000 106.200 ;
        RECT 489.800 102.200 490.600 105.600 ;
        RECT 494.000 102.200 494.800 106.000 ;
        RECT 497.200 102.200 498.000 106.000 ;
        RECT 498.800 102.200 499.600 106.200 ;
        RECT 502.000 105.600 503.800 106.200 ;
        RECT 503.000 102.200 503.800 105.600 ;
        RECT 505.200 102.200 506.000 119.800 ;
        RECT 511.000 112.400 511.800 119.800 ;
        RECT 512.400 113.600 513.200 114.400 ;
        RECT 512.600 112.400 513.200 113.600 ;
        RECT 518.600 112.800 519.400 119.800 ;
        RECT 522.800 115.000 523.600 119.000 ;
        RECT 510.000 111.600 512.000 112.400 ;
        RECT 512.600 111.800 514.000 112.400 ;
        RECT 513.200 111.600 514.000 111.800 ;
        RECT 517.800 112.200 519.400 112.800 ;
        RECT 506.800 110.300 507.600 110.400 ;
        RECT 510.000 110.300 510.800 110.400 ;
        RECT 506.800 109.700 510.800 110.300 ;
        RECT 506.800 109.600 507.600 109.700 ;
        RECT 510.000 108.800 510.800 109.700 ;
        RECT 511.400 108.400 512.000 111.600 ;
        RECT 514.800 110.300 515.600 110.400 ;
        RECT 516.400 110.300 517.200 111.200 ;
        RECT 514.800 109.700 517.200 110.300 ;
        RECT 514.800 109.600 515.600 109.700 ;
        RECT 516.400 109.600 517.200 109.700 ;
        RECT 517.800 110.400 518.400 112.200 ;
        RECT 523.000 111.600 523.600 115.000 ;
        RECT 527.000 112.400 527.800 119.800 ;
        RECT 528.400 113.600 529.200 114.400 ;
        RECT 528.600 112.400 529.200 113.600 ;
        RECT 531.600 113.600 532.400 114.400 ;
        RECT 531.600 112.400 532.200 113.600 ;
        RECT 533.000 112.400 533.800 119.800 ;
        RECT 527.000 111.800 528.000 112.400 ;
        RECT 528.600 111.800 530.000 112.400 ;
        RECT 519.800 111.000 523.600 111.600 ;
        RECT 517.800 109.600 518.800 110.400 ;
        RECT 517.800 108.400 518.400 109.600 ;
        RECT 519.800 109.000 520.400 111.000 ;
        RECT 508.400 108.200 509.200 108.400 ;
        RECT 508.400 107.600 510.000 108.200 ;
        RECT 511.400 107.600 514.000 108.400 ;
        RECT 516.400 107.600 518.400 108.400 ;
        RECT 519.000 108.200 520.400 109.000 ;
        RECT 521.200 108.800 522.000 110.400 ;
        RECT 522.800 108.800 523.600 110.400 ;
        RECT 526.000 108.800 526.800 110.400 ;
        RECT 527.400 108.400 528.000 111.800 ;
        RECT 529.200 111.600 530.000 111.800 ;
        RECT 530.800 111.800 532.200 112.400 ;
        RECT 532.800 111.800 533.800 112.400 ;
        RECT 530.800 111.600 531.600 111.800 ;
        RECT 529.300 110.300 529.900 111.600 ;
        RECT 532.800 110.300 533.400 111.800 ;
        RECT 537.200 111.200 538.000 119.800 ;
        RECT 541.400 115.800 542.600 119.800 ;
        RECT 546.000 115.800 546.800 119.800 ;
        RECT 550.400 116.400 551.200 119.800 ;
        RECT 550.400 115.800 552.400 116.400 ;
        RECT 542.000 115.000 542.800 115.800 ;
        RECT 546.200 115.200 546.800 115.800 ;
        RECT 545.400 114.600 549.000 115.200 ;
        RECT 551.600 115.000 552.400 115.800 ;
        RECT 545.400 114.400 546.200 114.600 ;
        RECT 548.200 114.400 549.000 114.600 ;
        RECT 541.200 113.200 542.600 114.000 ;
        RECT 542.000 112.200 542.600 113.200 ;
        RECT 544.200 113.000 546.400 113.600 ;
        RECT 544.200 112.800 545.000 113.000 ;
        RECT 542.000 111.600 544.400 112.200 ;
        RECT 537.200 110.600 541.400 111.200 ;
        RECT 529.300 109.700 533.400 110.300 ;
        RECT 532.800 108.400 533.400 109.700 ;
        RECT 534.000 108.800 534.800 110.400 ;
        RECT 509.200 107.200 510.000 107.600 ;
        RECT 506.800 104.800 507.600 106.400 ;
        RECT 508.600 106.200 512.200 106.600 ;
        RECT 513.200 106.200 513.800 107.600 ;
        RECT 517.800 107.000 518.400 107.600 ;
        RECT 519.400 107.800 520.400 108.200 ;
        RECT 524.400 108.200 525.200 108.400 ;
        RECT 519.400 107.200 523.600 107.800 ;
        RECT 524.400 107.600 526.000 108.200 ;
        RECT 527.400 107.600 530.000 108.400 ;
        RECT 530.800 107.600 533.400 108.400 ;
        RECT 535.600 108.200 536.400 108.400 ;
        RECT 534.800 107.600 536.400 108.200 ;
        RECT 525.200 107.200 526.000 107.600 ;
        RECT 517.800 106.600 518.600 107.000 ;
        RECT 508.400 106.000 512.400 106.200 ;
        RECT 508.400 102.200 509.200 106.000 ;
        RECT 511.600 102.200 512.400 106.000 ;
        RECT 513.200 102.200 514.000 106.200 ;
        RECT 517.800 106.000 519.400 106.600 ;
        RECT 518.600 103.000 519.400 106.000 ;
        RECT 523.000 105.000 523.600 107.200 ;
        RECT 524.600 106.200 528.200 106.600 ;
        RECT 529.200 106.200 529.800 107.600 ;
        RECT 531.000 106.200 531.600 107.600 ;
        RECT 534.800 107.200 535.600 107.600 ;
        RECT 537.200 107.200 538.000 110.600 ;
        RECT 540.600 110.400 541.400 110.600 ;
        RECT 539.000 109.800 539.800 110.000 ;
        RECT 539.000 109.200 542.800 109.800 ;
        RECT 542.000 109.000 542.800 109.200 ;
        RECT 543.800 108.400 544.400 111.600 ;
        RECT 545.800 111.800 546.400 113.000 ;
        RECT 547.000 113.000 547.800 113.200 ;
        RECT 551.600 113.000 552.400 113.200 ;
        RECT 547.000 112.400 552.400 113.000 ;
        RECT 545.800 111.400 550.600 111.800 ;
        RECT 554.800 111.400 555.600 119.800 ;
        RECT 556.400 112.400 557.200 119.800 ;
        RECT 559.600 112.800 560.400 119.800 ;
        RECT 556.400 111.800 559.000 112.400 ;
        RECT 559.600 111.800 560.600 112.800 ;
        RECT 565.400 112.400 566.200 119.800 ;
        RECT 566.800 114.300 567.600 114.400 ;
        RECT 570.800 114.300 571.600 119.800 ;
        RECT 574.000 115.200 574.800 119.800 ;
        RECT 566.800 113.700 571.600 114.300 ;
        RECT 566.800 113.600 567.600 113.700 ;
        RECT 567.000 112.400 567.600 113.600 ;
        RECT 565.400 111.800 566.400 112.400 ;
        RECT 567.000 111.800 568.400 112.400 ;
        RECT 570.800 112.000 571.600 113.700 ;
        RECT 545.800 111.200 555.600 111.400 ;
        RECT 549.800 111.000 555.600 111.200 ;
        RECT 550.000 110.800 555.600 111.000 ;
        RECT 548.400 110.200 549.200 110.400 ;
        RECT 548.400 109.600 553.400 110.200 ;
        RECT 556.400 109.600 557.400 110.400 ;
        RECT 552.600 109.400 553.400 109.600 ;
        RECT 556.600 108.800 557.400 109.600 ;
        RECT 558.400 109.800 559.000 111.800 ;
        RECT 558.400 109.000 559.400 109.800 ;
        RECT 551.000 108.400 551.800 108.600 ;
        RECT 543.800 107.800 554.800 108.400 ;
        RECT 544.200 107.600 545.000 107.800 ;
        RECT 537.200 106.600 541.000 107.200 ;
        RECT 532.600 106.200 536.200 106.600 ;
        RECT 522.800 103.000 523.600 105.000 ;
        RECT 524.400 106.000 528.400 106.200 ;
        RECT 524.400 102.200 525.200 106.000 ;
        RECT 527.600 102.200 528.400 106.000 ;
        RECT 529.200 102.200 530.000 106.200 ;
        RECT 530.800 102.200 531.600 106.200 ;
        RECT 532.400 106.000 536.400 106.200 ;
        RECT 532.400 102.200 533.200 106.000 ;
        RECT 535.600 102.200 536.400 106.000 ;
        RECT 537.200 102.200 538.000 106.600 ;
        RECT 540.200 106.400 541.000 106.600 ;
        RECT 550.000 105.600 550.600 107.800 ;
        RECT 553.200 107.600 554.800 107.800 ;
        RECT 558.400 107.400 559.000 109.000 ;
        RECT 560.000 108.400 560.600 111.800 ;
        RECT 564.400 108.800 565.200 110.400 ;
        RECT 565.800 110.300 566.400 111.800 ;
        RECT 567.600 111.600 568.400 111.800 ;
        RECT 570.600 111.200 571.600 112.000 ;
        RECT 572.200 114.600 574.800 115.200 ;
        RECT 572.200 113.000 572.800 114.600 ;
        RECT 577.200 114.400 578.000 119.800 ;
        RECT 580.400 117.000 581.200 119.800 ;
        RECT 582.000 117.000 582.800 119.800 ;
        RECT 583.600 117.000 584.400 119.800 ;
        RECT 578.600 114.400 582.800 115.200 ;
        RECT 575.400 113.600 578.000 114.400 ;
        RECT 585.200 113.600 586.000 119.800 ;
        RECT 588.400 115.000 589.200 119.800 ;
        RECT 591.600 115.000 592.400 119.800 ;
        RECT 593.200 117.000 594.000 119.800 ;
        RECT 594.800 117.000 595.600 119.800 ;
        RECT 598.000 115.200 598.800 119.800 ;
        RECT 601.200 116.400 602.000 119.800 ;
        RECT 601.200 115.800 602.200 116.400 ;
        RECT 601.600 115.200 602.200 115.800 ;
        RECT 596.800 114.400 601.000 115.200 ;
        RECT 601.600 114.600 603.600 115.200 ;
        RECT 588.400 113.600 591.000 114.400 ;
        RECT 591.600 113.800 597.400 114.400 ;
        RECT 600.400 114.000 601.000 114.400 ;
        RECT 580.400 113.000 581.200 113.200 ;
        RECT 572.200 112.400 581.200 113.000 ;
        RECT 583.600 113.000 584.400 113.200 ;
        RECT 591.600 113.000 592.200 113.800 ;
        RECT 598.000 113.200 599.400 113.800 ;
        RECT 600.400 113.200 602.000 114.000 ;
        RECT 583.600 112.400 592.200 113.000 ;
        RECT 593.200 113.000 599.400 113.200 ;
        RECT 593.200 112.600 598.600 113.000 ;
        RECT 593.200 112.400 594.000 112.600 ;
        RECT 569.200 110.300 570.000 110.400 ;
        RECT 565.800 109.700 570.000 110.300 ;
        RECT 565.800 108.400 566.400 109.700 ;
        RECT 569.200 109.600 570.000 109.700 ;
        RECT 559.600 108.300 560.600 108.400 ;
        RECT 562.800 108.300 563.600 108.400 ;
        RECT 559.600 108.200 563.600 108.300 ;
        RECT 559.600 107.700 564.400 108.200 ;
        RECT 559.600 107.600 560.600 107.700 ;
        RECT 562.800 107.600 564.400 107.700 ;
        RECT 565.800 107.600 568.400 108.400 ;
        RECT 548.200 105.400 549.000 105.600 ;
        RECT 542.000 104.200 542.800 105.000 ;
        RECT 546.200 104.800 549.000 105.400 ;
        RECT 550.000 104.800 550.800 105.600 ;
        RECT 546.200 104.200 546.800 104.800 ;
        RECT 551.600 104.200 552.400 105.000 ;
        RECT 541.400 103.600 542.800 104.200 ;
        RECT 541.400 102.200 542.600 103.600 ;
        RECT 546.000 102.200 546.800 104.200 ;
        RECT 550.400 103.600 552.400 104.200 ;
        RECT 550.400 102.200 551.200 103.600 ;
        RECT 554.800 102.200 555.600 107.000 ;
        RECT 556.400 106.800 559.000 107.400 ;
        RECT 556.400 102.200 557.200 106.800 ;
        RECT 560.000 106.200 560.600 107.600 ;
        RECT 563.600 107.200 564.400 107.600 ;
        RECT 563.000 106.200 566.600 106.600 ;
        RECT 567.600 106.200 568.200 107.600 ;
        RECT 570.600 106.800 571.400 111.200 ;
        RECT 572.200 110.600 572.800 112.400 ;
        RECT 572.000 110.000 572.800 110.600 ;
        RECT 578.800 110.000 602.200 110.600 ;
        RECT 572.000 108.000 572.600 110.000 ;
        RECT 578.800 109.400 579.600 110.000 ;
        RECT 596.400 109.600 597.200 110.000 ;
        RECT 598.000 109.600 598.800 110.000 ;
        RECT 601.400 109.800 602.200 110.000 ;
        RECT 573.200 108.600 577.000 109.400 ;
        RECT 572.000 107.400 573.200 108.000 ;
        RECT 559.600 105.600 560.600 106.200 ;
        RECT 562.800 106.000 566.800 106.200 ;
        RECT 559.600 102.200 560.400 105.600 ;
        RECT 562.800 102.200 563.600 106.000 ;
        RECT 566.000 102.200 566.800 106.000 ;
        RECT 567.600 102.200 568.400 106.200 ;
        RECT 570.600 106.000 571.600 106.800 ;
        RECT 570.800 102.200 571.600 106.000 ;
        RECT 572.400 102.200 573.200 107.400 ;
        RECT 576.200 107.400 577.000 108.600 ;
        RECT 576.200 106.800 578.000 107.400 ;
        RECT 577.200 106.200 578.000 106.800 ;
        RECT 582.000 106.400 582.800 109.200 ;
        RECT 585.200 108.600 588.400 109.400 ;
        RECT 592.200 108.600 594.200 109.400 ;
        RECT 602.800 109.000 603.600 114.600 ;
        RECT 605.200 113.600 606.000 114.400 ;
        RECT 605.200 112.400 605.800 113.600 ;
        RECT 606.600 112.400 607.400 119.800 ;
        RECT 604.400 111.800 605.800 112.400 ;
        RECT 606.400 111.800 607.400 112.400 ;
        RECT 604.400 111.600 605.200 111.800 ;
        RECT 584.800 107.800 585.600 108.000 ;
        RECT 584.800 107.200 589.200 107.800 ;
        RECT 588.400 107.000 589.200 107.200 ;
        RECT 590.000 106.800 590.800 108.400 ;
        RECT 577.200 105.400 579.600 106.200 ;
        RECT 582.000 105.600 583.000 106.400 ;
        RECT 586.000 105.600 587.600 106.400 ;
        RECT 588.400 106.200 589.200 106.400 ;
        RECT 592.200 106.200 593.000 108.600 ;
        RECT 594.800 108.200 603.600 109.000 ;
        RECT 606.400 108.400 607.000 111.800 ;
        RECT 607.600 108.800 608.400 110.400 ;
        RECT 598.200 106.800 601.200 107.600 ;
        RECT 598.200 106.200 599.000 106.800 ;
        RECT 588.400 105.600 593.000 106.200 ;
        RECT 578.800 102.200 579.600 105.400 ;
        RECT 596.400 105.400 599.000 106.200 ;
        RECT 580.400 102.200 581.200 105.000 ;
        RECT 582.000 102.200 582.800 105.000 ;
        RECT 583.600 102.200 584.400 105.000 ;
        RECT 585.200 102.200 586.000 105.000 ;
        RECT 588.400 102.200 589.200 105.000 ;
        RECT 591.600 102.200 592.400 105.000 ;
        RECT 593.200 102.200 594.000 105.000 ;
        RECT 594.800 102.200 595.600 105.000 ;
        RECT 596.400 102.200 597.200 105.400 ;
        RECT 602.800 102.200 603.600 108.200 ;
        RECT 604.400 107.600 607.000 108.400 ;
        RECT 609.200 108.200 610.000 108.400 ;
        RECT 608.400 107.600 610.000 108.200 ;
        RECT 604.600 106.200 605.200 107.600 ;
        RECT 608.400 107.200 609.200 107.600 ;
        RECT 606.200 106.200 609.800 106.600 ;
        RECT 604.400 102.200 605.200 106.200 ;
        RECT 606.000 106.000 610.000 106.200 ;
        RECT 606.000 102.200 606.800 106.000 ;
        RECT 609.200 102.200 610.000 106.000 ;
        RECT 1.200 95.400 2.000 99.800 ;
        RECT 5.400 98.400 6.600 99.800 ;
        RECT 5.400 97.800 6.800 98.400 ;
        RECT 10.000 97.800 10.800 99.800 ;
        RECT 14.400 98.400 15.200 99.800 ;
        RECT 14.400 97.800 16.400 98.400 ;
        RECT 6.000 97.000 6.800 97.800 ;
        RECT 10.200 97.200 10.800 97.800 ;
        RECT 10.200 96.600 13.000 97.200 ;
        RECT 12.200 96.400 13.000 96.600 ;
        RECT 14.000 96.400 14.800 97.200 ;
        RECT 15.600 97.000 16.400 97.800 ;
        RECT 4.200 95.400 5.000 95.600 ;
        RECT 1.200 94.800 5.000 95.400 ;
        RECT 1.200 91.400 2.000 94.800 ;
        RECT 8.200 94.200 9.000 94.400 ;
        RECT 12.400 94.200 13.200 94.400 ;
        RECT 14.000 94.200 14.600 96.400 ;
        RECT 18.800 95.000 19.600 99.800 ;
        RECT 20.400 95.800 21.200 99.800 ;
        RECT 22.000 96.000 22.800 99.800 ;
        RECT 25.200 96.000 26.000 99.800 ;
        RECT 22.000 95.800 26.000 96.000 ;
        RECT 26.800 96.000 27.600 99.800 ;
        RECT 30.000 96.000 30.800 99.800 ;
        RECT 26.800 95.800 30.800 96.000 ;
        RECT 31.600 95.800 32.400 99.800 ;
        RECT 37.000 96.000 37.800 99.000 ;
        RECT 41.200 97.000 42.000 99.000 ;
        RECT 20.600 94.400 21.200 95.800 ;
        RECT 22.200 95.400 25.800 95.800 ;
        RECT 27.000 95.400 30.600 95.800 ;
        RECT 24.400 94.400 25.200 94.800 ;
        RECT 27.600 94.400 28.400 94.800 ;
        RECT 31.600 94.400 32.200 95.800 ;
        RECT 36.200 95.400 37.800 96.000 ;
        RECT 36.200 95.000 37.000 95.400 ;
        RECT 36.200 94.400 36.800 95.000 ;
        RECT 41.400 94.800 42.000 97.000 ;
        RECT 42.800 95.800 43.600 99.800 ;
        RECT 44.400 96.000 45.200 99.800 ;
        RECT 47.600 96.000 48.400 99.800 ;
        RECT 44.400 95.800 48.400 96.000 ;
        RECT 17.200 94.200 18.800 94.400 ;
        RECT 7.800 93.600 18.800 94.200 ;
        RECT 20.400 93.600 23.000 94.400 ;
        RECT 24.400 93.800 26.000 94.400 ;
        RECT 25.200 93.600 26.000 93.800 ;
        RECT 26.800 93.800 28.400 94.400 ;
        RECT 26.800 93.600 27.600 93.800 ;
        RECT 29.800 93.600 32.400 94.400 ;
        RECT 34.800 93.600 36.800 94.400 ;
        RECT 37.800 94.200 42.000 94.800 ;
        RECT 43.000 94.400 43.600 95.800 ;
        RECT 44.600 95.400 48.200 95.800 ;
        RECT 49.200 95.000 50.000 99.800 ;
        RECT 53.600 98.400 54.400 99.800 ;
        RECT 52.400 97.800 54.400 98.400 ;
        RECT 58.000 97.800 58.800 99.800 ;
        RECT 62.200 98.400 63.400 99.800 ;
        RECT 62.000 97.800 63.400 98.400 ;
        RECT 52.400 97.000 53.200 97.800 ;
        RECT 58.000 97.200 58.600 97.800 ;
        RECT 54.000 96.400 54.800 97.200 ;
        RECT 55.800 96.600 58.600 97.200 ;
        RECT 62.000 97.000 62.800 97.800 ;
        RECT 55.800 96.400 56.600 96.600 ;
        RECT 46.800 94.400 47.600 94.800 ;
        RECT 37.800 93.800 38.800 94.200 ;
        RECT 6.000 92.800 6.800 93.000 ;
        RECT 3.000 92.200 6.800 92.800 ;
        RECT 3.000 92.000 3.800 92.200 ;
        RECT 4.600 91.400 5.400 91.600 ;
        RECT 1.200 90.800 5.400 91.400 ;
        RECT 1.200 82.200 2.000 90.800 ;
        RECT 7.800 90.400 8.400 93.600 ;
        RECT 15.000 93.400 15.800 93.600 ;
        RECT 14.000 92.400 14.800 92.600 ;
        RECT 16.600 92.400 17.400 92.600 ;
        RECT 12.400 91.800 17.400 92.400 ;
        RECT 12.400 91.600 13.200 91.800 ;
        RECT 14.000 91.000 19.600 91.200 ;
        RECT 13.800 90.800 19.600 91.000 ;
        RECT 6.000 89.800 8.400 90.400 ;
        RECT 9.800 90.600 19.600 90.800 ;
        RECT 9.800 90.200 14.600 90.600 ;
        RECT 6.000 88.800 6.600 89.800 ;
        RECT 5.200 88.000 6.600 88.800 ;
        RECT 8.200 89.000 9.000 89.200 ;
        RECT 9.800 89.000 10.400 90.200 ;
        RECT 8.200 88.400 10.400 89.000 ;
        RECT 11.000 89.000 16.400 89.600 ;
        RECT 11.000 88.800 11.800 89.000 ;
        RECT 15.600 88.800 16.400 89.000 ;
        RECT 9.400 87.400 10.200 87.600 ;
        RECT 12.200 87.400 13.000 87.600 ;
        RECT 6.000 86.200 6.800 87.000 ;
        RECT 9.400 86.800 13.000 87.400 ;
        RECT 10.200 86.200 10.800 86.800 ;
        RECT 15.600 86.200 16.400 87.000 ;
        RECT 5.400 82.200 6.600 86.200 ;
        RECT 10.000 82.200 10.800 86.200 ;
        RECT 14.400 85.600 16.400 86.200 ;
        RECT 14.400 82.200 15.200 85.600 ;
        RECT 18.800 82.200 19.600 90.600 ;
        RECT 20.400 90.200 21.200 90.400 ;
        RECT 22.400 90.200 23.000 93.600 ;
        RECT 23.600 91.600 24.400 93.200 ;
        RECT 28.400 91.600 29.200 93.200 ;
        RECT 29.800 90.400 30.400 93.600 ;
        RECT 36.200 92.400 36.800 93.600 ;
        RECT 37.400 93.000 38.800 93.800 ;
        RECT 42.800 93.600 45.400 94.400 ;
        RECT 46.800 93.800 48.400 94.400 ;
        RECT 47.600 93.600 48.400 93.800 ;
        RECT 50.000 94.200 51.600 94.400 ;
        RECT 54.200 94.200 54.800 96.400 ;
        RECT 63.800 95.400 64.600 95.600 ;
        RECT 66.800 95.400 67.600 99.800 ;
        RECT 68.400 95.600 69.200 99.800 ;
        RECT 70.000 96.000 70.800 99.800 ;
        RECT 73.200 96.000 74.000 99.800 ;
        RECT 70.000 95.800 74.000 96.000 ;
        RECT 74.800 97.000 75.600 99.000 ;
        RECT 63.800 94.800 67.600 95.400 ;
        RECT 55.600 94.200 56.400 94.400 ;
        RECT 59.800 94.200 60.600 94.400 ;
        RECT 50.000 93.600 61.000 94.200 ;
        RECT 34.800 90.800 35.600 92.400 ;
        RECT 36.200 91.600 37.200 92.400 ;
        RECT 20.400 89.600 21.800 90.200 ;
        RECT 22.400 89.600 23.400 90.200 ;
        RECT 28.400 89.600 30.400 90.400 ;
        RECT 31.600 90.200 32.400 90.400 ;
        RECT 31.000 89.600 32.400 90.200 ;
        RECT 36.200 89.800 36.800 91.600 ;
        RECT 38.200 91.000 38.800 93.000 ;
        RECT 39.600 91.600 40.400 93.200 ;
        RECT 41.200 91.600 42.000 93.200 ;
        RECT 38.200 90.400 42.000 91.000 ;
        RECT 21.200 88.400 21.800 89.600 ;
        RECT 21.200 87.600 22.000 88.400 ;
        RECT 22.600 84.400 23.400 89.600 ;
        RECT 22.600 83.600 24.400 84.400 ;
        RECT 22.600 82.200 23.400 83.600 ;
        RECT 29.400 82.200 30.200 89.600 ;
        RECT 31.000 88.400 31.600 89.600 ;
        RECT 36.200 89.200 37.800 89.800 ;
        RECT 30.800 87.600 31.600 88.400 ;
        RECT 37.000 82.200 37.800 89.200 ;
        RECT 41.400 87.000 42.000 90.400 ;
        RECT 42.800 90.200 43.600 90.400 ;
        RECT 44.800 90.200 45.400 93.600 ;
        RECT 53.000 93.400 53.800 93.600 ;
        RECT 46.000 91.600 46.800 93.200 ;
        RECT 51.400 92.400 52.200 92.600 ;
        RECT 51.400 92.300 56.400 92.400 ;
        RECT 58.800 92.300 59.600 92.400 ;
        RECT 51.400 91.800 59.600 92.300 ;
        RECT 55.600 91.700 59.600 91.800 ;
        RECT 55.600 91.600 56.400 91.700 ;
        RECT 58.800 91.600 59.600 91.700 ;
        RECT 49.200 91.000 54.800 91.200 ;
        RECT 49.200 90.800 55.000 91.000 ;
        RECT 49.200 90.600 59.000 90.800 ;
        RECT 42.800 89.600 44.200 90.200 ;
        RECT 44.800 89.600 45.800 90.200 ;
        RECT 43.600 88.400 44.200 89.600 ;
        RECT 43.600 87.600 44.400 88.400 ;
        RECT 41.200 83.000 42.000 87.000 ;
        RECT 45.000 82.200 45.800 89.600 ;
        RECT 49.200 82.200 50.000 90.600 ;
        RECT 54.200 90.200 59.000 90.600 ;
        RECT 52.400 89.000 57.800 89.600 ;
        RECT 52.400 88.800 53.200 89.000 ;
        RECT 57.000 88.800 57.800 89.000 ;
        RECT 58.400 89.000 59.000 90.200 ;
        RECT 60.400 90.400 61.000 93.600 ;
        RECT 62.000 92.800 62.800 93.000 ;
        RECT 62.000 92.200 65.800 92.800 ;
        RECT 65.000 92.000 65.800 92.200 ;
        RECT 63.400 91.400 64.200 91.600 ;
        RECT 66.800 91.400 67.600 94.800 ;
        RECT 68.600 94.400 69.200 95.600 ;
        RECT 70.200 95.400 73.800 95.800 ;
        RECT 74.800 94.800 75.400 97.000 ;
        RECT 79.000 96.400 79.800 99.000 ;
        RECT 79.000 96.000 80.400 96.400 ;
        RECT 79.000 95.400 80.600 96.000 ;
        RECT 84.400 95.800 85.200 99.800 ;
        RECT 86.000 96.000 86.800 99.800 ;
        RECT 89.200 96.000 90.000 99.800 ;
        RECT 86.000 95.800 90.000 96.000 ;
        RECT 79.800 95.000 80.600 95.400 ;
        RECT 72.400 94.400 73.200 94.800 ;
        RECT 68.400 93.600 71.000 94.400 ;
        RECT 72.400 93.800 74.000 94.400 ;
        RECT 74.800 94.200 79.000 94.800 ;
        RECT 73.200 93.600 74.000 93.800 ;
        RECT 78.000 93.800 79.000 94.200 ;
        RECT 80.000 94.400 80.600 95.000 ;
        RECT 84.600 94.400 85.200 95.800 ;
        RECT 86.200 95.400 89.800 95.800 ;
        RECT 88.400 94.400 89.200 94.800 ;
        RECT 63.400 90.800 67.600 91.400 ;
        RECT 60.400 89.800 62.800 90.400 ;
        RECT 59.800 89.000 60.600 89.200 ;
        RECT 58.400 88.400 60.600 89.000 ;
        RECT 62.200 88.800 62.800 89.800 ;
        RECT 62.200 88.000 63.600 88.800 ;
        RECT 55.800 87.400 56.600 87.600 ;
        RECT 58.600 87.400 59.400 87.600 ;
        RECT 52.400 86.200 53.200 87.000 ;
        RECT 55.800 86.800 59.400 87.400 ;
        RECT 58.000 86.200 58.600 86.800 ;
        RECT 62.000 86.200 62.800 87.000 ;
        RECT 52.400 85.600 54.400 86.200 ;
        RECT 53.600 82.200 54.400 85.600 ;
        RECT 58.000 82.200 58.800 86.200 ;
        RECT 62.200 82.200 63.400 86.200 ;
        RECT 66.800 82.200 67.600 90.800 ;
        RECT 68.400 90.200 69.200 90.400 ;
        RECT 70.400 90.200 71.000 93.600 ;
        RECT 71.600 91.600 72.400 93.200 ;
        RECT 74.800 91.600 75.600 93.200 ;
        RECT 76.400 91.600 77.200 93.200 ;
        RECT 78.000 93.000 79.400 93.800 ;
        RECT 80.000 93.600 82.000 94.400 ;
        RECT 84.400 93.600 87.000 94.400 ;
        RECT 88.400 93.800 90.000 94.400 ;
        RECT 94.400 94.200 95.200 99.800 ;
        RECT 97.200 95.800 98.000 99.800 ;
        RECT 98.800 96.000 99.600 99.800 ;
        RECT 102.000 96.000 102.800 99.800 ;
        RECT 98.800 95.800 102.800 96.000 ;
        RECT 97.400 94.400 98.000 95.800 ;
        RECT 99.000 95.400 102.600 95.800 ;
        RECT 101.200 94.400 102.000 94.800 ;
        RECT 94.400 93.800 96.200 94.200 ;
        RECT 89.200 93.600 90.000 93.800 ;
        RECT 94.600 93.600 96.200 93.800 ;
        RECT 97.200 93.600 99.800 94.400 ;
        RECT 101.200 93.800 102.800 94.400 ;
        RECT 107.200 94.200 108.000 99.800 ;
        RECT 111.600 97.800 112.400 99.800 ;
        RECT 111.600 94.400 112.200 97.800 ;
        RECT 113.200 95.600 114.000 97.200 ;
        RECT 114.800 95.800 115.600 99.800 ;
        RECT 116.400 96.000 117.200 99.800 ;
        RECT 119.600 96.000 120.400 99.800 ;
        RECT 121.800 98.400 122.600 99.800 ;
        RECT 121.200 97.600 122.600 98.400 ;
        RECT 116.400 95.800 120.400 96.000 ;
        RECT 121.800 96.400 122.600 97.600 ;
        RECT 121.800 95.800 123.600 96.400 ;
        RECT 129.800 96.000 130.600 99.000 ;
        RECT 134.000 97.000 134.800 99.000 ;
        RECT 115.000 94.400 115.600 95.800 ;
        RECT 116.600 95.400 120.200 95.800 ;
        RECT 118.800 94.400 119.600 94.800 ;
        RECT 107.200 93.800 109.000 94.200 ;
        RECT 102.000 93.600 102.800 93.800 ;
        RECT 107.400 93.600 109.000 93.800 ;
        RECT 78.000 91.000 78.600 93.000 ;
        RECT 74.800 90.400 78.600 91.000 ;
        RECT 68.400 89.600 69.800 90.200 ;
        RECT 70.400 89.600 71.400 90.200 ;
        RECT 69.200 88.400 69.800 89.600 ;
        RECT 69.200 87.600 70.000 88.400 ;
        RECT 70.600 82.200 71.400 89.600 ;
        RECT 74.800 87.000 75.400 90.400 ;
        RECT 80.000 89.800 80.600 93.600 ;
        RECT 81.200 92.300 82.000 92.400 ;
        RECT 86.400 92.300 87.000 93.600 ;
        RECT 81.200 91.700 87.000 92.300 ;
        RECT 81.200 90.800 82.000 91.700 ;
        RECT 79.000 89.200 80.600 89.800 ;
        RECT 84.400 90.200 85.200 90.400 ;
        RECT 86.400 90.200 87.000 91.700 ;
        RECT 87.600 91.600 88.400 93.200 ;
        RECT 92.400 91.600 94.000 92.400 ;
        RECT 84.400 89.600 85.800 90.200 ;
        RECT 86.400 89.600 87.400 90.200 ;
        RECT 90.800 89.600 91.600 91.200 ;
        RECT 95.600 90.400 96.200 93.600 ;
        RECT 95.600 90.300 96.400 90.400 ;
        RECT 97.200 90.300 98.000 90.400 ;
        RECT 95.600 90.200 98.000 90.300 ;
        RECT 99.200 90.200 99.800 93.600 ;
        RECT 100.400 91.600 101.200 93.200 ;
        RECT 105.200 91.600 106.800 92.400 ;
        RECT 95.600 89.700 98.600 90.200 ;
        RECT 95.600 89.600 96.400 89.700 ;
        RECT 97.200 89.600 98.600 89.700 ;
        RECT 99.200 89.600 100.200 90.200 ;
        RECT 103.600 89.600 104.400 91.200 ;
        RECT 108.400 90.400 109.000 93.600 ;
        RECT 111.600 93.600 112.400 94.400 ;
        RECT 114.800 93.600 117.400 94.400 ;
        RECT 118.800 93.800 120.400 94.400 ;
        RECT 119.600 93.600 120.400 93.800 ;
        RECT 110.000 90.800 110.800 92.400 ;
        RECT 111.600 90.400 112.200 93.600 ;
        RECT 108.400 89.600 109.200 90.400 ;
        RECT 111.600 90.200 112.400 90.400 ;
        RECT 74.800 83.000 75.600 87.000 ;
        RECT 79.000 82.200 79.800 89.200 ;
        RECT 85.200 88.400 85.800 89.600 ;
        RECT 85.200 87.600 86.000 88.400 ;
        RECT 86.600 84.400 87.400 89.600 ;
        RECT 94.000 87.600 94.800 89.200 ;
        RECT 95.600 87.000 96.200 89.600 ;
        RECT 98.000 88.400 98.600 89.600 ;
        RECT 98.000 87.600 98.800 88.400 ;
        RECT 92.600 86.400 96.200 87.000 ;
        RECT 92.600 86.200 93.200 86.400 ;
        RECT 86.600 83.600 88.400 84.400 ;
        RECT 86.600 82.200 87.400 83.600 ;
        RECT 92.400 82.200 93.200 86.200 ;
        RECT 95.600 86.200 96.200 86.400 ;
        RECT 95.600 82.200 96.400 86.200 ;
        RECT 99.400 82.200 100.200 89.600 ;
        RECT 106.800 87.600 107.600 89.200 ;
        RECT 108.400 88.400 109.000 89.600 ;
        RECT 110.600 89.400 112.400 90.200 ;
        RECT 114.800 90.200 115.600 90.400 ;
        RECT 116.800 90.200 117.400 93.600 ;
        RECT 118.000 91.600 118.800 93.200 ;
        RECT 114.800 89.600 116.200 90.200 ;
        RECT 116.800 89.600 117.800 90.200 ;
        RECT 108.400 87.600 109.200 88.400 ;
        RECT 108.400 87.000 109.000 87.600 ;
        RECT 105.400 86.400 109.000 87.000 ;
        RECT 105.400 86.200 106.000 86.400 ;
        RECT 105.200 82.200 106.000 86.200 ;
        RECT 108.400 86.200 109.000 86.400 ;
        RECT 108.400 82.200 109.200 86.200 ;
        RECT 110.600 82.200 111.400 89.400 ;
        RECT 115.600 88.400 116.200 89.600 ;
        RECT 115.600 87.600 116.400 88.400 ;
        RECT 117.000 82.200 117.800 89.600 ;
        RECT 121.200 88.800 122.000 90.400 ;
        RECT 122.800 82.200 123.600 95.800 ;
        RECT 129.000 95.400 130.600 96.000 ;
        RECT 124.400 93.600 125.200 95.200 ;
        RECT 129.000 95.000 129.800 95.400 ;
        RECT 129.000 94.400 129.600 95.000 ;
        RECT 134.200 94.800 134.800 97.000 ;
        RECT 135.600 96.000 136.400 99.800 ;
        RECT 138.800 96.000 139.600 99.800 ;
        RECT 135.600 95.800 139.600 96.000 ;
        RECT 140.400 95.800 141.200 99.800 ;
        RECT 142.600 98.400 143.400 99.800 ;
        RECT 142.600 97.600 144.400 98.400 ;
        RECT 142.600 96.400 143.400 97.600 ;
        RECT 142.600 95.800 144.400 96.400 ;
        RECT 135.800 95.400 139.400 95.800 ;
        RECT 127.600 93.600 129.600 94.400 ;
        RECT 130.600 94.200 134.800 94.800 ;
        RECT 136.400 94.400 137.200 94.800 ;
        RECT 140.400 94.400 141.000 95.800 ;
        RECT 130.600 93.800 131.600 94.200 ;
        RECT 126.000 92.300 126.800 92.400 ;
        RECT 127.600 92.300 128.400 92.400 ;
        RECT 126.000 91.700 128.400 92.300 ;
        RECT 126.000 91.600 126.800 91.700 ;
        RECT 127.600 90.800 128.400 91.700 ;
        RECT 129.000 89.800 129.600 93.600 ;
        RECT 130.200 93.000 131.600 93.800 ;
        RECT 135.600 93.800 137.200 94.400 ;
        RECT 135.600 93.600 136.400 93.800 ;
        RECT 138.600 93.600 141.200 94.400 ;
        RECT 131.000 91.000 131.600 93.000 ;
        RECT 132.400 91.600 133.200 93.200 ;
        RECT 134.000 92.300 134.800 93.200 ;
        RECT 135.600 92.300 136.400 92.400 ;
        RECT 134.000 91.700 136.400 92.300 ;
        RECT 134.000 91.600 134.800 91.700 ;
        RECT 135.600 91.600 136.400 91.700 ;
        RECT 137.200 91.600 138.000 93.200 ;
        RECT 131.000 90.400 134.800 91.000 ;
        RECT 129.000 89.200 130.600 89.800 ;
        RECT 129.800 84.400 130.600 89.200 ;
        RECT 134.200 87.000 134.800 90.400 ;
        RECT 138.600 90.200 139.200 93.600 ;
        RECT 140.400 90.200 141.200 90.400 ;
        RECT 129.800 83.600 131.600 84.400 ;
        RECT 129.800 82.200 130.600 83.600 ;
        RECT 134.000 83.000 134.800 87.000 ;
        RECT 138.200 89.600 139.200 90.200 ;
        RECT 139.800 89.600 141.200 90.200 ;
        RECT 138.200 82.200 139.000 89.600 ;
        RECT 139.800 88.400 140.400 89.600 ;
        RECT 142.000 88.800 142.800 90.400 ;
        RECT 139.600 87.600 140.400 88.400 ;
        RECT 143.600 82.200 144.400 95.800 ;
        RECT 145.200 93.600 146.000 95.200 ;
        RECT 148.000 94.200 148.800 99.800 ;
        RECT 147.000 93.800 148.800 94.200 ;
        RECT 158.000 95.400 158.800 99.800 ;
        RECT 162.200 98.400 163.400 99.800 ;
        RECT 162.200 97.800 163.600 98.400 ;
        RECT 166.800 97.800 167.600 99.800 ;
        RECT 171.200 98.400 172.000 99.800 ;
        RECT 171.200 97.800 173.200 98.400 ;
        RECT 162.800 97.000 163.600 97.800 ;
        RECT 167.000 97.200 167.600 97.800 ;
        RECT 167.000 96.600 169.800 97.200 ;
        RECT 169.000 96.400 169.800 96.600 ;
        RECT 170.800 96.400 171.600 97.200 ;
        RECT 172.400 97.000 173.200 97.800 ;
        RECT 161.000 95.400 161.800 95.600 ;
        RECT 158.000 94.800 161.800 95.400 ;
        RECT 147.000 93.600 148.600 93.800 ;
        RECT 147.000 90.400 147.600 93.600 ;
        RECT 149.200 91.600 150.800 92.400 ;
        RECT 158.000 91.400 158.800 94.800 ;
        RECT 165.000 94.200 165.800 94.400 ;
        RECT 169.200 94.200 170.000 94.400 ;
        RECT 170.800 94.200 171.400 96.400 ;
        RECT 175.600 95.000 176.400 99.800 ;
        RECT 174.000 94.200 175.600 94.400 ;
        RECT 164.600 93.600 175.600 94.200 ;
        RECT 177.200 93.800 178.000 99.800 ;
        RECT 183.600 96.600 184.400 99.800 ;
        RECT 185.200 97.000 186.000 99.800 ;
        RECT 186.800 97.000 187.600 99.800 ;
        RECT 188.400 97.000 189.200 99.800 ;
        RECT 191.600 97.000 192.400 99.800 ;
        RECT 194.800 97.000 195.600 99.800 ;
        RECT 196.400 97.000 197.200 99.800 ;
        RECT 198.000 97.000 198.800 99.800 ;
        RECT 199.600 97.000 200.400 99.800 ;
        RECT 181.800 95.800 184.400 96.600 ;
        RECT 201.200 96.600 202.000 99.800 ;
        RECT 187.800 95.800 192.400 96.400 ;
        RECT 181.800 95.200 182.600 95.800 ;
        RECT 179.600 94.400 182.600 95.200 ;
        RECT 162.800 92.800 163.600 93.000 ;
        RECT 159.800 92.200 163.600 92.800 ;
        RECT 159.800 92.000 160.600 92.200 ;
        RECT 161.400 91.400 162.200 91.600 ;
        RECT 146.800 89.600 147.600 90.400 ;
        RECT 151.600 90.300 152.400 91.200 ;
        RECT 158.000 90.800 162.200 91.400 ;
        RECT 158.000 90.300 158.800 90.800 ;
        RECT 164.600 90.400 165.200 93.600 ;
        RECT 171.800 93.400 172.600 93.600 ;
        RECT 177.200 93.000 186.000 93.800 ;
        RECT 187.800 93.400 188.600 95.800 ;
        RECT 191.600 95.600 192.400 95.800 ;
        RECT 193.200 95.600 194.800 96.400 ;
        RECT 197.800 95.600 198.800 96.400 ;
        RECT 201.200 95.800 203.600 96.600 ;
        RECT 190.000 93.600 190.800 95.200 ;
        RECT 191.600 94.800 192.400 95.000 ;
        RECT 191.600 94.200 196.000 94.800 ;
        RECT 195.200 94.000 196.000 94.200 ;
        RECT 170.800 92.400 171.600 92.600 ;
        RECT 173.400 92.400 174.200 92.600 ;
        RECT 169.200 91.800 174.200 92.400 ;
        RECT 169.200 91.600 170.000 91.800 ;
        RECT 170.800 91.000 176.400 91.200 ;
        RECT 170.600 90.800 176.400 91.000 ;
        RECT 151.600 89.700 158.800 90.300 ;
        RECT 151.600 89.600 152.400 89.700 ;
        RECT 147.000 88.400 147.600 89.600 ;
        RECT 146.800 87.600 147.600 88.400 ;
        RECT 148.400 87.600 149.200 89.200 ;
        RECT 147.000 87.000 147.600 87.600 ;
        RECT 147.000 86.400 150.600 87.000 ;
        RECT 147.000 86.200 147.600 86.400 ;
        RECT 146.800 82.200 147.600 86.200 ;
        RECT 150.000 86.200 150.600 86.400 ;
        RECT 150.000 82.200 150.800 86.200 ;
        RECT 158.000 82.200 158.800 89.700 ;
        RECT 162.800 89.800 165.200 90.400 ;
        RECT 166.600 90.600 176.400 90.800 ;
        RECT 166.600 90.200 171.400 90.600 ;
        RECT 162.800 88.800 163.400 89.800 ;
        RECT 162.000 88.000 163.400 88.800 ;
        RECT 165.000 89.000 165.800 89.200 ;
        RECT 166.600 89.000 167.200 90.200 ;
        RECT 165.000 88.400 167.200 89.000 ;
        RECT 167.800 89.000 173.200 89.600 ;
        RECT 167.800 88.800 168.600 89.000 ;
        RECT 172.400 88.800 173.200 89.000 ;
        RECT 166.200 87.400 167.000 87.600 ;
        RECT 169.000 87.400 169.800 87.600 ;
        RECT 162.800 86.200 163.600 87.000 ;
        RECT 166.200 86.800 169.800 87.400 ;
        RECT 167.000 86.200 167.600 86.800 ;
        RECT 172.400 86.200 173.200 87.000 ;
        RECT 162.200 82.200 163.400 86.200 ;
        RECT 166.800 82.200 167.600 86.200 ;
        RECT 171.200 85.600 173.200 86.200 ;
        RECT 171.200 82.200 172.000 85.600 ;
        RECT 175.600 82.200 176.400 90.600 ;
        RECT 177.200 87.400 178.000 93.000 ;
        RECT 186.600 92.600 188.600 93.400 ;
        RECT 192.400 92.600 195.600 93.400 ;
        RECT 198.000 92.800 198.800 95.600 ;
        RECT 202.800 95.200 203.600 95.800 ;
        RECT 202.800 94.600 204.600 95.200 ;
        RECT 203.800 93.400 204.600 94.600 ;
        RECT 207.600 94.600 208.400 99.800 ;
        RECT 209.200 96.000 210.000 99.800 ;
        RECT 209.200 95.200 210.200 96.000 ;
        RECT 212.400 95.800 213.200 99.800 ;
        RECT 214.000 96.000 214.800 99.800 ;
        RECT 217.200 96.000 218.000 99.800 ;
        RECT 221.400 96.400 222.200 99.800 ;
        RECT 224.200 98.400 225.000 99.800 ;
        RECT 223.600 97.600 225.000 98.400 ;
        RECT 214.000 95.800 218.000 96.000 ;
        RECT 220.400 95.800 222.200 96.400 ;
        RECT 224.200 96.400 225.000 97.600 ;
        RECT 229.000 96.800 229.800 99.800 ;
        RECT 224.200 95.800 226.000 96.400 ;
        RECT 207.600 94.000 208.800 94.600 ;
        RECT 203.800 92.600 207.600 93.400 ;
        RECT 178.600 92.000 179.400 92.200 ;
        RECT 182.000 92.000 182.800 92.400 ;
        RECT 183.600 92.000 184.400 92.400 ;
        RECT 201.200 92.000 202.000 92.600 ;
        RECT 208.200 92.000 208.800 94.000 ;
        RECT 178.600 91.400 202.000 92.000 ;
        RECT 208.000 91.400 208.800 92.000 ;
        RECT 208.000 89.600 208.600 91.400 ;
        RECT 209.400 90.800 210.200 95.200 ;
        RECT 212.600 94.400 213.200 95.800 ;
        RECT 214.200 95.400 217.800 95.800 ;
        RECT 216.400 94.400 217.200 94.800 ;
        RECT 212.400 93.600 215.000 94.400 ;
        RECT 216.400 93.800 218.000 94.400 ;
        RECT 217.200 93.600 218.000 93.800 ;
        RECT 218.800 93.600 219.600 95.200 ;
        RECT 186.800 89.400 187.600 89.600 ;
        RECT 182.200 89.000 187.600 89.400 ;
        RECT 181.400 88.800 187.600 89.000 ;
        RECT 188.600 89.000 197.200 89.600 ;
        RECT 178.800 88.000 180.400 88.800 ;
        RECT 181.400 88.200 182.800 88.800 ;
        RECT 188.600 88.200 189.200 89.000 ;
        RECT 196.400 88.800 197.200 89.000 ;
        RECT 199.600 89.000 208.600 89.600 ;
        RECT 199.600 88.800 200.400 89.000 ;
        RECT 179.800 87.600 180.400 88.000 ;
        RECT 183.400 87.600 189.200 88.200 ;
        RECT 189.800 87.600 192.400 88.400 ;
        RECT 177.200 86.800 179.200 87.400 ;
        RECT 179.800 86.800 184.000 87.600 ;
        RECT 178.600 86.200 179.200 86.800 ;
        RECT 178.600 85.600 179.600 86.200 ;
        RECT 178.800 82.200 179.600 85.600 ;
        RECT 182.000 82.200 182.800 86.800 ;
        RECT 185.200 82.200 186.000 85.000 ;
        RECT 186.800 82.200 187.600 85.000 ;
        RECT 188.400 82.200 189.200 87.000 ;
        RECT 191.600 82.200 192.400 87.000 ;
        RECT 194.800 82.200 195.600 88.400 ;
        RECT 202.800 87.600 205.400 88.400 ;
        RECT 198.000 86.800 202.200 87.600 ;
        RECT 196.400 82.200 197.200 85.000 ;
        RECT 198.000 82.200 198.800 85.000 ;
        RECT 199.600 82.200 200.400 85.000 ;
        RECT 202.800 82.200 203.600 87.600 ;
        RECT 208.000 87.400 208.600 89.000 ;
        RECT 206.000 86.800 208.600 87.400 ;
        RECT 209.200 90.000 210.200 90.800 ;
        RECT 214.400 90.400 215.000 93.600 ;
        RECT 215.600 91.600 216.400 93.200 ;
        RECT 220.400 92.300 221.200 95.800 ;
        RECT 220.400 91.700 224.300 92.300 ;
        RECT 212.400 90.200 213.200 90.400 ;
        RECT 206.000 82.200 206.800 86.800 ;
        RECT 209.200 82.200 210.000 90.000 ;
        RECT 212.400 89.600 213.800 90.200 ;
        RECT 214.400 89.600 216.400 90.400 ;
        RECT 213.200 88.400 213.800 89.600 ;
        RECT 213.200 87.600 214.000 88.400 ;
        RECT 214.600 82.200 215.400 89.600 ;
        RECT 220.400 82.200 221.200 91.700 ;
        RECT 223.700 90.400 224.300 91.700 ;
        RECT 222.000 88.800 222.800 90.400 ;
        RECT 223.600 88.800 224.400 90.400 ;
        RECT 225.200 82.200 226.000 95.800 ;
        RECT 228.400 95.800 229.800 96.800 ;
        RECT 233.200 95.800 234.000 99.800 ;
        RECT 235.400 96.400 236.200 99.800 ;
        RECT 235.400 95.800 237.200 96.400 ;
        RECT 239.600 96.000 240.400 99.800 ;
        RECT 242.800 96.000 243.600 99.800 ;
        RECT 239.600 95.800 243.600 96.000 ;
        RECT 244.400 96.300 245.200 99.800 ;
        RECT 246.000 96.300 246.800 97.200 ;
        RECT 226.800 93.600 227.600 95.200 ;
        RECT 228.400 92.400 229.000 95.800 ;
        RECT 233.200 95.600 233.800 95.800 ;
        RECT 232.000 95.200 233.800 95.600 ;
        RECT 229.600 95.000 233.800 95.200 ;
        RECT 229.600 94.600 232.600 95.000 ;
        RECT 229.600 94.400 230.400 94.600 ;
        RECT 226.800 92.300 227.600 92.400 ;
        RECT 228.400 92.300 229.200 92.400 ;
        RECT 226.800 91.700 229.200 92.300 ;
        RECT 226.800 91.600 227.600 91.700 ;
        RECT 228.400 91.600 229.200 91.700 ;
        RECT 228.400 90.200 229.000 91.600 ;
        RECT 229.800 91.000 230.400 94.400 ;
        RECT 233.200 94.300 234.000 94.400 ;
        RECT 234.800 94.300 235.600 94.400 ;
        RECT 231.200 93.200 232.400 94.000 ;
        RECT 233.200 93.700 235.600 94.300 ;
        RECT 231.600 92.400 232.200 93.200 ;
        RECT 233.200 92.800 234.000 93.700 ;
        RECT 234.800 93.600 235.600 93.700 ;
        RECT 231.600 91.600 232.400 92.400 ;
        RECT 236.400 92.300 237.200 95.800 ;
        RECT 239.800 95.400 243.400 95.800 ;
        RECT 244.400 95.700 246.800 96.300 ;
        RECT 238.000 93.600 238.800 95.200 ;
        RECT 240.400 94.400 241.200 94.800 ;
        RECT 244.400 94.400 245.000 95.700 ;
        RECT 246.000 95.600 246.800 95.700 ;
        RECT 239.600 93.800 241.200 94.400 ;
        RECT 239.600 93.600 240.400 93.800 ;
        RECT 242.600 93.600 245.200 94.400 ;
        RECT 239.600 92.300 240.400 92.400 ;
        RECT 236.400 91.700 240.400 92.300 ;
        RECT 229.800 90.400 232.200 91.000 ;
        RECT 228.400 82.200 229.200 90.200 ;
        RECT 231.600 86.200 232.200 90.400 ;
        RECT 234.800 88.800 235.600 90.400 ;
        RECT 231.600 82.200 232.400 86.200 ;
        RECT 236.400 82.200 237.200 91.700 ;
        RECT 239.600 91.600 240.400 91.700 ;
        RECT 241.200 91.600 242.000 93.200 ;
        RECT 242.600 90.200 243.200 93.600 ;
        RECT 244.400 90.200 245.200 90.400 ;
        RECT 242.200 89.600 243.200 90.200 ;
        RECT 243.800 89.600 245.200 90.200 ;
        RECT 242.200 82.200 243.000 89.600 ;
        RECT 243.800 88.400 244.400 89.600 ;
        RECT 243.600 87.600 244.400 88.400 ;
        RECT 247.600 82.200 248.400 99.800 ;
        RECT 250.800 96.000 251.600 99.800 ;
        RECT 250.600 95.200 251.600 96.000 ;
        RECT 250.600 90.800 251.400 95.200 ;
        RECT 252.400 94.600 253.200 99.800 ;
        RECT 258.800 96.600 259.600 99.800 ;
        RECT 260.400 97.000 261.200 99.800 ;
        RECT 262.000 97.000 262.800 99.800 ;
        RECT 263.600 97.000 264.400 99.800 ;
        RECT 265.200 97.000 266.000 99.800 ;
        RECT 268.400 97.000 269.200 99.800 ;
        RECT 271.600 97.000 272.400 99.800 ;
        RECT 273.200 97.000 274.000 99.800 ;
        RECT 274.800 97.000 275.600 99.800 ;
        RECT 257.200 95.800 259.600 96.600 ;
        RECT 276.400 96.600 277.200 99.800 ;
        RECT 257.200 95.200 258.000 95.800 ;
        RECT 252.000 94.000 253.200 94.600 ;
        RECT 256.200 94.600 258.000 95.200 ;
        RECT 262.000 95.600 263.000 96.400 ;
        RECT 266.000 95.600 267.600 96.400 ;
        RECT 268.400 95.800 273.000 96.400 ;
        RECT 276.400 95.800 279.000 96.600 ;
        RECT 268.400 95.600 269.200 95.800 ;
        RECT 252.000 92.000 252.600 94.000 ;
        RECT 256.200 93.400 257.000 94.600 ;
        RECT 253.200 92.600 257.000 93.400 ;
        RECT 262.000 92.800 262.800 95.600 ;
        RECT 268.400 94.800 269.200 95.000 ;
        RECT 264.800 94.200 269.200 94.800 ;
        RECT 264.800 94.000 265.600 94.200 ;
        RECT 270.000 93.600 270.800 95.200 ;
        RECT 272.200 93.400 273.000 95.800 ;
        RECT 278.200 95.200 279.000 95.800 ;
        RECT 278.200 94.400 281.200 95.200 ;
        RECT 282.800 93.800 283.600 99.800 ;
        RECT 265.200 92.600 268.400 93.400 ;
        RECT 272.200 92.600 274.200 93.400 ;
        RECT 274.800 93.000 283.600 93.800 ;
        RECT 258.800 92.000 259.600 92.600 ;
        RECT 276.400 92.000 277.200 92.400 ;
        RECT 279.600 92.000 280.400 92.400 ;
        RECT 281.400 92.000 282.200 92.200 ;
        RECT 252.000 91.400 252.800 92.000 ;
        RECT 258.800 91.400 282.200 92.000 ;
        RECT 250.600 90.000 251.600 90.800 ;
        RECT 250.800 82.200 251.600 90.000 ;
        RECT 252.200 89.600 252.800 91.400 ;
        RECT 252.200 89.000 261.200 89.600 ;
        RECT 252.200 87.400 252.800 89.000 ;
        RECT 260.400 88.800 261.200 89.000 ;
        RECT 263.600 89.000 272.200 89.600 ;
        RECT 263.600 88.800 264.400 89.000 ;
        RECT 255.400 87.600 258.000 88.400 ;
        RECT 252.200 86.800 254.800 87.400 ;
        RECT 254.000 82.200 254.800 86.800 ;
        RECT 257.200 82.200 258.000 87.600 ;
        RECT 258.600 86.800 262.800 87.600 ;
        RECT 260.400 82.200 261.200 85.000 ;
        RECT 262.000 82.200 262.800 85.000 ;
        RECT 263.600 82.200 264.400 85.000 ;
        RECT 265.200 82.200 266.000 88.400 ;
        RECT 268.400 87.600 271.000 88.400 ;
        RECT 271.600 88.200 272.200 89.000 ;
        RECT 273.200 89.400 274.000 89.600 ;
        RECT 273.200 89.000 278.600 89.400 ;
        RECT 273.200 88.800 279.400 89.000 ;
        RECT 278.000 88.200 279.400 88.800 ;
        RECT 271.600 87.600 277.400 88.200 ;
        RECT 280.400 88.000 282.000 88.800 ;
        RECT 280.400 87.600 281.000 88.000 ;
        RECT 268.400 82.200 269.200 87.000 ;
        RECT 271.600 82.200 272.400 87.000 ;
        RECT 276.800 86.800 281.000 87.600 ;
        RECT 282.800 87.400 283.600 93.000 ;
        RECT 281.600 86.800 283.600 87.400 ;
        RECT 284.400 93.800 285.200 99.800 ;
        RECT 290.800 96.600 291.600 99.800 ;
        RECT 292.400 97.000 293.200 99.800 ;
        RECT 294.000 97.000 294.800 99.800 ;
        RECT 295.600 97.000 296.400 99.800 ;
        RECT 298.800 97.000 299.600 99.800 ;
        RECT 302.000 97.000 302.800 99.800 ;
        RECT 303.600 97.000 304.400 99.800 ;
        RECT 305.200 97.000 306.000 99.800 ;
        RECT 306.800 97.000 307.600 99.800 ;
        RECT 289.000 95.800 291.600 96.600 ;
        RECT 308.400 96.600 309.200 99.800 ;
        RECT 295.000 95.800 299.600 96.400 ;
        RECT 289.000 95.200 289.800 95.800 ;
        RECT 286.800 94.400 289.800 95.200 ;
        RECT 284.400 93.000 293.200 93.800 ;
        RECT 295.000 93.400 295.800 95.800 ;
        RECT 298.800 95.600 299.600 95.800 ;
        RECT 300.400 95.600 302.000 96.400 ;
        RECT 305.000 95.600 306.000 96.400 ;
        RECT 308.400 95.800 310.800 96.600 ;
        RECT 297.200 93.600 298.000 95.200 ;
        RECT 298.800 94.800 299.600 95.000 ;
        RECT 298.800 94.200 303.200 94.800 ;
        RECT 302.400 94.000 303.200 94.200 ;
        RECT 284.400 87.400 285.200 93.000 ;
        RECT 293.800 92.600 295.800 93.400 ;
        RECT 299.600 92.600 302.800 93.400 ;
        RECT 305.200 92.800 306.000 95.600 ;
        RECT 310.000 95.200 310.800 95.800 ;
        RECT 310.000 94.600 311.800 95.200 ;
        RECT 311.000 93.400 311.800 94.600 ;
        RECT 314.800 94.600 315.600 99.800 ;
        RECT 316.400 96.000 317.200 99.800 ;
        RECT 326.000 96.400 326.800 99.800 ;
        RECT 316.400 95.200 317.400 96.000 ;
        RECT 314.800 94.000 316.000 94.600 ;
        RECT 311.000 92.600 314.800 93.400 ;
        RECT 286.000 92.200 286.800 92.400 ;
        RECT 285.800 92.000 286.800 92.200 ;
        RECT 287.600 92.000 288.400 92.400 ;
        RECT 290.800 92.000 291.600 92.400 ;
        RECT 308.400 92.000 309.200 92.600 ;
        RECT 315.400 92.000 316.000 94.000 ;
        RECT 285.800 91.400 309.200 92.000 ;
        RECT 315.200 91.400 316.000 92.000 ;
        RECT 315.200 89.600 315.800 91.400 ;
        RECT 316.600 90.800 317.400 95.200 ;
        RECT 294.000 89.400 294.800 89.600 ;
        RECT 289.400 89.000 294.800 89.400 ;
        RECT 288.600 88.800 294.800 89.000 ;
        RECT 295.800 89.000 304.400 89.600 ;
        RECT 286.000 88.000 287.600 88.800 ;
        RECT 288.600 88.200 290.000 88.800 ;
        RECT 295.800 88.200 296.400 89.000 ;
        RECT 303.600 88.800 304.400 89.000 ;
        RECT 306.800 89.000 315.800 89.600 ;
        RECT 306.800 88.800 307.600 89.000 ;
        RECT 287.000 87.600 287.600 88.000 ;
        RECT 290.600 87.600 296.400 88.200 ;
        RECT 297.000 87.600 299.600 88.400 ;
        RECT 284.400 86.800 286.400 87.400 ;
        RECT 287.000 86.800 291.200 87.600 ;
        RECT 273.200 82.200 274.000 85.000 ;
        RECT 274.800 82.200 275.600 85.000 ;
        RECT 278.000 82.200 278.800 86.800 ;
        RECT 281.600 86.200 282.200 86.800 ;
        RECT 281.200 85.600 282.200 86.200 ;
        RECT 285.800 86.200 286.400 86.800 ;
        RECT 285.800 85.600 286.800 86.200 ;
        RECT 281.200 82.200 282.000 85.600 ;
        RECT 286.000 82.200 286.800 85.600 ;
        RECT 289.200 82.200 290.000 86.800 ;
        RECT 292.400 82.200 293.200 85.000 ;
        RECT 294.000 82.200 294.800 85.000 ;
        RECT 295.600 82.200 296.400 87.000 ;
        RECT 298.800 82.200 299.600 87.000 ;
        RECT 302.000 82.200 302.800 88.400 ;
        RECT 310.000 87.600 312.600 88.400 ;
        RECT 305.200 86.800 309.400 87.600 ;
        RECT 303.600 82.200 304.400 85.000 ;
        RECT 305.200 82.200 306.000 85.000 ;
        RECT 306.800 82.200 307.600 85.000 ;
        RECT 310.000 82.200 310.800 87.600 ;
        RECT 315.200 87.400 315.800 89.000 ;
        RECT 313.200 86.800 315.800 87.400 ;
        RECT 316.400 90.000 317.400 90.800 ;
        RECT 325.800 95.800 326.800 96.400 ;
        RECT 325.800 94.400 326.400 95.800 ;
        RECT 329.200 95.200 330.000 99.800 ;
        RECT 332.400 96.000 333.200 99.800 ;
        RECT 327.400 94.600 330.000 95.200 ;
        RECT 332.200 95.200 333.200 96.000 ;
        RECT 325.800 93.600 326.800 94.400 ;
        RECT 325.800 90.200 326.400 93.600 ;
        RECT 327.400 93.000 328.000 94.600 ;
        RECT 327.000 92.200 328.000 93.000 ;
        RECT 327.400 90.200 328.000 92.200 ;
        RECT 329.000 92.400 329.800 93.200 ;
        RECT 329.000 92.300 330.000 92.400 ;
        RECT 332.200 92.300 333.000 95.200 ;
        RECT 334.000 94.600 334.800 99.800 ;
        RECT 340.400 96.600 341.200 99.800 ;
        RECT 342.000 97.000 342.800 99.800 ;
        RECT 343.600 97.000 344.400 99.800 ;
        RECT 345.200 97.000 346.000 99.800 ;
        RECT 346.800 97.000 347.600 99.800 ;
        RECT 350.000 97.000 350.800 99.800 ;
        RECT 353.200 97.000 354.000 99.800 ;
        RECT 354.800 97.000 355.600 99.800 ;
        RECT 356.400 97.000 357.200 99.800 ;
        RECT 338.800 95.800 341.200 96.600 ;
        RECT 358.000 96.600 358.800 99.800 ;
        RECT 338.800 95.200 339.600 95.800 ;
        RECT 329.000 91.700 333.000 92.300 ;
        RECT 329.000 91.600 330.000 91.700 ;
        RECT 332.200 90.800 333.000 91.700 ;
        RECT 333.600 94.000 334.800 94.600 ;
        RECT 337.800 94.600 339.600 95.200 ;
        RECT 343.600 95.600 344.600 96.400 ;
        RECT 347.600 95.600 349.200 96.400 ;
        RECT 350.000 95.800 354.600 96.400 ;
        RECT 358.000 95.800 360.600 96.600 ;
        RECT 350.000 95.600 350.800 95.800 ;
        RECT 333.600 92.000 334.200 94.000 ;
        RECT 337.800 93.400 338.600 94.600 ;
        RECT 334.800 92.600 338.600 93.400 ;
        RECT 343.600 92.800 344.400 95.600 ;
        RECT 350.000 94.800 350.800 95.000 ;
        RECT 346.400 94.200 350.800 94.800 ;
        RECT 346.400 94.000 347.200 94.200 ;
        RECT 351.600 93.600 352.400 95.200 ;
        RECT 353.800 93.400 354.600 95.800 ;
        RECT 359.800 95.200 360.600 95.800 ;
        RECT 359.800 94.400 362.800 95.200 ;
        RECT 364.400 93.800 365.200 99.800 ;
        RECT 346.800 92.600 350.000 93.400 ;
        RECT 353.800 92.600 355.800 93.400 ;
        RECT 356.400 93.000 365.200 93.800 ;
        RECT 333.600 91.400 334.400 92.000 ;
        RECT 313.200 82.200 314.000 86.800 ;
        RECT 316.400 82.200 317.200 90.000 ;
        RECT 325.800 89.200 326.800 90.200 ;
        RECT 327.400 89.600 330.000 90.200 ;
        RECT 332.200 90.000 333.200 90.800 ;
        RECT 326.000 82.200 326.800 89.200 ;
        RECT 329.200 82.200 330.000 89.600 ;
        RECT 332.400 82.200 333.200 90.000 ;
        RECT 333.800 89.600 334.400 91.400 ;
        RECT 335.000 90.800 335.800 91.000 ;
        RECT 335.000 90.200 362.000 90.800 ;
        RECT 357.800 90.000 358.800 90.200 ;
        RECT 361.200 89.600 362.000 90.200 ;
        RECT 333.800 89.000 342.800 89.600 ;
        RECT 333.800 87.400 334.400 89.000 ;
        RECT 342.000 88.800 342.800 89.000 ;
        RECT 345.200 89.000 353.800 89.600 ;
        RECT 345.200 88.800 346.000 89.000 ;
        RECT 337.000 87.600 339.600 88.400 ;
        RECT 333.800 86.800 336.400 87.400 ;
        RECT 335.600 82.200 336.400 86.800 ;
        RECT 338.800 82.200 339.600 87.600 ;
        RECT 340.200 86.800 344.400 87.600 ;
        RECT 342.000 82.200 342.800 85.000 ;
        RECT 343.600 82.200 344.400 85.000 ;
        RECT 345.200 82.200 346.000 85.000 ;
        RECT 346.800 82.200 347.600 88.400 ;
        RECT 350.000 87.600 352.600 88.400 ;
        RECT 353.200 88.200 353.800 89.000 ;
        RECT 354.800 89.400 355.600 89.600 ;
        RECT 354.800 89.000 360.200 89.400 ;
        RECT 354.800 88.800 361.000 89.000 ;
        RECT 359.600 88.200 361.000 88.800 ;
        RECT 353.200 87.600 359.000 88.200 ;
        RECT 362.000 88.000 363.600 88.800 ;
        RECT 362.000 87.600 362.600 88.000 ;
        RECT 350.000 82.200 350.800 87.000 ;
        RECT 353.200 82.200 354.000 87.000 ;
        RECT 358.400 86.800 362.600 87.600 ;
        RECT 364.400 87.400 365.200 93.000 ;
        RECT 363.200 86.800 365.200 87.400 ;
        RECT 366.000 93.800 366.800 99.800 ;
        RECT 372.400 96.600 373.200 99.800 ;
        RECT 374.000 97.000 374.800 99.800 ;
        RECT 375.600 97.000 376.400 99.800 ;
        RECT 377.200 97.000 378.000 99.800 ;
        RECT 380.400 97.000 381.200 99.800 ;
        RECT 383.600 97.000 384.400 99.800 ;
        RECT 385.200 97.000 386.000 99.800 ;
        RECT 386.800 97.000 387.600 99.800 ;
        RECT 388.400 97.000 389.200 99.800 ;
        RECT 370.600 95.800 373.200 96.600 ;
        RECT 390.000 96.600 390.800 99.800 ;
        RECT 376.600 95.800 381.200 96.400 ;
        RECT 370.600 95.200 371.400 95.800 ;
        RECT 368.400 94.400 371.400 95.200 ;
        RECT 366.000 93.000 374.800 93.800 ;
        RECT 376.600 93.400 377.400 95.800 ;
        RECT 380.400 95.600 381.200 95.800 ;
        RECT 382.000 95.600 383.600 96.400 ;
        RECT 386.600 95.600 387.600 96.400 ;
        RECT 390.000 95.800 392.400 96.600 ;
        RECT 378.800 93.600 379.600 95.200 ;
        RECT 380.400 94.800 381.200 95.000 ;
        RECT 380.400 94.200 384.800 94.800 ;
        RECT 384.000 94.000 384.800 94.200 ;
        RECT 366.000 87.400 366.800 93.000 ;
        RECT 375.400 92.600 377.400 93.400 ;
        RECT 381.200 92.600 384.400 93.400 ;
        RECT 386.800 92.800 387.600 95.600 ;
        RECT 391.600 95.200 392.400 95.800 ;
        RECT 391.600 94.600 393.400 95.200 ;
        RECT 392.600 93.400 393.400 94.600 ;
        RECT 396.400 94.600 397.200 99.800 ;
        RECT 398.000 96.000 398.800 99.800 ;
        RECT 398.000 95.200 399.000 96.000 ;
        RECT 401.200 95.800 402.000 99.800 ;
        RECT 402.800 96.000 403.600 99.800 ;
        RECT 406.000 96.000 406.800 99.800 ;
        RECT 402.800 95.800 406.800 96.000 ;
        RECT 396.400 94.000 397.600 94.600 ;
        RECT 392.600 92.600 396.400 93.400 ;
        RECT 367.400 92.000 368.200 92.200 ;
        RECT 369.200 92.000 370.000 92.400 ;
        RECT 372.400 92.000 373.200 92.400 ;
        RECT 390.000 92.000 390.800 92.600 ;
        RECT 397.000 92.000 397.600 94.000 ;
        RECT 367.400 91.400 390.800 92.000 ;
        RECT 396.800 91.400 397.600 92.000 ;
        RECT 396.800 89.600 397.400 91.400 ;
        RECT 398.200 90.800 399.000 95.200 ;
        RECT 401.400 94.400 402.000 95.800 ;
        RECT 403.000 95.400 406.600 95.800 ;
        RECT 407.600 95.600 408.400 97.200 ;
        RECT 405.200 94.400 406.000 94.800 ;
        RECT 401.200 93.600 403.800 94.400 ;
        RECT 405.200 94.300 406.800 94.400 ;
        RECT 407.600 94.300 408.400 94.400 ;
        RECT 405.200 93.800 408.400 94.300 ;
        RECT 406.000 93.700 408.400 93.800 ;
        RECT 406.000 93.600 406.800 93.700 ;
        RECT 407.600 93.600 408.400 93.700 ;
        RECT 409.200 94.300 410.000 99.800 ;
        RECT 410.800 96.000 411.600 99.800 ;
        RECT 414.000 96.000 414.800 99.800 ;
        RECT 410.800 95.800 414.800 96.000 ;
        RECT 415.600 95.800 416.400 99.800 ;
        RECT 421.000 98.400 421.800 99.000 ;
        RECT 421.000 97.600 422.800 98.400 ;
        RECT 421.000 96.000 421.800 97.600 ;
        RECT 425.200 97.000 426.000 99.000 ;
        RECT 411.000 95.400 414.600 95.800 ;
        RECT 411.600 94.400 412.400 94.800 ;
        RECT 415.600 94.400 416.200 95.800 ;
        RECT 420.200 95.400 421.800 96.000 ;
        RECT 420.200 95.000 421.000 95.400 ;
        RECT 420.200 94.400 420.800 95.000 ;
        RECT 425.400 94.800 426.000 97.000 ;
        RECT 410.800 94.300 412.400 94.400 ;
        RECT 409.200 93.800 412.400 94.300 ;
        RECT 409.200 93.700 411.600 93.800 ;
        RECT 375.600 89.400 376.400 89.600 ;
        RECT 371.000 89.000 376.400 89.400 ;
        RECT 370.200 88.800 376.400 89.000 ;
        RECT 377.400 89.000 386.000 89.600 ;
        RECT 367.600 88.000 369.200 88.800 ;
        RECT 370.200 88.200 371.600 88.800 ;
        RECT 377.400 88.200 378.000 89.000 ;
        RECT 385.200 88.800 386.000 89.000 ;
        RECT 388.400 89.000 397.400 89.600 ;
        RECT 388.400 88.800 389.200 89.000 ;
        RECT 368.600 87.600 369.200 88.000 ;
        RECT 372.200 87.600 378.000 88.200 ;
        RECT 378.600 87.600 381.200 88.400 ;
        RECT 366.000 86.800 368.000 87.400 ;
        RECT 368.600 86.800 372.800 87.600 ;
        RECT 354.800 82.200 355.600 85.000 ;
        RECT 356.400 82.200 357.200 85.000 ;
        RECT 359.600 82.200 360.400 86.800 ;
        RECT 363.200 86.200 363.800 86.800 ;
        RECT 362.800 85.600 363.800 86.200 ;
        RECT 367.400 86.200 368.000 86.800 ;
        RECT 367.400 85.600 368.400 86.200 ;
        RECT 362.800 82.200 363.600 85.600 ;
        RECT 367.600 82.200 368.400 85.600 ;
        RECT 370.800 82.200 371.600 86.800 ;
        RECT 374.000 82.200 374.800 85.000 ;
        RECT 375.600 82.200 376.400 85.000 ;
        RECT 377.200 82.200 378.000 87.000 ;
        RECT 380.400 82.200 381.200 87.000 ;
        RECT 383.600 82.200 384.400 88.400 ;
        RECT 391.600 87.600 394.200 88.400 ;
        RECT 386.800 86.800 391.000 87.600 ;
        RECT 385.200 82.200 386.000 85.000 ;
        RECT 386.800 82.200 387.600 85.000 ;
        RECT 388.400 82.200 389.200 85.000 ;
        RECT 391.600 82.200 392.400 87.600 ;
        RECT 396.800 87.400 397.400 89.000 ;
        RECT 394.800 86.800 397.400 87.400 ;
        RECT 398.000 90.000 399.000 90.800 ;
        RECT 401.200 90.200 402.000 90.400 ;
        RECT 403.200 90.200 403.800 93.600 ;
        RECT 404.400 91.600 405.200 93.200 ;
        RECT 394.800 82.200 395.600 86.800 ;
        RECT 398.000 82.200 398.800 90.000 ;
        RECT 401.200 89.600 402.600 90.200 ;
        RECT 403.200 89.600 404.200 90.200 ;
        RECT 402.000 88.400 402.600 89.600 ;
        RECT 402.000 87.600 402.800 88.400 ;
        RECT 403.400 82.200 404.200 89.600 ;
        RECT 409.200 82.200 410.000 93.700 ;
        RECT 410.800 93.600 411.600 93.700 ;
        RECT 413.800 93.600 416.400 94.400 ;
        RECT 418.800 93.600 420.800 94.400 ;
        RECT 421.800 94.200 426.000 94.800 ;
        RECT 428.400 97.600 429.200 99.800 ;
        RECT 428.400 94.400 429.000 97.600 ;
        RECT 430.000 95.600 430.800 97.200 ;
        RECT 433.200 96.400 434.000 99.800 ;
        RECT 433.000 95.800 434.000 96.400 ;
        RECT 433.000 94.400 433.600 95.800 ;
        RECT 436.400 95.200 437.200 99.800 ;
        RECT 438.000 96.000 438.800 99.800 ;
        RECT 441.200 96.000 442.000 99.800 ;
        RECT 438.000 95.800 442.000 96.000 ;
        RECT 442.800 95.800 443.600 99.800 ;
        RECT 446.000 97.800 446.800 99.800 ;
        RECT 438.200 95.400 441.800 95.800 ;
        RECT 434.600 94.600 437.200 95.200 ;
        RECT 421.800 93.800 422.800 94.200 ;
        RECT 412.400 91.600 413.200 93.200 ;
        RECT 413.800 90.200 414.400 93.600 ;
        RECT 418.800 90.800 419.600 92.400 ;
        RECT 415.600 90.200 416.400 90.400 ;
        RECT 413.400 89.600 414.400 90.200 ;
        RECT 415.000 89.600 416.400 90.200 ;
        RECT 420.200 89.800 420.800 93.600 ;
        RECT 421.400 93.000 422.800 93.800 ;
        RECT 428.400 93.600 429.200 94.400 ;
        RECT 433.000 93.600 434.000 94.400 ;
        RECT 422.200 91.000 422.800 93.000 ;
        RECT 423.600 91.600 424.400 93.200 ;
        RECT 425.200 91.600 426.000 93.200 ;
        RECT 422.200 90.400 426.000 91.000 ;
        RECT 426.800 90.800 427.600 92.400 ;
        RECT 413.400 82.200 414.200 89.600 ;
        RECT 415.000 88.400 415.600 89.600 ;
        RECT 420.200 89.200 421.800 89.800 ;
        RECT 414.800 87.600 415.600 88.400 ;
        RECT 421.000 82.200 421.800 89.200 ;
        RECT 425.400 87.000 426.000 90.400 ;
        RECT 428.400 90.200 429.000 93.600 ;
        RECT 433.000 90.200 433.600 93.600 ;
        RECT 434.600 93.000 435.200 94.600 ;
        RECT 438.800 94.400 439.600 94.800 ;
        RECT 442.800 94.400 443.400 95.800 ;
        RECT 446.000 94.400 446.600 97.800 ;
        RECT 447.600 95.600 448.400 97.200 ;
        RECT 449.200 95.800 450.000 99.800 ;
        RECT 450.800 96.000 451.600 99.800 ;
        RECT 454.000 96.000 454.800 99.800 ;
        RECT 450.800 95.800 454.800 96.000 ;
        RECT 456.200 96.400 457.000 99.800 ;
        RECT 465.200 97.000 466.000 99.000 ;
        RECT 456.200 95.800 458.000 96.400 ;
        RECT 449.400 94.400 450.000 95.800 ;
        RECT 451.000 95.400 454.600 95.800 ;
        RECT 453.200 94.400 454.000 94.800 ;
        RECT 438.000 93.800 439.600 94.400 ;
        RECT 438.000 93.600 438.800 93.800 ;
        RECT 441.000 93.600 443.600 94.400 ;
        RECT 446.000 93.600 446.800 94.400 ;
        RECT 449.200 93.600 451.800 94.400 ;
        RECT 453.200 94.300 454.800 94.400 ;
        RECT 455.600 94.300 456.400 94.400 ;
        RECT 453.200 93.800 456.400 94.300 ;
        RECT 454.000 93.700 456.400 93.800 ;
        RECT 454.000 93.600 454.800 93.700 ;
        RECT 455.600 93.600 456.400 93.700 ;
        RECT 434.200 92.200 435.200 93.000 ;
        RECT 434.600 90.200 435.200 92.200 ;
        RECT 436.200 92.400 437.000 93.200 ;
        RECT 436.200 91.600 437.200 92.400 ;
        RECT 439.600 91.600 440.400 93.200 ;
        RECT 441.000 90.200 441.600 93.600 ;
        RECT 444.400 90.800 445.200 92.400 ;
        RECT 446.000 92.300 446.600 93.600 ;
        RECT 449.200 92.300 450.000 92.400 ;
        RECT 446.000 91.700 450.000 92.300 ;
        RECT 442.800 90.200 443.600 90.400 ;
        RECT 446.000 90.200 446.600 91.700 ;
        RECT 449.200 91.600 450.000 91.700 ;
        RECT 449.200 90.200 450.000 90.400 ;
        RECT 451.200 90.200 451.800 93.600 ;
        RECT 452.400 91.600 453.200 93.200 ;
        RECT 425.200 83.000 426.000 87.000 ;
        RECT 427.400 89.400 429.200 90.200 ;
        RECT 427.400 82.200 428.200 89.400 ;
        RECT 433.000 89.200 434.000 90.200 ;
        RECT 434.600 89.600 437.200 90.200 ;
        RECT 433.200 82.200 434.000 89.200 ;
        RECT 436.400 82.200 437.200 89.600 ;
        RECT 440.600 89.600 441.600 90.200 ;
        RECT 442.200 89.600 443.600 90.200 ;
        RECT 440.600 84.400 441.400 89.600 ;
        RECT 442.200 88.400 442.800 89.600 ;
        RECT 442.000 87.600 442.800 88.400 ;
        RECT 445.000 89.400 446.800 90.200 ;
        RECT 449.200 89.600 450.600 90.200 ;
        RECT 451.200 89.600 452.200 90.200 ;
        RECT 439.600 83.600 441.400 84.400 ;
        RECT 440.600 82.200 441.400 83.600 ;
        RECT 445.000 82.200 445.800 89.400 ;
        RECT 450.000 88.400 450.600 89.600 ;
        RECT 450.000 87.600 450.800 88.400 ;
        RECT 451.400 82.200 452.200 89.600 ;
        RECT 455.600 88.800 456.400 90.400 ;
        RECT 457.200 82.200 458.000 95.800 ;
        RECT 458.800 93.600 459.600 95.200 ;
        RECT 465.200 94.800 465.800 97.000 ;
        RECT 469.400 96.000 470.200 99.000 ;
        RECT 469.400 95.400 471.000 96.000 ;
        RECT 470.200 95.000 471.000 95.400 ;
        RECT 465.200 94.200 469.400 94.800 ;
        RECT 468.400 93.800 469.400 94.200 ;
        RECT 470.400 94.400 471.000 95.000 ;
        RECT 465.200 91.600 466.000 93.200 ;
        RECT 466.800 91.600 467.600 93.200 ;
        RECT 468.400 93.000 469.800 93.800 ;
        RECT 470.400 93.600 472.400 94.400 ;
        RECT 473.200 94.300 474.000 94.400 ;
        RECT 474.800 94.300 475.600 99.800 ;
        RECT 476.400 95.600 477.200 97.200 ;
        RECT 479.600 96.400 480.400 99.800 ;
        RECT 479.400 95.800 480.400 96.400 ;
        RECT 473.200 93.700 475.600 94.300 ;
        RECT 473.200 93.600 474.000 93.700 ;
        RECT 468.400 91.000 469.000 93.000 ;
        RECT 465.200 90.400 469.000 91.000 ;
        RECT 465.200 87.000 465.800 90.400 ;
        RECT 470.400 89.800 471.000 93.600 ;
        RECT 471.600 90.800 472.400 92.400 ;
        RECT 469.400 89.200 471.000 89.800 ;
        RECT 465.200 83.000 466.000 87.000 ;
        RECT 469.400 84.400 470.200 89.200 ;
        RECT 469.400 83.600 470.800 84.400 ;
        RECT 469.400 82.200 470.200 83.600 ;
        RECT 474.800 82.200 475.600 93.700 ;
        RECT 479.400 94.400 480.000 95.800 ;
        RECT 482.800 95.200 483.600 99.800 ;
        RECT 481.000 94.600 483.600 95.200 ;
        RECT 484.400 95.200 485.200 99.800 ;
        RECT 487.600 96.400 488.400 99.800 ;
        RECT 487.600 95.800 488.600 96.400 ;
        RECT 490.800 96.000 491.600 99.800 ;
        RECT 494.000 96.000 494.800 99.800 ;
        RECT 490.800 95.800 494.800 96.000 ;
        RECT 495.600 95.800 496.400 99.800 ;
        RECT 497.200 97.000 498.000 99.000 ;
        RECT 484.400 94.600 487.000 95.200 ;
        RECT 479.400 93.600 480.400 94.400 ;
        RECT 479.400 90.200 480.000 93.600 ;
        RECT 481.000 93.000 481.600 94.600 ;
        RECT 480.600 92.200 481.600 93.000 ;
        RECT 481.000 90.200 481.600 92.200 ;
        RECT 482.600 92.400 483.400 93.200 ;
        RECT 484.600 92.400 485.400 93.200 ;
        RECT 482.600 92.300 483.600 92.400 ;
        RECT 484.400 92.300 485.400 92.400 ;
        RECT 482.600 91.700 485.400 92.300 ;
        RECT 482.600 91.600 483.600 91.700 ;
        RECT 484.400 91.600 485.400 91.700 ;
        RECT 486.400 93.000 487.000 94.600 ;
        RECT 488.000 94.400 488.600 95.800 ;
        RECT 491.000 95.400 494.600 95.800 ;
        RECT 491.600 94.400 492.400 94.800 ;
        RECT 495.600 94.400 496.200 95.800 ;
        RECT 497.200 94.800 497.800 97.000 ;
        RECT 501.400 96.000 502.200 99.000 ;
        RECT 501.400 95.400 503.000 96.000 ;
        RECT 502.200 95.000 503.000 95.400 ;
        RECT 487.600 93.600 488.600 94.400 ;
        RECT 490.800 93.800 492.400 94.400 ;
        RECT 490.800 93.600 491.600 93.800 ;
        RECT 493.800 93.600 496.400 94.400 ;
        RECT 497.200 94.200 501.400 94.800 ;
        RECT 500.400 93.800 501.400 94.200 ;
        RECT 502.400 94.400 503.000 95.000 ;
        RECT 506.800 95.200 507.600 99.800 ;
        RECT 510.000 96.400 510.800 99.800 ;
        RECT 515.800 98.400 516.600 99.800 ;
        RECT 515.800 97.600 517.200 98.400 ;
        RECT 515.800 96.400 516.600 97.600 ;
        RECT 510.000 95.600 511.000 96.400 ;
        RECT 506.800 94.600 509.400 95.200 ;
        RECT 486.400 92.200 487.400 93.000 ;
        RECT 486.400 90.200 487.000 92.200 ;
        RECT 488.000 90.200 488.600 93.600 ;
        RECT 490.800 92.300 491.600 92.400 ;
        RECT 492.400 92.300 493.200 93.200 ;
        RECT 490.800 91.700 493.200 92.300 ;
        RECT 490.800 91.600 491.600 91.700 ;
        RECT 492.400 91.600 493.200 91.700 ;
        RECT 493.800 90.200 494.400 93.600 ;
        RECT 497.200 91.600 498.000 93.200 ;
        RECT 498.800 91.600 499.600 93.200 ;
        RECT 500.400 93.000 501.800 93.800 ;
        RECT 502.400 93.600 504.400 94.400 ;
        RECT 500.400 91.000 501.000 93.000 ;
        RECT 497.200 90.400 501.000 91.000 ;
        RECT 495.600 90.200 496.400 90.400 ;
        RECT 479.400 89.200 480.400 90.200 ;
        RECT 481.000 89.600 483.600 90.200 ;
        RECT 479.600 82.200 480.400 89.200 ;
        RECT 482.800 82.200 483.600 89.600 ;
        RECT 484.400 89.600 487.000 90.200 ;
        RECT 484.400 82.200 485.200 89.600 ;
        RECT 487.600 89.200 488.600 90.200 ;
        RECT 493.400 89.600 494.400 90.200 ;
        RECT 495.000 89.600 496.400 90.200 ;
        RECT 487.600 82.200 488.400 89.200 ;
        RECT 493.400 84.400 494.200 89.600 ;
        RECT 495.000 88.400 495.600 89.600 ;
        RECT 494.800 87.600 495.600 88.400 ;
        RECT 492.400 83.600 494.200 84.400 ;
        RECT 493.400 82.200 494.200 83.600 ;
        RECT 497.200 87.000 497.800 90.400 ;
        RECT 502.400 89.800 503.000 93.600 ;
        RECT 507.000 92.400 507.800 93.200 ;
        RECT 503.600 90.800 504.400 92.400 ;
        RECT 506.800 91.600 507.800 92.400 ;
        RECT 508.800 93.000 509.400 94.600 ;
        RECT 510.400 94.400 511.000 95.600 ;
        RECT 514.800 95.800 516.600 96.400 ;
        RECT 518.000 97.000 518.800 99.000 ;
        RECT 510.000 93.600 511.000 94.400 ;
        RECT 511.600 94.300 512.400 94.400 ;
        RECT 513.200 94.300 514.000 95.200 ;
        RECT 511.600 93.700 514.000 94.300 ;
        RECT 511.600 93.600 512.400 93.700 ;
        RECT 513.200 93.600 514.000 93.700 ;
        RECT 508.800 92.200 509.800 93.000 ;
        RECT 508.800 90.200 509.400 92.200 ;
        RECT 510.400 90.200 511.000 93.600 ;
        RECT 501.400 89.200 503.000 89.800 ;
        RECT 506.800 89.600 509.400 90.200 ;
        RECT 497.200 83.000 498.000 87.000 ;
        RECT 501.400 84.400 502.200 89.200 ;
        RECT 501.400 83.600 502.800 84.400 ;
        RECT 501.400 82.200 502.200 83.600 ;
        RECT 506.800 82.200 507.600 89.600 ;
        RECT 510.000 89.200 511.000 90.200 ;
        RECT 510.000 82.200 510.800 89.200 ;
        RECT 514.800 82.200 515.600 95.800 ;
        RECT 518.000 94.800 518.600 97.000 ;
        RECT 522.200 96.000 523.000 99.000 ;
        RECT 527.600 96.000 528.400 99.800 ;
        RECT 530.800 96.000 531.600 99.800 ;
        RECT 522.200 95.400 523.800 96.000 ;
        RECT 527.600 95.800 531.600 96.000 ;
        RECT 532.400 95.800 533.200 99.800 ;
        RECT 534.000 95.800 534.800 99.800 ;
        RECT 535.600 96.000 536.400 99.800 ;
        RECT 538.800 96.000 539.600 99.800 ;
        RECT 543.000 98.400 543.800 99.800 ;
        RECT 542.000 97.600 543.800 98.400 ;
        RECT 543.000 96.400 543.800 97.600 ;
        RECT 535.600 95.800 539.600 96.000 ;
        RECT 542.000 95.800 543.800 96.400 ;
        RECT 527.800 95.400 531.400 95.800 ;
        RECT 523.000 95.000 523.800 95.400 ;
        RECT 518.000 94.200 522.200 94.800 ;
        RECT 521.200 93.800 522.200 94.200 ;
        RECT 523.200 94.400 523.800 95.000 ;
        RECT 528.400 94.400 529.200 94.800 ;
        RECT 532.400 94.400 533.000 95.800 ;
        RECT 534.200 94.400 534.800 95.800 ;
        RECT 535.800 95.400 539.400 95.800 ;
        RECT 538.000 94.400 538.800 94.800 ;
        RECT 523.200 94.300 525.200 94.400 ;
        RECT 518.000 91.600 518.800 93.200 ;
        RECT 519.600 91.600 520.400 93.200 ;
        RECT 521.200 93.000 522.600 93.800 ;
        RECT 523.200 93.700 526.700 94.300 ;
        RECT 523.200 93.600 525.200 93.700 ;
        RECT 521.200 91.000 521.800 93.000 ;
        RECT 518.000 90.400 521.800 91.000 ;
        RECT 516.400 87.600 517.200 90.400 ;
        RECT 518.000 87.000 518.600 90.400 ;
        RECT 523.200 89.800 523.800 93.600 ;
        RECT 524.400 90.800 525.200 92.400 ;
        RECT 526.100 92.300 526.700 93.700 ;
        RECT 527.600 93.800 529.200 94.400 ;
        RECT 527.600 93.600 528.400 93.800 ;
        RECT 530.600 93.600 533.200 94.400 ;
        RECT 534.000 93.600 536.600 94.400 ;
        RECT 538.000 93.800 539.600 94.400 ;
        RECT 538.800 93.600 539.600 93.800 ;
        RECT 540.400 93.600 541.200 95.200 ;
        RECT 529.200 92.300 530.000 93.200 ;
        RECT 526.100 91.700 530.000 92.300 ;
        RECT 529.200 91.600 530.000 91.700 ;
        RECT 530.600 90.200 531.200 93.600 ;
        RECT 536.000 92.300 536.600 93.600 ;
        RECT 532.500 91.700 536.600 92.300 ;
        RECT 532.500 90.400 533.100 91.700 ;
        RECT 532.400 90.200 533.200 90.400 ;
        RECT 522.200 89.200 523.800 89.800 ;
        RECT 530.200 89.600 531.200 90.200 ;
        RECT 531.800 89.600 533.200 90.200 ;
        RECT 534.000 90.200 534.800 90.400 ;
        RECT 536.000 90.200 536.600 91.700 ;
        RECT 537.200 91.600 538.000 93.200 ;
        RECT 534.000 89.600 535.400 90.200 ;
        RECT 536.000 89.600 537.000 90.200 ;
        RECT 518.000 83.000 518.800 87.000 ;
        RECT 522.200 82.200 523.000 89.200 ;
        RECT 530.200 82.200 531.000 89.600 ;
        RECT 531.800 88.400 532.400 89.600 ;
        RECT 531.600 87.600 532.400 88.400 ;
        RECT 534.800 88.400 535.400 89.600 ;
        RECT 534.800 87.600 535.600 88.400 ;
        RECT 536.200 82.200 537.000 89.600 ;
        RECT 542.000 82.200 542.800 95.800 ;
        RECT 545.200 95.400 546.000 99.800 ;
        RECT 549.400 98.400 550.600 99.800 ;
        RECT 549.400 97.800 550.800 98.400 ;
        RECT 554.000 97.800 554.800 99.800 ;
        RECT 558.400 98.400 559.200 99.800 ;
        RECT 558.400 97.800 560.400 98.400 ;
        RECT 550.000 97.000 550.800 97.800 ;
        RECT 554.200 97.200 554.800 97.800 ;
        RECT 554.200 96.600 557.000 97.200 ;
        RECT 556.200 96.400 557.000 96.600 ;
        RECT 558.000 96.400 558.800 97.200 ;
        RECT 559.600 97.000 560.400 97.800 ;
        RECT 548.200 95.400 549.000 95.600 ;
        RECT 545.200 94.800 549.000 95.400 ;
        RECT 545.200 91.400 546.000 94.800 ;
        RECT 552.200 94.200 553.000 94.400 ;
        RECT 558.000 94.200 558.600 96.400 ;
        RECT 562.800 95.000 563.600 99.800 ;
        RECT 567.000 98.400 567.800 99.800 ;
        RECT 566.000 97.600 567.800 98.400 ;
        RECT 567.000 96.400 567.800 97.600 ;
        RECT 566.000 95.800 567.800 96.400 ;
        RECT 569.200 96.000 570.000 99.800 ;
        RECT 572.400 96.000 573.200 99.800 ;
        RECT 569.200 95.800 573.200 96.000 ;
        RECT 574.000 95.800 574.800 99.800 ;
        RECT 561.200 94.200 562.800 94.400 ;
        RECT 551.800 93.600 562.800 94.200 ;
        RECT 564.400 93.600 565.200 95.200 ;
        RECT 550.000 92.800 550.800 93.000 ;
        RECT 547.000 92.200 550.800 92.800 ;
        RECT 547.000 92.000 547.800 92.200 ;
        RECT 548.600 91.400 549.400 91.600 ;
        RECT 545.200 90.800 549.400 91.400 ;
        RECT 543.600 87.600 544.400 90.400 ;
        RECT 545.200 82.200 546.000 90.800 ;
        RECT 551.800 90.400 552.400 93.600 ;
        RECT 559.000 93.400 559.800 93.600 ;
        RECT 560.600 92.400 561.400 92.600 ;
        RECT 556.400 91.800 561.400 92.400 ;
        RECT 556.400 91.600 557.200 91.800 ;
        RECT 558.000 91.000 563.600 91.200 ;
        RECT 557.800 90.800 563.600 91.000 ;
        RECT 550.000 89.800 552.400 90.400 ;
        RECT 553.800 90.600 563.600 90.800 ;
        RECT 553.800 90.200 558.600 90.600 ;
        RECT 550.000 88.800 550.600 89.800 ;
        RECT 549.200 88.000 550.600 88.800 ;
        RECT 552.200 89.000 553.000 89.200 ;
        RECT 553.800 89.000 554.400 90.200 ;
        RECT 552.200 88.400 554.400 89.000 ;
        RECT 555.000 89.000 560.400 89.600 ;
        RECT 555.000 88.800 555.800 89.000 ;
        RECT 559.600 88.800 560.400 89.000 ;
        RECT 553.400 87.400 554.200 87.600 ;
        RECT 556.200 87.400 557.000 87.600 ;
        RECT 550.000 86.200 550.800 87.000 ;
        RECT 553.400 86.800 557.000 87.400 ;
        RECT 554.200 86.200 554.800 86.800 ;
        RECT 559.600 86.200 560.400 87.000 ;
        RECT 549.400 82.200 550.600 86.200 ;
        RECT 554.000 82.200 554.800 86.200 ;
        RECT 558.400 85.600 560.400 86.200 ;
        RECT 558.400 82.200 559.200 85.600 ;
        RECT 562.800 82.200 563.600 90.600 ;
        RECT 566.000 82.200 566.800 95.800 ;
        RECT 569.400 95.400 573.000 95.800 ;
        RECT 570.000 94.400 570.800 94.800 ;
        RECT 574.000 94.400 574.600 95.800 ;
        RECT 569.200 93.800 570.800 94.400 ;
        RECT 569.200 93.600 570.000 93.800 ;
        RECT 572.200 93.600 574.800 94.400 ;
        RECT 575.600 93.800 576.400 99.800 ;
        RECT 582.000 96.600 582.800 99.800 ;
        RECT 583.600 97.000 584.400 99.800 ;
        RECT 585.200 97.000 586.000 99.800 ;
        RECT 586.800 97.000 587.600 99.800 ;
        RECT 590.000 97.000 590.800 99.800 ;
        RECT 593.200 97.000 594.000 99.800 ;
        RECT 594.800 97.000 595.600 99.800 ;
        RECT 596.400 97.000 597.200 99.800 ;
        RECT 598.000 97.000 598.800 99.800 ;
        RECT 580.200 95.800 582.800 96.600 ;
        RECT 599.600 96.600 600.400 99.800 ;
        RECT 586.200 95.800 590.800 96.400 ;
        RECT 580.200 95.200 581.000 95.800 ;
        RECT 578.000 94.400 581.000 95.200 ;
        RECT 570.800 91.600 571.600 93.200 ;
        RECT 567.600 88.800 568.400 90.400 ;
        RECT 572.200 90.200 572.800 93.600 ;
        RECT 575.600 93.000 584.400 93.800 ;
        RECT 586.200 93.400 587.000 95.800 ;
        RECT 590.000 95.600 590.800 95.800 ;
        RECT 591.600 95.600 593.200 96.400 ;
        RECT 596.200 95.600 597.200 96.400 ;
        RECT 599.600 95.800 602.000 96.600 ;
        RECT 588.400 93.600 589.200 95.200 ;
        RECT 590.000 94.800 590.800 95.000 ;
        RECT 590.000 94.200 594.400 94.800 ;
        RECT 593.600 94.000 594.400 94.200 ;
        RECT 574.000 90.200 574.800 90.400 ;
        RECT 571.800 89.600 572.800 90.200 ;
        RECT 573.400 89.600 574.800 90.200 ;
        RECT 571.800 84.400 572.600 89.600 ;
        RECT 573.400 88.400 574.000 89.600 ;
        RECT 573.200 87.600 574.000 88.400 ;
        RECT 575.600 87.400 576.400 93.000 ;
        RECT 585.000 92.600 587.000 93.400 ;
        RECT 590.800 92.600 594.000 93.400 ;
        RECT 596.400 92.800 597.200 95.600 ;
        RECT 601.200 95.200 602.000 95.800 ;
        RECT 601.200 94.600 603.000 95.200 ;
        RECT 602.200 93.400 603.000 94.600 ;
        RECT 606.000 94.600 606.800 99.800 ;
        RECT 607.600 96.000 608.400 99.800 ;
        RECT 607.600 95.200 608.600 96.000 ;
        RECT 606.000 94.000 607.200 94.600 ;
        RECT 602.200 92.600 606.000 93.400 ;
        RECT 577.000 92.000 577.800 92.200 ;
        RECT 578.800 92.000 579.600 92.400 ;
        RECT 582.000 92.000 582.800 92.400 ;
        RECT 588.400 92.000 589.200 92.400 ;
        RECT 599.600 92.000 600.400 92.600 ;
        RECT 606.600 92.000 607.200 94.000 ;
        RECT 577.000 91.400 600.400 92.000 ;
        RECT 606.400 91.400 607.200 92.000 ;
        RECT 606.400 89.600 607.000 91.400 ;
        RECT 607.800 90.800 608.600 95.200 ;
        RECT 585.200 89.400 586.000 89.600 ;
        RECT 580.600 89.000 586.000 89.400 ;
        RECT 579.800 88.800 586.000 89.000 ;
        RECT 587.000 89.000 595.600 89.600 ;
        RECT 577.200 88.000 578.800 88.800 ;
        RECT 579.800 88.200 581.200 88.800 ;
        RECT 587.000 88.200 587.600 89.000 ;
        RECT 594.800 88.800 595.600 89.000 ;
        RECT 598.000 89.000 607.000 89.600 ;
        RECT 598.000 88.800 598.800 89.000 ;
        RECT 578.200 87.600 578.800 88.000 ;
        RECT 581.800 87.600 587.600 88.200 ;
        RECT 588.200 87.600 590.800 88.400 ;
        RECT 575.600 86.800 577.600 87.400 ;
        RECT 578.200 86.800 582.400 87.600 ;
        RECT 577.000 86.200 577.600 86.800 ;
        RECT 577.000 85.600 578.000 86.200 ;
        RECT 570.800 83.600 572.600 84.400 ;
        RECT 571.800 82.200 572.600 83.600 ;
        RECT 577.200 82.200 578.000 85.600 ;
        RECT 580.400 82.200 581.200 86.800 ;
        RECT 583.600 82.200 584.400 85.000 ;
        RECT 585.200 82.200 586.000 85.000 ;
        RECT 586.800 82.200 587.600 87.000 ;
        RECT 590.000 82.200 590.800 87.000 ;
        RECT 593.200 82.200 594.000 88.400 ;
        RECT 601.200 87.600 603.800 88.400 ;
        RECT 596.400 86.800 600.600 87.600 ;
        RECT 594.800 82.200 595.600 85.000 ;
        RECT 596.400 82.200 597.200 85.000 ;
        RECT 598.000 82.200 598.800 85.000 ;
        RECT 601.200 82.200 602.000 87.600 ;
        RECT 606.400 87.400 607.000 89.000 ;
        RECT 604.400 86.800 607.000 87.400 ;
        RECT 607.600 90.000 608.600 90.800 ;
        RECT 604.400 82.200 605.200 86.800 ;
        RECT 607.600 82.200 608.400 90.000 ;
        RECT 2.800 68.300 3.600 79.800 ;
        RECT 7.000 72.400 7.800 79.800 ;
        RECT 8.400 73.600 9.200 74.400 ;
        RECT 8.600 72.400 9.200 73.600 ;
        RECT 11.600 73.600 12.400 74.400 ;
        RECT 11.600 72.400 12.200 73.600 ;
        RECT 13.000 72.400 13.800 79.800 ;
        RECT 18.800 74.300 19.600 79.800 ;
        RECT 20.400 74.300 21.200 74.400 ;
        RECT 18.800 73.700 21.200 74.300 ;
        RECT 7.000 71.800 8.000 72.400 ;
        RECT 8.600 71.800 10.000 72.400 ;
        RECT 6.000 68.800 6.800 70.400 ;
        RECT 7.400 68.400 8.000 71.800 ;
        RECT 9.200 71.600 10.000 71.800 ;
        RECT 10.800 71.800 12.200 72.400 ;
        RECT 12.800 71.800 13.800 72.400 ;
        RECT 10.800 71.600 11.600 71.800 ;
        RECT 9.300 70.300 9.900 71.600 ;
        RECT 12.800 70.300 13.400 71.800 ;
        RECT 17.200 71.600 18.000 73.200 ;
        RECT 9.300 69.700 13.400 70.300 ;
        RECT 12.800 68.400 13.400 69.700 ;
        RECT 14.000 68.800 14.800 70.400 ;
        RECT 4.400 68.300 5.200 68.400 ;
        RECT 2.800 68.200 5.200 68.300 ;
        RECT 2.800 67.700 6.000 68.200 ;
        RECT 2.800 62.200 3.600 67.700 ;
        RECT 4.400 67.600 6.000 67.700 ;
        RECT 7.400 67.600 10.000 68.400 ;
        RECT 10.800 67.600 13.400 68.400 ;
        RECT 15.600 68.200 16.400 68.400 ;
        RECT 14.800 67.600 16.400 68.200 ;
        RECT 5.200 67.200 6.000 67.600 ;
        RECT 4.600 66.200 8.200 66.600 ;
        RECT 9.200 66.200 9.800 67.600 ;
        RECT 11.000 66.200 11.600 67.600 ;
        RECT 14.800 67.200 15.600 67.600 ;
        RECT 12.600 66.200 16.200 66.600 ;
        RECT 18.800 66.200 19.600 73.700 ;
        RECT 20.400 73.600 21.200 73.700 ;
        RECT 25.800 72.800 26.600 79.800 ;
        RECT 30.000 75.000 30.800 79.000 ;
        RECT 25.000 72.200 26.600 72.800 ;
        RECT 23.600 69.600 24.400 71.200 ;
        RECT 25.000 70.400 25.600 72.200 ;
        RECT 30.200 71.600 30.800 75.000 ;
        RECT 34.200 72.400 35.000 79.800 ;
        RECT 35.600 73.600 36.400 74.400 ;
        RECT 35.800 72.400 36.400 73.600 ;
        RECT 38.800 73.600 39.600 74.400 ;
        RECT 38.800 72.400 39.400 73.600 ;
        RECT 40.200 72.400 41.000 79.800 ;
        RECT 34.200 71.800 35.200 72.400 ;
        RECT 35.800 71.800 37.200 72.400 ;
        RECT 27.000 71.000 30.800 71.600 ;
        RECT 25.000 69.600 26.000 70.400 ;
        RECT 25.000 68.400 25.600 69.600 ;
        RECT 27.000 69.000 27.600 71.000 ;
        RECT 20.400 68.300 21.200 68.400 ;
        RECT 22.000 68.300 22.800 68.400 ;
        RECT 20.400 67.700 22.800 68.300 ;
        RECT 20.400 66.800 21.200 67.700 ;
        RECT 22.000 67.600 22.800 67.700 ;
        RECT 23.600 67.600 25.600 68.400 ;
        RECT 26.200 68.200 27.600 69.000 ;
        RECT 28.400 68.800 29.200 70.400 ;
        RECT 30.000 68.800 30.800 70.400 ;
        RECT 33.200 68.800 34.000 70.400 ;
        RECT 34.600 68.400 35.200 71.800 ;
        RECT 36.400 71.600 37.200 71.800 ;
        RECT 38.000 71.800 39.400 72.400 ;
        RECT 40.000 71.800 41.000 72.400 ;
        RECT 38.000 71.600 38.800 71.800 ;
        RECT 36.500 70.300 37.100 71.600 ;
        RECT 40.000 70.300 40.600 71.800 ;
        RECT 44.400 71.400 45.200 79.800 ;
        RECT 48.800 76.400 49.600 79.800 ;
        RECT 47.600 75.800 49.600 76.400 ;
        RECT 53.200 75.800 54.000 79.800 ;
        RECT 57.400 75.800 58.600 79.800 ;
        RECT 47.600 75.000 48.400 75.800 ;
        RECT 53.200 75.200 53.800 75.800 ;
        RECT 51.000 74.600 54.600 75.200 ;
        RECT 57.200 75.000 58.000 75.800 ;
        RECT 51.000 74.400 51.800 74.600 ;
        RECT 53.800 74.400 54.600 74.600 ;
        RECT 47.600 73.000 48.400 73.200 ;
        RECT 52.200 73.000 53.000 73.200 ;
        RECT 47.600 72.400 53.000 73.000 ;
        RECT 53.600 73.000 55.800 73.600 ;
        RECT 53.600 71.800 54.200 73.000 ;
        RECT 55.000 72.800 55.800 73.000 ;
        RECT 57.400 73.200 58.800 74.000 ;
        RECT 57.400 72.200 58.000 73.200 ;
        RECT 49.400 71.400 54.200 71.800 ;
        RECT 44.400 71.200 54.200 71.400 ;
        RECT 55.600 71.600 58.000 72.200 ;
        RECT 44.400 71.000 50.200 71.200 ;
        RECT 44.400 70.800 50.000 71.000 ;
        RECT 55.600 70.400 56.200 71.600 ;
        RECT 62.000 71.200 62.800 79.800 ;
        RECT 66.200 78.400 67.000 79.800 ;
        RECT 65.200 77.600 67.000 78.400 ;
        RECT 66.200 72.400 67.000 77.600 ;
        RECT 67.600 73.600 68.400 74.400 ;
        RECT 67.800 72.400 68.400 73.600 ;
        RECT 72.600 72.400 73.400 79.800 ;
        RECT 78.600 74.400 79.400 79.800 ;
        RECT 82.800 75.000 83.600 79.000 ;
        RECT 74.000 73.600 74.800 74.400 ;
        RECT 74.200 72.400 74.800 73.600 ;
        RECT 77.200 73.600 78.000 74.400 ;
        RECT 78.600 73.600 80.400 74.400 ;
        RECT 77.200 72.400 77.800 73.600 ;
        RECT 78.600 72.400 79.400 73.600 ;
        RECT 66.200 71.800 67.200 72.400 ;
        RECT 67.800 71.800 69.200 72.400 ;
        RECT 72.600 71.800 73.600 72.400 ;
        RECT 74.200 71.800 75.600 72.400 ;
        RECT 58.600 70.600 62.800 71.200 ;
        RECT 58.600 70.400 59.400 70.600 ;
        RECT 36.500 69.700 40.600 70.300 ;
        RECT 40.000 68.400 40.600 69.700 ;
        RECT 41.200 68.800 42.000 70.400 ;
        RECT 50.800 70.200 51.600 70.400 ;
        RECT 46.600 69.600 51.600 70.200 ;
        RECT 55.600 69.600 56.400 70.400 ;
        RECT 60.200 69.800 61.000 70.000 ;
        RECT 46.600 69.400 47.400 69.600 ;
        RECT 49.200 69.400 50.000 69.600 ;
        RECT 48.200 68.400 49.000 68.600 ;
        RECT 55.600 68.400 56.200 69.600 ;
        RECT 57.200 69.200 61.000 69.800 ;
        RECT 57.200 69.000 58.000 69.200 ;
        RECT 25.000 67.000 25.600 67.600 ;
        RECT 26.600 67.800 27.600 68.200 ;
        RECT 31.600 68.200 32.400 68.400 ;
        RECT 26.600 67.200 30.800 67.800 ;
        RECT 31.600 67.600 33.200 68.200 ;
        RECT 34.600 67.600 37.200 68.400 ;
        RECT 38.000 67.600 40.600 68.400 ;
        RECT 42.800 68.200 43.600 68.400 ;
        RECT 42.000 67.600 43.600 68.200 ;
        RECT 45.200 67.800 56.200 68.400 ;
        RECT 45.200 67.600 46.800 67.800 ;
        RECT 32.400 67.200 33.200 67.600 ;
        RECT 4.400 66.000 8.400 66.200 ;
        RECT 4.400 62.200 5.200 66.000 ;
        RECT 7.600 62.200 8.400 66.000 ;
        RECT 9.200 62.200 10.000 66.200 ;
        RECT 10.800 62.200 11.600 66.200 ;
        RECT 12.400 66.000 16.400 66.200 ;
        RECT 12.400 62.200 13.200 66.000 ;
        RECT 15.600 62.200 16.400 66.000 ;
        RECT 17.800 65.600 19.600 66.200 ;
        RECT 25.000 66.600 25.800 67.000 ;
        RECT 25.000 66.000 26.600 66.600 ;
        RECT 17.800 62.200 18.600 65.600 ;
        RECT 25.800 63.000 26.600 66.000 ;
        RECT 30.200 65.000 30.800 67.200 ;
        RECT 31.800 66.200 35.400 66.600 ;
        RECT 36.400 66.200 37.000 67.600 ;
        RECT 38.200 66.200 38.800 67.600 ;
        RECT 42.000 67.200 42.800 67.600 ;
        RECT 39.800 66.200 43.400 66.600 ;
        RECT 30.000 63.000 30.800 65.000 ;
        RECT 31.600 66.000 35.600 66.200 ;
        RECT 31.600 62.200 32.400 66.000 ;
        RECT 34.800 62.200 35.600 66.000 ;
        RECT 36.400 62.200 37.200 66.200 ;
        RECT 38.000 62.200 38.800 66.200 ;
        RECT 39.600 66.000 43.600 66.200 ;
        RECT 39.600 62.200 40.400 66.000 ;
        RECT 42.800 62.200 43.600 66.000 ;
        RECT 44.400 62.200 45.200 67.000 ;
        RECT 49.400 66.400 50.000 67.800 ;
        RECT 55.000 67.600 55.800 67.800 ;
        RECT 62.000 67.200 62.800 70.600 ;
        RECT 65.200 68.800 66.000 70.400 ;
        RECT 66.600 68.400 67.200 71.800 ;
        RECT 68.400 71.600 69.200 71.800 ;
        RECT 71.600 68.800 72.400 70.400 ;
        RECT 73.000 70.300 73.600 71.800 ;
        RECT 74.800 71.600 75.600 71.800 ;
        RECT 76.400 71.800 77.800 72.400 ;
        RECT 78.400 71.800 79.400 72.400 ;
        RECT 76.400 71.600 77.200 71.800 ;
        RECT 76.500 70.300 77.100 71.600 ;
        RECT 73.000 69.700 77.100 70.300 ;
        RECT 73.000 68.400 73.600 69.700 ;
        RECT 78.400 68.400 79.000 71.800 ;
        RECT 82.800 71.600 83.400 75.000 ;
        RECT 87.000 72.800 87.800 79.800 ;
        RECT 94.000 72.800 94.800 79.800 ;
        RECT 87.000 72.200 88.600 72.800 ;
        RECT 82.800 71.000 86.600 71.600 ;
        RECT 79.600 68.800 80.400 70.400 ;
        RECT 82.800 68.800 83.600 70.400 ;
        RECT 84.400 68.800 85.200 70.400 ;
        RECT 86.000 69.000 86.600 71.000 ;
        RECT 63.600 68.200 64.400 68.400 ;
        RECT 63.600 67.600 65.200 68.200 ;
        RECT 66.600 67.600 69.200 68.400 ;
        RECT 70.000 68.200 70.800 68.400 ;
        RECT 70.000 67.600 71.600 68.200 ;
        RECT 73.000 67.600 75.600 68.400 ;
        RECT 76.400 67.600 79.000 68.400 ;
        RECT 81.200 68.200 82.000 68.400 ;
        RECT 80.400 67.600 82.000 68.200 ;
        RECT 86.000 68.200 87.400 69.000 ;
        RECT 88.000 68.400 88.600 72.200 ;
        RECT 93.800 71.800 94.800 72.800 ;
        RECT 97.200 72.400 98.000 79.800 ;
        RECT 95.400 71.800 98.000 72.400 ;
        RECT 89.200 70.300 90.000 71.200 ;
        RECT 92.400 70.300 93.200 70.400 ;
        RECT 89.200 69.700 93.200 70.300 ;
        RECT 89.200 69.600 90.000 69.700 ;
        RECT 92.400 69.600 93.200 69.700 ;
        RECT 93.800 68.400 94.400 71.800 ;
        RECT 95.400 69.800 96.000 71.800 ;
        RECT 95.000 69.000 96.000 69.800 ;
        RECT 86.000 67.800 87.000 68.200 ;
        RECT 64.400 67.200 65.200 67.600 ;
        RECT 59.000 66.600 62.800 67.200 ;
        RECT 59.000 66.400 59.800 66.600 ;
        RECT 47.600 64.200 48.400 65.000 ;
        RECT 49.200 64.800 50.000 66.400 ;
        RECT 51.000 65.400 51.800 65.600 ;
        RECT 51.000 64.800 53.800 65.400 ;
        RECT 53.200 64.200 53.800 64.800 ;
        RECT 57.200 64.200 58.000 65.000 ;
        RECT 47.600 63.600 49.600 64.200 ;
        RECT 48.800 62.200 49.600 63.600 ;
        RECT 53.200 62.200 54.000 64.200 ;
        RECT 57.200 63.600 58.600 64.200 ;
        RECT 57.400 62.200 58.600 63.600 ;
        RECT 62.000 62.200 62.800 66.600 ;
        RECT 63.800 66.200 67.400 66.600 ;
        RECT 68.400 66.200 69.000 67.600 ;
        RECT 70.800 67.200 71.600 67.600 ;
        RECT 70.200 66.200 73.800 66.600 ;
        RECT 74.800 66.200 75.400 67.600 ;
        RECT 76.600 66.200 77.200 67.600 ;
        RECT 80.400 67.200 81.200 67.600 ;
        RECT 82.800 67.200 87.000 67.800 ;
        RECT 88.000 67.600 90.000 68.400 ;
        RECT 90.800 68.300 91.600 68.400 ;
        RECT 93.800 68.300 94.800 68.400 ;
        RECT 90.800 67.700 94.800 68.300 ;
        RECT 90.800 67.600 91.600 67.700 ;
        RECT 93.800 67.600 94.800 67.700 ;
        RECT 78.200 66.200 81.800 66.600 ;
        RECT 63.600 66.000 67.600 66.200 ;
        RECT 63.600 62.200 64.400 66.000 ;
        RECT 66.800 62.200 67.600 66.000 ;
        RECT 68.400 62.200 69.200 66.200 ;
        RECT 70.000 66.000 74.000 66.200 ;
        RECT 70.000 62.200 70.800 66.000 ;
        RECT 73.200 62.200 74.000 66.000 ;
        RECT 74.800 62.200 75.600 66.200 ;
        RECT 76.400 62.200 77.200 66.200 ;
        RECT 78.000 66.000 82.000 66.200 ;
        RECT 78.000 62.200 78.800 66.000 ;
        RECT 81.200 62.200 82.000 66.000 ;
        RECT 82.800 65.000 83.400 67.200 ;
        RECT 88.000 67.000 88.600 67.600 ;
        RECT 87.800 66.600 88.600 67.000 ;
        RECT 87.000 66.400 88.600 66.600 ;
        RECT 86.000 66.000 88.600 66.400 ;
        RECT 93.800 66.200 94.400 67.600 ;
        RECT 95.400 67.400 96.000 69.000 ;
        RECT 97.000 70.300 98.000 70.400 ;
        RECT 98.800 70.300 99.600 70.400 ;
        RECT 97.000 69.700 99.600 70.300 ;
        RECT 97.000 69.600 98.000 69.700 ;
        RECT 98.800 69.600 99.600 69.700 ;
        RECT 97.000 68.800 97.800 69.600 ;
        RECT 95.400 66.800 98.000 67.400 ;
        RECT 86.000 65.600 87.800 66.000 ;
        RECT 93.800 65.600 94.800 66.200 ;
        RECT 82.800 63.000 83.600 65.000 ;
        RECT 87.000 63.000 87.800 65.600 ;
        RECT 94.000 62.200 94.800 65.600 ;
        RECT 97.200 62.200 98.000 66.800 ;
        RECT 98.800 64.800 99.600 66.400 ;
        RECT 100.400 62.200 101.200 79.800 ;
        RECT 102.000 64.800 102.800 66.400 ;
        RECT 103.600 62.200 104.400 79.800 ;
        RECT 105.200 64.800 106.000 66.400 ;
        RECT 106.800 62.200 107.600 79.800 ;
        RECT 108.400 71.200 109.200 79.800 ;
        RECT 112.600 75.800 113.800 79.800 ;
        RECT 117.200 75.800 118.000 79.800 ;
        RECT 121.600 76.400 122.400 79.800 ;
        RECT 121.600 75.800 123.600 76.400 ;
        RECT 113.200 75.000 114.000 75.800 ;
        RECT 117.400 75.200 118.000 75.800 ;
        RECT 116.600 74.600 120.200 75.200 ;
        RECT 122.800 75.000 123.600 75.800 ;
        RECT 116.600 74.400 117.400 74.600 ;
        RECT 119.400 74.400 120.200 74.600 ;
        RECT 112.400 73.200 113.800 74.000 ;
        RECT 113.200 72.200 113.800 73.200 ;
        RECT 115.400 73.000 117.600 73.600 ;
        RECT 115.400 72.800 116.200 73.000 ;
        RECT 113.200 71.600 115.600 72.200 ;
        RECT 108.400 70.600 112.600 71.200 ;
        RECT 108.400 67.200 109.200 70.600 ;
        RECT 111.800 70.400 112.600 70.600 ;
        RECT 110.200 69.800 111.000 70.000 ;
        RECT 110.200 69.200 114.000 69.800 ;
        RECT 113.200 69.000 114.000 69.200 ;
        RECT 115.000 68.400 115.600 71.600 ;
        RECT 117.000 71.800 117.600 73.000 ;
        RECT 118.200 73.000 119.000 73.200 ;
        RECT 122.800 73.000 123.600 73.200 ;
        RECT 118.200 72.400 123.600 73.000 ;
        RECT 117.000 71.400 121.800 71.800 ;
        RECT 126.000 71.400 126.800 79.800 ;
        RECT 117.000 71.200 126.800 71.400 ;
        RECT 121.000 71.000 126.800 71.200 ;
        RECT 121.200 70.800 126.800 71.000 ;
        RECT 119.600 70.200 120.400 70.400 ;
        RECT 119.600 69.600 124.600 70.200 ;
        RECT 123.800 69.400 124.600 69.600 ;
        RECT 122.200 68.400 123.000 68.600 ;
        RECT 115.000 67.800 126.000 68.400 ;
        RECT 115.400 67.600 116.200 67.800 ;
        RECT 118.000 67.600 118.800 67.800 ;
        RECT 108.400 66.600 112.200 67.200 ;
        RECT 108.400 62.200 109.200 66.600 ;
        RECT 111.400 66.400 112.200 66.600 ;
        RECT 121.200 65.600 121.800 67.800 ;
        RECT 124.400 67.600 126.000 67.800 ;
        RECT 119.400 65.400 120.200 65.600 ;
        RECT 113.200 64.200 114.000 65.000 ;
        RECT 117.400 64.800 120.200 65.400 ;
        RECT 121.200 64.800 122.000 65.600 ;
        RECT 117.400 64.200 118.000 64.800 ;
        RECT 122.800 64.200 123.600 65.000 ;
        RECT 112.600 63.600 114.000 64.200 ;
        RECT 112.600 62.200 113.800 63.600 ;
        RECT 117.200 62.200 118.000 64.200 ;
        RECT 121.600 63.600 123.600 64.200 ;
        RECT 121.600 62.200 122.400 63.600 ;
        RECT 126.000 62.200 126.800 67.000 ;
        RECT 127.600 62.200 128.400 79.800 ;
        RECT 129.200 64.800 130.000 66.400 ;
        RECT 130.800 64.800 131.600 66.400 ;
        RECT 132.400 62.200 133.200 79.800 ;
        RECT 134.000 72.400 134.800 79.800 ;
        RECT 137.200 72.800 138.000 79.800 ;
        RECT 134.000 71.800 136.600 72.400 ;
        RECT 137.200 71.800 138.200 72.800 ;
        RECT 143.000 72.400 143.800 79.800 ;
        RECT 144.400 73.600 145.200 74.400 ;
        RECT 144.600 72.400 145.200 73.600 ;
        RECT 147.600 73.600 148.400 74.400 ;
        RECT 147.600 72.400 148.200 73.600 ;
        RECT 149.000 72.400 149.800 79.800 ;
        RECT 143.000 71.800 144.000 72.400 ;
        RECT 144.600 71.800 146.000 72.400 ;
        RECT 134.000 69.600 135.000 70.400 ;
        RECT 134.200 68.800 135.000 69.600 ;
        RECT 136.000 69.800 136.600 71.800 ;
        RECT 136.000 69.000 137.000 69.800 ;
        RECT 136.000 67.400 136.600 69.000 ;
        RECT 137.600 68.400 138.200 71.800 ;
        RECT 142.000 70.300 142.800 70.400 ;
        RECT 137.200 68.300 138.200 68.400 ;
        RECT 138.900 69.700 142.800 70.300 ;
        RECT 138.900 68.300 139.500 69.700 ;
        RECT 142.000 68.800 142.800 69.700 ;
        RECT 143.400 70.300 144.000 71.800 ;
        RECT 145.200 71.600 146.000 71.800 ;
        RECT 146.800 71.800 148.200 72.400 ;
        RECT 148.800 71.800 149.800 72.400 ;
        RECT 146.800 71.600 147.600 71.800 ;
        RECT 146.900 70.300 147.500 71.600 ;
        RECT 143.400 69.700 147.500 70.300 ;
        RECT 143.400 68.400 144.000 69.700 ;
        RECT 148.800 68.400 149.400 71.800 ;
        RECT 158.000 71.400 158.800 79.800 ;
        RECT 162.400 76.400 163.200 79.800 ;
        RECT 161.200 75.800 163.200 76.400 ;
        RECT 166.800 75.800 167.600 79.800 ;
        RECT 171.000 75.800 172.200 79.800 ;
        RECT 161.200 75.000 162.000 75.800 ;
        RECT 166.800 75.200 167.400 75.800 ;
        RECT 164.600 74.600 168.200 75.200 ;
        RECT 170.800 75.000 171.600 75.800 ;
        RECT 164.600 74.400 165.400 74.600 ;
        RECT 167.400 74.400 168.200 74.600 ;
        RECT 161.200 73.000 162.000 73.200 ;
        RECT 165.800 73.000 166.600 73.200 ;
        RECT 161.200 72.400 166.600 73.000 ;
        RECT 167.200 73.000 169.400 73.600 ;
        RECT 167.200 71.800 167.800 73.000 ;
        RECT 168.600 72.800 169.400 73.000 ;
        RECT 171.000 73.200 172.400 74.000 ;
        RECT 171.000 72.200 171.600 73.200 ;
        RECT 163.000 71.400 167.800 71.800 ;
        RECT 158.000 71.200 167.800 71.400 ;
        RECT 169.200 71.600 171.600 72.200 ;
        RECT 158.000 71.000 163.800 71.200 ;
        RECT 158.000 70.800 163.600 71.000 ;
        RECT 150.000 68.800 150.800 70.400 ;
        RECT 164.400 70.200 165.200 70.400 ;
        RECT 160.200 69.600 165.200 70.200 ;
        RECT 160.200 69.400 161.000 69.600 ;
        RECT 162.800 69.400 163.600 69.600 ;
        RECT 161.800 68.400 162.600 68.600 ;
        RECT 169.200 68.400 169.800 71.600 ;
        RECT 175.600 71.200 176.400 79.800 ;
        RECT 179.800 72.400 180.600 79.800 ;
        RECT 185.800 78.400 186.600 79.800 ;
        RECT 185.800 77.600 187.600 78.400 ;
        RECT 181.200 73.600 182.000 74.400 ;
        RECT 181.400 72.400 182.000 73.600 ;
        RECT 184.400 73.600 185.200 74.400 ;
        RECT 184.400 72.400 185.000 73.600 ;
        RECT 185.800 72.400 186.600 77.600 ;
        RECT 179.800 71.800 180.800 72.400 ;
        RECT 181.400 71.800 182.800 72.400 ;
        RECT 172.200 70.600 176.400 71.200 ;
        RECT 172.200 70.400 173.000 70.600 ;
        RECT 173.800 69.800 174.600 70.000 ;
        RECT 170.800 69.200 174.600 69.800 ;
        RECT 170.800 69.000 171.600 69.200 ;
        RECT 137.200 67.700 139.500 68.300 ;
        RECT 140.400 68.200 141.200 68.400 ;
        RECT 137.200 67.600 138.200 67.700 ;
        RECT 140.400 67.600 142.000 68.200 ;
        RECT 143.400 67.600 146.000 68.400 ;
        RECT 146.800 67.600 149.400 68.400 ;
        RECT 151.600 68.300 152.400 68.400 ;
        RECT 156.400 68.300 157.200 68.400 ;
        RECT 151.600 68.200 157.200 68.300 ;
        RECT 150.800 67.700 157.200 68.200 ;
        RECT 150.800 67.600 152.400 67.700 ;
        RECT 156.400 67.600 157.200 67.700 ;
        RECT 158.800 67.800 169.800 68.400 ;
        RECT 158.800 67.600 160.400 67.800 ;
        RECT 134.000 66.800 136.600 67.400 ;
        RECT 134.000 62.200 134.800 66.800 ;
        RECT 137.600 66.200 138.200 67.600 ;
        RECT 141.200 67.200 142.000 67.600 ;
        RECT 140.600 66.200 144.200 66.600 ;
        RECT 145.200 66.200 145.800 67.600 ;
        RECT 147.000 66.200 147.600 67.600 ;
        RECT 150.800 67.200 151.600 67.600 ;
        RECT 148.600 66.200 152.200 66.600 ;
        RECT 137.200 65.600 138.200 66.200 ;
        RECT 140.400 66.000 144.400 66.200 ;
        RECT 137.200 62.200 138.000 65.600 ;
        RECT 140.400 62.200 141.200 66.000 ;
        RECT 143.600 62.200 144.400 66.000 ;
        RECT 145.200 62.200 146.000 66.200 ;
        RECT 146.800 62.200 147.600 66.200 ;
        RECT 148.400 66.000 152.400 66.200 ;
        RECT 148.400 62.200 149.200 66.000 ;
        RECT 151.600 62.200 152.400 66.000 ;
        RECT 158.000 62.200 158.800 67.000 ;
        RECT 163.000 66.400 163.600 67.800 ;
        RECT 168.600 67.600 169.400 67.800 ;
        RECT 175.600 67.200 176.400 70.600 ;
        RECT 178.800 68.800 179.600 70.400 ;
        RECT 180.200 70.300 180.800 71.800 ;
        RECT 182.000 71.600 182.800 71.800 ;
        RECT 183.600 71.800 185.000 72.400 ;
        RECT 185.600 71.800 186.600 72.400 ;
        RECT 190.000 75.000 190.800 79.000 ;
        RECT 183.600 71.600 184.400 71.800 ;
        RECT 183.700 70.300 184.300 71.600 ;
        RECT 180.200 69.700 184.300 70.300 ;
        RECT 180.200 68.400 180.800 69.700 ;
        RECT 185.600 68.400 186.200 71.800 ;
        RECT 190.000 71.600 190.600 75.000 ;
        RECT 194.200 72.800 195.000 79.800 ;
        RECT 194.200 72.200 195.800 72.800 ;
        RECT 190.000 71.000 193.800 71.600 ;
        RECT 186.800 68.800 187.600 70.400 ;
        RECT 190.000 68.800 190.800 70.400 ;
        RECT 191.600 68.800 192.400 70.400 ;
        RECT 193.200 69.000 193.800 71.000 ;
        RECT 177.200 68.200 178.000 68.400 ;
        RECT 177.200 67.600 178.800 68.200 ;
        RECT 180.200 67.600 182.800 68.400 ;
        RECT 183.600 67.600 186.200 68.400 ;
        RECT 188.400 68.200 189.200 68.400 ;
        RECT 187.600 67.600 189.200 68.200 ;
        RECT 193.200 68.200 194.600 69.000 ;
        RECT 195.200 68.400 195.800 72.200 ;
        RECT 199.600 71.600 200.400 73.200 ;
        RECT 196.400 69.600 197.200 71.200 ;
        RECT 193.200 67.800 194.200 68.200 ;
        RECT 178.000 67.200 178.800 67.600 ;
        RECT 172.600 66.600 176.400 67.200 ;
        RECT 172.600 66.400 173.400 66.600 ;
        RECT 161.200 64.200 162.000 65.000 ;
        RECT 162.800 64.800 163.600 66.400 ;
        RECT 164.600 65.400 165.400 65.600 ;
        RECT 164.600 64.800 167.400 65.400 ;
        RECT 166.800 64.200 167.400 64.800 ;
        RECT 170.800 64.200 171.600 65.000 ;
        RECT 161.200 63.600 163.200 64.200 ;
        RECT 162.400 62.200 163.200 63.600 ;
        RECT 166.800 62.200 167.600 64.200 ;
        RECT 170.800 63.600 172.200 64.200 ;
        RECT 171.000 62.200 172.200 63.600 ;
        RECT 175.600 62.200 176.400 66.600 ;
        RECT 177.400 66.200 181.000 66.600 ;
        RECT 182.000 66.200 182.600 67.600 ;
        RECT 183.800 66.200 184.400 67.600 ;
        RECT 187.600 67.200 188.400 67.600 ;
        RECT 190.000 67.200 194.200 67.800 ;
        RECT 195.200 67.600 197.200 68.400 ;
        RECT 185.400 66.200 189.000 66.600 ;
        RECT 177.200 66.000 181.200 66.200 ;
        RECT 177.200 62.200 178.000 66.000 ;
        RECT 180.400 62.200 181.200 66.000 ;
        RECT 182.000 62.200 182.800 66.200 ;
        RECT 183.600 62.200 184.400 66.200 ;
        RECT 185.200 66.000 189.200 66.200 ;
        RECT 185.200 62.200 186.000 66.000 ;
        RECT 188.400 62.200 189.200 66.000 ;
        RECT 190.000 65.000 190.600 67.200 ;
        RECT 195.200 67.000 195.800 67.600 ;
        RECT 195.000 66.600 195.800 67.000 ;
        RECT 194.200 66.400 195.800 66.600 ;
        RECT 193.200 66.000 195.800 66.400 ;
        RECT 201.200 66.200 202.000 79.800 ;
        RECT 206.000 76.400 206.800 79.800 ;
        RECT 205.800 75.800 206.800 76.400 ;
        RECT 205.800 75.200 206.400 75.800 ;
        RECT 209.200 75.200 210.000 79.800 ;
        RECT 212.400 77.000 213.200 79.800 ;
        RECT 214.000 77.000 214.800 79.800 ;
        RECT 204.400 74.600 206.400 75.200 ;
        RECT 204.400 69.000 205.200 74.600 ;
        RECT 207.000 74.400 211.200 75.200 ;
        RECT 215.600 75.000 216.400 79.800 ;
        RECT 218.800 75.000 219.600 79.800 ;
        RECT 207.000 74.000 207.600 74.400 ;
        RECT 206.000 73.200 207.600 74.000 ;
        RECT 210.600 73.800 216.400 74.400 ;
        RECT 208.600 73.200 210.000 73.800 ;
        RECT 208.600 73.000 214.800 73.200 ;
        RECT 209.400 72.600 214.800 73.000 ;
        RECT 214.000 72.400 214.800 72.600 ;
        RECT 215.800 73.000 216.400 73.800 ;
        RECT 217.000 73.600 219.600 74.400 ;
        RECT 222.000 73.600 222.800 79.800 ;
        RECT 223.600 77.000 224.400 79.800 ;
        RECT 225.200 77.000 226.000 79.800 ;
        RECT 226.800 77.000 227.600 79.800 ;
        RECT 225.200 74.400 229.400 75.200 ;
        RECT 230.000 74.400 230.800 79.800 ;
        RECT 233.200 75.200 234.000 79.800 ;
        RECT 233.200 74.600 235.800 75.200 ;
        RECT 230.000 73.600 232.600 74.400 ;
        RECT 223.600 73.000 224.400 73.200 ;
        RECT 215.800 72.400 224.400 73.000 ;
        RECT 226.800 73.000 227.600 73.200 ;
        RECT 235.200 73.000 235.800 74.600 ;
        RECT 226.800 72.400 235.800 73.000 ;
        RECT 235.200 70.600 235.800 72.400 ;
        RECT 236.400 74.300 237.200 79.800 ;
        RECT 240.400 74.300 241.200 74.400 ;
        RECT 236.400 73.700 241.200 74.300 ;
        RECT 236.400 72.000 237.200 73.700 ;
        RECT 240.400 73.600 241.200 73.700 ;
        RECT 240.400 72.400 241.000 73.600 ;
        RECT 241.800 72.400 242.600 79.800 ;
        RECT 236.400 71.200 237.400 72.000 ;
        RECT 239.600 71.800 241.000 72.400 ;
        RECT 241.600 71.800 242.600 72.400 ;
        RECT 248.600 72.400 249.400 79.800 ;
        RECT 250.000 74.300 250.800 74.400 ;
        RECT 252.400 74.300 253.200 74.400 ;
        RECT 250.000 73.700 253.200 74.300 ;
        RECT 250.000 73.600 250.800 73.700 ;
        RECT 252.400 73.600 253.200 73.700 ;
        RECT 250.200 72.400 250.800 73.600 ;
        RECT 248.600 71.800 249.600 72.400 ;
        RECT 250.200 71.800 251.600 72.400 ;
        RECT 239.600 71.600 240.400 71.800 ;
        RECT 205.800 70.000 229.200 70.600 ;
        RECT 235.200 70.000 236.000 70.600 ;
        RECT 205.800 69.800 206.600 70.000 ;
        RECT 207.600 69.600 208.400 70.000 ;
        RECT 210.800 69.600 211.600 70.000 ;
        RECT 228.400 69.400 229.200 70.000 ;
        RECT 202.800 66.800 203.600 68.400 ;
        RECT 204.400 68.200 213.200 69.000 ;
        RECT 213.800 68.600 215.800 69.400 ;
        RECT 219.600 68.600 222.800 69.400 ;
        RECT 193.200 65.600 195.000 66.000 ;
        RECT 190.000 63.000 190.800 65.000 ;
        RECT 194.200 63.000 195.000 65.600 ;
        RECT 200.200 65.600 202.000 66.200 ;
        RECT 200.200 62.200 201.000 65.600 ;
        RECT 204.400 62.200 205.200 68.200 ;
        RECT 206.800 66.800 209.800 67.600 ;
        RECT 209.000 66.200 209.800 66.800 ;
        RECT 215.000 66.200 215.800 68.600 ;
        RECT 217.200 66.800 218.000 68.400 ;
        RECT 222.400 67.800 223.200 68.000 ;
        RECT 218.800 67.200 223.200 67.800 ;
        RECT 218.800 67.000 219.600 67.200 ;
        RECT 225.200 66.400 226.000 69.200 ;
        RECT 231.000 68.600 234.800 69.400 ;
        RECT 231.000 67.400 231.800 68.600 ;
        RECT 235.400 68.000 236.000 70.000 ;
        RECT 218.800 66.200 219.600 66.400 ;
        RECT 209.000 65.400 211.600 66.200 ;
        RECT 215.000 65.600 219.600 66.200 ;
        RECT 220.400 65.600 222.000 66.400 ;
        RECT 225.000 65.600 226.000 66.400 ;
        RECT 230.000 66.800 231.800 67.400 ;
        RECT 234.800 67.400 236.000 68.000 ;
        RECT 230.000 66.200 230.800 66.800 ;
        RECT 210.800 62.200 211.600 65.400 ;
        RECT 228.400 65.400 230.800 66.200 ;
        RECT 212.400 62.200 213.200 65.000 ;
        RECT 214.000 62.200 214.800 65.000 ;
        RECT 215.600 62.200 216.400 65.000 ;
        RECT 218.800 62.200 219.600 65.000 ;
        RECT 222.000 62.200 222.800 65.000 ;
        RECT 223.600 62.200 224.400 65.000 ;
        RECT 225.200 62.200 226.000 65.000 ;
        RECT 226.800 62.200 227.600 65.000 ;
        RECT 228.400 62.200 229.200 65.400 ;
        RECT 234.800 62.200 235.600 67.400 ;
        RECT 236.600 66.800 237.400 71.200 ;
        RECT 238.000 70.300 238.800 70.400 ;
        RECT 241.600 70.300 242.200 71.800 ;
        RECT 238.000 69.700 242.200 70.300 ;
        RECT 238.000 69.600 238.800 69.700 ;
        RECT 241.600 68.400 242.200 69.700 ;
        RECT 242.800 70.300 243.600 70.400 ;
        RECT 247.600 70.300 248.400 70.400 ;
        RECT 242.800 69.700 248.400 70.300 ;
        RECT 242.800 68.800 243.600 69.700 ;
        RECT 247.600 68.800 248.400 69.700 ;
        RECT 249.000 68.400 249.600 71.800 ;
        RECT 250.800 71.600 251.600 71.800 ;
        RECT 239.600 67.600 242.200 68.400 ;
        RECT 244.400 68.300 245.200 68.400 ;
        RECT 246.000 68.300 246.800 68.400 ;
        RECT 244.400 68.200 246.800 68.300 ;
        RECT 249.000 68.300 251.600 68.400 ;
        RECT 252.400 68.300 253.200 68.400 ;
        RECT 243.600 67.700 247.600 68.200 ;
        RECT 243.600 67.600 245.200 67.700 ;
        RECT 246.000 67.600 247.600 67.700 ;
        RECT 249.000 67.700 253.200 68.300 ;
        RECT 249.000 67.600 251.600 67.700 ;
        RECT 236.400 66.000 237.400 66.800 ;
        RECT 239.800 66.200 240.400 67.600 ;
        RECT 243.600 67.200 244.400 67.600 ;
        RECT 246.800 67.200 247.600 67.600 ;
        RECT 241.400 66.200 245.000 66.600 ;
        RECT 246.200 66.200 249.800 66.600 ;
        RECT 250.800 66.200 251.400 67.600 ;
        RECT 252.400 66.800 253.200 67.700 ;
        RECT 254.000 68.300 254.800 79.800 ;
        RECT 255.600 71.600 256.400 73.200 ;
        RECT 258.800 72.000 259.600 79.800 ;
        RECT 262.000 75.200 262.800 79.800 ;
        RECT 258.600 71.200 259.600 72.000 ;
        RECT 260.200 74.600 262.800 75.200 ;
        RECT 260.200 73.000 260.800 74.600 ;
        RECT 265.200 74.400 266.000 79.800 ;
        RECT 268.400 77.000 269.200 79.800 ;
        RECT 270.000 77.000 270.800 79.800 ;
        RECT 271.600 77.000 272.400 79.800 ;
        RECT 266.600 74.400 270.800 75.200 ;
        RECT 263.400 73.600 266.000 74.400 ;
        RECT 273.200 73.600 274.000 79.800 ;
        RECT 276.400 75.000 277.200 79.800 ;
        RECT 279.600 75.000 280.400 79.800 ;
        RECT 281.200 77.000 282.000 79.800 ;
        RECT 282.800 77.000 283.600 79.800 ;
        RECT 286.000 75.200 286.800 79.800 ;
        RECT 289.200 76.400 290.000 79.800 ;
        RECT 289.200 75.800 290.200 76.400 ;
        RECT 289.600 75.200 290.200 75.800 ;
        RECT 284.800 74.400 289.000 75.200 ;
        RECT 289.600 74.600 291.600 75.200 ;
        RECT 276.400 73.600 279.000 74.400 ;
        RECT 279.600 73.800 285.400 74.400 ;
        RECT 288.400 74.000 289.000 74.400 ;
        RECT 268.400 73.000 269.200 73.200 ;
        RECT 260.200 72.400 269.200 73.000 ;
        RECT 271.600 73.000 272.400 73.200 ;
        RECT 279.600 73.000 280.200 73.800 ;
        RECT 286.000 73.200 287.400 73.800 ;
        RECT 288.400 73.200 290.000 74.000 ;
        RECT 271.600 72.400 280.200 73.000 ;
        RECT 281.200 73.000 287.400 73.200 ;
        RECT 281.200 72.600 286.600 73.000 ;
        RECT 281.200 72.400 282.000 72.600 ;
        RECT 257.200 68.300 258.000 68.400 ;
        RECT 254.000 67.700 258.000 68.300 ;
        RECT 254.000 66.200 254.800 67.700 ;
        RECT 257.200 67.600 258.000 67.700 ;
        RECT 258.600 66.800 259.400 71.200 ;
        RECT 260.200 70.600 260.800 72.400 ;
        RECT 260.000 70.000 260.800 70.600 ;
        RECT 266.800 70.000 290.200 70.600 ;
        RECT 260.000 68.000 260.600 70.000 ;
        RECT 266.800 69.400 267.600 70.000 ;
        RECT 284.400 69.600 285.200 70.000 ;
        RECT 286.000 69.600 286.800 70.000 ;
        RECT 289.400 69.800 290.200 70.000 ;
        RECT 261.200 68.600 265.000 69.400 ;
        RECT 260.000 67.400 261.200 68.000 ;
        RECT 236.400 62.200 237.200 66.000 ;
        RECT 239.600 62.200 240.400 66.200 ;
        RECT 241.200 66.000 245.200 66.200 ;
        RECT 241.200 62.200 242.000 66.000 ;
        RECT 244.400 62.200 245.200 66.000 ;
        RECT 246.000 66.000 250.000 66.200 ;
        RECT 246.000 62.200 246.800 66.000 ;
        RECT 249.200 62.200 250.000 66.000 ;
        RECT 250.800 62.200 251.600 66.200 ;
        RECT 254.000 65.600 255.800 66.200 ;
        RECT 258.600 66.000 259.600 66.800 ;
        RECT 255.000 62.200 255.800 65.600 ;
        RECT 258.800 62.200 259.600 66.000 ;
        RECT 260.400 62.200 261.200 67.400 ;
        RECT 264.200 67.400 265.000 68.600 ;
        RECT 264.200 66.800 266.000 67.400 ;
        RECT 265.200 66.200 266.000 66.800 ;
        RECT 270.000 66.400 270.800 69.200 ;
        RECT 273.200 68.600 276.400 69.400 ;
        RECT 280.200 68.600 282.200 69.400 ;
        RECT 290.800 69.000 291.600 74.600 ;
        RECT 272.800 67.800 273.600 68.000 ;
        RECT 272.800 67.200 277.200 67.800 ;
        RECT 276.400 67.000 277.200 67.200 ;
        RECT 278.000 66.800 278.800 68.400 ;
        RECT 265.200 65.400 267.600 66.200 ;
        RECT 270.000 65.600 271.000 66.400 ;
        RECT 274.000 65.600 275.600 66.400 ;
        RECT 276.400 66.200 277.200 66.400 ;
        RECT 280.200 66.200 281.000 68.600 ;
        RECT 282.800 68.200 291.600 69.000 ;
        RECT 286.200 66.800 289.200 67.600 ;
        RECT 286.200 66.200 287.000 66.800 ;
        RECT 276.400 65.600 281.000 66.200 ;
        RECT 266.800 62.200 267.600 65.400 ;
        RECT 284.400 65.400 287.000 66.200 ;
        RECT 268.400 62.200 269.200 65.000 ;
        RECT 270.000 62.200 270.800 65.000 ;
        RECT 271.600 62.200 272.400 65.000 ;
        RECT 273.200 62.200 274.000 65.000 ;
        RECT 276.400 62.200 277.200 65.000 ;
        RECT 279.600 62.200 280.400 65.000 ;
        RECT 281.200 62.200 282.000 65.000 ;
        RECT 282.800 62.200 283.600 65.000 ;
        RECT 284.400 62.200 285.200 65.400 ;
        RECT 290.800 62.200 291.600 68.200 ;
        RECT 292.400 66.800 293.200 68.400 ;
        RECT 294.000 66.200 294.800 79.800 ;
        RECT 295.600 72.300 296.400 73.200 ;
        RECT 303.600 72.300 304.400 79.800 ;
        RECT 306.800 75.200 307.600 79.800 ;
        RECT 295.600 71.700 304.400 72.300 ;
        RECT 295.600 71.600 296.400 71.700 ;
        RECT 303.400 71.200 304.400 71.700 ;
        RECT 305.000 74.600 307.600 75.200 ;
        RECT 305.000 73.000 305.600 74.600 ;
        RECT 310.000 74.400 310.800 79.800 ;
        RECT 313.200 77.000 314.000 79.800 ;
        RECT 314.800 77.000 315.600 79.800 ;
        RECT 316.400 77.000 317.200 79.800 ;
        RECT 311.400 74.400 315.600 75.200 ;
        RECT 308.200 73.600 310.800 74.400 ;
        RECT 318.000 73.600 318.800 79.800 ;
        RECT 321.200 75.000 322.000 79.800 ;
        RECT 324.400 75.000 325.200 79.800 ;
        RECT 326.000 77.000 326.800 79.800 ;
        RECT 327.600 77.000 328.400 79.800 ;
        RECT 330.800 75.200 331.600 79.800 ;
        RECT 334.000 76.400 334.800 79.800 ;
        RECT 334.000 75.800 335.000 76.400 ;
        RECT 334.400 75.200 335.000 75.800 ;
        RECT 329.600 74.400 333.800 75.200 ;
        RECT 334.400 74.600 336.400 75.200 ;
        RECT 321.200 73.600 323.800 74.400 ;
        RECT 324.400 73.800 330.200 74.400 ;
        RECT 333.200 74.000 333.800 74.400 ;
        RECT 313.200 73.000 314.000 73.200 ;
        RECT 305.000 72.400 314.000 73.000 ;
        RECT 316.400 73.000 317.200 73.200 ;
        RECT 324.400 73.000 325.000 73.800 ;
        RECT 330.800 73.200 332.200 73.800 ;
        RECT 333.200 73.200 334.800 74.000 ;
        RECT 316.400 72.400 325.000 73.000 ;
        RECT 326.000 73.000 332.200 73.200 ;
        RECT 326.000 72.600 331.400 73.000 ;
        RECT 326.000 72.400 326.800 72.600 ;
        RECT 303.400 66.800 304.200 71.200 ;
        RECT 305.000 70.600 305.600 72.400 ;
        RECT 304.800 70.000 305.600 70.600 ;
        RECT 311.600 70.000 335.000 70.600 ;
        RECT 304.800 68.000 305.400 70.000 ;
        RECT 311.600 69.400 312.400 70.000 ;
        RECT 322.800 69.600 323.600 70.000 ;
        RECT 329.200 69.600 330.000 70.000 ;
        RECT 334.200 69.800 335.000 70.000 ;
        RECT 306.000 68.600 309.800 69.400 ;
        RECT 304.800 67.400 306.000 68.000 ;
        RECT 294.000 65.600 295.800 66.200 ;
        RECT 303.400 66.000 304.400 66.800 ;
        RECT 295.000 64.400 295.800 65.600 ;
        RECT 294.000 63.600 295.800 64.400 ;
        RECT 295.000 62.200 295.800 63.600 ;
        RECT 303.600 62.200 304.400 66.000 ;
        RECT 305.200 62.200 306.000 67.400 ;
        RECT 309.000 67.400 309.800 68.600 ;
        RECT 309.000 66.800 310.800 67.400 ;
        RECT 310.000 66.200 310.800 66.800 ;
        RECT 314.800 66.400 315.600 69.200 ;
        RECT 318.000 68.600 321.200 69.400 ;
        RECT 325.000 68.600 327.000 69.400 ;
        RECT 335.600 69.000 336.400 74.600 ;
        RECT 339.800 72.400 340.600 79.800 ;
        RECT 341.200 73.600 342.000 74.400 ;
        RECT 341.400 72.400 342.000 73.600 ;
        RECT 343.600 72.400 344.400 79.800 ;
        RECT 345.400 72.400 346.200 72.600 ;
        RECT 339.800 71.800 340.800 72.400 ;
        RECT 341.400 71.800 342.800 72.400 ;
        RECT 343.600 71.800 346.200 72.400 ;
        RECT 348.000 71.800 349.600 79.800 ;
        RECT 351.600 72.400 352.400 72.600 ;
        RECT 353.200 72.400 354.000 79.800 ;
        RECT 354.800 73.600 356.400 74.400 ;
        RECT 355.600 72.400 356.200 73.600 ;
        RECT 357.000 72.400 357.800 79.800 ;
        RECT 351.600 71.800 354.000 72.400 ;
        RECT 354.800 71.800 356.200 72.400 ;
        RECT 356.800 71.800 357.800 72.400 ;
        RECT 317.600 67.800 318.400 68.000 ;
        RECT 317.600 67.200 322.000 67.800 ;
        RECT 321.200 67.000 322.000 67.200 ;
        RECT 322.800 66.800 323.600 68.400 ;
        RECT 310.000 65.400 312.400 66.200 ;
        RECT 314.800 65.600 315.800 66.400 ;
        RECT 318.800 65.600 320.400 66.400 ;
        RECT 321.200 66.200 322.000 66.400 ;
        RECT 325.000 66.200 325.800 68.600 ;
        RECT 327.600 68.200 336.400 69.000 ;
        RECT 338.800 68.800 339.600 70.400 ;
        RECT 340.200 68.400 340.800 71.800 ;
        RECT 342.000 71.600 342.800 71.800 ;
        RECT 346.600 70.400 347.400 70.600 ;
        RECT 348.600 70.400 349.200 71.800 ;
        RECT 354.800 71.600 355.600 71.800 ;
        RECT 345.800 69.800 347.400 70.400 ;
        RECT 345.800 69.600 346.600 69.800 ;
        RECT 348.400 69.600 349.200 70.400 ;
        RECT 347.200 68.600 348.000 68.800 ;
        RECT 345.200 68.400 348.000 68.600 ;
        RECT 331.000 66.800 334.000 67.600 ;
        RECT 331.000 66.200 331.800 66.800 ;
        RECT 321.200 65.600 325.800 66.200 ;
        RECT 311.600 62.200 312.400 65.400 ;
        RECT 329.200 65.400 331.800 66.200 ;
        RECT 313.200 62.200 314.000 65.000 ;
        RECT 314.800 62.200 315.600 65.000 ;
        RECT 316.400 62.200 317.200 65.000 ;
        RECT 318.000 62.200 318.800 65.000 ;
        RECT 321.200 62.200 322.000 65.000 ;
        RECT 324.400 62.200 325.200 65.000 ;
        RECT 326.000 62.200 326.800 65.000 ;
        RECT 327.600 62.200 328.400 65.000 ;
        RECT 329.200 62.200 330.000 65.400 ;
        RECT 335.600 62.200 336.400 68.200 ;
        RECT 337.200 68.200 338.000 68.400 ;
        RECT 340.200 68.300 342.800 68.400 ;
        RECT 343.600 68.300 348.000 68.400 ;
        RECT 337.200 67.600 338.800 68.200 ;
        RECT 340.200 68.000 348.000 68.300 ;
        RECT 348.600 68.400 349.200 69.600 ;
        RECT 356.800 68.400 357.400 71.800 ;
        RECT 358.000 68.800 358.800 70.400 ;
        RECT 340.200 67.800 345.800 68.000 ;
        RECT 348.600 67.800 349.600 68.400 ;
        RECT 340.200 67.700 345.200 67.800 ;
        RECT 340.200 67.600 342.800 67.700 ;
        RECT 343.600 67.600 345.200 67.700 ;
        RECT 338.000 67.200 338.800 67.600 ;
        RECT 337.400 66.200 341.000 66.600 ;
        RECT 342.000 66.200 342.600 67.600 ;
        RECT 345.400 66.800 346.200 67.000 ;
        RECT 343.600 66.200 346.200 66.800 ;
        RECT 346.800 66.400 348.400 67.200 ;
        RECT 337.200 66.000 341.200 66.200 ;
        RECT 337.200 62.200 338.000 66.000 ;
        RECT 340.400 62.200 341.200 66.000 ;
        RECT 342.000 62.200 342.800 66.200 ;
        RECT 343.600 62.200 344.400 66.200 ;
        RECT 349.000 65.800 349.600 67.800 ;
        RECT 350.400 67.600 351.200 68.400 ;
        RECT 352.400 67.600 354.000 68.400 ;
        RECT 354.800 67.600 357.400 68.400 ;
        RECT 359.600 68.200 360.400 68.400 ;
        RECT 358.800 67.600 360.400 68.200 ;
        RECT 350.400 67.200 351.000 67.600 ;
        RECT 350.200 66.400 351.000 67.200 ;
        RECT 351.600 66.800 352.400 67.000 ;
        RECT 351.600 66.200 354.000 66.800 ;
        RECT 355.000 66.200 355.600 67.600 ;
        RECT 358.800 67.200 359.600 67.600 ;
        RECT 361.200 66.800 362.000 68.400 ;
        RECT 356.600 66.200 360.200 66.600 ;
        RECT 362.800 66.200 363.600 79.800 ;
        RECT 364.400 71.600 365.200 73.200 ;
        RECT 366.000 71.200 366.800 79.800 ;
        RECT 370.200 72.400 371.000 79.800 ;
        RECT 375.000 72.600 375.800 79.800 ;
        RECT 370.200 71.800 371.600 72.400 ;
        RECT 366.000 70.800 370.000 71.200 ;
        RECT 366.000 70.600 370.200 70.800 ;
        RECT 369.400 70.000 370.200 70.600 ;
        RECT 371.000 70.400 371.600 71.800 ;
        RECT 374.000 71.800 375.800 72.600 ;
        RECT 379.800 72.400 380.600 79.800 ;
        RECT 381.200 73.600 382.000 74.400 ;
        RECT 381.400 72.400 382.000 73.600 ;
        RECT 379.800 71.800 380.800 72.400 ;
        RECT 381.400 71.800 382.800 72.400 ;
        RECT 374.000 71.600 374.800 71.800 ;
        RECT 368.000 68.400 368.800 69.200 ;
        RECT 367.600 67.600 368.600 68.400 ;
        RECT 369.600 67.000 370.200 70.000 ;
        RECT 370.800 69.600 371.600 70.400 ;
        RECT 367.800 66.400 370.200 67.000 ;
        RECT 348.000 64.400 349.600 65.800 ;
        RECT 346.800 63.600 349.600 64.400 ;
        RECT 348.000 62.200 349.600 63.600 ;
        RECT 353.200 62.200 354.000 66.200 ;
        RECT 354.800 62.200 355.600 66.200 ;
        RECT 356.400 66.000 360.400 66.200 ;
        RECT 356.400 62.200 357.200 66.000 ;
        RECT 359.600 62.200 360.400 66.000 ;
        RECT 362.800 65.600 364.600 66.200 ;
        RECT 363.800 62.200 364.600 65.600 ;
        RECT 366.000 64.800 366.800 66.400 ;
        RECT 367.800 64.200 368.400 66.400 ;
        RECT 371.000 66.200 371.600 69.600 ;
        RECT 374.200 68.400 374.800 71.600 ;
        RECT 375.600 69.600 376.400 71.200 ;
        RECT 378.800 68.800 379.600 70.400 ;
        RECT 380.200 68.400 380.800 71.800 ;
        RECT 382.000 71.600 382.800 71.800 ;
        RECT 374.000 67.600 374.800 68.400 ;
        RECT 377.200 68.200 378.000 68.400 ;
        RECT 380.200 68.300 382.800 68.400 ;
        RECT 383.600 68.300 384.400 68.400 ;
        RECT 377.200 67.600 378.800 68.200 ;
        RECT 380.200 67.700 384.400 68.300 ;
        RECT 380.200 67.600 382.800 67.700 ;
        RECT 367.600 62.200 368.400 64.200 ;
        RECT 370.800 62.200 371.600 66.200 ;
        RECT 372.400 64.800 373.200 66.400 ;
        RECT 374.200 64.200 374.800 67.600 ;
        RECT 378.000 67.200 378.800 67.600 ;
        RECT 377.400 66.200 381.000 66.600 ;
        RECT 382.000 66.200 382.600 67.600 ;
        RECT 383.600 66.800 384.400 67.700 ;
        RECT 385.200 66.200 386.000 79.800 ;
        RECT 391.000 74.400 391.800 79.800 ;
        RECT 390.000 73.600 391.800 74.400 ;
        RECT 392.400 73.600 393.200 74.400 ;
        RECT 386.800 71.600 387.600 73.200 ;
        RECT 391.000 72.400 391.800 73.600 ;
        RECT 392.600 72.400 393.200 73.600 ;
        RECT 394.800 72.400 395.600 79.800 ;
        RECT 399.200 78.400 400.800 79.800 ;
        RECT 398.000 77.600 400.800 78.400 ;
        RECT 396.200 72.400 397.000 72.600 ;
        RECT 391.000 71.800 392.000 72.400 ;
        RECT 392.600 71.800 394.000 72.400 ;
        RECT 394.800 71.800 397.000 72.400 ;
        RECT 399.200 72.400 400.800 77.600 ;
        RECT 402.800 72.400 403.600 72.600 ;
        RECT 404.400 72.400 405.200 79.800 ;
        RECT 399.200 71.800 401.200 72.400 ;
        RECT 402.800 71.800 405.200 72.400 ;
        RECT 390.000 68.800 390.800 70.400 ;
        RECT 391.400 68.400 392.000 71.800 ;
        RECT 393.200 71.600 394.000 71.800 ;
        RECT 396.400 71.200 397.000 71.800 ;
        RECT 396.400 70.600 399.800 71.200 ;
        RECT 399.000 70.400 399.800 70.600 ;
        RECT 400.600 70.400 401.200 71.800 ;
        RECT 396.800 69.800 397.600 70.000 ;
        RECT 400.600 69.800 402.000 70.400 ;
        RECT 407.600 70.300 408.400 79.800 ;
        RECT 411.800 74.400 412.600 79.800 ;
        RECT 410.800 73.600 412.600 74.400 ;
        RECT 413.200 73.600 414.000 74.400 ;
        RECT 411.800 72.400 412.600 73.600 ;
        RECT 413.400 72.400 414.000 73.600 ;
        RECT 418.200 72.400 419.000 79.800 ;
        RECT 419.600 73.600 420.400 74.400 ;
        RECT 419.800 72.400 420.400 73.600 ;
        RECT 411.800 71.800 412.800 72.400 ;
        RECT 413.400 71.800 414.800 72.400 ;
        RECT 396.800 69.200 399.400 69.800 ;
        RECT 398.800 68.600 399.400 69.200 ;
        RECT 400.200 69.600 402.000 69.800 ;
        RECT 404.500 69.700 408.400 70.300 ;
        RECT 400.200 69.200 401.200 69.600 ;
        RECT 388.400 68.200 389.200 68.400 ;
        RECT 388.400 67.600 390.000 68.200 ;
        RECT 391.400 67.600 394.000 68.400 ;
        RECT 394.800 68.200 396.400 68.400 ;
        RECT 394.800 67.600 398.200 68.200 ;
        RECT 398.800 67.800 399.600 68.600 ;
        RECT 389.200 67.200 390.000 67.600 ;
        RECT 388.600 66.200 392.200 66.600 ;
        RECT 393.200 66.200 393.800 67.600 ;
        RECT 397.600 67.200 398.200 67.600 ;
        RECT 396.200 66.800 397.000 67.000 ;
        RECT 394.800 66.200 397.000 66.800 ;
        RECT 397.600 66.600 399.600 67.200 ;
        RECT 398.000 66.400 399.600 66.600 ;
        RECT 374.000 62.200 374.800 64.200 ;
        RECT 377.200 66.000 381.200 66.200 ;
        RECT 377.200 62.200 378.000 66.000 ;
        RECT 380.400 62.200 381.200 66.000 ;
        RECT 382.000 62.200 382.800 66.200 ;
        RECT 385.200 65.600 387.000 66.200 ;
        RECT 386.200 64.400 387.000 65.600 ;
        RECT 385.200 63.600 387.000 64.400 ;
        RECT 386.200 62.200 387.000 63.600 ;
        RECT 388.400 66.000 392.400 66.200 ;
        RECT 388.400 62.200 389.200 66.000 ;
        RECT 391.600 62.200 392.400 66.000 ;
        RECT 393.200 62.200 394.000 66.200 ;
        RECT 394.800 62.200 395.600 66.200 ;
        RECT 400.200 65.800 400.800 69.200 ;
        RECT 404.500 68.400 405.100 69.700 ;
        RECT 401.600 67.600 402.400 68.400 ;
        RECT 403.600 67.600 405.200 68.400 ;
        RECT 401.600 67.200 402.200 67.600 ;
        RECT 401.400 66.400 402.200 67.200 ;
        RECT 402.800 66.800 403.600 67.000 ;
        RECT 406.000 66.800 406.800 68.400 ;
        RECT 402.800 66.200 405.200 66.800 ;
        RECT 399.200 62.200 400.800 65.800 ;
        RECT 404.400 62.200 405.200 66.200 ;
        RECT 407.600 62.200 408.400 69.700 ;
        RECT 410.800 68.800 411.600 70.400 ;
        RECT 412.200 68.400 412.800 71.800 ;
        RECT 414.000 71.600 414.800 71.800 ;
        RECT 417.200 71.600 419.200 72.400 ;
        RECT 419.800 71.800 421.200 72.400 ;
        RECT 420.400 71.600 421.200 71.800 ;
        RECT 422.000 71.600 422.800 73.200 ;
        RECT 417.200 68.800 418.000 70.400 ;
        RECT 418.600 68.400 419.200 71.600 ;
        RECT 409.200 68.200 410.000 68.400 ;
        RECT 409.200 67.600 410.800 68.200 ;
        RECT 412.200 67.600 414.800 68.400 ;
        RECT 415.600 68.200 416.400 68.400 ;
        RECT 415.600 67.600 417.200 68.200 ;
        RECT 418.600 67.600 421.200 68.400 ;
        RECT 410.000 67.200 410.800 67.600 ;
        RECT 409.400 66.200 413.000 66.600 ;
        RECT 414.000 66.200 414.600 67.600 ;
        RECT 416.400 67.200 417.200 67.600 ;
        RECT 415.800 66.200 419.400 66.600 ;
        RECT 420.400 66.200 421.000 67.600 ;
        RECT 423.600 66.200 424.400 79.800 ;
        RECT 428.400 75.800 429.200 79.800 ;
        RECT 428.600 75.600 429.200 75.800 ;
        RECT 431.600 75.800 432.400 79.800 ;
        RECT 431.600 75.600 432.200 75.800 ;
        RECT 428.600 75.000 432.200 75.600 ;
        RECT 425.200 74.300 426.000 74.400 ;
        RECT 430.000 74.300 430.800 74.400 ;
        RECT 425.200 73.700 430.800 74.300 ;
        RECT 425.200 73.600 426.000 73.700 ;
        RECT 426.800 70.800 427.600 72.400 ;
        RECT 430.000 71.600 430.800 73.700 ;
        RECT 431.600 72.400 432.200 75.000 ;
        RECT 434.800 72.800 435.600 79.800 ;
        RECT 431.600 71.600 432.400 72.400 ;
        RECT 434.600 71.800 435.600 72.800 ;
        RECT 438.000 72.400 438.800 79.800 ;
        RECT 442.200 78.400 443.000 79.800 ;
        RECT 441.200 77.600 443.000 78.400 ;
        RECT 436.200 71.800 438.800 72.400 ;
        RECT 442.200 72.400 443.000 77.600 ;
        RECT 443.600 73.600 444.400 74.400 ;
        RECT 443.800 72.400 444.400 73.600 ;
        RECT 446.800 73.600 447.600 74.400 ;
        RECT 446.800 72.400 447.400 73.600 ;
        RECT 448.200 72.400 449.000 79.800 ;
        RECT 454.600 76.400 455.400 79.800 ;
        RECT 454.600 75.600 456.400 76.400 ;
        RECT 453.200 73.600 454.000 74.400 ;
        RECT 453.200 72.400 453.800 73.600 ;
        RECT 454.600 72.400 455.400 75.600 ;
        RECT 442.200 71.800 443.200 72.400 ;
        RECT 443.800 71.800 445.200 72.400 ;
        RECT 428.400 69.600 430.000 70.400 ;
        RECT 431.600 68.400 432.200 71.600 ;
        RECT 425.200 66.800 426.000 68.400 ;
        RECT 430.600 68.200 432.200 68.400 ;
        RECT 430.400 67.800 432.200 68.200 ;
        RECT 434.600 68.400 435.200 71.800 ;
        RECT 436.200 69.800 436.800 71.800 ;
        RECT 435.800 69.000 436.800 69.800 ;
        RECT 409.200 66.000 413.200 66.200 ;
        RECT 409.200 62.200 410.000 66.000 ;
        RECT 412.400 62.200 413.200 66.000 ;
        RECT 414.000 62.200 414.800 66.200 ;
        RECT 415.600 66.000 419.600 66.200 ;
        RECT 415.600 62.200 416.400 66.000 ;
        RECT 418.800 62.200 419.600 66.000 ;
        RECT 420.400 62.200 421.200 66.200 ;
        RECT 422.600 65.600 424.400 66.200 ;
        RECT 422.600 64.400 423.400 65.600 ;
        RECT 422.600 63.600 424.400 64.400 ;
        RECT 422.600 62.200 423.400 63.600 ;
        RECT 430.400 62.200 431.200 67.800 ;
        RECT 434.600 67.600 435.600 68.400 ;
        RECT 434.600 66.200 435.200 67.600 ;
        RECT 436.200 67.400 436.800 69.000 ;
        RECT 437.800 69.600 438.800 70.400 ;
        RECT 437.800 68.800 438.600 69.600 ;
        RECT 441.200 68.800 442.000 70.400 ;
        RECT 442.600 68.400 443.200 71.800 ;
        RECT 444.400 71.600 445.200 71.800 ;
        RECT 446.000 71.800 447.400 72.400 ;
        RECT 448.000 71.800 449.000 72.400 ;
        RECT 452.400 71.800 453.800 72.400 ;
        RECT 454.400 71.800 455.400 72.400 ;
        RECT 446.000 71.600 446.800 71.800 ;
        RECT 444.400 70.300 445.200 70.400 ;
        RECT 448.000 70.300 448.600 71.800 ;
        RECT 452.400 71.600 453.200 71.800 ;
        RECT 444.400 69.700 448.600 70.300 ;
        RECT 444.400 69.600 445.200 69.700 ;
        RECT 448.000 68.400 448.600 69.700 ;
        RECT 449.200 68.800 450.000 70.400 ;
        RECT 454.400 68.400 455.000 71.800 ;
        RECT 463.600 71.200 464.400 79.800 ;
        RECT 467.800 75.800 469.000 79.800 ;
        RECT 472.400 75.800 473.200 79.800 ;
        RECT 476.800 76.400 477.600 79.800 ;
        RECT 476.800 75.800 478.800 76.400 ;
        RECT 468.400 75.000 469.200 75.800 ;
        RECT 472.600 75.200 473.200 75.800 ;
        RECT 471.800 74.600 475.400 75.200 ;
        RECT 478.000 75.000 478.800 75.800 ;
        RECT 471.800 74.400 472.600 74.600 ;
        RECT 474.600 74.400 475.400 74.600 ;
        RECT 467.600 73.200 469.000 74.000 ;
        RECT 468.400 72.200 469.000 73.200 ;
        RECT 470.600 73.000 472.800 73.600 ;
        RECT 470.600 72.800 471.400 73.000 ;
        RECT 468.400 71.600 470.800 72.200 ;
        RECT 463.600 70.600 467.800 71.200 ;
        RECT 455.600 70.300 456.400 70.400 ;
        RECT 457.200 70.300 458.000 70.400 ;
        RECT 455.600 69.700 458.000 70.300 ;
        RECT 455.600 68.800 456.400 69.700 ;
        RECT 457.200 69.600 458.000 69.700 ;
        RECT 439.600 68.200 440.400 68.400 ;
        RECT 439.600 67.600 441.200 68.200 ;
        RECT 442.600 67.600 445.200 68.400 ;
        RECT 446.000 67.600 448.600 68.400 ;
        RECT 450.800 68.200 451.600 68.400 ;
        RECT 450.000 67.600 451.600 68.200 ;
        RECT 452.400 67.600 455.000 68.400 ;
        RECT 457.200 68.300 458.000 68.400 ;
        RECT 458.800 68.300 459.600 68.400 ;
        RECT 457.200 68.200 459.600 68.300 ;
        RECT 456.400 67.700 459.600 68.200 ;
        RECT 456.400 67.600 458.000 67.700 ;
        RECT 458.800 67.600 459.600 67.700 ;
        RECT 436.200 66.800 438.800 67.400 ;
        RECT 440.400 67.200 441.200 67.600 ;
        RECT 434.600 65.600 435.600 66.200 ;
        RECT 434.800 62.200 435.600 65.600 ;
        RECT 438.000 62.200 438.800 66.800 ;
        RECT 439.800 66.200 443.400 66.600 ;
        RECT 444.400 66.200 445.000 67.600 ;
        RECT 446.200 66.200 446.800 67.600 ;
        RECT 450.000 67.200 450.800 67.600 ;
        RECT 447.800 66.200 451.400 66.600 ;
        RECT 452.600 66.200 453.200 67.600 ;
        RECT 456.400 67.200 457.200 67.600 ;
        RECT 463.600 67.200 464.400 70.600 ;
        RECT 467.000 70.400 467.800 70.600 ;
        RECT 465.400 69.800 466.200 70.000 ;
        RECT 465.400 69.200 469.200 69.800 ;
        RECT 468.400 69.000 469.200 69.200 ;
        RECT 470.200 68.400 470.800 71.600 ;
        RECT 472.200 71.800 472.800 73.000 ;
        RECT 473.400 73.000 474.200 73.200 ;
        RECT 478.000 73.000 478.800 73.200 ;
        RECT 473.400 72.400 478.800 73.000 ;
        RECT 472.200 71.400 477.000 71.800 ;
        RECT 481.200 71.400 482.000 79.800 ;
        RECT 485.400 72.400 486.200 79.800 ;
        RECT 486.800 73.600 487.600 74.400 ;
        RECT 487.000 72.400 487.600 73.600 ;
        RECT 490.000 73.600 490.800 74.400 ;
        RECT 490.000 72.400 490.600 73.600 ;
        RECT 491.400 72.400 492.200 79.800 ;
        RECT 485.400 71.800 486.400 72.400 ;
        RECT 487.000 71.800 488.400 72.400 ;
        RECT 472.200 71.200 482.000 71.400 ;
        RECT 476.200 71.000 482.000 71.200 ;
        RECT 476.400 70.800 482.000 71.000 ;
        RECT 474.800 70.200 475.600 70.400 ;
        RECT 474.800 69.600 479.800 70.200 ;
        RECT 479.000 69.400 479.800 69.600 ;
        RECT 484.400 68.800 485.200 70.400 ;
        RECT 477.400 68.400 478.200 68.600 ;
        RECT 485.800 68.400 486.400 71.800 ;
        RECT 487.600 71.600 488.400 71.800 ;
        RECT 489.200 71.800 490.600 72.400 ;
        RECT 491.200 71.800 492.200 72.400 ;
        RECT 498.200 72.400 499.000 79.800 ;
        RECT 499.600 73.600 500.400 74.400 ;
        RECT 499.800 72.400 500.400 73.600 ;
        RECT 502.800 73.600 503.600 74.400 ;
        RECT 502.800 72.400 503.400 73.600 ;
        RECT 504.200 72.400 505.000 79.800 ;
        RECT 511.000 72.400 511.800 79.800 ;
        RECT 512.400 73.600 513.200 74.400 ;
        RECT 512.600 72.400 513.200 73.600 ;
        RECT 498.200 71.800 499.200 72.400 ;
        RECT 499.800 71.800 501.200 72.400 ;
        RECT 489.200 71.600 490.000 71.800 ;
        RECT 487.700 70.300 488.300 71.600 ;
        RECT 491.200 70.300 491.800 71.800 ;
        RECT 487.700 69.700 491.800 70.300 ;
        RECT 491.200 68.400 491.800 69.700 ;
        RECT 492.400 70.300 493.200 70.400 ;
        RECT 497.200 70.300 498.000 70.400 ;
        RECT 492.400 69.700 498.000 70.300 ;
        RECT 492.400 68.800 493.200 69.700 ;
        RECT 497.200 68.800 498.000 69.700 ;
        RECT 498.600 70.300 499.200 71.800 ;
        RECT 500.400 71.600 501.200 71.800 ;
        RECT 502.000 71.800 503.400 72.400 ;
        RECT 502.000 71.600 502.800 71.800 ;
        RECT 504.000 71.600 506.000 72.400 ;
        RECT 511.000 71.800 512.000 72.400 ;
        RECT 512.600 71.800 514.000 72.400 ;
        RECT 502.100 70.300 502.700 71.600 ;
        RECT 498.600 69.700 502.700 70.300 ;
        RECT 498.600 68.400 499.200 69.700 ;
        RECT 504.000 68.400 504.600 71.600 ;
        RECT 505.200 68.800 506.000 70.400 ;
        RECT 508.400 70.300 509.200 70.400 ;
        RECT 510.000 70.300 510.800 70.400 ;
        RECT 508.400 69.700 510.800 70.300 ;
        RECT 508.400 69.600 509.200 69.700 ;
        RECT 510.000 68.800 510.800 69.700 ;
        RECT 511.400 68.400 512.000 71.800 ;
        RECT 513.200 71.600 514.000 71.800 ;
        RECT 514.800 71.200 515.600 79.800 ;
        RECT 519.000 75.800 520.200 79.800 ;
        RECT 523.600 75.800 524.400 79.800 ;
        RECT 528.000 76.400 528.800 79.800 ;
        RECT 528.000 75.800 530.000 76.400 ;
        RECT 519.600 75.000 520.400 75.800 ;
        RECT 523.800 75.200 524.400 75.800 ;
        RECT 523.000 74.600 526.600 75.200 ;
        RECT 529.200 75.000 530.000 75.800 ;
        RECT 523.000 74.400 523.800 74.600 ;
        RECT 525.800 74.400 526.600 74.600 ;
        RECT 518.800 73.200 520.200 74.000 ;
        RECT 519.600 72.200 520.200 73.200 ;
        RECT 521.800 73.000 524.000 73.600 ;
        RECT 521.800 72.800 522.600 73.000 ;
        RECT 519.600 71.600 522.000 72.200 ;
        RECT 514.800 70.600 519.000 71.200 ;
        RECT 470.200 67.800 481.200 68.400 ;
        RECT 470.600 67.600 471.400 67.800 ;
        RECT 473.200 67.600 474.000 67.800 ;
        RECT 463.600 66.600 467.400 67.200 ;
        RECT 454.200 66.200 457.800 66.600 ;
        RECT 439.600 66.000 443.600 66.200 ;
        RECT 439.600 62.200 440.400 66.000 ;
        RECT 442.800 62.200 443.600 66.000 ;
        RECT 444.400 62.200 445.200 66.200 ;
        RECT 446.000 62.200 446.800 66.200 ;
        RECT 447.600 66.000 451.600 66.200 ;
        RECT 447.600 62.200 448.400 66.000 ;
        RECT 450.800 62.200 451.600 66.000 ;
        RECT 452.400 62.200 453.200 66.200 ;
        RECT 454.000 66.000 458.000 66.200 ;
        RECT 454.000 62.200 454.800 66.000 ;
        RECT 457.200 62.200 458.000 66.000 ;
        RECT 463.600 62.200 464.400 66.600 ;
        RECT 466.600 66.400 467.400 66.600 ;
        RECT 476.400 65.600 477.000 67.800 ;
        RECT 479.600 67.600 481.200 67.800 ;
        RECT 482.800 68.200 483.600 68.400 ;
        RECT 482.800 67.600 484.400 68.200 ;
        RECT 485.800 67.600 488.400 68.400 ;
        RECT 489.200 67.600 491.800 68.400 ;
        RECT 494.000 68.300 494.800 68.400 ;
        RECT 495.600 68.300 496.400 68.400 ;
        RECT 494.000 68.200 496.400 68.300 ;
        RECT 493.200 67.700 497.200 68.200 ;
        RECT 493.200 67.600 494.800 67.700 ;
        RECT 495.600 67.600 497.200 67.700 ;
        RECT 498.600 67.600 501.200 68.400 ;
        RECT 502.000 67.600 504.600 68.400 ;
        RECT 506.800 68.200 507.600 68.400 ;
        RECT 506.000 67.600 507.600 68.200 ;
        RECT 508.400 68.200 509.200 68.400 ;
        RECT 508.400 67.600 510.000 68.200 ;
        RECT 511.400 67.600 514.000 68.400 ;
        RECT 483.600 67.200 484.400 67.600 ;
        RECT 474.600 65.400 475.400 65.600 ;
        RECT 468.400 64.200 469.200 65.000 ;
        RECT 472.600 64.800 475.400 65.400 ;
        RECT 476.400 64.800 477.200 65.600 ;
        RECT 472.600 64.200 473.200 64.800 ;
        RECT 478.000 64.200 478.800 65.000 ;
        RECT 467.800 63.600 469.200 64.200 ;
        RECT 467.800 62.200 469.000 63.600 ;
        RECT 472.400 62.200 473.200 64.200 ;
        RECT 476.800 63.600 478.800 64.200 ;
        RECT 476.800 62.200 477.600 63.600 ;
        RECT 481.200 62.200 482.000 67.000 ;
        RECT 483.000 66.200 486.600 66.600 ;
        RECT 487.600 66.200 488.200 67.600 ;
        RECT 489.400 66.200 490.000 67.600 ;
        RECT 493.200 67.200 494.000 67.600 ;
        RECT 496.400 67.200 497.200 67.600 ;
        RECT 491.000 66.200 494.600 66.600 ;
        RECT 495.800 66.200 499.400 66.600 ;
        RECT 500.400 66.200 501.000 67.600 ;
        RECT 502.200 66.200 502.800 67.600 ;
        RECT 506.000 67.200 506.800 67.600 ;
        RECT 509.200 67.200 510.000 67.600 ;
        RECT 503.800 66.200 507.400 66.600 ;
        RECT 508.600 66.200 512.200 66.600 ;
        RECT 513.200 66.200 513.800 67.600 ;
        RECT 514.800 67.200 515.600 70.600 ;
        RECT 518.200 70.400 519.000 70.600 ;
        RECT 516.600 69.800 517.400 70.000 ;
        RECT 516.600 69.200 520.400 69.800 ;
        RECT 519.600 69.000 520.400 69.200 ;
        RECT 521.400 68.400 522.000 71.600 ;
        RECT 523.400 71.800 524.000 73.000 ;
        RECT 524.600 73.000 525.400 73.200 ;
        RECT 529.200 73.000 530.000 73.200 ;
        RECT 524.600 72.400 530.000 73.000 ;
        RECT 523.400 71.400 528.200 71.800 ;
        RECT 532.400 71.400 533.200 79.800 ;
        RECT 536.600 74.400 537.400 79.800 ;
        RECT 535.600 73.600 537.400 74.400 ;
        RECT 538.000 73.600 538.800 74.400 ;
        RECT 536.600 72.400 537.400 73.600 ;
        RECT 538.200 72.400 538.800 73.600 ;
        RECT 536.600 71.800 537.600 72.400 ;
        RECT 538.200 72.300 539.600 72.400 ;
        RECT 542.000 72.300 542.800 79.800 ;
        RECT 538.200 71.800 542.800 72.300 ;
        RECT 523.400 71.200 533.200 71.400 ;
        RECT 527.400 71.000 533.200 71.200 ;
        RECT 527.600 70.800 533.200 71.000 ;
        RECT 526.000 70.200 526.800 70.400 ;
        RECT 526.000 69.600 531.000 70.200 ;
        RECT 530.200 69.400 531.000 69.600 ;
        RECT 535.600 68.800 536.400 70.400 ;
        RECT 528.600 68.400 529.400 68.600 ;
        RECT 537.000 68.400 537.600 71.800 ;
        RECT 538.800 71.700 542.800 71.800 ;
        RECT 538.800 71.600 539.600 71.700 ;
        RECT 521.400 67.800 532.400 68.400 ;
        RECT 521.800 67.600 522.600 67.800 ;
        RECT 526.000 67.600 526.800 67.800 ;
        RECT 514.800 66.600 518.600 67.200 ;
        RECT 482.800 66.000 486.800 66.200 ;
        RECT 482.800 62.200 483.600 66.000 ;
        RECT 486.000 62.200 486.800 66.000 ;
        RECT 487.600 62.200 488.400 66.200 ;
        RECT 489.200 62.200 490.000 66.200 ;
        RECT 490.800 66.000 494.800 66.200 ;
        RECT 490.800 62.200 491.600 66.000 ;
        RECT 494.000 62.200 494.800 66.000 ;
        RECT 495.600 66.000 499.600 66.200 ;
        RECT 495.600 62.200 496.400 66.000 ;
        RECT 498.800 62.200 499.600 66.000 ;
        RECT 500.400 62.200 501.200 66.200 ;
        RECT 502.000 62.200 502.800 66.200 ;
        RECT 503.600 66.000 507.600 66.200 ;
        RECT 503.600 62.200 504.400 66.000 ;
        RECT 506.800 62.200 507.600 66.000 ;
        RECT 508.400 66.000 512.400 66.200 ;
        RECT 508.400 62.200 509.200 66.000 ;
        RECT 511.600 62.200 512.400 66.000 ;
        RECT 513.200 62.200 514.000 66.200 ;
        RECT 514.800 62.200 515.600 66.600 ;
        RECT 517.800 66.400 518.600 66.600 ;
        RECT 527.600 65.600 528.200 67.800 ;
        RECT 530.800 67.600 532.400 67.800 ;
        RECT 534.000 68.200 534.800 68.400 ;
        RECT 534.000 67.600 535.600 68.200 ;
        RECT 537.000 67.600 539.600 68.400 ;
        RECT 534.800 67.200 535.600 67.600 ;
        RECT 525.800 65.400 526.600 65.600 ;
        RECT 519.600 64.200 520.400 65.000 ;
        RECT 523.800 64.800 526.600 65.400 ;
        RECT 527.600 64.800 528.400 65.600 ;
        RECT 523.800 64.200 524.400 64.800 ;
        RECT 529.200 64.200 530.000 65.000 ;
        RECT 519.000 63.600 520.400 64.200 ;
        RECT 519.000 62.200 520.200 63.600 ;
        RECT 523.600 62.200 524.400 64.200 ;
        RECT 528.000 63.600 530.000 64.200 ;
        RECT 528.000 62.200 528.800 63.600 ;
        RECT 532.400 62.200 533.200 67.000 ;
        RECT 534.200 66.200 537.800 66.600 ;
        RECT 538.800 66.200 539.400 67.600 ;
        RECT 540.400 66.800 541.200 68.400 ;
        RECT 542.000 66.200 542.800 71.700 ;
        RECT 543.600 72.300 544.400 73.200 ;
        RECT 545.200 72.300 546.000 73.200 ;
        RECT 543.600 71.700 546.000 72.300 ;
        RECT 543.600 71.600 544.400 71.700 ;
        RECT 545.200 71.600 546.000 71.700 ;
        RECT 546.800 66.400 547.600 79.800 ;
        RECT 550.000 72.400 550.800 79.800 ;
        RECT 553.200 72.800 554.000 79.800 ;
        RECT 559.000 74.400 559.800 79.800 ;
        RECT 562.800 75.000 563.600 79.000 ;
        RECT 558.000 73.600 559.800 74.400 ;
        RECT 560.400 73.600 561.200 74.400 ;
        RECT 550.000 71.800 552.600 72.400 ;
        RECT 553.200 71.800 554.200 72.800 ;
        RECT 559.000 72.400 559.800 73.600 ;
        RECT 560.600 72.400 561.200 73.600 ;
        RECT 559.000 71.800 560.000 72.400 ;
        RECT 560.600 71.800 562.000 72.400 ;
        RECT 548.400 70.300 549.200 70.400 ;
        RECT 550.000 70.300 551.000 70.400 ;
        RECT 548.400 69.700 551.000 70.300 ;
        RECT 548.400 69.600 549.200 69.700 ;
        RECT 550.000 69.600 551.000 69.700 ;
        RECT 550.200 68.800 551.000 69.600 ;
        RECT 552.000 69.800 552.600 71.800 ;
        RECT 552.000 69.000 553.000 69.800 ;
        RECT 548.400 66.800 549.200 68.400 ;
        RECT 552.000 67.400 552.600 69.000 ;
        RECT 553.600 68.400 554.200 71.800 ;
        RECT 554.800 70.300 555.600 70.400 ;
        RECT 558.000 70.300 558.800 70.400 ;
        RECT 554.800 69.700 558.800 70.300 ;
        RECT 554.800 69.600 555.600 69.700 ;
        RECT 558.000 68.800 558.800 69.700 ;
        RECT 559.400 68.400 560.000 71.800 ;
        RECT 561.200 71.600 562.000 71.800 ;
        RECT 562.800 71.600 563.400 75.000 ;
        RECT 567.000 72.800 567.800 79.800 ;
        RECT 574.600 74.400 575.400 79.800 ;
        RECT 573.200 73.600 574.000 74.400 ;
        RECT 574.600 73.600 576.400 74.400 ;
        RECT 567.000 72.200 568.600 72.800 ;
        RECT 573.200 72.400 573.800 73.600 ;
        RECT 574.600 72.400 575.400 73.600 ;
        RECT 562.800 71.000 566.600 71.600 ;
        RECT 561.200 70.300 562.000 70.400 ;
        RECT 562.800 70.300 563.600 70.400 ;
        RECT 561.200 69.700 563.600 70.300 ;
        RECT 561.200 69.600 562.000 69.700 ;
        RECT 562.800 68.800 563.600 69.700 ;
        RECT 564.400 68.800 565.200 70.400 ;
        RECT 566.000 69.000 566.600 71.000 ;
        RECT 553.200 67.600 554.200 68.400 ;
        RECT 556.400 68.200 557.200 68.400 ;
        RECT 556.400 67.600 558.000 68.200 ;
        RECT 559.400 67.600 562.000 68.400 ;
        RECT 566.000 68.200 567.400 69.000 ;
        RECT 568.000 68.400 568.600 72.200 ;
        RECT 572.400 71.800 573.800 72.400 ;
        RECT 574.400 71.800 575.400 72.400 ;
        RECT 572.400 71.600 573.200 71.800 ;
        RECT 569.200 69.600 570.000 71.200 ;
        RECT 574.400 68.400 575.000 71.800 ;
        RECT 578.800 71.400 579.600 79.800 ;
        RECT 583.200 76.400 584.000 79.800 ;
        RECT 582.000 75.800 584.000 76.400 ;
        RECT 587.600 75.800 588.400 79.800 ;
        RECT 591.800 75.800 593.000 79.800 ;
        RECT 582.000 75.000 582.800 75.800 ;
        RECT 587.600 75.200 588.200 75.800 ;
        RECT 585.400 74.600 589.000 75.200 ;
        RECT 591.600 75.000 592.400 75.800 ;
        RECT 585.400 74.400 586.200 74.600 ;
        RECT 588.200 74.400 589.000 74.600 ;
        RECT 582.000 73.000 582.800 73.200 ;
        RECT 586.600 73.000 587.400 73.200 ;
        RECT 582.000 72.400 587.400 73.000 ;
        RECT 588.000 73.000 590.200 73.600 ;
        RECT 588.000 71.800 588.600 73.000 ;
        RECT 589.400 72.800 590.200 73.000 ;
        RECT 591.800 73.200 593.200 74.000 ;
        RECT 591.800 72.200 592.400 73.200 ;
        RECT 583.800 71.400 588.600 71.800 ;
        RECT 578.800 71.200 588.600 71.400 ;
        RECT 590.000 71.600 592.400 72.200 ;
        RECT 578.800 71.000 584.600 71.200 ;
        RECT 578.800 70.800 584.400 71.000 ;
        RECT 575.600 68.800 576.400 70.400 ;
        RECT 585.200 70.200 586.000 70.400 ;
        RECT 581.000 69.600 586.000 70.200 ;
        RECT 581.000 69.400 581.800 69.600 ;
        RECT 583.600 69.400 584.400 69.600 ;
        RECT 582.600 68.400 583.400 68.600 ;
        RECT 590.000 68.400 590.600 71.600 ;
        RECT 596.400 71.200 597.200 79.800 ;
        RECT 593.000 70.600 597.200 71.200 ;
        RECT 593.000 70.400 593.800 70.600 ;
        RECT 594.600 69.800 595.400 70.000 ;
        RECT 591.600 69.200 595.400 69.800 ;
        RECT 591.600 69.000 592.400 69.200 ;
        RECT 568.000 68.300 570.000 68.400 ;
        RECT 570.800 68.300 571.600 68.400 ;
        RECT 566.000 67.800 567.000 68.200 ;
        RECT 550.000 66.800 552.600 67.400 ;
        RECT 534.000 66.000 538.000 66.200 ;
        RECT 534.000 62.200 534.800 66.000 ;
        RECT 537.200 62.200 538.000 66.000 ;
        RECT 538.800 62.200 539.600 66.200 ;
        RECT 542.000 65.600 543.800 66.200 ;
        RECT 545.200 65.600 547.600 66.400 ;
        RECT 543.000 62.200 543.800 65.600 ;
        RECT 545.800 62.200 546.600 65.600 ;
        RECT 550.000 62.200 550.800 66.800 ;
        RECT 553.600 66.200 554.200 67.600 ;
        RECT 557.200 67.200 558.000 67.600 ;
        RECT 556.600 66.200 560.200 66.600 ;
        RECT 561.200 66.200 561.800 67.600 ;
        RECT 562.800 67.200 567.000 67.800 ;
        RECT 568.000 67.700 571.600 68.300 ;
        RECT 568.000 67.600 570.000 67.700 ;
        RECT 570.800 67.600 571.600 67.700 ;
        RECT 572.400 67.600 575.000 68.400 ;
        RECT 577.200 68.200 578.000 68.400 ;
        RECT 576.400 67.600 578.000 68.200 ;
        RECT 579.600 67.800 590.600 68.400 ;
        RECT 579.600 67.600 581.200 67.800 ;
        RECT 553.200 65.600 554.200 66.200 ;
        RECT 556.400 66.000 560.400 66.200 ;
        RECT 553.200 62.200 554.000 65.600 ;
        RECT 556.400 62.200 557.200 66.000 ;
        RECT 559.600 62.200 560.400 66.000 ;
        RECT 561.200 62.200 562.000 66.200 ;
        RECT 562.800 65.000 563.400 67.200 ;
        RECT 568.000 67.000 568.600 67.600 ;
        RECT 567.800 66.600 568.600 67.000 ;
        RECT 567.000 66.000 568.600 66.600 ;
        RECT 572.600 66.200 573.200 67.600 ;
        RECT 576.400 67.200 577.200 67.600 ;
        RECT 574.200 66.200 577.800 66.600 ;
        RECT 562.800 63.000 563.600 65.000 ;
        RECT 567.000 63.000 567.800 66.000 ;
        RECT 572.400 62.200 573.200 66.200 ;
        RECT 574.000 66.000 578.000 66.200 ;
        RECT 574.000 62.200 574.800 66.000 ;
        RECT 577.200 62.200 578.000 66.000 ;
        RECT 578.800 62.200 579.600 67.000 ;
        RECT 583.800 65.600 584.400 67.800 ;
        RECT 589.400 67.600 590.200 67.800 ;
        RECT 596.400 67.200 597.200 70.600 ;
        RECT 593.400 66.600 597.200 67.200 ;
        RECT 598.000 66.800 598.800 68.400 ;
        RECT 593.400 66.400 594.200 66.600 ;
        RECT 582.000 64.200 582.800 65.000 ;
        RECT 583.600 64.800 584.400 65.600 ;
        RECT 585.400 65.400 586.200 65.600 ;
        RECT 585.400 64.800 588.200 65.400 ;
        RECT 587.600 64.200 588.200 64.800 ;
        RECT 591.600 64.200 592.400 65.000 ;
        RECT 582.000 63.600 584.000 64.200 ;
        RECT 583.200 62.200 584.000 63.600 ;
        RECT 587.600 62.200 588.400 64.200 ;
        RECT 591.600 63.600 593.000 64.200 ;
        RECT 591.800 62.200 593.000 63.600 ;
        RECT 596.400 62.200 597.200 66.600 ;
        RECT 599.600 66.200 600.400 79.800 ;
        RECT 603.600 73.600 604.400 74.400 ;
        RECT 601.200 71.600 602.000 73.200 ;
        RECT 603.600 72.400 604.200 73.600 ;
        RECT 605.000 72.400 605.800 79.800 ;
        RECT 602.800 71.800 604.200 72.400 ;
        RECT 604.800 71.800 605.800 72.400 ;
        RECT 602.800 71.600 603.600 71.800 ;
        RECT 604.800 68.400 605.400 71.800 ;
        RECT 606.000 68.800 606.800 70.400 ;
        RECT 602.800 67.600 605.400 68.400 ;
        RECT 607.600 68.200 608.400 68.400 ;
        RECT 606.800 67.600 608.400 68.200 ;
        RECT 603.000 66.200 603.600 67.600 ;
        RECT 606.800 67.200 607.600 67.600 ;
        RECT 604.600 66.200 608.200 66.600 ;
        RECT 599.600 65.600 601.400 66.200 ;
        RECT 600.600 62.200 601.400 65.600 ;
        RECT 602.800 62.200 603.600 66.200 ;
        RECT 604.400 66.000 608.400 66.200 ;
        RECT 604.400 62.200 605.200 66.000 ;
        RECT 607.600 62.200 608.400 66.000 ;
        RECT 1.200 53.800 2.000 59.800 ;
        RECT 7.600 56.600 8.400 59.800 ;
        RECT 9.200 57.000 10.000 59.800 ;
        RECT 10.800 57.000 11.600 59.800 ;
        RECT 12.400 57.000 13.200 59.800 ;
        RECT 15.600 57.000 16.400 59.800 ;
        RECT 18.800 57.000 19.600 59.800 ;
        RECT 20.400 57.000 21.200 59.800 ;
        RECT 22.000 57.000 22.800 59.800 ;
        RECT 23.600 57.000 24.400 59.800 ;
        RECT 5.800 55.800 8.400 56.600 ;
        RECT 25.200 56.600 26.000 59.800 ;
        RECT 11.800 55.800 16.400 56.400 ;
        RECT 5.800 55.200 6.600 55.800 ;
        RECT 3.600 54.400 6.600 55.200 ;
        RECT 1.200 53.000 10.000 53.800 ;
        RECT 11.800 53.400 12.600 55.800 ;
        RECT 15.600 55.600 16.400 55.800 ;
        RECT 17.200 55.600 18.800 56.400 ;
        RECT 21.800 55.600 22.800 56.400 ;
        RECT 25.200 55.800 27.600 56.600 ;
        RECT 14.000 53.600 14.800 55.200 ;
        RECT 15.600 54.800 16.400 55.000 ;
        RECT 15.600 54.200 20.000 54.800 ;
        RECT 19.200 54.000 20.000 54.200 ;
        RECT 1.200 47.400 2.000 53.000 ;
        RECT 10.600 52.600 12.600 53.400 ;
        RECT 16.400 52.600 19.600 53.400 ;
        RECT 22.000 52.800 22.800 55.600 ;
        RECT 26.800 55.200 27.600 55.800 ;
        RECT 26.800 54.600 28.600 55.200 ;
        RECT 27.800 53.400 28.600 54.600 ;
        RECT 31.600 54.600 32.400 59.800 ;
        RECT 33.200 56.000 34.000 59.800 ;
        RECT 36.400 56.000 37.200 59.800 ;
        RECT 39.600 56.000 40.400 59.800 ;
        RECT 33.200 55.200 34.200 56.000 ;
        RECT 36.400 55.800 40.400 56.000 ;
        RECT 41.200 55.800 42.000 59.800 ;
        RECT 43.400 58.400 44.200 59.800 ;
        RECT 43.400 57.600 45.200 58.400 ;
        RECT 43.400 56.400 44.200 57.600 ;
        RECT 43.400 55.800 45.200 56.400 ;
        RECT 36.600 55.400 40.200 55.800 ;
        RECT 31.600 54.000 32.800 54.600 ;
        RECT 27.800 52.600 31.600 53.400 ;
        RECT 2.600 52.000 3.400 52.200 ;
        RECT 7.600 52.000 8.400 52.400 ;
        RECT 25.200 52.000 26.000 52.600 ;
        RECT 32.200 52.000 32.800 54.000 ;
        RECT 2.600 51.400 26.000 52.000 ;
        RECT 32.000 51.400 32.800 52.000 ;
        RECT 32.000 49.600 32.600 51.400 ;
        RECT 33.400 50.800 34.200 55.200 ;
        RECT 37.200 54.400 38.000 54.800 ;
        RECT 41.200 54.400 41.800 55.800 ;
        RECT 36.400 53.800 38.000 54.400 ;
        RECT 36.400 53.600 37.200 53.800 ;
        RECT 39.400 53.600 42.000 54.400 ;
        RECT 34.800 52.300 35.600 52.400 ;
        RECT 38.000 52.300 38.800 53.200 ;
        RECT 34.800 51.700 38.800 52.300 ;
        RECT 34.800 51.600 35.600 51.700 ;
        RECT 38.000 51.600 38.800 51.700 ;
        RECT 10.800 49.400 11.600 49.600 ;
        RECT 6.200 49.000 11.600 49.400 ;
        RECT 5.400 48.800 11.600 49.000 ;
        RECT 12.600 49.000 21.200 49.600 ;
        RECT 2.800 48.000 4.400 48.800 ;
        RECT 5.400 48.200 6.800 48.800 ;
        RECT 12.600 48.200 13.200 49.000 ;
        RECT 20.400 48.800 21.200 49.000 ;
        RECT 23.600 49.000 32.600 49.600 ;
        RECT 23.600 48.800 24.400 49.000 ;
        RECT 3.800 47.600 4.400 48.000 ;
        RECT 7.400 47.600 13.200 48.200 ;
        RECT 13.800 47.600 16.400 48.400 ;
        RECT 1.200 46.800 3.200 47.400 ;
        RECT 3.800 46.800 8.000 47.600 ;
        RECT 2.600 46.200 3.200 46.800 ;
        RECT 2.600 45.600 3.600 46.200 ;
        RECT 2.800 42.200 3.600 45.600 ;
        RECT 6.000 42.200 6.800 46.800 ;
        RECT 9.200 42.200 10.000 45.000 ;
        RECT 10.800 42.200 11.600 45.000 ;
        RECT 12.400 42.200 13.200 47.000 ;
        RECT 15.600 42.200 16.400 47.000 ;
        RECT 18.800 42.200 19.600 48.400 ;
        RECT 26.800 47.600 29.400 48.400 ;
        RECT 22.000 46.800 26.200 47.600 ;
        RECT 20.400 42.200 21.200 45.000 ;
        RECT 22.000 42.200 22.800 45.000 ;
        RECT 23.600 42.200 24.400 45.000 ;
        RECT 26.800 42.200 27.600 47.600 ;
        RECT 32.000 47.400 32.600 49.000 ;
        RECT 30.000 46.800 32.600 47.400 ;
        RECT 33.200 50.000 34.200 50.800 ;
        RECT 39.400 50.200 40.000 53.600 ;
        RECT 41.200 50.200 42.000 50.400 ;
        RECT 30.000 42.200 30.800 46.800 ;
        RECT 33.200 42.200 34.000 50.000 ;
        RECT 39.000 49.600 40.000 50.200 ;
        RECT 40.600 49.600 42.000 50.200 ;
        RECT 39.000 44.400 39.800 49.600 ;
        RECT 40.600 48.400 41.200 49.600 ;
        RECT 40.400 47.600 41.200 48.400 ;
        RECT 42.800 47.600 43.600 50.400 ;
        RECT 38.000 43.600 39.800 44.400 ;
        RECT 39.000 42.200 39.800 43.600 ;
        RECT 44.400 42.200 45.200 55.800 ;
        RECT 49.200 55.200 50.000 59.800 ;
        RECT 52.400 55.200 53.200 59.800 ;
        RECT 55.600 55.200 56.400 59.800 ;
        RECT 58.800 55.200 59.600 59.800 ;
        RECT 65.800 56.000 66.600 59.000 ;
        RECT 70.000 57.000 70.800 59.000 ;
        RECT 46.000 53.600 46.800 55.200 ;
        RECT 47.600 54.400 50.000 55.200 ;
        RECT 51.000 54.400 53.200 55.200 ;
        RECT 54.200 54.400 56.400 55.200 ;
        RECT 57.800 54.400 59.600 55.200 ;
        RECT 65.000 55.400 66.600 56.000 ;
        RECT 65.000 55.000 65.800 55.400 ;
        RECT 65.000 54.400 65.600 55.000 ;
        RECT 70.200 54.800 70.800 57.000 ;
        RECT 72.200 58.400 73.000 59.800 ;
        RECT 72.200 57.600 74.000 58.400 ;
        RECT 72.200 56.400 73.000 57.600 ;
        RECT 76.400 57.000 77.200 59.000 ;
        RECT 72.200 55.800 74.000 56.400 ;
        RECT 47.600 51.600 48.400 54.400 ;
        RECT 51.000 53.800 51.800 54.400 ;
        RECT 54.200 53.800 55.000 54.400 ;
        RECT 57.800 53.800 58.600 54.400 ;
        RECT 60.400 53.800 61.200 54.400 ;
        RECT 49.200 53.000 51.800 53.800 ;
        RECT 52.600 53.000 55.000 53.800 ;
        RECT 56.000 53.000 58.600 53.800 ;
        RECT 59.400 53.000 61.200 53.800 ;
        RECT 63.600 53.600 65.600 54.400 ;
        RECT 66.600 54.200 70.800 54.800 ;
        RECT 66.600 53.800 67.600 54.200 ;
        RECT 51.000 51.600 51.800 53.000 ;
        RECT 54.200 51.600 55.000 53.000 ;
        RECT 57.800 51.600 58.600 53.000 ;
        RECT 47.600 50.800 50.000 51.600 ;
        RECT 51.000 50.800 53.200 51.600 ;
        RECT 54.200 50.800 56.400 51.600 ;
        RECT 57.800 50.800 59.600 51.600 ;
        RECT 63.600 50.800 64.400 52.400 ;
        RECT 49.200 42.200 50.000 50.800 ;
        RECT 52.400 42.200 53.200 50.800 ;
        RECT 55.600 42.200 56.400 50.800 ;
        RECT 58.800 42.200 59.600 50.800 ;
        RECT 65.000 49.800 65.600 53.600 ;
        RECT 66.200 53.000 67.600 53.800 ;
        RECT 67.000 51.000 67.600 53.000 ;
        RECT 68.400 51.600 69.200 53.200 ;
        RECT 70.000 52.300 70.800 53.200 ;
        RECT 71.600 52.300 72.400 52.400 ;
        RECT 70.000 51.700 72.400 52.300 ;
        RECT 70.000 51.600 70.800 51.700 ;
        RECT 71.600 51.600 72.400 51.700 ;
        RECT 67.000 50.400 70.800 51.000 ;
        RECT 65.000 49.200 66.600 49.800 ;
        RECT 65.800 44.400 66.600 49.200 ;
        RECT 70.200 47.000 70.800 50.400 ;
        RECT 71.600 48.800 72.400 50.400 ;
        RECT 65.200 43.600 66.600 44.400 ;
        RECT 65.800 42.200 66.600 43.600 ;
        RECT 70.000 43.000 70.800 47.000 ;
        RECT 73.200 42.200 74.000 55.800 ;
        RECT 74.800 53.600 75.600 55.200 ;
        RECT 76.400 54.800 77.000 57.000 ;
        RECT 80.600 56.000 81.400 59.000 ;
        RECT 89.800 56.000 90.600 59.000 ;
        RECT 94.000 57.000 94.800 59.000 ;
        RECT 80.600 55.400 82.200 56.000 ;
        RECT 81.400 55.000 82.200 55.400 ;
        RECT 76.400 54.200 80.600 54.800 ;
        RECT 79.600 53.800 80.600 54.200 ;
        RECT 81.600 54.400 82.200 55.000 ;
        RECT 89.000 55.400 90.600 56.000 ;
        RECT 89.000 55.000 89.800 55.400 ;
        RECT 89.000 54.400 89.600 55.000 ;
        RECT 94.200 54.800 94.800 57.000 ;
        RECT 95.600 55.600 96.400 57.200 ;
        RECT 76.400 51.600 77.200 53.200 ;
        RECT 78.000 51.600 78.800 53.200 ;
        RECT 79.600 53.000 81.000 53.800 ;
        RECT 81.600 53.600 83.600 54.400 ;
        RECT 87.600 53.600 89.600 54.400 ;
        RECT 90.600 54.200 94.800 54.800 ;
        RECT 90.600 53.800 91.600 54.200 ;
        RECT 79.600 51.000 80.200 53.000 ;
        RECT 76.400 50.400 80.200 51.000 ;
        RECT 76.400 47.000 77.000 50.400 ;
        RECT 81.600 49.800 82.200 53.600 ;
        RECT 82.800 52.300 83.600 52.400 ;
        RECT 86.000 52.300 86.800 52.400 ;
        RECT 82.800 51.700 86.800 52.300 ;
        RECT 82.800 50.800 83.600 51.700 ;
        RECT 86.000 51.600 86.800 51.700 ;
        RECT 87.600 50.800 88.400 52.400 ;
        RECT 80.600 49.200 82.200 49.800 ;
        RECT 89.000 49.800 89.600 53.600 ;
        RECT 90.200 53.000 91.600 53.800 ;
        RECT 91.000 51.000 91.600 53.000 ;
        RECT 92.400 51.600 93.200 53.200 ;
        RECT 94.000 51.600 94.800 53.200 ;
        RECT 91.000 50.400 94.800 51.000 ;
        RECT 89.000 49.200 90.600 49.800 ;
        RECT 76.400 43.000 77.200 47.000 ;
        RECT 80.600 44.400 81.400 49.200 ;
        RECT 79.600 43.600 81.400 44.400 ;
        RECT 80.600 42.200 81.400 43.600 ;
        RECT 89.800 44.400 90.600 49.200 ;
        RECT 94.200 47.000 94.800 50.400 ;
        RECT 89.800 43.600 91.600 44.400 ;
        RECT 89.800 42.200 90.600 43.600 ;
        RECT 94.000 43.000 94.800 47.000 ;
        RECT 97.200 42.200 98.000 59.800 ;
        RECT 100.400 55.200 101.200 59.800 ;
        RECT 103.600 55.200 104.400 59.800 ;
        RECT 106.800 55.200 107.600 59.800 ;
        RECT 110.000 55.200 110.800 59.800 ;
        RECT 117.000 56.000 117.800 59.000 ;
        RECT 121.200 57.000 122.000 59.000 ;
        RECT 98.800 54.400 101.200 55.200 ;
        RECT 102.200 54.400 104.400 55.200 ;
        RECT 105.400 54.400 107.600 55.200 ;
        RECT 109.000 54.400 110.800 55.200 ;
        RECT 116.200 55.400 117.800 56.000 ;
        RECT 116.200 55.000 117.000 55.400 ;
        RECT 116.200 54.400 116.800 55.000 ;
        RECT 121.400 54.800 122.000 57.000 ;
        RECT 98.800 51.600 99.600 54.400 ;
        RECT 102.200 53.800 103.000 54.400 ;
        RECT 105.400 53.800 106.200 54.400 ;
        RECT 109.000 53.800 109.800 54.400 ;
        RECT 111.600 53.800 112.400 54.400 ;
        RECT 100.400 53.000 103.000 53.800 ;
        RECT 103.800 53.000 106.200 53.800 ;
        RECT 107.200 53.000 109.800 53.800 ;
        RECT 110.600 53.000 112.400 53.800 ;
        RECT 114.800 53.600 116.800 54.400 ;
        RECT 117.800 54.200 122.000 54.800 ;
        RECT 122.800 57.000 123.600 59.000 ;
        RECT 122.800 54.800 123.400 57.000 ;
        RECT 127.000 56.000 127.800 59.000 ;
        RECT 134.000 56.400 134.800 59.800 ;
        RECT 127.000 55.400 128.600 56.000 ;
        RECT 127.800 55.000 128.600 55.400 ;
        RECT 122.800 54.200 127.000 54.800 ;
        RECT 117.800 53.800 118.800 54.200 ;
        RECT 102.200 51.600 103.000 53.000 ;
        RECT 105.400 51.600 106.200 53.000 ;
        RECT 109.000 51.600 109.800 53.000 ;
        RECT 113.200 52.300 114.000 52.400 ;
        RECT 114.800 52.300 115.600 52.400 ;
        RECT 113.200 51.700 115.600 52.300 ;
        RECT 113.200 51.600 114.000 51.700 ;
        RECT 98.800 50.800 101.200 51.600 ;
        RECT 102.200 50.800 104.400 51.600 ;
        RECT 105.400 50.800 107.600 51.600 ;
        RECT 109.000 50.800 110.800 51.600 ;
        RECT 114.800 50.800 115.600 51.700 ;
        RECT 100.400 42.200 101.200 50.800 ;
        RECT 103.600 42.200 104.400 50.800 ;
        RECT 106.800 42.200 107.600 50.800 ;
        RECT 110.000 42.200 110.800 50.800 ;
        RECT 116.200 49.800 116.800 53.600 ;
        RECT 117.400 53.000 118.800 53.800 ;
        RECT 126.000 53.800 127.000 54.200 ;
        RECT 128.000 54.400 128.600 55.000 ;
        RECT 133.800 55.800 134.800 56.400 ;
        RECT 133.800 54.400 134.400 55.800 ;
        RECT 137.200 55.200 138.000 59.800 ;
        RECT 142.600 56.400 143.400 59.000 ;
        RECT 146.800 57.000 147.600 59.000 ;
        RECT 142.600 56.000 144.400 56.400 ;
        RECT 135.400 54.600 138.000 55.200 ;
        RECT 141.800 55.600 144.400 56.000 ;
        RECT 141.800 55.400 143.400 55.600 ;
        RECT 141.800 55.000 142.600 55.400 ;
        RECT 118.200 51.000 118.800 53.000 ;
        RECT 119.600 51.600 120.400 53.200 ;
        RECT 121.200 52.300 122.000 53.200 ;
        RECT 122.800 52.300 123.600 53.200 ;
        RECT 121.200 51.700 123.600 52.300 ;
        RECT 121.200 51.600 122.000 51.700 ;
        RECT 122.800 51.600 123.600 51.700 ;
        RECT 124.400 51.600 125.200 53.200 ;
        RECT 126.000 53.000 127.400 53.800 ;
        RECT 128.000 53.600 130.000 54.400 ;
        RECT 133.800 53.600 134.800 54.400 ;
        RECT 126.000 51.000 126.600 53.000 ;
        RECT 118.200 50.400 122.000 51.000 ;
        RECT 116.200 49.200 117.800 49.800 ;
        RECT 117.000 44.400 117.800 49.200 ;
        RECT 121.400 47.000 122.000 50.400 ;
        RECT 117.000 43.600 118.800 44.400 ;
        RECT 117.000 42.200 117.800 43.600 ;
        RECT 121.200 43.000 122.000 47.000 ;
        RECT 122.800 50.400 126.600 51.000 ;
        RECT 122.800 47.000 123.400 50.400 ;
        RECT 128.000 49.800 128.600 53.600 ;
        RECT 129.200 50.800 130.000 52.400 ;
        RECT 127.000 49.200 128.600 49.800 ;
        RECT 133.800 50.200 134.400 53.600 ;
        RECT 135.400 53.000 136.000 54.600 ;
        RECT 141.800 54.400 142.400 55.000 ;
        RECT 147.000 54.800 147.600 57.000 ;
        RECT 153.200 56.000 154.000 59.800 ;
        RECT 156.400 56.000 157.200 59.800 ;
        RECT 153.200 55.800 157.200 56.000 ;
        RECT 158.000 55.800 158.800 59.800 ;
        RECT 159.600 55.800 160.400 59.800 ;
        RECT 161.200 56.000 162.000 59.800 ;
        RECT 164.400 56.000 165.200 59.800 ;
        RECT 161.200 55.800 165.200 56.000 ;
        RECT 153.400 55.400 157.000 55.800 ;
        RECT 140.400 53.600 142.400 54.400 ;
        RECT 143.400 54.200 147.600 54.800 ;
        RECT 154.000 54.400 154.800 54.800 ;
        RECT 158.000 54.400 158.600 55.800 ;
        RECT 159.800 54.400 160.400 55.800 ;
        RECT 161.400 55.400 165.000 55.800 ;
        RECT 167.600 55.200 168.400 59.800 ;
        RECT 170.800 55.200 171.600 59.800 ;
        RECT 174.000 55.200 174.800 59.800 ;
        RECT 177.200 55.200 178.000 59.800 ;
        RECT 163.600 54.400 164.400 54.800 ;
        RECT 167.600 54.400 169.400 55.200 ;
        RECT 170.800 54.400 173.000 55.200 ;
        RECT 174.000 54.400 176.200 55.200 ;
        RECT 177.200 54.400 179.600 55.200 ;
        RECT 143.400 53.800 144.400 54.200 ;
        RECT 135.000 52.200 136.000 53.000 ;
        RECT 135.400 50.200 136.000 52.200 ;
        RECT 137.000 52.400 137.800 53.200 ;
        RECT 137.000 52.300 138.000 52.400 ;
        RECT 138.800 52.300 139.600 52.400 ;
        RECT 137.000 51.700 139.600 52.300 ;
        RECT 137.000 51.600 138.000 51.700 ;
        RECT 138.800 51.600 139.600 51.700 ;
        RECT 140.400 50.800 141.200 52.400 ;
        RECT 133.800 49.200 134.800 50.200 ;
        RECT 135.400 49.600 138.000 50.200 ;
        RECT 122.800 43.000 123.600 47.000 ;
        RECT 127.000 44.400 127.800 49.200 ;
        RECT 126.000 43.600 127.800 44.400 ;
        RECT 127.000 42.200 127.800 43.600 ;
        RECT 134.000 42.200 134.800 49.200 ;
        RECT 137.200 42.200 138.000 49.600 ;
        RECT 141.800 49.800 142.400 53.600 ;
        RECT 143.000 53.000 144.400 53.800 ;
        RECT 153.200 53.800 154.800 54.400 ;
        RECT 153.200 53.600 154.000 53.800 ;
        RECT 156.200 53.600 158.800 54.400 ;
        RECT 159.600 53.600 162.200 54.400 ;
        RECT 163.600 53.800 165.200 54.400 ;
        RECT 164.400 53.600 165.200 53.800 ;
        RECT 166.000 53.800 166.800 54.400 ;
        RECT 168.600 53.800 169.400 54.400 ;
        RECT 172.200 53.800 173.000 54.400 ;
        RECT 175.400 53.800 176.200 54.400 ;
        RECT 143.800 51.000 144.400 53.000 ;
        RECT 145.200 51.600 146.000 53.200 ;
        RECT 146.800 51.600 147.600 53.200 ;
        RECT 154.800 51.600 155.600 53.200 ;
        RECT 156.200 52.400 156.800 53.600 ;
        RECT 156.200 51.600 157.200 52.400 ;
        RECT 161.600 52.300 162.200 53.600 ;
        RECT 158.100 51.700 162.200 52.300 ;
        RECT 143.800 50.400 147.600 51.000 ;
        RECT 141.800 49.200 143.400 49.800 ;
        RECT 142.600 42.200 143.400 49.200 ;
        RECT 147.000 47.000 147.600 50.400 ;
        RECT 156.200 50.200 156.800 51.600 ;
        RECT 158.100 50.400 158.700 51.700 ;
        RECT 158.000 50.200 158.800 50.400 ;
        RECT 146.800 43.000 147.600 47.000 ;
        RECT 155.800 49.600 156.800 50.200 ;
        RECT 157.400 49.600 158.800 50.200 ;
        RECT 159.600 50.200 160.400 50.400 ;
        RECT 161.600 50.200 162.200 51.700 ;
        RECT 162.800 51.600 163.600 53.200 ;
        RECT 166.000 53.000 167.800 53.800 ;
        RECT 168.600 53.000 171.200 53.800 ;
        RECT 172.200 53.000 174.600 53.800 ;
        RECT 175.400 53.000 178.000 53.800 ;
        RECT 168.600 51.600 169.400 53.000 ;
        RECT 172.200 51.600 173.000 53.000 ;
        RECT 175.400 51.600 176.200 53.000 ;
        RECT 178.800 51.600 179.600 54.400 ;
        RECT 167.600 50.800 169.400 51.600 ;
        RECT 170.800 50.800 173.000 51.600 ;
        RECT 174.000 50.800 176.200 51.600 ;
        RECT 177.200 50.800 179.600 51.600 ;
        RECT 180.400 53.800 181.200 59.800 ;
        RECT 186.800 56.600 187.600 59.800 ;
        RECT 188.400 57.000 189.200 59.800 ;
        RECT 190.000 57.000 190.800 59.800 ;
        RECT 191.600 57.000 192.400 59.800 ;
        RECT 194.800 57.000 195.600 59.800 ;
        RECT 198.000 57.000 198.800 59.800 ;
        RECT 199.600 57.000 200.400 59.800 ;
        RECT 201.200 57.000 202.000 59.800 ;
        RECT 202.800 57.000 203.600 59.800 ;
        RECT 185.000 55.800 187.600 56.600 ;
        RECT 204.400 56.600 205.200 59.800 ;
        RECT 191.000 55.800 195.600 56.400 ;
        RECT 185.000 55.200 185.800 55.800 ;
        RECT 182.800 54.400 185.800 55.200 ;
        RECT 180.400 53.000 189.200 53.800 ;
        RECT 191.000 53.400 191.800 55.800 ;
        RECT 194.800 55.600 195.600 55.800 ;
        RECT 196.400 55.600 198.000 56.400 ;
        RECT 201.000 55.600 202.000 56.400 ;
        RECT 204.400 55.800 206.800 56.600 ;
        RECT 193.200 53.600 194.000 55.200 ;
        RECT 194.800 54.800 195.600 55.000 ;
        RECT 194.800 54.200 199.200 54.800 ;
        RECT 198.400 54.000 199.200 54.200 ;
        RECT 159.600 49.600 161.000 50.200 ;
        RECT 161.600 49.600 162.600 50.200 ;
        RECT 155.800 42.200 156.600 49.600 ;
        RECT 157.400 48.400 158.000 49.600 ;
        RECT 157.200 47.600 158.000 48.400 ;
        RECT 160.400 48.400 161.000 49.600 ;
        RECT 160.400 47.600 161.200 48.400 ;
        RECT 161.800 42.200 162.600 49.600 ;
        RECT 167.600 42.200 168.400 50.800 ;
        RECT 170.800 42.200 171.600 50.800 ;
        RECT 174.000 42.200 174.800 50.800 ;
        RECT 177.200 42.200 178.000 50.800 ;
        RECT 180.400 47.400 181.200 53.000 ;
        RECT 189.800 52.600 191.800 53.400 ;
        RECT 195.600 52.600 198.800 53.400 ;
        RECT 201.200 52.800 202.000 55.600 ;
        RECT 206.000 55.200 206.800 55.800 ;
        RECT 206.000 54.600 207.800 55.200 ;
        RECT 207.000 53.400 207.800 54.600 ;
        RECT 210.800 54.600 211.600 59.800 ;
        RECT 212.400 56.000 213.200 59.800 ;
        RECT 218.200 56.400 219.000 59.800 ;
        RECT 212.400 55.200 213.400 56.000 ;
        RECT 217.200 55.800 219.000 56.400 ;
        RECT 210.800 54.000 212.000 54.600 ;
        RECT 207.000 52.600 210.800 53.400 ;
        RECT 181.800 52.000 182.600 52.200 ;
        RECT 185.200 52.000 186.000 52.400 ;
        RECT 186.800 52.000 187.600 52.400 ;
        RECT 204.400 52.000 205.200 52.600 ;
        RECT 211.400 52.000 212.000 54.000 ;
        RECT 181.800 51.400 205.200 52.000 ;
        RECT 211.200 51.400 212.000 52.000 ;
        RECT 211.200 49.600 211.800 51.400 ;
        RECT 212.600 50.800 213.400 55.200 ;
        RECT 215.600 53.600 216.400 55.200 ;
        RECT 190.000 49.400 190.800 49.600 ;
        RECT 185.400 49.000 190.800 49.400 ;
        RECT 184.600 48.800 190.800 49.000 ;
        RECT 191.800 49.000 200.400 49.600 ;
        RECT 182.000 48.000 183.600 48.800 ;
        RECT 184.600 48.200 186.000 48.800 ;
        RECT 191.800 48.200 192.400 49.000 ;
        RECT 199.600 48.800 200.400 49.000 ;
        RECT 202.800 49.000 211.800 49.600 ;
        RECT 202.800 48.800 203.600 49.000 ;
        RECT 183.000 47.600 183.600 48.000 ;
        RECT 186.600 47.600 192.400 48.200 ;
        RECT 193.000 47.600 195.600 48.400 ;
        RECT 180.400 46.800 182.400 47.400 ;
        RECT 183.000 46.800 187.200 47.600 ;
        RECT 181.800 46.200 182.400 46.800 ;
        RECT 181.800 45.600 182.800 46.200 ;
        RECT 182.000 42.200 182.800 45.600 ;
        RECT 185.200 42.200 186.000 46.800 ;
        RECT 188.400 42.200 189.200 45.000 ;
        RECT 190.000 42.200 190.800 45.000 ;
        RECT 191.600 42.200 192.400 47.000 ;
        RECT 194.800 42.200 195.600 47.000 ;
        RECT 198.000 42.200 198.800 48.400 ;
        RECT 206.000 47.600 208.600 48.400 ;
        RECT 201.200 46.800 205.400 47.600 ;
        RECT 199.600 42.200 200.400 45.000 ;
        RECT 201.200 42.200 202.000 45.000 ;
        RECT 202.800 42.200 203.600 45.000 ;
        RECT 206.000 42.200 206.800 47.600 ;
        RECT 211.200 47.400 211.800 49.000 ;
        RECT 209.200 46.800 211.800 47.400 ;
        RECT 212.400 50.000 213.400 50.800 ;
        RECT 209.200 42.200 210.000 46.800 ;
        RECT 212.400 42.200 213.200 50.000 ;
        RECT 217.200 42.200 218.000 55.800 ;
        RECT 218.800 48.800 219.600 50.400 ;
        RECT 220.400 42.200 221.200 59.800 ;
        RECT 222.000 55.600 222.800 57.200 ;
        RECT 226.200 56.400 227.000 59.800 ;
        RECT 231.000 56.400 231.800 59.800 ;
        RECT 225.200 55.800 227.000 56.400 ;
        RECT 230.000 55.800 231.800 56.400 ;
        RECT 233.200 55.800 234.000 59.800 ;
        RECT 234.800 56.000 235.600 59.800 ;
        RECT 238.000 56.000 238.800 59.800 ;
        RECT 234.800 55.800 238.800 56.000 ;
        RECT 223.600 53.600 224.400 55.200 ;
        RECT 223.600 48.300 224.400 48.400 ;
        RECT 225.200 48.300 226.000 55.800 ;
        RECT 228.400 53.600 229.200 55.200 ;
        RECT 230.000 52.300 230.800 55.800 ;
        RECT 233.400 54.400 234.000 55.800 ;
        RECT 235.000 55.400 238.600 55.800 ;
        RECT 237.200 54.400 238.000 54.800 ;
        RECT 233.200 53.600 235.800 54.400 ;
        RECT 237.200 53.800 238.800 54.400 ;
        RECT 238.000 53.600 238.800 53.800 ;
        RECT 230.000 51.700 233.900 52.300 ;
        RECT 226.800 48.800 227.600 50.400 ;
        RECT 223.600 47.700 226.000 48.300 ;
        RECT 223.600 47.600 224.400 47.700 ;
        RECT 225.200 42.200 226.000 47.700 ;
        RECT 230.000 42.200 230.800 51.700 ;
        RECT 233.300 50.400 233.900 51.700 ;
        RECT 235.200 50.400 235.800 53.600 ;
        RECT 236.400 52.300 237.200 53.200 ;
        RECT 239.600 52.300 240.400 59.800 ;
        RECT 241.200 55.600 242.000 57.200 ;
        RECT 236.400 51.700 240.400 52.300 ;
        RECT 236.400 51.600 237.200 51.700 ;
        RECT 231.600 48.800 232.400 50.400 ;
        RECT 233.200 50.200 234.000 50.400 ;
        RECT 233.200 49.600 234.600 50.200 ;
        RECT 235.200 49.600 237.200 50.400 ;
        RECT 234.000 48.400 234.600 49.600 ;
        RECT 234.000 47.600 234.800 48.400 ;
        RECT 235.400 42.200 236.200 49.600 ;
        RECT 239.600 42.200 240.400 51.700 ;
        RECT 242.800 53.800 243.600 59.800 ;
        RECT 249.200 56.600 250.000 59.800 ;
        RECT 250.800 57.000 251.600 59.800 ;
        RECT 252.400 57.000 253.200 59.800 ;
        RECT 254.000 57.000 254.800 59.800 ;
        RECT 257.200 57.000 258.000 59.800 ;
        RECT 260.400 57.000 261.200 59.800 ;
        RECT 262.000 57.000 262.800 59.800 ;
        RECT 263.600 57.000 264.400 59.800 ;
        RECT 265.200 57.000 266.000 59.800 ;
        RECT 247.400 55.800 250.000 56.600 ;
        RECT 266.800 56.600 267.600 59.800 ;
        RECT 253.400 55.800 258.000 56.400 ;
        RECT 247.400 55.200 248.200 55.800 ;
        RECT 245.200 54.400 248.200 55.200 ;
        RECT 242.800 53.000 251.600 53.800 ;
        RECT 253.400 53.400 254.200 55.800 ;
        RECT 257.200 55.600 258.000 55.800 ;
        RECT 258.800 55.600 260.400 56.400 ;
        RECT 263.400 55.600 264.400 56.400 ;
        RECT 266.800 55.800 269.200 56.600 ;
        RECT 255.600 53.600 256.400 55.200 ;
        RECT 257.200 54.800 258.000 55.000 ;
        RECT 257.200 54.200 261.600 54.800 ;
        RECT 260.800 54.000 261.600 54.200 ;
        RECT 242.800 47.400 243.600 53.000 ;
        RECT 252.200 52.600 254.200 53.400 ;
        RECT 258.000 52.600 261.200 53.400 ;
        RECT 263.600 52.800 264.400 55.600 ;
        RECT 268.400 55.200 269.200 55.800 ;
        RECT 268.400 54.600 270.200 55.200 ;
        RECT 269.400 53.400 270.200 54.600 ;
        RECT 273.200 54.600 274.000 59.800 ;
        RECT 274.800 56.000 275.600 59.800 ;
        RECT 278.000 56.000 278.800 59.800 ;
        RECT 281.200 56.000 282.000 59.800 ;
        RECT 274.800 55.200 275.800 56.000 ;
        RECT 278.000 55.800 282.000 56.000 ;
        RECT 282.800 55.800 283.600 59.800 ;
        RECT 284.400 55.800 285.200 59.800 ;
        RECT 286.000 56.000 286.800 59.800 ;
        RECT 289.200 56.000 290.000 59.800 ;
        RECT 286.000 55.800 290.000 56.000 ;
        RECT 278.200 55.400 281.800 55.800 ;
        RECT 273.200 54.000 274.400 54.600 ;
        RECT 269.400 52.600 273.200 53.400 ;
        RECT 244.200 52.000 245.000 52.200 ;
        RECT 246.000 52.000 246.800 52.400 ;
        RECT 249.200 52.000 250.000 52.400 ;
        RECT 266.800 52.000 267.600 52.600 ;
        RECT 273.800 52.000 274.400 54.000 ;
        RECT 244.200 51.400 267.600 52.000 ;
        RECT 273.600 51.400 274.400 52.000 ;
        RECT 273.600 49.600 274.200 51.400 ;
        RECT 275.000 50.800 275.800 55.200 ;
        RECT 278.800 54.400 279.600 54.800 ;
        RECT 282.800 54.400 283.400 55.800 ;
        RECT 284.600 54.400 285.200 55.800 ;
        RECT 286.200 55.400 289.800 55.800 ;
        RECT 288.400 54.400 289.200 54.800 ;
        RECT 278.000 53.800 279.600 54.400 ;
        RECT 278.000 53.600 278.800 53.800 ;
        RECT 281.000 53.600 283.600 54.400 ;
        RECT 284.400 53.600 287.000 54.400 ;
        RECT 288.400 53.800 290.000 54.400 ;
        RECT 289.200 53.600 290.000 53.800 ;
        RECT 295.600 53.800 296.400 59.800 ;
        RECT 302.000 56.600 302.800 59.800 ;
        RECT 303.600 57.000 304.400 59.800 ;
        RECT 305.200 57.000 306.000 59.800 ;
        RECT 306.800 57.000 307.600 59.800 ;
        RECT 310.000 57.000 310.800 59.800 ;
        RECT 313.200 57.000 314.000 59.800 ;
        RECT 314.800 57.000 315.600 59.800 ;
        RECT 316.400 57.000 317.200 59.800 ;
        RECT 318.000 57.000 318.800 59.800 ;
        RECT 300.200 55.800 302.800 56.600 ;
        RECT 319.600 56.600 320.400 59.800 ;
        RECT 306.200 55.800 310.800 56.400 ;
        RECT 300.200 55.200 301.000 55.800 ;
        RECT 298.000 54.400 301.000 55.200 ;
        RECT 279.600 51.600 280.400 53.200 ;
        RECT 252.400 49.400 253.200 49.600 ;
        RECT 247.800 49.000 253.200 49.400 ;
        RECT 247.000 48.800 253.200 49.000 ;
        RECT 254.200 49.000 262.800 49.600 ;
        RECT 244.400 48.000 246.000 48.800 ;
        RECT 247.000 48.200 248.400 48.800 ;
        RECT 254.200 48.200 254.800 49.000 ;
        RECT 262.000 48.800 262.800 49.000 ;
        RECT 265.200 49.000 274.200 49.600 ;
        RECT 265.200 48.800 266.000 49.000 ;
        RECT 245.400 47.600 246.000 48.000 ;
        RECT 249.000 47.600 254.800 48.200 ;
        RECT 255.400 47.600 258.000 48.400 ;
        RECT 242.800 46.800 244.800 47.400 ;
        RECT 245.400 46.800 249.600 47.600 ;
        RECT 244.200 46.200 244.800 46.800 ;
        RECT 244.200 45.600 245.200 46.200 ;
        RECT 244.400 42.200 245.200 45.600 ;
        RECT 247.600 42.200 248.400 46.800 ;
        RECT 250.800 42.200 251.600 45.000 ;
        RECT 252.400 42.200 253.200 45.000 ;
        RECT 254.000 42.200 254.800 47.000 ;
        RECT 257.200 42.200 258.000 47.000 ;
        RECT 260.400 42.200 261.200 48.400 ;
        RECT 268.400 47.600 271.000 48.400 ;
        RECT 263.600 46.800 267.800 47.600 ;
        RECT 262.000 42.200 262.800 45.000 ;
        RECT 263.600 42.200 264.400 45.000 ;
        RECT 265.200 42.200 266.000 45.000 ;
        RECT 268.400 42.200 269.200 47.600 ;
        RECT 273.600 47.400 274.200 49.000 ;
        RECT 271.600 46.800 274.200 47.400 ;
        RECT 274.800 50.000 275.800 50.800 ;
        RECT 281.000 50.200 281.600 53.600 ;
        RECT 282.800 50.200 283.600 50.400 ;
        RECT 271.600 42.200 272.400 46.800 ;
        RECT 274.800 42.200 275.600 50.000 ;
        RECT 280.600 49.600 281.600 50.200 ;
        RECT 282.200 49.600 283.600 50.200 ;
        RECT 284.400 50.200 285.200 50.400 ;
        RECT 286.400 50.200 287.000 53.600 ;
        RECT 287.600 52.300 288.400 53.200 ;
        RECT 295.600 53.000 304.400 53.800 ;
        RECT 306.200 53.400 307.000 55.800 ;
        RECT 310.000 55.600 310.800 55.800 ;
        RECT 311.600 55.600 313.200 56.400 ;
        RECT 316.200 55.600 317.200 56.400 ;
        RECT 319.600 55.800 322.000 56.600 ;
        RECT 308.400 53.600 309.200 55.200 ;
        RECT 310.000 54.800 310.800 55.000 ;
        RECT 310.000 54.200 314.400 54.800 ;
        RECT 313.600 54.000 314.400 54.200 ;
        RECT 289.200 52.300 290.000 52.400 ;
        RECT 287.600 51.700 290.000 52.300 ;
        RECT 287.600 51.600 288.400 51.700 ;
        RECT 289.200 51.600 290.000 51.700 ;
        RECT 284.400 49.600 285.800 50.200 ;
        RECT 286.400 49.600 287.400 50.200 ;
        RECT 280.600 44.400 281.400 49.600 ;
        RECT 282.200 48.400 282.800 49.600 ;
        RECT 282.000 47.600 282.800 48.400 ;
        RECT 285.200 48.400 285.800 49.600 ;
        RECT 285.200 47.600 286.000 48.400 ;
        RECT 279.600 43.600 281.400 44.400 ;
        RECT 280.600 42.200 281.400 43.600 ;
        RECT 286.600 44.400 287.400 49.600 ;
        RECT 295.600 47.400 296.400 53.000 ;
        RECT 305.000 52.600 307.000 53.400 ;
        RECT 310.800 52.600 314.000 53.400 ;
        RECT 316.400 52.800 317.200 55.600 ;
        RECT 321.200 55.200 322.000 55.800 ;
        RECT 321.200 54.600 323.000 55.200 ;
        RECT 322.200 53.400 323.000 54.600 ;
        RECT 326.000 54.600 326.800 59.800 ;
        RECT 327.600 56.000 328.400 59.800 ;
        RECT 334.600 56.000 335.400 59.000 ;
        RECT 338.800 57.000 339.600 59.000 ;
        RECT 327.600 55.200 328.600 56.000 ;
        RECT 326.000 54.000 327.200 54.600 ;
        RECT 322.200 52.600 326.000 53.400 ;
        RECT 297.200 52.200 298.000 52.400 ;
        RECT 297.000 52.000 298.000 52.200 ;
        RECT 302.000 52.000 302.800 52.400 ;
        RECT 319.600 52.000 320.400 52.600 ;
        RECT 326.600 52.000 327.200 54.000 ;
        RECT 297.000 51.400 320.400 52.000 ;
        RECT 326.400 51.400 327.200 52.000 ;
        RECT 326.400 49.600 327.000 51.400 ;
        RECT 327.800 50.800 328.600 55.200 ;
        RECT 333.800 55.400 335.400 56.000 ;
        RECT 333.800 55.000 334.600 55.400 ;
        RECT 333.800 54.400 334.400 55.000 ;
        RECT 339.000 54.800 339.600 57.000 ;
        RECT 343.000 56.400 343.800 59.800 ;
        RECT 342.000 55.800 343.800 56.400 ;
        RECT 345.800 56.400 346.600 59.800 ;
        RECT 345.800 55.800 347.600 56.400 ;
        RECT 332.400 53.600 334.400 54.400 ;
        RECT 335.400 54.200 339.600 54.800 ;
        RECT 335.400 53.800 336.400 54.200 ;
        RECT 330.800 52.300 331.600 52.400 ;
        RECT 332.400 52.300 333.200 52.400 ;
        RECT 330.800 51.700 333.200 52.300 ;
        RECT 330.800 51.600 331.600 51.700 ;
        RECT 332.400 50.800 333.200 51.700 ;
        RECT 305.200 49.400 306.000 49.600 ;
        RECT 300.600 49.000 306.000 49.400 ;
        RECT 299.800 48.800 306.000 49.000 ;
        RECT 307.000 49.000 315.600 49.600 ;
        RECT 297.200 48.000 298.800 48.800 ;
        RECT 299.800 48.200 301.200 48.800 ;
        RECT 307.000 48.200 307.600 49.000 ;
        RECT 314.800 48.800 315.600 49.000 ;
        RECT 318.000 49.000 327.000 49.600 ;
        RECT 318.000 48.800 318.800 49.000 ;
        RECT 298.200 47.600 298.800 48.000 ;
        RECT 301.800 47.600 307.600 48.200 ;
        RECT 308.200 47.600 310.800 48.400 ;
        RECT 295.600 46.800 297.600 47.400 ;
        RECT 298.200 46.800 302.400 47.600 ;
        RECT 297.000 46.200 297.600 46.800 ;
        RECT 297.000 45.600 298.000 46.200 ;
        RECT 286.600 43.600 288.400 44.400 ;
        RECT 286.600 42.200 287.400 43.600 ;
        RECT 297.200 42.200 298.000 45.600 ;
        RECT 300.400 42.200 301.200 46.800 ;
        RECT 303.600 42.200 304.400 45.000 ;
        RECT 305.200 42.200 306.000 45.000 ;
        RECT 306.800 42.200 307.600 47.000 ;
        RECT 310.000 42.200 310.800 47.000 ;
        RECT 313.200 42.200 314.000 48.400 ;
        RECT 321.200 47.600 323.800 48.400 ;
        RECT 316.400 46.800 320.600 47.600 ;
        RECT 314.800 42.200 315.600 45.000 ;
        RECT 316.400 42.200 317.200 45.000 ;
        RECT 318.000 42.200 318.800 45.000 ;
        RECT 321.200 42.200 322.000 47.600 ;
        RECT 326.400 47.400 327.000 49.000 ;
        RECT 324.400 46.800 327.000 47.400 ;
        RECT 327.600 50.000 328.600 50.800 ;
        RECT 324.400 42.200 325.200 46.800 ;
        RECT 327.600 42.200 328.400 50.000 ;
        RECT 333.800 49.800 334.400 53.600 ;
        RECT 335.000 53.000 336.400 53.800 ;
        RECT 340.400 53.600 341.200 55.200 ;
        RECT 335.800 51.000 336.400 53.000 ;
        RECT 337.200 51.600 338.000 53.200 ;
        RECT 338.800 51.600 339.600 53.200 ;
        RECT 342.000 52.300 342.800 55.800 ;
        RECT 346.800 52.300 347.600 55.800 ;
        RECT 353.200 55.800 354.000 59.800 ;
        RECT 354.600 56.400 355.400 57.200 ;
        RECT 348.400 53.600 349.200 55.200 ;
        RECT 351.600 52.800 352.400 54.400 ;
        RECT 350.000 52.300 350.800 52.400 ;
        RECT 342.000 51.700 345.900 52.300 ;
        RECT 335.800 50.400 339.600 51.000 ;
        RECT 333.800 49.200 335.400 49.800 ;
        RECT 334.600 44.400 335.400 49.200 ;
        RECT 339.000 47.000 339.600 50.400 ;
        RECT 334.000 43.600 335.400 44.400 ;
        RECT 334.600 42.200 335.400 43.600 ;
        RECT 338.800 43.000 339.600 47.000 ;
        RECT 342.000 42.200 342.800 51.700 ;
        RECT 345.300 50.400 345.900 51.700 ;
        RECT 346.800 52.200 350.800 52.300 ;
        RECT 353.200 52.200 353.800 55.800 ;
        RECT 354.800 55.600 355.600 56.400 ;
        RECT 356.400 56.000 357.200 59.800 ;
        RECT 359.600 56.000 360.400 59.800 ;
        RECT 356.400 55.800 360.400 56.000 ;
        RECT 356.600 55.400 360.200 55.800 ;
        RECT 361.200 55.600 362.000 59.800 ;
        RECT 362.800 55.800 363.600 59.800 ;
        RECT 367.000 58.400 367.800 59.800 ;
        RECT 367.000 57.600 368.400 58.400 ;
        RECT 367.000 56.800 367.800 57.600 ;
        RECT 367.000 55.800 368.400 56.800 ;
        RECT 363.000 55.600 363.600 55.800 ;
        RECT 357.200 54.400 358.000 54.800 ;
        RECT 361.200 54.400 361.800 55.600 ;
        RECT 363.000 55.200 364.800 55.600 ;
        RECT 363.000 55.000 367.200 55.200 ;
        RECT 364.200 54.600 367.200 55.000 ;
        RECT 366.400 54.400 367.200 54.600 ;
        RECT 354.800 54.300 355.600 54.400 ;
        RECT 356.400 54.300 358.000 54.400 ;
        RECT 354.800 53.800 358.000 54.300 ;
        RECT 354.800 53.700 357.200 53.800 ;
        RECT 354.800 53.600 355.600 53.700 ;
        RECT 356.400 53.600 357.200 53.700 ;
        RECT 359.400 53.600 362.000 54.400 ;
        RECT 354.800 52.200 355.600 52.400 ;
        RECT 346.800 51.700 351.600 52.200 ;
        RECT 343.600 48.800 344.400 50.400 ;
        RECT 345.200 48.800 346.000 50.400 ;
        RECT 346.800 42.200 347.600 51.700 ;
        RECT 350.000 51.600 351.600 51.700 ;
        RECT 353.200 51.600 355.600 52.200 ;
        RECT 358.000 51.600 358.800 53.200 ;
        RECT 350.800 51.200 351.600 51.600 ;
        RECT 354.800 50.200 355.400 51.600 ;
        RECT 359.400 50.200 360.000 53.600 ;
        RECT 362.800 52.800 363.600 54.400 ;
        RECT 364.800 53.800 365.600 54.000 ;
        RECT 364.600 53.200 365.600 53.800 ;
        RECT 364.600 52.400 365.200 53.200 ;
        RECT 364.400 51.600 365.200 52.400 ;
        RECT 366.400 51.000 367.000 54.400 ;
        RECT 367.800 52.400 368.400 55.800 ;
        RECT 369.200 55.600 370.000 57.200 ;
        RECT 367.600 51.600 368.400 52.400 ;
        RECT 364.600 50.400 367.000 51.000 ;
        RECT 361.200 50.200 362.000 50.400 ;
        RECT 350.000 49.600 354.000 50.200 ;
        RECT 350.000 42.200 350.800 49.600 ;
        RECT 353.200 42.200 354.000 49.600 ;
        RECT 354.800 42.200 355.600 50.200 ;
        RECT 359.000 49.600 360.000 50.200 ;
        RECT 360.600 49.600 362.000 50.200 ;
        RECT 359.000 42.200 359.800 49.600 ;
        RECT 360.600 48.400 361.200 49.600 ;
        RECT 360.400 47.600 361.200 48.400 ;
        RECT 364.600 46.200 365.200 50.400 ;
        RECT 367.800 50.200 368.400 51.600 ;
        RECT 364.400 42.200 365.200 46.200 ;
        RECT 367.600 42.200 368.400 50.200 ;
        RECT 370.800 42.200 371.600 59.800 ;
        RECT 372.400 53.800 373.200 59.800 ;
        RECT 378.800 56.600 379.600 59.800 ;
        RECT 380.400 57.000 381.200 59.800 ;
        RECT 382.000 57.000 382.800 59.800 ;
        RECT 383.600 57.000 384.400 59.800 ;
        RECT 386.800 57.000 387.600 59.800 ;
        RECT 390.000 57.000 390.800 59.800 ;
        RECT 391.600 57.000 392.400 59.800 ;
        RECT 393.200 57.000 394.000 59.800 ;
        RECT 394.800 57.000 395.600 59.800 ;
        RECT 377.000 55.800 379.600 56.600 ;
        RECT 396.400 56.600 397.200 59.800 ;
        RECT 383.000 55.800 387.600 56.400 ;
        RECT 377.000 55.200 377.800 55.800 ;
        RECT 374.800 54.400 377.800 55.200 ;
        RECT 372.400 53.000 381.200 53.800 ;
        RECT 383.000 53.400 383.800 55.800 ;
        RECT 386.800 55.600 387.600 55.800 ;
        RECT 388.400 55.600 390.000 56.400 ;
        RECT 393.000 55.600 394.000 56.400 ;
        RECT 396.400 55.800 398.800 56.600 ;
        RECT 385.200 53.600 386.000 55.200 ;
        RECT 386.800 54.800 387.600 55.000 ;
        RECT 386.800 54.200 391.200 54.800 ;
        RECT 390.400 54.000 391.200 54.200 ;
        RECT 372.400 47.400 373.200 53.000 ;
        RECT 381.800 52.600 383.800 53.400 ;
        RECT 387.600 52.600 390.800 53.400 ;
        RECT 393.200 52.800 394.000 55.600 ;
        RECT 398.000 55.200 398.800 55.800 ;
        RECT 398.000 54.600 399.800 55.200 ;
        RECT 399.000 53.400 399.800 54.600 ;
        RECT 402.800 54.600 403.600 59.800 ;
        RECT 404.400 56.000 405.200 59.800 ;
        RECT 404.400 55.200 405.400 56.000 ;
        RECT 402.800 54.000 404.000 54.600 ;
        RECT 399.000 52.600 402.800 53.400 ;
        RECT 373.800 52.000 374.600 52.200 ;
        RECT 375.600 52.000 376.400 52.400 ;
        RECT 378.800 52.000 379.600 52.400 ;
        RECT 385.200 52.000 386.000 52.400 ;
        RECT 396.400 52.000 397.200 52.600 ;
        RECT 403.400 52.000 404.000 54.000 ;
        RECT 373.800 51.400 397.200 52.000 ;
        RECT 403.200 51.400 404.000 52.000 ;
        RECT 403.200 49.600 403.800 51.400 ;
        RECT 404.600 50.800 405.400 55.200 ;
        RECT 407.600 55.000 408.400 59.800 ;
        RECT 412.000 58.400 412.800 59.800 ;
        RECT 410.800 57.800 412.800 58.400 ;
        RECT 416.400 57.800 417.200 59.800 ;
        RECT 420.600 58.400 421.800 59.800 ;
        RECT 420.400 57.800 421.800 58.400 ;
        RECT 410.800 57.000 411.600 57.800 ;
        RECT 416.400 57.200 417.000 57.800 ;
        RECT 412.400 56.400 413.200 57.200 ;
        RECT 414.200 56.600 417.000 57.200 ;
        RECT 420.400 57.000 421.200 57.800 ;
        RECT 414.200 56.400 415.000 56.600 ;
        RECT 408.400 54.200 410.000 54.400 ;
        RECT 412.600 54.200 413.200 56.400 ;
        RECT 422.200 55.400 423.000 55.600 ;
        RECT 425.200 55.400 426.000 59.800 ;
        RECT 426.800 55.600 427.600 57.200 ;
        RECT 422.200 54.800 426.000 55.400 ;
        RECT 418.200 54.200 419.000 54.400 ;
        RECT 408.400 53.600 419.400 54.200 ;
        RECT 411.400 53.400 412.200 53.600 ;
        RECT 409.800 52.400 410.600 52.600 ;
        RECT 418.800 52.400 419.400 53.600 ;
        RECT 420.400 52.800 421.200 53.000 ;
        RECT 409.800 51.800 414.800 52.400 ;
        RECT 414.000 51.600 414.800 51.800 ;
        RECT 418.800 51.600 419.600 52.400 ;
        RECT 420.400 52.200 424.200 52.800 ;
        RECT 423.400 52.000 424.200 52.200 ;
        RECT 382.000 49.400 382.800 49.600 ;
        RECT 377.400 49.000 382.800 49.400 ;
        RECT 376.600 48.800 382.800 49.000 ;
        RECT 383.800 49.000 392.400 49.600 ;
        RECT 374.000 48.000 375.600 48.800 ;
        RECT 376.600 48.200 378.000 48.800 ;
        RECT 383.800 48.200 384.400 49.000 ;
        RECT 391.600 48.800 392.400 49.000 ;
        RECT 394.800 49.000 403.800 49.600 ;
        RECT 394.800 48.800 395.600 49.000 ;
        RECT 375.000 47.600 375.600 48.000 ;
        RECT 378.600 47.600 384.400 48.200 ;
        RECT 385.000 47.600 387.600 48.400 ;
        RECT 372.400 46.800 374.400 47.400 ;
        RECT 375.000 46.800 379.200 47.600 ;
        RECT 373.800 46.200 374.400 46.800 ;
        RECT 373.800 45.600 374.800 46.200 ;
        RECT 374.000 42.200 374.800 45.600 ;
        RECT 377.200 42.200 378.000 46.800 ;
        RECT 380.400 42.200 381.200 45.000 ;
        RECT 382.000 42.200 382.800 45.000 ;
        RECT 383.600 42.200 384.400 47.000 ;
        RECT 386.800 42.200 387.600 47.000 ;
        RECT 390.000 42.200 390.800 48.400 ;
        RECT 398.000 47.600 400.600 48.400 ;
        RECT 393.200 46.800 397.400 47.600 ;
        RECT 391.600 42.200 392.400 45.000 ;
        RECT 393.200 42.200 394.000 45.000 ;
        RECT 394.800 42.200 395.600 45.000 ;
        RECT 398.000 42.200 398.800 47.600 ;
        RECT 403.200 47.400 403.800 49.000 ;
        RECT 401.200 46.800 403.800 47.400 ;
        RECT 404.400 50.000 405.400 50.800 ;
        RECT 407.600 51.000 413.200 51.200 ;
        RECT 407.600 50.800 413.400 51.000 ;
        RECT 407.600 50.600 417.400 50.800 ;
        RECT 401.200 42.200 402.000 46.800 ;
        RECT 404.400 42.200 405.200 50.000 ;
        RECT 407.600 42.200 408.400 50.600 ;
        RECT 412.600 50.200 417.400 50.600 ;
        RECT 410.800 49.000 416.200 49.600 ;
        RECT 410.800 48.800 411.600 49.000 ;
        RECT 415.400 48.800 416.200 49.000 ;
        RECT 416.800 49.000 417.400 50.200 ;
        RECT 418.800 50.400 419.400 51.600 ;
        RECT 421.800 51.400 422.600 51.600 ;
        RECT 425.200 51.400 426.000 54.800 ;
        RECT 421.800 50.800 426.000 51.400 ;
        RECT 418.800 49.800 421.200 50.400 ;
        RECT 418.200 49.000 419.000 49.200 ;
        RECT 416.800 48.400 419.000 49.000 ;
        RECT 420.600 48.800 421.200 49.800 ;
        RECT 420.600 48.000 422.000 48.800 ;
        RECT 414.200 47.400 415.000 47.600 ;
        RECT 417.000 47.400 417.800 47.600 ;
        RECT 410.800 46.200 411.600 47.000 ;
        RECT 414.200 46.800 417.800 47.400 ;
        RECT 416.400 46.200 417.000 46.800 ;
        RECT 420.400 46.200 421.200 47.000 ;
        RECT 410.800 45.600 412.800 46.200 ;
        RECT 412.000 42.200 412.800 45.600 ;
        RECT 416.400 42.200 417.200 46.200 ;
        RECT 420.600 42.200 421.800 46.200 ;
        RECT 425.200 42.200 426.000 50.800 ;
        RECT 428.400 54.300 429.200 59.800 ;
        RECT 430.000 56.000 430.800 59.800 ;
        RECT 433.200 56.000 434.000 59.800 ;
        RECT 430.000 55.800 434.000 56.000 ;
        RECT 434.800 55.800 435.600 59.800 ;
        RECT 436.400 55.800 437.200 59.800 ;
        RECT 438.000 56.000 438.800 59.800 ;
        RECT 441.200 56.000 442.000 59.800 ;
        RECT 438.000 55.800 442.000 56.000 ;
        RECT 430.200 55.400 433.800 55.800 ;
        RECT 430.800 54.400 431.600 54.800 ;
        RECT 434.800 54.400 435.400 55.800 ;
        RECT 436.600 54.400 437.200 55.800 ;
        RECT 438.200 55.400 441.800 55.800 ;
        RECT 442.800 55.600 443.600 59.800 ;
        RECT 444.400 56.000 445.200 59.800 ;
        RECT 447.600 56.000 448.400 59.800 ;
        RECT 453.000 56.400 453.800 59.000 ;
        RECT 457.200 57.000 458.000 59.000 ;
        RECT 458.800 58.300 459.600 58.400 ;
        RECT 463.600 58.300 464.400 59.800 ;
        RECT 458.800 57.700 464.400 58.300 ;
        RECT 458.800 57.600 459.600 57.700 ;
        RECT 452.400 56.000 453.800 56.400 ;
        RECT 444.400 55.800 448.400 56.000 ;
        RECT 440.400 54.400 441.200 54.800 ;
        RECT 443.000 54.400 443.600 55.600 ;
        RECT 444.600 55.400 448.200 55.800 ;
        RECT 452.200 55.400 453.800 56.000 ;
        RECT 452.200 55.000 453.000 55.400 ;
        RECT 446.800 54.400 447.600 54.800 ;
        RECT 452.200 54.400 452.800 55.000 ;
        RECT 457.400 54.800 458.000 57.000 ;
        RECT 463.600 55.800 464.400 57.700 ;
        RECT 465.200 56.000 466.000 59.800 ;
        RECT 468.400 56.000 469.200 59.800 ;
        RECT 465.200 55.800 469.200 56.000 ;
        RECT 430.000 54.300 431.600 54.400 ;
        RECT 428.400 53.800 431.600 54.300 ;
        RECT 428.400 53.700 430.800 53.800 ;
        RECT 428.400 42.200 429.200 53.700 ;
        RECT 430.000 53.600 430.800 53.700 ;
        RECT 433.000 53.600 435.600 54.400 ;
        RECT 436.400 53.600 439.000 54.400 ;
        RECT 440.400 53.800 442.000 54.400 ;
        RECT 441.200 53.600 442.000 53.800 ;
        RECT 442.800 53.600 445.400 54.400 ;
        RECT 446.800 53.800 448.400 54.400 ;
        RECT 447.600 53.600 448.400 53.800 ;
        RECT 450.800 53.600 452.800 54.400 ;
        RECT 453.800 54.200 458.000 54.800 ;
        RECT 463.800 54.400 464.400 55.800 ;
        RECT 465.400 55.400 469.000 55.800 ;
        RECT 467.600 54.400 468.400 54.800 ;
        RECT 453.800 53.800 454.800 54.200 ;
        RECT 431.600 51.600 432.400 53.200 ;
        RECT 433.000 50.200 433.600 53.600 ;
        RECT 438.400 50.400 439.000 53.600 ;
        RECT 439.600 51.600 440.400 53.200 ;
        RECT 434.800 50.200 435.600 50.400 ;
        RECT 432.600 49.600 433.600 50.200 ;
        RECT 434.200 49.600 435.600 50.200 ;
        RECT 436.400 50.200 437.200 50.400 ;
        RECT 436.400 49.600 437.800 50.200 ;
        RECT 438.400 49.600 440.400 50.400 ;
        RECT 442.800 50.200 443.600 50.400 ;
        RECT 444.800 50.200 445.400 53.600 ;
        RECT 446.000 51.600 446.800 53.200 ;
        RECT 447.600 52.300 448.400 52.400 ;
        RECT 450.800 52.300 451.600 52.400 ;
        RECT 447.600 51.700 451.600 52.300 ;
        RECT 447.600 51.600 448.400 51.700 ;
        RECT 450.800 50.800 451.600 51.700 ;
        RECT 442.800 49.600 444.200 50.200 ;
        RECT 444.800 49.600 445.800 50.200 ;
        RECT 432.600 42.200 433.400 49.600 ;
        RECT 434.200 48.400 434.800 49.600 ;
        RECT 434.000 47.600 434.800 48.400 ;
        RECT 437.200 48.400 437.800 49.600 ;
        RECT 437.200 47.600 438.000 48.400 ;
        RECT 438.600 42.200 439.400 49.600 ;
        RECT 443.600 48.400 444.200 49.600 ;
        RECT 443.600 47.600 444.400 48.400 ;
        RECT 445.000 42.200 445.800 49.600 ;
        RECT 452.200 49.800 452.800 53.600 ;
        RECT 453.400 53.000 454.800 53.800 ;
        RECT 463.600 53.600 466.200 54.400 ;
        RECT 467.600 54.300 469.200 54.400 ;
        RECT 470.000 54.300 470.800 59.800 ;
        RECT 471.600 55.600 472.400 57.200 ;
        RECT 473.200 57.000 474.000 59.000 ;
        RECT 467.600 53.800 470.800 54.300 ;
        RECT 473.200 54.800 473.800 57.000 ;
        RECT 477.400 56.000 478.200 59.000 ;
        RECT 477.400 55.400 479.000 56.000 ;
        RECT 478.200 55.000 479.000 55.400 ;
        RECT 482.800 55.000 483.600 59.800 ;
        RECT 487.200 58.400 488.000 59.800 ;
        RECT 486.000 57.800 488.000 58.400 ;
        RECT 491.600 57.800 492.400 59.800 ;
        RECT 495.800 58.400 497.000 59.800 ;
        RECT 495.600 57.800 497.000 58.400 ;
        RECT 486.000 57.000 486.800 57.800 ;
        RECT 491.600 57.200 492.200 57.800 ;
        RECT 487.600 56.400 488.400 57.200 ;
        RECT 489.400 56.600 492.200 57.200 ;
        RECT 495.600 57.000 496.400 57.800 ;
        RECT 489.400 56.400 490.200 56.600 ;
        RECT 473.200 54.200 477.400 54.800 ;
        RECT 468.400 53.700 470.800 53.800 ;
        RECT 468.400 53.600 469.200 53.700 ;
        RECT 454.200 51.000 454.800 53.000 ;
        RECT 455.600 51.600 456.400 53.200 ;
        RECT 457.200 52.300 458.000 53.200 ;
        RECT 463.600 52.300 464.400 52.400 ;
        RECT 457.200 51.700 464.400 52.300 ;
        RECT 457.200 51.600 458.000 51.700 ;
        RECT 463.600 51.600 464.400 51.700 ;
        RECT 454.200 50.400 458.000 51.000 ;
        RECT 452.200 49.200 453.800 49.800 ;
        RECT 453.000 42.200 453.800 49.200 ;
        RECT 457.400 47.000 458.000 50.400 ;
        RECT 463.600 50.200 464.400 50.400 ;
        RECT 465.600 50.200 466.200 53.600 ;
        RECT 466.800 51.600 467.600 53.200 ;
        RECT 463.600 49.600 465.000 50.200 ;
        RECT 465.600 49.600 466.600 50.200 ;
        RECT 464.400 48.400 465.000 49.600 ;
        RECT 464.400 47.600 465.200 48.400 ;
        RECT 457.200 43.000 458.000 47.000 ;
        RECT 465.800 42.200 466.600 49.600 ;
        RECT 470.000 42.200 470.800 53.700 ;
        RECT 476.400 53.800 477.400 54.200 ;
        RECT 478.400 54.400 479.000 55.000 ;
        RECT 473.200 51.600 474.000 53.200 ;
        RECT 474.800 51.600 475.600 53.200 ;
        RECT 476.400 53.000 477.800 53.800 ;
        RECT 478.400 53.600 480.400 54.400 ;
        RECT 483.600 54.200 485.200 54.400 ;
        RECT 487.800 54.200 488.400 56.400 ;
        RECT 497.400 55.400 498.200 55.600 ;
        RECT 500.400 55.400 501.200 59.800 ;
        RECT 502.000 55.600 502.800 57.200 ;
        RECT 497.400 54.800 501.200 55.400 ;
        RECT 493.400 54.200 494.200 54.400 ;
        RECT 483.600 53.600 494.600 54.200 ;
        RECT 476.400 51.000 477.000 53.000 ;
        RECT 473.200 50.400 477.000 51.000 ;
        RECT 473.200 47.000 473.800 50.400 ;
        RECT 478.400 49.800 479.000 53.600 ;
        RECT 486.600 53.400 487.400 53.600 ;
        RECT 485.000 52.400 485.800 52.600 ;
        RECT 487.600 52.400 488.400 52.600 ;
        RECT 479.600 50.800 480.400 52.400 ;
        RECT 485.000 51.800 490.000 52.400 ;
        RECT 489.200 51.600 490.000 51.800 ;
        RECT 482.800 51.000 488.400 51.200 ;
        RECT 482.800 50.800 488.600 51.000 ;
        RECT 477.400 49.200 479.000 49.800 ;
        RECT 482.800 50.600 492.600 50.800 ;
        RECT 473.200 43.000 474.000 47.000 ;
        RECT 477.400 44.400 478.200 49.200 ;
        RECT 477.400 43.600 478.800 44.400 ;
        RECT 477.400 42.200 478.200 43.600 ;
        RECT 482.800 42.200 483.600 50.600 ;
        RECT 487.800 50.200 492.600 50.600 ;
        RECT 486.000 49.000 491.400 49.600 ;
        RECT 486.000 48.800 486.800 49.000 ;
        RECT 490.600 48.800 491.400 49.000 ;
        RECT 492.000 49.000 492.600 50.200 ;
        RECT 494.000 50.400 494.600 53.600 ;
        RECT 495.600 52.800 496.400 53.000 ;
        RECT 495.600 52.200 499.400 52.800 ;
        RECT 498.600 52.000 499.400 52.200 ;
        RECT 497.000 51.400 497.800 51.600 ;
        RECT 500.400 51.400 501.200 54.800 ;
        RECT 497.000 50.800 501.200 51.400 ;
        RECT 494.000 49.800 496.400 50.400 ;
        RECT 493.400 49.000 494.200 49.200 ;
        RECT 492.000 48.400 494.200 49.000 ;
        RECT 495.800 48.800 496.400 49.800 ;
        RECT 495.800 48.000 497.200 48.800 ;
        RECT 489.400 47.400 490.200 47.600 ;
        RECT 492.200 47.400 493.000 47.600 ;
        RECT 486.000 46.200 486.800 47.000 ;
        RECT 489.400 46.800 493.000 47.400 ;
        RECT 491.600 46.200 492.200 46.800 ;
        RECT 495.600 46.200 496.400 47.000 ;
        RECT 486.000 45.600 488.000 46.200 ;
        RECT 487.200 42.200 488.000 45.600 ;
        RECT 491.600 42.200 492.400 46.200 ;
        RECT 495.800 42.200 497.000 46.200 ;
        RECT 500.400 42.200 501.200 50.800 ;
        RECT 503.600 42.200 504.400 59.800 ;
        RECT 505.200 57.000 506.000 59.000 ;
        RECT 505.200 54.800 505.800 57.000 ;
        RECT 509.400 56.000 510.200 59.000 ;
        RECT 516.400 56.400 517.200 59.800 ;
        RECT 509.400 55.400 511.000 56.000 ;
        RECT 510.200 55.000 511.000 55.400 ;
        RECT 505.200 54.200 509.400 54.800 ;
        RECT 508.400 53.800 509.400 54.200 ;
        RECT 510.400 54.400 511.000 55.000 ;
        RECT 516.200 55.800 517.200 56.400 ;
        RECT 516.200 54.400 516.800 55.800 ;
        RECT 519.600 55.200 520.400 59.800 ;
        RECT 525.000 56.000 525.800 59.000 ;
        RECT 529.200 57.000 530.000 59.000 ;
        RECT 517.800 54.600 520.400 55.200 ;
        RECT 524.200 55.400 525.800 56.000 ;
        RECT 524.200 55.000 525.000 55.400 ;
        RECT 505.200 51.600 506.000 53.200 ;
        RECT 506.800 51.600 507.600 53.200 ;
        RECT 508.400 53.000 509.800 53.800 ;
        RECT 510.400 53.600 512.400 54.400 ;
        RECT 516.200 53.600 517.200 54.400 ;
        RECT 508.400 51.000 509.000 53.000 ;
        RECT 505.200 50.400 509.000 51.000 ;
        RECT 505.200 47.000 505.800 50.400 ;
        RECT 510.400 49.800 511.000 53.600 ;
        RECT 511.600 52.300 512.400 52.400 ;
        RECT 514.800 52.300 515.600 52.400 ;
        RECT 511.600 51.700 515.600 52.300 ;
        RECT 511.600 50.800 512.400 51.700 ;
        RECT 514.800 51.600 515.600 51.700 ;
        RECT 509.400 49.200 511.000 49.800 ;
        RECT 516.200 50.200 516.800 53.600 ;
        RECT 517.800 53.000 518.400 54.600 ;
        RECT 524.200 54.400 524.800 55.000 ;
        RECT 529.400 54.800 530.000 57.000 ;
        RECT 530.800 56.000 531.600 59.800 ;
        RECT 534.000 56.000 534.800 59.800 ;
        RECT 530.800 55.800 534.800 56.000 ;
        RECT 535.600 55.800 536.400 59.800 ;
        RECT 537.200 55.800 538.000 59.800 ;
        RECT 538.800 56.000 539.600 59.800 ;
        RECT 542.000 56.000 542.800 59.800 ;
        RECT 538.800 55.800 542.800 56.000 ;
        RECT 531.000 55.400 534.600 55.800 ;
        RECT 522.800 53.600 524.800 54.400 ;
        RECT 525.800 54.200 530.000 54.800 ;
        RECT 531.600 54.400 532.400 54.800 ;
        RECT 535.600 54.400 536.200 55.800 ;
        RECT 537.400 54.400 538.000 55.800 ;
        RECT 539.000 55.400 542.600 55.800 ;
        RECT 543.600 55.400 544.400 59.800 ;
        RECT 547.800 58.400 549.000 59.800 ;
        RECT 547.800 57.800 549.200 58.400 ;
        RECT 552.400 57.800 553.200 59.800 ;
        RECT 556.800 58.400 557.600 59.800 ;
        RECT 556.800 57.800 558.800 58.400 ;
        RECT 548.400 57.000 549.200 57.800 ;
        RECT 552.600 57.200 553.200 57.800 ;
        RECT 552.600 56.600 555.400 57.200 ;
        RECT 554.600 56.400 555.400 56.600 ;
        RECT 556.400 56.400 557.200 57.200 ;
        RECT 558.000 57.000 558.800 57.800 ;
        RECT 546.600 55.400 547.400 55.600 ;
        RECT 543.600 54.800 547.400 55.400 ;
        RECT 541.200 54.400 542.000 54.800 ;
        RECT 525.800 53.800 526.800 54.200 ;
        RECT 517.400 52.200 518.400 53.000 ;
        RECT 517.800 50.200 518.400 52.200 ;
        RECT 519.400 52.400 520.200 53.200 ;
        RECT 519.400 52.300 520.400 52.400 ;
        RECT 521.200 52.300 522.000 52.400 ;
        RECT 519.400 51.700 522.000 52.300 ;
        RECT 519.400 51.600 520.400 51.700 ;
        RECT 521.200 51.600 522.000 51.700 ;
        RECT 522.800 50.800 523.600 52.400 ;
        RECT 524.200 50.400 524.800 53.600 ;
        RECT 525.400 53.000 526.800 53.800 ;
        RECT 530.800 53.800 532.400 54.400 ;
        RECT 530.800 53.600 531.600 53.800 ;
        RECT 533.800 53.600 536.400 54.400 ;
        RECT 537.200 53.600 539.800 54.400 ;
        RECT 541.200 53.800 542.800 54.400 ;
        RECT 542.000 53.600 542.800 53.800 ;
        RECT 526.200 51.000 526.800 53.000 ;
        RECT 527.600 51.600 528.400 53.200 ;
        RECT 529.200 51.600 530.000 53.200 ;
        RECT 532.400 51.600 533.200 53.200 ;
        RECT 533.800 52.300 534.400 53.600 ;
        RECT 533.800 51.700 537.900 52.300 ;
        RECT 526.200 50.400 530.000 51.000 ;
        RECT 516.200 49.200 517.200 50.200 ;
        RECT 517.800 49.600 520.400 50.200 ;
        RECT 505.200 43.000 506.000 47.000 ;
        RECT 509.400 44.400 510.200 49.200 ;
        RECT 509.400 43.600 510.800 44.400 ;
        RECT 509.400 42.200 510.200 43.600 ;
        RECT 516.400 42.200 517.200 49.200 ;
        RECT 519.600 42.200 520.400 49.600 ;
        RECT 524.200 49.800 525.200 50.400 ;
        RECT 524.200 49.200 525.800 49.800 ;
        RECT 525.000 42.200 525.800 49.200 ;
        RECT 529.400 47.000 530.000 50.400 ;
        RECT 533.800 50.200 534.400 51.700 ;
        RECT 537.300 50.400 537.900 51.700 ;
        RECT 535.600 50.200 536.400 50.400 ;
        RECT 529.200 43.000 530.000 47.000 ;
        RECT 533.400 49.600 534.400 50.200 ;
        RECT 535.000 49.600 536.400 50.200 ;
        RECT 537.200 50.200 538.000 50.400 ;
        RECT 539.200 50.200 539.800 53.600 ;
        RECT 540.400 51.600 541.200 53.200 ;
        RECT 543.600 51.400 544.400 54.800 ;
        RECT 550.600 54.200 551.400 54.400 ;
        RECT 556.400 54.200 557.000 56.400 ;
        RECT 561.200 55.000 562.000 59.800 ;
        RECT 564.400 55.200 565.200 59.800 ;
        RECT 567.600 55.200 568.400 59.800 ;
        RECT 570.800 55.200 571.600 59.800 ;
        RECT 574.000 55.200 574.800 59.800 ;
        RECT 578.800 56.000 579.600 59.800 ;
        RECT 562.800 54.400 565.200 55.200 ;
        RECT 566.200 54.400 568.400 55.200 ;
        RECT 569.400 54.400 571.600 55.200 ;
        RECT 573.000 54.400 574.800 55.200 ;
        RECT 578.600 55.200 579.600 56.000 ;
        RECT 559.600 54.200 561.200 54.400 ;
        RECT 550.200 53.600 561.200 54.200 ;
        RECT 548.400 52.800 549.200 53.000 ;
        RECT 545.400 52.200 549.200 52.800 ;
        RECT 550.200 52.400 550.800 53.600 ;
        RECT 557.400 53.400 558.200 53.600 ;
        RECT 559.000 52.400 559.800 52.600 ;
        RECT 545.400 52.000 546.200 52.200 ;
        RECT 550.000 51.600 550.800 52.400 ;
        RECT 551.600 52.300 552.400 52.400 ;
        RECT 554.800 52.300 559.800 52.400 ;
        RECT 551.600 51.800 559.800 52.300 ;
        RECT 551.600 51.700 555.600 51.800 ;
        RECT 551.600 51.600 552.400 51.700 ;
        RECT 554.800 51.600 555.600 51.700 ;
        RECT 562.800 51.600 563.600 54.400 ;
        RECT 566.200 53.800 567.000 54.400 ;
        RECT 569.400 53.800 570.200 54.400 ;
        RECT 573.000 53.800 573.800 54.400 ;
        RECT 575.600 53.800 576.400 54.400 ;
        RECT 564.400 53.000 567.000 53.800 ;
        RECT 567.800 53.000 570.200 53.800 ;
        RECT 571.200 53.000 573.800 53.800 ;
        RECT 574.600 53.000 576.400 53.800 ;
        RECT 566.200 51.600 567.000 53.000 ;
        RECT 569.400 51.600 570.200 53.000 ;
        RECT 573.000 51.600 573.800 53.000 ;
        RECT 547.000 51.400 547.800 51.600 ;
        RECT 543.600 50.800 547.800 51.400 ;
        RECT 537.200 49.600 538.600 50.200 ;
        RECT 539.200 49.600 540.200 50.200 ;
        RECT 533.400 42.200 534.200 49.600 ;
        RECT 535.000 48.400 535.600 49.600 ;
        RECT 534.800 47.600 535.600 48.400 ;
        RECT 538.000 48.400 538.600 49.600 ;
        RECT 539.400 48.400 540.200 49.600 ;
        RECT 538.000 47.600 538.800 48.400 ;
        RECT 539.400 47.600 541.200 48.400 ;
        RECT 539.400 42.200 540.200 47.600 ;
        RECT 543.600 42.200 544.400 50.800 ;
        RECT 550.200 50.400 550.800 51.600 ;
        RECT 556.400 51.000 562.000 51.200 ;
        RECT 556.200 50.800 562.000 51.000 ;
        RECT 562.800 50.800 565.200 51.600 ;
        RECT 566.200 50.800 568.400 51.600 ;
        RECT 569.400 50.800 571.600 51.600 ;
        RECT 573.000 50.800 574.800 51.600 ;
        RECT 548.400 49.800 550.800 50.400 ;
        RECT 552.200 50.600 562.000 50.800 ;
        RECT 552.200 50.200 557.000 50.600 ;
        RECT 548.400 48.800 549.000 49.800 ;
        RECT 547.600 48.000 549.000 48.800 ;
        RECT 550.600 49.000 551.400 49.200 ;
        RECT 552.200 49.000 552.800 50.200 ;
        RECT 550.600 48.400 552.800 49.000 ;
        RECT 553.400 49.000 558.800 49.600 ;
        RECT 553.400 48.800 554.200 49.000 ;
        RECT 558.000 48.800 558.800 49.000 ;
        RECT 551.800 47.400 552.600 47.600 ;
        RECT 554.600 47.400 555.400 47.600 ;
        RECT 548.400 46.200 549.200 47.000 ;
        RECT 551.800 46.800 555.400 47.400 ;
        RECT 552.600 46.200 553.200 46.800 ;
        RECT 558.000 46.200 558.800 47.000 ;
        RECT 547.800 42.200 549.000 46.200 ;
        RECT 552.400 42.200 553.200 46.200 ;
        RECT 556.800 45.600 558.800 46.200 ;
        RECT 556.800 42.200 557.600 45.600 ;
        RECT 561.200 42.200 562.000 50.600 ;
        RECT 564.400 42.200 565.200 50.800 ;
        RECT 567.600 42.200 568.400 50.800 ;
        RECT 570.800 42.200 571.600 50.800 ;
        RECT 574.000 42.200 574.800 50.800 ;
        RECT 578.600 50.800 579.400 55.200 ;
        RECT 580.400 54.600 581.200 59.800 ;
        RECT 586.800 56.600 587.600 59.800 ;
        RECT 588.400 57.000 589.200 59.800 ;
        RECT 590.000 57.000 590.800 59.800 ;
        RECT 591.600 57.000 592.400 59.800 ;
        RECT 593.200 57.000 594.000 59.800 ;
        RECT 596.400 57.000 597.200 59.800 ;
        RECT 599.600 57.000 600.400 59.800 ;
        RECT 601.200 57.000 602.000 59.800 ;
        RECT 602.800 57.000 603.600 59.800 ;
        RECT 585.200 55.800 587.600 56.600 ;
        RECT 604.400 56.600 605.200 59.800 ;
        RECT 585.200 55.200 586.000 55.800 ;
        RECT 580.000 54.000 581.200 54.600 ;
        RECT 584.200 54.600 586.000 55.200 ;
        RECT 590.000 55.600 591.000 56.400 ;
        RECT 594.000 55.600 595.600 56.400 ;
        RECT 596.400 55.800 601.000 56.400 ;
        RECT 604.400 55.800 607.000 56.600 ;
        RECT 596.400 55.600 597.200 55.800 ;
        RECT 580.000 52.000 580.600 54.000 ;
        RECT 584.200 53.400 585.000 54.600 ;
        RECT 581.200 52.600 585.000 53.400 ;
        RECT 590.000 52.800 590.800 55.600 ;
        RECT 596.400 54.800 597.200 55.000 ;
        RECT 592.800 54.200 597.200 54.800 ;
        RECT 592.800 54.000 593.600 54.200 ;
        RECT 598.000 53.600 598.800 55.200 ;
        RECT 600.200 53.400 601.000 55.800 ;
        RECT 606.200 55.200 607.000 55.800 ;
        RECT 606.200 54.400 609.200 55.200 ;
        RECT 610.800 53.800 611.600 59.800 ;
        RECT 593.200 52.600 596.400 53.400 ;
        RECT 600.200 52.600 602.200 53.400 ;
        RECT 602.800 53.000 611.600 53.800 ;
        RECT 586.800 52.000 587.600 52.600 ;
        RECT 598.000 52.000 598.800 52.400 ;
        RECT 604.400 52.000 605.200 52.400 ;
        RECT 609.400 52.000 610.200 52.200 ;
        RECT 580.000 51.400 580.800 52.000 ;
        RECT 586.800 51.400 610.200 52.000 ;
        RECT 578.600 50.000 579.600 50.800 ;
        RECT 578.800 42.200 579.600 50.000 ;
        RECT 580.200 49.600 580.800 51.400 ;
        RECT 580.200 49.000 589.200 49.600 ;
        RECT 580.200 47.400 580.800 49.000 ;
        RECT 588.400 48.800 589.200 49.000 ;
        RECT 591.600 49.000 600.200 49.600 ;
        RECT 591.600 48.800 592.400 49.000 ;
        RECT 583.400 47.600 586.000 48.400 ;
        RECT 580.200 46.800 582.800 47.400 ;
        RECT 582.000 42.200 582.800 46.800 ;
        RECT 585.200 42.200 586.000 47.600 ;
        RECT 586.600 46.800 590.800 47.600 ;
        RECT 588.400 42.200 589.200 45.000 ;
        RECT 590.000 42.200 590.800 45.000 ;
        RECT 591.600 42.200 592.400 45.000 ;
        RECT 593.200 42.200 594.000 48.400 ;
        RECT 596.400 47.600 599.000 48.400 ;
        RECT 599.600 48.200 600.200 49.000 ;
        RECT 601.200 49.400 602.000 49.600 ;
        RECT 601.200 49.000 606.600 49.400 ;
        RECT 601.200 48.800 607.400 49.000 ;
        RECT 606.000 48.200 607.400 48.800 ;
        RECT 599.600 47.600 605.400 48.200 ;
        RECT 608.400 48.000 610.000 48.800 ;
        RECT 608.400 47.600 609.000 48.000 ;
        RECT 596.400 42.200 597.200 47.000 ;
        RECT 599.600 42.200 600.400 47.000 ;
        RECT 604.800 46.800 609.000 47.600 ;
        RECT 610.800 47.400 611.600 53.000 ;
        RECT 609.600 46.800 611.600 47.400 ;
        RECT 601.200 42.200 602.000 45.000 ;
        RECT 602.800 42.200 603.600 45.000 ;
        RECT 606.000 42.200 606.800 46.800 ;
        RECT 609.600 46.200 610.200 46.800 ;
        RECT 609.200 45.600 610.200 46.200 ;
        RECT 609.200 42.200 610.000 45.600 ;
        RECT 4.400 32.400 5.200 39.800 ;
        RECT 7.600 36.400 8.400 39.800 ;
        RECT 7.400 35.800 8.400 36.400 ;
        RECT 7.400 35.200 8.000 35.800 ;
        RECT 10.800 35.200 11.600 39.800 ;
        RECT 14.000 37.000 14.800 39.800 ;
        RECT 15.600 37.000 16.400 39.800 ;
        RECT 3.000 31.800 5.200 32.400 ;
        RECT 6.000 34.600 8.000 35.200 ;
        RECT 3.000 31.200 3.600 31.800 ;
        RECT 2.400 30.400 3.600 31.200 ;
        RECT 3.000 27.400 3.600 30.400 ;
        RECT 4.400 28.800 5.200 30.400 ;
        RECT 6.000 29.000 6.800 34.600 ;
        RECT 8.600 34.400 12.800 35.200 ;
        RECT 17.200 35.000 18.000 39.800 ;
        RECT 20.400 35.000 21.200 39.800 ;
        RECT 8.600 34.000 9.200 34.400 ;
        RECT 7.600 33.200 9.200 34.000 ;
        RECT 12.200 33.800 18.000 34.400 ;
        RECT 10.200 33.200 11.600 33.800 ;
        RECT 10.200 33.000 16.400 33.200 ;
        RECT 11.000 32.600 16.400 33.000 ;
        RECT 15.600 32.400 16.400 32.600 ;
        RECT 17.400 33.000 18.000 33.800 ;
        RECT 18.600 33.600 21.200 34.400 ;
        RECT 23.600 33.600 24.400 39.800 ;
        RECT 25.200 37.000 26.000 39.800 ;
        RECT 26.800 37.000 27.600 39.800 ;
        RECT 28.400 37.000 29.200 39.800 ;
        RECT 26.800 34.400 31.000 35.200 ;
        RECT 31.600 34.400 32.400 39.800 ;
        RECT 34.800 35.200 35.600 39.800 ;
        RECT 34.800 34.600 37.400 35.200 ;
        RECT 31.600 33.600 34.200 34.400 ;
        RECT 25.200 33.000 26.000 33.200 ;
        RECT 17.400 32.400 26.000 33.000 ;
        RECT 28.400 33.000 29.200 33.200 ;
        RECT 36.800 33.000 37.400 34.600 ;
        RECT 28.400 32.400 37.400 33.000 ;
        RECT 36.800 30.600 37.400 32.400 ;
        RECT 38.000 32.000 38.800 39.800 ;
        RECT 42.000 33.600 42.800 34.400 ;
        RECT 42.000 32.400 42.600 33.600 ;
        RECT 43.400 32.400 44.200 39.800 ;
        RECT 38.000 31.200 39.000 32.000 ;
        RECT 41.200 31.800 42.600 32.400 ;
        RECT 43.200 31.800 44.200 32.400 ;
        RECT 41.200 31.600 42.000 31.800 ;
        RECT 7.400 30.000 30.800 30.600 ;
        RECT 36.800 30.000 37.600 30.600 ;
        RECT 7.400 29.800 8.200 30.000 ;
        RECT 9.200 29.600 10.000 30.000 ;
        RECT 12.400 29.600 13.200 30.000 ;
        RECT 30.000 29.400 30.800 30.000 ;
        RECT 6.000 28.200 14.800 29.000 ;
        RECT 15.400 28.600 17.400 29.400 ;
        RECT 21.200 28.600 24.400 29.400 ;
        RECT 3.000 26.800 5.200 27.400 ;
        RECT 4.400 22.200 5.200 26.800 ;
        RECT 6.000 22.200 6.800 28.200 ;
        RECT 8.400 26.800 11.400 27.600 ;
        RECT 10.600 26.200 11.400 26.800 ;
        RECT 16.600 26.200 17.400 28.600 ;
        RECT 18.800 26.800 19.600 28.400 ;
        RECT 24.000 27.800 24.800 28.000 ;
        RECT 20.400 27.200 24.800 27.800 ;
        RECT 20.400 27.000 21.200 27.200 ;
        RECT 26.800 26.400 27.600 29.200 ;
        RECT 32.600 28.600 36.400 29.400 ;
        RECT 32.600 27.400 33.400 28.600 ;
        RECT 37.000 28.000 37.600 30.000 ;
        RECT 20.400 26.200 21.200 26.400 ;
        RECT 10.600 25.400 13.200 26.200 ;
        RECT 16.600 25.600 21.200 26.200 ;
        RECT 22.000 25.600 23.600 26.400 ;
        RECT 26.600 25.600 27.600 26.400 ;
        RECT 31.600 26.800 33.400 27.400 ;
        RECT 36.400 27.400 37.600 28.000 ;
        RECT 31.600 26.200 32.400 26.800 ;
        RECT 12.400 22.200 13.200 25.400 ;
        RECT 30.000 25.400 32.400 26.200 ;
        RECT 14.000 22.200 14.800 25.000 ;
        RECT 15.600 22.200 16.400 25.000 ;
        RECT 17.200 22.200 18.000 25.000 ;
        RECT 20.400 22.200 21.200 25.000 ;
        RECT 23.600 22.200 24.400 25.000 ;
        RECT 25.200 22.200 26.000 25.000 ;
        RECT 26.800 22.200 27.600 25.000 ;
        RECT 28.400 22.200 29.200 25.000 ;
        RECT 30.000 22.200 30.800 25.400 ;
        RECT 36.400 22.200 37.200 27.400 ;
        RECT 38.200 26.800 39.000 31.200 ;
        RECT 43.200 28.400 43.800 31.800 ;
        RECT 44.400 28.800 45.200 30.400 ;
        RECT 39.600 28.300 40.400 28.400 ;
        RECT 41.200 28.300 43.800 28.400 ;
        RECT 39.600 27.700 43.800 28.300 ;
        RECT 46.000 28.300 46.800 28.400 ;
        RECT 47.600 28.300 48.400 39.800 ;
        RECT 53.400 32.400 54.200 39.800 ;
        RECT 54.800 33.600 55.600 34.400 ;
        RECT 55.000 32.400 55.600 33.600 ;
        RECT 58.000 33.600 58.800 34.400 ;
        RECT 58.000 32.400 58.600 33.600 ;
        RECT 59.400 32.400 60.200 39.800 ;
        RECT 53.400 31.800 54.400 32.400 ;
        RECT 55.000 31.800 56.400 32.400 ;
        RECT 52.400 28.800 53.200 30.400 ;
        RECT 53.800 30.300 54.400 31.800 ;
        RECT 55.600 31.600 56.400 31.800 ;
        RECT 57.200 31.800 58.600 32.400 ;
        RECT 59.200 31.800 60.200 32.400 ;
        RECT 57.200 31.600 58.000 31.800 ;
        RECT 57.300 30.300 57.900 31.600 ;
        RECT 53.800 29.700 57.900 30.300 ;
        RECT 53.800 28.400 54.400 29.700 ;
        RECT 59.200 28.400 59.800 31.800 ;
        RECT 63.600 31.200 64.400 39.800 ;
        RECT 67.800 35.800 69.000 39.800 ;
        RECT 72.400 35.800 73.200 39.800 ;
        RECT 76.800 36.400 77.600 39.800 ;
        RECT 76.800 35.800 78.800 36.400 ;
        RECT 68.400 35.000 69.200 35.800 ;
        RECT 72.600 35.200 73.200 35.800 ;
        RECT 71.800 34.600 75.400 35.200 ;
        RECT 78.000 35.000 78.800 35.800 ;
        RECT 71.800 34.400 72.600 34.600 ;
        RECT 74.600 34.400 75.400 34.600 ;
        RECT 67.600 33.200 69.000 34.000 ;
        RECT 68.400 32.200 69.000 33.200 ;
        RECT 70.600 33.000 72.800 33.600 ;
        RECT 70.600 32.800 71.400 33.000 ;
        RECT 68.400 31.600 70.800 32.200 ;
        RECT 63.600 30.600 67.800 31.200 ;
        RECT 60.400 28.800 61.200 30.400 ;
        RECT 46.000 28.200 48.400 28.300 ;
        RECT 39.600 27.600 40.400 27.700 ;
        RECT 41.200 27.600 43.800 27.700 ;
        RECT 45.200 27.700 48.400 28.200 ;
        RECT 45.200 27.600 46.800 27.700 ;
        RECT 38.000 26.000 39.000 26.800 ;
        RECT 41.400 26.200 42.000 27.600 ;
        RECT 45.200 27.200 46.000 27.600 ;
        RECT 43.000 26.200 46.600 26.600 ;
        RECT 38.000 22.200 38.800 26.000 ;
        RECT 41.200 22.200 42.000 26.200 ;
        RECT 42.800 26.000 46.800 26.200 ;
        RECT 42.800 22.200 43.600 26.000 ;
        RECT 46.000 22.200 46.800 26.000 ;
        RECT 47.600 22.200 48.400 27.700 ;
        RECT 50.800 28.200 51.600 28.400 ;
        RECT 50.800 27.600 52.400 28.200 ;
        RECT 53.800 27.600 56.400 28.400 ;
        RECT 57.200 27.600 59.800 28.400 ;
        RECT 62.000 28.200 62.800 28.400 ;
        RECT 61.200 27.600 62.800 28.200 ;
        RECT 51.600 27.200 52.400 27.600 ;
        RECT 51.000 26.200 54.600 26.600 ;
        RECT 55.600 26.200 56.200 27.600 ;
        RECT 57.400 26.200 58.000 27.600 ;
        RECT 61.200 27.200 62.000 27.600 ;
        RECT 63.600 27.200 64.400 30.600 ;
        RECT 67.000 30.400 67.800 30.600 ;
        RECT 65.400 29.800 66.200 30.000 ;
        RECT 65.400 29.200 69.200 29.800 ;
        RECT 68.400 29.000 69.200 29.200 ;
        RECT 70.200 28.400 70.800 31.600 ;
        RECT 72.200 31.800 72.800 33.000 ;
        RECT 73.400 33.000 74.200 33.200 ;
        RECT 78.000 33.000 78.800 33.200 ;
        RECT 73.400 32.400 78.800 33.000 ;
        RECT 72.200 31.400 77.000 31.800 ;
        RECT 81.200 31.400 82.000 39.800 ;
        RECT 85.400 32.400 86.200 39.800 ;
        RECT 86.800 33.600 87.600 34.400 ;
        RECT 87.000 32.400 87.600 33.600 ;
        RECT 90.000 33.600 90.800 34.400 ;
        RECT 90.000 32.400 90.600 33.600 ;
        RECT 91.400 32.400 92.200 39.800 ;
        RECT 84.400 31.600 86.400 32.400 ;
        RECT 87.000 31.800 88.400 32.400 ;
        RECT 87.600 31.600 88.400 31.800 ;
        RECT 89.200 31.800 90.600 32.400 ;
        RECT 91.200 31.800 92.200 32.400 ;
        RECT 89.200 31.600 90.000 31.800 ;
        RECT 72.200 31.200 82.000 31.400 ;
        RECT 76.200 31.000 82.000 31.200 ;
        RECT 76.400 30.800 82.000 31.000 ;
        RECT 74.800 30.200 75.600 30.400 ;
        RECT 74.800 29.600 79.800 30.200 ;
        RECT 76.400 29.400 77.200 29.600 ;
        RECT 79.000 29.400 79.800 29.600 ;
        RECT 84.400 28.800 85.200 30.400 ;
        RECT 77.400 28.400 78.200 28.600 ;
        RECT 85.800 28.400 86.400 31.600 ;
        RECT 87.700 30.300 88.300 31.600 ;
        RECT 91.200 30.300 91.800 31.800 ;
        RECT 95.600 31.400 96.400 39.800 ;
        RECT 100.000 36.400 100.800 39.800 ;
        RECT 98.800 35.800 100.800 36.400 ;
        RECT 104.400 35.800 105.200 39.800 ;
        RECT 108.600 35.800 109.800 39.800 ;
        RECT 98.800 35.000 99.600 35.800 ;
        RECT 104.400 35.200 105.000 35.800 ;
        RECT 102.200 34.600 105.800 35.200 ;
        RECT 108.400 35.000 109.200 35.800 ;
        RECT 102.200 34.400 103.000 34.600 ;
        RECT 105.000 34.400 105.800 34.600 ;
        RECT 98.800 33.000 99.600 33.200 ;
        RECT 103.400 33.000 104.200 33.200 ;
        RECT 98.800 32.400 104.200 33.000 ;
        RECT 104.800 33.000 107.000 33.600 ;
        RECT 104.800 31.800 105.400 33.000 ;
        RECT 106.200 32.800 107.000 33.000 ;
        RECT 108.600 33.200 110.000 34.000 ;
        RECT 108.600 32.200 109.200 33.200 ;
        RECT 100.600 31.400 105.400 31.800 ;
        RECT 95.600 31.200 105.400 31.400 ;
        RECT 106.800 31.600 109.200 32.200 ;
        RECT 95.600 31.000 101.400 31.200 ;
        RECT 95.600 30.800 101.200 31.000 ;
        RECT 87.700 29.700 91.800 30.300 ;
        RECT 91.200 28.400 91.800 29.700 ;
        RECT 92.400 28.800 93.200 30.400 ;
        RECT 102.000 30.200 102.800 30.400 ;
        RECT 97.800 29.600 102.800 30.200 ;
        RECT 97.800 29.400 98.600 29.600 ;
        RECT 99.400 28.400 100.200 28.600 ;
        RECT 106.800 28.400 107.400 31.600 ;
        RECT 113.200 31.200 114.000 39.800 ;
        RECT 117.400 32.400 118.200 39.800 ;
        RECT 118.800 33.600 119.600 34.400 ;
        RECT 119.000 32.400 119.600 33.600 ;
        RECT 122.000 33.600 122.800 34.400 ;
        RECT 122.000 32.400 122.600 33.600 ;
        RECT 123.400 32.400 124.200 39.800 ;
        RECT 116.400 31.600 118.400 32.400 ;
        RECT 119.000 31.800 120.400 32.400 ;
        RECT 119.600 31.600 120.400 31.800 ;
        RECT 121.200 31.800 122.600 32.400 ;
        RECT 123.200 31.800 124.200 32.400 ;
        RECT 130.200 32.400 131.000 39.800 ;
        RECT 131.600 33.600 132.400 34.400 ;
        RECT 131.800 32.400 132.400 33.600 ;
        RECT 134.800 33.600 135.600 34.400 ;
        RECT 134.800 32.400 135.400 33.600 ;
        RECT 136.200 32.400 137.000 39.800 ;
        RECT 130.200 31.800 131.200 32.400 ;
        RECT 131.800 31.800 133.200 32.400 ;
        RECT 121.200 31.600 122.000 31.800 ;
        RECT 109.800 30.600 114.000 31.200 ;
        RECT 109.800 30.400 110.600 30.600 ;
        RECT 111.400 29.800 112.200 30.000 ;
        RECT 108.400 29.200 112.200 29.800 ;
        RECT 108.400 29.000 109.200 29.200 ;
        RECT 70.200 27.800 81.200 28.400 ;
        RECT 70.600 27.600 71.400 27.800 ;
        RECT 63.600 26.600 67.400 27.200 ;
        RECT 59.000 26.200 62.600 26.600 ;
        RECT 50.800 26.000 54.800 26.200 ;
        RECT 50.800 22.200 51.600 26.000 ;
        RECT 54.000 22.200 54.800 26.000 ;
        RECT 55.600 22.200 56.400 26.200 ;
        RECT 57.200 22.200 58.000 26.200 ;
        RECT 58.800 26.000 62.800 26.200 ;
        RECT 58.800 22.200 59.600 26.000 ;
        RECT 62.000 22.200 62.800 26.000 ;
        RECT 63.600 22.200 64.400 26.600 ;
        RECT 66.600 26.400 67.400 26.600 ;
        RECT 76.400 26.400 77.000 27.800 ;
        RECT 79.600 27.600 81.200 27.800 ;
        RECT 82.800 28.200 83.600 28.400 ;
        RECT 82.800 27.600 84.400 28.200 ;
        RECT 85.800 27.600 88.400 28.400 ;
        RECT 89.200 27.600 91.800 28.400 ;
        RECT 94.000 28.200 94.800 28.400 ;
        RECT 93.200 27.600 94.800 28.200 ;
        RECT 96.400 27.800 107.400 28.400 ;
        RECT 96.400 27.600 98.000 27.800 ;
        RECT 100.400 27.600 101.200 27.800 ;
        RECT 106.200 27.600 107.000 27.800 ;
        RECT 83.600 27.200 84.400 27.600 ;
        RECT 74.600 25.400 75.400 25.600 ;
        RECT 68.400 24.200 69.200 25.000 ;
        RECT 72.600 24.800 75.400 25.400 ;
        RECT 76.400 24.800 77.200 26.400 ;
        RECT 72.600 24.200 73.200 24.800 ;
        RECT 78.000 24.200 78.800 25.000 ;
        RECT 67.800 23.600 69.200 24.200 ;
        RECT 67.800 22.200 69.000 23.600 ;
        RECT 72.400 22.200 73.200 24.200 ;
        RECT 76.800 23.600 78.800 24.200 ;
        RECT 76.800 22.200 77.600 23.600 ;
        RECT 81.200 22.200 82.000 27.000 ;
        RECT 83.000 26.200 86.600 26.600 ;
        RECT 87.600 26.200 88.200 27.600 ;
        RECT 89.400 26.200 90.000 27.600 ;
        RECT 93.200 27.200 94.000 27.600 ;
        RECT 91.000 26.200 94.600 26.600 ;
        RECT 82.800 26.000 86.800 26.200 ;
        RECT 82.800 22.200 83.600 26.000 ;
        RECT 86.000 22.200 86.800 26.000 ;
        RECT 87.600 22.200 88.400 26.200 ;
        RECT 89.200 22.200 90.000 26.200 ;
        RECT 90.800 26.000 94.800 26.200 ;
        RECT 90.800 22.200 91.600 26.000 ;
        RECT 94.000 22.200 94.800 26.000 ;
        RECT 95.600 22.200 96.400 27.000 ;
        RECT 100.600 25.600 101.200 27.600 ;
        RECT 113.200 27.200 114.000 30.600 ;
        RECT 116.400 28.800 117.200 30.400 ;
        RECT 117.800 28.400 118.400 31.600 ;
        RECT 119.700 30.300 120.300 31.600 ;
        RECT 123.200 30.300 123.800 31.800 ;
        RECT 119.700 29.700 123.800 30.300 ;
        RECT 123.200 28.400 123.800 29.700 ;
        RECT 124.400 28.800 125.200 30.400 ;
        RECT 126.000 30.300 126.800 30.400 ;
        RECT 129.200 30.300 130.000 30.400 ;
        RECT 126.000 29.700 130.000 30.300 ;
        RECT 126.000 29.600 126.800 29.700 ;
        RECT 129.200 28.800 130.000 29.700 ;
        RECT 130.600 28.400 131.200 31.800 ;
        RECT 132.400 31.600 133.200 31.800 ;
        RECT 134.000 31.800 135.400 32.400 ;
        RECT 136.000 31.800 137.000 32.400 ;
        RECT 134.000 31.600 134.800 31.800 ;
        RECT 132.500 30.300 133.100 31.600 ;
        RECT 136.000 30.300 136.600 31.800 ;
        RECT 140.400 31.200 141.200 39.800 ;
        RECT 144.600 35.800 145.800 39.800 ;
        RECT 149.200 35.800 150.000 39.800 ;
        RECT 153.600 36.400 154.400 39.800 ;
        RECT 153.600 35.800 155.600 36.400 ;
        RECT 145.200 35.000 146.000 35.800 ;
        RECT 149.400 35.200 150.000 35.800 ;
        RECT 148.600 34.600 152.200 35.200 ;
        RECT 154.800 35.000 155.600 35.800 ;
        RECT 148.600 34.400 149.400 34.600 ;
        RECT 151.400 34.400 152.200 34.600 ;
        RECT 144.400 33.200 145.800 34.000 ;
        RECT 145.200 32.200 145.800 33.200 ;
        RECT 147.400 33.000 149.600 33.600 ;
        RECT 147.400 32.800 148.200 33.000 ;
        RECT 145.200 31.600 147.600 32.200 ;
        RECT 140.400 30.600 144.600 31.200 ;
        RECT 132.500 29.700 136.600 30.300 ;
        RECT 136.000 28.400 136.600 29.700 ;
        RECT 137.200 28.800 138.000 30.400 ;
        RECT 114.800 28.200 115.600 28.400 ;
        RECT 114.800 27.600 116.400 28.200 ;
        RECT 117.800 27.600 120.400 28.400 ;
        RECT 121.200 27.600 123.800 28.400 ;
        RECT 126.000 28.200 126.800 28.400 ;
        RECT 125.200 27.600 126.800 28.200 ;
        RECT 127.600 28.200 128.400 28.400 ;
        RECT 127.600 27.600 129.200 28.200 ;
        RECT 130.600 27.600 133.200 28.400 ;
        RECT 134.000 27.600 136.600 28.400 ;
        RECT 138.800 28.200 139.600 28.400 ;
        RECT 138.000 27.600 139.600 28.200 ;
        RECT 115.600 27.200 116.400 27.600 ;
        RECT 110.200 26.600 114.000 27.200 ;
        RECT 110.200 26.400 111.000 26.600 ;
        RECT 98.800 24.200 99.600 25.000 ;
        RECT 100.400 24.800 101.200 25.600 ;
        RECT 102.200 25.400 103.000 25.600 ;
        RECT 102.200 24.800 105.000 25.400 ;
        RECT 104.400 24.200 105.000 24.800 ;
        RECT 108.400 24.200 109.200 25.000 ;
        RECT 98.800 23.600 100.800 24.200 ;
        RECT 100.000 22.200 100.800 23.600 ;
        RECT 104.400 22.200 105.200 24.200 ;
        RECT 108.400 23.600 109.800 24.200 ;
        RECT 108.600 22.200 109.800 23.600 ;
        RECT 113.200 22.200 114.000 26.600 ;
        RECT 115.000 26.200 118.600 26.600 ;
        RECT 119.600 26.200 120.200 27.600 ;
        RECT 121.400 26.200 122.000 27.600 ;
        RECT 125.200 27.200 126.000 27.600 ;
        RECT 128.400 27.200 129.200 27.600 ;
        RECT 123.000 26.200 126.600 26.600 ;
        RECT 127.800 26.200 131.400 26.600 ;
        RECT 132.400 26.200 133.000 27.600 ;
        RECT 134.200 26.200 134.800 27.600 ;
        RECT 138.000 27.200 138.800 27.600 ;
        RECT 140.400 27.200 141.200 30.600 ;
        RECT 143.800 30.400 144.600 30.600 ;
        RECT 147.000 30.400 147.600 31.600 ;
        RECT 149.000 31.800 149.600 33.000 ;
        RECT 150.200 33.000 151.000 33.200 ;
        RECT 154.800 33.000 155.600 33.200 ;
        RECT 150.200 32.400 155.600 33.000 ;
        RECT 149.000 31.400 153.800 31.800 ;
        RECT 158.000 31.400 158.800 39.800 ;
        RECT 149.000 31.200 158.800 31.400 ;
        RECT 153.000 31.000 158.800 31.200 ;
        RECT 153.200 30.800 158.800 31.000 ;
        RECT 142.200 29.800 143.000 30.000 ;
        RECT 142.200 29.200 146.000 29.800 ;
        RECT 146.800 29.600 147.600 30.400 ;
        RECT 151.600 30.200 152.400 30.400 ;
        RECT 166.000 30.300 166.800 39.800 ;
        RECT 170.200 32.400 171.000 39.800 ;
        RECT 171.600 33.600 172.400 34.400 ;
        RECT 171.800 32.400 172.400 33.600 ;
        RECT 170.200 31.800 171.200 32.400 ;
        RECT 171.800 31.800 173.200 32.400 ;
        RECT 169.200 30.300 170.000 30.400 ;
        RECT 151.600 29.600 156.600 30.200 ;
        RECT 145.200 29.000 146.000 29.200 ;
        RECT 147.000 28.400 147.600 29.600 ;
        RECT 153.200 29.400 154.000 29.600 ;
        RECT 155.800 29.400 156.600 29.600 ;
        RECT 166.000 29.700 170.000 30.300 ;
        RECT 154.200 28.400 155.000 28.600 ;
        RECT 147.000 28.300 158.000 28.400 ;
        RECT 161.200 28.300 162.000 28.400 ;
        RECT 147.000 27.800 162.000 28.300 ;
        RECT 147.400 27.600 148.200 27.800 ;
        RECT 140.400 26.600 144.200 27.200 ;
        RECT 135.800 26.200 139.400 26.600 ;
        RECT 114.800 26.000 118.800 26.200 ;
        RECT 114.800 22.200 115.600 26.000 ;
        RECT 118.000 22.200 118.800 26.000 ;
        RECT 119.600 22.200 120.400 26.200 ;
        RECT 121.200 22.200 122.000 26.200 ;
        RECT 122.800 26.000 126.800 26.200 ;
        RECT 122.800 22.200 123.600 26.000 ;
        RECT 126.000 22.200 126.800 26.000 ;
        RECT 127.600 26.000 131.600 26.200 ;
        RECT 127.600 22.200 128.400 26.000 ;
        RECT 130.800 22.200 131.600 26.000 ;
        RECT 132.400 22.200 133.200 26.200 ;
        RECT 134.000 22.200 134.800 26.200 ;
        RECT 135.600 26.000 139.600 26.200 ;
        RECT 135.600 22.200 136.400 26.000 ;
        RECT 138.800 22.200 139.600 26.000 ;
        RECT 140.400 22.200 141.200 26.600 ;
        RECT 143.400 26.400 144.200 26.600 ;
        RECT 153.200 25.600 153.800 27.800 ;
        RECT 156.400 27.700 162.000 27.800 ;
        RECT 156.400 27.600 158.000 27.700 ;
        RECT 161.200 27.600 162.000 27.700 ;
        RECT 151.400 25.400 152.200 25.600 ;
        RECT 145.200 24.200 146.000 25.000 ;
        RECT 149.400 24.800 152.200 25.400 ;
        RECT 153.200 24.800 154.000 25.600 ;
        RECT 149.400 24.200 150.000 24.800 ;
        RECT 154.800 24.200 155.600 25.000 ;
        RECT 144.600 23.600 146.000 24.200 ;
        RECT 144.600 22.200 145.800 23.600 ;
        RECT 149.200 22.200 150.000 24.200 ;
        RECT 153.600 23.600 155.600 24.200 ;
        RECT 153.600 22.200 154.400 23.600 ;
        RECT 158.000 22.200 158.800 27.000 ;
        RECT 162.800 26.300 163.600 26.400 ;
        RECT 164.400 26.300 165.200 26.400 ;
        RECT 162.800 25.700 165.200 26.300 ;
        RECT 162.800 25.600 163.600 25.700 ;
        RECT 164.400 24.800 165.200 25.700 ;
        RECT 166.000 22.200 166.800 29.700 ;
        RECT 169.200 28.800 170.000 29.700 ;
        RECT 170.600 28.400 171.200 31.800 ;
        RECT 172.400 31.600 173.200 31.800 ;
        RECT 174.000 31.600 174.800 33.200 ;
        RECT 172.500 30.300 173.100 31.600 ;
        RECT 175.600 30.300 176.400 39.800 ;
        RECT 180.400 32.000 181.200 39.800 ;
        RECT 183.600 35.200 184.400 39.800 ;
        RECT 172.500 29.700 176.400 30.300 ;
        RECT 167.600 28.200 168.400 28.400 ;
        RECT 167.600 27.600 169.200 28.200 ;
        RECT 170.600 27.600 173.200 28.400 ;
        RECT 168.400 27.200 169.200 27.600 ;
        RECT 167.800 26.200 171.400 26.600 ;
        RECT 172.400 26.200 173.000 27.600 ;
        RECT 175.600 26.200 176.400 29.700 ;
        RECT 180.200 31.200 181.200 32.000 ;
        RECT 181.800 34.600 184.400 35.200 ;
        RECT 181.800 33.000 182.400 34.600 ;
        RECT 186.800 34.400 187.600 39.800 ;
        RECT 190.000 37.000 190.800 39.800 ;
        RECT 191.600 37.000 192.400 39.800 ;
        RECT 193.200 37.000 194.000 39.800 ;
        RECT 188.200 34.400 192.400 35.200 ;
        RECT 185.000 33.600 187.600 34.400 ;
        RECT 194.800 33.600 195.600 39.800 ;
        RECT 198.000 35.000 198.800 39.800 ;
        RECT 201.200 35.000 202.000 39.800 ;
        RECT 202.800 37.000 203.600 39.800 ;
        RECT 204.400 37.000 205.200 39.800 ;
        RECT 207.600 35.200 208.400 39.800 ;
        RECT 210.800 36.400 211.600 39.800 ;
        RECT 210.800 35.800 211.800 36.400 ;
        RECT 211.200 35.200 211.800 35.800 ;
        RECT 206.400 34.400 210.600 35.200 ;
        RECT 211.200 34.600 213.200 35.200 ;
        RECT 198.000 33.600 200.600 34.400 ;
        RECT 201.200 33.800 207.000 34.400 ;
        RECT 210.000 34.000 210.600 34.400 ;
        RECT 190.000 33.000 190.800 33.200 ;
        RECT 181.800 32.400 190.800 33.000 ;
        RECT 193.200 33.000 194.000 33.200 ;
        RECT 201.200 33.000 201.800 33.800 ;
        RECT 207.600 33.200 209.000 33.800 ;
        RECT 210.000 33.200 211.600 34.000 ;
        RECT 193.200 32.400 201.800 33.000 ;
        RECT 202.800 33.000 209.000 33.200 ;
        RECT 202.800 32.600 208.200 33.000 ;
        RECT 202.800 32.400 203.600 32.600 ;
        RECT 177.200 28.300 178.000 28.400 ;
        RECT 180.200 28.300 181.000 31.200 ;
        RECT 181.800 30.600 182.400 32.400 ;
        RECT 177.200 27.700 181.000 28.300 ;
        RECT 177.200 26.800 178.000 27.700 ;
        RECT 180.200 26.800 181.000 27.700 ;
        RECT 181.600 30.000 182.400 30.600 ;
        RECT 188.400 30.000 211.800 30.600 ;
        RECT 181.600 28.000 182.200 30.000 ;
        RECT 188.400 29.400 189.200 30.000 ;
        RECT 206.000 29.600 206.800 30.000 ;
        RECT 211.000 29.800 211.800 30.000 ;
        RECT 182.800 28.600 186.600 29.400 ;
        RECT 181.600 27.400 182.800 28.000 ;
        RECT 167.600 26.000 171.600 26.200 ;
        RECT 167.600 22.200 168.400 26.000 ;
        RECT 170.800 22.200 171.600 26.000 ;
        RECT 172.400 22.200 173.200 26.200 ;
        RECT 174.600 25.600 176.400 26.200 ;
        RECT 180.200 26.000 181.200 26.800 ;
        RECT 174.600 22.200 175.400 25.600 ;
        RECT 180.400 22.200 181.200 26.000 ;
        RECT 182.000 22.200 182.800 27.400 ;
        RECT 185.800 27.400 186.600 28.600 ;
        RECT 185.800 26.800 187.600 27.400 ;
        RECT 186.800 26.200 187.600 26.800 ;
        RECT 191.600 26.400 192.400 29.200 ;
        RECT 194.800 28.600 198.000 29.400 ;
        RECT 201.800 28.600 203.800 29.400 ;
        RECT 212.400 29.000 213.200 34.600 ;
        RECT 194.400 27.800 195.200 28.000 ;
        RECT 194.400 27.200 198.800 27.800 ;
        RECT 198.000 27.000 198.800 27.200 ;
        RECT 199.600 26.800 200.400 28.400 ;
        RECT 186.800 25.400 189.200 26.200 ;
        RECT 191.600 25.600 192.600 26.400 ;
        RECT 195.600 25.600 197.200 26.400 ;
        RECT 198.000 26.200 198.800 26.400 ;
        RECT 201.800 26.200 202.600 28.600 ;
        RECT 204.400 28.200 213.200 29.000 ;
        RECT 207.800 26.800 210.800 27.600 ;
        RECT 207.800 26.200 208.600 26.800 ;
        RECT 198.000 25.600 202.600 26.200 ;
        RECT 188.400 22.200 189.200 25.400 ;
        RECT 206.000 25.400 208.600 26.200 ;
        RECT 190.000 22.200 190.800 25.000 ;
        RECT 191.600 22.200 192.400 25.000 ;
        RECT 193.200 22.200 194.000 25.000 ;
        RECT 194.800 22.200 195.600 25.000 ;
        RECT 198.000 22.200 198.800 25.000 ;
        RECT 201.200 22.200 202.000 25.000 ;
        RECT 202.800 22.200 203.600 25.000 ;
        RECT 204.400 22.200 205.200 25.000 ;
        RECT 206.000 22.200 206.800 25.400 ;
        RECT 212.400 22.200 213.200 28.200 ;
        RECT 214.000 30.300 214.800 39.800 ;
        RECT 218.000 33.600 218.800 34.400 ;
        RECT 218.000 32.400 218.600 33.600 ;
        RECT 219.400 32.400 220.200 39.800 ;
        RECT 224.400 33.600 225.200 34.400 ;
        RECT 224.400 32.400 225.000 33.600 ;
        RECT 225.800 32.400 226.600 39.800 ;
        RECT 217.200 31.800 218.600 32.400 ;
        RECT 219.200 31.800 220.200 32.400 ;
        RECT 223.600 31.800 225.000 32.400 ;
        RECT 225.600 31.800 226.600 32.400 ;
        RECT 217.200 31.600 218.000 31.800 ;
        RECT 217.200 30.300 218.000 30.400 ;
        RECT 214.000 29.700 218.000 30.300 ;
        RECT 214.000 22.200 214.800 29.700 ;
        RECT 217.200 29.600 218.000 29.700 ;
        RECT 219.200 28.400 219.800 31.800 ;
        RECT 223.600 31.600 224.400 31.800 ;
        RECT 220.400 28.800 221.200 30.400 ;
        RECT 225.600 28.400 226.200 31.800 ;
        RECT 226.800 30.300 227.600 30.400 ;
        RECT 230.000 30.300 230.800 39.800 ;
        RECT 234.800 36.400 235.600 39.800 ;
        RECT 234.600 35.800 235.600 36.400 ;
        RECT 234.600 35.200 235.200 35.800 ;
        RECT 238.000 35.200 238.800 39.800 ;
        RECT 241.200 37.000 242.000 39.800 ;
        RECT 242.800 37.000 243.600 39.800 ;
        RECT 226.800 29.700 230.800 30.300 ;
        RECT 226.800 28.800 227.600 29.700 ;
        RECT 217.200 27.600 219.800 28.400 ;
        RECT 222.000 28.200 222.800 28.400 ;
        RECT 221.200 27.600 222.800 28.200 ;
        RECT 223.600 27.600 226.200 28.400 ;
        RECT 228.400 28.200 229.200 28.400 ;
        RECT 227.600 27.600 229.200 28.200 ;
        RECT 215.600 24.800 216.400 26.400 ;
        RECT 217.400 26.200 218.000 27.600 ;
        RECT 221.200 27.200 222.000 27.600 ;
        RECT 219.000 26.200 222.600 26.600 ;
        RECT 223.800 26.200 224.400 27.600 ;
        RECT 227.600 27.200 228.400 27.600 ;
        RECT 225.400 26.200 229.000 26.600 ;
        RECT 217.200 22.200 218.000 26.200 ;
        RECT 218.800 26.000 222.800 26.200 ;
        RECT 218.800 22.200 219.600 26.000 ;
        RECT 222.000 22.200 222.800 26.000 ;
        RECT 223.600 22.200 224.400 26.200 ;
        RECT 225.200 26.000 229.200 26.200 ;
        RECT 225.200 22.200 226.000 26.000 ;
        RECT 228.400 22.200 229.200 26.000 ;
        RECT 230.000 22.200 230.800 29.700 ;
        RECT 233.200 34.600 235.200 35.200 ;
        RECT 233.200 29.000 234.000 34.600 ;
        RECT 235.800 34.400 240.000 35.200 ;
        RECT 244.400 35.000 245.200 39.800 ;
        RECT 247.600 35.000 248.400 39.800 ;
        RECT 235.800 34.000 236.400 34.400 ;
        RECT 234.800 33.200 236.400 34.000 ;
        RECT 239.400 33.800 245.200 34.400 ;
        RECT 237.400 33.200 238.800 33.800 ;
        RECT 237.400 33.000 243.600 33.200 ;
        RECT 238.200 32.600 243.600 33.000 ;
        RECT 242.800 32.400 243.600 32.600 ;
        RECT 244.600 33.000 245.200 33.800 ;
        RECT 245.800 33.600 248.400 34.400 ;
        RECT 250.800 33.600 251.600 39.800 ;
        RECT 252.400 37.000 253.200 39.800 ;
        RECT 254.000 37.000 254.800 39.800 ;
        RECT 255.600 37.000 256.400 39.800 ;
        RECT 254.000 34.400 258.200 35.200 ;
        RECT 258.800 34.400 259.600 39.800 ;
        RECT 262.000 35.200 262.800 39.800 ;
        RECT 262.000 34.600 264.600 35.200 ;
        RECT 258.800 33.600 261.400 34.400 ;
        RECT 252.400 33.000 253.200 33.200 ;
        RECT 244.600 32.400 253.200 33.000 ;
        RECT 255.600 33.000 256.400 33.200 ;
        RECT 264.000 33.000 264.600 34.600 ;
        RECT 255.600 32.400 264.600 33.000 ;
        RECT 264.000 30.600 264.600 32.400 ;
        RECT 265.200 32.000 266.000 39.800 ;
        RECT 265.200 31.200 266.200 32.000 ;
        RECT 234.600 30.000 258.000 30.600 ;
        RECT 264.000 30.000 264.800 30.600 ;
        RECT 234.600 29.800 235.400 30.000 ;
        RECT 239.600 29.600 240.400 30.000 ;
        RECT 257.200 29.400 258.000 30.000 ;
        RECT 233.200 28.200 242.000 29.000 ;
        RECT 242.600 28.600 244.600 29.400 ;
        RECT 248.400 28.600 251.600 29.400 ;
        RECT 231.600 24.800 232.400 26.400 ;
        RECT 233.200 22.200 234.000 28.200 ;
        RECT 235.600 26.800 238.600 27.600 ;
        RECT 237.800 26.200 238.600 26.800 ;
        RECT 243.800 26.200 244.600 28.600 ;
        RECT 246.000 26.800 246.800 28.400 ;
        RECT 251.200 27.800 252.000 28.000 ;
        RECT 247.600 27.200 252.000 27.800 ;
        RECT 247.600 27.000 248.400 27.200 ;
        RECT 254.000 26.400 254.800 29.200 ;
        RECT 259.800 28.600 263.600 29.400 ;
        RECT 259.800 27.400 260.600 28.600 ;
        RECT 264.200 28.000 264.800 30.000 ;
        RECT 247.600 26.200 248.400 26.400 ;
        RECT 237.800 25.400 240.400 26.200 ;
        RECT 243.800 25.600 248.400 26.200 ;
        RECT 249.200 25.600 250.800 26.400 ;
        RECT 253.800 25.600 254.800 26.400 ;
        RECT 258.800 26.800 260.600 27.400 ;
        RECT 263.600 27.400 264.800 28.000 ;
        RECT 258.800 26.200 259.600 26.800 ;
        RECT 239.600 22.200 240.400 25.400 ;
        RECT 257.200 25.400 259.600 26.200 ;
        RECT 241.200 22.200 242.000 25.000 ;
        RECT 242.800 22.200 243.600 25.000 ;
        RECT 244.400 22.200 245.200 25.000 ;
        RECT 247.600 22.200 248.400 25.000 ;
        RECT 250.800 22.200 251.600 25.000 ;
        RECT 252.400 22.200 253.200 25.000 ;
        RECT 254.000 22.200 254.800 25.000 ;
        RECT 255.600 22.200 256.400 25.000 ;
        RECT 257.200 22.200 258.000 25.400 ;
        RECT 263.600 22.200 264.400 27.400 ;
        RECT 265.400 26.800 266.200 31.200 ;
        RECT 265.200 26.300 266.200 26.800 ;
        RECT 268.400 26.300 269.200 26.400 ;
        RECT 265.200 25.700 269.200 26.300 ;
        RECT 265.200 22.200 266.000 25.700 ;
        RECT 268.400 24.800 269.200 25.700 ;
        RECT 270.000 22.200 270.800 39.800 ;
        RECT 273.200 36.400 274.000 39.800 ;
        RECT 273.000 35.800 274.000 36.400 ;
        RECT 273.000 35.200 273.600 35.800 ;
        RECT 276.400 35.200 277.200 39.800 ;
        RECT 279.600 37.000 280.400 39.800 ;
        RECT 281.200 37.000 282.000 39.800 ;
        RECT 271.600 34.600 273.600 35.200 ;
        RECT 271.600 29.000 272.400 34.600 ;
        RECT 274.200 34.400 278.400 35.200 ;
        RECT 282.800 35.000 283.600 39.800 ;
        RECT 286.000 35.000 286.800 39.800 ;
        RECT 274.200 34.000 274.800 34.400 ;
        RECT 273.200 33.200 274.800 34.000 ;
        RECT 277.800 33.800 283.600 34.400 ;
        RECT 275.800 33.200 277.200 33.800 ;
        RECT 275.800 33.000 282.000 33.200 ;
        RECT 276.600 32.600 282.000 33.000 ;
        RECT 281.200 32.400 282.000 32.600 ;
        RECT 283.000 33.000 283.600 33.800 ;
        RECT 284.200 33.600 286.800 34.400 ;
        RECT 289.200 33.600 290.000 39.800 ;
        RECT 290.800 37.000 291.600 39.800 ;
        RECT 292.400 37.000 293.200 39.800 ;
        RECT 294.000 37.000 294.800 39.800 ;
        RECT 292.400 34.400 296.600 35.200 ;
        RECT 297.200 34.400 298.000 39.800 ;
        RECT 300.400 35.200 301.200 39.800 ;
        RECT 300.400 34.600 303.000 35.200 ;
        RECT 297.200 33.600 299.800 34.400 ;
        RECT 290.800 33.000 291.600 33.200 ;
        RECT 283.000 32.400 291.600 33.000 ;
        RECT 294.000 33.000 294.800 33.200 ;
        RECT 302.400 33.000 303.000 34.600 ;
        RECT 294.000 32.400 303.000 33.000 ;
        RECT 302.400 30.600 303.000 32.400 ;
        RECT 303.600 32.000 304.400 39.800 ;
        RECT 303.600 31.200 304.600 32.000 ;
        RECT 273.000 30.000 296.400 30.600 ;
        RECT 302.400 30.000 303.200 30.600 ;
        RECT 273.000 29.800 273.800 30.000 ;
        RECT 278.000 29.600 278.800 30.000 ;
        RECT 295.600 29.400 296.400 30.000 ;
        RECT 271.600 28.200 280.400 29.000 ;
        RECT 281.000 28.600 283.000 29.400 ;
        RECT 286.800 28.600 290.000 29.400 ;
        RECT 271.600 22.200 272.400 28.200 ;
        RECT 274.000 26.800 277.000 27.600 ;
        RECT 276.200 26.200 277.000 26.800 ;
        RECT 282.200 26.200 283.000 28.600 ;
        RECT 284.400 26.800 285.200 28.400 ;
        RECT 289.600 27.800 290.400 28.000 ;
        RECT 286.000 27.200 290.400 27.800 ;
        RECT 286.000 27.000 286.800 27.200 ;
        RECT 292.400 26.400 293.200 29.200 ;
        RECT 298.200 28.600 302.000 29.400 ;
        RECT 298.200 27.400 299.000 28.600 ;
        RECT 302.600 28.000 303.200 30.000 ;
        RECT 286.000 26.200 286.800 26.400 ;
        RECT 276.200 25.400 278.800 26.200 ;
        RECT 282.200 25.600 286.800 26.200 ;
        RECT 287.600 25.600 289.200 26.400 ;
        RECT 292.200 25.600 293.200 26.400 ;
        RECT 297.200 26.800 299.000 27.400 ;
        RECT 302.000 27.400 303.200 28.000 ;
        RECT 297.200 26.200 298.000 26.800 ;
        RECT 278.000 22.200 278.800 25.400 ;
        RECT 295.600 25.400 298.000 26.200 ;
        RECT 279.600 22.200 280.400 25.000 ;
        RECT 281.200 22.200 282.000 25.000 ;
        RECT 282.800 22.200 283.600 25.000 ;
        RECT 286.000 22.200 286.800 25.000 ;
        RECT 289.200 22.200 290.000 25.000 ;
        RECT 290.800 22.200 291.600 25.000 ;
        RECT 292.400 22.200 293.200 25.000 ;
        RECT 294.000 22.200 294.800 25.000 ;
        RECT 295.600 22.200 296.400 25.400 ;
        RECT 302.000 22.200 302.800 27.400 ;
        RECT 303.800 26.800 304.600 31.200 ;
        RECT 303.600 26.000 304.600 26.800 ;
        RECT 310.000 26.300 310.800 26.400 ;
        RECT 311.600 26.300 312.400 26.400 ;
        RECT 303.600 22.200 304.400 26.000 ;
        RECT 310.000 25.700 312.400 26.300 ;
        RECT 310.000 25.600 310.800 25.700 ;
        RECT 311.600 24.800 312.400 25.700 ;
        RECT 313.200 22.200 314.000 39.800 ;
        RECT 314.800 32.400 315.600 39.800 ;
        RECT 316.400 32.400 317.200 32.600 ;
        RECT 319.200 32.400 320.800 39.800 ;
        RECT 314.800 31.800 317.200 32.400 ;
        RECT 318.800 31.800 320.800 32.400 ;
        RECT 323.000 32.400 323.800 32.600 ;
        RECT 324.400 32.400 325.200 39.800 ;
        RECT 323.000 31.800 325.200 32.400 ;
        RECT 326.000 35.000 326.800 39.000 ;
        RECT 330.200 38.400 331.000 39.800 ;
        RECT 330.200 37.600 331.600 38.400 ;
        RECT 318.800 30.400 319.400 31.800 ;
        RECT 323.000 31.200 323.600 31.800 ;
        RECT 320.200 30.600 323.600 31.200 ;
        RECT 326.000 31.600 326.600 35.000 ;
        RECT 330.200 32.800 331.000 37.600 ;
        RECT 330.200 32.200 331.800 32.800 ;
        RECT 326.000 31.000 329.800 31.600 ;
        RECT 320.200 30.400 321.000 30.600 ;
        RECT 314.800 30.300 315.600 30.400 ;
        RECT 318.000 30.300 319.400 30.400 ;
        RECT 326.000 30.300 326.800 30.400 ;
        RECT 314.800 29.800 319.400 30.300 ;
        RECT 322.400 29.800 323.200 30.000 ;
        RECT 314.800 29.700 319.800 29.800 ;
        RECT 314.800 29.600 315.600 29.700 ;
        RECT 318.000 29.600 319.800 29.700 ;
        RECT 318.800 29.200 319.800 29.600 ;
        RECT 314.800 27.600 316.400 28.400 ;
        RECT 317.600 27.600 318.400 28.400 ;
        RECT 317.800 27.200 318.400 27.600 ;
        RECT 316.400 26.800 317.200 27.000 ;
        RECT 314.800 26.200 317.200 26.800 ;
        RECT 317.800 26.400 318.600 27.200 ;
        RECT 314.800 22.200 315.600 26.200 ;
        RECT 319.200 25.800 319.800 29.200 ;
        RECT 320.600 29.200 323.200 29.800 ;
        RECT 324.500 29.700 326.800 30.300 ;
        RECT 320.600 28.600 321.200 29.200 ;
        RECT 320.400 27.800 321.200 28.600 ;
        RECT 324.500 28.400 325.100 29.700 ;
        RECT 326.000 28.800 326.800 29.700 ;
        RECT 327.600 28.800 328.400 30.400 ;
        RECT 329.200 29.000 329.800 31.000 ;
        RECT 323.600 28.200 325.200 28.400 ;
        RECT 321.800 27.600 325.200 28.200 ;
        RECT 329.200 28.200 330.600 29.000 ;
        RECT 331.200 28.400 331.800 32.200 ;
        RECT 335.600 32.400 336.400 39.800 ;
        RECT 340.000 38.400 341.600 39.800 ;
        RECT 338.800 37.600 341.600 38.400 ;
        RECT 337.400 32.400 338.200 32.600 ;
        RECT 335.600 31.800 338.200 32.400 ;
        RECT 340.000 31.800 341.600 37.600 ;
        RECT 343.600 32.400 344.400 32.600 ;
        RECT 345.200 32.400 346.000 39.800 ;
        RECT 348.400 35.800 349.200 39.800 ;
        RECT 348.600 35.600 349.200 35.800 ;
        RECT 351.600 35.800 352.400 39.800 ;
        RECT 355.800 38.400 356.600 39.800 ;
        RECT 355.800 37.600 357.200 38.400 ;
        RECT 351.600 35.600 352.200 35.800 ;
        RECT 348.600 35.000 352.200 35.600 ;
        RECT 350.000 32.800 350.800 34.400 ;
        RECT 351.600 32.400 352.200 35.000 ;
        RECT 355.800 32.600 356.600 37.600 ;
        RECT 343.600 31.800 346.000 32.400 ;
        RECT 332.400 30.300 333.200 31.200 ;
        RECT 338.600 30.400 339.400 30.600 ;
        RECT 340.600 30.400 341.200 31.800 ;
        RECT 346.800 30.800 347.600 32.400 ;
        RECT 351.600 31.600 352.400 32.400 ;
        RECT 354.800 31.800 356.600 32.600 ;
        RECT 359.600 32.000 360.400 39.800 ;
        RECT 362.800 35.200 363.600 39.800 ;
        RECT 332.400 29.700 336.300 30.300 ;
        RECT 332.400 29.600 333.200 29.700 ;
        RECT 335.700 28.400 336.300 29.700 ;
        RECT 337.800 29.800 339.400 30.400 ;
        RECT 337.800 29.600 338.600 29.800 ;
        RECT 340.400 29.600 341.200 30.400 ;
        RECT 348.400 29.600 350.000 30.400 ;
        RECT 339.200 28.600 340.000 28.800 ;
        RECT 337.200 28.400 340.000 28.600 ;
        RECT 329.200 27.800 330.200 28.200 ;
        RECT 321.800 27.200 322.400 27.600 ;
        RECT 320.400 26.600 322.400 27.200 ;
        RECT 326.000 27.200 330.200 27.800 ;
        RECT 331.200 27.600 333.200 28.400 ;
        RECT 335.600 28.000 340.000 28.400 ;
        RECT 340.600 28.400 341.200 29.600 ;
        RECT 351.600 28.400 352.200 31.600 ;
        RECT 355.000 28.400 355.600 31.800 ;
        RECT 359.400 31.200 360.400 32.000 ;
        RECT 361.000 34.600 363.600 35.200 ;
        RECT 361.000 33.000 361.600 34.600 ;
        RECT 366.000 34.400 366.800 39.800 ;
        RECT 369.200 37.000 370.000 39.800 ;
        RECT 370.800 37.000 371.600 39.800 ;
        RECT 372.400 37.000 373.200 39.800 ;
        RECT 367.400 34.400 371.600 35.200 ;
        RECT 364.200 33.600 366.800 34.400 ;
        RECT 374.000 33.600 374.800 39.800 ;
        RECT 377.200 35.000 378.000 39.800 ;
        RECT 380.400 35.000 381.200 39.800 ;
        RECT 382.000 37.000 382.800 39.800 ;
        RECT 383.600 37.000 384.400 39.800 ;
        RECT 386.800 35.200 387.600 39.800 ;
        RECT 390.000 36.400 390.800 39.800 ;
        RECT 390.000 35.800 391.000 36.400 ;
        RECT 390.400 35.200 391.000 35.800 ;
        RECT 385.600 34.400 389.800 35.200 ;
        RECT 390.400 34.600 392.400 35.200 ;
        RECT 377.200 33.600 379.800 34.400 ;
        RECT 380.400 33.800 386.200 34.400 ;
        RECT 389.200 34.000 389.800 34.400 ;
        RECT 369.200 33.000 370.000 33.200 ;
        RECT 361.000 32.400 370.000 33.000 ;
        RECT 372.400 33.000 373.200 33.200 ;
        RECT 380.400 33.000 381.000 33.800 ;
        RECT 386.800 33.200 388.200 33.800 ;
        RECT 389.200 33.200 390.800 34.000 ;
        RECT 372.400 32.400 381.000 33.000 ;
        RECT 382.000 33.000 388.200 33.200 ;
        RECT 382.000 32.600 387.400 33.000 ;
        RECT 382.000 32.400 382.800 32.600 ;
        RECT 356.400 29.600 357.200 31.200 ;
        RECT 335.600 27.800 337.800 28.000 ;
        RECT 340.600 27.800 341.600 28.400 ;
        RECT 335.600 27.600 337.200 27.800 ;
        RECT 323.000 26.800 323.800 27.000 ;
        RECT 320.400 26.400 322.000 26.600 ;
        RECT 323.000 26.200 325.200 26.800 ;
        RECT 319.200 22.200 320.800 25.800 ;
        RECT 324.400 22.200 325.200 26.200 ;
        RECT 326.000 25.000 326.600 27.200 ;
        RECT 331.200 27.000 331.800 27.600 ;
        RECT 331.000 26.600 331.800 27.000 ;
        RECT 337.400 26.800 338.200 27.000 ;
        RECT 330.200 26.000 331.800 26.600 ;
        RECT 335.600 26.200 338.200 26.800 ;
        RECT 338.800 26.400 340.400 27.200 ;
        RECT 326.000 23.000 326.800 25.000 ;
        RECT 330.200 23.000 331.000 26.000 ;
        RECT 335.600 22.200 336.400 26.200 ;
        RECT 341.000 25.800 341.600 27.800 ;
        RECT 342.400 27.600 343.200 28.400 ;
        RECT 344.400 27.600 346.000 28.400 ;
        RECT 350.600 28.200 352.200 28.400 ;
        RECT 350.400 27.800 352.200 28.200 ;
        RECT 342.400 27.200 343.000 27.600 ;
        RECT 342.200 26.400 343.000 27.200 ;
        RECT 343.600 26.800 344.400 27.000 ;
        RECT 343.600 26.200 346.000 26.800 ;
        RECT 340.000 22.200 341.600 25.800 ;
        RECT 345.200 22.200 346.000 26.200 ;
        RECT 350.400 22.200 351.200 27.800 ;
        RECT 354.800 27.600 355.600 28.400 ;
        RECT 353.200 24.800 354.000 26.400 ;
        RECT 355.000 24.200 355.600 27.600 ;
        RECT 359.400 26.800 360.200 31.200 ;
        RECT 361.000 30.600 361.600 32.400 ;
        RECT 360.800 30.000 361.600 30.600 ;
        RECT 367.600 30.000 391.000 30.600 ;
        RECT 360.800 28.000 361.400 30.000 ;
        RECT 367.600 29.400 368.400 30.000 ;
        RECT 385.200 29.600 386.000 30.000 ;
        RECT 390.200 29.800 391.000 30.000 ;
        RECT 362.000 28.600 365.800 29.400 ;
        RECT 360.800 27.400 362.000 28.000 ;
        RECT 359.400 26.000 360.400 26.800 ;
        RECT 354.800 22.200 355.600 24.200 ;
        RECT 359.600 22.200 360.400 26.000 ;
        RECT 361.200 22.200 362.000 27.400 ;
        RECT 365.000 27.400 365.800 28.600 ;
        RECT 365.000 26.800 366.800 27.400 ;
        RECT 366.000 26.200 366.800 26.800 ;
        RECT 370.800 26.400 371.600 29.200 ;
        RECT 374.000 28.600 377.200 29.400 ;
        RECT 381.000 28.600 383.000 29.400 ;
        RECT 391.600 29.000 392.400 34.600 ;
        RECT 394.800 31.200 395.600 39.800 ;
        RECT 398.000 31.200 398.800 39.800 ;
        RECT 401.200 31.200 402.000 39.800 ;
        RECT 404.400 31.200 405.200 39.800 ;
        RECT 373.600 27.800 374.400 28.000 ;
        RECT 373.600 27.200 378.000 27.800 ;
        RECT 377.200 27.000 378.000 27.200 ;
        RECT 378.800 26.800 379.600 28.400 ;
        RECT 366.000 25.400 368.400 26.200 ;
        RECT 370.800 25.600 371.800 26.400 ;
        RECT 374.800 25.600 376.400 26.400 ;
        RECT 377.200 26.200 378.000 26.400 ;
        RECT 381.000 26.200 381.800 28.600 ;
        RECT 383.600 28.200 392.400 29.000 ;
        RECT 387.000 26.800 390.000 27.600 ;
        RECT 387.000 26.200 387.800 26.800 ;
        RECT 377.200 25.600 381.800 26.200 ;
        RECT 367.600 22.200 368.400 25.400 ;
        RECT 385.200 25.400 387.800 26.200 ;
        RECT 369.200 22.200 370.000 25.000 ;
        RECT 370.800 22.200 371.600 25.000 ;
        RECT 372.400 22.200 373.200 25.000 ;
        RECT 374.000 22.200 374.800 25.000 ;
        RECT 377.200 22.200 378.000 25.000 ;
        RECT 380.400 22.200 381.200 25.000 ;
        RECT 382.000 22.200 382.800 25.000 ;
        RECT 383.600 22.200 384.400 25.000 ;
        RECT 385.200 22.200 386.000 25.400 ;
        RECT 391.600 22.200 392.400 28.200 ;
        RECT 393.200 30.400 395.600 31.200 ;
        RECT 396.600 30.400 398.800 31.200 ;
        RECT 399.800 30.400 402.000 31.200 ;
        RECT 403.400 30.400 405.200 31.200 ;
        RECT 409.200 31.200 410.000 39.800 ;
        RECT 412.400 31.200 413.200 39.800 ;
        RECT 415.600 31.200 416.400 39.800 ;
        RECT 418.800 31.200 419.600 39.800 ;
        RECT 424.600 32.400 425.400 39.800 ;
        RECT 428.400 35.800 429.200 39.800 ;
        RECT 428.600 35.600 429.200 35.800 ;
        RECT 431.600 35.800 432.400 39.800 ;
        RECT 431.600 35.600 432.200 35.800 ;
        RECT 428.600 35.000 432.200 35.600 ;
        RECT 426.000 33.600 426.800 34.400 ;
        RECT 426.200 32.400 426.800 33.600 ;
        RECT 428.600 32.400 429.200 35.000 ;
        RECT 430.000 32.800 430.800 34.400 ;
        RECT 435.600 33.600 436.400 34.400 ;
        RECT 435.600 32.400 436.200 33.600 ;
        RECT 437.000 32.400 437.800 39.800 ;
        RECT 441.200 35.800 442.000 39.800 ;
        RECT 441.400 35.600 442.000 35.800 ;
        RECT 444.400 35.800 445.200 39.800 ;
        RECT 444.400 35.600 445.000 35.800 ;
        RECT 441.400 35.000 445.000 35.600 ;
        RECT 441.400 32.400 442.000 35.000 ;
        RECT 442.800 32.800 443.600 34.400 ;
        RECT 448.400 33.600 449.200 34.400 ;
        RECT 448.400 32.400 449.000 33.600 ;
        RECT 449.800 32.400 450.600 39.800 ;
        RECT 424.600 31.800 425.600 32.400 ;
        RECT 426.200 31.800 427.600 32.400 ;
        RECT 409.200 30.400 411.000 31.200 ;
        RECT 412.400 30.400 414.600 31.200 ;
        RECT 415.600 30.400 417.800 31.200 ;
        RECT 418.800 30.400 421.200 31.200 ;
        RECT 393.200 27.600 394.000 30.400 ;
        RECT 396.600 29.000 397.400 30.400 ;
        RECT 399.800 29.000 400.600 30.400 ;
        RECT 403.400 29.000 404.200 30.400 ;
        RECT 410.200 29.000 411.000 30.400 ;
        RECT 413.800 29.000 414.600 30.400 ;
        RECT 417.000 29.000 417.800 30.400 ;
        RECT 394.800 28.200 397.400 29.000 ;
        RECT 398.200 28.200 400.600 29.000 ;
        RECT 401.600 28.200 404.200 29.000 ;
        RECT 405.000 28.300 406.800 29.000 ;
        RECT 407.600 28.300 409.400 29.000 ;
        RECT 405.000 28.200 409.400 28.300 ;
        RECT 410.200 28.200 412.800 29.000 ;
        RECT 413.800 28.200 416.200 29.000 ;
        RECT 417.000 28.200 419.600 29.000 ;
        RECT 396.600 27.600 397.400 28.200 ;
        RECT 399.800 27.600 400.600 28.200 ;
        RECT 403.400 27.600 404.200 28.200 ;
        RECT 406.000 27.700 408.400 28.200 ;
        RECT 406.000 27.600 406.800 27.700 ;
        RECT 407.600 27.600 408.400 27.700 ;
        RECT 410.200 27.600 411.000 28.200 ;
        RECT 413.800 27.600 414.600 28.200 ;
        RECT 417.000 27.600 417.800 28.200 ;
        RECT 420.400 27.600 421.200 30.400 ;
        RECT 423.600 28.800 424.400 30.400 ;
        RECT 425.000 28.400 425.600 31.800 ;
        RECT 426.800 31.600 427.600 31.800 ;
        RECT 428.400 31.600 429.200 32.400 ;
        RECT 428.600 28.400 429.200 31.600 ;
        RECT 433.200 32.300 434.000 32.400 ;
        RECT 434.800 32.300 436.200 32.400 ;
        RECT 433.200 31.800 436.200 32.300 ;
        RECT 436.800 31.800 437.800 32.400 ;
        RECT 433.200 31.700 435.600 31.800 ;
        RECT 433.200 30.800 434.000 31.700 ;
        RECT 434.800 31.600 435.600 31.700 ;
        RECT 436.800 30.400 437.400 31.800 ;
        RECT 441.200 31.600 442.000 32.400 ;
        RECT 430.800 29.600 432.400 30.400 ;
        RECT 436.400 29.600 437.400 30.400 ;
        RECT 436.800 28.400 437.400 29.600 ;
        RECT 438.000 28.800 438.800 30.400 ;
        RECT 441.400 28.400 442.000 31.600 ;
        RECT 446.000 32.300 446.800 32.400 ;
        RECT 447.600 32.300 449.000 32.400 ;
        RECT 446.000 31.800 449.000 32.300 ;
        RECT 449.600 31.800 450.600 32.400 ;
        RECT 446.000 31.700 448.400 31.800 ;
        RECT 446.000 30.800 446.800 31.700 ;
        RECT 447.600 31.600 448.400 31.700 ;
        RECT 443.600 29.600 445.200 30.400 ;
        RECT 449.600 28.400 450.200 31.800 ;
        RECT 458.800 31.400 459.600 39.800 ;
        RECT 463.200 36.400 464.000 39.800 ;
        RECT 462.000 35.800 464.000 36.400 ;
        RECT 467.600 35.800 468.400 39.800 ;
        RECT 471.800 35.800 473.000 39.800 ;
        RECT 462.000 35.000 462.800 35.800 ;
        RECT 467.600 35.200 468.200 35.800 ;
        RECT 465.400 34.600 469.000 35.200 ;
        RECT 471.600 35.000 472.400 35.800 ;
        RECT 465.400 34.400 466.200 34.600 ;
        RECT 468.200 34.400 469.000 34.600 ;
        RECT 462.000 33.000 462.800 33.200 ;
        RECT 466.600 33.000 467.400 33.200 ;
        RECT 462.000 32.400 467.400 33.000 ;
        RECT 468.000 33.000 470.200 33.600 ;
        RECT 468.000 31.800 468.600 33.000 ;
        RECT 469.400 32.800 470.200 33.000 ;
        RECT 471.800 33.200 473.200 34.000 ;
        RECT 471.800 32.200 472.400 33.200 ;
        RECT 463.800 31.400 468.600 31.800 ;
        RECT 458.800 31.200 468.600 31.400 ;
        RECT 470.000 31.600 472.400 32.200 ;
        RECT 458.800 31.000 464.600 31.200 ;
        RECT 458.800 30.800 464.400 31.000 ;
        RECT 470.000 30.400 470.600 31.600 ;
        RECT 476.400 31.200 477.200 39.800 ;
        RECT 480.600 32.400 481.400 39.800 ;
        RECT 482.000 33.600 482.800 34.400 ;
        RECT 482.200 32.400 482.800 33.600 ;
        RECT 485.200 33.600 486.000 34.400 ;
        RECT 485.200 32.400 485.800 33.600 ;
        RECT 486.600 32.400 487.400 39.800 ;
        RECT 480.600 31.800 481.600 32.400 ;
        RECT 482.200 31.800 483.600 32.400 ;
        RECT 473.000 30.600 477.200 31.200 ;
        RECT 473.000 30.400 473.800 30.600 ;
        RECT 450.800 28.800 451.600 30.400 ;
        RECT 465.200 30.200 466.000 30.400 ;
        RECT 461.000 29.600 466.000 30.200 ;
        RECT 470.000 29.600 470.800 30.400 ;
        RECT 474.600 29.800 475.400 30.000 ;
        RECT 461.000 29.400 461.800 29.600 ;
        RECT 462.600 28.400 463.400 28.600 ;
        RECT 470.000 28.400 470.600 29.600 ;
        RECT 471.600 29.200 475.400 29.800 ;
        RECT 471.600 29.000 472.400 29.200 ;
        RECT 422.000 28.200 422.800 28.400 ;
        RECT 422.000 27.600 423.600 28.200 ;
        RECT 425.000 27.600 427.600 28.400 ;
        RECT 428.600 28.200 430.200 28.400 ;
        RECT 428.600 27.800 430.400 28.200 ;
        RECT 393.200 26.800 395.600 27.600 ;
        RECT 396.600 26.800 398.800 27.600 ;
        RECT 399.800 26.800 402.000 27.600 ;
        RECT 403.400 26.800 405.200 27.600 ;
        RECT 394.800 22.200 395.600 26.800 ;
        RECT 398.000 22.200 398.800 26.800 ;
        RECT 401.200 22.200 402.000 26.800 ;
        RECT 404.400 22.200 405.200 26.800 ;
        RECT 409.200 26.800 411.000 27.600 ;
        RECT 412.400 26.800 414.600 27.600 ;
        RECT 415.600 26.800 417.800 27.600 ;
        RECT 418.800 26.800 421.200 27.600 ;
        RECT 422.800 27.200 423.600 27.600 ;
        RECT 409.200 22.200 410.000 26.800 ;
        RECT 412.400 22.200 413.200 26.800 ;
        RECT 415.600 22.200 416.400 26.800 ;
        RECT 418.800 22.200 419.600 26.800 ;
        RECT 422.200 26.200 425.800 26.600 ;
        RECT 426.800 26.200 427.400 27.600 ;
        RECT 422.000 26.000 426.000 26.200 ;
        RECT 422.000 22.200 422.800 26.000 ;
        RECT 425.200 22.200 426.000 26.000 ;
        RECT 426.800 22.200 427.600 26.200 ;
        RECT 429.600 22.200 430.400 27.800 ;
        RECT 434.800 27.600 437.400 28.400 ;
        RECT 439.600 28.200 440.400 28.400 ;
        RECT 438.800 27.600 440.400 28.200 ;
        RECT 441.400 28.200 443.000 28.400 ;
        RECT 441.400 27.800 443.200 28.200 ;
        RECT 435.000 26.200 435.600 27.600 ;
        RECT 438.800 27.200 439.600 27.600 ;
        RECT 436.600 26.200 440.200 26.600 ;
        RECT 434.800 22.200 435.600 26.200 ;
        RECT 436.400 26.000 440.400 26.200 ;
        RECT 436.400 22.200 437.200 26.000 ;
        RECT 439.600 22.200 440.400 26.000 ;
        RECT 442.400 22.200 443.200 27.800 ;
        RECT 447.600 27.600 450.200 28.400 ;
        RECT 452.400 28.200 453.200 28.400 ;
        RECT 451.600 27.600 453.200 28.200 ;
        RECT 459.600 27.800 470.600 28.400 ;
        RECT 459.600 27.600 461.200 27.800 ;
        RECT 447.800 26.200 448.400 27.600 ;
        RECT 451.600 27.200 452.400 27.600 ;
        RECT 449.400 26.200 453.000 26.600 ;
        RECT 447.600 22.200 448.400 26.200 ;
        RECT 449.200 26.000 453.200 26.200 ;
        RECT 449.200 22.200 450.000 26.000 ;
        RECT 452.400 22.200 453.200 26.000 ;
        RECT 458.800 22.200 459.600 27.000 ;
        RECT 463.800 25.600 464.400 27.800 ;
        RECT 469.400 27.600 470.200 27.800 ;
        RECT 476.400 27.200 477.200 30.600 ;
        RECT 481.000 30.400 481.600 31.800 ;
        RECT 482.800 31.600 483.600 31.800 ;
        RECT 484.400 31.800 485.800 32.400 ;
        RECT 486.400 31.800 487.400 32.400 ;
        RECT 484.400 31.600 485.200 31.800 ;
        RECT 478.000 30.300 478.800 30.400 ;
        RECT 479.600 30.300 480.400 30.400 ;
        RECT 478.000 29.700 480.400 30.300 ;
        RECT 478.000 29.600 478.800 29.700 ;
        RECT 479.600 28.800 480.400 29.700 ;
        RECT 481.000 29.600 482.000 30.400 ;
        RECT 482.900 30.300 483.500 31.600 ;
        RECT 486.400 30.300 487.000 31.800 ;
        RECT 490.800 31.400 491.600 39.800 ;
        RECT 495.200 36.400 496.000 39.800 ;
        RECT 494.000 35.800 496.000 36.400 ;
        RECT 499.600 35.800 500.400 39.800 ;
        RECT 503.800 35.800 505.000 39.800 ;
        RECT 494.000 35.000 494.800 35.800 ;
        RECT 499.600 35.200 500.200 35.800 ;
        RECT 497.400 34.600 501.000 35.200 ;
        RECT 503.600 35.000 504.400 35.800 ;
        RECT 497.400 34.400 498.200 34.600 ;
        RECT 500.200 34.400 501.000 34.600 ;
        RECT 494.000 33.000 494.800 33.200 ;
        RECT 498.600 33.000 499.400 33.200 ;
        RECT 494.000 32.400 499.400 33.000 ;
        RECT 500.000 33.000 502.200 33.600 ;
        RECT 500.000 31.800 500.600 33.000 ;
        RECT 501.400 32.800 502.200 33.000 ;
        RECT 503.800 33.200 505.200 34.000 ;
        RECT 503.800 32.200 504.400 33.200 ;
        RECT 495.800 31.400 500.600 31.800 ;
        RECT 490.800 31.200 500.600 31.400 ;
        RECT 502.000 31.600 504.400 32.200 ;
        RECT 490.800 31.000 496.600 31.200 ;
        RECT 490.800 30.800 496.400 31.000 ;
        RECT 502.000 30.400 502.600 31.600 ;
        RECT 508.400 31.200 509.200 39.800 ;
        RECT 512.600 32.400 513.400 39.800 ;
        RECT 514.000 33.600 514.800 34.400 ;
        RECT 514.200 32.400 514.800 33.600 ;
        RECT 517.200 33.600 518.000 34.400 ;
        RECT 517.200 32.400 517.800 33.600 ;
        RECT 518.600 32.400 519.400 39.800 ;
        RECT 512.600 31.800 513.600 32.400 ;
        RECT 514.200 31.800 515.600 32.400 ;
        RECT 505.000 30.600 509.200 31.200 ;
        RECT 505.000 30.400 505.800 30.600 ;
        RECT 482.900 29.700 487.000 30.300 ;
        RECT 481.000 28.400 481.600 29.600 ;
        RECT 486.400 28.400 487.000 29.700 ;
        RECT 487.600 30.300 488.400 30.400 ;
        RECT 489.200 30.300 490.000 30.400 ;
        RECT 487.600 29.700 490.000 30.300 ;
        RECT 497.200 30.200 498.000 30.400 ;
        RECT 487.600 28.800 488.400 29.700 ;
        RECT 489.200 29.600 490.000 29.700 ;
        RECT 493.000 29.600 498.000 30.200 ;
        RECT 502.000 29.600 502.800 30.400 ;
        RECT 506.600 29.800 507.400 30.000 ;
        RECT 493.000 29.400 493.800 29.600 ;
        RECT 494.600 28.400 495.400 28.600 ;
        RECT 502.000 28.400 502.600 29.600 ;
        RECT 503.600 29.200 507.400 29.800 ;
        RECT 503.600 29.000 504.400 29.200 ;
        RECT 478.000 28.200 478.800 28.400 ;
        RECT 478.000 27.600 479.600 28.200 ;
        RECT 481.000 27.600 483.600 28.400 ;
        RECT 484.400 27.600 487.000 28.400 ;
        RECT 489.200 28.200 490.000 28.400 ;
        RECT 488.400 27.600 490.000 28.200 ;
        RECT 491.600 27.800 502.600 28.400 ;
        RECT 491.600 27.600 493.200 27.800 ;
        RECT 478.800 27.200 479.600 27.600 ;
        RECT 473.400 26.600 477.200 27.200 ;
        RECT 473.400 26.400 474.200 26.600 ;
        RECT 462.000 24.200 462.800 25.000 ;
        RECT 463.600 24.800 464.400 25.600 ;
        RECT 465.400 25.400 466.200 25.600 ;
        RECT 465.400 24.800 468.200 25.400 ;
        RECT 467.600 24.200 468.200 24.800 ;
        RECT 471.600 24.200 472.400 25.000 ;
        RECT 462.000 23.600 464.000 24.200 ;
        RECT 463.200 22.200 464.000 23.600 ;
        RECT 467.600 22.200 468.400 24.200 ;
        RECT 471.600 23.600 473.000 24.200 ;
        RECT 471.800 22.200 473.000 23.600 ;
        RECT 476.400 22.200 477.200 26.600 ;
        RECT 478.200 26.200 481.800 26.600 ;
        RECT 482.800 26.200 483.400 27.600 ;
        RECT 484.600 26.200 485.200 27.600 ;
        RECT 488.400 27.200 489.200 27.600 ;
        RECT 486.200 26.200 489.800 26.600 ;
        RECT 478.000 26.000 482.000 26.200 ;
        RECT 478.000 22.200 478.800 26.000 ;
        RECT 481.200 22.200 482.000 26.000 ;
        RECT 482.800 22.200 483.600 26.200 ;
        RECT 484.400 22.200 485.200 26.200 ;
        RECT 486.000 26.000 490.000 26.200 ;
        RECT 486.000 22.200 486.800 26.000 ;
        RECT 489.200 22.200 490.000 26.000 ;
        RECT 490.800 22.200 491.600 27.000 ;
        RECT 495.800 25.600 496.400 27.800 ;
        RECT 501.400 27.600 502.200 27.800 ;
        RECT 508.400 27.200 509.200 30.600 ;
        RECT 513.000 30.400 513.600 31.800 ;
        RECT 514.800 31.600 515.600 31.800 ;
        RECT 516.400 31.800 517.800 32.400 ;
        RECT 518.400 31.800 519.400 32.400 ;
        RECT 516.400 31.600 517.200 31.800 ;
        RECT 510.000 30.300 510.800 30.400 ;
        RECT 511.600 30.300 512.400 30.400 ;
        RECT 510.000 29.700 512.400 30.300 ;
        RECT 510.000 29.600 510.800 29.700 ;
        RECT 511.600 28.800 512.400 29.700 ;
        RECT 513.000 29.600 514.000 30.400 ;
        RECT 514.900 30.300 515.500 31.600 ;
        RECT 518.400 30.300 519.000 31.800 ;
        RECT 524.400 31.200 525.200 39.800 ;
        RECT 527.600 31.200 528.400 39.800 ;
        RECT 530.800 31.200 531.600 39.800 ;
        RECT 534.000 31.200 534.800 39.800 ;
        RECT 522.800 30.400 525.200 31.200 ;
        RECT 526.200 30.400 528.400 31.200 ;
        RECT 529.400 30.400 531.600 31.200 ;
        RECT 533.000 30.400 534.800 31.200 ;
        RECT 514.900 29.700 519.000 30.300 ;
        RECT 513.000 28.400 513.600 29.600 ;
        RECT 518.400 28.400 519.000 29.700 ;
        RECT 519.600 28.800 520.400 30.400 ;
        RECT 510.000 28.200 510.800 28.400 ;
        RECT 510.000 27.600 511.600 28.200 ;
        RECT 513.000 27.600 515.600 28.400 ;
        RECT 516.400 27.600 519.000 28.400 ;
        RECT 521.200 28.200 522.000 28.400 ;
        RECT 520.400 27.600 522.000 28.200 ;
        RECT 522.800 27.600 523.600 30.400 ;
        RECT 526.200 29.000 527.000 30.400 ;
        RECT 529.400 29.000 530.200 30.400 ;
        RECT 533.000 29.000 533.800 30.400 ;
        RECT 524.400 28.200 527.000 29.000 ;
        RECT 527.800 28.200 530.200 29.000 ;
        RECT 531.200 28.200 533.800 29.000 ;
        RECT 534.600 28.200 536.400 29.000 ;
        RECT 526.200 27.600 527.000 28.200 ;
        RECT 529.400 27.600 530.200 28.200 ;
        RECT 533.000 27.600 533.800 28.200 ;
        RECT 535.600 27.600 536.400 28.200 ;
        RECT 510.800 27.200 511.600 27.600 ;
        RECT 505.400 26.600 509.200 27.200 ;
        RECT 505.400 26.400 506.200 26.600 ;
        RECT 494.000 24.200 494.800 25.000 ;
        RECT 495.600 24.800 496.400 25.600 ;
        RECT 497.400 25.400 498.200 25.600 ;
        RECT 497.400 24.800 500.200 25.400 ;
        RECT 499.600 24.200 500.200 24.800 ;
        RECT 503.600 24.200 504.400 25.000 ;
        RECT 494.000 23.600 496.000 24.200 ;
        RECT 495.200 22.200 496.000 23.600 ;
        RECT 499.600 22.200 500.400 24.200 ;
        RECT 503.600 23.600 505.000 24.200 ;
        RECT 503.800 22.200 505.000 23.600 ;
        RECT 508.400 22.200 509.200 26.600 ;
        RECT 510.200 26.200 513.800 26.600 ;
        RECT 514.800 26.200 515.400 27.600 ;
        RECT 516.600 26.200 517.200 27.600 ;
        RECT 520.400 27.200 521.200 27.600 ;
        RECT 522.800 26.800 525.200 27.600 ;
        RECT 526.200 26.800 528.400 27.600 ;
        RECT 529.400 26.800 531.600 27.600 ;
        RECT 533.000 26.800 534.800 27.600 ;
        RECT 518.200 26.200 521.800 26.600 ;
        RECT 510.000 26.000 514.000 26.200 ;
        RECT 510.000 22.200 510.800 26.000 ;
        RECT 513.200 22.200 514.000 26.000 ;
        RECT 514.800 22.200 515.600 26.200 ;
        RECT 516.400 22.200 517.200 26.200 ;
        RECT 518.000 26.000 522.000 26.200 ;
        RECT 518.000 22.200 518.800 26.000 ;
        RECT 521.200 22.200 522.000 26.000 ;
        RECT 524.400 22.200 525.200 26.800 ;
        RECT 527.600 22.200 528.400 26.800 ;
        RECT 530.800 22.200 531.600 26.800 ;
        RECT 534.000 22.200 534.800 26.800 ;
        RECT 537.200 22.200 538.000 39.800 ;
        RECT 542.600 34.400 543.400 39.800 ;
        RECT 541.200 33.600 542.000 34.400 ;
        RECT 542.600 33.600 544.400 34.400 ;
        RECT 541.200 32.400 541.800 33.600 ;
        RECT 542.600 32.400 543.400 33.600 ;
        RECT 538.800 32.300 539.600 32.400 ;
        RECT 540.400 32.300 541.800 32.400 ;
        RECT 538.800 31.800 541.800 32.300 ;
        RECT 542.400 31.800 543.400 32.400 ;
        RECT 549.400 32.400 550.200 39.800 ;
        RECT 550.800 33.600 551.600 34.400 ;
        RECT 551.000 32.400 551.600 33.600 ;
        RECT 554.000 33.600 554.800 34.400 ;
        RECT 554.000 32.400 554.600 33.600 ;
        RECT 555.400 32.400 556.200 39.800 ;
        RECT 560.400 33.600 561.200 34.400 ;
        RECT 560.400 32.400 561.000 33.600 ;
        RECT 561.800 32.400 562.600 39.800 ;
        RECT 549.400 31.800 550.400 32.400 ;
        RECT 551.000 31.800 552.400 32.400 ;
        RECT 538.800 31.700 541.200 31.800 ;
        RECT 538.800 31.600 539.600 31.700 ;
        RECT 540.400 31.600 541.200 31.700 ;
        RECT 542.400 28.400 543.000 31.800 ;
        RECT 543.600 30.300 544.400 30.400 ;
        RECT 548.400 30.300 549.200 30.400 ;
        RECT 543.600 29.700 549.200 30.300 ;
        RECT 543.600 28.800 544.400 29.700 ;
        RECT 548.400 28.800 549.200 29.700 ;
        RECT 549.800 28.400 550.400 31.800 ;
        RECT 551.600 31.600 552.400 31.800 ;
        RECT 553.200 31.800 554.600 32.400 ;
        RECT 555.200 31.800 556.200 32.400 ;
        RECT 559.600 31.800 561.000 32.400 ;
        RECT 561.600 31.800 562.600 32.400 ;
        RECT 553.200 31.600 554.000 31.800 ;
        RECT 555.200 28.400 555.800 31.800 ;
        RECT 559.600 31.600 560.400 31.800 ;
        RECT 556.400 28.800 557.200 30.400 ;
        RECT 561.600 28.400 562.200 31.800 ;
        RECT 562.800 28.800 563.600 30.400 ;
        RECT 540.400 27.600 543.000 28.400 ;
        RECT 545.200 28.300 546.000 28.400 ;
        RECT 546.800 28.300 547.600 28.400 ;
        RECT 545.200 28.200 547.600 28.300 ;
        RECT 544.400 27.700 548.400 28.200 ;
        RECT 544.400 27.600 546.000 27.700 ;
        RECT 546.800 27.600 548.400 27.700 ;
        RECT 549.800 27.600 552.400 28.400 ;
        RECT 553.200 27.600 555.800 28.400 ;
        RECT 558.000 28.200 558.800 28.400 ;
        RECT 557.200 27.600 558.800 28.200 ;
        RECT 559.600 27.600 562.200 28.400 ;
        RECT 564.400 28.300 565.200 28.400 ;
        RECT 566.000 28.300 566.800 39.800 ;
        RECT 570.800 32.000 571.600 39.800 ;
        RECT 574.000 35.200 574.800 39.800 ;
        RECT 564.400 28.200 566.800 28.300 ;
        RECT 563.600 27.700 566.800 28.200 ;
        RECT 563.600 27.600 565.200 27.700 ;
        RECT 538.800 24.800 539.600 26.400 ;
        RECT 540.600 26.200 541.200 27.600 ;
        RECT 544.400 27.200 545.200 27.600 ;
        RECT 547.600 27.200 548.400 27.600 ;
        RECT 542.200 26.200 545.800 26.600 ;
        RECT 547.000 26.200 550.600 26.600 ;
        RECT 551.600 26.200 552.200 27.600 ;
        RECT 553.400 26.200 554.000 27.600 ;
        RECT 557.200 27.200 558.000 27.600 ;
        RECT 555.000 26.200 558.600 26.600 ;
        RECT 559.800 26.200 560.400 27.600 ;
        RECT 563.600 27.200 564.400 27.600 ;
        RECT 561.400 26.200 565.000 26.600 ;
        RECT 540.400 22.200 541.200 26.200 ;
        RECT 542.000 26.000 546.000 26.200 ;
        RECT 542.000 22.200 542.800 26.000 ;
        RECT 545.200 22.200 546.000 26.000 ;
        RECT 546.800 26.000 550.800 26.200 ;
        RECT 546.800 22.200 547.600 26.000 ;
        RECT 550.000 22.200 550.800 26.000 ;
        RECT 551.600 22.200 552.400 26.200 ;
        RECT 553.200 22.200 554.000 26.200 ;
        RECT 554.800 26.000 558.800 26.200 ;
        RECT 554.800 22.200 555.600 26.000 ;
        RECT 558.000 22.200 558.800 26.000 ;
        RECT 559.600 22.200 560.400 26.200 ;
        RECT 561.200 26.000 565.200 26.200 ;
        RECT 561.200 22.200 562.000 26.000 ;
        RECT 564.400 22.200 565.200 26.000 ;
        RECT 566.000 22.200 566.800 27.700 ;
        RECT 570.600 31.200 571.600 32.000 ;
        RECT 572.200 34.600 574.800 35.200 ;
        RECT 572.200 33.000 572.800 34.600 ;
        RECT 577.200 34.400 578.000 39.800 ;
        RECT 580.400 37.000 581.200 39.800 ;
        RECT 582.000 37.000 582.800 39.800 ;
        RECT 583.600 37.000 584.400 39.800 ;
        RECT 578.600 34.400 582.800 35.200 ;
        RECT 575.400 33.600 578.000 34.400 ;
        RECT 585.200 33.600 586.000 39.800 ;
        RECT 588.400 35.000 589.200 39.800 ;
        RECT 591.600 35.000 592.400 39.800 ;
        RECT 593.200 37.000 594.000 39.800 ;
        RECT 594.800 37.000 595.600 39.800 ;
        RECT 598.000 35.200 598.800 39.800 ;
        RECT 601.200 36.400 602.000 39.800 ;
        RECT 601.200 35.800 602.200 36.400 ;
        RECT 601.600 35.200 602.200 35.800 ;
        RECT 596.800 34.400 601.000 35.200 ;
        RECT 601.600 34.600 603.600 35.200 ;
        RECT 588.400 33.600 591.000 34.400 ;
        RECT 591.600 33.800 597.400 34.400 ;
        RECT 600.400 34.000 601.000 34.400 ;
        RECT 580.400 33.000 581.200 33.200 ;
        RECT 572.200 32.400 581.200 33.000 ;
        RECT 583.600 33.000 584.400 33.200 ;
        RECT 591.600 33.000 592.200 33.800 ;
        RECT 598.000 33.200 599.400 33.800 ;
        RECT 600.400 33.200 602.000 34.000 ;
        RECT 583.600 32.400 592.200 33.000 ;
        RECT 593.200 33.000 599.400 33.200 ;
        RECT 593.200 32.600 598.600 33.000 ;
        RECT 593.200 32.400 594.000 32.600 ;
        RECT 570.600 26.800 571.400 31.200 ;
        RECT 572.200 30.600 572.800 32.400 ;
        RECT 572.000 30.000 572.800 30.600 ;
        RECT 578.800 30.000 602.200 30.600 ;
        RECT 572.000 28.000 572.600 30.000 ;
        RECT 578.800 29.400 579.600 30.000 ;
        RECT 596.400 29.600 597.200 30.000 ;
        RECT 598.000 29.600 598.800 30.000 ;
        RECT 601.200 29.800 602.200 30.000 ;
        RECT 601.200 29.600 602.000 29.800 ;
        RECT 573.200 28.600 577.000 29.400 ;
        RECT 572.000 27.400 573.200 28.000 ;
        RECT 570.600 26.000 571.600 26.800 ;
        RECT 570.800 22.200 571.600 26.000 ;
        RECT 572.400 22.200 573.200 27.400 ;
        RECT 576.200 27.400 577.000 28.600 ;
        RECT 576.200 26.800 578.000 27.400 ;
        RECT 577.200 26.200 578.000 26.800 ;
        RECT 582.000 26.400 582.800 29.200 ;
        RECT 585.200 28.600 588.400 29.400 ;
        RECT 592.200 28.600 594.200 29.400 ;
        RECT 602.800 29.000 603.600 34.600 ;
        RECT 584.800 27.800 585.600 28.000 ;
        RECT 584.800 27.200 589.200 27.800 ;
        RECT 588.400 27.000 589.200 27.200 ;
        RECT 590.000 26.800 590.800 28.400 ;
        RECT 577.200 25.400 579.600 26.200 ;
        RECT 582.000 25.600 583.000 26.400 ;
        RECT 586.000 25.600 587.600 26.400 ;
        RECT 588.400 26.200 589.200 26.400 ;
        RECT 592.200 26.200 593.000 28.600 ;
        RECT 594.800 28.200 603.600 29.000 ;
        RECT 598.200 26.800 601.200 27.600 ;
        RECT 598.200 26.200 599.000 26.800 ;
        RECT 588.400 25.600 593.000 26.200 ;
        RECT 578.800 22.200 579.600 25.400 ;
        RECT 596.400 25.400 599.000 26.200 ;
        RECT 580.400 22.200 581.200 25.000 ;
        RECT 582.000 22.200 582.800 25.000 ;
        RECT 583.600 22.200 584.400 25.000 ;
        RECT 585.200 22.200 586.000 25.000 ;
        RECT 588.400 22.200 589.200 25.000 ;
        RECT 591.600 22.200 592.400 25.000 ;
        RECT 593.200 22.200 594.000 25.000 ;
        RECT 594.800 22.200 595.600 25.000 ;
        RECT 596.400 22.200 597.200 25.400 ;
        RECT 602.800 22.200 603.600 28.200 ;
        RECT 604.400 22.200 605.200 39.800 ;
        RECT 607.600 32.400 608.400 39.800 ;
        RECT 607.600 31.800 609.800 32.400 ;
        RECT 609.200 31.200 609.800 31.800 ;
        RECT 609.200 30.400 610.400 31.200 ;
        RECT 606.000 30.300 606.800 30.400 ;
        RECT 607.600 30.300 608.400 30.400 ;
        RECT 606.000 29.700 608.400 30.300 ;
        RECT 606.000 29.600 606.800 29.700 ;
        RECT 607.600 28.800 608.400 29.700 ;
        RECT 609.200 27.400 609.800 30.400 ;
        RECT 607.600 26.800 609.800 27.400 ;
        RECT 607.600 22.200 608.400 26.800 ;
        RECT 1.200 13.800 2.000 19.800 ;
        RECT 7.600 16.600 8.400 19.800 ;
        RECT 9.200 17.000 10.000 19.800 ;
        RECT 10.800 17.000 11.600 19.800 ;
        RECT 12.400 17.000 13.200 19.800 ;
        RECT 15.600 17.000 16.400 19.800 ;
        RECT 18.800 17.000 19.600 19.800 ;
        RECT 20.400 17.000 21.200 19.800 ;
        RECT 22.000 17.000 22.800 19.800 ;
        RECT 23.600 17.000 24.400 19.800 ;
        RECT 5.800 15.800 8.400 16.600 ;
        RECT 25.200 16.600 26.000 19.800 ;
        RECT 11.800 15.800 16.400 16.400 ;
        RECT 5.800 15.200 6.600 15.800 ;
        RECT 3.600 14.400 6.600 15.200 ;
        RECT 1.200 13.000 10.000 13.800 ;
        RECT 11.800 13.400 12.600 15.800 ;
        RECT 15.600 15.600 16.400 15.800 ;
        RECT 17.200 15.600 18.800 16.400 ;
        RECT 21.800 15.600 22.800 16.400 ;
        RECT 25.200 15.800 27.600 16.600 ;
        RECT 14.000 13.600 14.800 15.200 ;
        RECT 15.600 14.800 16.400 15.000 ;
        RECT 15.600 14.200 20.000 14.800 ;
        RECT 19.200 14.000 20.000 14.200 ;
        RECT 1.200 7.400 2.000 13.000 ;
        RECT 10.600 12.600 12.600 13.400 ;
        RECT 16.400 12.600 19.600 13.400 ;
        RECT 22.000 12.800 22.800 15.600 ;
        RECT 26.800 15.200 27.600 15.800 ;
        RECT 26.800 14.600 28.600 15.200 ;
        RECT 27.800 13.400 28.600 14.600 ;
        RECT 31.600 14.600 32.400 19.800 ;
        RECT 33.200 16.000 34.000 19.800 ;
        RECT 36.400 16.000 37.200 19.800 ;
        RECT 39.600 16.000 40.400 19.800 ;
        RECT 33.200 15.200 34.200 16.000 ;
        RECT 36.400 15.800 40.400 16.000 ;
        RECT 41.200 15.800 42.000 19.800 ;
        RECT 42.800 15.800 43.600 19.800 ;
        RECT 44.400 16.000 45.200 19.800 ;
        RECT 47.600 16.000 48.400 19.800 ;
        RECT 44.400 15.800 48.400 16.000 ;
        RECT 36.600 15.400 40.200 15.800 ;
        RECT 31.600 14.000 32.800 14.600 ;
        RECT 27.800 12.600 31.600 13.400 ;
        RECT 2.600 12.000 3.400 12.200 ;
        RECT 7.600 12.000 8.400 12.400 ;
        RECT 25.200 12.000 26.000 12.600 ;
        RECT 32.200 12.000 32.800 14.000 ;
        RECT 2.600 11.400 26.000 12.000 ;
        RECT 32.000 11.400 32.800 12.000 ;
        RECT 32.000 9.600 32.600 11.400 ;
        RECT 33.400 10.800 34.200 15.200 ;
        RECT 37.200 14.400 38.000 14.800 ;
        RECT 41.200 14.400 41.800 15.800 ;
        RECT 43.000 14.400 43.600 15.800 ;
        RECT 44.600 15.400 48.200 15.800 ;
        RECT 46.800 14.400 47.600 14.800 ;
        RECT 36.400 13.800 38.000 14.400 ;
        RECT 36.400 13.600 37.200 13.800 ;
        RECT 39.400 13.600 42.000 14.400 ;
        RECT 42.800 13.600 45.400 14.400 ;
        RECT 46.800 14.300 48.400 14.400 ;
        RECT 49.200 14.300 50.000 19.800 ;
        RECT 52.400 15.000 53.200 19.800 ;
        RECT 56.800 18.400 57.600 19.800 ;
        RECT 55.600 17.800 57.600 18.400 ;
        RECT 61.200 17.800 62.000 19.800 ;
        RECT 65.400 18.400 66.600 19.800 ;
        RECT 65.200 17.800 66.600 18.400 ;
        RECT 55.600 17.000 56.400 17.800 ;
        RECT 61.200 17.200 61.800 17.800 ;
        RECT 57.200 16.400 58.000 17.200 ;
        RECT 59.000 16.600 61.800 17.200 ;
        RECT 65.200 17.000 66.000 17.800 ;
        RECT 59.000 16.400 59.800 16.600 ;
        RECT 46.800 13.800 50.000 14.300 ;
        RECT 47.600 13.700 50.000 13.800 ;
        RECT 47.600 13.600 48.400 13.700 ;
        RECT 38.000 11.600 38.800 13.200 ;
        RECT 39.400 12.300 40.000 13.600 ;
        RECT 39.400 11.700 43.500 12.300 ;
        RECT 10.800 9.400 11.600 9.600 ;
        RECT 6.200 9.000 11.600 9.400 ;
        RECT 5.400 8.800 11.600 9.000 ;
        RECT 12.600 9.000 21.200 9.600 ;
        RECT 2.800 8.000 4.400 8.800 ;
        RECT 5.400 8.200 6.800 8.800 ;
        RECT 12.600 8.200 13.200 9.000 ;
        RECT 20.400 8.800 21.200 9.000 ;
        RECT 23.600 9.000 32.600 9.600 ;
        RECT 23.600 8.800 24.400 9.000 ;
        RECT 3.800 7.600 4.400 8.000 ;
        RECT 7.400 7.600 13.200 8.200 ;
        RECT 13.800 7.600 16.400 8.400 ;
        RECT 1.200 6.800 3.200 7.400 ;
        RECT 3.800 6.800 8.000 7.600 ;
        RECT 2.600 6.200 3.200 6.800 ;
        RECT 2.600 5.600 3.600 6.200 ;
        RECT 2.800 2.200 3.600 5.600 ;
        RECT 6.000 2.200 6.800 6.800 ;
        RECT 9.200 2.200 10.000 5.000 ;
        RECT 10.800 2.200 11.600 5.000 ;
        RECT 12.400 2.200 13.200 7.000 ;
        RECT 15.600 2.200 16.400 7.000 ;
        RECT 18.800 2.200 19.600 8.400 ;
        RECT 26.800 7.600 29.400 8.400 ;
        RECT 22.000 6.800 26.200 7.600 ;
        RECT 20.400 2.200 21.200 5.000 ;
        RECT 22.000 2.200 22.800 5.000 ;
        RECT 23.600 2.200 24.400 5.000 ;
        RECT 26.800 2.200 27.600 7.600 ;
        RECT 32.000 7.400 32.600 9.000 ;
        RECT 30.000 6.800 32.600 7.400 ;
        RECT 33.200 10.000 34.200 10.800 ;
        RECT 39.400 10.200 40.000 11.700 ;
        RECT 42.900 10.400 43.500 11.700 ;
        RECT 41.200 10.200 42.000 10.400 ;
        RECT 30.000 2.200 30.800 6.800 ;
        RECT 33.200 2.200 34.000 10.000 ;
        RECT 39.000 9.600 40.000 10.200 ;
        RECT 40.600 9.600 42.000 10.200 ;
        RECT 42.800 10.200 43.600 10.400 ;
        RECT 44.800 10.200 45.400 13.600 ;
        RECT 46.000 11.600 46.800 13.200 ;
        RECT 42.800 9.600 44.200 10.200 ;
        RECT 44.800 9.600 45.800 10.200 ;
        RECT 39.000 2.200 39.800 9.600 ;
        RECT 40.600 8.400 41.200 9.600 ;
        RECT 40.400 7.600 41.200 8.400 ;
        RECT 43.600 8.400 44.200 9.600 ;
        RECT 43.600 7.600 44.400 8.400 ;
        RECT 45.000 2.200 45.800 9.600 ;
        RECT 49.200 2.200 50.000 13.700 ;
        RECT 53.200 14.200 54.800 14.400 ;
        RECT 57.400 14.200 58.000 16.400 ;
        RECT 67.000 15.400 67.800 15.600 ;
        RECT 70.000 15.400 70.800 19.800 ;
        RECT 73.200 16.400 74.000 19.800 ;
        RECT 67.000 14.800 70.800 15.400 ;
        RECT 63.000 14.200 63.800 14.400 ;
        RECT 53.200 13.600 64.200 14.200 ;
        RECT 56.200 13.400 57.000 13.600 ;
        RECT 54.600 12.400 55.400 12.600 ;
        RECT 57.200 12.400 58.000 12.600 ;
        RECT 54.600 11.800 59.600 12.400 ;
        RECT 58.800 11.600 59.600 11.800 ;
        RECT 52.400 11.000 58.000 11.200 ;
        RECT 52.400 10.800 58.200 11.000 ;
        RECT 52.400 10.600 62.200 10.800 ;
        RECT 52.400 2.200 53.200 10.600 ;
        RECT 57.400 10.200 62.200 10.600 ;
        RECT 55.600 9.000 61.000 9.600 ;
        RECT 55.600 8.800 56.400 9.000 ;
        RECT 60.200 8.800 61.000 9.000 ;
        RECT 61.600 9.000 62.200 10.200 ;
        RECT 63.600 10.400 64.200 13.600 ;
        RECT 65.200 12.800 66.000 13.000 ;
        RECT 65.200 12.200 69.000 12.800 ;
        RECT 68.200 12.000 69.000 12.200 ;
        RECT 66.600 11.400 67.400 11.600 ;
        RECT 70.000 11.400 70.800 14.800 ;
        RECT 66.600 10.800 70.800 11.400 ;
        RECT 63.600 9.800 66.000 10.400 ;
        RECT 63.000 9.000 63.800 9.200 ;
        RECT 61.600 8.400 63.800 9.000 ;
        RECT 65.400 8.800 66.000 9.800 ;
        RECT 65.400 8.000 66.800 8.800 ;
        RECT 59.000 7.400 59.800 7.600 ;
        RECT 61.800 7.400 62.600 7.600 ;
        RECT 55.600 6.200 56.400 7.000 ;
        RECT 59.000 6.800 62.600 7.400 ;
        RECT 61.200 6.200 61.800 6.800 ;
        RECT 65.200 6.200 66.000 7.000 ;
        RECT 55.600 5.600 57.600 6.200 ;
        RECT 56.800 2.200 57.600 5.600 ;
        RECT 61.200 2.200 62.000 6.200 ;
        RECT 65.400 2.200 66.600 6.200 ;
        RECT 70.000 2.200 70.800 10.800 ;
        RECT 73.000 15.800 74.000 16.400 ;
        RECT 73.000 14.400 73.600 15.800 ;
        RECT 76.400 15.200 77.200 19.800 ;
        RECT 78.000 16.000 78.800 19.800 ;
        RECT 81.200 16.000 82.000 19.800 ;
        RECT 78.000 15.800 82.000 16.000 ;
        RECT 82.800 15.800 83.600 19.800 ;
        RECT 84.400 15.800 85.200 19.800 ;
        RECT 86.000 16.000 86.800 19.800 ;
        RECT 89.200 16.000 90.000 19.800 ;
        RECT 86.000 15.800 90.000 16.000 ;
        RECT 78.200 15.400 81.800 15.800 ;
        RECT 74.600 14.600 77.200 15.200 ;
        RECT 73.000 13.600 74.000 14.400 ;
        RECT 73.000 10.200 73.600 13.600 ;
        RECT 74.600 13.000 75.200 14.600 ;
        RECT 78.800 14.400 79.600 14.800 ;
        RECT 82.800 14.400 83.400 15.800 ;
        RECT 84.600 14.400 85.200 15.800 ;
        RECT 86.200 15.400 89.800 15.800 ;
        RECT 90.800 15.400 91.600 19.800 ;
        RECT 95.000 18.400 96.200 19.800 ;
        RECT 95.000 17.800 96.400 18.400 ;
        RECT 99.600 17.800 100.400 19.800 ;
        RECT 104.000 18.400 104.800 19.800 ;
        RECT 104.000 17.800 106.000 18.400 ;
        RECT 95.600 17.000 96.400 17.800 ;
        RECT 99.800 17.200 100.400 17.800 ;
        RECT 99.800 16.600 102.600 17.200 ;
        RECT 101.800 16.400 102.600 16.600 ;
        RECT 103.600 16.400 104.400 17.200 ;
        RECT 105.200 17.000 106.000 17.800 ;
        RECT 93.800 15.400 94.600 15.600 ;
        RECT 90.800 14.800 94.600 15.400 ;
        RECT 88.400 14.400 89.200 14.800 ;
        RECT 78.000 13.800 79.600 14.400 ;
        RECT 78.000 13.600 78.800 13.800 ;
        RECT 81.000 13.600 83.600 14.400 ;
        RECT 84.400 13.600 87.000 14.400 ;
        RECT 88.400 13.800 90.000 14.400 ;
        RECT 89.200 13.600 90.000 13.800 ;
        RECT 74.200 12.200 75.200 13.000 ;
        RECT 74.600 10.200 75.200 12.200 ;
        RECT 76.200 12.400 77.000 13.200 ;
        RECT 76.200 12.300 77.200 12.400 ;
        RECT 78.000 12.300 78.800 12.400 ;
        RECT 76.200 11.700 78.800 12.300 ;
        RECT 76.200 11.600 77.200 11.700 ;
        RECT 78.000 11.600 78.800 11.700 ;
        RECT 79.600 11.600 80.400 13.200 ;
        RECT 81.000 10.200 81.600 13.600 ;
        RECT 86.400 12.300 87.000 13.600 ;
        RECT 82.900 11.700 87.000 12.300 ;
        RECT 82.900 10.400 83.500 11.700 ;
        RECT 82.800 10.200 83.600 10.400 ;
        RECT 73.000 9.200 74.000 10.200 ;
        RECT 74.600 9.600 77.200 10.200 ;
        RECT 73.200 2.200 74.000 9.200 ;
        RECT 76.400 2.200 77.200 9.600 ;
        RECT 80.600 9.600 81.600 10.200 ;
        RECT 82.200 9.600 83.600 10.200 ;
        RECT 84.400 10.200 85.200 10.400 ;
        RECT 86.400 10.200 87.000 11.700 ;
        RECT 87.600 11.600 88.400 13.200 ;
        RECT 90.800 11.400 91.600 14.800 ;
        RECT 97.800 14.200 98.600 14.400 ;
        RECT 100.400 14.200 101.200 14.400 ;
        RECT 103.600 14.200 104.200 16.400 ;
        RECT 108.400 15.000 109.200 19.800 ;
        RECT 110.000 15.400 110.800 19.800 ;
        RECT 114.200 18.400 115.400 19.800 ;
        RECT 114.200 17.800 115.600 18.400 ;
        RECT 118.800 17.800 119.600 19.800 ;
        RECT 123.200 18.400 124.000 19.800 ;
        RECT 123.200 17.800 125.200 18.400 ;
        RECT 114.800 17.000 115.600 17.800 ;
        RECT 119.000 17.200 119.600 17.800 ;
        RECT 119.000 16.600 121.800 17.200 ;
        RECT 121.000 16.400 121.800 16.600 ;
        RECT 122.800 16.400 123.600 17.200 ;
        RECT 124.400 17.000 125.200 17.800 ;
        RECT 113.000 15.400 113.800 15.600 ;
        RECT 110.000 14.800 113.800 15.400 ;
        RECT 106.800 14.200 108.400 14.400 ;
        RECT 97.400 13.600 108.400 14.200 ;
        RECT 95.600 12.800 96.400 13.000 ;
        RECT 92.600 12.200 96.400 12.800 ;
        RECT 92.600 12.000 93.400 12.200 ;
        RECT 94.200 11.400 95.000 11.600 ;
        RECT 90.800 10.800 95.000 11.400 ;
        RECT 84.400 9.600 85.800 10.200 ;
        RECT 86.400 9.600 87.400 10.200 ;
        RECT 80.600 2.200 81.400 9.600 ;
        RECT 82.200 8.400 82.800 9.600 ;
        RECT 82.000 7.600 82.800 8.400 ;
        RECT 85.200 8.400 85.800 9.600 ;
        RECT 85.200 7.600 86.000 8.400 ;
        RECT 86.600 2.200 87.400 9.600 ;
        RECT 90.800 2.200 91.600 10.800 ;
        RECT 97.400 10.400 98.000 13.600 ;
        RECT 104.600 13.400 105.400 13.600 ;
        RECT 106.200 12.400 107.000 12.600 ;
        RECT 102.000 11.800 107.000 12.400 ;
        RECT 102.000 11.600 102.800 11.800 ;
        RECT 110.000 11.400 110.800 14.800 ;
        RECT 117.000 14.200 117.800 14.400 ;
        RECT 122.800 14.200 123.400 16.400 ;
        RECT 127.600 15.000 128.400 19.800 ;
        RECT 130.800 16.400 131.600 19.800 ;
        RECT 130.600 15.800 131.600 16.400 ;
        RECT 130.600 14.400 131.200 15.800 ;
        RECT 134.000 15.200 134.800 19.800 ;
        RECT 138.800 15.200 139.600 19.800 ;
        RECT 146.800 16.000 147.600 19.800 ;
        RECT 132.200 14.600 134.800 15.200 ;
        RECT 137.400 14.600 139.600 15.200 ;
        RECT 146.600 15.200 147.600 16.000 ;
        RECT 126.000 14.300 127.600 14.400 ;
        RECT 129.200 14.300 130.000 14.400 ;
        RECT 126.000 14.200 130.000 14.300 ;
        RECT 116.600 13.700 130.000 14.200 ;
        RECT 116.600 13.600 127.600 13.700 ;
        RECT 129.200 13.600 130.000 13.700 ;
        RECT 130.600 13.600 131.600 14.400 ;
        RECT 114.800 12.800 115.600 13.000 ;
        RECT 111.800 12.200 115.600 12.800 ;
        RECT 116.600 12.400 117.200 13.600 ;
        RECT 123.800 13.400 124.600 13.600 ;
        RECT 122.800 12.400 123.600 12.600 ;
        RECT 125.400 12.400 126.200 12.600 ;
        RECT 111.800 12.000 112.600 12.200 ;
        RECT 116.400 11.600 117.200 12.400 ;
        RECT 121.200 11.800 126.200 12.400 ;
        RECT 121.200 11.600 122.000 11.800 ;
        RECT 113.400 11.400 114.200 11.600 ;
        RECT 103.600 11.000 109.200 11.200 ;
        RECT 103.400 10.800 109.200 11.000 ;
        RECT 95.600 9.800 98.000 10.400 ;
        RECT 99.400 10.600 109.200 10.800 ;
        RECT 99.400 10.200 104.200 10.600 ;
        RECT 95.600 8.800 96.200 9.800 ;
        RECT 94.800 8.000 96.200 8.800 ;
        RECT 97.800 9.000 98.600 9.200 ;
        RECT 99.400 9.000 100.000 10.200 ;
        RECT 97.800 8.400 100.000 9.000 ;
        RECT 100.600 9.000 106.000 9.600 ;
        RECT 100.600 8.800 101.400 9.000 ;
        RECT 105.200 8.800 106.000 9.000 ;
        RECT 99.000 7.400 99.800 7.600 ;
        RECT 101.800 7.400 102.600 7.600 ;
        RECT 95.600 6.200 96.400 7.000 ;
        RECT 99.000 6.800 102.600 7.400 ;
        RECT 99.800 6.200 100.400 6.800 ;
        RECT 105.200 6.200 106.000 7.000 ;
        RECT 95.000 2.200 96.200 6.200 ;
        RECT 99.600 2.200 100.400 6.200 ;
        RECT 104.000 5.600 106.000 6.200 ;
        RECT 104.000 2.200 104.800 5.600 ;
        RECT 108.400 2.200 109.200 10.600 ;
        RECT 110.000 10.800 114.200 11.400 ;
        RECT 110.000 2.200 110.800 10.800 ;
        RECT 116.600 10.400 117.200 11.600 ;
        RECT 122.800 11.000 128.400 11.200 ;
        RECT 122.600 10.800 128.400 11.000 ;
        RECT 114.800 9.800 117.200 10.400 ;
        RECT 118.600 10.600 128.400 10.800 ;
        RECT 118.600 10.200 123.400 10.600 ;
        RECT 114.800 8.800 115.400 9.800 ;
        RECT 114.000 8.000 115.400 8.800 ;
        RECT 117.000 9.000 117.800 9.200 ;
        RECT 118.600 9.000 119.200 10.200 ;
        RECT 117.000 8.400 119.200 9.000 ;
        RECT 119.800 9.000 125.200 9.600 ;
        RECT 119.800 8.800 120.600 9.000 ;
        RECT 124.400 8.800 125.200 9.000 ;
        RECT 118.200 7.400 119.000 7.600 ;
        RECT 121.000 7.400 121.800 7.600 ;
        RECT 114.800 6.200 115.600 7.000 ;
        RECT 118.200 6.800 121.800 7.400 ;
        RECT 119.000 6.200 119.600 6.800 ;
        RECT 124.400 6.200 125.200 7.000 ;
        RECT 114.200 2.200 115.400 6.200 ;
        RECT 118.800 2.200 119.600 6.200 ;
        RECT 123.200 5.600 125.200 6.200 ;
        RECT 123.200 2.200 124.000 5.600 ;
        RECT 127.600 2.200 128.400 10.600 ;
        RECT 130.600 10.200 131.200 13.600 ;
        RECT 132.200 13.000 132.800 14.600 ;
        RECT 131.800 12.200 132.800 13.000 ;
        RECT 132.200 10.200 132.800 12.200 ;
        RECT 133.800 12.400 134.600 13.200 ;
        RECT 133.800 11.600 134.800 12.400 ;
        RECT 137.400 11.600 138.000 14.600 ;
        RECT 138.800 12.300 139.600 13.200 ;
        RECT 146.600 12.300 147.400 15.200 ;
        RECT 148.400 14.600 149.200 19.800 ;
        RECT 154.800 16.600 155.600 19.800 ;
        RECT 156.400 17.000 157.200 19.800 ;
        RECT 158.000 17.000 158.800 19.800 ;
        RECT 159.600 17.000 160.400 19.800 ;
        RECT 161.200 17.000 162.000 19.800 ;
        RECT 164.400 17.000 165.200 19.800 ;
        RECT 167.600 17.000 168.400 19.800 ;
        RECT 169.200 17.000 170.000 19.800 ;
        RECT 170.800 17.000 171.600 19.800 ;
        RECT 153.200 15.800 155.600 16.600 ;
        RECT 172.400 16.600 173.200 19.800 ;
        RECT 153.200 15.200 154.000 15.800 ;
        RECT 138.800 11.700 147.400 12.300 ;
        RECT 138.800 11.600 139.600 11.700 ;
        RECT 136.800 10.800 138.000 11.600 ;
        RECT 137.400 10.200 138.000 10.800 ;
        RECT 146.600 10.800 147.400 11.700 ;
        RECT 148.000 14.000 149.200 14.600 ;
        RECT 152.200 14.600 154.000 15.200 ;
        RECT 158.000 15.600 159.000 16.400 ;
        RECT 162.000 15.600 163.600 16.400 ;
        RECT 164.400 15.800 169.000 16.400 ;
        RECT 172.400 15.800 175.000 16.600 ;
        RECT 164.400 15.600 165.200 15.800 ;
        RECT 148.000 12.000 148.600 14.000 ;
        RECT 152.200 13.400 153.000 14.600 ;
        RECT 149.200 12.600 153.000 13.400 ;
        RECT 158.000 12.800 158.800 15.600 ;
        RECT 164.400 14.800 165.200 15.000 ;
        RECT 160.800 14.200 165.200 14.800 ;
        RECT 160.800 14.000 161.600 14.200 ;
        RECT 166.000 13.600 166.800 15.200 ;
        RECT 168.200 13.400 169.000 15.800 ;
        RECT 174.200 15.200 175.000 15.800 ;
        RECT 174.200 14.400 177.200 15.200 ;
        RECT 178.800 13.800 179.600 19.800 ;
        RECT 161.200 12.600 164.400 13.400 ;
        RECT 168.200 12.600 170.200 13.400 ;
        RECT 170.800 13.000 179.600 13.800 ;
        RECT 154.800 12.000 155.600 12.600 ;
        RECT 172.400 12.000 173.200 12.400 ;
        RECT 177.200 12.200 178.000 12.400 ;
        RECT 177.200 12.000 178.200 12.200 ;
        RECT 148.000 11.400 148.800 12.000 ;
        RECT 154.800 11.400 178.200 12.000 ;
        RECT 130.600 9.200 131.600 10.200 ;
        RECT 132.200 9.600 134.800 10.200 ;
        RECT 137.400 9.600 139.600 10.200 ;
        RECT 146.600 10.000 147.600 10.800 ;
        RECT 130.800 2.200 131.600 9.200 ;
        RECT 134.000 2.200 134.800 9.600 ;
        RECT 138.800 2.200 139.600 9.600 ;
        RECT 146.800 2.200 147.600 10.000 ;
        RECT 148.200 9.600 148.800 11.400 ;
        RECT 148.200 9.000 157.200 9.600 ;
        RECT 148.200 7.400 148.800 9.000 ;
        RECT 156.400 8.800 157.200 9.000 ;
        RECT 159.600 9.000 168.200 9.600 ;
        RECT 159.600 8.800 160.400 9.000 ;
        RECT 151.400 7.600 154.000 8.400 ;
        RECT 148.200 6.800 150.800 7.400 ;
        RECT 150.000 2.200 150.800 6.800 ;
        RECT 153.200 2.200 154.000 7.600 ;
        RECT 154.600 6.800 158.800 7.600 ;
        RECT 156.400 2.200 157.200 5.000 ;
        RECT 158.000 2.200 158.800 5.000 ;
        RECT 159.600 2.200 160.400 5.000 ;
        RECT 161.200 2.200 162.000 8.400 ;
        RECT 164.400 7.600 167.000 8.400 ;
        RECT 167.600 8.200 168.200 9.000 ;
        RECT 169.200 9.400 170.000 9.600 ;
        RECT 169.200 9.000 174.600 9.400 ;
        RECT 169.200 8.800 175.400 9.000 ;
        RECT 174.000 8.200 175.400 8.800 ;
        RECT 167.600 7.600 173.400 8.200 ;
        RECT 176.400 8.000 178.000 8.800 ;
        RECT 176.400 7.600 177.000 8.000 ;
        RECT 164.400 2.200 165.200 7.000 ;
        RECT 167.600 2.200 168.400 7.000 ;
        RECT 172.800 6.800 177.000 7.600 ;
        RECT 178.800 7.400 179.600 13.000 ;
        RECT 177.600 6.800 179.600 7.400 ;
        RECT 180.400 13.800 181.200 19.800 ;
        RECT 186.800 16.600 187.600 19.800 ;
        RECT 188.400 17.000 189.200 19.800 ;
        RECT 190.000 17.000 190.800 19.800 ;
        RECT 191.600 17.000 192.400 19.800 ;
        RECT 194.800 17.000 195.600 19.800 ;
        RECT 198.000 17.000 198.800 19.800 ;
        RECT 199.600 17.000 200.400 19.800 ;
        RECT 201.200 17.000 202.000 19.800 ;
        RECT 202.800 17.000 203.600 19.800 ;
        RECT 185.000 15.800 187.600 16.600 ;
        RECT 204.400 16.600 205.200 19.800 ;
        RECT 191.000 15.800 195.600 16.400 ;
        RECT 185.000 15.200 185.800 15.800 ;
        RECT 182.800 14.400 185.800 15.200 ;
        RECT 180.400 13.000 189.200 13.800 ;
        RECT 191.000 13.400 191.800 15.800 ;
        RECT 194.800 15.600 195.600 15.800 ;
        RECT 196.400 15.600 198.000 16.400 ;
        RECT 201.000 15.600 202.000 16.400 ;
        RECT 204.400 15.800 206.800 16.600 ;
        RECT 193.200 13.600 194.000 15.200 ;
        RECT 194.800 14.800 195.600 15.000 ;
        RECT 194.800 14.200 199.200 14.800 ;
        RECT 198.400 14.000 199.200 14.200 ;
        RECT 180.400 7.400 181.200 13.000 ;
        RECT 189.800 12.600 191.800 13.400 ;
        RECT 195.600 12.600 198.800 13.400 ;
        RECT 201.200 12.800 202.000 15.600 ;
        RECT 206.000 15.200 206.800 15.800 ;
        RECT 206.000 14.600 207.800 15.200 ;
        RECT 207.000 13.400 207.800 14.600 ;
        RECT 210.800 14.600 211.600 19.800 ;
        RECT 212.400 16.000 213.200 19.800 ;
        RECT 212.400 15.200 213.400 16.000 ;
        RECT 210.800 14.000 212.000 14.600 ;
        RECT 207.000 12.600 210.800 13.400 ;
        RECT 181.800 12.000 182.600 12.200 ;
        RECT 183.600 12.000 184.400 12.400 ;
        RECT 186.800 12.000 187.600 12.400 ;
        RECT 204.400 12.000 205.200 12.600 ;
        RECT 211.400 12.000 212.000 14.000 ;
        RECT 181.800 11.400 205.200 12.000 ;
        RECT 211.200 11.400 212.000 12.000 ;
        RECT 212.600 12.300 213.400 15.200 ;
        RECT 215.600 15.200 216.400 19.800 ;
        RECT 215.600 14.600 217.800 15.200 ;
        RECT 215.600 12.300 216.400 13.200 ;
        RECT 212.600 11.700 216.400 12.300 ;
        RECT 211.200 9.600 211.800 11.400 ;
        RECT 212.600 10.800 213.400 11.700 ;
        RECT 215.600 11.600 216.400 11.700 ;
        RECT 217.200 11.600 217.800 14.600 ;
        RECT 220.400 13.800 221.200 19.800 ;
        RECT 226.800 16.600 227.600 19.800 ;
        RECT 228.400 17.000 229.200 19.800 ;
        RECT 230.000 17.000 230.800 19.800 ;
        RECT 231.600 17.000 232.400 19.800 ;
        RECT 234.800 17.000 235.600 19.800 ;
        RECT 238.000 17.000 238.800 19.800 ;
        RECT 239.600 17.000 240.400 19.800 ;
        RECT 241.200 17.000 242.000 19.800 ;
        RECT 242.800 17.000 243.600 19.800 ;
        RECT 225.000 15.800 227.600 16.600 ;
        RECT 244.400 16.600 245.200 19.800 ;
        RECT 231.000 15.800 235.600 16.400 ;
        RECT 225.000 15.200 225.800 15.800 ;
        RECT 222.800 14.400 225.800 15.200 ;
        RECT 220.400 13.000 229.200 13.800 ;
        RECT 231.000 13.400 231.800 15.800 ;
        RECT 234.800 15.600 235.600 15.800 ;
        RECT 236.400 15.600 238.000 16.400 ;
        RECT 241.000 15.600 242.000 16.400 ;
        RECT 244.400 15.800 246.800 16.600 ;
        RECT 233.200 13.600 234.000 15.200 ;
        RECT 234.800 14.800 235.600 15.000 ;
        RECT 234.800 14.200 239.200 14.800 ;
        RECT 238.400 14.000 239.200 14.200 ;
        RECT 190.000 9.400 190.800 9.600 ;
        RECT 185.400 9.000 190.800 9.400 ;
        RECT 184.600 8.800 190.800 9.000 ;
        RECT 191.800 9.000 200.400 9.600 ;
        RECT 182.000 8.000 183.600 8.800 ;
        RECT 184.600 8.200 186.000 8.800 ;
        RECT 191.800 8.200 192.400 9.000 ;
        RECT 199.600 8.800 200.400 9.000 ;
        RECT 202.800 9.000 211.800 9.600 ;
        RECT 202.800 8.800 203.600 9.000 ;
        RECT 183.000 7.600 183.600 8.000 ;
        RECT 186.600 7.600 192.400 8.200 ;
        RECT 193.000 7.600 195.600 8.400 ;
        RECT 180.400 6.800 182.400 7.400 ;
        RECT 183.000 6.800 187.200 7.600 ;
        RECT 169.200 2.200 170.000 5.000 ;
        RECT 170.800 2.200 171.600 5.000 ;
        RECT 174.000 2.200 174.800 6.800 ;
        RECT 177.600 6.200 178.200 6.800 ;
        RECT 177.200 5.600 178.200 6.200 ;
        RECT 181.800 6.200 182.400 6.800 ;
        RECT 181.800 5.600 182.800 6.200 ;
        RECT 177.200 2.200 178.000 5.600 ;
        RECT 182.000 2.200 182.800 5.600 ;
        RECT 185.200 2.200 186.000 6.800 ;
        RECT 188.400 2.200 189.200 5.000 ;
        RECT 190.000 2.200 190.800 5.000 ;
        RECT 191.600 2.200 192.400 7.000 ;
        RECT 194.800 2.200 195.600 7.000 ;
        RECT 198.000 2.200 198.800 8.400 ;
        RECT 206.000 7.600 208.600 8.400 ;
        RECT 201.200 6.800 205.400 7.600 ;
        RECT 199.600 2.200 200.400 5.000 ;
        RECT 201.200 2.200 202.000 5.000 ;
        RECT 202.800 2.200 203.600 5.000 ;
        RECT 206.000 2.200 206.800 7.600 ;
        RECT 211.200 7.400 211.800 9.000 ;
        RECT 209.200 6.800 211.800 7.400 ;
        RECT 212.400 10.000 213.400 10.800 ;
        RECT 217.200 10.800 218.400 11.600 ;
        RECT 217.200 10.200 217.800 10.800 ;
        RECT 209.200 2.200 210.000 6.800 ;
        RECT 212.400 2.200 213.200 10.000 ;
        RECT 215.600 9.600 217.800 10.200 ;
        RECT 215.600 2.200 216.400 9.600 ;
        RECT 220.400 7.400 221.200 13.000 ;
        RECT 229.800 12.600 231.800 13.400 ;
        RECT 235.600 12.600 238.800 13.400 ;
        RECT 241.200 12.800 242.000 15.600 ;
        RECT 246.000 15.200 246.800 15.800 ;
        RECT 246.000 14.600 247.800 15.200 ;
        RECT 247.000 13.400 247.800 14.600 ;
        RECT 250.800 14.600 251.600 19.800 ;
        RECT 252.400 16.000 253.200 19.800 ;
        RECT 252.400 15.200 253.400 16.000 ;
        RECT 250.800 14.000 252.000 14.600 ;
        RECT 247.000 12.600 250.800 13.400 ;
        RECT 221.800 12.000 222.600 12.200 ;
        RECT 223.600 12.000 224.400 12.400 ;
        RECT 226.800 12.000 227.600 12.400 ;
        RECT 244.400 12.000 245.200 12.600 ;
        RECT 251.400 12.000 252.000 14.000 ;
        RECT 221.800 11.400 245.200 12.000 ;
        RECT 251.200 11.400 252.000 12.000 ;
        RECT 252.600 12.300 253.400 15.200 ;
        RECT 255.600 15.200 256.400 19.800 ;
        RECT 260.400 15.200 261.200 19.800 ;
        RECT 265.200 15.200 266.000 19.800 ;
        RECT 255.600 14.600 257.800 15.200 ;
        RECT 260.400 14.600 262.600 15.200 ;
        RECT 265.200 14.600 267.400 15.200 ;
        RECT 255.600 12.300 256.400 13.200 ;
        RECT 252.600 11.700 256.400 12.300 ;
        RECT 251.200 9.600 251.800 11.400 ;
        RECT 252.600 10.800 253.400 11.700 ;
        RECT 255.600 11.600 256.400 11.700 ;
        RECT 257.200 11.600 257.800 14.600 ;
        RECT 260.400 11.600 261.200 13.200 ;
        RECT 262.000 11.600 262.600 14.600 ;
        RECT 265.200 11.600 266.000 13.200 ;
        RECT 266.800 11.600 267.400 14.600 ;
        RECT 270.000 13.800 270.800 19.800 ;
        RECT 276.400 16.600 277.200 19.800 ;
        RECT 278.000 17.000 278.800 19.800 ;
        RECT 279.600 17.000 280.400 19.800 ;
        RECT 281.200 17.000 282.000 19.800 ;
        RECT 284.400 17.000 285.200 19.800 ;
        RECT 287.600 17.000 288.400 19.800 ;
        RECT 289.200 17.000 290.000 19.800 ;
        RECT 290.800 17.000 291.600 19.800 ;
        RECT 292.400 17.000 293.200 19.800 ;
        RECT 274.600 15.800 277.200 16.600 ;
        RECT 294.000 16.600 294.800 19.800 ;
        RECT 280.600 15.800 285.200 16.400 ;
        RECT 274.600 15.200 275.400 15.800 ;
        RECT 272.400 14.400 275.400 15.200 ;
        RECT 270.000 13.000 278.800 13.800 ;
        RECT 280.600 13.400 281.400 15.800 ;
        RECT 284.400 15.600 285.200 15.800 ;
        RECT 286.000 15.600 287.600 16.400 ;
        RECT 290.600 15.600 291.600 16.400 ;
        RECT 294.000 15.800 296.400 16.600 ;
        RECT 282.800 13.600 283.600 15.200 ;
        RECT 284.400 14.800 285.200 15.000 ;
        RECT 284.400 14.200 288.800 14.800 ;
        RECT 288.000 14.000 288.800 14.200 ;
        RECT 230.000 9.400 230.800 9.600 ;
        RECT 225.400 9.000 230.800 9.400 ;
        RECT 224.600 8.800 230.800 9.000 ;
        RECT 231.800 9.000 240.400 9.600 ;
        RECT 222.000 8.000 223.600 8.800 ;
        RECT 224.600 8.200 226.000 8.800 ;
        RECT 231.800 8.200 232.400 9.000 ;
        RECT 239.600 8.800 240.400 9.000 ;
        RECT 242.800 9.000 251.800 9.600 ;
        RECT 242.800 8.800 243.600 9.000 ;
        RECT 223.000 7.600 223.600 8.000 ;
        RECT 226.600 7.600 232.400 8.200 ;
        RECT 233.000 7.600 235.600 8.400 ;
        RECT 220.400 6.800 222.400 7.400 ;
        RECT 223.000 6.800 227.200 7.600 ;
        RECT 221.800 6.200 222.400 6.800 ;
        RECT 221.800 5.600 222.800 6.200 ;
        RECT 222.000 2.200 222.800 5.600 ;
        RECT 225.200 2.200 226.000 6.800 ;
        RECT 228.400 2.200 229.200 5.000 ;
        RECT 230.000 2.200 230.800 5.000 ;
        RECT 231.600 2.200 232.400 7.000 ;
        RECT 234.800 2.200 235.600 7.000 ;
        RECT 238.000 2.200 238.800 8.400 ;
        RECT 246.000 7.600 248.600 8.400 ;
        RECT 241.200 6.800 245.400 7.600 ;
        RECT 239.600 2.200 240.400 5.000 ;
        RECT 241.200 2.200 242.000 5.000 ;
        RECT 242.800 2.200 243.600 5.000 ;
        RECT 246.000 2.200 246.800 7.600 ;
        RECT 251.200 7.400 251.800 9.000 ;
        RECT 249.200 6.800 251.800 7.400 ;
        RECT 252.400 10.000 253.400 10.800 ;
        RECT 257.200 10.800 258.400 11.600 ;
        RECT 262.000 10.800 263.200 11.600 ;
        RECT 266.800 10.800 268.000 11.600 ;
        RECT 257.200 10.200 257.800 10.800 ;
        RECT 262.000 10.200 262.600 10.800 ;
        RECT 266.800 10.200 267.400 10.800 ;
        RECT 249.200 2.200 250.000 6.800 ;
        RECT 252.400 2.200 253.200 10.000 ;
        RECT 255.600 9.600 257.800 10.200 ;
        RECT 260.400 9.600 262.600 10.200 ;
        RECT 265.200 9.600 267.400 10.200 ;
        RECT 255.600 2.200 256.400 9.600 ;
        RECT 260.400 2.200 261.200 9.600 ;
        RECT 265.200 2.200 266.000 9.600 ;
        RECT 270.000 7.400 270.800 13.000 ;
        RECT 279.400 12.600 281.400 13.400 ;
        RECT 285.200 12.600 288.400 13.400 ;
        RECT 290.800 12.800 291.600 15.600 ;
        RECT 295.600 15.200 296.400 15.800 ;
        RECT 295.600 14.600 297.400 15.200 ;
        RECT 296.600 13.400 297.400 14.600 ;
        RECT 300.400 14.600 301.200 19.800 ;
        RECT 302.000 16.000 302.800 19.800 ;
        RECT 302.000 15.200 303.000 16.000 ;
        RECT 300.400 14.000 301.600 14.600 ;
        RECT 296.600 12.600 300.400 13.400 ;
        RECT 271.400 12.000 272.200 12.200 ;
        RECT 273.200 12.000 274.000 12.400 ;
        RECT 276.400 12.000 277.200 12.400 ;
        RECT 294.000 12.000 294.800 12.600 ;
        RECT 301.000 12.000 301.600 14.000 ;
        RECT 271.400 11.400 294.800 12.000 ;
        RECT 300.800 11.400 301.600 12.000 ;
        RECT 302.200 12.300 303.000 15.200 ;
        RECT 310.000 15.200 310.800 19.800 ;
        RECT 310.000 14.600 312.200 15.200 ;
        RECT 310.000 12.300 310.800 13.200 ;
        RECT 302.200 11.700 310.800 12.300 ;
        RECT 300.800 9.600 301.400 11.400 ;
        RECT 302.200 10.800 303.000 11.700 ;
        RECT 310.000 11.600 310.800 11.700 ;
        RECT 311.600 11.600 312.200 14.600 ;
        RECT 314.800 13.800 315.600 19.800 ;
        RECT 321.200 16.600 322.000 19.800 ;
        RECT 322.800 17.000 323.600 19.800 ;
        RECT 324.400 17.000 325.200 19.800 ;
        RECT 326.000 17.000 326.800 19.800 ;
        RECT 329.200 17.000 330.000 19.800 ;
        RECT 332.400 17.000 333.200 19.800 ;
        RECT 334.000 17.000 334.800 19.800 ;
        RECT 335.600 17.000 336.400 19.800 ;
        RECT 337.200 17.000 338.000 19.800 ;
        RECT 319.400 15.800 322.000 16.600 ;
        RECT 338.800 16.600 339.600 19.800 ;
        RECT 325.400 15.800 330.000 16.400 ;
        RECT 319.400 15.200 320.200 15.800 ;
        RECT 317.200 14.400 320.200 15.200 ;
        RECT 314.800 13.000 323.600 13.800 ;
        RECT 325.400 13.400 326.200 15.800 ;
        RECT 329.200 15.600 330.000 15.800 ;
        RECT 330.800 15.600 332.400 16.400 ;
        RECT 335.400 15.600 336.400 16.400 ;
        RECT 338.800 15.800 341.200 16.600 ;
        RECT 327.600 13.600 328.400 15.200 ;
        RECT 329.200 14.800 330.000 15.000 ;
        RECT 329.200 14.200 333.600 14.800 ;
        RECT 332.800 14.000 333.600 14.200 ;
        RECT 279.600 9.400 280.400 9.600 ;
        RECT 275.000 9.000 280.400 9.400 ;
        RECT 274.200 8.800 280.400 9.000 ;
        RECT 281.400 9.000 290.000 9.600 ;
        RECT 271.600 8.000 273.200 8.800 ;
        RECT 274.200 8.200 275.600 8.800 ;
        RECT 281.400 8.200 282.000 9.000 ;
        RECT 289.200 8.800 290.000 9.000 ;
        RECT 292.400 9.000 301.400 9.600 ;
        RECT 292.400 8.800 293.200 9.000 ;
        RECT 272.600 7.600 273.200 8.000 ;
        RECT 276.200 7.600 282.000 8.200 ;
        RECT 282.600 7.600 285.200 8.400 ;
        RECT 270.000 6.800 272.000 7.400 ;
        RECT 272.600 6.800 276.800 7.600 ;
        RECT 271.400 6.200 272.000 6.800 ;
        RECT 271.400 5.600 272.400 6.200 ;
        RECT 271.600 2.200 272.400 5.600 ;
        RECT 274.800 2.200 275.600 6.800 ;
        RECT 278.000 2.200 278.800 5.000 ;
        RECT 279.600 2.200 280.400 5.000 ;
        RECT 281.200 2.200 282.000 7.000 ;
        RECT 284.400 2.200 285.200 7.000 ;
        RECT 287.600 2.200 288.400 8.400 ;
        RECT 295.600 7.600 298.200 8.400 ;
        RECT 290.800 6.800 295.000 7.600 ;
        RECT 289.200 2.200 290.000 5.000 ;
        RECT 290.800 2.200 291.600 5.000 ;
        RECT 292.400 2.200 293.200 5.000 ;
        RECT 295.600 2.200 296.400 7.600 ;
        RECT 300.800 7.400 301.400 9.000 ;
        RECT 298.800 6.800 301.400 7.400 ;
        RECT 302.000 10.000 303.000 10.800 ;
        RECT 311.600 10.800 312.800 11.600 ;
        RECT 311.600 10.200 312.200 10.800 ;
        RECT 298.800 2.200 299.600 6.800 ;
        RECT 302.000 2.200 302.800 10.000 ;
        RECT 310.000 9.600 312.200 10.200 ;
        RECT 310.000 2.200 310.800 9.600 ;
        RECT 314.800 7.400 315.600 13.000 ;
        RECT 324.200 12.600 326.200 13.400 ;
        RECT 330.000 12.600 333.200 13.400 ;
        RECT 335.600 12.800 336.400 15.600 ;
        RECT 340.400 15.200 341.200 15.800 ;
        RECT 340.400 14.600 342.200 15.200 ;
        RECT 341.400 13.400 342.200 14.600 ;
        RECT 345.200 14.600 346.000 19.800 ;
        RECT 346.800 16.300 347.600 19.800 ;
        RECT 351.600 17.800 352.400 19.800 ;
        RECT 350.000 16.300 350.800 17.200 ;
        RECT 346.800 15.700 350.800 16.300 ;
        RECT 346.800 15.200 347.800 15.700 ;
        RECT 350.000 15.600 350.800 15.700 ;
        RECT 351.800 15.600 352.400 17.800 ;
        RECT 354.800 16.300 355.600 19.800 ;
        RECT 358.000 17.800 358.800 19.800 ;
        RECT 356.400 16.300 357.200 16.400 ;
        RECT 354.800 15.800 357.200 16.300 ;
        RECT 354.900 15.700 357.200 15.800 ;
        RECT 345.200 14.000 346.400 14.600 ;
        RECT 341.400 12.600 345.200 13.400 ;
        RECT 316.200 12.000 317.000 12.200 ;
        RECT 318.000 12.000 318.800 12.400 ;
        RECT 321.200 12.000 322.000 12.400 ;
        RECT 338.800 12.000 339.600 12.600 ;
        RECT 345.800 12.000 346.400 14.000 ;
        RECT 316.200 11.400 339.600 12.000 ;
        RECT 345.600 11.400 346.400 12.000 ;
        RECT 345.600 9.600 346.200 11.400 ;
        RECT 347.000 10.800 347.800 15.200 ;
        RECT 351.800 15.000 354.200 15.600 ;
        RECT 348.400 14.300 349.200 14.400 ;
        RECT 351.600 14.300 352.600 14.400 ;
        RECT 348.400 13.700 352.600 14.300 ;
        RECT 348.400 13.600 349.200 13.700 ;
        RECT 351.600 13.600 352.600 13.700 ;
        RECT 352.000 12.800 352.800 13.600 ;
        RECT 353.600 12.000 354.200 15.000 ;
        RECT 355.000 12.400 355.600 15.700 ;
        RECT 356.400 15.600 357.200 15.700 ;
        RECT 358.000 14.400 358.600 17.800 ;
        RECT 359.600 16.300 360.400 17.200 ;
        RECT 361.200 16.300 362.000 19.800 ;
        RECT 359.600 15.700 362.000 16.300 ;
        RECT 359.600 15.600 360.400 15.700 ;
        RECT 358.000 14.300 358.800 14.400 ;
        RECT 359.600 14.300 360.400 14.400 ;
        RECT 358.000 13.700 360.400 14.300 ;
        RECT 358.000 13.600 358.800 13.700 ;
        RECT 359.600 13.600 360.400 13.700 ;
        RECT 353.400 11.400 354.200 12.000 ;
        RECT 354.800 12.300 355.600 12.400 ;
        RECT 356.400 12.300 357.200 12.400 ;
        RECT 354.800 11.700 357.200 12.300 ;
        RECT 354.800 11.600 355.600 11.700 ;
        RECT 324.400 9.400 325.200 9.600 ;
        RECT 319.800 9.000 325.200 9.400 ;
        RECT 319.000 8.800 325.200 9.000 ;
        RECT 326.200 9.000 334.800 9.600 ;
        RECT 316.400 8.000 318.000 8.800 ;
        RECT 319.000 8.200 320.400 8.800 ;
        RECT 326.200 8.200 326.800 9.000 ;
        RECT 334.000 8.800 334.800 9.000 ;
        RECT 337.200 9.000 346.200 9.600 ;
        RECT 337.200 8.800 338.000 9.000 ;
        RECT 317.400 7.600 318.000 8.000 ;
        RECT 321.000 7.600 326.800 8.200 ;
        RECT 327.400 7.600 330.000 8.400 ;
        RECT 314.800 6.800 316.800 7.400 ;
        RECT 317.400 6.800 321.600 7.600 ;
        RECT 316.200 6.200 316.800 6.800 ;
        RECT 316.200 5.600 317.200 6.200 ;
        RECT 316.400 2.200 317.200 5.600 ;
        RECT 319.600 2.200 320.400 6.800 ;
        RECT 322.800 2.200 323.600 5.000 ;
        RECT 324.400 2.200 325.200 5.000 ;
        RECT 326.000 2.200 326.800 7.000 ;
        RECT 329.200 2.200 330.000 7.000 ;
        RECT 332.400 2.200 333.200 8.400 ;
        RECT 340.400 7.600 343.000 8.400 ;
        RECT 335.600 6.800 339.800 7.600 ;
        RECT 334.000 2.200 334.800 5.000 ;
        RECT 335.600 2.200 336.400 5.000 ;
        RECT 337.200 2.200 338.000 5.000 ;
        RECT 340.400 2.200 341.200 7.600 ;
        RECT 345.600 7.400 346.200 9.000 ;
        RECT 343.600 6.800 346.200 7.400 ;
        RECT 346.800 10.000 347.800 10.800 ;
        RECT 350.000 11.200 354.200 11.400 ;
        RECT 350.000 10.800 354.000 11.200 ;
        RECT 343.600 2.200 344.400 6.800 ;
        RECT 346.800 2.200 347.600 10.000 ;
        RECT 350.000 2.200 350.800 10.800 ;
        RECT 355.000 10.200 355.600 11.600 ;
        RECT 356.400 10.800 357.200 11.700 ;
        RECT 358.000 10.200 358.600 13.600 ;
        RECT 354.200 9.600 355.600 10.200 ;
        RECT 354.200 2.200 355.000 9.600 ;
        RECT 357.000 9.400 358.800 10.200 ;
        RECT 357.000 2.200 357.800 9.400 ;
        RECT 361.200 2.200 362.000 15.700 ;
        RECT 362.800 15.600 363.600 17.200 ;
        RECT 364.400 13.800 365.200 19.800 ;
        RECT 370.800 16.600 371.600 19.800 ;
        RECT 372.400 17.000 373.200 19.800 ;
        RECT 374.000 17.000 374.800 19.800 ;
        RECT 375.600 17.000 376.400 19.800 ;
        RECT 378.800 17.000 379.600 19.800 ;
        RECT 382.000 17.000 382.800 19.800 ;
        RECT 383.600 17.000 384.400 19.800 ;
        RECT 385.200 17.000 386.000 19.800 ;
        RECT 386.800 17.000 387.600 19.800 ;
        RECT 369.000 15.800 371.600 16.600 ;
        RECT 388.400 16.600 389.200 19.800 ;
        RECT 375.000 15.800 379.600 16.400 ;
        RECT 369.000 15.200 369.800 15.800 ;
        RECT 366.800 14.400 369.800 15.200 ;
        RECT 364.400 13.000 373.200 13.800 ;
        RECT 375.000 13.400 375.800 15.800 ;
        RECT 378.800 15.600 379.600 15.800 ;
        RECT 380.400 15.600 382.000 16.400 ;
        RECT 385.000 15.600 386.000 16.400 ;
        RECT 388.400 15.800 390.800 16.600 ;
        RECT 377.200 13.600 378.000 15.200 ;
        RECT 378.800 14.800 379.600 15.000 ;
        RECT 378.800 14.200 383.200 14.800 ;
        RECT 382.400 14.000 383.200 14.200 ;
        RECT 364.400 7.400 365.200 13.000 ;
        RECT 373.800 12.600 375.800 13.400 ;
        RECT 379.600 12.600 382.800 13.400 ;
        RECT 385.200 12.800 386.000 15.600 ;
        RECT 390.000 15.200 390.800 15.800 ;
        RECT 390.000 14.600 391.800 15.200 ;
        RECT 391.000 13.400 391.800 14.600 ;
        RECT 394.800 14.600 395.600 19.800 ;
        RECT 396.400 16.000 397.200 19.800 ;
        RECT 396.400 15.200 397.400 16.000 ;
        RECT 394.800 14.000 396.000 14.600 ;
        RECT 391.000 12.600 394.800 13.400 ;
        RECT 365.800 12.000 366.600 12.200 ;
        RECT 367.600 12.000 368.400 12.400 ;
        RECT 370.800 12.000 371.600 12.400 ;
        RECT 388.400 12.000 389.200 12.600 ;
        RECT 395.400 12.000 396.000 14.000 ;
        RECT 365.800 11.400 389.200 12.000 ;
        RECT 395.200 11.400 396.000 12.000 ;
        RECT 395.200 9.600 395.800 11.400 ;
        RECT 396.600 10.800 397.400 15.200 ;
        RECT 399.600 15.200 400.400 19.800 ;
        RECT 399.600 14.600 401.800 15.200 ;
        RECT 404.400 15.000 405.200 19.800 ;
        RECT 408.800 18.400 409.600 19.800 ;
        RECT 407.600 17.800 409.600 18.400 ;
        RECT 413.200 17.800 414.000 19.800 ;
        RECT 417.400 18.400 418.600 19.800 ;
        RECT 417.200 17.800 418.600 18.400 ;
        RECT 407.600 17.000 408.400 17.800 ;
        RECT 413.200 17.200 413.800 17.800 ;
        RECT 409.200 15.600 410.000 17.200 ;
        RECT 411.000 16.600 413.800 17.200 ;
        RECT 417.200 17.000 418.000 17.800 ;
        RECT 411.000 16.400 411.800 16.600 ;
        RECT 399.600 11.600 400.400 13.200 ;
        RECT 401.200 11.600 401.800 14.600 ;
        RECT 405.200 14.200 406.800 14.400 ;
        RECT 409.400 14.200 410.000 15.600 ;
        RECT 419.000 15.400 419.800 15.600 ;
        RECT 422.000 15.400 422.800 19.800 ;
        RECT 419.000 14.800 422.800 15.400 ;
        RECT 415.000 14.200 415.800 14.400 ;
        RECT 405.200 13.600 416.200 14.200 ;
        RECT 408.200 13.400 409.000 13.600 ;
        RECT 406.600 12.400 407.400 12.600 ;
        RECT 406.600 11.800 411.600 12.400 ;
        RECT 410.800 11.600 411.600 11.800 ;
        RECT 374.000 9.400 374.800 9.600 ;
        RECT 369.400 9.000 374.800 9.400 ;
        RECT 368.600 8.800 374.800 9.000 ;
        RECT 375.800 9.000 384.400 9.600 ;
        RECT 366.000 8.000 367.600 8.800 ;
        RECT 368.600 8.200 370.000 8.800 ;
        RECT 375.800 8.200 376.400 9.000 ;
        RECT 383.600 8.800 384.400 9.000 ;
        RECT 386.800 9.000 395.800 9.600 ;
        RECT 386.800 8.800 387.600 9.000 ;
        RECT 367.000 7.600 367.600 8.000 ;
        RECT 370.600 7.600 376.400 8.200 ;
        RECT 377.000 7.600 379.600 8.400 ;
        RECT 364.400 6.800 366.400 7.400 ;
        RECT 367.000 6.800 371.200 7.600 ;
        RECT 365.800 6.200 366.400 6.800 ;
        RECT 365.800 5.600 366.800 6.200 ;
        RECT 366.000 2.200 366.800 5.600 ;
        RECT 369.200 2.200 370.000 6.800 ;
        RECT 372.400 2.200 373.200 5.000 ;
        RECT 374.000 2.200 374.800 5.000 ;
        RECT 375.600 2.200 376.400 7.000 ;
        RECT 378.800 2.200 379.600 7.000 ;
        RECT 382.000 2.200 382.800 8.400 ;
        RECT 390.000 7.600 392.600 8.400 ;
        RECT 385.200 6.800 389.400 7.600 ;
        RECT 383.600 2.200 384.400 5.000 ;
        RECT 385.200 2.200 386.000 5.000 ;
        RECT 386.800 2.200 387.600 5.000 ;
        RECT 390.000 2.200 390.800 7.600 ;
        RECT 395.200 7.400 395.800 9.000 ;
        RECT 393.200 6.800 395.800 7.400 ;
        RECT 396.400 10.000 397.400 10.800 ;
        RECT 401.200 10.800 402.400 11.600 ;
        RECT 404.400 11.000 410.000 11.200 ;
        RECT 404.400 10.800 410.200 11.000 ;
        RECT 401.200 10.200 401.800 10.800 ;
        RECT 393.200 2.200 394.000 6.800 ;
        RECT 396.400 2.200 397.200 10.000 ;
        RECT 399.600 9.600 401.800 10.200 ;
        RECT 404.400 10.600 414.200 10.800 ;
        RECT 399.600 2.200 400.400 9.600 ;
        RECT 404.400 2.200 405.200 10.600 ;
        RECT 409.400 10.200 414.200 10.600 ;
        RECT 407.600 9.000 413.000 9.600 ;
        RECT 407.600 8.800 408.400 9.000 ;
        RECT 412.200 8.800 413.000 9.000 ;
        RECT 413.600 9.000 414.200 10.200 ;
        RECT 415.600 10.400 416.200 13.600 ;
        RECT 417.200 12.800 418.000 13.000 ;
        RECT 417.200 12.200 421.000 12.800 ;
        RECT 420.200 12.000 421.000 12.200 ;
        RECT 418.600 11.400 419.400 11.600 ;
        RECT 422.000 11.400 422.800 14.800 ;
        RECT 423.600 17.000 424.400 19.000 ;
        RECT 427.800 18.400 428.600 19.000 ;
        RECT 426.800 17.600 428.600 18.400 ;
        RECT 423.600 14.800 424.200 17.000 ;
        RECT 427.800 16.000 428.600 17.600 ;
        RECT 427.800 15.400 429.400 16.000 ;
        RECT 428.600 15.000 429.400 15.400 ;
        RECT 423.600 14.200 427.800 14.800 ;
        RECT 426.800 13.800 427.800 14.200 ;
        RECT 428.800 14.400 429.400 15.000 ;
        RECT 433.200 15.400 434.000 19.800 ;
        RECT 437.400 18.400 438.600 19.800 ;
        RECT 437.400 17.800 438.800 18.400 ;
        RECT 442.000 17.800 442.800 19.800 ;
        RECT 446.400 18.400 447.200 19.800 ;
        RECT 446.400 17.800 448.400 18.400 ;
        RECT 438.000 17.000 438.800 17.800 ;
        RECT 442.200 17.200 442.800 17.800 ;
        RECT 442.200 16.600 445.000 17.200 ;
        RECT 444.200 16.400 445.000 16.600 ;
        RECT 446.000 15.600 446.800 17.200 ;
        RECT 447.600 17.000 448.400 17.800 ;
        RECT 436.200 15.400 437.000 15.600 ;
        RECT 433.200 14.800 437.000 15.400 ;
        RECT 423.600 11.600 424.400 13.200 ;
        RECT 425.200 11.600 426.000 13.200 ;
        RECT 426.800 13.000 428.200 13.800 ;
        RECT 428.800 13.600 430.800 14.400 ;
        RECT 418.600 10.800 422.800 11.400 ;
        RECT 426.800 11.000 427.400 13.000 ;
        RECT 415.600 9.800 418.000 10.400 ;
        RECT 415.000 9.000 415.800 9.200 ;
        RECT 413.600 8.400 415.800 9.000 ;
        RECT 417.400 8.800 418.000 9.800 ;
        RECT 417.400 8.000 418.800 8.800 ;
        RECT 411.000 7.400 411.800 7.600 ;
        RECT 413.800 7.400 414.600 7.600 ;
        RECT 407.600 6.200 408.400 7.000 ;
        RECT 411.000 6.800 414.600 7.400 ;
        RECT 413.200 6.200 413.800 6.800 ;
        RECT 417.200 6.200 418.000 7.000 ;
        RECT 407.600 5.600 409.600 6.200 ;
        RECT 408.800 2.200 409.600 5.600 ;
        RECT 413.200 2.200 414.000 6.200 ;
        RECT 417.400 2.200 418.600 6.200 ;
        RECT 422.000 2.200 422.800 10.800 ;
        RECT 423.600 10.400 427.400 11.000 ;
        RECT 423.600 7.000 424.200 10.400 ;
        RECT 428.800 9.800 429.400 13.600 ;
        RECT 430.000 10.800 430.800 12.400 ;
        RECT 433.200 11.400 434.000 14.800 ;
        RECT 440.200 14.200 441.000 14.400 ;
        RECT 446.000 14.200 446.600 15.600 ;
        RECT 450.800 15.000 451.600 19.800 ;
        RECT 452.400 15.800 453.200 19.800 ;
        RECT 454.000 16.000 454.800 19.800 ;
        RECT 457.200 16.000 458.000 19.800 ;
        RECT 454.000 15.800 458.000 16.000 ;
        RECT 463.600 17.000 464.400 19.000 ;
        RECT 452.600 14.400 453.200 15.800 ;
        RECT 454.200 15.400 457.800 15.800 ;
        RECT 463.600 14.800 464.200 17.000 ;
        RECT 467.800 16.400 468.600 19.000 ;
        RECT 466.800 16.000 468.600 16.400 ;
        RECT 477.000 16.400 477.800 19.000 ;
        RECT 481.200 17.000 482.000 19.000 ;
        RECT 477.000 16.000 478.800 16.400 ;
        RECT 466.800 15.600 469.400 16.000 ;
        RECT 467.800 15.400 469.400 15.600 ;
        RECT 468.600 15.000 469.400 15.400 ;
        RECT 456.400 14.400 457.200 14.800 ;
        RECT 449.200 14.200 450.800 14.400 ;
        RECT 439.800 13.600 450.800 14.200 ;
        RECT 452.400 13.600 455.000 14.400 ;
        RECT 456.400 13.800 458.000 14.400 ;
        RECT 463.600 14.200 467.800 14.800 ;
        RECT 457.200 13.600 458.000 13.800 ;
        RECT 466.800 13.800 467.800 14.200 ;
        RECT 468.800 14.400 469.400 15.000 ;
        RECT 476.200 15.600 478.800 16.000 ;
        RECT 476.200 15.400 477.800 15.600 ;
        RECT 476.200 15.000 477.000 15.400 ;
        RECT 476.200 14.400 476.800 15.000 ;
        RECT 481.400 14.800 482.000 17.000 ;
        RECT 482.800 16.000 483.600 19.800 ;
        RECT 486.000 16.000 486.800 19.800 ;
        RECT 482.800 15.800 486.800 16.000 ;
        RECT 487.600 15.800 488.400 19.800 ;
        RECT 489.200 15.800 490.000 19.800 ;
        RECT 490.800 16.000 491.600 19.800 ;
        RECT 494.000 16.000 494.800 19.800 ;
        RECT 490.800 15.800 494.800 16.000 ;
        RECT 483.000 15.400 486.600 15.800 ;
        RECT 438.000 12.800 438.800 13.000 ;
        RECT 435.000 12.200 438.800 12.800 ;
        RECT 435.000 12.000 435.800 12.200 ;
        RECT 436.600 11.400 437.400 11.600 ;
        RECT 433.200 10.800 437.400 11.400 ;
        RECT 427.800 9.200 429.400 9.800 ;
        RECT 423.600 3.000 424.400 7.000 ;
        RECT 427.800 2.200 428.600 9.200 ;
        RECT 433.200 2.200 434.000 10.800 ;
        RECT 439.800 10.400 440.400 13.600 ;
        RECT 447.000 13.400 447.800 13.600 ;
        RECT 446.000 12.400 446.800 12.600 ;
        RECT 448.600 12.400 449.400 12.600 ;
        RECT 444.400 11.800 449.400 12.400 ;
        RECT 444.400 11.600 445.200 11.800 ;
        RECT 446.000 11.000 451.600 11.200 ;
        RECT 445.800 10.800 451.600 11.000 ;
        RECT 438.000 9.800 440.400 10.400 ;
        RECT 441.800 10.600 451.600 10.800 ;
        RECT 441.800 10.200 446.600 10.600 ;
        RECT 438.000 8.800 438.600 9.800 ;
        RECT 437.200 8.000 438.600 8.800 ;
        RECT 440.200 9.000 441.000 9.200 ;
        RECT 441.800 9.000 442.400 10.200 ;
        RECT 440.200 8.400 442.400 9.000 ;
        RECT 443.000 9.000 448.400 9.600 ;
        RECT 443.000 8.800 443.800 9.000 ;
        RECT 447.600 8.800 448.400 9.000 ;
        RECT 441.400 7.400 442.200 7.600 ;
        RECT 444.200 7.400 445.000 7.600 ;
        RECT 438.000 6.200 438.800 7.000 ;
        RECT 441.400 6.800 445.000 7.400 ;
        RECT 442.200 6.200 442.800 6.800 ;
        RECT 447.600 6.200 448.400 7.000 ;
        RECT 437.400 2.200 438.600 6.200 ;
        RECT 442.000 2.200 442.800 6.200 ;
        RECT 446.400 5.600 448.400 6.200 ;
        RECT 446.400 2.200 447.200 5.600 ;
        RECT 450.800 2.200 451.600 10.600 ;
        RECT 452.400 10.200 453.200 10.400 ;
        RECT 454.400 10.200 455.000 13.600 ;
        RECT 455.600 11.600 456.400 13.200 ;
        RECT 463.600 11.600 464.400 13.200 ;
        RECT 465.200 11.600 466.000 13.200 ;
        RECT 466.800 13.000 468.200 13.800 ;
        RECT 468.800 13.600 470.800 14.400 ;
        RECT 474.800 13.600 476.800 14.400 ;
        RECT 477.800 14.200 482.000 14.800 ;
        RECT 483.600 14.400 484.400 14.800 ;
        RECT 487.600 14.400 488.200 15.800 ;
        RECT 489.400 14.400 490.000 15.800 ;
        RECT 491.000 15.400 494.600 15.800 ;
        RECT 495.600 15.000 496.400 19.800 ;
        RECT 500.000 18.400 500.800 19.800 ;
        RECT 498.800 17.800 500.800 18.400 ;
        RECT 504.400 17.800 505.200 19.800 ;
        RECT 508.600 18.400 509.800 19.800 ;
        RECT 508.400 17.800 509.800 18.400 ;
        RECT 498.800 17.000 499.600 17.800 ;
        RECT 504.400 17.200 505.000 17.800 ;
        RECT 500.400 16.400 501.200 17.200 ;
        RECT 502.200 16.600 505.000 17.200 ;
        RECT 508.400 17.000 509.200 17.800 ;
        RECT 502.200 16.400 503.000 16.600 ;
        RECT 493.200 14.400 494.000 14.800 ;
        RECT 477.800 13.800 478.800 14.200 ;
        RECT 466.800 11.000 467.400 13.000 ;
        RECT 463.600 10.400 467.400 11.000 ;
        RECT 452.400 9.600 453.800 10.200 ;
        RECT 454.400 9.600 455.400 10.200 ;
        RECT 453.200 8.400 453.800 9.600 ;
        RECT 453.200 7.600 454.000 8.400 ;
        RECT 454.600 2.200 455.400 9.600 ;
        RECT 463.600 7.000 464.200 10.400 ;
        RECT 468.800 9.800 469.400 13.600 ;
        RECT 470.000 12.300 470.800 12.400 ;
        RECT 473.200 12.300 474.000 12.400 ;
        RECT 470.000 11.700 474.000 12.300 ;
        RECT 470.000 10.800 470.800 11.700 ;
        RECT 473.200 11.600 474.000 11.700 ;
        RECT 474.800 10.800 475.600 12.400 ;
        RECT 467.800 9.200 469.400 9.800 ;
        RECT 476.200 9.800 476.800 13.600 ;
        RECT 477.400 13.000 478.800 13.800 ;
        RECT 482.800 13.800 484.400 14.400 ;
        RECT 482.800 13.600 483.600 13.800 ;
        RECT 485.800 13.600 488.400 14.400 ;
        RECT 489.200 13.600 491.800 14.400 ;
        RECT 493.200 13.800 494.800 14.400 ;
        RECT 494.000 13.600 494.800 13.800 ;
        RECT 496.400 14.200 498.000 14.400 ;
        RECT 500.600 14.200 501.200 16.400 ;
        RECT 510.200 15.400 511.000 15.600 ;
        RECT 513.200 15.400 514.000 19.800 ;
        RECT 518.600 16.000 519.400 19.000 ;
        RECT 522.800 17.000 523.600 19.000 ;
        RECT 510.200 14.800 514.000 15.400 ;
        RECT 502.000 14.200 502.800 14.400 ;
        RECT 506.200 14.200 507.000 14.400 ;
        RECT 496.400 13.600 507.400 14.200 ;
        RECT 478.200 11.000 478.800 13.000 ;
        RECT 479.600 11.600 480.400 13.200 ;
        RECT 481.200 11.600 482.000 13.200 ;
        RECT 484.400 11.600 485.200 13.200 ;
        RECT 478.200 10.400 482.000 11.000 ;
        RECT 476.200 9.200 477.800 9.800 ;
        RECT 463.600 3.000 464.400 7.000 ;
        RECT 467.800 2.200 468.600 9.200 ;
        RECT 477.000 2.200 477.800 9.200 ;
        RECT 481.400 7.000 482.000 10.400 ;
        RECT 485.800 10.200 486.400 13.600 ;
        RECT 491.200 12.300 491.800 13.600 ;
        RECT 499.400 13.400 500.200 13.600 ;
        RECT 487.700 11.700 491.800 12.300 ;
        RECT 487.700 10.400 488.300 11.700 ;
        RECT 487.600 10.200 488.400 10.400 ;
        RECT 481.200 3.000 482.000 7.000 ;
        RECT 485.400 9.600 486.400 10.200 ;
        RECT 487.000 9.600 488.400 10.200 ;
        RECT 489.200 10.200 490.000 10.400 ;
        RECT 491.200 10.200 491.800 11.700 ;
        RECT 492.400 11.600 493.200 13.200 ;
        RECT 497.800 12.400 498.600 12.600 ;
        RECT 500.400 12.400 501.200 12.600 ;
        RECT 497.800 11.800 502.800 12.400 ;
        RECT 502.000 11.600 502.800 11.800 ;
        RECT 495.600 11.000 501.200 11.200 ;
        RECT 495.600 10.800 501.400 11.000 ;
        RECT 495.600 10.600 505.400 10.800 ;
        RECT 489.200 9.600 490.600 10.200 ;
        RECT 491.200 9.600 492.200 10.200 ;
        RECT 485.400 2.200 486.200 9.600 ;
        RECT 487.000 8.400 487.600 9.600 ;
        RECT 486.800 7.600 487.600 8.400 ;
        RECT 490.000 8.400 490.600 9.600 ;
        RECT 490.000 7.600 490.800 8.400 ;
        RECT 491.400 2.200 492.200 9.600 ;
        RECT 495.600 2.200 496.400 10.600 ;
        RECT 500.600 10.200 505.400 10.600 ;
        RECT 498.800 9.000 504.200 9.600 ;
        RECT 498.800 8.800 499.600 9.000 ;
        RECT 503.400 8.800 504.200 9.000 ;
        RECT 504.800 9.000 505.400 10.200 ;
        RECT 506.800 10.400 507.400 13.600 ;
        RECT 508.400 12.800 509.200 13.000 ;
        RECT 508.400 12.200 512.200 12.800 ;
        RECT 511.400 12.000 512.200 12.200 ;
        RECT 509.800 11.400 510.600 11.600 ;
        RECT 513.200 11.400 514.000 14.800 ;
        RECT 517.800 15.400 519.400 16.000 ;
        RECT 517.800 15.000 518.600 15.400 ;
        RECT 517.800 14.400 518.400 15.000 ;
        RECT 523.000 14.800 523.600 17.000 ;
        RECT 524.400 16.000 525.200 19.800 ;
        RECT 527.600 16.000 528.400 19.800 ;
        RECT 524.400 15.800 528.400 16.000 ;
        RECT 529.200 15.800 530.000 19.800 ;
        RECT 530.800 15.800 531.600 19.800 ;
        RECT 532.400 16.000 533.200 19.800 ;
        RECT 535.600 16.000 536.400 19.800 ;
        RECT 538.800 16.400 539.600 19.800 ;
        RECT 532.400 15.800 536.400 16.000 ;
        RECT 538.600 15.800 539.600 16.400 ;
        RECT 524.600 15.400 528.200 15.800 ;
        RECT 516.400 13.600 518.400 14.400 ;
        RECT 519.400 14.200 523.600 14.800 ;
        RECT 525.200 14.400 526.000 14.800 ;
        RECT 529.200 14.400 529.800 15.800 ;
        RECT 531.000 14.400 531.600 15.800 ;
        RECT 532.600 15.400 536.200 15.800 ;
        RECT 534.800 14.400 535.600 14.800 ;
        RECT 538.600 14.400 539.200 15.800 ;
        RECT 542.000 15.200 542.800 19.800 ;
        RECT 540.200 14.600 542.800 15.200 ;
        RECT 543.600 15.400 544.400 19.800 ;
        RECT 547.800 18.400 549.000 19.800 ;
        RECT 547.800 17.800 549.200 18.400 ;
        RECT 552.400 17.800 553.200 19.800 ;
        RECT 556.800 18.400 557.600 19.800 ;
        RECT 556.800 17.800 558.800 18.400 ;
        RECT 548.400 17.000 549.200 17.800 ;
        RECT 552.600 17.200 553.200 17.800 ;
        RECT 552.600 16.600 555.400 17.200 ;
        RECT 554.600 16.400 555.400 16.600 ;
        RECT 556.400 16.400 557.200 17.200 ;
        RECT 558.000 17.000 558.800 17.800 ;
        RECT 546.600 15.400 547.400 15.600 ;
        RECT 543.600 14.800 547.400 15.400 ;
        RECT 519.400 13.800 520.400 14.200 ;
        RECT 514.800 12.300 515.600 12.400 ;
        RECT 516.400 12.300 517.200 12.400 ;
        RECT 514.800 11.700 517.200 12.300 ;
        RECT 514.800 11.600 515.600 11.700 ;
        RECT 509.800 10.800 514.000 11.400 ;
        RECT 516.400 10.800 517.200 11.700 ;
        RECT 506.800 9.800 509.200 10.400 ;
        RECT 506.200 9.000 507.000 9.200 ;
        RECT 504.800 8.400 507.000 9.000 ;
        RECT 508.600 8.800 509.200 9.800 ;
        RECT 508.600 8.000 510.000 8.800 ;
        RECT 502.200 7.400 503.000 7.600 ;
        RECT 505.000 7.400 505.800 7.600 ;
        RECT 498.800 6.200 499.600 7.000 ;
        RECT 502.200 6.800 505.800 7.400 ;
        RECT 504.400 6.200 505.000 6.800 ;
        RECT 508.400 6.200 509.200 7.000 ;
        RECT 498.800 5.600 500.800 6.200 ;
        RECT 500.000 2.200 500.800 5.600 ;
        RECT 504.400 2.200 505.200 6.200 ;
        RECT 508.600 2.200 509.800 6.200 ;
        RECT 513.200 2.200 514.000 10.800 ;
        RECT 517.800 10.400 518.400 13.600 ;
        RECT 519.000 13.000 520.400 13.800 ;
        RECT 524.400 13.800 526.000 14.400 ;
        RECT 524.400 13.600 525.200 13.800 ;
        RECT 527.400 13.600 530.000 14.400 ;
        RECT 530.800 13.600 533.400 14.400 ;
        RECT 534.800 14.300 536.400 14.400 ;
        RECT 538.600 14.300 539.600 14.400 ;
        RECT 534.800 13.800 539.600 14.300 ;
        RECT 535.600 13.700 539.600 13.800 ;
        RECT 535.600 13.600 536.400 13.700 ;
        RECT 538.600 13.600 539.600 13.700 ;
        RECT 519.800 11.000 520.400 13.000 ;
        RECT 521.200 11.600 522.000 13.200 ;
        RECT 522.800 11.600 523.600 13.200 ;
        RECT 526.000 11.600 526.800 13.200 ;
        RECT 519.800 10.400 523.600 11.000 ;
        RECT 517.800 9.800 518.800 10.400 ;
        RECT 517.800 9.200 519.400 9.800 ;
        RECT 518.600 2.200 519.400 9.200 ;
        RECT 523.000 7.000 523.600 10.400 ;
        RECT 527.400 10.200 528.000 13.600 ;
        RECT 532.800 12.300 533.400 13.600 ;
        RECT 529.300 11.700 533.400 12.300 ;
        RECT 529.300 10.400 529.900 11.700 ;
        RECT 529.200 10.200 530.000 10.400 ;
        RECT 522.800 3.000 523.600 7.000 ;
        RECT 527.000 9.600 528.000 10.200 ;
        RECT 528.600 9.600 530.000 10.200 ;
        RECT 530.800 10.200 531.600 10.400 ;
        RECT 532.800 10.200 533.400 11.700 ;
        RECT 534.000 11.600 534.800 13.200 ;
        RECT 538.600 10.200 539.200 13.600 ;
        RECT 540.200 13.000 540.800 14.600 ;
        RECT 539.800 12.200 540.800 13.000 ;
        RECT 540.200 10.200 540.800 12.200 ;
        RECT 541.800 12.400 542.600 13.200 ;
        RECT 541.800 11.600 542.800 12.400 ;
        RECT 543.600 11.400 544.400 14.800 ;
        RECT 550.600 14.200 551.400 14.400 ;
        RECT 556.400 14.200 557.000 16.400 ;
        RECT 561.200 15.000 562.000 19.800 ;
        RECT 559.600 14.200 561.200 14.400 ;
        RECT 550.200 13.600 561.200 14.200 ;
        RECT 548.400 12.800 549.200 13.000 ;
        RECT 545.400 12.200 549.200 12.800 ;
        RECT 545.400 12.000 546.200 12.200 ;
        RECT 547.000 11.400 547.800 11.600 ;
        RECT 543.600 10.800 547.800 11.400 ;
        RECT 530.800 9.600 532.200 10.200 ;
        RECT 532.800 9.600 533.800 10.200 ;
        RECT 527.000 2.200 527.800 9.600 ;
        RECT 528.600 8.400 529.200 9.600 ;
        RECT 528.400 7.600 529.200 8.400 ;
        RECT 531.600 8.400 532.200 9.600 ;
        RECT 531.600 7.600 532.400 8.400 ;
        RECT 533.000 2.200 533.800 9.600 ;
        RECT 538.600 9.200 539.600 10.200 ;
        RECT 540.200 9.600 542.800 10.200 ;
        RECT 538.800 2.200 539.600 9.200 ;
        RECT 542.000 2.200 542.800 9.600 ;
        RECT 543.600 2.200 544.400 10.800 ;
        RECT 550.200 10.400 550.800 13.600 ;
        RECT 557.400 13.400 558.200 13.600 ;
        RECT 559.000 12.400 559.800 12.600 ;
        RECT 554.800 11.800 559.800 12.400 ;
        RECT 554.800 11.600 555.600 11.800 ;
        RECT 556.400 11.000 562.000 11.200 ;
        RECT 556.200 10.800 562.000 11.000 ;
        RECT 548.400 9.800 550.800 10.400 ;
        RECT 552.200 10.600 562.000 10.800 ;
        RECT 552.200 10.200 557.000 10.600 ;
        RECT 548.400 8.800 549.000 9.800 ;
        RECT 547.600 8.000 549.000 8.800 ;
        RECT 550.600 9.000 551.400 9.200 ;
        RECT 552.200 9.000 552.800 10.200 ;
        RECT 550.600 8.400 552.800 9.000 ;
        RECT 553.400 9.000 558.800 9.600 ;
        RECT 553.400 8.800 554.200 9.000 ;
        RECT 558.000 8.800 558.800 9.000 ;
        RECT 551.800 7.400 552.600 7.600 ;
        RECT 554.600 7.400 555.400 7.600 ;
        RECT 548.400 6.200 549.200 7.000 ;
        RECT 551.800 6.800 555.400 7.400 ;
        RECT 552.600 6.200 553.200 6.800 ;
        RECT 558.000 6.200 558.800 7.000 ;
        RECT 547.800 2.200 549.000 6.200 ;
        RECT 552.400 2.200 553.200 6.200 ;
        RECT 556.800 5.600 558.800 6.200 ;
        RECT 556.800 2.200 557.600 5.600 ;
        RECT 561.200 2.200 562.000 10.600 ;
        RECT 562.800 2.200 563.600 19.800 ;
        RECT 566.000 16.000 566.800 19.800 ;
        RECT 569.200 16.000 570.000 19.800 ;
        RECT 566.000 15.800 570.000 16.000 ;
        RECT 570.800 15.800 571.600 19.800 ;
        RECT 574.000 16.000 574.800 19.800 ;
        RECT 566.200 15.400 569.800 15.800 ;
        RECT 566.800 14.400 567.600 14.800 ;
        RECT 570.800 14.400 571.400 15.800 ;
        RECT 573.800 15.200 574.800 16.000 ;
        RECT 566.000 13.800 567.600 14.400 ;
        RECT 566.000 13.600 566.800 13.800 ;
        RECT 569.000 13.600 571.600 14.400 ;
        RECT 567.600 11.600 568.400 13.200 ;
        RECT 569.000 10.200 569.600 13.600 ;
        RECT 573.800 10.800 574.600 15.200 ;
        RECT 575.600 14.600 576.400 19.800 ;
        RECT 582.000 16.600 582.800 19.800 ;
        RECT 583.600 17.000 584.400 19.800 ;
        RECT 585.200 17.000 586.000 19.800 ;
        RECT 586.800 17.000 587.600 19.800 ;
        RECT 588.400 17.000 589.200 19.800 ;
        RECT 591.600 17.000 592.400 19.800 ;
        RECT 594.800 17.000 595.600 19.800 ;
        RECT 596.400 17.000 597.200 19.800 ;
        RECT 598.000 17.000 598.800 19.800 ;
        RECT 580.400 15.800 582.800 16.600 ;
        RECT 599.600 16.600 600.400 19.800 ;
        RECT 580.400 15.200 581.200 15.800 ;
        RECT 575.200 14.000 576.400 14.600 ;
        RECT 579.400 14.600 581.200 15.200 ;
        RECT 585.200 15.600 586.200 16.400 ;
        RECT 589.200 15.600 590.800 16.400 ;
        RECT 591.600 15.800 596.200 16.400 ;
        RECT 599.600 15.800 602.200 16.600 ;
        RECT 591.600 15.600 592.400 15.800 ;
        RECT 575.200 12.000 575.800 14.000 ;
        RECT 579.400 13.400 580.200 14.600 ;
        RECT 576.400 12.600 580.200 13.400 ;
        RECT 585.200 12.800 586.000 15.600 ;
        RECT 591.600 14.800 592.400 15.000 ;
        RECT 588.000 14.200 592.400 14.800 ;
        RECT 588.000 14.000 588.800 14.200 ;
        RECT 593.200 13.600 594.000 15.200 ;
        RECT 595.400 13.400 596.200 15.800 ;
        RECT 601.400 15.200 602.200 15.800 ;
        RECT 601.400 14.400 604.400 15.200 ;
        RECT 606.000 13.800 606.800 19.800 ;
        RECT 588.400 12.600 591.600 13.400 ;
        RECT 595.400 12.600 597.400 13.400 ;
        RECT 598.000 13.000 606.800 13.800 ;
        RECT 582.000 12.000 582.800 12.600 ;
        RECT 599.600 12.000 600.400 12.400 ;
        RECT 601.200 12.000 602.000 12.400 ;
        RECT 604.600 12.000 605.400 12.200 ;
        RECT 575.200 11.400 576.000 12.000 ;
        RECT 582.000 11.400 605.400 12.000 ;
        RECT 570.800 10.200 571.600 10.400 ;
        RECT 568.600 9.600 569.600 10.200 ;
        RECT 570.200 9.600 571.600 10.200 ;
        RECT 573.800 10.000 574.800 10.800 ;
        RECT 568.600 2.200 569.400 9.600 ;
        RECT 570.200 8.400 570.800 9.600 ;
        RECT 570.000 7.600 570.800 8.400 ;
        RECT 574.000 2.200 574.800 10.000 ;
        RECT 575.400 9.600 576.000 11.400 ;
        RECT 575.400 9.000 584.400 9.600 ;
        RECT 575.400 7.400 576.000 9.000 ;
        RECT 583.600 8.800 584.400 9.000 ;
        RECT 586.800 9.000 595.400 9.600 ;
        RECT 586.800 8.800 587.600 9.000 ;
        RECT 578.600 7.600 581.200 8.400 ;
        RECT 575.400 6.800 578.000 7.400 ;
        RECT 577.200 2.200 578.000 6.800 ;
        RECT 580.400 2.200 581.200 7.600 ;
        RECT 581.800 6.800 586.000 7.600 ;
        RECT 583.600 2.200 584.400 5.000 ;
        RECT 585.200 2.200 586.000 5.000 ;
        RECT 586.800 2.200 587.600 5.000 ;
        RECT 588.400 2.200 589.200 8.400 ;
        RECT 591.600 7.600 594.200 8.400 ;
        RECT 594.800 8.200 595.400 9.000 ;
        RECT 596.400 9.400 597.200 9.600 ;
        RECT 596.400 9.000 601.800 9.400 ;
        RECT 596.400 8.800 602.600 9.000 ;
        RECT 601.200 8.200 602.600 8.800 ;
        RECT 594.800 7.600 600.600 8.200 ;
        RECT 603.600 8.000 605.200 8.800 ;
        RECT 603.600 7.600 604.200 8.000 ;
        RECT 591.600 2.200 592.400 7.000 ;
        RECT 594.800 2.200 595.600 7.000 ;
        RECT 600.000 6.800 604.200 7.600 ;
        RECT 606.000 7.400 606.800 13.000 ;
        RECT 604.800 6.800 606.800 7.400 ;
        RECT 596.400 2.200 597.200 5.000 ;
        RECT 598.000 2.200 598.800 5.000 ;
        RECT 601.200 2.200 602.000 6.800 ;
        RECT 604.800 6.200 605.400 6.800 ;
        RECT 604.400 5.600 605.400 6.200 ;
        RECT 604.400 2.200 605.200 5.600 ;
        RECT 607.600 2.200 608.400 19.800 ;
      LAYER via1 ;
        RECT 22.000 555.000 22.800 555.800 ;
        RECT 18.800 553.600 19.600 554.400 ;
        RECT 23.600 552.400 24.400 553.200 ;
        RECT 28.400 549.600 29.200 550.400 ;
        RECT 12.400 548.200 13.200 549.000 ;
        RECT 22.000 548.600 22.800 549.400 ;
        RECT 2.800 545.600 3.600 546.400 ;
        RECT 17.200 547.600 18.000 548.400 ;
        RECT 12.400 544.200 13.200 545.000 ;
        RECT 14.000 544.200 14.800 545.000 ;
        RECT 15.600 544.200 16.400 545.000 ;
        RECT 18.800 544.200 19.600 545.000 ;
        RECT 22.000 544.200 22.800 545.000 ;
        RECT 23.600 544.200 24.400 545.000 ;
        RECT 25.200 544.200 26.000 545.000 ;
        RECT 26.800 544.200 27.600 545.000 ;
        RECT 44.400 547.600 45.200 548.400 ;
        RECT 47.600 553.600 48.400 554.400 ;
        RECT 60.400 549.600 61.200 550.400 ;
        RECT 78.000 554.400 78.800 555.200 ;
        RECT 81.200 555.000 82.000 555.800 ;
        RECT 76.400 552.400 77.200 553.200 ;
        RECT 57.200 547.600 58.000 548.400 ;
        RECT 74.800 549.600 75.600 550.400 ;
        RECT 86.000 547.600 86.800 548.400 ;
        RECT 82.800 545.600 83.600 546.400 ;
        RECT 76.400 544.200 77.200 545.000 ;
        RECT 78.000 544.200 78.800 545.000 ;
        RECT 79.600 544.200 80.400 545.000 ;
        RECT 81.200 544.200 82.000 545.000 ;
        RECT 84.400 544.200 85.200 545.000 ;
        RECT 87.600 544.200 88.400 545.000 ;
        RECT 89.200 544.200 90.000 545.000 ;
        RECT 90.800 544.200 91.600 545.000 ;
        RECT 102.000 547.600 102.800 548.400 ;
        RECT 100.400 546.200 101.200 547.000 ;
        RECT 111.600 547.600 112.400 548.400 ;
        RECT 121.200 547.600 122.000 548.400 ;
        RECT 118.000 543.600 118.800 544.400 ;
        RECT 119.600 546.200 120.400 547.000 ;
        RECT 137.200 543.600 138.000 544.400 ;
        RECT 161.200 555.000 162.000 555.800 ;
        RECT 158.000 553.600 158.800 554.400 ;
        RECT 162.800 552.400 163.600 553.200 ;
        RECT 167.600 549.600 168.400 550.400 ;
        RECT 151.600 548.200 152.400 549.000 ;
        RECT 161.200 548.600 162.000 549.400 ;
        RECT 156.400 547.600 157.200 548.400 ;
        RECT 175.800 547.600 176.600 548.400 ;
        RECT 151.600 544.200 152.400 545.000 ;
        RECT 153.200 544.200 154.000 545.000 ;
        RECT 154.800 544.200 155.600 545.000 ;
        RECT 158.000 544.200 158.800 545.000 ;
        RECT 161.200 544.200 162.000 545.000 ;
        RECT 162.800 544.200 163.600 545.000 ;
        RECT 164.400 544.200 165.200 545.000 ;
        RECT 166.000 544.200 166.800 545.000 ;
        RECT 190.000 553.600 190.800 554.400 ;
        RECT 183.600 545.600 184.400 546.400 ;
        RECT 190.000 549.600 190.800 550.400 ;
        RECT 193.200 547.600 194.000 548.400 ;
        RECT 201.200 549.600 202.000 550.400 ;
        RECT 220.400 555.000 221.200 555.800 ;
        RECT 217.200 553.600 218.000 554.400 ;
        RECT 222.000 552.400 222.800 553.200 ;
        RECT 226.800 549.600 227.600 550.400 ;
        RECT 210.800 548.200 211.600 549.000 ;
        RECT 220.400 548.600 221.200 549.400 ;
        RECT 215.600 547.600 216.400 548.400 ;
        RECT 210.800 544.200 211.600 545.000 ;
        RECT 212.400 544.200 213.200 545.000 ;
        RECT 214.000 544.200 214.800 545.000 ;
        RECT 217.200 544.200 218.000 545.000 ;
        RECT 220.400 544.200 221.200 545.000 ;
        RECT 222.000 544.200 222.800 545.000 ;
        RECT 223.600 544.200 224.400 545.000 ;
        RECT 225.200 544.200 226.000 545.000 ;
        RECT 238.000 545.600 238.800 546.400 ;
        RECT 244.400 549.600 245.200 550.400 ;
        RECT 247.600 547.600 248.400 548.400 ;
        RECT 255.600 549.600 256.400 550.400 ;
        RECT 274.800 555.000 275.600 555.800 ;
        RECT 271.600 553.600 272.400 554.400 ;
        RECT 276.400 552.400 277.200 553.200 ;
        RECT 265.200 548.200 266.000 549.000 ;
        RECT 274.800 548.600 275.600 549.400 ;
        RECT 270.000 547.600 270.800 548.400 ;
        RECT 314.800 554.400 315.600 555.200 ;
        RECT 318.000 555.000 318.800 555.800 ;
        RECT 313.200 552.400 314.000 553.200 ;
        RECT 265.200 544.200 266.000 545.000 ;
        RECT 266.800 544.200 267.600 545.000 ;
        RECT 268.400 544.200 269.200 545.000 ;
        RECT 271.600 544.200 272.400 545.000 ;
        RECT 274.800 544.200 275.600 545.000 ;
        RECT 276.400 544.200 277.200 545.000 ;
        RECT 278.000 544.200 278.800 545.000 ;
        RECT 279.600 544.200 280.400 545.000 ;
        RECT 289.200 543.600 290.000 544.400 ;
        RECT 322.800 547.600 323.600 548.400 ;
        RECT 319.600 545.600 320.400 546.400 ;
        RECT 313.200 544.200 314.000 545.000 ;
        RECT 314.800 544.200 315.600 545.000 ;
        RECT 316.400 544.200 317.200 545.000 ;
        RECT 318.000 544.200 318.800 545.000 ;
        RECT 321.200 544.200 322.000 545.000 ;
        RECT 324.400 544.200 325.200 545.000 ;
        RECT 326.000 544.200 326.800 545.000 ;
        RECT 327.600 544.200 328.400 545.000 ;
        RECT 342.000 549.600 342.800 550.400 ;
        RECT 350.000 549.600 350.800 550.400 ;
        RECT 343.600 547.600 344.400 548.400 ;
        RECT 351.600 547.600 352.400 548.400 ;
        RECT 358.000 549.600 358.800 550.400 ;
        RECT 364.400 549.600 365.200 550.400 ;
        RECT 382.000 554.400 382.800 555.200 ;
        RECT 385.200 555.000 386.000 555.800 ;
        RECT 380.400 552.400 381.200 553.200 ;
        RECT 370.800 543.600 371.600 544.400 ;
        RECT 406.000 553.600 406.800 554.400 ;
        RECT 390.000 547.600 390.800 548.400 ;
        RECT 386.800 545.600 387.600 546.400 ;
        RECT 380.400 544.200 381.200 545.000 ;
        RECT 382.000 544.200 382.800 545.000 ;
        RECT 383.600 544.200 384.400 545.000 ;
        RECT 385.200 544.200 386.000 545.000 ;
        RECT 388.400 544.200 389.200 545.000 ;
        RECT 391.600 544.200 392.400 545.000 ;
        RECT 393.200 544.200 394.000 545.000 ;
        RECT 394.800 544.200 395.600 545.000 ;
        RECT 433.200 552.400 434.000 553.200 ;
        RECT 436.400 551.000 437.200 551.800 ;
        RECT 439.600 549.600 440.400 550.400 ;
        RECT 441.200 549.600 442.000 550.400 ;
        RECT 447.600 549.600 448.400 550.400 ;
        RECT 436.400 546.200 437.200 547.000 ;
        RECT 449.200 547.600 450.000 548.400 ;
        RECT 476.400 552.400 477.200 553.200 ;
        RECT 479.600 551.000 480.400 551.800 ;
        RECT 482.800 549.600 483.600 550.400 ;
        RECT 494.000 553.600 494.800 554.400 ;
        RECT 490.800 549.600 491.600 550.400 ;
        RECT 418.800 543.600 419.600 544.400 ;
        RECT 450.800 543.600 451.600 544.400 ;
        RECT 455.600 545.600 456.400 546.400 ;
        RECT 486.000 547.600 486.800 548.400 ;
        RECT 479.600 546.200 480.400 547.000 ;
        RECT 492.400 547.600 493.200 548.400 ;
        RECT 508.400 552.400 509.200 553.200 ;
        RECT 511.600 551.000 512.400 551.800 ;
        RECT 514.800 549.600 515.600 550.400 ;
        RECT 519.600 549.600 520.400 550.400 ;
        RECT 521.200 549.600 522.000 550.400 ;
        RECT 518.000 547.600 518.800 548.400 ;
        RECT 532.400 551.600 533.200 552.400 ;
        RECT 532.400 549.600 533.200 550.400 ;
        RECT 511.600 546.200 512.400 547.000 ;
        RECT 534.000 547.600 534.800 548.400 ;
        RECT 537.200 543.600 538.000 544.400 ;
        RECT 553.200 552.400 554.000 553.200 ;
        RECT 556.400 551.000 557.200 551.800 ;
        RECT 570.800 554.400 571.600 555.200 ;
        RECT 574.000 555.000 574.800 555.800 ;
        RECT 569.200 552.400 570.000 553.200 ;
        RECT 556.400 546.200 557.200 547.000 ;
        RECT 538.800 543.600 539.600 544.400 ;
        RECT 559.600 543.600 560.400 544.400 ;
        RECT 578.800 547.600 579.600 548.400 ;
        RECT 575.600 545.600 576.400 546.400 ;
        RECT 569.200 544.200 570.000 545.000 ;
        RECT 570.800 544.200 571.600 545.000 ;
        RECT 572.400 544.200 573.200 545.000 ;
        RECT 574.000 544.200 574.800 545.000 ;
        RECT 577.200 544.200 578.000 545.000 ;
        RECT 580.400 544.200 581.200 545.000 ;
        RECT 582.000 544.200 582.800 545.000 ;
        RECT 583.600 544.200 584.400 545.000 ;
        RECT 607.600 555.600 608.400 556.400 ;
        RECT 593.200 547.600 594.000 548.400 ;
        RECT 594.800 545.600 595.600 546.400 ;
        RECT 9.200 533.000 10.000 533.800 ;
        RECT 18.800 532.600 19.600 533.400 ;
        RECT 33.200 537.600 34.000 538.400 ;
        RECT 6.000 531.600 6.800 532.400 ;
        RECT 10.800 528.800 11.600 529.600 ;
        RECT 15.600 527.600 16.400 528.400 ;
        RECT 12.400 526.200 13.200 527.000 ;
        RECT 9.200 524.200 10.000 525.000 ;
        RECT 10.800 524.200 11.600 525.000 ;
        RECT 15.600 526.200 16.400 527.000 ;
        RECT 18.800 526.200 19.600 527.000 ;
        RECT 20.400 524.200 21.200 525.000 ;
        RECT 22.000 524.200 22.800 525.000 ;
        RECT 23.600 524.200 24.400 525.000 ;
        RECT 42.800 529.600 43.600 530.400 ;
        RECT 55.600 533.600 56.400 534.400 ;
        RECT 81.200 535.600 82.000 536.400 ;
        RECT 82.800 534.200 83.600 535.000 ;
        RECT 103.600 537.600 104.400 538.400 ;
        RECT 118.000 537.600 118.800 538.400 ;
        RECT 108.400 533.600 109.200 534.400 ;
        RECT 127.600 534.800 128.400 535.600 ;
        RECT 94.000 531.600 94.800 532.400 ;
        RECT 55.600 529.600 56.400 530.400 ;
        RECT 65.200 523.600 66.000 524.400 ;
        RECT 76.400 526.800 77.200 527.600 ;
        RECT 79.600 526.200 80.400 527.000 ;
        RECT 74.800 524.200 75.600 525.000 ;
        RECT 76.400 524.200 77.200 525.000 ;
        RECT 78.000 524.200 78.800 525.000 ;
        RECT 82.800 526.200 83.600 527.000 ;
        RECT 86.000 526.200 86.800 527.000 ;
        RECT 87.600 524.200 88.400 525.000 ;
        RECT 89.200 524.200 90.000 525.000 ;
        RECT 103.600 529.600 104.400 530.400 ;
        RECT 110.000 529.600 110.800 530.400 ;
        RECT 116.400 529.600 117.200 530.400 ;
        RECT 158.000 535.600 158.800 536.400 ;
        RECT 159.600 534.200 160.400 535.000 ;
        RECT 167.600 531.600 168.400 532.400 ;
        RECT 142.000 523.600 142.800 524.400 ;
        RECT 153.200 526.800 154.000 527.600 ;
        RECT 156.400 526.200 157.200 527.000 ;
        RECT 151.600 524.200 152.400 525.000 ;
        RECT 153.200 524.200 154.000 525.000 ;
        RECT 154.800 524.200 155.600 525.000 ;
        RECT 159.600 526.200 160.400 527.000 ;
        RECT 162.800 526.200 163.600 527.000 ;
        RECT 183.600 533.000 184.400 533.800 ;
        RECT 193.200 532.600 194.000 533.400 ;
        RECT 207.600 537.600 208.400 538.400 ;
        RECT 177.200 531.600 178.000 532.400 ;
        RECT 199.600 531.600 200.400 532.400 ;
        RECT 185.200 528.800 186.000 529.600 ;
        RECT 190.000 527.600 190.800 528.400 ;
        RECT 164.400 524.200 165.200 525.000 ;
        RECT 166.000 524.200 166.800 525.000 ;
        RECT 186.800 526.200 187.600 527.000 ;
        RECT 183.600 524.200 184.400 525.000 ;
        RECT 185.200 524.200 186.000 525.000 ;
        RECT 190.000 526.200 190.800 527.000 ;
        RECT 193.200 526.200 194.000 527.000 ;
        RECT 194.800 524.200 195.600 525.000 ;
        RECT 196.400 524.200 197.200 525.000 ;
        RECT 198.000 524.200 198.800 525.000 ;
        RECT 226.800 537.600 227.600 538.400 ;
        RECT 217.200 533.600 218.000 534.400 ;
        RECT 220.400 529.600 221.200 530.400 ;
        RECT 242.800 535.600 243.600 536.400 ;
        RECT 244.400 534.200 245.200 535.000 ;
        RECT 252.400 531.600 253.200 532.400 ;
        RECT 226.800 523.600 227.600 524.400 ;
        RECT 238.000 526.800 238.800 527.600 ;
        RECT 241.200 526.200 242.000 527.000 ;
        RECT 236.400 524.200 237.200 525.000 ;
        RECT 238.000 524.200 238.800 525.000 ;
        RECT 239.600 524.200 240.400 525.000 ;
        RECT 244.400 526.200 245.200 527.000 ;
        RECT 247.600 526.200 248.400 527.000 ;
        RECT 268.400 533.000 269.200 533.800 ;
        RECT 278.000 532.600 278.800 533.400 ;
        RECT 292.400 537.600 293.200 538.400 ;
        RECT 263.600 531.600 264.400 532.400 ;
        RECT 270.000 528.800 270.800 529.600 ;
        RECT 274.800 527.600 275.600 528.400 ;
        RECT 249.200 524.200 250.000 525.000 ;
        RECT 250.800 524.200 251.600 525.000 ;
        RECT 271.600 526.200 272.400 527.000 ;
        RECT 268.400 524.200 269.200 525.000 ;
        RECT 270.000 524.200 270.800 525.000 ;
        RECT 274.800 526.200 275.600 527.000 ;
        RECT 278.000 526.200 278.800 527.000 ;
        RECT 279.600 524.200 280.400 525.000 ;
        RECT 281.200 524.200 282.000 525.000 ;
        RECT 282.800 524.200 283.600 525.000 ;
        RECT 302.000 533.600 302.800 534.400 ;
        RECT 332.400 535.600 333.200 536.400 ;
        RECT 334.000 534.200 334.800 535.000 ;
        RECT 345.200 531.600 346.000 532.400 ;
        RECT 313.200 529.600 314.000 530.400 ;
        RECT 316.400 523.600 317.200 524.400 ;
        RECT 327.600 526.800 328.400 527.600 ;
        RECT 330.800 526.200 331.600 527.000 ;
        RECT 326.000 524.200 326.800 525.000 ;
        RECT 327.600 524.200 328.400 525.000 ;
        RECT 329.200 524.200 330.000 525.000 ;
        RECT 334.000 526.200 334.800 527.000 ;
        RECT 337.200 526.200 338.000 527.000 ;
        RECT 338.800 524.200 339.600 525.000 ;
        RECT 340.400 524.200 341.200 525.000 ;
        RECT 370.800 529.600 371.600 530.400 ;
        RECT 399.600 535.600 400.400 536.400 ;
        RECT 401.200 534.200 402.000 535.000 ;
        RECT 391.600 531.600 392.400 532.400 ;
        RECT 412.400 531.600 413.200 532.400 ;
        RECT 380.400 529.600 381.200 530.400 ;
        RECT 383.600 527.600 384.400 528.400 ;
        RECT 394.800 526.800 395.600 527.600 ;
        RECT 398.000 526.200 398.800 527.000 ;
        RECT 393.200 524.200 394.000 525.000 ;
        RECT 394.800 524.200 395.600 525.000 ;
        RECT 396.400 524.200 397.200 525.000 ;
        RECT 401.200 526.200 402.000 527.000 ;
        RECT 404.400 526.200 405.200 527.000 ;
        RECT 417.200 533.600 418.000 534.400 ;
        RECT 430.000 533.600 430.800 534.400 ;
        RECT 406.000 524.200 406.800 525.000 ;
        RECT 407.600 524.200 408.400 525.000 ;
        RECT 436.400 532.200 437.200 533.000 ;
        RECT 444.400 531.800 445.200 532.600 ;
        RECT 449.200 530.200 450.000 531.000 ;
        RECT 431.600 523.600 432.400 524.400 ;
        RECT 478.000 533.600 478.800 534.400 ;
        RECT 492.400 533.600 493.200 534.400 ;
        RECT 502.000 533.600 502.800 534.400 ;
        RECT 505.200 531.800 506.000 532.600 ;
        RECT 500.400 530.200 501.200 531.000 ;
        RECT 519.600 529.600 520.400 530.400 ;
        RECT 518.000 527.600 518.800 528.400 ;
        RECT 527.600 537.600 528.400 538.400 ;
        RECT 534.000 537.600 534.800 538.400 ;
        RECT 561.200 535.600 562.000 536.400 ;
        RECT 562.800 534.200 563.600 535.000 ;
        RECT 586.800 537.600 587.600 538.400 ;
        RECT 572.400 531.600 573.200 532.400 ;
        RECT 521.200 523.600 522.000 524.400 ;
        RECT 545.200 523.600 546.000 524.400 ;
        RECT 556.400 526.800 557.200 527.600 ;
        RECT 559.600 526.200 560.400 527.000 ;
        RECT 554.800 524.200 555.600 525.000 ;
        RECT 556.400 524.200 557.200 525.000 ;
        RECT 558.000 524.200 558.800 525.000 ;
        RECT 562.800 526.200 563.600 527.000 ;
        RECT 566.000 526.200 566.800 527.000 ;
        RECT 582.000 531.600 582.800 532.400 ;
        RECT 598.000 533.600 598.800 534.400 ;
        RECT 567.600 524.200 568.400 525.000 ;
        RECT 569.200 524.200 570.000 525.000 ;
        RECT 583.600 527.600 584.400 528.400 ;
        RECT 1.200 506.200 2.000 507.000 ;
        RECT 26.800 509.600 27.600 510.400 ;
        RECT 22.000 507.600 22.800 508.400 ;
        RECT 18.800 503.600 19.600 504.400 ;
        RECT 20.400 506.200 21.200 507.000 ;
        RECT 41.200 509.600 42.000 510.400 ;
        RECT 42.800 509.600 43.600 510.400 ;
        RECT 46.000 509.600 46.800 510.400 ;
        RECT 47.600 509.600 48.400 510.400 ;
        RECT 71.600 511.600 72.400 512.400 ;
        RECT 71.600 509.600 72.400 510.400 ;
        RECT 25.200 505.600 26.000 506.400 ;
        RECT 38.000 503.600 38.800 504.400 ;
        RECT 73.200 507.600 74.000 508.400 ;
        RECT 74.800 506.200 75.600 507.000 ;
        RECT 100.400 509.600 101.200 510.400 ;
        RECT 92.400 503.600 93.200 504.400 ;
        RECT 94.000 506.200 94.800 507.000 ;
        RECT 111.600 503.600 112.400 504.400 ;
        RECT 114.800 505.600 115.600 506.400 ;
        RECT 116.400 505.600 117.200 506.400 ;
        RECT 113.200 503.600 114.000 504.400 ;
        RECT 126.000 509.600 126.800 510.400 ;
        RECT 127.600 509.600 128.400 510.400 ;
        RECT 130.800 509.600 131.600 510.400 ;
        RECT 118.000 503.600 118.800 504.400 ;
        RECT 138.800 505.600 139.600 506.400 ;
        RECT 140.400 503.600 141.200 504.400 ;
        RECT 153.200 513.600 154.000 514.400 ;
        RECT 175.600 511.800 176.400 512.600 ;
        RECT 166.000 505.600 166.800 506.400 ;
        RECT 167.600 505.600 168.400 506.400 ;
        RECT 169.200 505.600 170.000 506.400 ;
        RECT 175.600 506.200 176.400 507.000 ;
        RECT 183.600 507.600 184.400 508.400 ;
        RECT 180.400 506.400 181.200 507.200 ;
        RECT 217.200 515.000 218.000 515.800 ;
        RECT 214.000 513.600 214.800 514.400 ;
        RECT 218.800 512.400 219.600 513.200 ;
        RECT 242.800 517.600 243.600 518.400 ;
        RECT 223.600 509.600 224.400 510.400 ;
        RECT 207.600 508.200 208.400 509.000 ;
        RECT 217.200 508.600 218.000 509.400 ;
        RECT 196.400 503.600 197.200 504.400 ;
        RECT 212.400 507.600 213.200 508.400 ;
        RECT 207.600 504.200 208.400 505.000 ;
        RECT 209.200 504.200 210.000 505.000 ;
        RECT 210.800 504.200 211.600 505.000 ;
        RECT 214.000 504.200 214.800 505.000 ;
        RECT 217.200 504.200 218.000 505.000 ;
        RECT 218.800 504.200 219.600 505.000 ;
        RECT 220.400 504.200 221.200 505.000 ;
        RECT 222.000 504.200 222.800 505.000 ;
        RECT 238.000 509.600 238.800 510.400 ;
        RECT 239.600 507.600 240.400 508.400 ;
        RECT 241.200 507.600 242.000 508.400 ;
        RECT 247.600 507.600 248.400 508.400 ;
        RECT 231.600 503.600 232.400 504.400 ;
        RECT 246.000 505.600 246.800 506.400 ;
        RECT 266.800 515.000 267.600 515.800 ;
        RECT 263.600 513.600 264.400 514.400 ;
        RECT 281.200 517.600 282.000 518.400 ;
        RECT 268.400 512.400 269.200 513.200 ;
        RECT 257.200 508.200 258.000 509.000 ;
        RECT 266.800 508.600 267.600 509.400 ;
        RECT 262.000 507.600 262.800 508.400 ;
        RECT 257.200 504.200 258.000 505.000 ;
        RECT 258.800 504.200 259.600 505.000 ;
        RECT 260.400 504.200 261.200 505.000 ;
        RECT 263.600 504.200 264.400 505.000 ;
        RECT 266.800 504.200 267.600 505.000 ;
        RECT 268.400 504.200 269.200 505.000 ;
        RECT 270.000 504.200 270.800 505.000 ;
        RECT 271.600 504.200 272.400 505.000 ;
        RECT 302.000 515.000 302.800 515.800 ;
        RECT 298.800 513.600 299.600 514.400 ;
        RECT 303.600 512.400 304.400 513.200 ;
        RECT 292.400 508.200 293.200 509.000 ;
        RECT 302.000 508.600 302.800 509.400 ;
        RECT 281.200 503.600 282.000 504.400 ;
        RECT 297.200 507.600 298.000 508.400 ;
        RECT 316.600 509.600 317.400 510.400 ;
        RECT 292.400 504.200 293.200 505.000 ;
        RECT 294.000 504.200 294.800 505.000 ;
        RECT 295.600 504.200 296.400 505.000 ;
        RECT 298.800 504.200 299.600 505.000 ;
        RECT 302.000 504.200 302.800 505.000 ;
        RECT 303.600 504.200 304.400 505.000 ;
        RECT 305.200 504.200 306.000 505.000 ;
        RECT 306.800 504.200 307.600 505.000 ;
        RECT 329.200 513.600 330.000 514.400 ;
        RECT 327.600 507.600 328.400 508.400 ;
        RECT 332.400 507.600 333.200 508.400 ;
        RECT 335.600 507.600 336.400 508.400 ;
        RECT 334.000 506.200 334.800 507.000 ;
        RECT 330.800 503.600 331.600 504.400 ;
        RECT 353.200 507.600 354.000 508.400 ;
        RECT 356.400 513.600 357.200 514.400 ;
        RECT 372.400 513.600 373.200 514.400 ;
        RECT 375.600 513.600 376.400 514.400 ;
        RECT 364.400 509.600 365.200 510.400 ;
        RECT 358.000 506.200 358.800 507.000 ;
        RECT 351.600 503.600 352.400 504.400 ;
        RECT 377.200 509.600 378.000 510.400 ;
        RECT 378.800 509.600 379.600 510.400 ;
        RECT 393.200 513.600 394.000 514.400 ;
        RECT 390.000 509.600 390.800 510.400 ;
        RECT 406.000 517.600 406.800 518.400 ;
        RECT 396.400 507.600 397.200 508.400 ;
        RECT 409.200 509.600 410.000 510.400 ;
        RECT 410.800 505.600 411.600 506.400 ;
        RECT 420.400 509.600 421.200 510.400 ;
        RECT 422.000 509.600 422.800 510.400 ;
        RECT 425.200 509.600 426.000 510.400 ;
        RECT 434.800 509.600 435.600 510.400 ;
        RECT 452.400 517.600 453.200 518.400 ;
        RECT 428.400 503.600 429.200 504.400 ;
        RECT 431.600 503.600 432.400 504.400 ;
        RECT 439.600 507.600 440.400 508.400 ;
        RECT 454.000 509.600 454.800 510.400 ;
        RECT 455.600 509.600 456.400 510.400 ;
        RECT 444.400 503.600 445.200 504.400 ;
        RECT 463.600 505.600 464.400 506.400 ;
        RECT 474.800 517.600 475.600 518.400 ;
        RECT 470.000 509.600 470.800 510.400 ;
        RECT 471.600 509.600 472.400 510.400 ;
        RECT 468.400 507.600 469.200 508.400 ;
        RECT 479.600 507.600 480.400 508.400 ;
        RECT 489.200 517.600 490.000 518.400 ;
        RECT 482.800 513.600 483.600 514.400 ;
        RECT 490.800 509.600 491.600 510.400 ;
        RECT 498.800 509.600 499.600 510.400 ;
        RECT 500.400 507.600 501.200 508.400 ;
        RECT 495.600 503.600 496.400 504.400 ;
        RECT 503.600 513.600 504.400 514.400 ;
        RECT 518.000 511.600 518.800 512.400 ;
        RECT 503.600 503.600 504.400 504.400 ;
        RECT 508.400 503.600 509.200 504.400 ;
        RECT 516.400 503.600 517.200 504.400 ;
        RECT 521.200 509.600 522.000 510.400 ;
        RECT 522.800 509.600 523.600 510.400 ;
        RECT 538.800 509.600 539.600 510.400 ;
        RECT 545.200 509.600 546.000 510.400 ;
        RECT 519.600 505.600 520.400 506.400 ;
        RECT 535.600 505.600 536.400 506.400 ;
        RECT 564.400 512.400 565.200 513.200 ;
        RECT 567.600 511.000 568.400 511.800 ;
        RECT 567.600 506.200 568.400 507.000 ;
        RECT 575.600 517.600 576.400 518.400 ;
        RECT 586.800 514.400 587.600 515.200 ;
        RECT 590.000 515.000 590.800 515.800 ;
        RECT 585.200 512.400 586.000 513.200 ;
        RECT 572.400 507.600 573.200 508.400 ;
        RECT 583.600 509.600 584.400 510.400 ;
        RECT 570.800 503.600 571.600 504.400 ;
        RECT 594.800 507.600 595.600 508.400 ;
        RECT 591.600 505.600 592.400 506.400 ;
        RECT 585.200 504.200 586.000 505.000 ;
        RECT 586.800 504.200 587.600 505.000 ;
        RECT 588.400 504.200 589.200 505.000 ;
        RECT 590.000 504.200 590.800 505.000 ;
        RECT 593.200 504.200 594.000 505.000 ;
        RECT 596.400 504.200 597.200 505.000 ;
        RECT 598.000 504.200 598.800 505.000 ;
        RECT 599.600 504.200 600.400 505.000 ;
        RECT 1.200 497.600 2.000 498.400 ;
        RECT 41.200 497.600 42.000 498.400 ;
        RECT 9.200 491.600 10.000 492.400 ;
        RECT 25.200 493.600 26.000 494.400 ;
        RECT 23.600 490.200 24.400 491.000 ;
        RECT 46.000 491.600 46.800 492.400 ;
        RECT 38.000 487.600 38.800 488.400 ;
        RECT 47.600 489.600 48.400 490.400 ;
        RECT 71.600 493.600 72.400 494.400 ;
        RECT 71.600 491.600 72.400 492.400 ;
        RECT 78.000 489.600 78.800 490.400 ;
        RECT 82.800 489.600 83.600 490.400 ;
        RECT 81.200 487.600 82.000 488.400 ;
        RECT 94.000 497.600 94.800 498.400 ;
        RECT 86.000 483.600 86.800 484.400 ;
        RECT 92.400 489.600 93.200 490.400 ;
        RECT 103.600 485.600 104.400 486.400 ;
        RECT 111.600 483.600 112.400 484.400 ;
        RECT 130.800 497.600 131.600 498.400 ;
        RECT 124.400 491.600 125.200 492.400 ;
        RECT 146.800 495.600 147.600 496.400 ;
        RECT 148.400 494.200 149.200 495.000 ;
        RECT 159.600 491.600 160.400 492.400 ;
        RECT 116.400 483.600 117.200 484.400 ;
        RECT 121.200 483.600 122.000 484.400 ;
        RECT 142.000 486.800 142.800 487.600 ;
        RECT 145.200 486.200 146.000 487.000 ;
        RECT 140.400 484.200 141.200 485.000 ;
        RECT 142.000 484.200 142.800 485.000 ;
        RECT 143.600 484.200 144.400 485.000 ;
        RECT 148.400 486.200 149.200 487.000 ;
        RECT 151.600 486.200 152.400 487.000 ;
        RECT 169.200 491.600 170.000 492.400 ;
        RECT 191.600 495.600 192.400 496.400 ;
        RECT 193.200 494.200 194.000 495.000 ;
        RECT 183.600 491.600 184.400 492.400 ;
        RECT 204.400 491.600 205.200 492.400 ;
        RECT 153.200 484.200 154.000 485.000 ;
        RECT 154.800 484.200 155.600 485.000 ;
        RECT 170.800 483.600 171.600 484.400 ;
        RECT 175.600 483.600 176.400 484.400 ;
        RECT 186.800 486.800 187.600 487.600 ;
        RECT 190.000 486.200 190.800 487.000 ;
        RECT 185.200 484.200 186.000 485.000 ;
        RECT 186.800 484.200 187.600 485.000 ;
        RECT 188.400 484.200 189.200 485.000 ;
        RECT 193.200 486.200 194.000 487.000 ;
        RECT 196.400 486.200 197.200 487.000 ;
        RECT 226.800 495.600 227.600 496.400 ;
        RECT 228.400 494.200 229.200 495.000 ;
        RECT 247.600 497.600 248.400 498.400 ;
        RECT 238.000 491.600 238.800 492.400 ;
        RECT 198.000 484.200 198.800 485.000 ;
        RECT 199.600 484.200 200.400 485.000 ;
        RECT 222.000 486.800 222.800 487.600 ;
        RECT 225.200 486.200 226.000 487.000 ;
        RECT 220.400 484.200 221.200 485.000 ;
        RECT 222.000 484.200 222.800 485.000 ;
        RECT 223.600 484.200 224.400 485.000 ;
        RECT 228.400 486.200 229.200 487.000 ;
        RECT 231.600 486.200 232.400 487.000 ;
        RECT 289.200 497.600 290.000 498.400 ;
        RECT 250.800 493.600 251.600 494.400 ;
        RECT 263.600 493.600 264.400 494.400 ;
        RECT 265.200 493.600 266.000 494.400 ;
        RECT 278.000 493.600 278.800 494.400 ;
        RECT 281.200 493.600 282.000 494.400 ;
        RECT 233.200 484.200 234.000 485.000 ;
        RECT 234.800 484.200 235.600 485.000 ;
        RECT 252.400 483.600 253.200 484.400 ;
        RECT 319.600 495.600 320.400 496.400 ;
        RECT 329.200 497.600 330.000 498.400 ;
        RECT 289.200 489.600 290.000 490.400 ;
        RECT 295.600 489.600 296.400 490.400 ;
        RECT 310.000 491.600 310.800 492.400 ;
        RECT 311.600 491.600 312.400 492.400 ;
        RECT 302.000 489.600 302.800 490.400 ;
        RECT 322.800 491.600 323.600 492.400 ;
        RECT 329.200 489.600 330.000 490.400 ;
        RECT 334.000 491.600 334.800 492.400 ;
        RECT 404.400 497.600 405.200 498.400 ;
        RECT 351.600 491.600 352.400 492.400 ;
        RECT 345.200 487.600 346.000 488.400 ;
        RECT 374.000 491.600 374.800 492.400 ;
        RECT 418.800 493.600 419.600 494.400 ;
        RECT 385.200 492.200 386.000 493.000 ;
        RECT 398.000 490.200 398.800 491.000 ;
        RECT 380.400 487.600 381.200 488.400 ;
        RECT 412.400 490.200 413.200 491.000 ;
        RECT 433.200 491.600 434.000 492.400 ;
        RECT 430.000 487.600 430.800 488.400 ;
        RECT 446.000 489.600 446.800 490.400 ;
        RECT 470.000 489.600 470.800 490.400 ;
        RECT 482.800 492.200 483.600 493.000 ;
        RECT 495.600 490.200 496.400 491.000 ;
        RECT 478.000 483.600 478.800 484.400 ;
        RECT 503.600 491.600 504.400 492.400 ;
        RECT 524.400 492.200 525.200 493.000 ;
        RECT 537.200 490.200 538.000 491.000 ;
        RECT 578.800 497.600 579.600 498.400 ;
        RECT 567.600 493.600 568.400 494.400 ;
        RECT 556.400 492.200 557.200 493.000 ;
        RECT 519.600 487.600 520.400 488.400 ;
        RECT 543.600 489.600 544.400 490.400 ;
        RECT 569.200 490.200 570.000 491.000 ;
        RECT 551.600 483.600 552.400 484.400 ;
        RECT 594.800 495.600 595.600 496.400 ;
        RECT 596.400 494.200 597.200 495.000 ;
        RECT 606.000 491.600 606.800 492.400 ;
        RECT 578.800 483.600 579.600 484.400 ;
        RECT 590.000 486.800 590.800 487.600 ;
        RECT 593.200 486.200 594.000 487.000 ;
        RECT 588.400 484.200 589.200 485.000 ;
        RECT 590.000 484.200 590.800 485.000 ;
        RECT 591.600 484.200 592.400 485.000 ;
        RECT 596.400 486.200 597.200 487.000 ;
        RECT 599.600 486.200 600.400 487.000 ;
        RECT 601.200 484.200 602.000 485.000 ;
        RECT 602.800 484.200 603.600 485.000 ;
        RECT 18.800 473.600 19.600 474.400 ;
        RECT 7.600 469.600 8.400 470.400 ;
        RECT 1.200 466.200 2.000 467.000 ;
        RECT 50.800 475.600 51.600 476.400 ;
        RECT 22.000 469.600 22.800 470.400 ;
        RECT 23.600 469.600 24.400 470.400 ;
        RECT 30.000 469.600 30.800 470.400 ;
        RECT 39.600 469.600 40.400 470.400 ;
        RECT 31.600 467.600 32.400 468.400 ;
        RECT 33.200 466.200 34.000 467.000 ;
        RECT 54.000 469.600 54.800 470.400 ;
        RECT 62.000 469.600 62.800 470.400 ;
        RECT 74.800 473.600 75.600 474.400 ;
        RECT 63.600 467.600 64.400 468.400 ;
        RECT 71.600 469.600 72.400 470.400 ;
        RECT 73.200 469.600 74.000 470.400 ;
        RECT 90.800 477.600 91.600 478.400 ;
        RECT 78.000 467.600 78.800 468.400 ;
        RECT 86.000 469.600 86.800 470.400 ;
        RECT 87.600 469.600 88.400 470.400 ;
        RECT 94.000 469.600 94.800 470.400 ;
        RECT 102.000 469.600 102.800 470.400 ;
        RECT 103.600 469.600 104.400 470.400 ;
        RECT 124.400 475.600 125.200 476.400 ;
        RECT 118.000 473.600 118.800 474.400 ;
        RECT 114.800 471.600 115.600 472.400 ;
        RECT 113.200 469.600 114.000 470.400 ;
        RECT 106.800 463.600 107.600 464.400 ;
        RECT 111.600 465.600 112.400 466.400 ;
        RECT 130.800 471.600 131.600 472.400 ;
        RECT 130.800 469.600 131.600 470.400 ;
        RECT 135.600 469.600 136.400 470.400 ;
        RECT 146.800 469.600 147.600 470.400 ;
        RECT 126.000 467.600 126.800 468.400 ;
        RECT 132.400 467.600 133.200 468.400 ;
        RECT 140.400 465.600 141.200 466.400 ;
        RECT 166.000 469.600 166.800 470.400 ;
        RECT 169.200 469.600 170.000 470.400 ;
        RECT 170.800 469.600 171.600 470.400 ;
        RECT 185.200 473.600 186.000 474.400 ;
        RECT 180.400 469.600 181.200 470.400 ;
        RECT 182.000 469.600 182.800 470.400 ;
        RECT 142.000 463.600 142.800 464.400 ;
        RECT 177.200 467.600 178.000 468.400 ;
        RECT 199.600 472.400 200.400 473.200 ;
        RECT 202.800 471.000 203.600 471.800 ;
        RECT 204.400 467.600 205.200 468.400 ;
        RECT 202.800 466.200 203.600 467.000 ;
        RECT 210.800 471.600 211.600 472.400 ;
        RECT 209.200 467.600 210.000 468.400 ;
        RECT 214.000 469.600 214.800 470.400 ;
        RECT 230.000 477.600 230.800 478.400 ;
        RECT 226.800 471.800 227.600 472.600 ;
        RECT 222.000 469.600 222.800 470.400 ;
        RECT 223.600 467.600 224.400 468.400 ;
        RECT 226.800 466.200 227.600 467.000 ;
        RECT 239.600 469.600 240.400 470.400 ;
        RECT 234.800 467.600 235.600 468.400 ;
        RECT 231.600 466.400 232.400 467.200 ;
        RECT 241.200 467.600 242.000 468.400 ;
        RECT 236.400 463.600 237.200 464.400 ;
        RECT 246.000 465.600 246.800 466.400 ;
        RECT 271.600 475.000 272.400 475.800 ;
        RECT 268.400 473.600 269.200 474.400 ;
        RECT 273.200 472.400 274.000 473.200 ;
        RECT 257.200 471.600 258.000 472.400 ;
        RECT 262.000 468.200 262.800 469.000 ;
        RECT 271.600 468.600 272.400 469.400 ;
        RECT 266.800 467.600 267.600 468.400 ;
        RECT 262.000 464.200 262.800 465.000 ;
        RECT 263.600 464.200 264.400 465.000 ;
        RECT 265.200 464.200 266.000 465.000 ;
        RECT 268.400 464.200 269.200 465.000 ;
        RECT 271.600 464.200 272.400 465.000 ;
        RECT 273.200 464.200 274.000 465.000 ;
        RECT 274.800 464.200 275.600 465.000 ;
        RECT 276.400 464.200 277.200 465.000 ;
        RECT 289.200 467.600 290.000 468.400 ;
        RECT 300.400 477.600 301.200 478.400 ;
        RECT 327.600 473.600 328.400 474.400 ;
        RECT 286.000 463.600 286.800 464.400 ;
        RECT 297.200 465.600 298.000 466.400 ;
        RECT 303.600 469.600 304.400 470.400 ;
        RECT 316.400 469.600 317.200 470.400 ;
        RECT 354.800 475.600 355.600 476.400 ;
        RECT 292.400 463.600 293.200 464.400 ;
        RECT 295.600 463.600 296.400 464.400 ;
        RECT 310.000 466.200 310.800 467.000 ;
        RECT 332.400 469.600 333.200 470.400 ;
        RECT 314.800 465.600 315.600 466.400 ;
        RECT 340.400 463.600 341.200 464.400 ;
        RECT 346.800 469.600 347.600 470.400 ;
        RECT 354.800 469.600 355.600 470.400 ;
        RECT 385.200 475.600 386.000 476.400 ;
        RECT 364.400 469.600 365.200 470.400 ;
        RECT 366.000 469.600 366.800 470.400 ;
        RECT 374.000 469.600 374.800 470.400 ;
        RECT 367.600 466.200 368.400 467.000 ;
        RECT 391.600 469.600 392.400 470.400 ;
        RECT 396.400 469.600 397.200 470.400 ;
        RECT 388.400 463.600 389.200 464.400 ;
        RECT 398.000 467.600 398.800 468.400 ;
        RECT 393.200 463.600 394.000 464.400 ;
        RECT 399.600 465.600 400.400 466.400 ;
        RECT 409.200 469.600 410.000 470.400 ;
        RECT 404.400 467.600 405.200 468.400 ;
        RECT 401.200 463.600 402.000 464.400 ;
        RECT 402.800 466.200 403.600 467.000 ;
        RECT 422.000 467.600 422.800 468.400 ;
        RECT 433.200 469.600 434.000 470.400 ;
        RECT 434.800 469.600 435.600 470.400 ;
        RECT 441.200 469.600 442.000 470.400 ;
        RECT 444.400 469.600 445.200 470.400 ;
        RECT 446.000 469.600 446.800 470.400 ;
        RECT 442.800 467.600 443.600 468.400 ;
        RECT 465.200 469.600 466.000 470.400 ;
        RECT 466.800 469.600 467.600 470.400 ;
        RECT 420.400 463.600 421.200 464.400 ;
        RECT 430.000 463.600 430.800 464.400 ;
        RECT 468.400 467.600 469.200 468.400 ;
        RECT 474.800 469.600 475.600 470.400 ;
        RECT 481.200 471.600 482.000 472.400 ;
        RECT 484.400 469.600 485.200 470.400 ;
        RECT 486.000 469.600 486.800 470.400 ;
        RECT 487.600 469.600 488.400 470.400 ;
        RECT 478.000 463.600 478.800 464.400 ;
        RECT 495.600 465.600 496.400 466.400 ;
        RECT 506.800 477.600 507.600 478.400 ;
        RECT 500.400 469.600 501.200 470.400 ;
        RECT 502.000 469.600 502.800 470.400 ;
        RECT 505.200 467.600 506.000 468.400 ;
        RECT 511.600 477.600 512.400 478.400 ;
        RECT 524.400 477.600 525.200 478.400 ;
        RECT 519.600 469.600 520.400 470.400 ;
        RECT 521.200 469.600 522.000 470.400 ;
        RECT 497.200 463.600 498.000 464.400 ;
        RECT 514.800 465.600 515.600 466.400 ;
        RECT 538.800 471.800 539.600 472.600 ;
        RECT 535.600 465.600 536.400 466.400 ;
        RECT 538.800 466.200 539.600 467.000 ;
        RECT 553.200 471.600 554.000 472.400 ;
        RECT 557.800 471.800 558.600 472.600 ;
        RECT 569.000 471.800 569.800 472.600 ;
        RECT 543.600 466.400 544.400 467.200 ;
        RECT 543.600 463.600 544.400 464.400 ;
        RECT 591.600 474.400 592.400 475.200 ;
        RECT 594.800 475.000 595.600 475.800 ;
        RECT 590.000 472.400 590.800 473.200 ;
        RECT 554.800 465.600 555.600 466.400 ;
        RECT 557.800 466.200 558.600 467.000 ;
        RECT 566.000 467.600 566.800 468.400 ;
        RECT 562.800 463.600 563.600 464.400 ;
        RECT 569.000 466.200 569.800 467.000 ;
        RECT 577.200 467.600 578.000 468.400 ;
        RECT 588.400 469.600 589.200 470.400 ;
        RECT 599.600 467.600 600.400 468.400 ;
        RECT 596.400 465.600 597.200 466.400 ;
        RECT 590.000 464.200 590.800 465.000 ;
        RECT 591.600 464.200 592.400 465.000 ;
        RECT 593.200 464.200 594.000 465.000 ;
        RECT 594.800 464.200 595.600 465.000 ;
        RECT 598.000 464.200 598.800 465.000 ;
        RECT 601.200 464.200 602.000 465.000 ;
        RECT 602.800 464.200 603.600 465.000 ;
        RECT 604.400 464.200 605.200 465.000 ;
        RECT 38.000 457.600 38.800 458.400 ;
        RECT 17.200 453.600 18.000 454.400 ;
        RECT 6.000 452.200 6.800 453.000 ;
        RECT 14.000 451.800 14.800 452.600 ;
        RECT 23.600 451.600 24.400 452.400 ;
        RECT 28.400 451.600 29.200 452.400 ;
        RECT 18.800 450.200 19.600 451.000 ;
        RECT 1.200 443.600 2.000 444.400 ;
        RECT 25.200 449.600 26.000 450.400 ;
        RECT 41.200 457.600 42.000 458.400 ;
        RECT 47.600 453.600 48.400 454.400 ;
        RECT 54.000 453.600 54.800 454.400 ;
        RECT 44.400 451.600 45.200 452.400 ;
        RECT 52.400 450.200 53.200 451.000 ;
        RECT 95.600 457.600 96.400 458.400 ;
        RECT 70.000 447.600 70.800 448.400 ;
        RECT 130.800 457.600 131.600 458.400 ;
        RECT 98.800 451.600 99.600 452.400 ;
        RECT 105.200 449.600 106.000 450.400 ;
        RECT 121.200 451.600 122.000 452.400 ;
        RECT 118.000 443.600 118.800 444.400 ;
        RECT 143.600 449.600 144.400 450.400 ;
        RECT 177.200 457.600 178.000 458.400 ;
        RECT 156.400 451.600 157.200 452.400 ;
        RECT 148.400 449.600 149.200 450.400 ;
        RECT 174.000 453.600 174.800 454.400 ;
        RECT 167.600 451.600 168.400 452.400 ;
        RECT 193.200 453.600 194.000 454.400 ;
        RECT 182.000 452.200 182.800 453.000 ;
        RECT 167.600 443.600 168.400 444.400 ;
        RECT 175.600 449.600 176.400 450.400 ;
        RECT 194.800 450.200 195.600 451.000 ;
        RECT 177.200 443.600 178.000 444.400 ;
        RECT 207.600 457.600 208.400 458.400 ;
        RECT 201.200 443.600 202.000 444.400 ;
        RECT 222.000 455.600 222.800 456.400 ;
        RECT 210.800 453.600 211.600 454.400 ;
        RECT 225.200 449.600 226.000 450.400 ;
        RECT 254.000 455.600 254.800 456.400 ;
        RECT 255.600 454.200 256.400 455.000 ;
        RECT 246.000 451.600 246.800 452.400 ;
        RECT 233.200 443.600 234.000 444.400 ;
        RECT 238.000 443.600 238.800 444.400 ;
        RECT 249.200 446.800 250.000 447.600 ;
        RECT 252.400 446.200 253.200 447.000 ;
        RECT 247.600 444.200 248.400 445.000 ;
        RECT 249.200 444.200 250.000 445.000 ;
        RECT 250.800 444.200 251.600 445.000 ;
        RECT 255.600 446.200 256.400 447.000 ;
        RECT 258.800 446.200 259.600 447.000 ;
        RECT 289.200 457.600 290.000 458.400 ;
        RECT 274.800 453.600 275.600 454.400 ;
        RECT 260.400 444.200 261.200 445.000 ;
        RECT 262.000 444.200 262.800 445.000 ;
        RECT 313.200 455.600 314.000 456.400 ;
        RECT 314.800 454.200 315.600 455.000 ;
        RECT 305.200 451.600 306.000 452.400 ;
        RECT 281.200 443.600 282.000 444.400 ;
        RECT 297.200 443.600 298.000 444.400 ;
        RECT 308.400 446.800 309.200 447.600 ;
        RECT 311.600 446.200 312.400 447.000 ;
        RECT 306.800 444.200 307.600 445.000 ;
        RECT 308.400 444.200 309.200 445.000 ;
        RECT 310.000 444.200 310.800 445.000 ;
        RECT 314.800 446.200 315.600 447.000 ;
        RECT 318.000 446.200 318.800 447.000 ;
        RECT 335.600 452.200 336.400 453.000 ;
        RECT 343.600 451.800 344.400 452.600 ;
        RECT 348.400 450.200 349.200 451.000 ;
        RECT 330.800 447.600 331.600 448.400 ;
        RECT 319.600 444.200 320.400 445.000 ;
        RECT 321.200 444.200 322.000 445.000 ;
        RECT 362.800 451.600 363.600 452.400 ;
        RECT 351.600 447.600 352.400 448.400 ;
        RECT 364.400 449.600 365.200 450.400 ;
        RECT 372.400 451.600 373.200 452.400 ;
        RECT 382.000 453.600 382.800 454.400 ;
        RECT 390.000 453.600 390.800 454.400 ;
        RECT 398.000 453.600 398.800 454.400 ;
        RECT 390.000 449.600 390.800 450.400 ;
        RECT 391.600 450.200 392.400 451.000 ;
        RECT 439.600 453.600 440.400 454.400 ;
        RECT 409.200 443.600 410.000 444.400 ;
        RECT 434.800 449.600 435.600 450.400 ;
        RECT 420.400 443.600 421.200 444.400 ;
        RECT 426.800 443.600 427.600 444.400 ;
        RECT 441.200 449.600 442.000 450.400 ;
        RECT 444.400 443.600 445.200 444.400 ;
        RECT 450.800 443.600 451.600 444.400 ;
        RECT 468.400 449.600 469.200 450.400 ;
        RECT 474.800 449.600 475.600 450.400 ;
        RECT 494.000 453.600 494.800 454.400 ;
        RECT 540.400 457.600 541.200 458.400 ;
        RECT 489.200 451.600 490.000 452.400 ;
        RECT 505.200 451.600 506.000 452.400 ;
        RECT 503.600 449.600 504.400 450.400 ;
        RECT 513.200 451.600 514.000 452.400 ;
        RECT 513.200 445.600 514.000 446.400 ;
        RECT 529.200 443.600 530.000 444.400 ;
        RECT 556.400 455.600 557.200 456.400 ;
        RECT 558.000 454.200 558.800 455.000 ;
        RECT 559.600 451.600 560.400 452.400 ;
        RECT 535.600 443.600 536.400 444.400 ;
        RECT 551.600 446.800 552.400 447.600 ;
        RECT 554.800 446.200 555.600 447.000 ;
        RECT 550.000 444.200 550.800 445.000 ;
        RECT 551.600 444.200 552.400 445.000 ;
        RECT 553.200 444.200 554.000 445.000 ;
        RECT 558.000 446.200 558.800 447.000 ;
        RECT 561.200 446.200 562.000 447.000 ;
        RECT 591.600 455.600 592.400 456.400 ;
        RECT 593.200 454.200 594.000 455.000 ;
        RECT 583.600 451.600 584.400 452.400 ;
        RECT 562.800 444.200 563.600 445.000 ;
        RECT 564.400 444.200 565.200 445.000 ;
        RECT 575.600 443.600 576.400 444.400 ;
        RECT 586.800 446.800 587.600 447.600 ;
        RECT 590.000 446.200 590.800 447.000 ;
        RECT 585.200 444.200 586.000 445.000 ;
        RECT 586.800 444.200 587.600 445.000 ;
        RECT 588.400 444.200 589.200 445.000 ;
        RECT 593.200 446.200 594.000 447.000 ;
        RECT 596.400 446.200 597.200 447.000 ;
        RECT 598.000 444.200 598.800 445.000 ;
        RECT 599.600 444.200 600.400 445.000 ;
        RECT 6.000 429.600 6.800 430.400 ;
        RECT 22.000 437.600 22.800 438.400 ;
        RECT 28.400 437.600 29.200 438.400 ;
        RECT 7.600 427.600 8.400 428.400 ;
        RECT 28.400 429.600 29.200 430.400 ;
        RECT 66.800 433.600 67.600 434.400 ;
        RECT 70.000 433.600 70.800 434.400 ;
        RECT 31.600 425.600 32.400 426.400 ;
        RECT 54.000 427.600 54.800 428.400 ;
        RECT 52.400 426.200 53.200 427.000 ;
        RECT 71.600 429.600 72.400 430.400 ;
        RECT 73.200 429.600 74.000 430.400 ;
        RECT 84.400 429.600 85.200 430.400 ;
        RECT 90.800 429.600 91.600 430.400 ;
        RECT 57.200 425.600 58.000 426.400 ;
        RECT 92.400 427.600 93.200 428.400 ;
        RECT 94.000 427.600 94.800 428.400 ;
        RECT 98.800 429.600 99.600 430.400 ;
        RECT 100.400 429.600 101.200 430.400 ;
        RECT 110.000 429.600 110.800 430.400 ;
        RECT 118.000 429.600 118.800 430.400 ;
        RECT 113.200 427.600 114.000 428.400 ;
        RECT 119.600 427.600 120.400 428.400 ;
        RECT 132.400 437.600 133.200 438.400 ;
        RECT 126.000 429.600 126.800 430.400 ;
        RECT 121.200 425.600 122.000 426.400 ;
        RECT 130.800 425.600 131.600 426.400 ;
        RECT 129.200 423.600 130.000 424.400 ;
        RECT 134.000 433.600 134.800 434.400 ;
        RECT 148.400 432.400 149.200 433.200 ;
        RECT 167.600 433.600 168.400 434.400 ;
        RECT 151.600 431.000 152.400 431.800 ;
        RECT 180.400 437.600 181.200 438.400 ;
        RECT 183.600 437.600 184.400 438.400 ;
        RECT 167.600 429.600 168.400 430.400 ;
        RECT 172.400 429.600 173.200 430.400 ;
        RECT 180.400 429.600 181.200 430.400 ;
        RECT 151.600 426.200 152.400 427.000 ;
        RECT 169.200 427.600 170.000 428.400 ;
        RECT 182.000 427.600 182.800 428.400 ;
        RECT 198.000 432.400 198.800 433.200 ;
        RECT 201.200 431.000 202.000 431.800 ;
        RECT 204.400 429.600 205.200 430.400 ;
        RECT 210.800 429.600 211.600 430.400 ;
        RECT 201.200 426.200 202.000 427.000 ;
        RECT 223.600 429.600 224.400 430.400 ;
        RECT 218.800 427.600 219.600 428.400 ;
        RECT 233.200 427.600 234.000 428.400 ;
        RECT 238.000 427.600 238.800 428.400 ;
        RECT 246.000 429.600 246.800 430.400 ;
        RECT 273.200 437.600 274.000 438.400 ;
        RECT 255.600 429.600 256.400 430.400 ;
        RECT 258.800 429.600 259.600 430.400 ;
        RECT 260.400 429.600 261.200 430.400 ;
        RECT 214.000 423.600 214.800 424.400 ;
        RECT 257.200 427.600 258.000 428.400 ;
        RECT 268.400 429.600 269.200 430.400 ;
        RECT 270.000 429.600 270.800 430.400 ;
        RECT 265.200 427.600 266.000 428.400 ;
        RECT 284.400 437.600 285.200 438.400 ;
        RECT 281.200 427.600 282.000 428.400 ;
        RECT 282.800 425.600 283.600 426.400 ;
        RECT 279.600 423.600 280.400 424.400 ;
        RECT 287.600 433.600 288.400 434.400 ;
        RECT 298.800 434.400 299.600 435.200 ;
        RECT 302.000 435.000 302.800 435.800 ;
        RECT 327.600 437.600 328.400 438.400 ;
        RECT 297.200 432.400 298.000 433.200 ;
        RECT 295.600 429.600 296.400 430.400 ;
        RECT 306.800 427.600 307.600 428.400 ;
        RECT 303.600 425.600 304.400 426.400 ;
        RECT 297.200 424.200 298.000 425.000 ;
        RECT 298.800 424.200 299.600 425.000 ;
        RECT 300.400 424.200 301.200 425.000 ;
        RECT 302.000 424.200 302.800 425.000 ;
        RECT 305.200 424.200 306.000 425.000 ;
        RECT 308.400 424.200 309.200 425.000 ;
        RECT 310.000 424.200 310.800 425.000 ;
        RECT 311.600 424.200 312.400 425.000 ;
        RECT 326.000 425.600 326.800 426.400 ;
        RECT 346.800 433.600 347.600 434.400 ;
        RECT 335.600 429.600 336.400 430.400 ;
        RECT 329.200 426.200 330.000 427.000 ;
        RECT 348.400 429.600 349.200 430.400 ;
        RECT 350.000 429.600 350.800 430.400 ;
        RECT 361.200 429.600 362.000 430.400 ;
        RECT 367.600 429.600 368.400 430.400 ;
        RECT 369.200 427.600 370.000 428.400 ;
        RECT 377.200 429.600 378.000 430.400 ;
        RECT 378.800 429.600 379.600 430.400 ;
        RECT 382.000 429.600 382.800 430.400 ;
        RECT 398.000 431.600 398.800 432.400 ;
        RECT 393.200 429.600 394.000 430.400 ;
        RECT 396.400 425.600 397.200 426.400 ;
        RECT 415.600 433.600 416.400 434.400 ;
        RECT 402.800 429.600 403.600 430.400 ;
        RECT 406.000 429.600 406.800 430.400 ;
        RECT 407.600 429.600 408.400 430.400 ;
        RECT 410.800 429.600 411.600 430.400 ;
        RECT 430.000 432.400 430.800 433.200 ;
        RECT 433.200 431.000 434.000 431.800 ;
        RECT 439.600 429.600 440.400 430.400 ;
        RECT 462.000 433.600 462.800 434.400 ;
        RECT 471.600 437.600 472.400 438.400 ;
        RECT 470.000 433.600 470.800 434.400 ;
        RECT 433.200 426.200 434.000 427.000 ;
        RECT 434.800 425.600 435.600 426.400 ;
        RECT 446.000 427.600 446.800 428.400 ;
        RECT 444.400 426.200 445.200 427.000 ;
        RECT 442.800 423.600 443.600 424.400 ;
        RECT 487.600 434.400 488.400 435.200 ;
        RECT 490.800 435.000 491.600 435.800 ;
        RECT 511.600 437.600 512.400 438.400 ;
        RECT 486.000 432.400 486.800 433.200 ;
        RECT 471.600 429.600 472.400 430.400 ;
        RECT 495.600 427.600 496.400 428.400 ;
        RECT 492.400 425.600 493.200 426.400 ;
        RECT 486.000 424.200 486.800 425.000 ;
        RECT 487.600 424.200 488.400 425.000 ;
        RECT 489.200 424.200 490.000 425.000 ;
        RECT 490.800 424.200 491.600 425.000 ;
        RECT 494.000 424.200 494.800 425.000 ;
        RECT 497.200 424.200 498.000 425.000 ;
        RECT 498.800 424.200 499.600 425.000 ;
        RECT 500.400 424.200 501.200 425.000 ;
        RECT 522.800 434.400 523.600 435.200 ;
        RECT 526.000 435.000 526.800 435.800 ;
        RECT 521.200 432.400 522.000 433.200 ;
        RECT 519.600 429.600 520.400 430.400 ;
        RECT 559.600 437.600 560.400 438.400 ;
        RECT 530.800 427.600 531.600 428.400 ;
        RECT 527.600 425.600 528.400 426.400 ;
        RECT 545.200 429.600 546.000 430.400 ;
        RECT 546.800 429.600 547.600 430.400 ;
        RECT 521.200 424.200 522.000 425.000 ;
        RECT 522.800 424.200 523.600 425.000 ;
        RECT 524.400 424.200 525.200 425.000 ;
        RECT 526.000 424.200 526.800 425.000 ;
        RECT 529.200 424.200 530.000 425.000 ;
        RECT 532.400 424.200 533.200 425.000 ;
        RECT 534.000 424.200 534.800 425.000 ;
        RECT 535.600 424.200 536.400 425.000 ;
        RECT 554.800 429.600 555.600 430.400 ;
        RECT 556.400 429.600 557.200 430.400 ;
        RECT 577.200 434.400 578.000 435.200 ;
        RECT 580.400 435.000 581.200 435.800 ;
        RECT 575.600 432.400 576.400 433.200 ;
        RECT 574.000 429.600 574.800 430.400 ;
        RECT 566.000 423.600 566.800 424.400 ;
        RECT 585.200 427.600 586.000 428.400 ;
        RECT 582.000 425.600 582.800 426.400 ;
        RECT 575.600 424.200 576.400 425.000 ;
        RECT 577.200 424.200 578.000 425.000 ;
        RECT 578.800 424.200 579.600 425.000 ;
        RECT 580.400 424.200 581.200 425.000 ;
        RECT 583.600 424.200 584.400 425.000 ;
        RECT 586.800 424.200 587.600 425.000 ;
        RECT 588.400 424.200 589.200 425.000 ;
        RECT 590.000 424.200 590.800 425.000 ;
        RECT 601.200 423.600 602.000 424.400 ;
        RECT 9.200 413.000 10.000 413.800 ;
        RECT 18.800 412.600 19.600 413.400 ;
        RECT 36.400 417.600 37.200 418.400 ;
        RECT 25.200 411.600 26.000 412.400 ;
        RECT 10.800 408.800 11.600 409.600 ;
        RECT 15.600 407.600 16.400 408.400 ;
        RECT 12.400 406.200 13.200 407.000 ;
        RECT 9.200 404.200 10.000 405.000 ;
        RECT 10.800 404.200 11.600 405.000 ;
        RECT 15.600 406.200 16.400 407.000 ;
        RECT 18.800 406.200 19.600 407.000 ;
        RECT 20.400 404.200 21.200 405.000 ;
        RECT 22.000 404.200 22.800 405.000 ;
        RECT 23.600 404.200 24.400 405.000 ;
        RECT 55.600 413.600 56.400 414.400 ;
        RECT 66.800 413.600 67.600 414.400 ;
        RECT 100.400 417.600 101.200 418.400 ;
        RECT 47.600 409.600 48.400 410.400 ;
        RECT 55.600 411.600 56.400 412.400 ;
        RECT 70.000 411.800 70.800 412.600 ;
        RECT 65.200 410.200 66.000 411.000 ;
        RECT 82.800 407.600 83.600 408.400 ;
        RECT 116.400 417.600 117.200 418.400 ;
        RECT 110.000 413.600 110.800 414.400 ;
        RECT 100.400 409.600 101.200 410.400 ;
        RECT 106.800 409.600 107.600 410.400 ;
        RECT 124.400 417.600 125.200 418.400 ;
        RECT 113.200 411.600 114.000 412.400 ;
        RECT 119.600 411.600 120.400 412.400 ;
        RECT 129.200 415.600 130.000 416.400 ;
        RECT 135.600 409.600 136.400 410.400 ;
        RECT 172.400 417.600 173.200 418.400 ;
        RECT 167.600 413.600 168.400 414.400 ;
        RECT 148.400 409.600 149.200 410.400 ;
        RECT 142.000 403.600 142.800 404.400 ;
        RECT 150.000 409.600 150.800 410.400 ;
        RECT 161.200 409.600 162.000 410.400 ;
        RECT 167.600 409.600 168.400 410.400 ;
        RECT 190.000 413.000 190.800 413.800 ;
        RECT 180.400 409.600 181.200 410.400 ;
        RECT 199.600 412.600 200.400 413.400 ;
        RECT 194.800 411.600 195.600 412.400 ;
        RECT 191.600 408.800 192.400 409.600 ;
        RECT 196.400 407.600 197.200 408.400 ;
        RECT 193.200 406.200 194.000 407.000 ;
        RECT 190.000 404.200 190.800 405.000 ;
        RECT 191.600 404.200 192.400 405.000 ;
        RECT 196.400 406.200 197.200 407.000 ;
        RECT 199.600 406.200 200.400 407.000 ;
        RECT 201.200 404.200 202.000 405.000 ;
        RECT 202.800 404.200 203.600 405.000 ;
        RECT 204.400 404.200 205.200 405.000 ;
        RECT 226.800 417.600 227.600 418.400 ;
        RECT 223.600 411.600 224.400 412.400 ;
        RECT 230.000 411.600 230.800 412.400 ;
        RECT 234.800 411.600 235.600 412.400 ;
        RECT 254.000 417.600 254.800 418.400 ;
        RECT 273.200 417.600 274.000 418.400 ;
        RECT 218.800 407.600 219.600 408.400 ;
        RECT 242.800 409.600 243.600 410.400 ;
        RECT 258.800 413.600 259.600 414.400 ;
        RECT 262.000 413.600 262.800 414.400 ;
        RECT 276.400 413.600 277.200 414.400 ;
        RECT 281.200 413.600 282.000 414.400 ;
        RECT 282.800 407.600 283.600 408.400 ;
        RECT 308.400 413.000 309.200 413.800 ;
        RECT 294.000 409.600 294.800 410.400 ;
        RECT 318.000 412.600 318.800 413.400 ;
        RECT 303.600 411.600 304.400 412.400 ;
        RECT 353.200 417.600 354.000 418.400 ;
        RECT 337.200 413.600 338.000 414.400 ;
        RECT 310.000 408.800 310.800 409.600 ;
        RECT 314.800 407.600 315.600 408.400 ;
        RECT 311.600 406.200 312.400 407.000 ;
        RECT 308.400 404.200 309.200 405.000 ;
        RECT 310.000 404.200 310.800 405.000 ;
        RECT 314.800 406.200 315.600 407.000 ;
        RECT 318.000 406.200 318.800 407.000 ;
        RECT 319.600 404.200 320.400 405.000 ;
        RECT 321.200 404.200 322.000 405.000 ;
        RECT 322.800 404.200 323.600 405.000 ;
        RECT 335.600 410.200 336.400 411.000 ;
        RECT 332.400 407.600 333.200 408.400 ;
        RECT 369.200 415.600 370.000 416.400 ;
        RECT 350.000 407.600 350.800 408.400 ;
        RECT 359.600 409.600 360.400 410.400 ;
        RECT 375.600 409.600 376.400 410.400 ;
        RECT 380.400 403.600 381.200 404.400 ;
        RECT 410.800 417.600 411.600 418.400 ;
        RECT 391.600 409.600 392.400 410.400 ;
        RECT 394.800 405.600 395.600 406.400 ;
        RECT 410.800 409.600 411.600 410.400 ;
        RECT 436.400 415.600 437.200 416.400 ;
        RECT 420.400 409.600 421.200 410.400 ;
        RECT 426.800 409.600 427.600 410.400 ;
        RECT 433.200 409.600 434.000 410.400 ;
        RECT 447.600 409.600 448.400 410.400 ;
        RECT 481.200 417.600 482.000 418.400 ;
        RECT 481.200 414.800 482.000 415.600 ;
        RECT 484.400 413.600 485.200 414.400 ;
        RECT 465.200 405.600 466.000 406.400 ;
        RECT 471.600 403.600 472.400 404.400 ;
        RECT 495.600 413.200 496.400 414.000 ;
        RECT 502.000 413.600 502.800 414.400 ;
        RECT 489.200 403.600 490.000 404.400 ;
        RECT 513.200 409.600 514.000 410.400 ;
        RECT 542.000 417.600 542.800 418.400 ;
        RECT 532.400 413.600 533.200 414.400 ;
        RECT 566.000 417.600 566.800 418.400 ;
        RECT 545.200 413.600 546.000 414.400 ;
        RECT 516.400 405.600 517.200 406.400 ;
        RECT 551.600 409.600 552.400 410.400 ;
        RECT 569.200 413.600 570.000 414.400 ;
        RECT 558.000 409.600 558.800 410.400 ;
        RECT 583.600 413.000 584.400 413.800 ;
        RECT 574.000 409.600 574.800 410.400 ;
        RECT 593.200 412.600 594.000 413.400 ;
        RECT 578.800 411.600 579.600 412.400 ;
        RECT 599.600 411.600 600.400 412.400 ;
        RECT 585.200 408.800 586.000 409.600 ;
        RECT 590.000 407.600 590.800 408.400 ;
        RECT 572.400 403.600 573.200 404.400 ;
        RECT 586.800 406.200 587.600 407.000 ;
        RECT 583.600 404.200 584.400 405.000 ;
        RECT 585.200 404.200 586.000 405.000 ;
        RECT 590.000 406.200 590.800 407.000 ;
        RECT 593.200 406.200 594.000 407.000 ;
        RECT 594.800 404.200 595.600 405.000 ;
        RECT 596.400 404.200 597.200 405.000 ;
        RECT 598.000 404.200 598.800 405.000 ;
        RECT 607.600 403.600 608.400 404.400 ;
        RECT 18.800 395.000 19.600 395.800 ;
        RECT 15.600 393.600 16.400 394.400 ;
        RECT 20.400 392.400 21.200 393.200 ;
        RECT 36.400 393.600 37.200 394.400 ;
        RECT 25.200 389.600 26.000 390.400 ;
        RECT 9.200 388.200 10.000 389.000 ;
        RECT 18.800 388.600 19.600 389.400 ;
        RECT 14.000 387.600 14.800 388.400 ;
        RECT 9.200 384.200 10.000 385.000 ;
        RECT 10.800 384.200 11.600 385.000 ;
        RECT 12.400 384.200 13.200 385.000 ;
        RECT 15.600 384.200 16.400 385.000 ;
        RECT 18.800 384.200 19.600 385.000 ;
        RECT 20.400 384.200 21.200 385.000 ;
        RECT 22.000 384.200 22.800 385.000 ;
        RECT 23.600 384.200 24.400 385.000 ;
        RECT 42.800 397.600 43.600 398.400 ;
        RECT 65.200 397.600 66.000 398.400 ;
        RECT 39.600 387.600 40.400 388.400 ;
        RECT 46.000 389.600 46.800 390.400 ;
        RECT 54.000 389.600 54.800 390.400 ;
        RECT 38.000 383.600 38.800 384.400 ;
        RECT 42.800 383.600 43.600 384.400 ;
        RECT 47.600 386.200 48.400 387.000 ;
        RECT 78.000 387.600 78.800 388.400 ;
        RECT 86.000 389.600 86.800 390.400 ;
        RECT 98.800 397.600 99.600 398.400 ;
        RECT 95.600 389.600 96.400 390.400 ;
        RECT 97.200 389.600 98.000 390.400 ;
        RECT 70.000 383.600 70.800 384.400 ;
        RECT 130.800 393.600 131.600 394.400 ;
        RECT 100.400 385.600 101.200 386.400 ;
        RECT 106.800 389.600 107.600 390.400 ;
        RECT 119.600 389.600 120.400 390.400 ;
        RECT 103.600 383.600 104.400 384.400 ;
        RECT 111.600 385.600 112.400 386.400 ;
        RECT 113.200 386.200 114.000 387.000 ;
        RECT 134.000 389.600 134.800 390.400 ;
        RECT 158.000 397.600 158.800 398.400 ;
        RECT 142.000 389.600 142.800 390.400 ;
        RECT 143.600 387.600 144.400 388.400 ;
        RECT 161.200 397.600 162.000 398.400 ;
        RECT 167.600 397.600 168.400 398.400 ;
        RECT 178.800 394.400 179.600 395.200 ;
        RECT 182.000 395.000 182.800 395.800 ;
        RECT 202.800 397.600 203.600 398.400 ;
        RECT 177.200 392.400 178.000 393.200 ;
        RECT 161.200 383.600 162.000 384.400 ;
        RECT 186.800 387.600 187.600 388.400 ;
        RECT 183.600 385.600 184.400 386.400 ;
        RECT 177.200 384.200 178.000 385.000 ;
        RECT 178.800 384.200 179.600 385.000 ;
        RECT 180.400 384.200 181.200 385.000 ;
        RECT 182.000 384.200 182.800 385.000 ;
        RECT 185.200 384.200 186.000 385.000 ;
        RECT 188.400 384.200 189.200 385.000 ;
        RECT 190.000 384.200 190.800 385.000 ;
        RECT 191.600 384.200 192.400 385.000 ;
        RECT 201.200 385.600 202.000 386.400 ;
        RECT 231.600 395.000 232.400 395.800 ;
        RECT 228.400 393.600 229.200 394.400 ;
        RECT 233.200 392.400 234.000 393.200 ;
        RECT 246.000 393.600 246.800 394.400 ;
        RECT 207.600 387.600 208.400 388.400 ;
        RECT 210.800 387.600 211.600 388.400 ;
        RECT 212.400 387.600 213.200 388.400 ;
        RECT 222.000 388.200 222.800 389.000 ;
        RECT 231.600 388.600 232.400 389.400 ;
        RECT 226.800 387.600 227.600 388.400 ;
        RECT 222.000 384.200 222.800 385.000 ;
        RECT 223.600 384.200 224.400 385.000 ;
        RECT 225.200 384.200 226.000 385.000 ;
        RECT 228.400 384.200 229.200 385.000 ;
        RECT 231.600 384.200 232.400 385.000 ;
        RECT 233.200 384.200 234.000 385.000 ;
        RECT 234.800 384.200 235.600 385.000 ;
        RECT 236.400 384.200 237.200 385.000 ;
        RECT 249.200 387.600 250.000 388.400 ;
        RECT 257.200 389.600 258.000 390.400 ;
        RECT 252.400 383.600 253.200 384.400 ;
        RECT 263.600 389.600 264.400 390.400 ;
        RECT 282.800 395.000 283.600 395.800 ;
        RECT 279.600 393.600 280.400 394.400 ;
        RECT 297.200 397.600 298.000 398.400 ;
        RECT 284.400 392.400 285.200 393.200 ;
        RECT 289.200 389.600 290.000 390.400 ;
        RECT 273.200 388.200 274.000 389.000 ;
        RECT 282.800 388.600 283.600 389.400 ;
        RECT 260.400 383.600 261.200 384.400 ;
        RECT 278.000 387.600 278.800 388.400 ;
        RECT 273.200 384.200 274.000 385.000 ;
        RECT 274.800 384.200 275.600 385.000 ;
        RECT 276.400 384.200 277.200 385.000 ;
        RECT 279.600 384.200 280.400 385.000 ;
        RECT 282.800 384.200 283.600 385.000 ;
        RECT 284.400 384.200 285.200 385.000 ;
        RECT 286.000 384.200 286.800 385.000 ;
        RECT 287.600 384.200 288.400 385.000 ;
        RECT 322.800 395.000 323.600 395.800 ;
        RECT 319.600 393.600 320.400 394.400 ;
        RECT 337.200 397.600 338.000 398.400 ;
        RECT 324.400 392.400 325.200 393.200 ;
        RECT 342.000 397.600 342.800 398.400 ;
        RECT 313.200 388.200 314.000 389.000 ;
        RECT 322.800 388.600 323.600 389.400 ;
        RECT 318.000 387.600 318.800 388.400 ;
        RECT 313.200 384.200 314.000 385.000 ;
        RECT 314.800 384.200 315.600 385.000 ;
        RECT 316.400 384.200 317.200 385.000 ;
        RECT 319.600 384.200 320.400 385.000 ;
        RECT 322.800 384.200 323.600 385.000 ;
        RECT 324.400 384.200 325.200 385.000 ;
        RECT 326.000 384.200 326.800 385.000 ;
        RECT 327.600 384.200 328.400 385.000 ;
        RECT 353.200 394.400 354.000 395.200 ;
        RECT 356.400 395.000 357.200 395.800 ;
        RECT 351.600 392.400 352.400 393.200 ;
        RECT 337.200 383.600 338.000 384.400 ;
        RECT 393.200 397.600 394.000 398.400 ;
        RECT 361.200 387.600 362.000 388.400 ;
        RECT 358.000 385.600 358.800 386.400 ;
        RECT 351.600 384.200 352.400 385.000 ;
        RECT 353.200 384.200 354.000 385.000 ;
        RECT 354.800 384.200 355.600 385.000 ;
        RECT 356.400 384.200 357.200 385.000 ;
        RECT 359.600 384.200 360.400 385.000 ;
        RECT 362.800 384.200 363.600 385.000 ;
        RECT 364.400 384.200 365.200 385.000 ;
        RECT 366.000 384.200 366.800 385.000 ;
        RECT 375.600 386.200 376.400 387.000 ;
        RECT 396.400 397.600 397.200 398.400 ;
        RECT 394.800 385.600 395.600 386.400 ;
        RECT 399.600 397.600 400.400 398.400 ;
        RECT 398.000 385.600 398.800 386.400 ;
        RECT 409.200 393.600 410.000 394.400 ;
        RECT 420.400 394.400 421.200 395.200 ;
        RECT 423.600 395.000 424.400 395.800 ;
        RECT 418.800 392.400 419.600 393.200 ;
        RECT 404.400 383.600 405.200 384.400 ;
        RECT 409.200 383.600 410.000 384.400 ;
        RECT 428.400 387.600 429.200 388.400 ;
        RECT 425.200 385.600 426.000 386.400 ;
        RECT 418.800 384.200 419.600 385.000 ;
        RECT 420.400 384.200 421.200 385.000 ;
        RECT 422.000 384.200 422.800 385.000 ;
        RECT 423.600 384.200 424.400 385.000 ;
        RECT 426.800 384.200 427.600 385.000 ;
        RECT 430.000 384.200 430.800 385.000 ;
        RECT 431.600 384.200 432.400 385.000 ;
        RECT 433.200 384.200 434.000 385.000 ;
        RECT 450.800 389.600 451.600 390.400 ;
        RECT 476.400 395.000 477.200 395.800 ;
        RECT 473.200 393.600 474.000 394.400 ;
        RECT 490.800 397.600 491.600 398.400 ;
        RECT 478.000 392.400 478.800 393.200 ;
        RECT 510.000 397.600 510.800 398.400 ;
        RECT 482.800 389.600 483.600 390.400 ;
        RECT 452.400 387.600 453.200 388.400 ;
        RECT 466.800 388.200 467.600 389.000 ;
        RECT 476.400 388.600 477.200 389.400 ;
        RECT 471.600 387.600 472.400 388.400 ;
        RECT 466.800 384.200 467.600 385.000 ;
        RECT 468.400 384.200 469.200 385.000 ;
        RECT 470.000 384.200 470.800 385.000 ;
        RECT 473.200 384.200 474.000 385.000 ;
        RECT 476.400 384.200 477.200 385.000 ;
        RECT 478.000 384.200 478.800 385.000 ;
        RECT 479.600 384.200 480.400 385.000 ;
        RECT 481.200 384.200 482.000 385.000 ;
        RECT 535.600 395.000 536.400 395.800 ;
        RECT 532.400 393.600 533.200 394.400 ;
        RECT 537.200 392.400 538.000 393.200 ;
        RECT 561.200 393.600 562.000 394.400 ;
        RECT 542.000 389.600 542.800 390.400 ;
        RECT 514.800 387.600 515.600 388.400 ;
        RECT 511.600 385.600 512.400 386.400 ;
        RECT 516.400 387.600 517.200 388.400 ;
        RECT 526.000 388.200 526.800 389.000 ;
        RECT 535.600 388.600 536.400 389.400 ;
        RECT 530.800 387.600 531.600 388.400 ;
        RECT 550.200 389.600 551.000 390.400 ;
        RECT 526.000 384.200 526.800 385.000 ;
        RECT 527.600 384.200 528.400 385.000 ;
        RECT 529.200 384.200 530.000 385.000 ;
        RECT 532.400 384.200 533.200 385.000 ;
        RECT 535.600 384.200 536.400 385.000 ;
        RECT 537.200 384.200 538.000 385.000 ;
        RECT 538.800 384.200 539.600 385.000 ;
        RECT 540.400 384.200 541.200 385.000 ;
        RECT 561.200 389.600 562.000 390.400 ;
        RECT 556.400 385.600 557.200 386.400 ;
        RECT 554.800 383.600 555.600 384.400 ;
        RECT 566.000 385.600 566.800 386.400 ;
        RECT 591.600 395.000 592.400 395.800 ;
        RECT 588.400 393.600 589.200 394.400 ;
        RECT 606.000 397.600 606.800 398.400 ;
        RECT 593.200 392.400 594.000 393.200 ;
        RECT 570.800 387.600 571.600 388.400 ;
        RECT 582.000 388.200 582.800 389.000 ;
        RECT 591.600 388.600 592.400 389.400 ;
        RECT 572.400 385.600 573.200 386.400 ;
        RECT 586.800 387.600 587.600 388.400 ;
        RECT 582.000 384.200 582.800 385.000 ;
        RECT 583.600 384.200 584.400 385.000 ;
        RECT 585.200 384.200 586.000 385.000 ;
        RECT 588.400 384.200 589.200 385.000 ;
        RECT 591.600 384.200 592.400 385.000 ;
        RECT 593.200 384.200 594.000 385.000 ;
        RECT 594.800 384.200 595.600 385.000 ;
        RECT 596.400 384.200 597.200 385.000 ;
        RECT 12.400 377.600 13.200 378.400 ;
        RECT 6.000 373.600 6.800 374.400 ;
        RECT 39.600 377.600 40.400 378.400 ;
        RECT 12.400 369.600 13.200 370.400 ;
        RECT 31.600 369.600 32.400 370.400 ;
        RECT 46.000 369.600 46.800 370.400 ;
        RECT 92.400 377.600 93.200 378.400 ;
        RECT 52.400 373.600 53.200 374.400 ;
        RECT 63.600 371.600 64.400 372.400 ;
        RECT 108.400 373.600 109.200 374.400 ;
        RECT 97.200 372.200 98.000 373.000 ;
        RECT 84.400 369.600 85.200 370.400 ;
        RECT 89.200 369.600 90.000 370.400 ;
        RECT 110.000 370.200 110.800 371.000 ;
        RECT 114.800 377.600 115.600 378.400 ;
        RECT 142.000 377.600 142.800 378.400 ;
        RECT 172.400 377.600 173.200 378.400 ;
        RECT 156.400 373.600 157.200 374.400 ;
        RECT 166.000 373.600 166.800 374.400 ;
        RECT 126.000 369.600 126.800 370.400 ;
        RECT 132.400 367.600 133.200 368.400 ;
        RECT 142.000 369.600 142.800 370.400 ;
        RECT 159.600 371.800 160.400 372.600 ;
        RECT 148.400 369.600 149.200 370.400 ;
        RECT 154.800 370.200 155.600 371.000 ;
        RECT 182.000 373.000 182.800 373.800 ;
        RECT 191.600 372.600 192.400 373.400 ;
        RECT 214.000 377.600 214.800 378.400 ;
        RECT 231.600 377.600 232.400 378.400 ;
        RECT 198.000 371.600 198.800 372.400 ;
        RECT 183.600 368.800 184.400 369.600 ;
        RECT 188.400 367.600 189.200 368.400 ;
        RECT 185.200 366.200 186.000 367.000 ;
        RECT 182.000 364.200 182.800 365.000 ;
        RECT 183.600 364.200 184.400 365.000 ;
        RECT 188.400 366.200 189.200 367.000 ;
        RECT 191.600 366.200 192.400 367.000 ;
        RECT 193.200 364.200 194.000 365.000 ;
        RECT 194.800 364.200 195.600 365.000 ;
        RECT 196.400 364.200 197.200 365.000 ;
        RECT 206.000 369.600 206.800 370.400 ;
        RECT 209.200 369.600 210.000 370.400 ;
        RECT 250.800 375.600 251.600 376.400 ;
        RECT 252.400 374.200 253.200 375.000 ;
        RECT 263.600 371.600 264.400 372.400 ;
        RECT 210.800 363.600 211.600 364.400 ;
        RECT 231.600 367.600 232.400 368.400 ;
        RECT 246.000 366.800 246.800 367.600 ;
        RECT 249.200 366.200 250.000 367.000 ;
        RECT 244.400 364.200 245.200 365.000 ;
        RECT 246.000 364.200 246.800 365.000 ;
        RECT 247.600 364.200 248.400 365.000 ;
        RECT 252.400 366.200 253.200 367.000 ;
        RECT 255.600 366.200 256.400 367.000 ;
        RECT 286.000 377.600 286.800 378.400 ;
        RECT 300.400 377.600 301.200 378.400 ;
        RECT 313.200 377.600 314.000 378.400 ;
        RECT 270.000 373.600 270.800 374.400 ;
        RECT 274.800 373.600 275.600 374.400 ;
        RECT 289.200 373.600 290.000 374.400 ;
        RECT 257.200 364.200 258.000 365.000 ;
        RECT 258.800 364.200 259.600 365.000 ;
        RECT 286.000 363.600 286.800 364.400 ;
        RECT 321.200 377.600 322.000 378.400 ;
        RECT 351.600 373.000 352.400 373.800 ;
        RECT 361.200 372.600 362.000 373.400 ;
        RECT 375.600 377.600 376.400 378.400 ;
        RECT 346.800 371.600 347.600 372.400 ;
        RECT 367.600 371.600 368.400 372.400 ;
        RECT 353.200 368.800 354.000 369.600 ;
        RECT 358.000 367.600 358.800 368.400 ;
        RECT 354.800 366.200 355.600 367.000 ;
        RECT 351.600 364.200 352.400 365.000 ;
        RECT 353.200 364.200 354.000 365.000 ;
        RECT 358.000 366.200 358.800 367.000 ;
        RECT 361.200 366.200 362.000 367.000 ;
        RECT 362.800 364.200 363.600 365.000 ;
        RECT 364.400 364.200 365.200 365.000 ;
        RECT 366.000 364.200 366.800 365.000 ;
        RECT 396.400 375.600 397.200 376.400 ;
        RECT 398.000 374.200 398.800 375.000 ;
        RECT 407.600 371.600 408.400 372.400 ;
        RECT 380.400 369.600 381.200 370.400 ;
        RECT 391.600 366.800 392.400 367.600 ;
        RECT 394.800 366.200 395.600 367.000 ;
        RECT 390.000 364.200 390.800 365.000 ;
        RECT 391.600 364.200 392.400 365.000 ;
        RECT 393.200 364.200 394.000 365.000 ;
        RECT 398.000 366.200 398.800 367.000 ;
        RECT 401.200 366.200 402.000 367.000 ;
        RECT 402.800 364.200 403.600 365.000 ;
        RECT 404.400 364.200 405.200 365.000 ;
        RECT 420.400 369.600 421.200 370.400 ;
        RECT 465.200 375.600 466.000 376.400 ;
        RECT 466.800 374.200 467.600 375.000 ;
        RECT 457.200 371.600 458.000 372.400 ;
        RECT 478.000 371.600 478.800 372.400 ;
        RECT 449.200 369.600 450.000 370.400 ;
        RECT 460.400 366.800 461.200 367.600 ;
        RECT 463.600 366.200 464.400 367.000 ;
        RECT 458.800 364.200 459.600 365.000 ;
        RECT 460.400 364.200 461.200 365.000 ;
        RECT 462.000 364.200 462.800 365.000 ;
        RECT 466.800 366.200 467.600 367.000 ;
        RECT 470.000 366.200 470.800 367.000 ;
        RECT 471.600 364.200 472.400 365.000 ;
        RECT 473.200 364.200 474.000 365.000 ;
        RECT 508.400 377.600 509.200 378.400 ;
        RECT 498.800 373.600 499.600 374.400 ;
        RECT 482.800 363.600 483.600 364.400 ;
        RECT 514.800 377.600 515.600 378.400 ;
        RECT 505.200 371.600 506.000 372.400 ;
        RECT 511.600 371.600 512.400 372.400 ;
        RECT 537.200 375.600 538.000 376.400 ;
        RECT 538.800 374.200 539.600 375.000 ;
        RECT 546.800 370.000 547.600 370.800 ;
        RECT 521.200 363.600 522.000 364.400 ;
        RECT 532.400 366.800 533.200 367.600 ;
        RECT 535.600 366.200 536.400 367.000 ;
        RECT 530.800 364.200 531.600 365.000 ;
        RECT 532.400 364.200 533.200 365.000 ;
        RECT 534.000 364.200 534.800 365.000 ;
        RECT 538.800 366.200 539.600 367.000 ;
        RECT 542.000 366.200 542.800 367.000 ;
        RECT 562.800 375.600 563.600 376.400 ;
        RECT 543.600 364.200 544.400 365.000 ;
        RECT 545.200 364.200 546.000 365.000 ;
        RECT 561.200 369.600 562.000 370.400 ;
        RECT 569.200 373.600 570.000 374.400 ;
        RECT 590.000 375.600 590.800 376.400 ;
        RECT 591.600 374.200 592.400 375.000 ;
        RECT 582.000 371.600 582.800 372.400 ;
        RECT 570.800 367.600 571.600 368.400 ;
        RECT 585.200 366.800 586.000 367.600 ;
        RECT 588.400 366.200 589.200 367.000 ;
        RECT 583.600 364.200 584.400 365.000 ;
        RECT 585.200 364.200 586.000 365.000 ;
        RECT 586.800 364.200 587.600 365.000 ;
        RECT 591.600 366.200 592.400 367.000 ;
        RECT 594.800 366.200 595.600 367.000 ;
        RECT 596.400 364.200 597.200 365.000 ;
        RECT 598.000 364.200 598.800 365.000 ;
        RECT 6.000 349.600 6.800 350.400 ;
        RECT 28.400 355.000 29.200 355.800 ;
        RECT 25.200 353.600 26.000 354.400 ;
        RECT 30.000 352.400 30.800 353.200 ;
        RECT 42.800 353.600 43.600 354.400 ;
        RECT 47.600 357.600 48.400 358.400 ;
        RECT 18.800 348.200 19.600 349.000 ;
        RECT 28.400 348.600 29.200 349.400 ;
        RECT 9.200 343.600 10.000 344.400 ;
        RECT 23.600 347.600 24.400 348.400 ;
        RECT 18.800 344.200 19.600 345.000 ;
        RECT 20.400 344.200 21.200 345.000 ;
        RECT 22.000 344.200 22.800 345.000 ;
        RECT 25.200 344.200 26.000 345.000 ;
        RECT 28.400 344.200 29.200 345.000 ;
        RECT 30.000 344.200 30.800 345.000 ;
        RECT 31.600 344.200 32.400 345.000 ;
        RECT 33.200 344.200 34.000 345.000 ;
        RECT 49.200 357.600 50.000 358.400 ;
        RECT 57.200 357.600 58.000 358.400 ;
        RECT 50.800 345.600 51.600 346.400 ;
        RECT 55.600 347.600 56.400 348.400 ;
        RECT 78.000 357.600 78.800 358.400 ;
        RECT 58.800 345.600 59.600 346.400 ;
        RECT 60.400 346.200 61.200 347.000 ;
        RECT 79.600 357.600 80.400 358.400 ;
        RECT 97.200 353.600 98.000 354.400 ;
        RECT 81.200 345.600 82.000 346.400 ;
        RECT 90.800 351.600 91.600 352.400 ;
        RECT 90.800 349.600 91.600 350.400 ;
        RECT 86.000 347.600 86.800 348.400 ;
        RECT 92.400 347.600 93.200 348.400 ;
        RECT 98.800 347.600 99.600 348.400 ;
        RECT 103.600 349.600 104.400 350.400 ;
        RECT 105.200 349.600 106.000 350.400 ;
        RECT 114.800 349.600 115.600 350.400 ;
        RECT 122.800 349.600 123.600 350.400 ;
        RECT 129.200 349.600 130.000 350.400 ;
        RECT 132.400 349.600 133.200 350.400 ;
        RECT 134.000 349.600 134.800 350.400 ;
        RECT 102.000 345.600 102.800 346.400 ;
        RECT 116.400 347.600 117.200 348.400 ;
        RECT 124.400 347.600 125.200 348.400 ;
        RECT 127.600 347.600 128.400 348.400 ;
        RECT 130.800 347.600 131.600 348.400 ;
        RECT 153.200 357.600 154.000 358.400 ;
        RECT 153.200 343.600 154.000 344.400 ;
        RECT 170.800 349.600 171.600 350.400 ;
        RECT 172.400 349.600 173.200 350.400 ;
        RECT 174.000 349.600 174.800 350.400 ;
        RECT 169.200 343.600 170.000 344.400 ;
        RECT 196.400 355.000 197.200 355.800 ;
        RECT 193.200 353.600 194.000 354.400 ;
        RECT 210.800 357.600 211.600 358.400 ;
        RECT 198.000 352.400 198.800 353.200 ;
        RECT 202.800 349.600 203.600 350.400 ;
        RECT 186.800 348.200 187.600 349.000 ;
        RECT 196.400 348.600 197.200 349.400 ;
        RECT 191.600 347.600 192.400 348.400 ;
        RECT 186.800 344.200 187.600 345.000 ;
        RECT 188.400 344.200 189.200 345.000 ;
        RECT 190.000 344.200 190.800 345.000 ;
        RECT 193.200 344.200 194.000 345.000 ;
        RECT 196.400 344.200 197.200 345.000 ;
        RECT 198.000 344.200 198.800 345.000 ;
        RECT 199.600 344.200 200.400 345.000 ;
        RECT 201.200 344.200 202.000 345.000 ;
        RECT 222.000 357.600 222.800 358.400 ;
        RECT 218.800 349.600 219.600 350.400 ;
        RECT 252.400 355.000 253.200 355.800 ;
        RECT 249.200 353.600 250.000 354.400 ;
        RECT 266.800 357.600 267.600 358.400 ;
        RECT 254.000 352.400 254.800 353.200 ;
        RECT 258.800 349.600 259.600 350.400 ;
        RECT 242.800 348.200 243.600 349.000 ;
        RECT 252.400 348.600 253.200 349.400 ;
        RECT 247.600 347.600 248.400 348.400 ;
        RECT 242.800 344.200 243.600 345.000 ;
        RECT 244.400 344.200 245.200 345.000 ;
        RECT 246.000 344.200 246.800 345.000 ;
        RECT 249.200 344.200 250.000 345.000 ;
        RECT 252.400 344.200 253.200 345.000 ;
        RECT 254.000 344.200 254.800 345.000 ;
        RECT 255.600 344.200 256.400 345.000 ;
        RECT 257.200 344.200 258.000 345.000 ;
        RECT 270.000 349.600 270.800 350.400 ;
        RECT 271.600 349.600 272.400 350.400 ;
        RECT 284.400 357.600 285.200 358.400 ;
        RECT 281.200 345.600 282.000 346.400 ;
        RECT 282.800 345.600 283.600 346.400 ;
        RECT 303.600 355.000 304.400 355.800 ;
        RECT 300.400 353.600 301.200 354.400 ;
        RECT 305.200 352.400 306.000 353.200 ;
        RECT 310.000 349.600 310.800 350.400 ;
        RECT 294.000 348.200 294.800 349.000 ;
        RECT 303.600 348.600 304.400 349.400 ;
        RECT 298.800 347.600 299.600 348.400 ;
        RECT 318.200 349.600 319.000 350.400 ;
        RECT 294.000 344.200 294.800 345.000 ;
        RECT 295.600 344.200 296.400 345.000 ;
        RECT 297.200 344.200 298.000 345.000 ;
        RECT 300.400 344.200 301.200 345.000 ;
        RECT 303.600 344.200 304.400 345.000 ;
        RECT 305.200 344.200 306.000 345.000 ;
        RECT 306.800 344.200 307.600 345.000 ;
        RECT 308.400 344.200 309.200 345.000 ;
        RECT 327.600 349.600 328.400 350.400 ;
        RECT 356.400 355.000 357.200 355.800 ;
        RECT 353.200 353.600 354.000 354.400 ;
        RECT 358.000 352.400 358.800 353.200 ;
        RECT 362.800 349.600 363.600 350.400 ;
        RECT 346.800 348.200 347.600 349.000 ;
        RECT 356.400 348.600 357.200 349.400 ;
        RECT 337.200 345.600 338.000 346.400 ;
        RECT 351.600 347.600 352.400 348.400 ;
        RECT 346.800 344.200 347.600 345.000 ;
        RECT 348.400 344.200 349.200 345.000 ;
        RECT 350.000 344.200 350.800 345.000 ;
        RECT 353.200 344.200 354.000 345.000 ;
        RECT 356.400 344.200 357.200 345.000 ;
        RECT 358.000 344.200 358.800 345.000 ;
        RECT 359.600 344.200 360.400 345.000 ;
        RECT 361.200 344.200 362.000 345.000 ;
        RECT 374.000 345.600 374.800 346.400 ;
        RECT 370.800 343.600 371.600 344.400 ;
        RECT 394.800 351.600 395.600 352.400 ;
        RECT 388.400 349.600 389.200 350.400 ;
        RECT 390.000 349.600 390.800 350.400 ;
        RECT 398.000 349.600 398.800 350.400 ;
        RECT 399.600 349.600 400.400 350.400 ;
        RECT 380.400 343.600 381.200 344.400 ;
        RECT 404.400 347.600 405.200 348.400 ;
        RECT 402.800 343.600 403.600 344.400 ;
        RECT 409.200 347.600 410.000 348.400 ;
        RECT 407.600 345.600 408.400 346.400 ;
        RECT 426.800 354.400 427.600 355.200 ;
        RECT 430.000 355.000 430.800 355.800 ;
        RECT 425.200 352.400 426.000 353.200 ;
        RECT 423.600 349.600 424.400 350.400 ;
        RECT 415.600 345.600 416.400 346.400 ;
        RECT 434.800 347.600 435.600 348.400 ;
        RECT 431.600 345.600 432.400 346.400 ;
        RECT 471.600 354.400 472.400 355.200 ;
        RECT 474.800 355.000 475.600 355.800 ;
        RECT 470.000 352.400 470.800 353.200 ;
        RECT 425.200 344.200 426.000 345.000 ;
        RECT 426.800 344.200 427.600 345.000 ;
        RECT 428.400 344.200 429.200 345.000 ;
        RECT 430.000 344.200 430.800 345.000 ;
        RECT 433.200 344.200 434.000 345.000 ;
        RECT 436.400 344.200 437.200 345.000 ;
        RECT 438.000 344.200 438.800 345.000 ;
        RECT 439.600 344.200 440.400 345.000 ;
        RECT 449.200 345.600 450.000 346.400 ;
        RECT 460.200 347.600 461.000 348.400 ;
        RECT 479.600 347.600 480.400 348.400 ;
        RECT 476.400 345.600 477.200 346.400 ;
        RECT 470.000 344.200 470.800 345.000 ;
        RECT 471.600 344.200 472.400 345.000 ;
        RECT 473.200 344.200 474.000 345.000 ;
        RECT 474.800 344.200 475.600 345.000 ;
        RECT 478.000 344.200 478.800 345.000 ;
        RECT 481.200 344.200 482.000 345.000 ;
        RECT 482.800 344.200 483.600 345.000 ;
        RECT 484.400 344.200 485.200 345.000 ;
        RECT 511.600 355.000 512.400 355.800 ;
        RECT 508.400 353.600 509.200 354.400 ;
        RECT 513.200 352.400 514.000 353.200 ;
        RECT 518.000 349.600 518.800 350.400 ;
        RECT 502.000 348.200 502.800 349.000 ;
        RECT 511.600 348.600 512.400 349.400 ;
        RECT 506.800 347.600 507.600 348.400 ;
        RECT 502.000 344.200 502.800 345.000 ;
        RECT 503.600 344.200 504.400 345.000 ;
        RECT 505.200 344.200 506.000 345.000 ;
        RECT 508.400 344.200 509.200 345.000 ;
        RECT 511.600 344.200 512.400 345.000 ;
        RECT 513.200 344.200 514.000 345.000 ;
        RECT 514.800 344.200 515.600 345.000 ;
        RECT 516.400 344.200 517.200 345.000 ;
        RECT 529.200 347.600 530.000 348.400 ;
        RECT 538.800 349.600 539.600 350.400 ;
        RECT 551.600 357.600 552.400 358.400 ;
        RECT 526.000 343.600 526.800 344.400 ;
        RECT 535.600 343.600 536.400 344.400 ;
        RECT 583.600 355.000 584.400 355.800 ;
        RECT 580.400 353.600 581.200 354.400 ;
        RECT 585.200 352.400 586.000 353.200 ;
        RECT 590.000 349.600 590.800 350.400 ;
        RECT 558.000 347.600 558.800 348.400 ;
        RECT 574.000 348.200 574.800 349.000 ;
        RECT 583.600 348.600 584.400 349.400 ;
        RECT 578.800 347.600 579.600 348.400 ;
        RECT 598.200 349.600 599.000 350.400 ;
        RECT 574.000 344.200 574.800 345.000 ;
        RECT 575.600 344.200 576.400 345.000 ;
        RECT 577.200 344.200 578.000 345.000 ;
        RECT 580.400 344.200 581.200 345.000 ;
        RECT 583.600 344.200 584.400 345.000 ;
        RECT 585.200 344.200 586.000 345.000 ;
        RECT 586.800 344.200 587.600 345.000 ;
        RECT 588.400 344.200 589.200 345.000 ;
        RECT 9.200 333.000 10.000 333.800 ;
        RECT 18.800 332.600 19.600 333.400 ;
        RECT 7.600 331.600 8.400 332.400 ;
        RECT 10.800 328.800 11.600 329.600 ;
        RECT 15.600 327.600 16.400 328.400 ;
        RECT 12.400 326.200 13.200 327.000 ;
        RECT 9.200 324.200 10.000 325.000 ;
        RECT 10.800 324.200 11.600 325.000 ;
        RECT 15.600 326.200 16.400 327.000 ;
        RECT 18.800 326.200 19.600 327.000 ;
        RECT 20.400 324.200 21.200 325.000 ;
        RECT 22.000 324.200 22.800 325.000 ;
        RECT 23.600 324.200 24.400 325.000 ;
        RECT 38.000 323.600 38.800 324.400 ;
        RECT 60.400 337.600 61.200 338.400 ;
        RECT 76.400 335.600 77.200 336.400 ;
        RECT 78.000 334.200 78.800 335.000 ;
        RECT 79.600 331.600 80.400 332.400 ;
        RECT 57.200 323.600 58.000 324.400 ;
        RECT 71.600 326.800 72.400 327.600 ;
        RECT 74.800 326.200 75.600 327.000 ;
        RECT 70.000 324.200 70.800 325.000 ;
        RECT 71.600 324.200 72.400 325.000 ;
        RECT 73.200 324.200 74.000 325.000 ;
        RECT 78.000 326.200 78.800 327.000 ;
        RECT 81.200 326.200 82.000 327.000 ;
        RECT 124.400 337.600 125.200 338.400 ;
        RECT 82.800 324.200 83.600 325.000 ;
        RECT 84.400 324.200 85.200 325.000 ;
        RECT 108.400 333.600 109.200 334.400 ;
        RECT 143.600 337.600 144.400 338.400 ;
        RECT 106.800 330.200 107.600 331.000 ;
        RECT 134.000 333.600 134.800 334.400 ;
        RECT 130.800 331.800 131.600 332.600 ;
        RECT 126.000 330.200 126.800 331.000 ;
        RECT 145.200 337.600 146.000 338.400 ;
        RECT 154.800 337.600 155.600 338.400 ;
        RECT 170.800 335.600 171.600 336.400 ;
        RECT 172.400 334.200 173.200 335.000 ;
        RECT 180.400 331.600 181.200 332.400 ;
        RECT 183.600 331.600 184.400 332.400 ;
        RECT 166.000 326.800 166.800 327.600 ;
        RECT 169.200 326.200 170.000 327.000 ;
        RECT 164.400 324.200 165.200 325.000 ;
        RECT 166.000 324.200 166.800 325.000 ;
        RECT 167.600 324.200 168.400 325.000 ;
        RECT 172.400 326.200 173.200 327.000 ;
        RECT 175.600 326.200 176.400 327.000 ;
        RECT 177.200 324.200 178.000 325.000 ;
        RECT 178.800 324.200 179.600 325.000 ;
        RECT 202.800 333.000 203.600 333.800 ;
        RECT 212.400 332.600 213.200 333.400 ;
        RECT 226.800 337.600 227.600 338.400 ;
        RECT 218.800 331.600 219.600 332.400 ;
        RECT 234.800 337.600 235.600 338.400 ;
        RECT 204.400 328.800 205.200 329.600 ;
        RECT 209.200 327.600 210.000 328.400 ;
        RECT 206.000 326.200 206.800 327.000 ;
        RECT 202.800 324.200 203.600 325.000 ;
        RECT 204.400 324.200 205.200 325.000 ;
        RECT 209.200 326.200 210.000 327.000 ;
        RECT 212.400 326.200 213.200 327.000 ;
        RECT 214.000 324.200 214.800 325.000 ;
        RECT 215.600 324.200 216.400 325.000 ;
        RECT 217.200 324.200 218.000 325.000 ;
        RECT 249.200 333.000 250.000 333.800 ;
        RECT 258.800 332.600 259.600 333.400 ;
        RECT 273.200 335.600 274.000 336.400 ;
        RECT 254.000 331.600 254.800 332.400 ;
        RECT 250.800 328.800 251.600 329.600 ;
        RECT 255.600 327.600 256.400 328.400 ;
        RECT 239.600 323.600 240.400 324.400 ;
        RECT 252.400 326.200 253.200 327.000 ;
        RECT 249.200 324.200 250.000 325.000 ;
        RECT 250.800 324.200 251.600 325.000 ;
        RECT 255.600 326.200 256.400 327.000 ;
        RECT 258.800 326.200 259.600 327.000 ;
        RECT 260.400 324.200 261.200 325.000 ;
        RECT 262.000 324.200 262.800 325.000 ;
        RECT 263.600 324.200 264.400 325.000 ;
        RECT 314.800 331.600 315.600 332.400 ;
        RECT 327.600 333.600 328.400 334.400 ;
        RECT 276.400 323.600 277.200 324.400 ;
        RECT 279.600 323.600 280.400 324.400 ;
        RECT 289.200 323.600 290.000 324.400 ;
        RECT 295.600 323.600 296.400 324.400 ;
        RECT 302.000 323.600 302.800 324.400 ;
        RECT 353.200 335.600 354.000 336.400 ;
        RECT 354.800 334.200 355.600 335.000 ;
        RECT 378.800 337.600 379.600 338.400 ;
        RECT 377.200 333.600 378.000 334.400 ;
        RECT 362.800 331.600 363.600 332.400 ;
        RECT 337.200 329.600 338.000 330.400 ;
        RECT 348.400 326.800 349.200 327.600 ;
        RECT 351.600 326.200 352.400 327.000 ;
        RECT 346.800 324.200 347.600 325.000 ;
        RECT 348.400 324.200 349.200 325.000 ;
        RECT 350.000 324.200 350.800 325.000 ;
        RECT 354.800 326.200 355.600 327.000 ;
        RECT 358.000 326.200 358.800 327.000 ;
        RECT 374.000 327.600 374.800 328.400 ;
        RECT 359.600 324.200 360.400 325.000 ;
        RECT 361.200 324.200 362.000 325.000 ;
        RECT 385.200 329.600 386.000 330.400 ;
        RECT 391.600 333.600 392.400 334.400 ;
        RECT 414.000 335.600 414.800 336.400 ;
        RECT 415.600 334.200 416.400 335.000 ;
        RECT 423.600 331.600 424.400 332.400 ;
        RECT 398.000 323.600 398.800 324.400 ;
        RECT 409.200 326.800 410.000 327.600 ;
        RECT 412.400 326.200 413.200 327.000 ;
        RECT 407.600 324.200 408.400 325.000 ;
        RECT 409.200 324.200 410.000 325.000 ;
        RECT 410.800 324.200 411.600 325.000 ;
        RECT 415.600 326.200 416.400 327.000 ;
        RECT 418.800 326.200 419.600 327.000 ;
        RECT 431.600 329.600 432.400 330.400 ;
        RECT 420.400 324.200 421.200 325.000 ;
        RECT 422.000 324.200 422.800 325.000 ;
        RECT 433.200 323.600 434.000 324.400 ;
        RECT 450.800 333.600 451.600 334.400 ;
        RECT 444.400 329.600 445.200 330.400 ;
        RECT 450.800 329.600 451.600 330.400 ;
        RECT 455.600 329.600 456.400 330.400 ;
        RECT 471.600 331.600 472.400 332.400 ;
        RECT 466.800 327.600 467.600 328.400 ;
        RECT 474.800 323.600 475.600 324.400 ;
        RECT 490.800 335.600 491.600 336.400 ;
        RECT 487.600 329.600 488.400 330.400 ;
        RECT 486.000 323.600 486.800 324.400 ;
        RECT 500.400 331.600 501.200 332.400 ;
        RECT 522.800 335.600 523.600 336.400 ;
        RECT 524.400 334.200 525.200 335.000 ;
        RECT 535.600 331.600 536.400 332.400 ;
        RECT 490.800 323.600 491.600 324.400 ;
        RECT 498.800 323.600 499.600 324.400 ;
        RECT 502.000 323.600 502.800 324.400 ;
        RECT 506.800 323.600 507.600 324.400 ;
        RECT 518.000 326.800 518.800 327.600 ;
        RECT 521.200 326.200 522.000 327.000 ;
        RECT 516.400 324.200 517.200 325.000 ;
        RECT 518.000 324.200 518.800 325.000 ;
        RECT 519.600 324.200 520.400 325.000 ;
        RECT 524.400 326.200 525.200 327.000 ;
        RECT 527.600 326.200 528.400 327.000 ;
        RECT 548.400 333.000 549.200 333.800 ;
        RECT 558.000 332.600 558.800 333.400 ;
        RECT 572.400 337.600 573.200 338.400 ;
        RECT 580.400 337.600 581.200 338.400 ;
        RECT 543.600 331.600 544.400 332.400 ;
        RECT 550.000 328.800 550.800 329.600 ;
        RECT 554.800 327.600 555.600 328.400 ;
        RECT 529.200 324.200 530.000 325.000 ;
        RECT 530.800 324.200 531.600 325.000 ;
        RECT 551.600 326.200 552.400 327.000 ;
        RECT 548.400 324.200 549.200 325.000 ;
        RECT 550.000 324.200 550.800 325.000 ;
        RECT 554.800 326.200 555.600 327.000 ;
        RECT 558.000 326.200 558.800 327.000 ;
        RECT 559.600 324.200 560.400 325.000 ;
        RECT 561.200 324.200 562.000 325.000 ;
        RECT 562.800 324.200 563.600 325.000 ;
        RECT 593.200 329.600 594.000 330.400 ;
        RECT 606.000 337.600 606.800 338.400 ;
        RECT 591.600 323.600 592.400 324.400 ;
        RECT 12.400 317.600 13.200 318.400 ;
        RECT 33.200 315.000 34.000 315.800 ;
        RECT 30.000 313.600 30.800 314.400 ;
        RECT 47.600 317.600 48.400 318.400 ;
        RECT 34.800 312.400 35.600 313.200 ;
        RECT 52.400 317.600 53.200 318.400 ;
        RECT 23.600 308.200 24.400 309.000 ;
        RECT 33.200 308.600 34.000 309.400 ;
        RECT 28.400 307.600 29.200 308.400 ;
        RECT 23.600 304.200 24.400 305.000 ;
        RECT 25.200 304.200 26.000 305.000 ;
        RECT 26.800 304.200 27.600 305.000 ;
        RECT 30.000 304.200 30.800 305.000 ;
        RECT 33.200 304.200 34.000 305.000 ;
        RECT 34.800 304.200 35.600 305.000 ;
        RECT 36.400 304.200 37.200 305.000 ;
        RECT 38.000 304.200 38.800 305.000 ;
        RECT 63.600 314.400 64.400 315.200 ;
        RECT 66.800 315.000 67.600 315.800 ;
        RECT 62.000 312.400 62.800 313.200 ;
        RECT 71.600 307.600 72.400 308.400 ;
        RECT 68.400 305.600 69.200 306.400 ;
        RECT 62.000 304.200 62.800 305.000 ;
        RECT 63.600 304.200 64.400 305.000 ;
        RECT 65.200 304.200 66.000 305.000 ;
        RECT 66.800 304.200 67.600 305.000 ;
        RECT 70.000 304.200 70.800 305.000 ;
        RECT 73.200 304.200 74.000 305.000 ;
        RECT 74.800 304.200 75.600 305.000 ;
        RECT 76.400 304.200 77.200 305.000 ;
        RECT 92.400 309.600 93.200 310.400 ;
        RECT 95.600 309.600 96.400 310.400 ;
        RECT 97.200 309.600 98.000 310.400 ;
        RECT 110.000 317.600 110.800 318.400 ;
        RECT 121.200 314.400 122.000 315.200 ;
        RECT 124.400 315.000 125.200 315.800 ;
        RECT 119.600 312.400 120.400 313.200 ;
        RECT 118.000 309.600 118.800 310.400 ;
        RECT 161.200 317.600 162.000 318.400 ;
        RECT 129.200 307.600 130.000 308.400 ;
        RECT 126.000 305.600 126.800 306.400 ;
        RECT 172.400 314.400 173.200 315.200 ;
        RECT 175.600 315.000 176.400 315.800 ;
        RECT 196.400 317.600 197.200 318.400 ;
        RECT 170.800 312.400 171.600 313.200 ;
        RECT 119.600 304.200 120.400 305.000 ;
        RECT 121.200 304.200 122.000 305.000 ;
        RECT 122.800 304.200 123.600 305.000 ;
        RECT 124.400 304.200 125.200 305.000 ;
        RECT 127.600 304.200 128.400 305.000 ;
        RECT 130.800 304.200 131.600 305.000 ;
        RECT 132.400 304.200 133.200 305.000 ;
        RECT 134.000 304.200 134.800 305.000 ;
        RECT 143.600 305.600 144.400 306.400 ;
        RECT 169.200 309.600 170.000 310.400 ;
        RECT 154.800 303.600 155.600 304.400 ;
        RECT 161.200 303.600 162.000 304.400 ;
        RECT 194.800 311.600 195.600 312.400 ;
        RECT 180.400 307.600 181.200 308.400 ;
        RECT 177.200 305.600 178.000 306.400 ;
        RECT 170.800 304.200 171.600 305.000 ;
        RECT 172.400 304.200 173.200 305.000 ;
        RECT 174.000 304.200 174.800 305.000 ;
        RECT 175.600 304.200 176.400 305.000 ;
        RECT 178.800 304.200 179.600 305.000 ;
        RECT 182.000 304.200 182.800 305.000 ;
        RECT 183.600 304.200 184.400 305.000 ;
        RECT 185.200 304.200 186.000 305.000 ;
        RECT 218.800 315.000 219.600 315.800 ;
        RECT 215.600 313.600 216.400 314.400 ;
        RECT 220.400 312.400 221.200 313.200 ;
        RECT 236.400 317.600 237.200 318.400 ;
        RECT 209.200 308.200 210.000 309.000 ;
        RECT 218.800 308.600 219.600 309.400 ;
        RECT 214.000 307.600 214.800 308.400 ;
        RECT 233.400 309.600 234.200 310.400 ;
        RECT 209.200 304.200 210.000 305.000 ;
        RECT 210.800 304.200 211.600 305.000 ;
        RECT 212.400 304.200 213.200 305.000 ;
        RECT 215.600 304.200 216.400 305.000 ;
        RECT 218.800 304.200 219.600 305.000 ;
        RECT 220.400 304.200 221.200 305.000 ;
        RECT 222.000 304.200 222.800 305.000 ;
        RECT 223.600 304.200 224.400 305.000 ;
        RECT 238.000 307.600 238.800 308.400 ;
        RECT 262.000 309.600 262.800 310.400 ;
        RECT 265.200 309.600 266.000 310.400 ;
        RECT 266.800 309.600 267.600 310.400 ;
        RECT 278.000 309.600 278.800 310.400 ;
        RECT 279.600 307.600 280.400 308.400 ;
        RECT 282.800 307.600 283.600 308.400 ;
        RECT 310.000 314.400 310.800 315.200 ;
        RECT 313.200 315.000 314.000 315.800 ;
        RECT 308.400 312.400 309.200 313.200 ;
        RECT 287.600 307.600 288.400 308.400 ;
        RECT 298.600 307.600 299.400 308.400 ;
        RECT 306.800 309.600 307.600 310.400 ;
        RECT 289.200 303.600 290.000 304.400 ;
        RECT 318.000 307.600 318.800 308.400 ;
        RECT 314.800 305.600 315.600 306.400 ;
        RECT 308.400 304.200 309.200 305.000 ;
        RECT 310.000 304.200 310.800 305.000 ;
        RECT 311.600 304.200 312.400 305.000 ;
        RECT 313.200 304.200 314.000 305.000 ;
        RECT 316.400 304.200 317.200 305.000 ;
        RECT 319.600 304.200 320.400 305.000 ;
        RECT 321.200 304.200 322.000 305.000 ;
        RECT 322.800 304.200 323.600 305.000 ;
        RECT 332.400 307.600 333.200 308.400 ;
        RECT 351.600 309.600 352.400 310.400 ;
        RECT 346.800 307.600 347.600 308.400 ;
        RECT 372.400 313.600 373.200 314.400 ;
        RECT 356.400 305.600 357.200 306.400 ;
        RECT 385.200 311.600 386.000 312.400 ;
        RECT 383.600 307.600 384.400 308.400 ;
        RECT 398.000 309.600 398.800 310.400 ;
        RECT 404.400 309.600 405.200 310.400 ;
        RECT 415.600 309.600 416.400 310.400 ;
        RECT 420.400 309.600 421.200 310.400 ;
        RECT 442.800 315.000 443.600 315.800 ;
        RECT 439.600 313.600 440.400 314.400 ;
        RECT 457.200 315.600 458.000 316.400 ;
        RECT 444.400 312.400 445.200 313.200 ;
        RECT 449.200 309.600 450.000 310.400 ;
        RECT 409.200 307.600 410.000 308.400 ;
        RECT 393.200 303.600 394.000 304.400 ;
        RECT 410.800 305.600 411.600 306.400 ;
        RECT 417.200 307.600 418.000 308.400 ;
        RECT 433.200 308.200 434.000 309.000 ;
        RECT 442.800 308.600 443.600 309.400 ;
        RECT 412.400 303.600 413.200 304.400 ;
        RECT 438.000 307.600 438.800 308.400 ;
        RECT 433.200 304.200 434.000 305.000 ;
        RECT 434.800 304.200 435.600 305.000 ;
        RECT 436.400 304.200 437.200 305.000 ;
        RECT 439.600 304.200 440.400 305.000 ;
        RECT 442.800 304.200 443.600 305.000 ;
        RECT 444.400 304.200 445.200 305.000 ;
        RECT 446.000 304.200 446.800 305.000 ;
        RECT 447.600 304.200 448.400 305.000 ;
        RECT 466.800 309.600 467.600 310.400 ;
        RECT 476.400 309.600 477.200 310.400 ;
        RECT 484.400 309.600 485.200 310.400 ;
        RECT 457.200 303.600 458.000 304.400 ;
        RECT 471.600 305.600 472.400 306.400 ;
        RECT 479.600 305.600 480.400 306.400 ;
        RECT 486.000 307.600 486.800 308.400 ;
        RECT 492.400 307.600 493.200 308.400 ;
        RECT 481.200 303.600 482.000 304.400 ;
        RECT 487.600 303.600 488.400 304.400 ;
        RECT 502.000 309.600 502.800 310.400 ;
        RECT 508.400 309.600 509.200 310.400 ;
        RECT 516.400 307.600 517.200 308.400 ;
        RECT 526.000 317.600 526.800 318.400 ;
        RECT 532.400 313.600 533.200 314.400 ;
        RECT 526.000 309.600 526.800 310.400 ;
        RECT 529.200 309.600 530.000 310.400 ;
        RECT 521.200 307.600 522.000 308.400 ;
        RECT 527.600 307.600 528.400 308.400 ;
        RECT 534.000 307.600 534.800 308.400 ;
        RECT 546.800 317.600 547.600 318.400 ;
        RECT 537.200 303.600 538.000 304.400 ;
        RECT 542.000 303.600 542.800 304.400 ;
        RECT 546.800 303.600 547.600 304.400 ;
        RECT 567.600 315.000 568.400 315.800 ;
        RECT 564.400 313.600 565.200 314.400 ;
        RECT 569.200 312.400 570.000 313.200 ;
        RECT 574.000 309.600 574.800 310.400 ;
        RECT 558.000 308.200 558.800 309.000 ;
        RECT 567.600 308.600 568.400 309.400 ;
        RECT 562.800 307.600 563.600 308.400 ;
        RECT 558.000 304.200 558.800 305.000 ;
        RECT 559.600 304.200 560.400 305.000 ;
        RECT 561.200 304.200 562.000 305.000 ;
        RECT 564.400 304.200 565.200 305.000 ;
        RECT 567.600 304.200 568.400 305.000 ;
        RECT 569.200 304.200 570.000 305.000 ;
        RECT 570.800 304.200 571.600 305.000 ;
        RECT 572.400 304.200 573.200 305.000 ;
        RECT 582.000 305.600 582.800 306.400 ;
        RECT 590.000 307.600 590.800 308.400 ;
        RECT 593.200 305.600 594.000 306.400 ;
        RECT 599.600 307.600 600.400 308.400 ;
        RECT 594.800 303.600 595.600 304.400 ;
        RECT 604.400 309.600 605.200 310.400 ;
        RECT 602.800 305.600 603.600 306.400 ;
        RECT 1.200 293.600 2.000 294.400 ;
        RECT 14.000 293.600 14.800 294.400 ;
        RECT 23.600 293.000 24.400 293.800 ;
        RECT 33.200 292.600 34.000 293.400 ;
        RECT 18.800 291.600 19.600 292.400 ;
        RECT 28.400 291.600 29.200 292.400 ;
        RECT 25.200 288.800 26.000 289.600 ;
        RECT 30.000 287.600 30.800 288.400 ;
        RECT 26.800 286.200 27.600 287.000 ;
        RECT 23.600 284.200 24.400 285.000 ;
        RECT 25.200 284.200 26.000 285.000 ;
        RECT 30.000 286.200 30.800 287.000 ;
        RECT 33.200 286.200 34.000 287.000 ;
        RECT 34.800 284.200 35.600 285.000 ;
        RECT 36.400 284.200 37.200 285.000 ;
        RECT 38.000 284.200 38.800 285.000 ;
        RECT 54.000 291.600 54.800 292.400 ;
        RECT 58.800 293.600 59.600 294.400 ;
        RECT 70.000 293.000 70.800 293.800 ;
        RECT 60.400 291.600 61.200 292.400 ;
        RECT 47.600 283.600 48.400 284.400 ;
        RECT 79.600 292.600 80.400 293.400 ;
        RECT 68.400 291.600 69.200 292.400 ;
        RECT 71.600 288.800 72.400 289.600 ;
        RECT 76.400 287.600 77.200 288.400 ;
        RECT 73.200 286.200 74.000 287.000 ;
        RECT 70.000 284.200 70.800 285.000 ;
        RECT 71.600 284.200 72.400 285.000 ;
        RECT 76.400 286.200 77.200 287.000 ;
        RECT 79.600 286.200 80.400 287.000 ;
        RECT 81.200 284.200 82.000 285.000 ;
        RECT 82.800 284.200 83.600 285.000 ;
        RECT 84.400 284.200 85.200 285.000 ;
        RECT 100.400 291.600 101.200 292.400 ;
        RECT 105.200 293.600 106.000 294.400 ;
        RECT 122.800 297.600 123.600 298.400 ;
        RECT 106.800 291.600 107.600 292.400 ;
        RECT 110.000 291.600 110.800 292.400 ;
        RECT 94.000 283.600 94.800 284.400 ;
        RECT 118.000 291.600 118.800 292.400 ;
        RECT 138.800 295.600 139.600 296.400 ;
        RECT 140.400 294.200 141.200 295.000 ;
        RECT 151.600 291.600 152.400 292.400 ;
        RECT 122.800 283.600 123.600 284.400 ;
        RECT 134.000 286.800 134.800 287.600 ;
        RECT 137.200 286.200 138.000 287.000 ;
        RECT 132.400 284.200 133.200 285.000 ;
        RECT 134.000 284.200 134.800 285.000 ;
        RECT 135.600 284.200 136.400 285.000 ;
        RECT 140.400 286.200 141.200 287.000 ;
        RECT 143.600 286.200 144.400 287.000 ;
        RECT 169.200 297.600 170.000 298.400 ;
        RECT 145.200 284.200 146.000 285.000 ;
        RECT 146.800 284.200 147.600 285.000 ;
        RECT 178.800 293.000 179.600 293.800 ;
        RECT 169.200 289.600 170.000 290.400 ;
        RECT 188.400 292.600 189.200 293.400 ;
        RECT 207.600 297.600 208.400 298.400 ;
        RECT 175.600 291.600 176.400 292.400 ;
        RECT 180.400 288.800 181.200 289.600 ;
        RECT 185.200 287.600 186.000 288.400 ;
        RECT 182.000 286.200 182.800 287.000 ;
        RECT 178.800 284.200 179.600 285.000 ;
        RECT 180.400 284.200 181.200 285.000 ;
        RECT 185.200 286.200 186.000 287.000 ;
        RECT 188.400 286.200 189.200 287.000 ;
        RECT 190.000 284.200 190.800 285.000 ;
        RECT 191.600 284.200 192.400 285.000 ;
        RECT 193.200 284.200 194.000 285.000 ;
        RECT 207.600 283.600 208.400 284.400 ;
        RECT 226.800 293.000 227.600 293.800 ;
        RECT 217.200 289.600 218.000 290.400 ;
        RECT 236.400 292.600 237.200 293.400 ;
        RECT 222.000 291.600 222.800 292.400 ;
        RECT 228.400 288.800 229.200 289.600 ;
        RECT 233.200 287.600 234.000 288.400 ;
        RECT 230.000 286.200 230.800 287.000 ;
        RECT 226.800 284.200 227.600 285.000 ;
        RECT 228.400 284.200 229.200 285.000 ;
        RECT 233.200 286.200 234.000 287.000 ;
        RECT 236.400 286.200 237.200 287.000 ;
        RECT 238.000 284.200 238.800 285.000 ;
        RECT 239.600 284.200 240.400 285.000 ;
        RECT 241.200 284.200 242.000 285.000 ;
        RECT 250.800 283.600 251.600 284.400 ;
        RECT 274.800 293.000 275.600 293.800 ;
        RECT 284.400 292.600 285.200 293.400 ;
        RECT 298.800 297.600 299.600 298.400 ;
        RECT 270.000 291.600 270.800 292.400 ;
        RECT 290.800 291.600 291.600 292.400 ;
        RECT 276.400 288.800 277.200 289.600 ;
        RECT 281.200 287.600 282.000 288.400 ;
        RECT 278.000 286.200 278.800 287.000 ;
        RECT 274.800 284.200 275.600 285.000 ;
        RECT 276.400 284.200 277.200 285.000 ;
        RECT 281.200 286.200 282.000 287.000 ;
        RECT 284.400 286.200 285.200 287.000 ;
        RECT 286.000 284.200 286.800 285.000 ;
        RECT 287.600 284.200 288.400 285.000 ;
        RECT 289.200 284.200 290.000 285.000 ;
        RECT 305.200 289.600 306.000 290.400 ;
        RECT 314.800 289.600 315.600 290.400 ;
        RECT 330.800 291.600 331.600 292.400 ;
        RECT 319.600 289.600 320.400 290.400 ;
        RECT 326.000 289.600 326.800 290.400 ;
        RECT 332.400 289.600 333.200 290.400 ;
        RECT 354.800 285.600 355.600 286.400 ;
        RECT 366.000 291.600 366.800 292.400 ;
        RECT 369.200 289.600 370.000 290.400 ;
        RECT 396.400 297.600 397.200 298.400 ;
        RECT 399.600 297.600 400.400 298.400 ;
        RECT 390.000 293.600 390.800 294.400 ;
        RECT 385.200 291.600 386.000 292.400 ;
        RECT 391.600 291.600 392.400 292.400 ;
        RECT 382.000 283.600 382.800 284.400 ;
        RECT 415.600 295.600 416.400 296.400 ;
        RECT 417.200 294.200 418.000 295.000 ;
        RECT 428.400 291.600 429.200 292.400 ;
        RECT 399.600 283.600 400.400 284.400 ;
        RECT 410.800 286.800 411.600 287.600 ;
        RECT 414.000 286.200 414.800 287.000 ;
        RECT 409.200 284.200 410.000 285.000 ;
        RECT 410.800 284.200 411.600 285.000 ;
        RECT 412.400 284.200 413.200 285.000 ;
        RECT 417.200 286.200 418.000 287.000 ;
        RECT 420.400 286.200 421.200 287.000 ;
        RECT 438.000 293.600 438.800 294.400 ;
        RECT 433.200 291.600 434.000 292.400 ;
        RECT 439.600 291.600 440.400 292.400 ;
        RECT 441.200 291.600 442.000 292.400 ;
        RECT 447.600 291.600 448.400 292.400 ;
        RECT 422.000 284.200 422.800 285.000 ;
        RECT 423.600 284.200 424.400 285.000 ;
        RECT 476.400 297.600 477.200 298.400 ;
        RECT 474.800 293.600 475.600 294.400 ;
        RECT 471.600 283.600 472.400 284.400 ;
        RECT 479.600 289.600 480.400 290.400 ;
        RECT 486.000 293.600 486.800 294.400 ;
        RECT 511.600 297.600 512.400 298.400 ;
        RECT 489.200 291.600 490.000 292.400 ;
        RECT 494.000 291.600 494.800 292.400 ;
        RECT 498.800 289.600 499.600 290.400 ;
        RECT 529.200 297.600 530.000 298.400 ;
        RECT 518.000 291.600 518.800 292.400 ;
        RECT 516.400 289.600 517.200 290.400 ;
        RECT 526.000 291.600 526.800 292.400 ;
        RECT 532.400 293.600 533.200 294.400 ;
        RECT 554.800 295.600 555.600 296.400 ;
        RECT 556.400 294.200 557.200 295.000 ;
        RECT 575.600 297.600 576.400 298.400 ;
        RECT 558.000 291.600 558.800 292.400 ;
        RECT 569.200 291.600 570.000 292.400 ;
        RECT 519.600 283.600 520.400 284.400 ;
        RECT 526.000 283.600 526.800 284.400 ;
        RECT 529.200 283.600 530.000 284.400 ;
        RECT 538.800 289.600 539.600 290.400 ;
        RECT 550.000 286.800 550.800 287.600 ;
        RECT 553.200 286.200 554.000 287.000 ;
        RECT 548.400 284.200 549.200 285.000 ;
        RECT 550.000 284.200 550.800 285.000 ;
        RECT 551.600 284.200 552.400 285.000 ;
        RECT 556.400 286.200 557.200 287.000 ;
        RECT 559.600 286.200 560.400 287.000 ;
        RECT 561.200 284.200 562.000 285.000 ;
        RECT 562.800 284.200 563.600 285.000 ;
        RECT 585.200 293.000 586.000 293.800 ;
        RECT 575.600 289.600 576.400 290.400 ;
        RECT 594.800 292.600 595.600 293.400 ;
        RECT 578.800 291.600 579.600 292.400 ;
        RECT 601.200 291.600 602.000 292.400 ;
        RECT 586.800 288.800 587.600 289.600 ;
        RECT 591.600 287.600 592.400 288.400 ;
        RECT 588.400 286.200 589.200 287.000 ;
        RECT 585.200 284.200 586.000 285.000 ;
        RECT 586.800 284.200 587.600 285.000 ;
        RECT 591.600 286.200 592.400 287.000 ;
        RECT 594.800 286.200 595.600 287.000 ;
        RECT 596.400 284.200 597.200 285.000 ;
        RECT 598.000 284.200 598.800 285.000 ;
        RECT 599.600 284.200 600.400 285.000 ;
        RECT 609.200 283.600 610.000 284.400 ;
        RECT 18.800 275.000 19.600 275.800 ;
        RECT 15.600 273.600 16.400 274.400 ;
        RECT 20.400 272.400 21.200 273.200 ;
        RECT 25.200 269.600 26.000 270.400 ;
        RECT 9.200 268.200 10.000 269.000 ;
        RECT 18.800 268.600 19.600 269.400 ;
        RECT 14.000 267.600 14.800 268.400 ;
        RECT 9.200 264.200 10.000 265.000 ;
        RECT 10.800 264.200 11.600 265.000 ;
        RECT 12.400 264.200 13.200 265.000 ;
        RECT 15.600 264.200 16.400 265.000 ;
        RECT 18.800 264.200 19.600 265.000 ;
        RECT 20.400 264.200 21.200 265.000 ;
        RECT 22.000 264.200 22.800 265.000 ;
        RECT 23.600 264.200 24.400 265.000 ;
        RECT 49.200 274.400 50.000 275.200 ;
        RECT 52.400 275.000 53.200 275.800 ;
        RECT 47.600 272.400 48.400 273.200 ;
        RECT 46.000 269.600 46.800 270.400 ;
        RECT 33.200 263.600 34.000 264.400 ;
        RECT 38.000 263.600 38.800 264.400 ;
        RECT 84.400 277.600 85.200 278.400 ;
        RECT 57.200 267.600 58.000 268.400 ;
        RECT 54.000 265.600 54.800 266.400 ;
        RECT 95.600 274.400 96.400 275.200 ;
        RECT 98.800 275.000 99.600 275.800 ;
        RECT 94.000 272.400 94.800 273.200 ;
        RECT 47.600 264.200 48.400 265.000 ;
        RECT 49.200 264.200 50.000 265.000 ;
        RECT 50.800 264.200 51.600 265.000 ;
        RECT 52.400 264.200 53.200 265.000 ;
        RECT 55.600 264.200 56.400 265.000 ;
        RECT 58.800 264.200 59.600 265.000 ;
        RECT 60.400 264.200 61.200 265.000 ;
        RECT 62.000 264.200 62.800 265.000 ;
        RECT 71.600 265.600 72.400 266.400 ;
        RECT 92.400 269.600 93.200 270.400 ;
        RECT 126.000 277.600 126.800 278.400 ;
        RECT 103.600 267.600 104.400 268.400 ;
        RECT 100.400 265.600 101.200 266.400 ;
        RECT 94.000 264.200 94.800 265.000 ;
        RECT 95.600 264.200 96.400 265.000 ;
        RECT 97.200 264.200 98.000 265.000 ;
        RECT 98.800 264.200 99.600 265.000 ;
        RECT 102.000 264.200 102.800 265.000 ;
        RECT 105.200 264.200 106.000 265.000 ;
        RECT 106.800 264.200 107.600 265.000 ;
        RECT 108.400 264.200 109.200 265.000 ;
        RECT 119.600 263.600 120.400 264.400 ;
        RECT 126.000 263.600 126.800 264.400 ;
        RECT 150.000 263.600 150.800 264.400 ;
        RECT 167.600 265.600 168.400 266.400 ;
        RECT 193.200 275.000 194.000 275.800 ;
        RECT 190.000 273.600 190.800 274.400 ;
        RECT 194.800 272.400 195.600 273.200 ;
        RECT 199.600 269.600 200.400 270.400 ;
        RECT 183.600 268.200 184.400 269.000 ;
        RECT 193.200 268.600 194.000 269.400 ;
        RECT 174.000 265.600 174.800 266.400 ;
        RECT 188.400 267.600 189.200 268.400 ;
        RECT 207.800 267.600 208.600 268.400 ;
        RECT 183.600 264.200 184.400 265.000 ;
        RECT 185.200 264.200 186.000 265.000 ;
        RECT 186.800 264.200 187.600 265.000 ;
        RECT 190.000 264.200 190.800 265.000 ;
        RECT 193.200 264.200 194.000 265.000 ;
        RECT 194.800 264.200 195.600 265.000 ;
        RECT 196.400 264.200 197.200 265.000 ;
        RECT 198.000 264.200 198.800 265.000 ;
        RECT 212.400 267.600 213.200 268.400 ;
        RECT 228.400 277.600 229.200 278.400 ;
        RECT 249.200 275.000 250.000 275.800 ;
        RECT 246.000 273.600 246.800 274.400 ;
        RECT 250.800 272.400 251.600 273.200 ;
        RECT 255.600 269.600 256.400 270.400 ;
        RECT 239.600 268.200 240.400 269.000 ;
        RECT 249.200 268.600 250.000 269.400 ;
        RECT 225.200 263.600 226.000 264.400 ;
        RECT 244.400 267.600 245.200 268.400 ;
        RECT 239.600 264.200 240.400 265.000 ;
        RECT 241.200 264.200 242.000 265.000 ;
        RECT 242.800 264.200 243.600 265.000 ;
        RECT 246.000 264.200 246.800 265.000 ;
        RECT 249.200 264.200 250.000 265.000 ;
        RECT 250.800 264.200 251.600 265.000 ;
        RECT 252.400 264.200 253.200 265.000 ;
        RECT 254.000 264.200 254.800 265.000 ;
        RECT 266.800 269.600 267.600 270.400 ;
        RECT 268.400 269.600 269.200 270.400 ;
        RECT 294.000 277.600 294.800 278.400 ;
        RECT 263.600 265.600 264.400 266.400 ;
        RECT 287.600 269.600 288.400 270.400 ;
        RECT 278.000 265.600 278.800 266.400 ;
        RECT 284.400 267.600 285.200 268.400 ;
        RECT 292.400 265.600 293.200 266.400 ;
        RECT 295.600 269.600 296.400 270.400 ;
        RECT 297.200 269.600 298.000 270.400 ;
        RECT 327.600 275.000 328.400 275.800 ;
        RECT 324.400 273.600 325.200 274.400 ;
        RECT 329.200 272.400 330.000 273.200 ;
        RECT 318.000 268.200 318.800 269.000 ;
        RECT 327.600 268.600 328.400 269.400 ;
        RECT 322.800 267.600 323.600 268.400 ;
        RECT 318.000 264.200 318.800 265.000 ;
        RECT 319.600 264.200 320.400 265.000 ;
        RECT 321.200 264.200 322.000 265.000 ;
        RECT 324.400 264.200 325.200 265.000 ;
        RECT 327.600 264.200 328.400 265.000 ;
        RECT 329.200 264.200 330.000 265.000 ;
        RECT 330.800 264.200 331.600 265.000 ;
        RECT 332.400 264.200 333.200 265.000 ;
        RECT 342.000 263.600 342.800 264.400 ;
        RECT 351.600 269.600 352.400 270.400 ;
        RECT 346.800 265.600 347.600 266.400 ;
        RECT 353.200 267.600 354.000 268.400 ;
        RECT 362.800 265.600 363.600 266.400 ;
        RECT 380.400 277.600 381.200 278.400 ;
        RECT 383.600 277.600 384.400 278.400 ;
        RECT 390.000 277.600 390.800 278.400 ;
        RECT 372.400 273.600 373.200 274.400 ;
        RECT 378.800 273.600 379.600 274.400 ;
        RECT 385.200 273.600 386.000 274.400 ;
        RECT 391.600 273.600 392.400 274.400 ;
        RECT 369.200 271.600 370.000 272.400 ;
        RECT 375.600 271.600 376.400 272.400 ;
        RECT 382.000 271.600 382.800 272.400 ;
        RECT 399.600 275.600 400.400 276.400 ;
        RECT 407.600 273.600 408.400 274.400 ;
        RECT 367.600 267.600 368.400 268.400 ;
        RECT 366.000 263.600 366.800 264.400 ;
        RECT 410.800 267.600 411.600 268.400 ;
        RECT 417.200 273.600 418.000 274.400 ;
        RECT 433.200 277.600 434.000 278.400 ;
        RECT 434.800 273.600 435.600 274.400 ;
        RECT 441.200 277.600 442.000 278.400 ;
        RECT 439.600 273.600 440.400 274.400 ;
        RECT 431.600 271.600 432.400 272.400 ;
        RECT 442.800 271.600 443.600 272.400 ;
        RECT 452.400 277.600 453.200 278.400 ;
        RECT 474.800 277.600 475.600 278.400 ;
        RECT 466.800 273.600 467.600 274.400 ;
        RECT 479.600 273.600 480.400 274.400 ;
        RECT 492.400 277.600 493.200 278.400 ;
        RECT 441.200 269.600 442.000 270.400 ;
        RECT 463.600 271.600 464.400 272.400 ;
        RECT 476.400 271.600 477.200 272.400 ;
        RECT 500.400 275.600 501.200 276.400 ;
        RECT 505.200 277.600 506.000 278.400 ;
        RECT 510.000 273.600 510.800 274.400 ;
        RECT 489.200 269.600 490.000 270.400 ;
        RECT 492.400 269.600 493.200 270.400 ;
        RECT 486.000 265.600 486.800 266.400 ;
        RECT 494.000 267.600 494.800 268.400 ;
        RECT 484.400 263.600 485.200 264.400 ;
        RECT 502.000 265.600 502.800 266.400 ;
        RECT 511.600 267.600 512.400 268.400 ;
        RECT 530.800 269.600 531.600 270.400 ;
        RECT 534.000 269.600 534.800 270.400 ;
        RECT 513.200 265.600 514.000 266.400 ;
        RECT 521.200 265.600 522.000 266.400 ;
        RECT 540.400 267.600 541.200 268.400 ;
        RECT 543.600 265.600 544.400 266.400 ;
        RECT 548.400 267.600 549.200 268.400 ;
        RECT 556.400 269.600 557.200 270.400 ;
        RECT 567.600 269.600 568.400 270.400 ;
        RECT 578.800 275.600 579.600 276.400 ;
        RECT 590.000 274.400 590.800 275.200 ;
        RECT 593.200 275.000 594.000 275.800 ;
        RECT 588.400 272.400 589.200 273.200 ;
        RECT 586.800 269.600 587.600 270.400 ;
        RECT 538.800 263.600 539.600 264.400 ;
        RECT 542.000 263.600 542.800 264.400 ;
        RECT 551.600 263.600 552.400 264.400 ;
        RECT 564.400 263.600 565.200 264.400 ;
        RECT 598.000 267.600 598.800 268.400 ;
        RECT 594.800 265.600 595.600 266.400 ;
        RECT 588.400 264.200 589.200 265.000 ;
        RECT 590.000 264.200 590.800 265.000 ;
        RECT 591.600 264.200 592.400 265.000 ;
        RECT 593.200 264.200 594.000 265.000 ;
        RECT 596.400 264.200 597.200 265.000 ;
        RECT 599.600 264.200 600.400 265.000 ;
        RECT 601.200 264.200 602.000 265.000 ;
        RECT 602.800 264.200 603.600 265.000 ;
        RECT 9.200 253.000 10.000 253.800 ;
        RECT 18.800 252.600 19.600 253.400 ;
        RECT 25.200 251.600 26.000 252.400 ;
        RECT 10.800 248.800 11.600 249.600 ;
        RECT 15.600 247.600 16.400 248.400 ;
        RECT 12.400 246.200 13.200 247.000 ;
        RECT 9.200 244.200 10.000 245.000 ;
        RECT 10.800 244.200 11.600 245.000 ;
        RECT 15.600 246.200 16.400 247.000 ;
        RECT 18.800 246.200 19.600 247.000 ;
        RECT 20.400 244.200 21.200 245.000 ;
        RECT 22.000 244.200 22.800 245.000 ;
        RECT 23.600 244.200 24.400 245.000 ;
        RECT 33.200 243.600 34.000 244.400 ;
        RECT 47.600 253.000 48.400 253.800 ;
        RECT 57.200 252.600 58.000 253.400 ;
        RECT 81.200 257.600 82.000 258.400 ;
        RECT 41.200 251.600 42.000 252.400 ;
        RECT 63.600 251.600 64.400 252.400 ;
        RECT 49.200 248.800 50.000 249.600 ;
        RECT 54.000 247.600 54.800 248.400 ;
        RECT 50.800 246.200 51.600 247.000 ;
        RECT 47.600 244.200 48.400 245.000 ;
        RECT 49.200 244.200 50.000 245.000 ;
        RECT 54.000 246.200 54.800 247.000 ;
        RECT 57.200 246.200 58.000 247.000 ;
        RECT 58.800 244.200 59.600 245.000 ;
        RECT 60.400 244.200 61.200 245.000 ;
        RECT 62.000 244.200 62.800 245.000 ;
        RECT 78.000 251.600 78.800 252.400 ;
        RECT 82.800 253.600 83.600 254.400 ;
        RECT 84.400 251.600 85.200 252.400 ;
        RECT 71.600 243.600 72.400 244.400 ;
        RECT 111.600 255.600 112.400 256.400 ;
        RECT 113.200 254.200 114.000 255.000 ;
        RECT 124.400 251.600 125.200 252.400 ;
        RECT 86.000 243.600 86.800 244.400 ;
        RECT 95.600 243.600 96.400 244.400 ;
        RECT 106.800 246.800 107.600 247.600 ;
        RECT 110.000 246.200 110.800 247.000 ;
        RECT 105.200 244.200 106.000 245.000 ;
        RECT 106.800 244.200 107.600 245.000 ;
        RECT 108.400 244.200 109.200 245.000 ;
        RECT 113.200 246.200 114.000 247.000 ;
        RECT 116.400 246.200 117.200 247.000 ;
        RECT 118.000 244.200 118.800 245.000 ;
        RECT 119.600 244.200 120.400 245.000 ;
        RECT 137.200 251.600 138.000 252.400 ;
        RECT 161.200 255.600 162.000 256.400 ;
        RECT 162.800 254.200 163.600 255.000 ;
        RECT 174.000 251.600 174.800 252.400 ;
        RECT 129.200 243.600 130.000 244.400 ;
        RECT 145.200 243.600 146.000 244.400 ;
        RECT 156.400 246.800 157.200 247.600 ;
        RECT 159.600 246.200 160.400 247.000 ;
        RECT 154.800 244.200 155.600 245.000 ;
        RECT 156.400 244.200 157.200 245.000 ;
        RECT 158.000 244.200 158.800 245.000 ;
        RECT 162.800 246.200 163.600 247.000 ;
        RECT 166.000 246.200 166.800 247.000 ;
        RECT 167.600 244.200 168.400 245.000 ;
        RECT 169.200 244.200 170.000 245.000 ;
        RECT 182.000 249.600 182.800 250.400 ;
        RECT 202.800 253.000 203.600 253.800 ;
        RECT 212.400 252.600 213.200 253.400 ;
        RECT 199.600 251.600 200.400 252.400 ;
        RECT 204.400 248.800 205.200 249.600 ;
        RECT 209.200 247.600 210.000 248.400 ;
        RECT 206.000 246.200 206.800 247.000 ;
        RECT 202.800 244.200 203.600 245.000 ;
        RECT 204.400 244.200 205.200 245.000 ;
        RECT 209.200 246.200 210.000 247.000 ;
        RECT 212.400 246.200 213.200 247.000 ;
        RECT 214.000 244.200 214.800 245.000 ;
        RECT 215.600 244.200 216.400 245.000 ;
        RECT 217.200 244.200 218.000 245.000 ;
        RECT 226.800 243.600 227.600 244.400 ;
        RECT 247.600 251.600 248.400 252.400 ;
        RECT 266.800 255.600 267.600 256.400 ;
        RECT 268.400 254.200 269.200 255.000 ;
        RECT 286.000 257.600 286.800 258.400 ;
        RECT 258.800 251.600 259.600 252.400 ;
        RECT 244.400 243.600 245.200 244.400 ;
        RECT 250.800 243.600 251.600 244.400 ;
        RECT 262.000 246.800 262.800 247.600 ;
        RECT 265.200 246.200 266.000 247.000 ;
        RECT 260.400 244.200 261.200 245.000 ;
        RECT 262.000 244.200 262.800 245.000 ;
        RECT 263.600 244.200 264.400 245.000 ;
        RECT 268.400 246.200 269.200 247.000 ;
        RECT 271.600 246.200 272.400 247.000 ;
        RECT 284.400 253.600 285.200 254.400 ;
        RECT 273.200 244.200 274.000 245.000 ;
        RECT 274.800 244.200 275.600 245.000 ;
        RECT 302.000 249.600 302.800 250.400 ;
        RECT 319.600 251.600 320.400 252.400 ;
        RECT 327.600 253.600 328.400 254.400 ;
        RECT 350.000 255.600 350.800 256.400 ;
        RECT 313.200 243.600 314.000 244.400 ;
        RECT 316.400 243.600 317.200 244.400 ;
        RECT 324.400 247.600 325.200 248.400 ;
        RECT 335.600 249.600 336.400 250.400 ;
        RECT 342.000 243.600 342.800 244.400 ;
        RECT 359.600 253.000 360.400 253.800 ;
        RECT 369.200 252.600 370.000 253.400 ;
        RECT 386.800 257.600 387.600 258.400 ;
        RECT 356.400 251.600 357.200 252.400 ;
        RECT 361.200 248.800 362.000 249.600 ;
        RECT 366.000 247.600 366.800 248.400 ;
        RECT 362.800 246.200 363.600 247.000 ;
        RECT 359.600 244.200 360.400 245.000 ;
        RECT 361.200 244.200 362.000 245.000 ;
        RECT 366.000 246.200 366.800 247.000 ;
        RECT 369.200 246.200 370.000 247.000 ;
        RECT 370.800 244.200 371.600 245.000 ;
        RECT 372.400 244.200 373.200 245.000 ;
        RECT 374.000 244.200 374.800 245.000 ;
        RECT 383.600 243.600 384.400 244.400 ;
        RECT 401.200 253.600 402.000 254.400 ;
        RECT 409.200 253.600 410.000 254.400 ;
        RECT 396.400 251.600 397.200 252.400 ;
        RECT 402.800 251.600 403.600 252.400 ;
        RECT 404.400 251.600 405.200 252.400 ;
        RECT 410.800 251.600 411.600 252.400 ;
        RECT 433.200 257.600 434.000 258.400 ;
        RECT 391.600 245.600 392.400 246.400 ;
        RECT 414.000 249.600 414.800 250.400 ;
        RECT 415.600 249.600 416.400 250.400 ;
        RECT 423.600 249.600 424.400 250.400 ;
        RECT 430.000 253.600 430.800 254.400 ;
        RECT 434.800 251.600 435.600 252.400 ;
        RECT 439.600 249.600 440.400 250.400 ;
        RECT 441.200 249.600 442.000 250.400 ;
        RECT 455.600 257.600 456.400 258.400 ;
        RECT 468.400 257.600 469.200 258.400 ;
        RECT 478.000 257.600 478.800 258.400 ;
        RECT 457.200 253.600 458.000 254.400 ;
        RECT 470.000 253.600 470.800 254.400 ;
        RECT 452.400 251.600 453.200 252.400 ;
        RECT 458.800 251.600 459.600 252.400 ;
        RECT 465.200 251.600 466.000 252.400 ;
        RECT 471.600 251.600 472.400 252.400 ;
        RECT 492.400 257.600 493.200 258.400 ;
        RECT 489.200 255.600 490.000 256.400 ;
        RECT 482.800 251.600 483.600 252.400 ;
        RECT 484.400 251.600 485.200 252.400 ;
        RECT 497.200 253.600 498.000 254.400 ;
        RECT 502.000 249.600 502.800 250.400 ;
        RECT 519.600 257.600 520.400 258.400 ;
        RECT 527.600 257.600 528.400 258.400 ;
        RECT 518.000 253.600 518.800 254.400 ;
        RECT 526.000 253.600 526.800 254.400 ;
        RECT 546.800 257.600 547.600 258.400 ;
        RECT 510.000 251.600 510.800 252.400 ;
        RECT 513.200 251.600 514.000 252.400 ;
        RECT 503.600 243.600 504.400 244.400 ;
        RECT 506.800 243.600 507.600 244.400 ;
        RECT 570.800 257.600 571.600 258.400 ;
        RECT 554.800 253.600 555.600 254.400 ;
        RECT 586.800 255.600 587.600 256.400 ;
        RECT 588.400 254.200 589.200 255.000 ;
        RECT 578.800 251.600 579.600 252.400 ;
        RECT 553.200 249.600 554.000 250.400 ;
        RECT 566.000 243.600 566.800 244.400 ;
        RECT 582.000 246.800 582.800 247.600 ;
        RECT 585.200 246.200 586.000 247.000 ;
        RECT 580.400 244.200 581.200 245.000 ;
        RECT 582.000 244.200 582.800 245.000 ;
        RECT 583.600 244.200 584.400 245.000 ;
        RECT 588.400 246.200 589.200 247.000 ;
        RECT 591.600 246.200 592.400 247.000 ;
        RECT 593.200 244.200 594.000 245.000 ;
        RECT 594.800 244.200 595.600 245.000 ;
        RECT 2.800 227.600 3.600 228.400 ;
        RECT 9.200 229.600 10.000 230.400 ;
        RECT 15.600 229.600 16.400 230.400 ;
        RECT 22.000 229.600 22.800 230.400 ;
        RECT 6.000 225.600 6.800 226.400 ;
        RECT 26.800 227.600 27.600 228.400 ;
        RECT 30.000 233.600 30.800 234.400 ;
        RECT 33.200 229.600 34.000 230.400 ;
        RECT 42.800 227.600 43.600 228.400 ;
        RECT 39.600 225.600 40.400 226.400 ;
        RECT 41.200 225.600 42.000 226.400 ;
        RECT 38.000 223.600 38.800 224.400 ;
        RECT 62.000 235.000 62.800 235.800 ;
        RECT 58.800 233.600 59.600 234.400 ;
        RECT 63.600 232.400 64.400 233.200 ;
        RECT 68.400 229.600 69.200 230.400 ;
        RECT 52.400 228.200 53.200 229.000 ;
        RECT 62.000 228.600 62.800 229.400 ;
        RECT 57.200 227.600 58.000 228.400 ;
        RECT 76.600 229.600 77.400 230.400 ;
        RECT 52.400 224.200 53.200 225.000 ;
        RECT 54.000 224.200 54.800 225.000 ;
        RECT 55.600 224.200 56.400 225.000 ;
        RECT 58.800 224.200 59.600 225.000 ;
        RECT 62.000 224.200 62.800 225.000 ;
        RECT 63.600 224.200 64.400 225.000 ;
        RECT 65.200 224.200 66.000 225.000 ;
        RECT 66.800 224.200 67.600 225.000 ;
        RECT 82.800 227.600 83.600 228.400 ;
        RECT 127.600 231.600 128.400 232.400 ;
        RECT 106.800 227.600 107.600 228.400 ;
        RECT 95.600 223.600 96.400 224.400 ;
        RECT 105.200 226.200 106.000 227.000 ;
        RECT 122.800 223.600 123.600 224.400 ;
        RECT 138.800 227.600 139.600 228.400 ;
        RECT 132.400 223.600 133.200 224.400 ;
        RECT 167.600 235.000 168.400 235.800 ;
        RECT 164.400 233.600 165.200 234.400 ;
        RECT 182.000 237.600 182.800 238.400 ;
        RECT 169.200 232.400 170.000 233.200 ;
        RECT 186.800 237.600 187.600 238.400 ;
        RECT 174.000 229.600 174.800 230.400 ;
        RECT 158.000 228.200 158.800 229.000 ;
        RECT 167.600 228.600 168.400 229.400 ;
        RECT 143.600 225.600 144.400 226.400 ;
        RECT 162.800 227.600 163.600 228.400 ;
        RECT 158.000 224.200 158.800 225.000 ;
        RECT 159.600 224.200 160.400 225.000 ;
        RECT 161.200 224.200 162.000 225.000 ;
        RECT 164.400 224.200 165.200 225.000 ;
        RECT 167.600 224.200 168.400 225.000 ;
        RECT 169.200 224.200 170.000 225.000 ;
        RECT 170.800 224.200 171.600 225.000 ;
        RECT 172.400 224.200 173.200 225.000 ;
        RECT 185.200 225.600 186.000 226.400 ;
        RECT 206.000 235.000 206.800 235.800 ;
        RECT 202.800 233.600 203.600 234.400 ;
        RECT 220.400 237.600 221.200 238.400 ;
        RECT 207.600 232.400 208.400 233.200 ;
        RECT 212.400 229.600 213.200 230.400 ;
        RECT 196.400 228.200 197.200 229.000 ;
        RECT 206.000 228.600 206.800 229.400 ;
        RECT 201.200 227.600 202.000 228.400 ;
        RECT 196.400 224.200 197.200 225.000 ;
        RECT 198.000 224.200 198.800 225.000 ;
        RECT 199.600 224.200 200.400 225.000 ;
        RECT 202.800 224.200 203.600 225.000 ;
        RECT 206.000 224.200 206.800 225.000 ;
        RECT 207.600 224.200 208.400 225.000 ;
        RECT 209.200 224.200 210.000 225.000 ;
        RECT 210.800 224.200 211.600 225.000 ;
        RECT 249.200 235.000 250.000 235.800 ;
        RECT 246.000 233.600 246.800 234.400 ;
        RECT 250.800 232.400 251.600 233.200 ;
        RECT 255.600 229.600 256.400 230.400 ;
        RECT 239.600 228.200 240.400 229.000 ;
        RECT 249.200 228.600 250.000 229.400 ;
        RECT 220.400 223.600 221.200 224.400 ;
        RECT 225.200 225.600 226.000 226.400 ;
        RECT 244.400 227.600 245.200 228.400 ;
        RECT 263.800 227.600 264.600 228.400 ;
        RECT 239.600 224.200 240.400 225.000 ;
        RECT 241.200 224.200 242.000 225.000 ;
        RECT 242.800 224.200 243.600 225.000 ;
        RECT 246.000 224.200 246.800 225.000 ;
        RECT 249.200 224.200 250.000 225.000 ;
        RECT 250.800 224.200 251.600 225.000 ;
        RECT 252.400 224.200 253.200 225.000 ;
        RECT 254.000 224.200 254.800 225.000 ;
        RECT 286.000 237.600 286.800 238.400 ;
        RECT 274.800 227.600 275.600 228.400 ;
        RECT 282.800 229.600 283.600 230.400 ;
        RECT 284.400 227.600 285.200 228.400 ;
        RECT 279.600 223.600 280.400 224.400 ;
        RECT 297.200 229.600 298.000 230.400 ;
        RECT 319.600 237.600 320.400 238.400 ;
        RECT 326.000 237.600 326.800 238.400 ;
        RECT 321.200 233.600 322.000 234.400 ;
        RECT 318.000 231.600 318.800 232.400 ;
        RECT 340.400 237.600 341.200 238.400 ;
        RECT 342.000 233.600 342.800 234.400 ;
        RECT 348.400 233.600 349.200 234.400 ;
        RECT 287.600 225.600 288.400 226.400 ;
        RECT 294.000 227.600 294.800 228.400 ;
        RECT 302.000 227.600 302.800 228.400 ;
        RECT 303.600 227.600 304.400 228.400 ;
        RECT 338.800 231.600 339.600 232.400 ;
        RECT 351.600 231.600 352.400 232.400 ;
        RECT 358.000 229.600 358.800 230.400 ;
        RECT 359.600 229.600 360.400 230.400 ;
        RECT 326.000 223.600 326.800 224.400 ;
        RECT 385.200 235.000 386.000 235.800 ;
        RECT 382.000 233.600 382.800 234.400 ;
        RECT 386.800 232.400 387.600 233.200 ;
        RECT 399.600 233.600 400.400 234.400 ;
        RECT 375.600 228.200 376.400 229.000 ;
        RECT 385.200 228.600 386.000 229.400 ;
        RECT 380.400 227.600 381.200 228.400 ;
        RECT 375.600 224.200 376.400 225.000 ;
        RECT 377.200 224.200 378.000 225.000 ;
        RECT 378.800 224.200 379.600 225.000 ;
        RECT 382.000 224.200 382.800 225.000 ;
        RECT 385.200 224.200 386.000 225.000 ;
        RECT 386.800 224.200 387.600 225.000 ;
        RECT 388.400 224.200 389.200 225.000 ;
        RECT 390.000 224.200 390.800 225.000 ;
        RECT 407.600 231.600 408.400 232.400 ;
        RECT 418.800 237.600 419.600 238.400 ;
        RECT 404.400 225.600 405.200 226.400 ;
        RECT 409.200 227.600 410.000 228.400 ;
        RECT 473.200 237.600 474.000 238.400 ;
        RECT 474.800 233.600 475.600 234.400 ;
        RECT 471.600 231.600 472.400 232.400 ;
        RECT 466.800 227.600 467.600 228.400 ;
        RECT 442.800 223.600 443.600 224.400 ;
        RECT 478.000 227.600 478.800 228.400 ;
        RECT 487.600 233.600 488.400 234.400 ;
        RECT 490.800 237.600 491.600 238.400 ;
        RECT 492.400 233.600 493.200 234.400 ;
        RECT 495.600 231.600 496.400 232.400 ;
        RECT 513.200 237.600 514.000 238.400 ;
        RECT 524.400 237.600 525.200 238.400 ;
        RECT 535.600 237.600 536.400 238.400 ;
        RECT 511.600 233.600 512.400 234.400 ;
        RECT 519.600 233.600 520.400 234.400 ;
        RECT 526.000 233.600 526.800 234.400 ;
        RECT 537.200 233.600 538.000 234.400 ;
        RECT 543.600 233.600 544.400 234.400 ;
        RECT 494.000 229.600 494.800 230.400 ;
        RECT 508.400 231.600 509.200 232.400 ;
        RECT 506.800 229.600 507.600 230.400 ;
        RECT 514.800 231.600 515.600 232.400 ;
        RECT 522.800 231.600 523.600 232.400 ;
        RECT 513.200 229.600 514.000 230.400 ;
        RECT 529.200 231.600 530.000 232.400 ;
        RECT 540.400 231.600 541.200 232.400 ;
        RECT 546.800 231.600 547.600 232.400 ;
        RECT 538.800 229.600 539.600 230.400 ;
        RECT 545.200 229.600 546.000 230.400 ;
        RECT 554.800 237.600 555.600 238.400 ;
        RECT 558.000 237.600 558.800 238.400 ;
        RECT 559.600 233.600 560.400 234.400 ;
        RECT 551.600 227.600 552.400 228.400 ;
        RECT 553.200 227.600 554.000 228.400 ;
        RECT 580.400 234.400 581.200 235.200 ;
        RECT 583.600 235.000 584.400 235.800 ;
        RECT 578.800 232.400 579.600 233.200 ;
        RECT 566.000 227.600 566.800 228.400 ;
        RECT 577.200 229.600 578.000 230.400 ;
        RECT 569.200 223.600 570.000 224.400 ;
        RECT 588.400 227.600 589.200 228.400 ;
        RECT 585.200 225.600 586.000 226.400 ;
        RECT 604.400 229.600 605.200 230.400 ;
        RECT 578.800 224.200 579.600 225.000 ;
        RECT 580.400 224.200 581.200 225.000 ;
        RECT 582.000 224.200 582.800 225.000 ;
        RECT 583.600 224.200 584.400 225.000 ;
        RECT 586.800 224.200 587.600 225.000 ;
        RECT 590.000 224.200 590.800 225.000 ;
        RECT 591.600 224.200 592.400 225.000 ;
        RECT 593.200 224.200 594.000 225.000 ;
        RECT 14.000 213.600 14.800 214.400 ;
        RECT 9.200 209.600 10.000 210.400 ;
        RECT 22.000 209.600 22.800 210.400 ;
        RECT 66.800 217.600 67.600 218.400 ;
        RECT 74.800 215.600 75.600 216.400 ;
        RECT 26.800 209.600 27.600 210.400 ;
        RECT 25.200 207.600 26.000 208.400 ;
        RECT 55.600 213.600 56.400 214.400 ;
        RECT 116.400 217.600 117.200 218.400 ;
        RECT 38.000 203.600 38.800 204.400 ;
        RECT 71.600 211.600 72.400 212.400 ;
        RECT 102.000 213.600 102.800 214.400 ;
        RECT 84.400 212.200 85.200 213.000 ;
        RECT 92.400 211.800 93.200 212.600 ;
        RECT 97.200 210.200 98.000 211.000 ;
        RECT 79.600 207.600 80.400 208.400 ;
        RECT 172.400 217.600 173.200 218.400 ;
        RECT 142.000 212.200 142.800 213.000 ;
        RECT 129.200 209.600 130.000 210.400 ;
        RECT 134.000 209.600 134.800 210.400 ;
        RECT 154.800 210.200 155.600 211.000 ;
        RECT 172.400 214.800 173.200 215.600 ;
        RECT 175.600 213.600 176.400 214.400 ;
        RECT 164.400 211.600 165.200 212.400 ;
        RECT 194.800 215.600 195.600 216.400 ;
        RECT 196.400 214.200 197.200 215.000 ;
        RECT 204.400 211.600 205.200 212.400 ;
        RECT 137.200 207.600 138.000 208.400 ;
        RECT 178.800 203.600 179.600 204.400 ;
        RECT 190.000 206.800 190.800 207.600 ;
        RECT 193.200 206.200 194.000 207.000 ;
        RECT 188.400 204.200 189.200 205.000 ;
        RECT 190.000 204.200 190.800 205.000 ;
        RECT 191.600 204.200 192.400 205.000 ;
        RECT 196.400 206.200 197.200 207.000 ;
        RECT 199.600 206.200 200.400 207.000 ;
        RECT 220.400 213.000 221.200 213.800 ;
        RECT 230.000 212.600 230.800 213.400 ;
        RECT 244.400 217.600 245.200 218.400 ;
        RECT 249.200 217.600 250.000 218.400 ;
        RECT 215.600 211.600 216.400 212.400 ;
        RECT 222.000 208.800 222.800 209.600 ;
        RECT 226.800 207.600 227.600 208.400 ;
        RECT 201.200 204.200 202.000 205.000 ;
        RECT 202.800 204.200 203.600 205.000 ;
        RECT 223.600 206.200 224.400 207.000 ;
        RECT 220.400 204.200 221.200 205.000 ;
        RECT 222.000 204.200 222.800 205.000 ;
        RECT 226.800 206.200 227.600 207.000 ;
        RECT 230.000 206.200 230.800 207.000 ;
        RECT 231.600 204.200 232.400 205.000 ;
        RECT 233.200 204.200 234.000 205.000 ;
        RECT 234.800 204.200 235.600 205.000 ;
        RECT 244.400 203.600 245.200 204.400 ;
        RECT 258.800 213.000 259.600 213.800 ;
        RECT 268.400 212.600 269.200 213.400 ;
        RECT 255.600 211.600 256.400 212.400 ;
        RECT 274.800 211.600 275.600 212.400 ;
        RECT 260.400 208.800 261.200 209.600 ;
        RECT 265.200 207.600 266.000 208.400 ;
        RECT 262.000 206.200 262.800 207.000 ;
        RECT 258.800 204.200 259.600 205.000 ;
        RECT 260.400 204.200 261.200 205.000 ;
        RECT 265.200 206.200 266.000 207.000 ;
        RECT 268.400 206.200 269.200 207.000 ;
        RECT 270.000 204.200 270.800 205.000 ;
        RECT 271.600 204.200 272.400 205.000 ;
        RECT 273.200 204.200 274.000 205.000 ;
        RECT 282.800 205.600 283.600 206.400 ;
        RECT 310.000 217.600 310.800 218.400 ;
        RECT 302.000 213.600 302.800 214.400 ;
        RECT 290.800 203.600 291.600 204.400 ;
        RECT 326.000 215.600 326.800 216.400 ;
        RECT 327.600 214.200 328.400 215.000 ;
        RECT 351.600 217.600 352.400 218.400 ;
        RECT 318.000 211.600 318.800 212.400 ;
        RECT 340.400 211.600 341.200 212.400 ;
        RECT 310.000 203.600 310.800 204.400 ;
        RECT 321.200 206.800 322.000 207.600 ;
        RECT 324.400 206.200 325.200 207.000 ;
        RECT 319.600 204.200 320.400 205.000 ;
        RECT 321.200 204.200 322.000 205.000 ;
        RECT 322.800 204.200 323.600 205.000 ;
        RECT 327.600 206.200 328.400 207.000 ;
        RECT 330.800 206.200 331.600 207.000 ;
        RECT 367.600 215.600 368.400 216.400 ;
        RECT 369.200 214.200 370.000 215.000 ;
        RECT 386.800 215.600 387.600 216.400 ;
        RECT 378.800 211.600 379.600 212.400 ;
        RECT 332.400 204.200 333.200 205.000 ;
        RECT 334.000 204.200 334.800 205.000 ;
        RECT 362.800 206.800 363.600 207.600 ;
        RECT 366.000 206.200 366.800 207.000 ;
        RECT 361.200 204.200 362.000 205.000 ;
        RECT 362.800 204.200 363.600 205.000 ;
        RECT 364.400 204.200 365.200 205.000 ;
        RECT 369.200 206.200 370.000 207.000 ;
        RECT 372.400 206.200 373.200 207.000 ;
        RECT 374.000 204.200 374.800 205.000 ;
        RECT 375.600 204.200 376.400 205.000 ;
        RECT 401.200 217.600 402.000 218.400 ;
        RECT 388.400 209.600 389.200 210.400 ;
        RECT 391.600 203.600 392.400 204.400 ;
        RECT 412.400 203.600 413.200 204.400 ;
        RECT 417.200 203.600 418.000 204.400 ;
        RECT 442.800 215.600 443.600 216.400 ;
        RECT 444.400 214.200 445.200 215.000 ;
        RECT 434.800 211.600 435.600 212.400 ;
        RECT 423.600 209.600 424.400 210.400 ;
        RECT 426.800 209.600 427.600 210.400 ;
        RECT 438.000 206.800 438.800 207.600 ;
        RECT 441.200 206.200 442.000 207.000 ;
        RECT 436.400 204.200 437.200 205.000 ;
        RECT 438.000 204.200 438.800 205.000 ;
        RECT 439.600 204.200 440.400 205.000 ;
        RECT 444.400 206.200 445.200 207.000 ;
        RECT 447.600 206.200 448.400 207.000 ;
        RECT 449.200 204.200 450.000 205.000 ;
        RECT 450.800 204.200 451.600 205.000 ;
        RECT 466.800 203.600 467.600 204.400 ;
        RECT 470.000 203.600 470.800 204.400 ;
        RECT 473.200 203.600 474.000 204.400 ;
        RECT 476.400 203.600 477.200 204.400 ;
        RECT 479.600 203.600 480.400 204.400 ;
        RECT 486.000 213.600 486.800 214.400 ;
        RECT 495.600 213.000 496.400 213.800 ;
        RECT 505.200 212.600 506.000 213.400 ;
        RECT 519.600 217.600 520.400 218.400 ;
        RECT 511.600 211.600 512.400 212.400 ;
        RECT 497.200 208.800 498.000 209.600 ;
        RECT 502.000 207.600 502.800 208.400 ;
        RECT 498.800 206.200 499.600 207.000 ;
        RECT 495.600 204.200 496.400 205.000 ;
        RECT 497.200 204.200 498.000 205.000 ;
        RECT 502.000 206.200 502.800 207.000 ;
        RECT 505.200 206.200 506.000 207.000 ;
        RECT 506.800 204.200 507.600 205.000 ;
        RECT 508.400 204.200 509.200 205.000 ;
        RECT 510.000 204.200 510.800 205.000 ;
        RECT 534.000 217.600 534.800 218.400 ;
        RECT 538.800 217.600 539.600 218.400 ;
        RECT 530.800 209.600 531.600 210.400 ;
        RECT 554.800 215.600 555.600 216.400 ;
        RECT 556.400 214.200 557.200 215.000 ;
        RECT 604.400 217.600 605.200 218.400 ;
        RECT 578.800 213.600 579.600 214.400 ;
        RECT 567.600 211.600 568.400 212.400 ;
        RECT 550.000 206.800 550.800 207.600 ;
        RECT 553.200 206.200 554.000 207.000 ;
        RECT 548.400 204.200 549.200 205.000 ;
        RECT 550.000 204.200 550.800 205.000 ;
        RECT 551.600 204.200 552.400 205.000 ;
        RECT 556.400 206.200 557.200 207.000 ;
        RECT 559.600 206.200 560.400 207.000 ;
        RECT 575.600 211.600 576.400 212.400 ;
        RECT 591.600 213.600 592.400 214.400 ;
        RECT 561.200 204.200 562.000 205.000 ;
        RECT 562.800 204.200 563.600 205.000 ;
        RECT 577.200 209.600 578.000 210.400 ;
        RECT 18.800 195.000 19.600 195.800 ;
        RECT 15.600 193.600 16.400 194.400 ;
        RECT 33.200 197.600 34.000 198.400 ;
        RECT 20.400 192.400 21.200 193.200 ;
        RECT 25.200 189.600 26.000 190.400 ;
        RECT 9.200 188.200 10.000 189.000 ;
        RECT 18.800 188.600 19.600 189.400 ;
        RECT 14.000 187.600 14.800 188.400 ;
        RECT 9.200 184.200 10.000 185.000 ;
        RECT 10.800 184.200 11.600 185.000 ;
        RECT 12.400 184.200 13.200 185.000 ;
        RECT 15.600 184.200 16.400 185.000 ;
        RECT 18.800 184.200 19.600 185.000 ;
        RECT 20.400 184.200 21.200 185.000 ;
        RECT 22.000 184.200 22.800 185.000 ;
        RECT 23.600 184.200 24.400 185.000 ;
        RECT 57.200 195.600 58.000 196.400 ;
        RECT 41.200 187.600 42.000 188.400 ;
        RECT 38.000 185.600 38.800 186.400 ;
        RECT 39.600 186.200 40.400 187.000 ;
        RECT 36.400 183.600 37.200 184.400 ;
        RECT 62.000 189.600 62.800 190.400 ;
        RECT 66.800 189.600 67.600 190.400 ;
        RECT 82.800 197.600 83.600 198.400 ;
        RECT 63.600 187.600 64.400 188.400 ;
        RECT 78.000 189.600 78.800 190.400 ;
        RECT 79.600 189.600 80.400 190.400 ;
        RECT 86.000 189.600 86.800 190.400 ;
        RECT 94.000 189.600 94.800 190.400 ;
        RECT 89.200 187.600 90.000 188.400 ;
        RECT 82.800 183.600 83.600 184.400 ;
        RECT 87.600 186.200 88.400 187.000 ;
        RECT 108.400 189.600 109.200 190.400 ;
        RECT 113.200 189.600 114.000 190.400 ;
        RECT 114.800 189.600 115.600 190.400 ;
        RECT 126.000 189.600 126.800 190.400 ;
        RECT 129.200 189.600 130.000 190.400 ;
        RECT 130.800 189.600 131.600 190.400 ;
        RECT 105.200 183.600 106.000 184.400 ;
        RECT 127.600 187.600 128.400 188.400 ;
        RECT 142.000 197.600 142.800 198.400 ;
        RECT 145.200 197.600 146.000 198.400 ;
        RECT 158.000 197.600 158.800 198.400 ;
        RECT 146.800 185.600 147.600 186.400 ;
        RECT 145.200 183.600 146.000 184.400 ;
        RECT 162.600 191.800 163.400 192.600 ;
        RECT 185.200 194.400 186.000 195.200 ;
        RECT 188.400 195.000 189.200 195.800 ;
        RECT 209.200 197.600 210.000 198.400 ;
        RECT 183.600 192.400 184.400 193.200 ;
        RECT 159.600 185.600 160.400 186.400 ;
        RECT 162.600 186.200 163.400 187.000 ;
        RECT 170.800 187.600 171.600 188.400 ;
        RECT 182.000 189.600 182.800 190.400 ;
        RECT 193.200 187.600 194.000 188.400 ;
        RECT 190.000 185.600 190.800 186.400 ;
        RECT 183.600 184.200 184.400 185.000 ;
        RECT 185.200 184.200 186.000 185.000 ;
        RECT 186.800 184.200 187.600 185.000 ;
        RECT 188.400 184.200 189.200 185.000 ;
        RECT 191.600 184.200 192.400 185.000 ;
        RECT 194.800 184.200 195.600 185.000 ;
        RECT 196.400 184.200 197.200 185.000 ;
        RECT 198.000 184.200 198.800 185.000 ;
        RECT 217.200 193.600 218.000 194.400 ;
        RECT 214.000 189.600 214.800 190.400 ;
        RECT 218.800 189.600 219.600 190.400 ;
        RECT 210.800 187.600 211.600 188.400 ;
        RECT 215.600 187.600 216.400 188.400 ;
        RECT 236.400 193.600 237.200 194.400 ;
        RECT 233.200 189.600 234.000 190.400 ;
        RECT 234.800 189.600 235.600 190.400 ;
        RECT 239.600 189.600 240.400 190.400 ;
        RECT 225.200 183.600 226.000 184.400 ;
        RECT 254.000 189.600 254.800 190.400 ;
        RECT 273.200 195.000 274.000 195.800 ;
        RECT 270.000 193.600 270.800 194.400 ;
        RECT 274.800 192.400 275.600 193.200 ;
        RECT 287.600 193.600 288.400 194.400 ;
        RECT 300.400 197.600 301.200 198.400 ;
        RECT 310.000 197.600 310.800 198.400 ;
        RECT 263.600 188.200 264.400 189.000 ;
        RECT 273.200 188.600 274.000 189.400 ;
        RECT 268.400 187.600 269.200 188.400 ;
        RECT 263.600 184.200 264.400 185.000 ;
        RECT 265.200 184.200 266.000 185.000 ;
        RECT 266.800 184.200 267.600 185.000 ;
        RECT 270.000 184.200 270.800 185.000 ;
        RECT 273.200 184.200 274.000 185.000 ;
        RECT 274.800 184.200 275.600 185.000 ;
        RECT 276.400 184.200 277.200 185.000 ;
        RECT 278.000 184.200 278.800 185.000 ;
        RECT 294.000 189.600 294.800 190.400 ;
        RECT 295.600 187.600 296.400 188.400 ;
        RECT 290.800 183.600 291.600 184.400 ;
        RECT 308.400 185.600 309.200 186.400 ;
        RECT 324.400 197.600 325.200 198.400 ;
        RECT 318.000 189.600 318.800 190.400 ;
        RECT 335.600 194.400 336.400 195.200 ;
        RECT 338.800 195.000 339.600 195.800 ;
        RECT 334.000 192.400 334.800 193.200 ;
        RECT 311.600 185.600 312.400 186.400 ;
        RECT 332.400 189.600 333.200 190.400 ;
        RECT 321.200 183.600 322.000 184.400 ;
        RECT 366.000 193.600 366.800 194.400 ;
        RECT 343.600 187.600 344.400 188.400 ;
        RECT 340.400 185.600 341.200 186.400 ;
        RECT 377.200 194.400 378.000 195.200 ;
        RECT 380.400 195.000 381.200 195.800 ;
        RECT 375.600 192.400 376.400 193.200 ;
        RECT 361.200 189.600 362.000 190.400 ;
        RECT 334.000 184.200 334.800 185.000 ;
        RECT 335.600 184.200 336.400 185.000 ;
        RECT 337.200 184.200 338.000 185.000 ;
        RECT 338.800 184.200 339.600 185.000 ;
        RECT 342.000 184.200 342.800 185.000 ;
        RECT 345.200 184.200 346.000 185.000 ;
        RECT 346.800 184.200 347.600 185.000 ;
        RECT 348.400 184.200 349.200 185.000 ;
        RECT 374.000 189.600 374.800 190.400 ;
        RECT 358.000 183.600 358.800 184.400 ;
        RECT 385.200 187.600 386.000 188.400 ;
        RECT 382.000 185.600 382.800 186.400 ;
        RECT 375.600 184.200 376.400 185.000 ;
        RECT 377.200 184.200 378.000 185.000 ;
        RECT 378.800 184.200 379.600 185.000 ;
        RECT 380.400 184.200 381.200 185.000 ;
        RECT 383.600 184.200 384.400 185.000 ;
        RECT 386.800 184.200 387.600 185.000 ;
        RECT 388.400 184.200 389.200 185.000 ;
        RECT 390.000 184.200 390.800 185.000 ;
        RECT 417.200 195.000 418.000 195.800 ;
        RECT 414.000 193.600 414.800 194.400 ;
        RECT 418.800 192.400 419.600 193.200 ;
        RECT 407.600 188.200 408.400 189.000 ;
        RECT 417.200 188.600 418.000 189.400 ;
        RECT 412.400 187.600 413.200 188.400 ;
        RECT 407.600 184.200 408.400 185.000 ;
        RECT 409.200 184.200 410.000 185.000 ;
        RECT 410.800 184.200 411.600 185.000 ;
        RECT 414.000 184.200 414.800 185.000 ;
        RECT 417.200 184.200 418.000 185.000 ;
        RECT 418.800 184.200 419.600 185.000 ;
        RECT 420.400 184.200 421.200 185.000 ;
        RECT 422.000 184.200 422.800 185.000 ;
        RECT 452.400 195.000 453.200 195.800 ;
        RECT 449.200 193.600 450.000 194.400 ;
        RECT 454.000 192.400 454.800 193.200 ;
        RECT 442.800 188.200 443.600 189.000 ;
        RECT 452.400 188.600 453.200 189.400 ;
        RECT 431.600 183.600 432.400 184.400 ;
        RECT 447.600 187.600 448.400 188.400 ;
        RECT 442.800 184.200 443.600 185.000 ;
        RECT 444.400 184.200 445.200 185.000 ;
        RECT 446.000 184.200 446.800 185.000 ;
        RECT 449.200 184.200 450.000 185.000 ;
        RECT 452.400 184.200 453.200 185.000 ;
        RECT 454.000 184.200 454.800 185.000 ;
        RECT 455.600 184.200 456.400 185.000 ;
        RECT 457.200 184.200 458.000 185.000 ;
        RECT 489.200 193.600 490.000 194.400 ;
        RECT 474.800 186.200 475.600 187.000 ;
        RECT 466.800 183.600 467.600 184.400 ;
        RECT 495.600 189.600 496.400 190.400 ;
        RECT 510.000 191.600 510.800 192.400 ;
        RECT 503.600 187.600 504.400 188.400 ;
        RECT 519.600 187.600 520.400 188.400 ;
        RECT 492.400 183.600 493.200 184.400 ;
        RECT 498.800 183.600 499.600 184.400 ;
        RECT 516.400 185.600 517.200 186.400 ;
        RECT 522.800 187.600 523.600 188.400 ;
        RECT 514.800 183.600 515.600 184.400 ;
        RECT 540.400 194.400 541.200 195.200 ;
        RECT 543.600 195.000 544.400 195.800 ;
        RECT 538.800 192.400 539.600 193.200 ;
        RECT 537.200 189.600 538.000 190.400 ;
        RECT 526.000 185.600 526.800 186.400 ;
        RECT 529.200 183.600 530.000 184.400 ;
        RECT 548.400 187.600 549.200 188.400 ;
        RECT 545.200 185.600 546.000 186.400 ;
        RECT 538.800 184.200 539.600 185.000 ;
        RECT 540.400 184.200 541.200 185.000 ;
        RECT 542.000 184.200 542.800 185.000 ;
        RECT 543.600 184.200 544.400 185.000 ;
        RECT 546.800 184.200 547.600 185.000 ;
        RECT 550.000 184.200 550.800 185.000 ;
        RECT 551.600 184.200 552.400 185.000 ;
        RECT 553.200 184.200 554.000 185.000 ;
        RECT 580.400 195.000 581.200 195.800 ;
        RECT 577.200 193.600 578.000 194.400 ;
        RECT 582.000 192.400 582.800 193.200 ;
        RECT 570.800 188.200 571.600 189.000 ;
        RECT 580.400 188.600 581.200 189.400 ;
        RECT 575.600 187.600 576.400 188.400 ;
        RECT 595.000 189.600 595.800 190.400 ;
        RECT 570.800 184.200 571.600 185.000 ;
        RECT 572.400 184.200 573.200 185.000 ;
        RECT 574.000 184.200 574.800 185.000 ;
        RECT 577.200 184.200 578.000 185.000 ;
        RECT 580.400 184.200 581.200 185.000 ;
        RECT 582.000 184.200 582.800 185.000 ;
        RECT 583.600 184.200 584.400 185.000 ;
        RECT 585.200 184.200 586.000 185.000 ;
        RECT 601.200 189.600 602.000 190.400 ;
        RECT 602.800 187.600 603.600 188.400 ;
        RECT 598.000 183.600 598.800 184.400 ;
        RECT 1.200 170.200 2.000 171.000 ;
        RECT 38.000 177.600 38.800 178.400 ;
        RECT 18.800 167.600 19.600 168.400 ;
        RECT 33.200 171.600 34.000 172.400 ;
        RECT 41.200 171.600 42.000 172.400 ;
        RECT 52.400 177.600 53.200 178.400 ;
        RECT 38.000 163.600 38.800 164.400 ;
        RECT 46.000 163.600 46.800 164.400 ;
        RECT 76.400 175.600 77.200 176.400 ;
        RECT 68.400 173.600 69.200 174.400 ;
        RECT 57.200 172.200 58.000 173.000 ;
        RECT 65.200 171.800 66.000 172.600 ;
        RECT 73.200 171.600 74.000 172.400 ;
        RECT 70.000 170.200 70.800 171.000 ;
        RECT 102.000 177.600 102.800 178.400 ;
        RECT 98.800 171.600 99.600 172.400 ;
        RECT 113.200 169.600 114.000 170.400 ;
        RECT 111.600 163.600 112.400 164.400 ;
        RECT 116.400 163.600 117.200 164.400 ;
        RECT 121.200 169.600 122.000 170.400 ;
        RECT 119.600 163.600 120.400 164.400 ;
        RECT 132.400 177.600 133.200 178.400 ;
        RECT 129.200 171.600 130.000 172.400 ;
        RECT 135.600 171.600 136.400 172.400 ;
        RECT 140.400 171.600 141.200 172.400 ;
        RECT 167.600 175.600 168.400 176.400 ;
        RECT 169.200 174.200 170.000 175.000 ;
        RECT 193.200 177.600 194.000 178.400 ;
        RECT 180.400 171.600 181.200 172.400 ;
        RECT 138.800 163.600 139.600 164.400 ;
        RECT 151.600 165.600 152.400 166.400 ;
        RECT 162.800 166.800 163.600 167.600 ;
        RECT 166.000 166.200 166.800 167.000 ;
        RECT 161.200 164.200 162.000 165.000 ;
        RECT 162.800 164.200 163.600 165.000 ;
        RECT 164.400 164.200 165.200 165.000 ;
        RECT 169.200 166.200 170.000 167.000 ;
        RECT 172.400 166.200 173.200 167.000 ;
        RECT 190.000 171.600 190.800 172.400 ;
        RECT 174.000 164.200 174.800 165.000 ;
        RECT 175.600 164.200 176.400 165.000 ;
        RECT 191.600 169.600 192.400 170.400 ;
        RECT 196.400 169.600 197.200 170.400 ;
        RECT 225.200 175.600 226.000 176.400 ;
        RECT 226.800 174.200 227.600 175.000 ;
        RECT 238.000 171.600 238.800 172.400 ;
        RECT 209.200 169.600 210.000 170.400 ;
        RECT 220.400 166.800 221.200 167.600 ;
        RECT 223.600 166.200 224.400 167.000 ;
        RECT 218.800 164.200 219.600 165.000 ;
        RECT 220.400 164.200 221.200 165.000 ;
        RECT 222.000 164.200 222.800 165.000 ;
        RECT 226.800 166.200 227.600 167.000 ;
        RECT 230.000 166.200 230.800 167.000 ;
        RECT 250.800 173.000 251.600 173.800 ;
        RECT 260.400 172.600 261.200 173.400 ;
        RECT 274.800 177.600 275.600 178.400 ;
        RECT 249.200 171.600 250.000 172.400 ;
        RECT 252.400 168.800 253.200 169.600 ;
        RECT 257.200 167.600 258.000 168.400 ;
        RECT 231.600 164.200 232.400 165.000 ;
        RECT 233.200 164.200 234.000 165.000 ;
        RECT 254.000 166.200 254.800 167.000 ;
        RECT 250.800 164.200 251.600 165.000 ;
        RECT 252.400 164.200 253.200 165.000 ;
        RECT 257.200 166.200 258.000 167.000 ;
        RECT 260.400 166.200 261.200 167.000 ;
        RECT 262.000 164.200 262.800 165.000 ;
        RECT 263.600 164.200 264.400 165.000 ;
        RECT 265.200 164.200 266.000 165.000 ;
        RECT 278.000 169.600 278.800 170.400 ;
        RECT 310.000 173.000 310.800 173.800 ;
        RECT 284.400 163.600 285.200 164.400 ;
        RECT 319.600 172.600 320.400 173.400 ;
        RECT 340.400 177.600 341.200 178.400 ;
        RECT 326.000 171.600 326.800 172.400 ;
        RECT 311.600 168.800 312.400 169.600 ;
        RECT 316.400 167.600 317.200 168.400 ;
        RECT 313.200 166.200 314.000 167.000 ;
        RECT 310.000 164.200 310.800 165.000 ;
        RECT 311.600 164.200 312.400 165.000 ;
        RECT 316.400 166.200 317.200 167.000 ;
        RECT 319.600 166.200 320.400 167.000 ;
        RECT 321.200 164.200 322.000 165.000 ;
        RECT 322.800 164.200 323.600 165.000 ;
        RECT 324.400 164.200 325.200 165.000 ;
        RECT 334.000 169.600 334.800 170.400 ;
        RECT 350.000 175.600 350.800 176.400 ;
        RECT 343.600 173.600 344.400 174.400 ;
        RECT 340.400 169.600 341.200 170.400 ;
        RECT 362.800 177.600 363.600 178.400 ;
        RECT 351.600 169.600 352.400 170.400 ;
        RECT 374.000 177.600 374.800 178.400 ;
        RECT 380.400 177.600 381.200 178.400 ;
        RECT 369.200 173.600 370.000 174.400 ;
        RECT 362.800 169.600 363.600 170.400 ;
        RECT 369.200 169.600 370.000 170.400 ;
        RECT 380.400 169.600 381.200 170.400 ;
        RECT 385.200 177.600 386.000 178.400 ;
        RECT 401.200 173.600 402.000 174.400 ;
        RECT 390.000 172.200 390.800 173.000 ;
        RECT 398.000 171.800 398.800 172.600 ;
        RECT 402.800 170.200 403.600 171.000 ;
        RECT 409.200 169.600 410.000 170.400 ;
        RECT 433.200 173.600 434.000 174.400 ;
        RECT 426.800 170.200 427.600 171.000 ;
        RECT 449.200 171.600 450.000 172.400 ;
        RECT 444.400 163.600 445.200 164.400 ;
        RECT 468.400 169.600 469.200 170.400 ;
        RECT 474.800 169.600 475.600 170.400 ;
        RECT 510.000 177.600 510.800 178.400 ;
        RECT 502.000 173.600 502.800 174.400 ;
        RECT 550.000 177.600 550.800 178.400 ;
        RECT 490.800 172.200 491.600 173.000 ;
        RECT 503.600 170.200 504.400 171.000 ;
        RECT 486.000 167.600 486.800 168.400 ;
        RECT 524.400 171.600 525.200 172.400 ;
        RECT 534.000 171.600 534.800 172.400 ;
        RECT 540.400 171.600 541.200 172.400 ;
        RECT 532.400 163.600 533.200 164.400 ;
        RECT 542.000 169.600 542.800 170.400 ;
        RECT 548.400 169.600 549.200 170.400 ;
        RECT 556.400 169.600 557.200 170.400 ;
        RECT 582.000 175.600 582.800 176.400 ;
        RECT 583.600 174.200 584.400 175.000 ;
        RECT 574.000 171.600 574.800 172.400 ;
        RECT 594.800 171.600 595.600 172.400 ;
        RECT 562.800 169.600 563.600 170.400 ;
        RECT 577.200 166.800 578.000 167.600 ;
        RECT 580.400 166.200 581.200 167.000 ;
        RECT 575.600 164.200 576.400 165.000 ;
        RECT 577.200 164.200 578.000 165.000 ;
        RECT 578.800 164.200 579.600 165.000 ;
        RECT 583.600 166.200 584.400 167.000 ;
        RECT 586.800 166.200 587.600 167.000 ;
        RECT 588.400 164.200 589.200 165.000 ;
        RECT 590.000 164.200 590.800 165.000 ;
        RECT 7.600 149.600 8.400 150.400 ;
        RECT 23.600 157.600 24.400 158.400 ;
        RECT 1.200 146.200 2.000 147.000 ;
        RECT 28.400 149.600 29.200 150.400 ;
        RECT 36.400 149.600 37.200 150.400 ;
        RECT 38.000 147.600 38.800 148.400 ;
        RECT 46.000 149.600 46.800 150.400 ;
        RECT 47.600 149.600 48.400 150.400 ;
        RECT 55.600 149.600 56.400 150.400 ;
        RECT 57.200 149.600 58.000 150.400 ;
        RECT 60.400 149.600 61.200 150.400 ;
        RECT 89.200 153.600 90.000 154.400 ;
        RECT 94.000 153.600 94.800 154.400 ;
        RECT 68.400 149.600 69.200 150.400 ;
        RECT 106.800 153.600 107.600 154.400 ;
        RECT 18.800 143.600 19.600 144.400 ;
        RECT 54.000 145.600 54.800 146.400 ;
        RECT 70.000 147.600 70.800 148.400 ;
        RECT 73.200 147.600 74.000 148.400 ;
        RECT 71.600 146.200 72.400 147.000 ;
        RECT 98.800 149.600 99.600 150.400 ;
        RECT 103.600 151.600 104.400 152.400 ;
        RECT 111.600 149.600 112.400 150.400 ;
        RECT 119.600 149.600 120.400 150.400 ;
        RECT 124.400 149.600 125.200 150.400 ;
        RECT 130.800 149.600 131.600 150.400 ;
        RECT 137.200 149.600 138.000 150.400 ;
        RECT 76.400 145.600 77.200 146.400 ;
        RECT 102.000 143.600 102.800 144.400 ;
        RECT 121.200 147.600 122.000 148.400 ;
        RECT 127.600 147.600 128.400 148.400 ;
        RECT 142.000 147.600 142.800 148.400 ;
        RECT 151.600 157.600 152.400 158.400 ;
        RECT 146.800 151.800 147.600 152.600 ;
        RECT 143.600 143.600 144.400 144.400 ;
        RECT 146.800 146.200 147.600 147.000 ;
        RECT 178.800 155.000 179.600 155.800 ;
        RECT 175.600 153.600 176.400 154.400 ;
        RECT 193.200 157.600 194.000 158.400 ;
        RECT 180.400 152.400 181.200 153.200 ;
        RECT 185.200 149.600 186.000 150.400 ;
        RECT 154.800 147.600 155.600 148.400 ;
        RECT 169.200 148.200 170.000 149.000 ;
        RECT 178.800 148.600 179.600 149.400 ;
        RECT 151.600 146.400 152.400 147.200 ;
        RECT 174.000 147.600 174.800 148.400 ;
        RECT 169.200 144.200 170.000 145.000 ;
        RECT 170.800 144.200 171.600 145.000 ;
        RECT 172.400 144.200 173.200 145.000 ;
        RECT 175.600 144.200 176.400 145.000 ;
        RECT 178.800 144.200 179.600 145.000 ;
        RECT 180.400 144.200 181.200 145.000 ;
        RECT 182.000 144.200 182.800 145.000 ;
        RECT 183.600 144.200 184.400 145.000 ;
        RECT 207.600 149.600 208.400 150.400 ;
        RECT 196.400 143.600 197.200 144.400 ;
        RECT 204.400 145.600 205.200 146.400 ;
        RECT 212.400 145.600 213.200 146.400 ;
        RECT 223.600 153.600 224.400 154.400 ;
        RECT 220.400 149.600 221.200 150.400 ;
        RECT 242.800 155.000 243.600 155.800 ;
        RECT 239.600 153.600 240.400 154.400 ;
        RECT 257.200 155.600 258.000 156.400 ;
        RECT 244.400 152.400 245.200 153.200 ;
        RECT 249.200 149.600 250.000 150.400 ;
        RECT 217.200 147.600 218.000 148.400 ;
        RECT 222.000 147.600 222.800 148.400 ;
        RECT 233.200 148.200 234.000 149.000 ;
        RECT 242.800 148.600 243.600 149.400 ;
        RECT 210.800 143.600 211.600 144.400 ;
        RECT 215.600 143.600 216.400 144.400 ;
        RECT 238.000 147.600 238.800 148.400 ;
        RECT 233.200 144.200 234.000 145.000 ;
        RECT 234.800 144.200 235.600 145.000 ;
        RECT 236.400 144.200 237.200 145.000 ;
        RECT 239.600 144.200 240.400 145.000 ;
        RECT 242.800 144.200 243.600 145.000 ;
        RECT 244.400 144.200 245.200 145.000 ;
        RECT 246.000 144.200 246.800 145.000 ;
        RECT 247.600 144.200 248.400 145.000 ;
        RECT 282.800 155.000 283.600 155.800 ;
        RECT 279.600 153.600 280.400 154.400 ;
        RECT 284.400 152.400 285.200 153.200 ;
        RECT 289.200 149.600 290.000 150.400 ;
        RECT 263.600 147.600 264.400 148.400 ;
        RECT 273.200 148.200 274.000 149.000 ;
        RECT 282.800 148.600 283.600 149.400 ;
        RECT 262.000 143.600 262.800 144.400 ;
        RECT 278.000 147.600 278.800 148.400 ;
        RECT 273.200 144.200 274.000 145.000 ;
        RECT 274.800 144.200 275.600 145.000 ;
        RECT 276.400 144.200 277.200 145.000 ;
        RECT 279.600 144.200 280.400 145.000 ;
        RECT 282.800 144.200 283.600 145.000 ;
        RECT 284.400 144.200 285.200 145.000 ;
        RECT 286.000 144.200 286.800 145.000 ;
        RECT 287.600 144.200 288.400 145.000 ;
        RECT 310.000 149.600 310.800 150.400 ;
        RECT 297.200 143.600 298.000 144.400 ;
        RECT 337.200 155.000 338.000 155.800 ;
        RECT 334.000 153.600 334.800 154.400 ;
        RECT 338.800 152.400 339.600 153.200 ;
        RECT 351.600 153.600 352.400 154.400 ;
        RECT 343.600 149.600 344.400 150.400 ;
        RECT 327.600 148.200 328.400 149.000 ;
        RECT 337.200 148.600 338.000 149.400 ;
        RECT 318.000 143.600 318.800 144.400 ;
        RECT 332.400 147.600 333.200 148.400 ;
        RECT 327.600 144.200 328.400 145.000 ;
        RECT 329.200 144.200 330.000 145.000 ;
        RECT 330.800 144.200 331.600 145.000 ;
        RECT 334.000 144.200 334.800 145.000 ;
        RECT 337.200 144.200 338.000 145.000 ;
        RECT 338.800 144.200 339.600 145.000 ;
        RECT 340.400 144.200 341.200 145.000 ;
        RECT 342.000 144.200 342.800 145.000 ;
        RECT 362.800 149.600 363.600 150.400 ;
        RECT 364.400 147.600 365.200 148.400 ;
        RECT 366.000 147.600 366.800 148.400 ;
        RECT 374.000 157.600 374.800 158.400 ;
        RECT 380.400 157.600 381.200 158.400 ;
        RECT 374.000 149.600 374.800 150.400 ;
        RECT 398.000 153.600 398.800 154.400 ;
        RECT 404.400 153.600 405.200 154.400 ;
        RECT 380.400 149.600 381.200 150.400 ;
        RECT 385.200 149.600 386.000 150.400 ;
        RECT 393.200 149.600 394.000 150.400 ;
        RECT 401.200 151.600 402.000 152.400 ;
        RECT 399.600 149.600 400.400 150.400 ;
        RECT 407.600 151.600 408.400 152.400 ;
        RECT 406.000 149.600 406.800 150.400 ;
        RECT 410.800 149.600 411.600 150.400 ;
        RECT 375.600 147.600 376.400 148.400 ;
        RECT 382.000 147.600 382.800 148.400 ;
        RECT 394.800 147.600 395.600 148.400 ;
        RECT 369.200 143.600 370.000 144.400 ;
        RECT 417.200 147.600 418.000 148.400 ;
        RECT 420.400 147.600 421.200 148.400 ;
        RECT 428.400 149.600 429.200 150.400 ;
        RECT 430.000 149.600 430.800 150.400 ;
        RECT 434.800 149.600 435.600 150.400 ;
        RECT 446.000 157.600 446.800 158.400 ;
        RECT 441.200 149.600 442.000 150.400 ;
        RECT 442.800 149.600 443.600 150.400 ;
        RECT 431.600 143.600 432.400 144.400 ;
        RECT 439.600 145.600 440.400 146.400 ;
        RECT 460.400 155.600 461.200 156.400 ;
        RECT 454.000 147.600 454.800 148.400 ;
        RECT 474.800 152.400 475.600 153.200 ;
        RECT 478.000 151.000 478.800 151.800 ;
        RECT 479.600 157.600 480.400 158.400 ;
        RECT 478.000 146.200 478.800 147.000 ;
        RECT 487.600 153.600 488.400 154.400 ;
        RECT 482.800 149.600 483.600 150.400 ;
        RECT 484.400 149.600 485.200 150.400 ;
        RECT 492.400 147.600 493.200 148.400 ;
        RECT 481.200 145.600 482.000 146.400 ;
        RECT 500.400 149.600 501.200 150.400 ;
        RECT 505.200 149.600 506.000 150.400 ;
        RECT 516.400 153.600 517.200 154.400 ;
        RECT 513.200 149.600 514.000 150.400 ;
        RECT 502.000 147.600 502.800 148.400 ;
        RECT 508.400 147.600 509.200 148.400 ;
        RECT 514.800 147.600 515.600 148.400 ;
        RECT 530.800 152.400 531.600 153.200 ;
        RECT 542.000 157.600 542.800 158.400 ;
        RECT 534.000 151.000 534.800 151.800 ;
        RECT 537.200 149.600 538.000 150.400 ;
        RECT 497.200 143.600 498.000 144.400 ;
        RECT 529.200 145.600 530.000 146.400 ;
        RECT 534.000 146.200 534.800 147.000 ;
        RECT 556.400 152.400 557.200 153.200 ;
        RECT 559.600 151.000 560.400 151.800 ;
        RECT 559.600 146.200 560.400 147.000 ;
        RECT 561.200 145.600 562.000 146.400 ;
        RECT 580.400 154.400 581.200 155.200 ;
        RECT 583.600 155.000 584.400 155.800 ;
        RECT 578.800 152.400 579.600 153.200 ;
        RECT 569.200 143.600 570.000 144.400 ;
        RECT 588.400 147.600 589.200 148.400 ;
        RECT 585.200 145.600 586.000 146.400 ;
        RECT 578.800 144.200 579.600 145.000 ;
        RECT 580.400 144.200 581.200 145.000 ;
        RECT 582.000 144.200 582.800 145.000 ;
        RECT 583.600 144.200 584.400 145.000 ;
        RECT 586.800 144.200 587.600 145.000 ;
        RECT 590.000 144.200 590.800 145.000 ;
        RECT 591.600 144.200 592.400 145.000 ;
        RECT 593.200 144.200 594.000 145.000 ;
        RECT 606.000 149.600 606.800 150.400 ;
        RECT 602.800 143.600 603.600 144.400 ;
        RECT 18.800 135.600 19.600 136.400 ;
        RECT 20.400 134.200 21.200 135.000 ;
        RECT 10.800 131.600 11.600 132.400 ;
        RECT 30.000 131.600 30.800 132.400 ;
        RECT 2.800 123.600 3.600 124.400 ;
        RECT 14.000 126.800 14.800 127.600 ;
        RECT 17.200 126.200 18.000 127.000 ;
        RECT 12.400 124.200 13.200 125.000 ;
        RECT 14.000 124.200 14.800 125.000 ;
        RECT 15.600 124.200 16.400 125.000 ;
        RECT 20.400 126.200 21.200 127.000 ;
        RECT 23.600 126.200 24.400 127.000 ;
        RECT 25.200 124.200 26.000 125.000 ;
        RECT 26.800 124.200 27.600 125.000 ;
        RECT 39.600 129.600 40.400 130.400 ;
        RECT 49.200 131.600 50.000 132.400 ;
        RECT 76.400 133.600 77.200 134.400 ;
        RECT 74.800 131.800 75.600 132.600 ;
        RECT 62.000 129.600 62.800 130.400 ;
        RECT 70.000 130.200 70.800 131.000 ;
        RECT 95.600 137.600 96.400 138.400 ;
        RECT 103.600 133.600 104.400 134.400 ;
        RECT 94.000 131.600 94.800 132.400 ;
        RECT 106.800 131.800 107.600 132.600 ;
        RECT 102.000 130.200 102.800 131.000 ;
        RECT 87.600 123.600 88.400 124.400 ;
        RECT 119.600 123.600 120.400 124.400 ;
        RECT 127.600 133.600 128.400 134.400 ;
        RECT 124.400 129.600 125.200 130.400 ;
        RECT 161.200 137.600 162.000 138.400 ;
        RECT 132.400 129.600 133.200 130.400 ;
        RECT 130.800 127.600 131.600 128.400 ;
        RECT 138.800 129.600 139.600 130.400 ;
        RECT 145.200 129.600 146.000 130.400 ;
        RECT 146.800 129.600 147.600 130.400 ;
        RECT 180.400 135.600 181.200 136.400 ;
        RECT 182.000 134.200 182.800 135.000 ;
        RECT 183.600 131.600 184.400 132.400 ;
        RECT 193.200 131.600 194.000 132.400 ;
        RECT 161.200 129.600 162.000 130.400 ;
        RECT 164.400 123.600 165.200 124.400 ;
        RECT 175.600 126.800 176.400 127.600 ;
        RECT 178.800 126.200 179.600 127.000 ;
        RECT 174.000 124.200 174.800 125.000 ;
        RECT 175.600 124.200 176.400 125.000 ;
        RECT 177.200 124.200 178.000 125.000 ;
        RECT 182.000 126.200 182.800 127.000 ;
        RECT 185.200 126.200 186.000 127.000 ;
        RECT 198.000 129.600 198.800 130.400 ;
        RECT 186.800 124.200 187.600 125.000 ;
        RECT 188.400 124.200 189.200 125.000 ;
        RECT 207.600 131.600 208.400 132.400 ;
        RECT 226.800 135.600 227.600 136.400 ;
        RECT 228.400 134.200 229.200 135.000 ;
        RECT 218.800 131.600 219.600 132.400 ;
        RECT 222.000 126.800 222.800 127.600 ;
        RECT 225.200 126.200 226.000 127.000 ;
        RECT 220.400 124.200 221.200 125.000 ;
        RECT 222.000 124.200 222.800 125.000 ;
        RECT 223.600 124.200 224.400 125.000 ;
        RECT 228.400 126.200 229.200 127.000 ;
        RECT 231.600 126.200 232.400 127.000 ;
        RECT 244.400 131.600 245.200 132.400 ;
        RECT 252.400 131.600 253.200 132.400 ;
        RECT 263.600 133.600 264.400 134.400 ;
        RECT 284.400 135.600 285.200 136.400 ;
        RECT 286.000 134.200 286.800 135.000 ;
        RECT 276.400 131.600 277.200 132.400 ;
        RECT 287.600 131.600 288.400 132.400 ;
        RECT 233.200 124.200 234.000 125.000 ;
        RECT 234.800 124.200 235.600 125.000 ;
        RECT 257.200 123.600 258.000 124.400 ;
        RECT 265.200 127.600 266.000 128.400 ;
        RECT 279.600 126.800 280.400 127.600 ;
        RECT 282.800 126.200 283.600 127.000 ;
        RECT 278.000 124.200 278.800 125.000 ;
        RECT 279.600 124.200 280.400 125.000 ;
        RECT 281.200 124.200 282.000 125.000 ;
        RECT 286.000 126.200 286.800 127.000 ;
        RECT 289.200 126.200 290.000 127.000 ;
        RECT 319.600 133.600 320.400 134.400 ;
        RECT 329.200 133.000 330.000 133.800 ;
        RECT 290.800 124.200 291.600 125.000 ;
        RECT 292.400 124.200 293.200 125.000 ;
        RECT 338.800 132.600 339.600 133.400 ;
        RECT 322.800 131.600 323.600 132.400 ;
        RECT 345.200 131.600 346.000 132.400 ;
        RECT 330.800 128.800 331.600 129.600 ;
        RECT 335.600 127.600 336.400 128.400 ;
        RECT 332.400 126.200 333.200 127.000 ;
        RECT 329.200 124.200 330.000 125.000 ;
        RECT 330.800 124.200 331.600 125.000 ;
        RECT 335.600 126.200 336.400 127.000 ;
        RECT 338.800 126.200 339.600 127.000 ;
        RECT 340.400 124.200 341.200 125.000 ;
        RECT 342.000 124.200 342.800 125.000 ;
        RECT 343.600 124.200 344.400 125.000 ;
        RECT 353.200 123.600 354.000 124.400 ;
        RECT 362.800 133.600 363.600 134.400 ;
        RECT 386.800 133.000 387.600 133.800 ;
        RECT 377.200 129.600 378.000 130.400 ;
        RECT 396.400 132.600 397.200 133.400 ;
        RECT 382.000 131.600 382.800 132.400 ;
        RECT 414.000 133.600 414.800 134.400 ;
        RECT 426.800 133.600 427.600 134.400 ;
        RECT 388.400 128.800 389.200 129.600 ;
        RECT 393.200 127.600 394.000 128.400 ;
        RECT 390.000 126.200 390.800 127.000 ;
        RECT 386.800 124.200 387.600 125.000 ;
        RECT 388.400 124.200 389.200 125.000 ;
        RECT 393.200 126.200 394.000 127.000 ;
        RECT 396.400 126.200 397.200 127.000 ;
        RECT 398.000 124.200 398.800 125.000 ;
        RECT 399.600 124.200 400.400 125.000 ;
        RECT 401.200 124.200 402.000 125.000 ;
        RECT 410.800 127.600 411.600 128.400 ;
        RECT 415.600 123.600 416.400 124.400 ;
        RECT 455.600 134.800 456.400 135.600 ;
        RECT 444.400 131.600 445.200 132.400 ;
        RECT 431.600 123.600 432.400 124.400 ;
        RECT 450.800 131.600 451.600 132.400 ;
        RECT 444.400 123.600 445.200 124.400 ;
        RECT 474.800 131.600 475.600 132.400 ;
        RECT 481.200 129.600 482.000 130.400 ;
        RECT 506.800 137.600 507.600 138.400 ;
        RECT 518.000 137.600 518.800 138.400 ;
        RECT 487.600 131.600 488.400 132.400 ;
        RECT 497.200 131.600 498.000 132.400 ;
        RECT 492.400 129.600 493.200 130.400 ;
        RECT 510.000 131.600 510.800 132.400 ;
        RECT 514.800 131.600 515.600 132.400 ;
        RECT 529.200 133.600 530.000 134.400 ;
        RECT 522.800 132.200 523.600 133.000 ;
        RECT 516.400 129.600 517.200 130.400 ;
        RECT 540.400 131.600 541.200 132.400 ;
        RECT 535.600 130.200 536.400 131.000 ;
        RECT 559.600 137.600 560.400 138.400 ;
        RECT 550.000 123.600 550.800 124.400 ;
        RECT 567.600 129.600 568.400 130.400 ;
        RECT 575.600 131.600 576.400 132.400 ;
        RECT 583.600 129.600 584.400 130.400 ;
        RECT 607.600 137.600 608.400 138.400 ;
        RECT 591.600 133.600 592.400 134.400 ;
        RECT 594.800 131.800 595.600 132.600 ;
        RECT 590.000 130.200 590.800 131.000 ;
        RECT 18.800 113.600 19.600 114.400 ;
        RECT 1.200 106.200 2.000 107.000 ;
        RECT 34.800 117.600 35.600 118.400 ;
        RECT 23.600 109.600 24.400 110.400 ;
        RECT 30.000 109.600 30.800 110.400 ;
        RECT 25.200 107.600 26.000 108.400 ;
        RECT 34.800 107.600 35.600 108.400 ;
        RECT 38.000 109.600 38.800 110.400 ;
        RECT 46.000 109.600 46.800 110.400 ;
        RECT 47.600 109.600 48.400 110.400 ;
        RECT 50.800 109.600 51.600 110.400 ;
        RECT 60.400 107.600 61.200 108.400 ;
        RECT 73.200 111.600 74.000 112.400 ;
        RECT 94.000 117.600 94.800 118.400 ;
        RECT 86.000 113.600 86.800 114.400 ;
        RECT 68.400 109.600 69.200 110.400 ;
        RECT 70.000 109.600 70.800 110.400 ;
        RECT 82.800 109.600 83.600 110.400 ;
        RECT 84.400 107.600 85.200 108.400 ;
        RECT 79.600 103.600 80.400 104.400 ;
        RECT 92.400 113.600 93.200 114.400 ;
        RECT 89.200 111.600 90.000 112.400 ;
        RECT 98.800 111.600 99.600 112.400 ;
        RECT 98.800 109.600 99.600 110.400 ;
        RECT 110.000 109.600 110.800 110.400 ;
        RECT 118.000 109.600 118.800 110.400 ;
        RECT 100.400 107.600 101.200 108.400 ;
        RECT 134.000 117.600 134.800 118.400 ;
        RECT 129.200 103.600 130.000 104.400 ;
        RECT 156.400 117.600 157.200 118.400 ;
        RECT 145.200 109.600 146.000 110.400 ;
        RECT 170.800 117.600 171.600 118.400 ;
        RECT 137.200 107.600 138.000 108.400 ;
        RECT 140.400 107.600 141.200 108.400 ;
        RECT 146.800 107.600 147.600 108.400 ;
        RECT 158.000 107.600 158.800 108.400 ;
        RECT 174.000 109.600 174.800 110.400 ;
        RECT 175.600 109.600 176.400 110.400 ;
        RECT 183.600 109.600 184.400 110.400 ;
        RECT 185.200 109.600 186.000 110.400 ;
        RECT 195.000 111.800 195.800 112.600 ;
        RECT 196.200 109.800 197.000 110.600 ;
        RECT 220.400 113.600 221.200 114.400 ;
        RECT 223.600 113.600 224.400 114.400 ;
        RECT 217.200 111.600 218.000 112.400 ;
        RECT 195.000 106.200 195.800 107.000 ;
        RECT 178.800 103.600 179.600 104.400 ;
        RECT 202.800 107.600 203.600 108.400 ;
        RECT 207.600 107.600 208.400 108.400 ;
        RECT 204.400 103.600 205.200 104.400 ;
        RECT 212.400 103.600 213.200 104.400 ;
        RECT 225.200 105.600 226.000 106.400 ;
        RECT 226.800 105.600 227.600 106.400 ;
        RECT 241.200 109.600 242.000 110.400 ;
        RECT 262.000 115.000 262.800 115.800 ;
        RECT 258.800 113.600 259.600 114.400 ;
        RECT 263.600 112.400 264.400 113.200 ;
        RECT 250.800 111.200 251.600 112.000 ;
        RECT 276.400 113.600 277.200 114.400 ;
        RECT 294.200 111.800 295.000 112.600 ;
        RECT 233.200 105.600 234.000 106.400 ;
        RECT 242.800 107.600 243.600 108.400 ;
        RECT 252.400 108.200 253.200 109.000 ;
        RECT 262.000 108.600 262.800 109.400 ;
        RECT 238.000 103.600 238.800 104.400 ;
        RECT 257.200 107.600 258.000 108.400 ;
        RECT 252.400 104.200 253.200 105.000 ;
        RECT 254.000 104.200 254.800 105.000 ;
        RECT 255.600 104.200 256.400 105.000 ;
        RECT 258.800 104.200 259.600 105.000 ;
        RECT 262.000 104.200 262.800 105.000 ;
        RECT 263.600 104.200 264.400 105.000 ;
        RECT 265.200 104.200 266.000 105.000 ;
        RECT 266.800 104.200 267.600 105.000 ;
        RECT 282.800 109.600 283.600 110.400 ;
        RECT 281.200 107.600 282.000 108.400 ;
        RECT 284.400 107.600 285.200 108.400 ;
        RECT 290.800 109.600 291.600 110.400 ;
        RECT 295.400 109.800 296.200 110.600 ;
        RECT 294.200 106.200 295.000 107.000 ;
        RECT 302.000 107.600 302.800 108.400 ;
        RECT 308.400 107.600 309.200 108.400 ;
        RECT 297.200 103.600 298.000 104.400 ;
        RECT 314.800 117.600 315.600 118.400 ;
        RECT 326.000 114.400 326.800 115.200 ;
        RECT 329.200 115.000 330.000 115.800 ;
        RECT 324.400 112.400 325.200 113.200 ;
        RECT 322.800 109.600 323.600 110.400 ;
        RECT 334.000 107.600 334.800 108.400 ;
        RECT 330.800 105.600 331.600 106.400 ;
        RECT 324.400 104.200 325.200 105.000 ;
        RECT 326.000 104.200 326.800 105.000 ;
        RECT 327.600 104.200 328.400 105.000 ;
        RECT 329.200 104.200 330.000 105.000 ;
        RECT 332.400 104.200 333.200 105.000 ;
        RECT 335.600 104.200 336.400 105.000 ;
        RECT 337.200 104.200 338.000 105.000 ;
        RECT 338.800 104.200 339.600 105.000 ;
        RECT 350.000 107.600 350.800 108.400 ;
        RECT 358.000 103.600 358.800 104.400 ;
        RECT 388.400 115.000 389.200 115.800 ;
        RECT 385.200 113.600 386.000 114.400 ;
        RECT 390.000 112.400 390.800 113.200 ;
        RECT 406.000 117.600 406.800 118.400 ;
        RECT 394.800 109.600 395.600 110.400 ;
        RECT 369.200 107.600 370.000 108.400 ;
        RECT 378.800 108.200 379.600 109.000 ;
        RECT 388.400 108.600 389.200 109.400 ;
        RECT 362.800 105.600 363.600 106.400 ;
        RECT 383.600 107.600 384.400 108.400 ;
        RECT 378.800 104.200 379.600 105.000 ;
        RECT 380.400 104.200 381.200 105.000 ;
        RECT 382.000 104.200 382.800 105.000 ;
        RECT 385.200 104.200 386.000 105.000 ;
        RECT 388.400 104.200 389.200 105.000 ;
        RECT 390.000 104.200 390.800 105.000 ;
        RECT 391.600 104.200 392.400 105.000 ;
        RECT 393.200 104.200 394.000 105.000 ;
        RECT 420.400 112.400 421.200 113.200 ;
        RECT 423.600 111.000 424.400 111.800 ;
        RECT 426.800 117.600 427.600 118.400 ;
        RECT 407.600 107.600 408.400 108.400 ;
        RECT 402.800 103.600 403.600 104.400 ;
        RECT 423.600 106.200 424.400 107.000 ;
        RECT 425.200 105.600 426.000 106.400 ;
        RECT 433.200 107.600 434.000 108.400 ;
        RECT 441.200 109.600 442.000 110.400 ;
        RECT 454.000 109.600 454.800 110.400 ;
        RECT 444.400 105.600 445.200 106.400 ;
        RECT 455.600 107.600 456.400 108.400 ;
        RECT 462.000 107.600 462.800 108.400 ;
        RECT 468.400 105.600 469.200 106.400 ;
        RECT 471.600 105.600 472.400 106.400 ;
        RECT 481.200 117.600 482.000 118.400 ;
        RECT 486.000 109.600 486.800 110.400 ;
        RECT 505.200 117.600 506.000 118.400 ;
        RECT 478.000 105.600 478.800 106.400 ;
        RECT 487.600 107.600 488.400 108.400 ;
        RECT 492.400 107.600 493.200 108.400 ;
        RECT 500.400 107.600 501.200 108.400 ;
        RECT 503.600 113.600 504.400 114.400 ;
        RECT 482.800 103.600 483.600 104.400 ;
        RECT 498.800 103.600 499.600 104.400 ;
        RECT 518.000 109.600 518.800 110.400 ;
        RECT 521.200 109.600 522.000 110.400 ;
        RECT 522.800 109.600 523.600 110.400 ;
        RECT 526.000 109.600 526.800 110.400 ;
        RECT 537.200 113.600 538.000 114.400 ;
        RECT 534.000 109.600 534.800 110.400 ;
        RECT 506.800 105.600 507.600 106.400 ;
        RECT 529.200 107.600 530.000 108.400 ;
        RECT 513.200 103.600 514.000 104.400 ;
        RECT 535.600 107.600 536.400 108.400 ;
        RECT 551.600 112.400 552.400 113.200 ;
        RECT 554.800 111.000 555.600 111.800 ;
        RECT 564.400 109.600 565.200 110.400 ;
        RECT 582.000 114.400 582.800 115.200 ;
        RECT 585.200 115.000 586.000 115.800 ;
        RECT 580.400 112.400 581.200 113.200 ;
        RECT 554.800 106.200 555.600 107.000 ;
        RECT 578.800 109.600 579.600 110.400 ;
        RECT 590.000 107.600 590.800 108.400 ;
        RECT 586.800 105.600 587.600 106.400 ;
        RECT 607.600 109.600 608.400 110.400 ;
        RECT 580.400 104.200 581.200 105.000 ;
        RECT 582.000 104.200 582.800 105.000 ;
        RECT 583.600 104.200 584.400 105.000 ;
        RECT 585.200 104.200 586.000 105.000 ;
        RECT 588.400 104.200 589.200 105.000 ;
        RECT 591.600 104.200 592.400 105.000 ;
        RECT 593.200 104.200 594.000 105.000 ;
        RECT 594.800 104.200 595.600 105.000 ;
        RECT 609.200 107.600 610.000 108.400 ;
        RECT 12.400 93.600 13.200 94.400 ;
        RECT 20.400 97.600 21.200 98.400 ;
        RECT 42.800 97.600 43.600 98.400 ;
        RECT 6.000 92.200 6.800 93.000 ;
        RECT 14.000 91.800 14.800 92.600 ;
        RECT 18.800 90.200 19.600 91.000 ;
        RECT 1.200 87.600 2.000 88.400 ;
        RECT 55.600 93.600 56.400 94.400 ;
        RECT 34.800 91.600 35.600 92.400 ;
        RECT 36.400 91.600 37.200 92.400 ;
        RECT 23.600 83.600 24.400 84.400 ;
        RECT 31.600 89.600 32.400 90.400 ;
        RECT 49.200 90.200 50.000 91.000 ;
        RECT 79.600 95.600 80.400 96.400 ;
        RECT 97.200 97.600 98.000 98.400 ;
        RECT 114.800 97.600 115.600 98.400 ;
        RECT 66.800 87.600 67.600 88.400 ;
        RECT 110.000 91.600 110.800 92.400 ;
        RECT 111.600 89.600 112.400 90.400 ;
        RECT 87.600 83.600 88.400 84.400 ;
        RECT 121.200 89.600 122.000 90.400 ;
        RECT 140.400 97.600 141.200 98.400 ;
        RECT 143.600 97.600 144.400 98.400 ;
        RECT 130.800 83.600 131.600 84.400 ;
        RECT 140.400 89.600 141.200 90.400 ;
        RECT 142.000 89.600 142.800 90.400 ;
        RECT 150.000 91.600 150.800 92.400 ;
        RECT 169.200 93.600 170.000 94.400 ;
        RECT 162.800 92.200 163.600 93.000 ;
        RECT 185.200 93.000 186.000 93.800 ;
        RECT 170.800 91.800 171.600 92.600 ;
        RECT 175.600 90.200 176.400 91.000 ;
        RECT 158.000 83.600 158.800 84.400 ;
        RECT 194.800 92.600 195.600 93.400 ;
        RECT 209.200 97.600 210.000 98.400 ;
        RECT 182.000 91.600 182.800 92.400 ;
        RECT 201.200 91.600 202.000 92.400 ;
        RECT 186.800 88.800 187.600 89.600 ;
        RECT 191.600 87.600 192.400 88.400 ;
        RECT 188.400 86.200 189.200 87.000 ;
        RECT 185.200 84.200 186.000 85.000 ;
        RECT 186.800 84.200 187.600 85.000 ;
        RECT 191.600 86.200 192.400 87.000 ;
        RECT 194.800 86.200 195.600 87.000 ;
        RECT 196.400 84.200 197.200 85.000 ;
        RECT 198.000 84.200 198.800 85.000 ;
        RECT 199.600 84.200 200.400 85.000 ;
        RECT 215.600 89.600 216.400 90.400 ;
        RECT 222.000 89.600 222.800 90.400 ;
        RECT 247.600 97.600 248.400 98.400 ;
        RECT 231.600 93.200 232.400 94.000 ;
        RECT 234.800 89.600 235.600 90.400 ;
        RECT 244.400 89.600 245.200 90.400 ;
        RECT 250.800 95.600 251.600 96.400 ;
        RECT 266.800 95.600 267.600 96.400 ;
        RECT 268.400 94.200 269.200 95.000 ;
        RECT 279.600 91.600 280.400 92.400 ;
        RECT 262.000 86.800 262.800 87.600 ;
        RECT 265.200 86.200 266.000 87.000 ;
        RECT 260.400 84.200 261.200 85.000 ;
        RECT 262.000 84.200 262.800 85.000 ;
        RECT 263.600 84.200 264.400 85.000 ;
        RECT 268.400 86.200 269.200 87.000 ;
        RECT 271.600 86.200 272.400 87.000 ;
        RECT 292.400 93.000 293.200 93.800 ;
        RECT 302.000 92.600 302.800 93.400 ;
        RECT 286.000 91.600 286.800 92.400 ;
        RECT 287.600 91.600 288.400 92.400 ;
        RECT 316.600 93.600 317.400 94.400 ;
        RECT 294.000 88.800 294.800 89.600 ;
        RECT 298.800 87.600 299.600 88.400 ;
        RECT 273.200 84.200 274.000 85.000 ;
        RECT 274.800 84.200 275.600 85.000 ;
        RECT 295.600 86.200 296.400 87.000 ;
        RECT 292.400 84.200 293.200 85.000 ;
        RECT 294.000 84.200 294.800 85.000 ;
        RECT 298.800 86.200 299.600 87.000 ;
        RECT 302.000 86.200 302.800 87.000 ;
        RECT 303.600 84.200 304.400 85.000 ;
        RECT 305.200 84.200 306.000 85.000 ;
        RECT 306.800 84.200 307.600 85.000 ;
        RECT 332.400 97.600 333.200 98.400 ;
        RECT 348.400 95.600 349.200 96.400 ;
        RECT 350.000 94.200 350.800 95.000 ;
        RECT 326.000 83.600 326.800 84.400 ;
        RECT 358.000 90.000 358.800 90.800 ;
        RECT 343.600 86.800 344.400 87.600 ;
        RECT 346.800 86.200 347.600 87.000 ;
        RECT 342.000 84.200 342.800 85.000 ;
        RECT 343.600 84.200 344.400 85.000 ;
        RECT 345.200 84.200 346.000 85.000 ;
        RECT 350.000 86.200 350.800 87.000 ;
        RECT 353.200 86.200 354.000 87.000 ;
        RECT 374.000 93.000 374.800 93.800 ;
        RECT 383.600 92.600 384.400 93.400 ;
        RECT 401.200 97.600 402.000 98.400 ;
        RECT 369.200 91.600 370.000 92.400 ;
        RECT 422.000 97.600 422.800 98.400 ;
        RECT 375.600 88.800 376.400 89.600 ;
        RECT 380.400 87.600 381.200 88.400 ;
        RECT 354.800 84.200 355.600 85.000 ;
        RECT 356.400 84.200 357.200 85.000 ;
        RECT 377.200 86.200 378.000 87.000 ;
        RECT 374.000 84.200 374.800 85.000 ;
        RECT 375.600 84.200 376.400 85.000 ;
        RECT 380.400 86.200 381.200 87.000 ;
        RECT 383.600 86.200 384.400 87.000 ;
        RECT 385.200 84.200 386.000 85.000 ;
        RECT 386.800 84.200 387.600 85.000 ;
        RECT 388.400 84.200 389.200 85.000 ;
        RECT 398.000 83.600 398.800 84.400 ;
        RECT 414.000 93.600 414.800 94.400 ;
        RECT 433.200 97.600 434.000 98.400 ;
        RECT 418.800 91.600 419.600 92.400 ;
        RECT 415.600 89.600 416.400 90.400 ;
        RECT 426.800 91.600 427.600 92.400 ;
        RECT 449.200 97.600 450.000 98.400 ;
        RECT 436.400 91.600 437.200 92.400 ;
        RECT 444.400 91.600 445.200 92.400 ;
        RECT 442.800 89.600 443.600 90.400 ;
        RECT 455.600 89.600 456.400 90.400 ;
        RECT 457.200 89.600 458.000 90.400 ;
        RECT 471.600 91.600 472.400 92.400 ;
        RECT 470.000 83.600 470.800 84.400 ;
        RECT 516.400 97.600 517.200 98.400 ;
        RECT 479.600 83.600 480.400 84.400 ;
        RECT 495.600 89.600 496.400 90.400 ;
        RECT 487.600 83.600 488.400 84.400 ;
        RECT 503.600 91.600 504.400 92.400 ;
        RECT 502.000 83.600 502.800 84.400 ;
        RECT 524.400 91.600 525.200 92.400 ;
        RECT 532.400 93.600 533.200 94.400 ;
        RECT 561.200 93.600 562.000 94.400 ;
        RECT 550.000 92.200 550.800 93.000 ;
        RECT 562.800 90.200 563.600 91.000 ;
        RECT 545.200 87.600 546.000 88.400 ;
        RECT 567.600 89.600 568.400 90.400 ;
        RECT 583.600 93.000 584.400 93.800 ;
        RECT 574.000 89.600 574.800 90.400 ;
        RECT 593.200 92.600 594.000 93.400 ;
        RECT 607.600 97.600 608.400 98.400 ;
        RECT 578.800 91.600 579.600 92.400 ;
        RECT 588.400 91.600 589.200 92.400 ;
        RECT 585.200 88.800 586.000 89.600 ;
        RECT 590.000 87.600 590.800 88.400 ;
        RECT 586.800 86.200 587.600 87.000 ;
        RECT 583.600 84.200 584.400 85.000 ;
        RECT 585.200 84.200 586.000 85.000 ;
        RECT 590.000 86.200 590.800 87.000 ;
        RECT 593.200 86.200 594.000 87.000 ;
        RECT 594.800 84.200 595.600 85.000 ;
        RECT 596.400 84.200 597.200 85.000 ;
        RECT 598.000 84.200 598.800 85.000 ;
        RECT 6.000 69.600 6.800 70.400 ;
        RECT 14.000 69.600 14.800 70.400 ;
        RECT 15.600 67.600 16.400 68.400 ;
        RECT 25.200 69.600 26.000 70.400 ;
        RECT 28.400 69.600 29.200 70.400 ;
        RECT 30.000 69.600 30.800 70.400 ;
        RECT 33.200 69.600 34.000 70.400 ;
        RECT 62.000 73.600 62.800 74.400 ;
        RECT 41.200 69.600 42.000 70.400 ;
        RECT 36.400 67.600 37.200 68.400 ;
        RECT 9.200 63.600 10.000 64.400 ;
        RECT 42.800 67.600 43.600 68.400 ;
        RECT 44.400 66.200 45.200 67.000 ;
        RECT 65.200 69.600 66.000 70.400 ;
        RECT 79.600 73.600 80.400 74.400 ;
        RECT 71.600 69.600 72.400 70.400 ;
        RECT 79.600 69.600 80.400 70.400 ;
        RECT 82.800 69.600 83.600 70.400 ;
        RECT 84.400 69.600 85.200 70.400 ;
        RECT 49.200 65.600 50.000 66.400 ;
        RECT 81.200 67.600 82.000 68.400 ;
        RECT 100.400 77.600 101.200 78.400 ;
        RECT 98.800 65.600 99.600 66.400 ;
        RECT 103.600 77.600 104.400 78.400 ;
        RECT 102.000 65.600 102.800 66.400 ;
        RECT 106.800 77.600 107.600 78.400 ;
        RECT 105.200 65.600 106.000 66.400 ;
        RECT 122.800 72.400 123.600 73.200 ;
        RECT 126.000 71.000 126.800 71.800 ;
        RECT 127.600 77.600 128.400 78.400 ;
        RECT 126.000 66.200 126.800 67.000 ;
        RECT 108.400 63.600 109.200 64.400 ;
        RECT 132.400 77.600 133.200 78.400 ;
        RECT 129.200 65.600 130.000 66.400 ;
        RECT 130.800 65.600 131.600 66.400 ;
        RECT 175.600 77.600 176.400 78.400 ;
        RECT 150.000 69.600 150.800 70.400 ;
        RECT 186.800 77.600 187.600 78.400 ;
        RECT 158.000 66.200 158.800 67.000 ;
        RECT 178.800 69.600 179.600 70.400 ;
        RECT 186.800 69.600 187.600 70.400 ;
        RECT 190.000 69.600 190.800 70.400 ;
        RECT 191.600 69.600 192.400 70.400 ;
        RECT 137.200 63.600 138.000 64.400 ;
        RECT 162.800 65.600 163.600 66.400 ;
        RECT 188.400 67.600 189.200 68.400 ;
        RECT 222.000 75.000 222.800 75.800 ;
        RECT 218.800 73.600 219.600 74.400 ;
        RECT 223.600 72.400 224.400 73.200 ;
        RECT 201.200 67.600 202.000 68.400 ;
        RECT 202.800 67.600 203.600 68.400 ;
        RECT 212.400 68.200 213.200 69.000 ;
        RECT 222.000 68.600 222.800 69.400 ;
        RECT 217.200 67.600 218.000 68.400 ;
        RECT 212.400 64.200 213.200 65.000 ;
        RECT 214.000 64.200 214.800 65.000 ;
        RECT 215.600 64.200 216.400 65.000 ;
        RECT 218.800 64.200 219.600 65.000 ;
        RECT 222.000 64.200 222.800 65.000 ;
        RECT 223.600 64.200 224.400 65.000 ;
        RECT 225.200 64.200 226.000 65.000 ;
        RECT 226.800 64.200 227.600 65.000 ;
        RECT 247.600 69.600 248.400 70.400 ;
        RECT 258.800 73.600 259.600 74.400 ;
        RECT 270.000 74.400 270.800 75.200 ;
        RECT 273.200 75.000 274.000 75.800 ;
        RECT 268.400 72.400 269.200 73.200 ;
        RECT 236.400 63.600 237.200 64.400 ;
        RECT 278.000 67.600 278.800 68.400 ;
        RECT 274.800 65.600 275.600 66.400 ;
        RECT 268.400 64.200 269.200 65.000 ;
        RECT 270.000 64.200 270.800 65.000 ;
        RECT 271.600 64.200 272.400 65.000 ;
        RECT 273.200 64.200 274.000 65.000 ;
        RECT 276.400 64.200 277.200 65.000 ;
        RECT 279.600 64.200 280.400 65.000 ;
        RECT 281.200 64.200 282.000 65.000 ;
        RECT 282.800 64.200 283.600 65.000 ;
        RECT 292.400 67.600 293.200 68.400 ;
        RECT 303.600 73.600 304.400 74.400 ;
        RECT 314.800 74.400 315.600 75.200 ;
        RECT 318.000 75.000 318.800 75.800 ;
        RECT 313.200 72.400 314.000 73.200 ;
        RECT 311.600 69.600 312.400 70.400 ;
        RECT 322.800 67.600 323.600 68.400 ;
        RECT 319.600 65.600 320.400 66.400 ;
        RECT 338.800 69.600 339.600 70.400 ;
        RECT 345.400 71.800 346.200 72.600 ;
        RECT 346.600 69.800 347.400 70.600 ;
        RECT 313.200 64.200 314.000 65.000 ;
        RECT 314.800 64.200 315.600 65.000 ;
        RECT 316.400 64.200 317.200 65.000 ;
        RECT 318.000 64.200 318.800 65.000 ;
        RECT 321.200 64.200 322.000 65.000 ;
        RECT 324.400 64.200 325.200 65.000 ;
        RECT 326.000 64.200 326.800 65.000 ;
        RECT 327.600 64.200 328.400 65.000 ;
        RECT 358.000 69.600 358.800 70.400 ;
        RECT 345.400 66.200 346.200 67.000 ;
        RECT 353.200 67.600 354.000 68.400 ;
        RECT 356.400 67.600 357.200 68.400 ;
        RECT 359.600 67.600 360.400 68.400 ;
        RECT 361.200 67.600 362.000 68.400 ;
        RECT 366.000 65.600 366.800 66.400 ;
        RECT 378.800 69.600 379.600 70.400 ;
        RECT 372.400 65.600 373.200 66.400 ;
        RECT 370.800 63.600 371.600 64.400 ;
        RECT 390.000 69.600 390.800 70.400 ;
        RECT 396.200 71.800 397.000 72.600 ;
        RECT 396.200 66.200 397.000 67.000 ;
        RECT 410.800 69.600 411.600 70.400 ;
        RECT 417.200 69.600 418.000 70.400 ;
        RECT 406.000 67.600 406.800 68.400 ;
        RECT 407.600 67.600 408.400 68.400 ;
        RECT 428.400 77.600 429.200 78.400 ;
        RECT 426.800 71.600 427.600 72.400 ;
        RECT 425.200 67.600 426.000 68.400 ;
        RECT 423.600 63.600 424.400 64.400 ;
        RECT 438.000 69.600 438.800 70.400 ;
        RECT 441.200 69.600 442.000 70.400 ;
        RECT 455.600 75.600 456.400 76.400 ;
        RECT 463.600 73.600 464.400 74.400 ;
        RECT 449.200 69.600 450.000 70.400 ;
        RECT 434.800 63.600 435.600 64.400 ;
        RECT 450.800 67.600 451.600 68.400 ;
        RECT 478.000 72.400 478.800 73.200 ;
        RECT 481.200 71.000 482.000 71.800 ;
        RECT 484.400 69.600 485.200 70.400 ;
        RECT 514.800 75.600 515.600 76.400 ;
        RECT 492.400 69.600 493.200 70.400 ;
        RECT 505.200 71.600 506.000 72.400 ;
        RECT 505.200 69.600 506.000 70.400 ;
        RECT 481.200 66.200 482.000 67.000 ;
        RECT 494.000 67.600 494.800 68.400 ;
        RECT 506.800 67.600 507.600 68.400 ;
        RECT 529.200 72.400 530.000 73.200 ;
        RECT 532.400 71.000 533.200 71.800 ;
        RECT 535.600 69.600 536.400 70.400 ;
        RECT 487.600 63.600 488.400 64.400 ;
        RECT 513.200 63.600 514.000 64.400 ;
        RECT 540.400 67.600 541.200 68.400 ;
        RECT 532.400 66.200 533.200 67.000 ;
        RECT 548.400 67.600 549.200 68.400 ;
        RECT 575.600 73.600 576.400 74.400 ;
        RECT 564.400 69.600 565.200 70.400 ;
        RECT 596.400 73.600 597.200 74.400 ;
        RECT 575.600 69.600 576.400 70.400 ;
        RECT 553.200 63.600 554.000 64.400 ;
        RECT 577.200 67.600 578.000 68.400 ;
        RECT 580.400 67.600 581.200 68.400 ;
        RECT 578.800 66.200 579.600 67.000 ;
        RECT 599.600 77.600 600.400 78.400 ;
        RECT 598.000 67.600 598.800 68.400 ;
        RECT 606.000 69.600 606.800 70.400 ;
        RECT 607.600 67.600 608.400 68.400 ;
        RECT 602.800 63.600 603.600 64.400 ;
        RECT 9.200 53.000 10.000 53.800 ;
        RECT 18.800 52.600 19.600 53.400 ;
        RECT 33.200 57.600 34.000 58.400 ;
        RECT 44.400 57.600 45.200 58.400 ;
        RECT 49.200 57.600 50.000 58.400 ;
        RECT 7.600 51.600 8.400 52.400 ;
        RECT 10.800 48.800 11.600 49.600 ;
        RECT 15.600 47.600 16.400 48.400 ;
        RECT 12.400 46.200 13.200 47.000 ;
        RECT 9.200 44.200 10.000 45.000 ;
        RECT 10.800 44.200 11.600 45.000 ;
        RECT 15.600 46.200 16.400 47.000 ;
        RECT 18.800 46.200 19.600 47.000 ;
        RECT 20.400 44.200 21.200 45.000 ;
        RECT 22.000 44.200 22.800 45.000 ;
        RECT 23.600 44.200 24.400 45.000 ;
        RECT 41.200 49.600 42.000 50.400 ;
        RECT 73.200 57.600 74.000 58.400 ;
        RECT 60.400 53.600 61.200 54.400 ;
        RECT 63.600 51.600 64.400 52.400 ;
        RECT 71.600 49.600 72.400 50.400 ;
        RECT 97.200 57.600 98.000 58.400 ;
        RECT 87.600 51.600 88.400 52.400 ;
        RECT 90.800 43.600 91.600 44.400 ;
        RECT 100.400 57.600 101.200 58.400 ;
        RECT 111.600 53.600 112.400 54.400 ;
        RECT 100.400 43.600 101.200 44.400 ;
        RECT 143.600 55.600 144.400 56.400 ;
        RECT 118.000 43.600 118.800 44.400 ;
        RECT 129.200 51.600 130.000 52.400 ;
        RECT 140.400 51.600 141.200 52.400 ;
        RECT 134.000 43.600 134.800 44.400 ;
        RECT 166.000 53.600 166.800 54.400 ;
        RECT 156.400 51.600 157.200 52.400 ;
        RECT 178.800 53.600 179.600 54.400 ;
        RECT 188.400 53.000 189.200 53.800 ;
        RECT 198.000 52.600 198.800 53.400 ;
        RECT 212.400 57.600 213.200 58.400 ;
        RECT 185.200 51.600 186.000 52.400 ;
        RECT 204.400 51.600 205.200 52.400 ;
        RECT 190.000 48.800 190.800 49.600 ;
        RECT 194.800 47.600 195.600 48.400 ;
        RECT 191.600 46.200 192.400 47.000 ;
        RECT 188.400 44.200 189.200 45.000 ;
        RECT 190.000 44.200 190.800 45.000 ;
        RECT 194.800 46.200 195.600 47.000 ;
        RECT 198.000 46.200 198.800 47.000 ;
        RECT 199.600 44.200 200.400 45.000 ;
        RECT 201.200 44.200 202.000 45.000 ;
        RECT 202.800 44.200 203.600 45.000 ;
        RECT 220.400 55.600 221.200 56.400 ;
        RECT 218.800 49.600 219.600 50.400 ;
        RECT 217.200 43.600 218.000 44.400 ;
        RECT 226.800 49.600 227.600 50.400 ;
        RECT 231.600 49.600 232.400 50.400 ;
        RECT 236.400 49.600 237.200 50.400 ;
        RECT 250.800 53.000 251.600 53.800 ;
        RECT 260.400 52.600 261.200 53.400 ;
        RECT 274.800 55.600 275.600 56.400 ;
        RECT 246.000 51.600 246.800 52.400 ;
        RECT 252.400 48.800 253.200 49.600 ;
        RECT 257.200 47.600 258.000 48.400 ;
        RECT 254.000 46.200 254.800 47.000 ;
        RECT 250.800 44.200 251.600 45.000 ;
        RECT 252.400 44.200 253.200 45.000 ;
        RECT 257.200 46.200 258.000 47.000 ;
        RECT 260.400 46.200 261.200 47.000 ;
        RECT 262.000 44.200 262.800 45.000 ;
        RECT 263.600 44.200 264.400 45.000 ;
        RECT 265.200 44.200 266.000 45.000 ;
        RECT 282.800 49.600 283.600 50.400 ;
        RECT 303.600 53.000 304.400 53.800 ;
        RECT 274.800 43.600 275.600 44.400 ;
        RECT 313.200 52.600 314.000 53.400 ;
        RECT 297.200 51.600 298.000 52.400 ;
        RECT 319.600 51.600 320.400 52.400 ;
        RECT 353.200 57.600 354.000 58.400 ;
        RECT 305.200 48.800 306.000 49.600 ;
        RECT 310.000 47.600 310.800 48.400 ;
        RECT 287.600 43.600 288.400 44.400 ;
        RECT 306.800 46.200 307.600 47.000 ;
        RECT 303.600 44.200 304.400 45.000 ;
        RECT 305.200 44.200 306.000 45.000 ;
        RECT 310.000 46.200 310.800 47.000 ;
        RECT 313.200 46.200 314.000 47.000 ;
        RECT 314.800 44.200 315.600 45.000 ;
        RECT 316.400 44.200 317.200 45.000 ;
        RECT 318.000 44.200 318.800 45.000 ;
        RECT 327.600 49.600 328.400 50.400 ;
        RECT 351.600 53.600 352.400 54.400 ;
        RECT 367.600 57.600 368.400 58.400 ;
        RECT 370.800 57.600 371.600 58.400 ;
        RECT 362.800 53.600 363.600 54.400 ;
        RECT 343.600 49.600 344.400 50.400 ;
        RECT 361.200 49.600 362.000 50.400 ;
        RECT 380.400 53.000 381.200 53.800 ;
        RECT 390.000 52.600 390.800 53.400 ;
        RECT 404.400 57.600 405.200 58.400 ;
        RECT 375.600 51.600 376.400 52.400 ;
        RECT 385.200 51.600 386.000 52.400 ;
        RECT 425.200 57.600 426.000 58.400 ;
        RECT 409.200 53.600 410.000 54.400 ;
        RECT 382.000 48.800 382.800 49.600 ;
        RECT 386.800 47.600 387.600 48.400 ;
        RECT 383.600 46.200 384.400 47.000 ;
        RECT 380.400 44.200 381.200 45.000 ;
        RECT 382.000 44.200 382.800 45.000 ;
        RECT 386.800 46.200 387.600 47.000 ;
        RECT 390.000 46.200 390.800 47.000 ;
        RECT 391.600 44.200 392.400 45.000 ;
        RECT 393.200 44.200 394.000 45.000 ;
        RECT 394.800 44.200 395.600 45.000 ;
        RECT 407.600 50.200 408.400 51.000 ;
        RECT 434.800 57.600 435.600 58.400 ;
        RECT 452.400 55.600 453.200 56.400 ;
        RECT 434.800 49.600 435.600 50.400 ;
        RECT 439.600 49.600 440.400 50.400 ;
        RECT 500.400 57.600 501.200 58.400 ;
        RECT 484.400 53.600 485.200 54.400 ;
        RECT 503.600 57.600 504.400 58.400 ;
        RECT 479.600 51.600 480.400 52.400 ;
        RECT 487.600 51.800 488.400 52.600 ;
        RECT 482.800 50.200 483.600 51.000 ;
        RECT 478.000 43.600 478.800 44.400 ;
        RECT 516.400 53.600 517.200 54.400 ;
        RECT 511.600 51.600 512.400 52.400 ;
        RECT 543.600 57.600 544.400 58.400 ;
        RECT 522.800 51.600 523.600 52.400 ;
        RECT 510.000 43.600 510.800 44.400 ;
        RECT 524.400 49.600 525.200 50.400 ;
        RECT 535.600 49.600 536.400 50.400 ;
        RECT 578.800 57.600 579.600 58.400 ;
        RECT 559.600 53.600 560.400 54.400 ;
        RECT 548.400 52.200 549.200 53.000 ;
        RECT 575.600 53.600 576.400 54.400 ;
        RECT 540.400 47.600 541.200 48.400 ;
        RECT 561.200 50.200 562.000 51.000 ;
        RECT 564.400 43.600 565.200 44.400 ;
        RECT 594.800 55.600 595.600 56.400 ;
        RECT 596.400 54.200 597.200 55.000 ;
        RECT 586.800 51.600 587.600 52.400 ;
        RECT 598.000 51.600 598.800 52.400 ;
        RECT 590.000 46.800 590.800 47.600 ;
        RECT 593.200 46.200 594.000 47.000 ;
        RECT 588.400 44.200 589.200 45.000 ;
        RECT 590.000 44.200 590.800 45.000 ;
        RECT 591.600 44.200 592.400 45.000 ;
        RECT 596.400 46.200 597.200 47.000 ;
        RECT 599.600 46.200 600.400 47.000 ;
        RECT 601.200 44.200 602.000 45.000 ;
        RECT 602.800 44.200 603.600 45.000 ;
        RECT 4.400 29.600 5.200 30.400 ;
        RECT 23.600 35.000 24.400 35.800 ;
        RECT 20.400 33.600 21.200 34.400 ;
        RECT 38.000 37.600 38.800 38.400 ;
        RECT 25.200 32.400 26.000 33.200 ;
        RECT 30.000 29.600 30.800 30.400 ;
        RECT 14.000 28.200 14.800 29.000 ;
        RECT 23.600 28.600 24.400 29.400 ;
        RECT 18.800 27.600 19.600 28.400 ;
        RECT 14.000 24.200 14.800 25.000 ;
        RECT 15.600 24.200 16.400 25.000 ;
        RECT 17.200 24.200 18.000 25.000 ;
        RECT 20.400 24.200 21.200 25.000 ;
        RECT 23.600 24.200 24.400 25.000 ;
        RECT 25.200 24.200 26.000 25.000 ;
        RECT 26.800 24.200 27.600 25.000 ;
        RECT 28.400 24.200 29.200 25.000 ;
        RECT 44.400 29.600 45.200 30.400 ;
        RECT 52.400 29.600 53.200 30.400 ;
        RECT 63.600 35.600 64.400 36.400 ;
        RECT 60.400 29.600 61.200 30.400 ;
        RECT 62.000 27.600 62.800 28.400 ;
        RECT 78.000 32.400 78.800 33.200 ;
        RECT 81.200 31.000 82.000 31.800 ;
        RECT 113.200 37.600 114.000 38.400 ;
        RECT 84.400 29.600 85.200 30.400 ;
        RECT 92.400 29.600 93.200 30.400 ;
        RECT 102.000 29.600 102.800 30.400 ;
        RECT 57.200 23.600 58.000 24.400 ;
        RECT 76.400 25.600 77.200 26.400 ;
        RECT 81.200 26.200 82.000 27.000 ;
        RECT 94.000 27.600 94.800 28.400 ;
        RECT 95.600 26.200 96.400 27.000 ;
        RECT 116.400 29.600 117.200 30.400 ;
        RECT 124.400 29.600 125.200 30.400 ;
        RECT 140.400 37.600 141.200 38.400 ;
        RECT 137.200 29.600 138.000 30.400 ;
        RECT 126.000 27.600 126.800 28.400 ;
        RECT 138.800 27.600 139.600 28.400 ;
        RECT 154.800 32.400 155.600 33.200 ;
        RECT 158.000 31.000 158.800 31.800 ;
        RECT 132.400 23.600 133.200 24.400 ;
        RECT 158.000 26.200 158.800 27.000 ;
        RECT 191.600 34.400 192.400 35.200 ;
        RECT 194.800 35.000 195.600 35.800 ;
        RECT 190.000 32.400 190.800 33.200 ;
        RECT 180.200 29.600 181.000 30.400 ;
        RECT 188.400 29.600 189.200 30.400 ;
        RECT 172.400 23.600 173.200 24.400 ;
        RECT 199.600 27.600 200.400 28.400 ;
        RECT 196.400 25.600 197.200 26.400 ;
        RECT 190.000 24.200 190.800 25.000 ;
        RECT 191.600 24.200 192.400 25.000 ;
        RECT 193.200 24.200 194.000 25.000 ;
        RECT 194.800 24.200 195.600 25.000 ;
        RECT 198.000 24.200 198.800 25.000 ;
        RECT 201.200 24.200 202.000 25.000 ;
        RECT 202.800 24.200 203.600 25.000 ;
        RECT 204.400 24.200 205.200 25.000 ;
        RECT 220.400 29.600 221.200 30.400 ;
        RECT 215.600 25.600 216.400 26.400 ;
        RECT 222.000 27.600 222.800 28.400 ;
        RECT 228.400 27.600 229.200 28.400 ;
        RECT 217.200 23.600 218.000 24.400 ;
        RECT 223.600 23.600 224.400 24.400 ;
        RECT 250.800 35.000 251.600 35.800 ;
        RECT 247.600 33.600 248.400 34.400 ;
        RECT 252.400 32.400 253.200 33.200 ;
        RECT 270.000 37.600 270.800 38.400 ;
        RECT 257.200 29.600 258.000 30.400 ;
        RECT 241.200 28.200 242.000 29.000 ;
        RECT 250.800 28.600 251.600 29.400 ;
        RECT 231.600 25.600 232.400 26.400 ;
        RECT 246.000 27.600 246.800 28.400 ;
        RECT 241.200 24.200 242.000 25.000 ;
        RECT 242.800 24.200 243.600 25.000 ;
        RECT 244.400 24.200 245.200 25.000 ;
        RECT 247.600 24.200 248.400 25.000 ;
        RECT 250.800 24.200 251.600 25.000 ;
        RECT 252.400 24.200 253.200 25.000 ;
        RECT 254.000 24.200 254.800 25.000 ;
        RECT 255.600 24.200 256.400 25.000 ;
        RECT 265.200 23.600 266.000 24.400 ;
        RECT 289.200 35.000 290.000 35.800 ;
        RECT 286.000 33.600 286.800 34.400 ;
        RECT 290.800 32.400 291.600 33.200 ;
        RECT 313.200 37.600 314.000 38.400 ;
        RECT 295.600 29.600 296.400 30.400 ;
        RECT 279.600 28.200 280.400 29.000 ;
        RECT 289.200 28.600 290.000 29.400 ;
        RECT 284.400 27.600 285.200 28.400 ;
        RECT 303.800 27.600 304.600 28.400 ;
        RECT 279.600 24.200 280.400 25.000 ;
        RECT 281.200 24.200 282.000 25.000 ;
        RECT 282.800 24.200 283.600 25.000 ;
        RECT 286.000 24.200 286.800 25.000 ;
        RECT 289.200 24.200 290.000 25.000 ;
        RECT 290.800 24.200 291.600 25.000 ;
        RECT 292.400 24.200 293.200 25.000 ;
        RECT 294.000 24.200 294.800 25.000 ;
        RECT 316.400 31.800 317.200 32.600 ;
        RECT 330.800 37.600 331.600 38.400 ;
        RECT 316.400 26.200 317.200 27.000 ;
        RECT 326.000 29.600 326.800 30.400 ;
        RECT 327.600 29.600 328.400 30.400 ;
        RECT 337.400 31.800 338.200 32.600 ;
        RECT 351.600 37.600 352.400 38.400 ;
        RECT 356.400 37.600 357.200 38.400 ;
        RECT 350.000 33.600 350.800 34.400 ;
        RECT 338.600 29.800 339.400 30.600 ;
        RECT 346.800 31.600 347.600 32.400 ;
        RECT 321.200 26.400 322.000 27.200 ;
        RECT 370.800 34.400 371.600 35.200 ;
        RECT 374.000 35.000 374.800 35.800 ;
        RECT 369.200 32.400 370.000 33.200 ;
        RECT 337.400 26.200 338.200 27.000 ;
        RECT 345.200 27.600 346.000 28.400 ;
        RECT 353.200 25.600 354.000 26.400 ;
        RECT 367.600 29.600 368.400 30.400 ;
        RECT 359.600 25.600 360.400 26.400 ;
        RECT 378.800 27.600 379.600 28.400 ;
        RECT 375.600 25.600 376.400 26.400 ;
        RECT 369.200 24.200 370.000 25.000 ;
        RECT 370.800 24.200 371.600 25.000 ;
        RECT 372.400 24.200 373.200 25.000 ;
        RECT 374.000 24.200 374.800 25.000 ;
        RECT 377.200 24.200 378.000 25.000 ;
        RECT 380.400 24.200 381.200 25.000 ;
        RECT 382.000 24.200 382.800 25.000 ;
        RECT 383.600 24.200 384.400 25.000 ;
        RECT 418.800 37.600 419.600 38.400 ;
        RECT 431.600 37.600 432.400 38.400 ;
        RECT 430.000 33.600 430.800 34.400 ;
        RECT 423.600 29.600 424.400 30.400 ;
        RECT 444.400 37.600 445.200 38.400 ;
        RECT 442.800 33.600 443.600 34.400 ;
        RECT 431.600 29.600 432.400 30.400 ;
        RECT 438.000 29.600 438.800 30.400 ;
        RECT 476.400 37.600 477.200 38.400 ;
        RECT 444.400 29.600 445.200 30.400 ;
        RECT 450.800 29.600 451.600 30.400 ;
        RECT 465.200 29.600 466.000 30.400 ;
        RECT 394.800 23.600 395.600 24.400 ;
        RECT 425.200 27.600 426.000 28.400 ;
        RECT 439.600 27.600 440.400 28.400 ;
        RECT 449.200 27.600 450.000 28.400 ;
        RECT 452.400 27.600 453.200 28.400 ;
        RECT 458.800 26.200 459.600 27.000 ;
        RECT 508.400 37.600 509.200 38.400 ;
        RECT 481.200 29.600 482.000 30.400 ;
        RECT 497.200 29.600 498.000 30.400 ;
        RECT 489.200 27.600 490.000 28.400 ;
        RECT 490.800 26.200 491.600 27.000 ;
        RECT 513.200 29.600 514.000 30.400 ;
        RECT 537.200 37.600 538.000 38.400 ;
        RECT 519.600 29.600 520.400 30.400 ;
        RECT 521.200 27.600 522.000 28.400 ;
        RECT 543.600 33.600 544.400 34.400 ;
        RECT 548.400 29.600 549.200 30.400 ;
        RECT 556.400 29.600 557.200 30.400 ;
        RECT 562.800 29.600 563.600 30.400 ;
        RECT 538.800 25.600 539.600 26.400 ;
        RECT 545.200 27.600 546.000 28.400 ;
        RECT 551.600 27.600 552.400 28.400 ;
        RECT 558.000 27.600 558.800 28.400 ;
        RECT 561.200 27.600 562.000 28.400 ;
        RECT 570.800 35.600 571.600 36.400 ;
        RECT 553.200 23.600 554.000 24.400 ;
        RECT 582.000 34.400 582.800 35.200 ;
        RECT 585.200 35.000 586.000 35.800 ;
        RECT 604.400 37.600 605.200 38.400 ;
        RECT 580.400 32.400 581.200 33.200 ;
        RECT 590.000 27.600 590.800 28.400 ;
        RECT 586.800 25.600 587.600 26.400 ;
        RECT 580.400 24.200 581.200 25.000 ;
        RECT 582.000 24.200 582.800 25.000 ;
        RECT 583.600 24.200 584.400 25.000 ;
        RECT 585.200 24.200 586.000 25.000 ;
        RECT 588.400 24.200 589.200 25.000 ;
        RECT 591.600 24.200 592.400 25.000 ;
        RECT 593.200 24.200 594.000 25.000 ;
        RECT 594.800 24.200 595.600 25.000 ;
        RECT 9.200 13.000 10.000 13.800 ;
        RECT 18.800 12.600 19.600 13.400 ;
        RECT 33.200 15.600 34.000 16.400 ;
        RECT 7.600 11.600 8.400 12.400 ;
        RECT 70.000 17.600 70.800 18.400 ;
        RECT 10.800 8.800 11.600 9.600 ;
        RECT 15.600 7.600 16.400 8.400 ;
        RECT 12.400 6.200 13.200 7.000 ;
        RECT 9.200 4.200 10.000 5.000 ;
        RECT 10.800 4.200 11.600 5.000 ;
        RECT 15.600 6.200 16.400 7.000 ;
        RECT 18.800 6.200 19.600 7.000 ;
        RECT 20.400 4.200 21.200 5.000 ;
        RECT 22.000 4.200 22.800 5.000 ;
        RECT 23.600 4.200 24.400 5.000 ;
        RECT 41.200 9.600 42.000 10.400 ;
        RECT 54.000 13.600 54.800 14.400 ;
        RECT 73.200 17.600 74.000 18.400 ;
        RECT 57.200 11.800 58.000 12.600 ;
        RECT 52.400 10.200 53.200 11.000 ;
        RECT 90.800 17.600 91.600 18.400 ;
        RECT 82.800 13.600 83.600 14.400 ;
        RECT 100.400 13.600 101.200 14.400 ;
        RECT 110.000 17.600 110.800 18.400 ;
        RECT 95.600 12.200 96.400 13.000 ;
        RECT 130.800 17.600 131.600 18.400 ;
        RECT 146.800 17.600 147.600 18.400 ;
        RECT 114.800 12.200 115.600 13.000 ;
        RECT 122.800 11.800 123.600 12.600 ;
        RECT 108.400 10.200 109.200 11.000 ;
        RECT 127.600 10.200 128.400 11.000 ;
        RECT 134.000 11.600 134.800 12.400 ;
        RECT 162.800 15.600 163.600 16.400 ;
        RECT 164.400 14.200 165.200 15.000 ;
        RECT 154.800 11.600 155.600 12.400 ;
        RECT 177.200 11.600 178.000 12.400 ;
        RECT 158.000 6.800 158.800 7.600 ;
        RECT 161.200 6.200 162.000 7.000 ;
        RECT 156.400 4.200 157.200 5.000 ;
        RECT 158.000 4.200 158.800 5.000 ;
        RECT 159.600 4.200 160.400 5.000 ;
        RECT 164.400 6.200 165.200 7.000 ;
        RECT 167.600 6.200 168.400 7.000 ;
        RECT 188.400 13.000 189.200 13.800 ;
        RECT 198.000 12.600 198.800 13.400 ;
        RECT 183.600 11.600 184.400 12.400 ;
        RECT 204.400 11.600 205.200 12.400 ;
        RECT 228.400 13.000 229.200 13.800 ;
        RECT 190.000 8.800 190.800 9.600 ;
        RECT 194.800 7.600 195.600 8.400 ;
        RECT 169.200 4.200 170.000 5.000 ;
        RECT 170.800 4.200 171.600 5.000 ;
        RECT 191.600 6.200 192.400 7.000 ;
        RECT 188.400 4.200 189.200 5.000 ;
        RECT 190.000 4.200 190.800 5.000 ;
        RECT 194.800 6.200 195.600 7.000 ;
        RECT 198.000 6.200 198.800 7.000 ;
        RECT 199.600 4.200 200.400 5.000 ;
        RECT 201.200 4.200 202.000 5.000 ;
        RECT 202.800 4.200 203.600 5.000 ;
        RECT 238.000 12.600 238.800 13.400 ;
        RECT 252.400 17.600 253.200 18.400 ;
        RECT 223.600 11.600 224.400 12.400 ;
        RECT 278.000 13.000 278.800 13.800 ;
        RECT 230.000 8.800 230.800 9.600 ;
        RECT 234.800 7.600 235.600 8.400 ;
        RECT 231.600 6.200 232.400 7.000 ;
        RECT 228.400 4.200 229.200 5.000 ;
        RECT 230.000 4.200 230.800 5.000 ;
        RECT 234.800 6.200 235.600 7.000 ;
        RECT 238.000 6.200 238.800 7.000 ;
        RECT 239.600 4.200 240.400 5.000 ;
        RECT 241.200 4.200 242.000 5.000 ;
        RECT 242.800 4.200 243.600 5.000 ;
        RECT 287.600 12.600 288.400 13.400 ;
        RECT 273.200 11.600 274.000 12.400 ;
        RECT 322.800 13.000 323.600 13.800 ;
        RECT 279.600 8.800 280.400 9.600 ;
        RECT 284.400 7.600 285.200 8.400 ;
        RECT 281.200 6.200 282.000 7.000 ;
        RECT 278.000 4.200 278.800 5.000 ;
        RECT 279.600 4.200 280.400 5.000 ;
        RECT 284.400 6.200 285.200 7.000 ;
        RECT 287.600 6.200 288.400 7.000 ;
        RECT 289.200 4.200 290.000 5.000 ;
        RECT 290.800 4.200 291.600 5.000 ;
        RECT 292.400 4.200 293.200 5.000 ;
        RECT 332.400 12.600 333.200 13.400 ;
        RECT 346.800 17.600 347.600 18.400 ;
        RECT 318.000 11.600 318.800 12.400 ;
        RECT 324.400 8.800 325.200 9.600 ;
        RECT 329.200 7.600 330.000 8.400 ;
        RECT 326.000 6.200 326.800 7.000 ;
        RECT 322.800 4.200 323.600 5.000 ;
        RECT 324.400 4.200 325.200 5.000 ;
        RECT 329.200 6.200 330.000 7.000 ;
        RECT 332.400 6.200 333.200 7.000 ;
        RECT 334.000 4.200 334.800 5.000 ;
        RECT 335.600 4.200 336.400 5.000 ;
        RECT 337.200 4.200 338.000 5.000 ;
        RECT 372.400 13.000 373.200 13.800 ;
        RECT 382.000 12.600 382.800 13.400 ;
        RECT 396.400 17.600 397.200 18.400 ;
        RECT 367.600 11.600 368.400 12.400 ;
        RECT 374.000 8.800 374.800 9.600 ;
        RECT 378.800 7.600 379.600 8.400 ;
        RECT 375.600 6.200 376.400 7.000 ;
        RECT 372.400 4.200 373.200 5.000 ;
        RECT 374.000 4.200 374.800 5.000 ;
        RECT 378.800 6.200 379.600 7.000 ;
        RECT 382.000 6.200 382.800 7.000 ;
        RECT 383.600 4.200 384.400 5.000 ;
        RECT 385.200 4.200 386.000 5.000 ;
        RECT 386.800 4.200 387.600 5.000 ;
        RECT 404.400 10.200 405.200 11.000 ;
        RECT 433.200 17.600 434.000 18.400 ;
        RECT 422.000 7.600 422.800 8.400 ;
        RECT 430.000 11.600 430.800 12.400 ;
        RECT 478.000 15.600 478.800 16.400 ;
        RECT 438.000 12.200 438.800 13.000 ;
        RECT 446.000 11.800 446.800 12.600 ;
        RECT 450.800 10.200 451.600 11.000 ;
        RECT 474.800 11.600 475.600 12.400 ;
        RECT 487.600 13.600 488.400 14.400 ;
        RECT 502.000 13.600 502.800 14.400 ;
        RECT 500.400 11.800 501.200 12.600 ;
        RECT 495.600 10.200 496.400 11.000 ;
        RECT 538.800 17.600 539.600 18.400 ;
        RECT 543.600 17.600 544.400 18.400 ;
        RECT 529.200 13.600 530.000 14.400 ;
        RECT 518.000 9.600 518.800 10.400 ;
        RECT 513.200 7.600 514.000 8.400 ;
        RECT 542.000 11.600 542.800 12.400 ;
        RECT 562.800 17.600 563.600 18.400 ;
        RECT 559.600 13.600 560.400 14.400 ;
        RECT 548.400 12.200 549.200 13.000 ;
        RECT 561.200 10.200 562.000 11.000 ;
        RECT 570.800 17.600 571.600 18.400 ;
        RECT 574.000 17.600 574.800 18.400 ;
        RECT 590.000 15.600 590.800 16.400 ;
        RECT 591.600 14.200 592.400 15.000 ;
        RECT 601.200 11.600 602.000 12.400 ;
        RECT 570.800 9.600 571.600 10.400 ;
        RECT 585.200 6.800 586.000 7.600 ;
        RECT 588.400 6.200 589.200 7.000 ;
        RECT 583.600 4.200 584.400 5.000 ;
        RECT 585.200 4.200 586.000 5.000 ;
        RECT 586.800 4.200 587.600 5.000 ;
        RECT 591.600 6.200 592.400 7.000 ;
        RECT 594.800 6.200 595.600 7.000 ;
        RECT 607.600 17.600 608.400 18.400 ;
        RECT 596.400 4.200 597.200 5.000 ;
        RECT 598.000 4.200 598.800 5.000 ;
      LAYER metal2 ;
        RECT 6.000 549.600 6.800 550.400 ;
        RECT 2.800 547.600 3.600 548.400 ;
        RECT 2.800 545.600 3.600 546.400 ;
        RECT 2.900 528.400 3.500 545.600 ;
        RECT 6.100 532.400 6.700 549.600 ;
        RECT 12.400 544.200 13.200 557.800 ;
        RECT 14.000 544.200 14.800 557.800 ;
        RECT 15.600 544.200 16.400 555.800 ;
        RECT 17.200 547.600 18.000 548.400 ;
        RECT 17.200 545.600 18.000 546.400 ;
        RECT 6.000 531.600 6.800 532.400 ;
        RECT 2.800 527.600 3.600 528.400 ;
        RECT 1.200 506.200 2.000 511.800 ;
        RECT 1.200 503.600 2.000 504.400 ;
        RECT 1.300 498.400 1.900 503.600 ;
        RECT 1.200 497.600 2.000 498.400 ;
        RECT 1.200 491.600 2.000 492.400 ;
        RECT 1.300 490.400 1.900 491.600 ;
        RECT 1.200 489.600 2.000 490.400 ;
        RECT 1.200 466.200 2.000 471.800 ;
        RECT 1.200 443.600 2.000 444.400 ;
        RECT 1.300 432.400 1.900 443.600 ;
        RECT 1.200 431.600 2.000 432.400 ;
        RECT 2.900 430.400 3.500 527.600 ;
        RECT 9.200 524.200 10.000 537.800 ;
        RECT 10.800 524.200 11.600 537.800 ;
        RECT 12.400 526.200 13.200 537.800 ;
        RECT 14.000 533.600 14.800 534.400 ;
        RECT 15.600 526.200 16.400 537.800 ;
        RECT 17.300 536.400 17.900 545.600 ;
        RECT 18.800 544.200 19.600 555.800 ;
        RECT 20.400 545.600 21.200 546.400 ;
        RECT 22.000 544.200 22.800 555.800 ;
        RECT 23.600 544.200 24.400 557.800 ;
        RECT 25.200 544.200 26.000 557.800 ;
        RECT 26.800 544.200 27.600 557.800 ;
        RECT 47.600 553.600 48.400 554.400 ;
        RECT 63.600 553.600 64.400 554.400 ;
        RECT 63.700 552.400 64.300 553.600 ;
        RECT 57.200 551.600 58.000 552.400 ;
        RECT 60.400 551.600 61.200 552.400 ;
        RECT 63.600 551.600 64.400 552.400 ;
        RECT 28.400 549.600 29.200 550.400 ;
        RECT 33.200 549.600 34.000 550.400 ;
        RECT 44.400 549.600 45.200 550.400 ;
        RECT 52.400 549.600 53.200 550.400 ;
        RECT 60.400 549.600 61.200 550.400 ;
        RECT 74.800 549.600 75.600 550.400 ;
        RECT 28.500 546.400 29.100 549.600 ;
        RECT 28.400 545.600 29.200 546.400 ;
        RECT 33.300 538.400 33.900 549.600 ;
        RECT 44.400 547.600 45.200 548.400 ;
        RECT 38.000 545.600 38.800 546.400 ;
        RECT 17.200 535.600 18.000 536.400 ;
        RECT 4.400 504.200 5.200 515.800 ;
        RECT 6.000 509.400 6.800 510.200 ;
        RECT 12.400 509.600 13.200 510.400 ;
        RECT 6.100 504.400 6.700 509.400 ;
        RECT 12.500 508.400 13.100 509.600 ;
        RECT 12.400 507.600 13.200 508.400 ;
        RECT 6.000 503.600 6.800 504.400 ;
        RECT 6.000 493.600 6.800 494.400 ;
        RECT 6.100 486.400 6.700 493.600 ;
        RECT 9.200 491.600 10.000 492.400 ;
        RECT 6.000 485.600 6.800 486.400 ;
        RECT 4.400 464.200 5.200 475.800 ;
        RECT 7.600 469.600 8.400 470.400 ;
        RECT 6.000 446.200 6.800 457.800 ;
        RECT 9.300 448.400 9.900 491.600 ;
        RECT 12.500 470.400 13.100 507.600 ;
        RECT 14.000 504.200 14.800 515.800 ;
        RECT 17.300 508.400 17.900 535.600 ;
        RECT 18.800 526.200 19.600 537.800 ;
        RECT 20.400 524.200 21.200 537.800 ;
        RECT 22.000 524.200 22.800 537.800 ;
        RECT 23.600 524.200 24.400 537.800 ;
        RECT 33.200 537.600 34.000 538.400 ;
        RECT 33.300 530.400 33.900 537.600 ;
        RECT 34.800 535.600 35.600 536.400 ;
        RECT 34.900 530.400 35.500 535.600 ;
        RECT 36.400 533.600 37.200 534.400 ;
        RECT 38.100 532.300 38.700 545.600 ;
        RECT 42.800 535.600 43.600 536.400 ;
        RECT 41.200 533.600 42.000 534.400 ;
        RECT 39.600 532.300 40.400 532.400 ;
        RECT 38.100 531.700 40.400 532.300 ;
        RECT 39.600 531.600 40.400 531.700 ;
        RECT 33.200 529.600 34.000 530.400 ;
        RECT 34.800 529.600 35.600 530.400 ;
        RECT 41.300 522.400 41.900 533.600 ;
        RECT 44.500 532.400 45.100 547.600 ;
        RECT 46.000 543.600 46.800 544.400 ;
        RECT 46.100 536.400 46.700 543.600 ;
        RECT 46.000 535.600 46.800 536.400 ;
        RECT 46.000 533.600 46.800 534.400 ;
        RECT 52.500 532.400 53.100 549.600 ;
        RECT 57.200 547.600 58.000 548.400 ;
        RECT 58.800 547.600 59.600 548.400 ;
        RECT 58.900 546.300 59.500 547.600 ;
        RECT 57.300 545.700 59.500 546.300 ;
        RECT 57.300 534.400 57.900 545.700 ;
        RECT 55.600 533.600 56.400 534.400 ;
        RECT 57.200 533.600 58.000 534.400 ;
        RECT 44.400 531.600 45.200 532.400 ;
        RECT 52.400 531.600 53.200 532.400 ;
        RECT 42.800 529.600 43.600 530.400 ;
        RECT 52.500 528.400 53.100 531.600 ;
        RECT 55.600 529.600 56.400 530.400 ;
        RECT 52.400 527.600 53.200 528.400 ;
        RECT 57.300 522.400 57.900 533.600 ;
        RECT 58.800 532.300 59.600 532.400 ;
        RECT 60.500 532.300 61.100 549.600 ;
        RECT 74.900 546.400 75.500 549.600 ;
        RECT 74.800 545.600 75.600 546.400 ;
        RECT 76.400 544.200 77.200 557.800 ;
        RECT 78.000 544.200 78.800 557.800 ;
        RECT 79.600 544.200 80.400 557.800 ;
        RECT 81.200 544.200 82.000 555.800 ;
        RECT 82.800 545.600 83.600 546.400 ;
        RECT 82.900 542.300 83.500 545.600 ;
        RECT 84.400 544.200 85.200 555.800 ;
        RECT 86.000 547.600 86.800 548.400 ;
        RECT 87.600 544.200 88.400 555.800 ;
        RECT 89.200 544.200 90.000 557.800 ;
        RECT 90.800 544.200 91.600 557.800 ;
        RECT 95.600 549.600 96.400 550.400 ;
        RECT 95.700 546.400 96.300 549.600 ;
        RECT 95.600 546.300 96.400 546.400 ;
        RECT 94.100 545.700 96.400 546.300 ;
        RECT 100.400 546.200 101.200 551.800 ;
        RECT 102.000 547.600 102.800 548.400 ;
        RECT 81.300 541.700 83.500 542.300 ;
        RECT 58.800 531.700 61.100 532.300 ;
        RECT 58.800 531.600 59.600 531.700 ;
        RECT 58.800 529.600 59.600 530.400 ;
        RECT 65.200 523.600 66.000 524.400 ;
        RECT 74.800 524.200 75.600 537.800 ;
        RECT 76.400 524.200 77.200 537.800 ;
        RECT 78.000 524.200 78.800 537.800 ;
        RECT 79.600 526.200 80.400 537.800 ;
        RECT 81.300 536.400 81.900 541.700 ;
        RECT 81.200 535.600 82.000 536.400 ;
        RECT 31.600 521.600 32.400 522.400 ;
        RECT 41.200 521.600 42.000 522.400 ;
        RECT 57.200 521.600 58.000 522.400 ;
        RECT 17.200 507.600 18.000 508.400 ;
        RECT 20.400 506.200 21.200 511.800 ;
        RECT 22.000 507.600 22.800 508.400 ;
        RECT 18.800 503.600 19.600 504.400 ;
        RECT 23.600 504.200 24.400 515.800 ;
        RECT 26.800 509.600 27.600 510.400 ;
        RECT 25.200 505.600 26.000 506.400 ;
        RECT 18.900 502.400 19.500 503.600 ;
        RECT 18.800 501.600 19.600 502.400 ;
        RECT 15.600 499.600 16.400 500.400 ;
        RECT 15.700 492.400 16.300 499.600 ;
        RECT 17.200 493.600 18.000 494.400 ;
        RECT 17.300 492.400 17.900 493.600 ;
        RECT 14.000 491.600 14.800 492.400 ;
        RECT 15.600 491.600 16.400 492.400 ;
        RECT 17.200 491.600 18.000 492.400 ;
        RECT 14.100 490.400 14.700 491.600 ;
        RECT 14.000 489.600 14.800 490.400 ;
        RECT 15.700 484.400 16.300 491.600 ;
        RECT 17.200 490.300 18.000 490.400 ;
        RECT 18.900 490.300 19.500 501.600 ;
        RECT 22.000 493.600 22.800 494.400 ;
        RECT 20.400 491.600 21.200 492.400 ;
        RECT 20.500 490.400 21.100 491.600 ;
        RECT 17.200 489.700 19.500 490.300 ;
        RECT 17.200 489.600 18.000 489.700 ;
        RECT 20.400 489.600 21.200 490.400 ;
        RECT 20.400 485.600 21.200 486.400 ;
        RECT 15.600 483.600 16.400 484.400 ;
        RECT 12.400 469.600 13.200 470.400 ;
        RECT 9.200 447.600 10.000 448.400 ;
        RECT 12.500 440.400 13.100 469.600 ;
        RECT 14.000 464.200 14.800 475.800 ;
        RECT 18.800 473.600 19.600 474.400 ;
        RECT 20.500 468.400 21.100 485.600 ;
        RECT 22.100 480.400 22.700 493.600 ;
        RECT 23.600 490.200 24.400 495.800 ;
        RECT 25.300 494.400 25.900 505.600 ;
        RECT 25.200 493.600 26.000 494.400 ;
        RECT 26.800 486.200 27.600 497.800 ;
        RECT 30.000 491.600 30.800 492.400 ;
        RECT 30.000 489.600 30.800 490.400 ;
        RECT 22.000 479.600 22.800 480.400 ;
        RECT 26.800 473.600 27.600 474.400 ;
        RECT 26.900 472.400 27.500 473.600 ;
        RECT 26.800 471.600 27.600 472.400 ;
        RECT 30.100 470.400 30.700 489.600 ;
        RECT 31.700 480.400 32.300 521.600 ;
        RECT 33.200 504.200 34.000 515.800 ;
        RECT 44.400 512.300 45.200 512.400 ;
        RECT 46.000 512.300 46.800 512.400 ;
        RECT 44.400 511.700 46.800 512.300 ;
        RECT 44.400 511.600 45.200 511.700 ;
        RECT 46.000 511.600 46.800 511.700 ;
        RECT 54.000 511.600 54.800 512.400 ;
        RECT 55.600 511.600 56.400 512.400 ;
        RECT 66.800 511.600 67.600 512.400 ;
        RECT 71.600 511.600 72.400 512.400 ;
        RECT 54.100 510.400 54.700 511.600 ;
        RECT 41.200 509.600 42.000 510.400 ;
        RECT 42.800 509.600 43.600 510.400 ;
        RECT 46.000 509.600 46.800 510.400 ;
        RECT 47.600 509.600 48.400 510.400 ;
        RECT 52.400 509.600 53.200 510.400 ;
        RECT 54.000 509.600 54.800 510.400 ;
        RECT 38.000 507.600 38.800 508.400 ;
        RECT 39.600 507.600 40.400 508.400 ;
        RECT 38.100 504.400 38.700 507.600 ;
        RECT 38.000 503.600 38.800 504.400 ;
        RECT 34.800 495.600 35.600 496.400 ;
        RECT 31.600 479.600 32.400 480.400 ;
        RECT 22.000 469.600 22.800 470.400 ;
        RECT 23.600 469.600 24.400 470.400 ;
        RECT 30.000 469.600 30.800 470.400 ;
        RECT 20.400 467.600 21.200 468.400 ;
        RECT 14.000 451.600 14.800 452.600 ;
        RECT 15.600 446.200 16.400 457.800 ;
        RECT 17.200 455.600 18.000 456.400 ;
        RECT 17.300 454.400 17.900 455.600 ;
        RECT 17.200 453.600 18.000 454.400 ;
        RECT 12.400 439.600 13.200 440.400 ;
        RECT 9.200 431.600 10.000 432.400 ;
        RECT 2.800 429.600 3.600 430.400 ;
        RECT 6.000 429.600 6.800 430.400 ;
        RECT 6.100 376.400 6.700 429.600 ;
        RECT 7.600 427.600 8.400 428.400 ;
        RECT 7.700 414.400 8.300 427.600 ;
        RECT 9.300 424.400 9.900 431.600 ;
        RECT 10.800 427.600 11.600 428.400 ;
        RECT 9.200 423.600 10.000 424.400 ;
        RECT 7.600 413.600 8.400 414.400 ;
        RECT 9.200 404.200 10.000 417.800 ;
        RECT 10.800 404.200 11.600 417.800 ;
        RECT 12.400 406.200 13.200 417.800 ;
        RECT 14.000 413.600 14.800 414.400 ;
        RECT 15.600 406.200 16.400 417.800 ;
        RECT 17.300 416.400 17.900 453.600 ;
        RECT 18.800 450.200 19.600 455.800 ;
        RECT 20.500 454.400 21.100 467.600 ;
        RECT 22.100 464.400 22.700 469.600 ;
        RECT 22.000 463.600 22.800 464.400 ;
        RECT 20.400 453.600 21.200 454.400 ;
        RECT 22.000 453.600 22.800 454.400 ;
        RECT 26.800 453.600 27.600 454.400 ;
        RECT 22.100 452.400 22.700 453.600 ;
        RECT 22.000 451.600 22.800 452.400 ;
        RECT 23.600 451.600 24.400 452.400 ;
        RECT 28.400 451.600 29.200 452.400 ;
        RECT 25.200 449.600 26.000 450.400 ;
        RECT 28.400 449.600 29.200 450.400 ;
        RECT 26.800 447.600 27.600 448.400 ;
        RECT 22.000 439.600 22.800 440.400 ;
        RECT 22.100 438.400 22.700 439.600 ;
        RECT 22.000 437.600 22.800 438.400 ;
        RECT 25.200 431.600 26.000 432.400 ;
        RECT 17.200 415.600 18.000 416.400 ;
        RECT 9.200 384.200 10.000 397.800 ;
        RECT 10.800 384.200 11.600 397.800 ;
        RECT 12.400 384.200 13.200 395.800 ;
        RECT 14.000 387.600 14.800 388.400 ;
        RECT 14.100 382.300 14.700 387.600 ;
        RECT 15.600 384.200 16.400 395.800 ;
        RECT 17.300 386.400 17.900 415.600 ;
        RECT 18.800 406.200 19.600 417.800 ;
        RECT 20.400 404.200 21.200 417.800 ;
        RECT 22.000 404.200 22.800 417.800 ;
        RECT 23.600 404.200 24.400 417.800 ;
        RECT 25.200 411.600 26.000 412.400 ;
        RECT 17.200 385.600 18.000 386.400 ;
        RECT 18.800 384.200 19.600 395.800 ;
        RECT 20.400 384.200 21.200 397.800 ;
        RECT 22.000 384.200 22.800 397.800 ;
        RECT 23.600 384.200 24.400 397.800 ;
        RECT 25.300 390.400 25.900 411.600 ;
        RECT 25.200 389.600 26.000 390.400 ;
        RECT 12.500 381.700 14.700 382.300 ;
        RECT 12.500 378.400 13.100 381.700 ;
        RECT 12.400 377.600 13.200 378.400 ;
        RECT 6.000 375.600 6.800 376.400 ;
        RECT 9.200 375.600 10.000 376.400 ;
        RECT 12.400 375.600 13.200 376.400 ;
        RECT 6.000 373.600 6.800 374.400 ;
        RECT 7.600 373.600 8.400 374.400 ;
        RECT 7.700 372.400 8.300 373.600 ;
        RECT 9.300 372.400 9.900 375.600 ;
        RECT 4.400 371.600 5.200 372.400 ;
        RECT 7.600 371.600 8.400 372.400 ;
        RECT 9.200 371.600 10.000 372.400 ;
        RECT 9.300 360.400 9.900 371.600 ;
        RECT 12.500 370.400 13.100 375.600 ;
        RECT 14.000 373.600 14.800 374.400 ;
        RECT 15.600 371.600 16.400 372.400 ;
        RECT 12.400 369.600 13.200 370.400 ;
        RECT 20.400 369.600 21.200 370.400 ;
        RECT 15.600 363.600 16.400 364.400 ;
        RECT 6.000 359.600 6.800 360.400 ;
        RECT 9.200 359.600 10.000 360.400 ;
        RECT 6.100 350.400 6.700 359.600 ;
        RECT 9.200 357.600 10.000 358.400 ;
        RECT 9.300 352.400 9.900 357.600 ;
        RECT 9.200 351.600 10.000 352.400 ;
        RECT 6.000 349.600 6.800 350.400 ;
        RECT 12.400 349.600 13.200 350.400 ;
        RECT 9.200 343.600 10.000 344.400 ;
        RECT 9.300 342.400 9.900 343.600 ;
        RECT 9.200 341.600 10.000 342.400 ;
        RECT 12.500 340.400 13.100 349.600 ;
        RECT 15.700 348.400 16.300 363.600 ;
        RECT 20.500 362.400 21.100 369.600 ;
        RECT 20.400 361.600 21.200 362.400 ;
        RECT 25.300 358.300 25.900 389.600 ;
        RECT 26.900 382.400 27.500 447.600 ;
        RECT 28.500 438.400 29.100 449.600 ;
        RECT 28.400 437.600 29.200 438.400 ;
        RECT 28.400 430.300 29.200 430.400 ;
        RECT 30.100 430.300 30.700 469.600 ;
        RECT 31.700 468.400 32.300 479.600 ;
        RECT 31.600 467.600 32.400 468.400 ;
        RECT 33.200 466.200 34.000 471.800 ;
        RECT 33.200 453.600 34.000 454.400 ;
        RECT 33.300 452.400 33.900 453.600 ;
        RECT 34.900 452.400 35.500 495.600 ;
        RECT 36.400 486.200 37.200 497.800 ;
        RECT 38.000 487.600 38.800 488.400 ;
        RECT 36.400 464.200 37.200 475.800 ;
        RECT 38.100 468.400 38.700 487.600 ;
        RECT 39.700 486.400 40.300 507.600 ;
        RECT 41.300 506.400 41.900 509.600 ;
        RECT 41.200 505.600 42.000 506.400 ;
        RECT 46.100 500.400 46.700 509.600 ;
        RECT 47.700 508.400 48.300 509.600 ;
        RECT 47.600 507.600 48.400 508.400 ;
        RECT 49.200 505.600 50.000 506.400 ;
        RECT 46.000 499.600 46.800 500.400 ;
        RECT 41.200 497.600 42.000 498.400 ;
        RECT 41.300 490.400 41.900 497.600 ;
        RECT 42.800 493.600 43.600 494.400 ;
        RECT 44.400 493.600 45.200 494.400 ;
        RECT 49.200 493.600 50.000 494.400 ;
        RECT 41.200 489.600 42.000 490.400 ;
        RECT 42.900 486.400 43.500 493.600 ;
        RECT 44.500 492.400 45.100 493.600 ;
        RECT 44.400 491.600 45.200 492.400 ;
        RECT 46.000 491.600 46.800 492.400 ;
        RECT 47.600 491.600 48.400 492.400 ;
        RECT 49.200 491.600 50.000 492.400 ;
        RECT 47.700 490.400 48.300 491.600 ;
        RECT 47.600 489.600 48.400 490.400 ;
        RECT 49.300 488.300 49.900 491.600 ;
        RECT 52.500 488.400 53.100 509.600 ;
        RECT 55.700 508.400 56.300 511.600 ;
        RECT 60.400 509.600 61.200 510.400 ;
        RECT 55.600 507.600 56.400 508.400 ;
        RECT 55.600 497.600 56.400 498.400 ;
        RECT 55.700 492.400 56.300 497.600 ;
        RECT 55.600 491.600 56.400 492.400 ;
        RECT 57.200 491.600 58.000 492.400 ;
        RECT 58.800 491.600 59.600 492.400 ;
        RECT 60.500 492.300 61.100 509.600 ;
        RECT 62.000 507.600 62.800 508.400 ;
        RECT 62.100 494.300 62.700 507.600 ;
        RECT 66.900 500.400 67.500 511.600 ;
        RECT 71.600 509.600 72.400 510.400 ;
        RECT 66.800 499.600 67.600 500.400 ;
        RECT 65.200 495.600 66.000 496.400 ;
        RECT 63.600 494.300 64.400 494.400 ;
        RECT 62.100 493.700 64.400 494.300 ;
        RECT 63.600 493.600 64.400 493.700 ;
        RECT 65.300 492.400 65.900 495.600 ;
        RECT 66.900 492.400 67.500 499.600 ;
        RECT 71.700 494.400 72.300 509.600 ;
        RECT 73.200 507.600 74.000 508.400 ;
        RECT 73.300 504.400 73.900 507.600 ;
        RECT 74.800 506.200 75.600 511.800 ;
        RECT 73.200 503.600 74.000 504.400 ;
        RECT 78.000 504.200 78.800 515.800 ;
        RECT 81.300 514.400 81.900 535.600 ;
        RECT 82.800 526.200 83.600 537.800 ;
        RECT 84.400 533.600 85.200 534.400 ;
        RECT 86.000 526.200 86.800 537.800 ;
        RECT 87.600 524.200 88.400 537.800 ;
        RECT 89.200 524.200 90.000 537.800 ;
        RECT 94.100 532.400 94.700 545.700 ;
        RECT 95.600 545.600 96.400 545.700 ;
        RECT 98.800 533.600 99.600 534.400 ;
        RECT 94.000 531.600 94.800 532.400 ;
        RECT 98.900 530.400 99.500 533.600 ;
        RECT 100.400 531.600 101.200 532.400 ;
        RECT 98.800 529.600 99.600 530.400 ;
        RECT 89.200 521.600 90.000 522.400 ;
        RECT 81.200 513.600 82.000 514.400 ;
        RECT 86.000 513.600 86.800 514.400 ;
        RECT 79.600 511.600 80.400 512.400 ;
        RECT 79.700 510.200 80.300 511.600 ;
        RECT 86.100 510.400 86.700 513.600 ;
        RECT 79.600 509.400 80.400 510.200 ;
        RECT 86.000 509.600 86.800 510.400 ;
        RECT 79.600 507.600 80.400 508.400 ;
        RECT 71.600 493.600 72.400 494.400 ;
        RECT 62.000 492.300 62.800 492.400 ;
        RECT 60.500 491.700 62.800 492.300 ;
        RECT 62.000 491.600 62.800 491.700 ;
        RECT 65.200 491.600 66.000 492.400 ;
        RECT 66.800 491.600 67.600 492.400 ;
        RECT 71.600 491.600 72.400 492.400 ;
        RECT 55.700 490.400 56.300 491.600 ;
        RECT 55.600 489.600 56.400 490.400 ;
        RECT 47.700 487.700 49.900 488.300 ;
        RECT 39.600 485.600 40.400 486.400 ;
        RECT 42.800 485.600 43.600 486.400 ;
        RECT 47.700 484.400 48.300 487.700 ;
        RECT 52.400 487.600 53.200 488.400 ;
        RECT 47.600 483.600 48.400 484.400 ;
        RECT 39.600 471.600 40.400 472.400 ;
        RECT 39.700 470.400 40.300 471.600 ;
        RECT 39.600 469.600 40.400 470.400 ;
        RECT 38.000 467.600 38.800 468.400 ;
        RECT 41.200 467.600 42.000 468.400 ;
        RECT 38.000 459.600 38.800 460.400 ;
        RECT 38.100 458.400 38.700 459.600 ;
        RECT 41.300 458.400 41.900 467.600 ;
        RECT 46.000 464.200 46.800 475.800 ;
        RECT 38.000 457.600 38.800 458.400 ;
        RECT 41.200 457.600 42.000 458.400 ;
        RECT 46.000 457.600 46.800 458.400 ;
        RECT 36.400 455.600 37.200 456.400 ;
        RECT 36.500 454.400 37.100 455.600 ;
        RECT 36.400 453.600 37.200 454.400 ;
        RECT 33.200 451.600 34.000 452.400 ;
        RECT 34.800 451.600 35.600 452.400 ;
        RECT 44.400 451.600 45.200 452.400 ;
        RECT 33.300 432.400 33.900 451.600 ;
        RECT 44.500 444.400 45.100 451.600 ;
        RECT 46.100 450.400 46.700 457.600 ;
        RECT 47.700 454.400 48.300 483.600 ;
        RECT 57.300 482.400 57.900 491.600 ;
        RECT 58.800 489.600 59.600 490.400 ;
        RECT 65.200 487.600 66.000 488.400 ;
        RECT 57.200 481.600 58.000 482.400 ;
        RECT 50.800 475.600 51.600 476.400 ;
        RECT 57.200 475.600 58.000 476.400 ;
        RECT 57.300 472.400 57.900 475.600 ;
        RECT 57.200 471.600 58.000 472.400 ;
        RECT 58.800 471.600 59.600 472.400 ;
        RECT 54.000 469.600 54.800 470.400 ;
        RECT 57.300 468.400 57.900 471.600 ;
        RECT 58.900 468.400 59.500 471.600 ;
        RECT 65.300 470.400 65.900 487.600 ;
        RECT 71.700 484.400 72.300 491.600 ;
        RECT 73.300 486.400 73.900 503.600 ;
        RECT 74.800 501.600 75.600 502.400 ;
        RECT 74.900 494.400 75.500 501.600 ;
        RECT 79.700 494.400 80.300 507.600 ;
        RECT 87.600 504.200 88.400 515.800 ;
        RECT 84.400 499.600 85.200 500.400 ;
        RECT 84.500 496.400 85.100 499.600 ;
        RECT 84.400 495.600 85.200 496.400 ;
        RECT 74.800 493.600 75.600 494.400 ;
        RECT 79.600 493.600 80.400 494.400 ;
        RECT 87.600 493.600 88.400 494.400 ;
        RECT 79.600 492.300 80.400 492.400 ;
        RECT 79.600 491.700 85.100 492.300 ;
        RECT 79.600 491.600 80.400 491.700 ;
        RECT 84.500 490.400 85.100 491.700 ;
        RECT 74.800 489.600 75.600 490.400 ;
        RECT 78.000 489.600 78.800 490.400 ;
        RECT 82.800 489.600 83.600 490.400 ;
        RECT 84.400 489.600 85.200 490.400 ;
        RECT 87.700 490.300 88.300 493.600 ;
        RECT 89.300 492.400 89.900 521.600 ;
        RECT 94.000 506.200 94.800 511.800 ;
        RECT 90.800 503.600 91.600 504.400 ;
        RECT 92.400 503.600 93.200 504.400 ;
        RECT 94.000 503.600 94.800 504.400 ;
        RECT 97.200 504.200 98.000 515.800 ;
        RECT 89.200 491.600 90.000 492.400 ;
        RECT 87.700 489.700 89.900 490.300 ;
        RECT 73.200 485.600 74.000 486.400 ;
        RECT 71.600 483.600 72.400 484.400 ;
        RECT 71.700 480.400 72.300 483.600 ;
        RECT 73.200 481.600 74.000 482.400 ;
        RECT 71.600 479.600 72.400 480.400 ;
        RECT 71.600 473.600 72.400 474.400 ;
        RECT 71.700 470.400 72.300 473.600 ;
        RECT 73.300 470.400 73.900 481.600 ;
        RECT 74.900 474.400 75.500 489.600 ;
        RECT 81.200 487.600 82.000 488.400 ;
        RECT 82.900 478.400 83.500 489.600 ;
        RECT 86.000 483.600 86.800 484.400 ;
        RECT 87.600 483.600 88.400 484.400 ;
        RECT 86.100 482.400 86.700 483.600 ;
        RECT 86.000 481.600 86.800 482.400 ;
        RECT 86.000 479.600 86.800 480.400 ;
        RECT 82.800 477.600 83.600 478.400 ;
        RECT 74.800 473.600 75.600 474.400 ;
        RECT 86.100 470.400 86.700 479.600 ;
        RECT 87.700 470.400 88.300 483.600 ;
        RECT 62.000 469.600 62.800 470.400 ;
        RECT 65.200 469.600 66.000 470.400 ;
        RECT 71.600 469.600 72.400 470.400 ;
        RECT 73.200 469.600 74.000 470.400 ;
        RECT 81.200 469.600 82.000 470.400 ;
        RECT 86.000 469.600 86.800 470.400 ;
        RECT 87.600 469.600 88.400 470.400 ;
        RECT 52.400 467.600 53.200 468.400 ;
        RECT 57.200 467.600 58.000 468.400 ;
        RECT 58.800 467.600 59.600 468.400 ;
        RECT 62.100 466.400 62.700 469.600 ;
        RECT 63.600 467.600 64.400 468.400 ;
        RECT 62.000 465.600 62.800 466.400 ;
        RECT 63.700 462.400 64.300 467.600 ;
        RECT 63.600 461.600 64.400 462.400 ;
        RECT 65.300 460.300 65.900 469.600 ;
        RECT 68.400 463.600 69.200 464.400 ;
        RECT 63.700 459.700 65.900 460.300 ;
        RECT 47.600 453.600 48.400 454.400 ;
        RECT 50.800 453.600 51.600 454.400 ;
        RECT 49.200 451.600 50.000 452.400 ;
        RECT 46.000 449.600 46.800 450.400 ;
        RECT 49.300 448.400 49.900 451.600 ;
        RECT 52.400 450.200 53.200 455.800 ;
        RECT 54.000 455.600 54.800 456.400 ;
        RECT 54.100 454.400 54.700 455.600 ;
        RECT 54.000 453.600 54.800 454.400 ;
        RECT 46.000 447.600 46.800 448.400 ;
        RECT 49.200 447.600 50.000 448.400 ;
        RECT 44.400 443.600 45.200 444.400 ;
        RECT 33.200 431.600 34.000 432.400 ;
        RECT 44.500 430.400 45.100 443.600 ;
        RECT 28.400 429.700 30.700 430.300 ;
        RECT 28.400 429.600 29.200 429.700 ;
        RECT 36.400 429.600 37.200 430.400 ;
        RECT 44.400 429.600 45.200 430.400 ;
        RECT 28.500 416.400 29.100 429.600 ;
        RECT 33.200 427.600 34.000 428.400 ;
        RECT 38.000 427.600 38.800 428.400 ;
        RECT 39.600 427.600 40.400 428.400 ;
        RECT 38.100 426.400 38.700 427.600 ;
        RECT 31.600 425.600 32.400 426.400 ;
        RECT 38.000 425.600 38.800 426.400 ;
        RECT 31.700 422.400 32.300 425.600 ;
        RECT 36.400 423.600 37.200 424.400 ;
        RECT 31.600 421.600 32.400 422.400 ;
        RECT 36.500 418.400 37.100 423.600 ;
        RECT 36.400 417.600 37.200 418.400 ;
        RECT 28.400 415.600 29.200 416.400 ;
        RECT 39.700 412.400 40.300 427.600 ;
        RECT 42.800 421.600 43.600 422.400 ;
        RECT 42.900 414.400 43.500 421.600 ;
        RECT 44.400 415.600 45.200 416.400 ;
        RECT 42.800 413.600 43.600 414.400 ;
        RECT 39.600 411.600 40.400 412.400 ;
        RECT 36.400 409.600 37.200 410.400 ;
        RECT 36.500 394.400 37.100 409.600 ;
        RECT 36.400 393.600 37.200 394.400 ;
        RECT 39.700 390.400 40.300 411.600 ;
        RECT 42.900 398.400 43.500 413.600 ;
        RECT 44.500 412.400 45.100 415.600 ;
        RECT 44.400 411.600 45.200 412.400 ;
        RECT 46.100 398.400 46.700 447.600 ;
        RECT 49.200 435.600 50.000 436.400 ;
        RECT 49.300 412.400 49.900 435.600 ;
        RECT 50.800 427.600 51.600 428.400 ;
        RECT 52.400 426.200 53.200 431.800 ;
        RECT 54.100 428.400 54.700 453.600 ;
        RECT 55.600 446.200 56.400 457.800 ;
        RECT 58.800 451.600 59.600 452.400 ;
        RECT 58.900 450.400 59.500 451.600 ;
        RECT 58.800 449.600 59.600 450.400 ;
        RECT 54.000 427.600 54.800 428.400 ;
        RECT 52.400 423.600 53.200 424.400 ;
        RECT 55.600 424.200 56.400 435.800 ;
        RECT 60.400 429.600 61.200 430.400 ;
        RECT 63.700 428.400 64.300 459.700 ;
        RECT 65.200 446.200 66.000 457.800 ;
        RECT 73.300 454.300 73.900 469.600 ;
        RECT 81.300 468.400 81.900 469.600 ;
        RECT 78.000 467.600 78.800 468.400 ;
        RECT 79.600 467.600 80.400 468.400 ;
        RECT 81.200 467.600 82.000 468.400 ;
        RECT 74.800 463.600 75.600 464.400 ;
        RECT 71.700 453.700 73.900 454.300 ;
        RECT 71.700 452.400 72.300 453.700 ;
        RECT 71.600 451.600 72.400 452.400 ;
        RECT 73.200 451.600 74.000 452.400 ;
        RECT 73.300 448.400 73.900 451.600 ;
        RECT 70.000 447.600 70.800 448.400 ;
        RECT 73.200 447.600 74.000 448.400 ;
        RECT 63.600 427.600 64.400 428.400 ;
        RECT 57.200 425.600 58.000 426.400 ;
        RECT 47.600 411.600 48.400 412.400 ;
        RECT 49.200 411.600 50.000 412.400 ;
        RECT 50.800 411.600 51.600 412.400 ;
        RECT 50.900 410.400 51.500 411.600 ;
        RECT 47.600 409.600 48.400 410.400 ;
        RECT 50.800 409.600 51.600 410.400 ;
        RECT 42.800 397.600 43.600 398.400 ;
        RECT 46.000 397.600 46.800 398.400 ;
        RECT 36.400 389.600 37.200 390.400 ;
        RECT 39.600 389.600 40.400 390.400 ;
        RECT 46.000 389.600 46.800 390.400 ;
        RECT 34.800 385.600 35.600 386.400 ;
        RECT 26.800 381.600 27.600 382.400 ;
        RECT 33.200 375.600 34.000 376.400 ;
        RECT 26.800 373.600 27.600 374.400 ;
        RECT 28.400 371.600 29.200 372.400 ;
        RECT 34.900 370.400 35.500 385.600 ;
        RECT 36.500 372.400 37.100 389.600 ;
        RECT 39.600 387.600 40.400 388.400 ;
        RECT 47.600 386.200 48.400 391.800 ;
        RECT 38.000 383.600 38.800 384.400 ;
        RECT 42.800 383.600 43.600 384.400 ;
        RECT 47.600 383.600 48.400 384.400 ;
        RECT 50.800 384.200 51.600 395.800 ;
        RECT 38.100 376.300 38.700 383.600 ;
        RECT 39.600 381.600 40.400 382.400 ;
        RECT 39.700 378.400 40.300 381.600 ;
        RECT 39.600 377.600 40.400 378.400 ;
        RECT 38.100 375.700 40.300 376.300 ;
        RECT 38.000 373.600 38.800 374.400 ;
        RECT 36.400 371.600 37.200 372.400 ;
        RECT 39.700 370.400 40.300 375.700 ;
        RECT 42.900 374.400 43.500 383.600 ;
        RECT 42.800 373.600 43.600 374.400 ;
        RECT 44.400 373.600 45.200 374.400 ;
        RECT 42.800 371.600 43.600 372.400 ;
        RECT 31.600 369.600 32.400 370.400 ;
        RECT 33.200 369.600 34.000 370.400 ;
        RECT 34.800 369.600 35.600 370.400 ;
        RECT 39.600 369.600 40.400 370.400 ;
        RECT 46.000 369.600 46.800 370.400 ;
        RECT 31.700 368.400 32.300 369.600 ;
        RECT 31.600 367.600 32.400 368.400 ;
        RECT 34.800 367.600 35.600 368.400 ;
        RECT 28.400 363.600 29.200 364.400 ;
        RECT 28.500 358.400 29.100 363.600 ;
        RECT 15.600 347.600 16.400 348.400 ;
        RECT 17.200 345.600 18.000 346.400 ;
        RECT 14.000 341.600 14.800 342.400 ;
        RECT 7.600 339.600 8.400 340.400 ;
        RECT 12.400 339.600 13.200 340.400 ;
        RECT 7.700 332.400 8.300 339.600 ;
        RECT 7.600 331.600 8.400 332.400 ;
        RECT 9.200 324.200 10.000 337.800 ;
        RECT 10.800 324.200 11.600 337.800 ;
        RECT 12.400 326.200 13.200 337.800 ;
        RECT 14.100 334.400 14.700 341.600 ;
        RECT 14.000 333.600 14.800 334.400 ;
        RECT 15.600 326.200 16.400 337.800 ;
        RECT 17.300 336.400 17.900 345.600 ;
        RECT 18.800 344.200 19.600 357.800 ;
        RECT 20.400 344.200 21.200 357.800 ;
        RECT 23.700 357.700 25.900 358.300 ;
        RECT 22.000 344.200 22.800 355.800 ;
        RECT 23.700 350.400 24.300 357.700 ;
        RECT 28.400 357.600 29.200 358.400 ;
        RECT 23.600 349.600 24.400 350.400 ;
        RECT 23.600 347.600 24.400 348.400 ;
        RECT 25.200 344.200 26.000 355.800 ;
        RECT 26.800 345.600 27.600 346.400 ;
        RECT 28.400 344.200 29.200 355.800 ;
        RECT 30.000 344.200 30.800 357.800 ;
        RECT 31.600 344.200 32.400 357.800 ;
        RECT 33.200 344.200 34.000 357.800 ;
        RECT 34.900 348.400 35.500 367.600 ;
        RECT 42.800 361.600 43.600 362.400 ;
        RECT 42.900 354.400 43.500 361.600 ;
        RECT 47.700 358.400 48.300 383.600 ;
        RECT 52.500 374.400 53.100 423.600 ;
        RECT 55.600 413.600 56.400 414.400 ;
        RECT 55.600 411.600 56.400 412.400 ;
        RECT 55.700 402.400 56.300 411.600 ;
        RECT 55.600 401.600 56.400 402.400 ;
        RECT 54.000 391.600 54.800 392.400 ;
        RECT 54.100 390.400 54.700 391.600 ;
        RECT 57.300 390.400 57.900 425.600 ;
        RECT 63.700 424.400 64.300 427.600 ;
        RECT 63.600 423.600 64.400 424.400 ;
        RECT 65.200 424.200 66.000 435.800 ;
        RECT 71.600 435.600 72.400 436.400 ;
        RECT 66.800 433.600 67.600 434.400 ;
        RECT 70.000 433.600 70.800 434.400 ;
        RECT 62.000 413.600 62.800 414.400 ;
        RECT 63.600 413.600 64.400 414.400 ;
        RECT 62.100 412.400 62.700 413.600 ;
        RECT 58.800 411.600 59.600 412.400 ;
        RECT 60.400 411.600 61.200 412.400 ;
        RECT 62.000 411.600 62.800 412.400 ;
        RECT 58.900 410.400 59.500 411.600 ;
        RECT 58.800 409.600 59.600 410.400 ;
        RECT 65.200 410.200 66.000 415.800 ;
        RECT 66.900 414.400 67.500 433.600 ;
        RECT 71.700 430.400 72.300 435.600 ;
        RECT 73.200 433.600 74.000 434.400 ;
        RECT 73.300 432.400 73.900 433.600 ;
        RECT 73.200 431.600 74.000 432.400 ;
        RECT 73.300 430.400 73.900 431.600 ;
        RECT 71.600 429.600 72.400 430.400 ;
        RECT 73.200 429.600 74.000 430.400 ;
        RECT 66.800 413.600 67.600 414.400 ;
        RECT 68.400 406.200 69.200 417.800 ;
        RECT 71.600 415.600 72.400 416.400 ;
        RECT 70.000 411.600 70.800 412.600 ;
        RECT 71.700 412.400 72.300 415.600 ;
        RECT 71.600 411.600 72.400 412.400 ;
        RECT 65.200 403.600 66.000 404.400 ;
        RECT 74.900 404.300 75.500 463.600 ;
        RECT 78.100 454.400 78.700 467.600 ;
        RECT 79.700 466.400 80.300 467.600 ;
        RECT 79.600 465.600 80.400 466.400 ;
        RECT 81.200 461.600 82.000 462.400 ;
        RECT 81.300 454.400 81.900 461.600 ;
        RECT 86.100 454.400 86.700 469.600 ;
        RECT 78.000 453.600 78.800 454.400 ;
        RECT 79.600 453.600 80.400 454.400 ;
        RECT 81.200 453.600 82.000 454.400 ;
        RECT 82.800 453.600 83.600 454.400 ;
        RECT 86.000 453.600 86.800 454.400 ;
        RECT 79.600 451.600 80.400 452.400 ;
        RECT 78.000 445.600 78.800 446.400 ;
        RECT 78.100 430.400 78.700 445.600 ;
        RECT 78.000 430.300 78.800 430.400 ;
        RECT 73.300 403.700 75.500 404.300 ;
        RECT 76.500 429.700 78.800 430.300 ;
        RECT 65.300 398.400 65.900 403.600 ;
        RECT 65.200 397.600 66.000 398.400 ;
        RECT 66.800 397.600 67.600 398.400 ;
        RECT 54.000 389.600 54.800 390.400 ;
        RECT 57.200 389.600 58.000 390.400 ;
        RECT 55.600 387.600 56.400 388.400 ;
        RECT 55.700 374.400 56.300 387.600 ;
        RECT 60.400 384.200 61.200 395.800 ;
        RECT 66.900 390.400 67.500 397.600 ;
        RECT 73.300 392.400 73.900 403.700 ;
        RECT 74.800 401.600 75.600 402.400 ;
        RECT 73.200 391.600 74.000 392.400 ;
        RECT 74.900 390.400 75.500 401.600 ;
        RECT 66.800 389.600 67.600 390.400 ;
        RECT 74.800 389.600 75.600 390.400 ;
        RECT 70.000 383.600 70.800 384.400 ;
        RECT 70.100 376.400 70.700 383.600 ;
        RECT 70.000 375.600 70.800 376.400 ;
        RECT 49.200 373.600 50.000 374.400 ;
        RECT 52.400 373.600 53.200 374.400 ;
        RECT 55.600 373.600 56.400 374.400 ;
        RECT 57.200 373.600 58.000 374.400 ;
        RECT 66.800 373.600 67.600 374.400 ;
        RECT 57.300 372.400 57.900 373.600 ;
        RECT 49.200 371.600 50.000 372.400 ;
        RECT 55.600 371.600 56.400 372.400 ;
        RECT 57.200 371.600 58.000 372.400 ;
        RECT 58.800 371.600 59.600 372.400 ;
        RECT 63.600 371.600 64.400 372.400 ;
        RECT 49.300 358.400 49.900 371.600 ;
        RECT 55.700 370.300 56.300 371.600 ;
        RECT 58.900 370.400 59.500 371.600 ;
        RECT 55.700 369.700 57.900 370.300 ;
        RECT 57.300 358.400 57.900 369.700 ;
        RECT 58.800 369.600 59.600 370.400 ;
        RECT 63.700 364.400 64.300 371.600 ;
        RECT 66.900 366.400 67.500 373.600 ;
        RECT 73.200 369.600 74.000 370.400 ;
        RECT 66.800 365.600 67.600 366.400 ;
        RECT 76.500 364.400 77.100 429.700 ;
        RECT 78.000 429.600 78.800 429.700 ;
        RECT 78.000 406.200 78.800 417.800 ;
        RECT 79.700 402.400 80.300 451.600 ;
        RECT 81.300 434.400 81.900 453.600 ;
        RECT 82.900 452.400 83.500 453.600 ;
        RECT 82.800 451.600 83.600 452.400 ;
        RECT 87.700 452.300 88.300 469.600 ;
        RECT 89.300 458.400 89.900 489.700 ;
        RECT 90.900 478.400 91.500 503.600 ;
        RECT 92.500 500.400 93.100 503.600 ;
        RECT 92.400 499.600 93.200 500.400 ;
        RECT 94.100 498.400 94.700 503.600 ;
        RECT 94.000 497.600 94.800 498.400 ;
        RECT 98.900 494.400 99.500 529.600 ;
        RECT 100.500 528.400 101.100 531.600 ;
        RECT 100.400 527.600 101.200 528.400 ;
        RECT 102.100 514.400 102.700 547.600 ;
        RECT 103.600 544.200 104.400 555.800 ;
        RECT 105.200 549.400 106.000 550.200 ;
        RECT 105.300 542.300 105.900 549.400 ;
        RECT 111.600 547.600 112.400 548.400 ;
        RECT 110.000 543.600 110.800 544.400 ;
        RECT 113.200 544.200 114.000 555.800 ;
        RECT 119.600 546.200 120.400 551.800 ;
        RECT 121.200 547.600 122.000 548.400 ;
        RECT 118.000 543.600 118.800 544.400 ;
        RECT 122.800 544.200 123.600 555.800 ;
        RECT 124.400 549.400 125.200 550.400 ;
        RECT 132.400 544.200 133.200 555.800 ;
        RECT 145.200 549.600 146.000 550.400 ;
        RECT 145.300 546.400 145.900 549.600 ;
        RECT 145.200 545.600 146.000 546.400 ;
        RECT 137.200 543.600 138.000 544.400 ;
        RECT 151.600 544.200 152.400 557.800 ;
        RECT 153.200 544.200 154.000 557.800 ;
        RECT 154.800 544.200 155.600 555.800 ;
        RECT 156.400 553.600 157.200 554.400 ;
        RECT 156.500 548.400 157.100 553.600 ;
        RECT 156.400 547.600 157.200 548.400 ;
        RECT 158.000 544.200 158.800 555.800 ;
        RECT 159.600 545.600 160.400 546.400 ;
        RECT 103.700 541.700 105.900 542.300 ;
        RECT 103.700 538.400 104.300 541.700 ;
        RECT 103.600 537.600 104.400 538.400 ;
        RECT 103.600 535.600 104.400 536.400 ;
        RECT 108.400 535.600 109.200 536.400 ;
        RECT 103.700 530.400 104.300 535.600 ;
        RECT 108.500 534.400 109.100 535.600 ;
        RECT 105.200 533.600 106.000 534.400 ;
        RECT 108.400 533.600 109.200 534.400 ;
        RECT 105.200 531.600 106.000 532.400 ;
        RECT 103.600 529.600 104.400 530.400 ;
        RECT 105.300 522.400 105.900 531.600 ;
        RECT 110.100 530.400 110.700 543.600 ;
        RECT 118.000 541.600 118.800 542.400 ;
        RECT 116.400 539.600 117.200 540.400 ;
        RECT 111.600 533.600 112.400 534.400 ;
        RECT 113.200 531.600 114.000 532.400 ;
        RECT 116.500 530.400 117.100 539.600 ;
        RECT 118.100 538.400 118.700 541.600 ;
        RECT 137.300 540.400 137.900 543.600 ;
        RECT 159.700 542.300 160.300 545.600 ;
        RECT 161.200 544.200 162.000 555.800 ;
        RECT 162.800 544.200 163.600 557.800 ;
        RECT 164.400 544.200 165.200 557.800 ;
        RECT 166.000 544.200 166.800 557.800 ;
        RECT 190.000 553.600 190.800 554.400 ;
        RECT 186.800 551.600 187.600 552.400 ;
        RECT 193.200 551.600 194.000 552.400 ;
        RECT 196.400 551.600 197.200 552.400 ;
        RECT 167.600 549.600 168.400 550.400 ;
        RECT 177.200 549.600 178.000 550.400 ;
        RECT 183.600 549.600 184.400 550.400 ;
        RECT 186.800 549.600 187.600 550.400 ;
        RECT 190.000 549.600 190.800 550.400 ;
        RECT 175.600 547.600 176.600 548.400 ;
        RECT 158.100 541.700 160.300 542.300 ;
        RECT 137.200 539.600 138.000 540.400 ;
        RECT 118.000 537.600 118.800 538.400 ;
        RECT 125.800 535.000 126.600 535.800 ;
        RECT 127.600 535.000 131.800 535.600 ;
        RECT 132.400 535.000 133.200 535.800 ;
        RECT 124.400 533.600 125.200 534.400 ;
        RECT 122.800 531.600 123.600 532.400 ;
        RECT 110.000 529.600 110.800 530.400 ;
        RECT 116.400 529.600 117.200 530.400 ;
        RECT 105.200 521.600 106.000 522.400 ;
        RECT 102.000 513.600 102.800 514.400 ;
        RECT 105.200 513.600 106.000 514.400 ;
        RECT 105.300 510.400 105.900 513.600 ;
        RECT 100.400 509.600 101.200 510.400 ;
        RECT 105.200 509.600 106.000 510.400 ;
        RECT 100.500 504.400 101.100 509.600 ;
        RECT 100.400 503.600 101.200 504.400 ;
        RECT 106.800 504.200 107.600 515.800 ;
        RECT 110.100 512.400 110.700 529.600 ;
        RECT 110.000 511.600 110.800 512.400 ;
        RECT 114.800 511.600 115.600 512.400 ;
        RECT 114.900 506.400 115.500 511.600 ;
        RECT 116.500 508.400 117.100 529.600 ;
        RECT 122.900 518.400 123.500 531.600 ;
        RECT 124.500 530.400 125.100 533.600 ;
        RECT 124.400 529.600 125.200 530.400 ;
        RECT 125.800 530.200 126.400 535.000 ;
        RECT 127.600 534.800 128.400 535.000 ;
        RECT 131.000 534.800 131.800 535.000 ;
        RECT 132.600 534.200 133.200 535.000 ;
        RECT 128.400 533.600 133.200 534.200 ;
        RECT 146.800 533.600 147.600 534.400 ;
        RECT 128.400 533.400 129.200 533.600 ;
        RECT 132.600 530.200 133.200 533.600 ;
        RECT 140.400 531.600 141.200 532.400 ;
        RECT 125.800 529.400 126.600 530.200 ;
        RECT 132.400 529.400 133.200 530.200 ;
        RECT 132.400 527.600 133.200 528.400 ;
        RECT 132.500 518.400 133.100 527.600 ;
        RECT 142.000 523.600 142.800 524.400 ;
        RECT 122.800 517.600 123.600 518.400 ;
        RECT 132.400 517.600 133.200 518.400 ;
        RECT 130.800 511.600 131.600 512.400 ;
        RECT 130.900 510.400 131.500 511.600 ;
        RECT 142.100 510.400 142.700 523.600 ;
        RECT 121.200 509.600 122.000 510.400 ;
        RECT 126.000 509.600 126.800 510.400 ;
        RECT 127.600 509.600 128.400 510.400 ;
        RECT 130.800 509.600 131.600 510.400 ;
        RECT 137.200 509.600 138.000 510.400 ;
        RECT 142.000 509.600 142.800 510.400 ;
        RECT 126.100 508.400 126.700 509.600 ;
        RECT 116.400 507.600 117.200 508.400 ;
        RECT 126.000 507.600 126.800 508.400 ;
        RECT 116.500 506.400 117.100 507.600 ;
        RECT 114.800 505.600 115.600 506.400 ;
        RECT 116.400 505.600 117.200 506.400 ;
        RECT 119.600 505.600 120.400 506.400 ;
        RECT 111.600 503.600 112.400 504.400 ;
        RECT 113.200 503.600 114.000 504.400 ;
        RECT 118.000 503.600 118.800 504.400 ;
        RECT 105.200 499.600 106.000 500.400 ;
        RECT 105.300 494.400 105.900 499.600 ;
        RECT 106.800 497.600 107.600 498.400 ;
        RECT 98.800 493.600 99.600 494.400 ;
        RECT 102.000 493.600 102.800 494.400 ;
        RECT 105.200 493.600 106.000 494.400 ;
        RECT 98.800 491.600 99.600 492.400 ;
        RECT 92.400 489.600 93.200 490.400 ;
        RECT 92.500 482.400 93.100 489.600 ;
        RECT 92.400 481.600 93.200 482.400 ;
        RECT 98.900 478.400 99.500 491.600 ;
        RECT 100.400 489.600 101.200 490.400 ;
        RECT 102.100 482.400 102.700 493.600 ;
        RECT 103.600 491.600 104.400 492.400 ;
        RECT 106.900 490.400 107.500 497.600 ;
        RECT 111.700 494.400 112.300 503.600 ;
        RECT 113.300 500.400 113.900 503.600 ;
        RECT 113.200 499.600 114.000 500.400 ;
        RECT 118.100 494.400 118.700 503.600 ;
        RECT 119.700 494.400 120.300 505.600 ;
        RECT 124.400 503.600 125.200 504.400 ;
        RECT 111.600 493.600 112.400 494.400 ;
        RECT 118.000 493.600 118.800 494.400 ;
        RECT 119.600 493.600 120.400 494.400 ;
        RECT 124.500 492.400 125.100 503.600 ;
        RECT 127.700 496.400 128.300 509.600 ;
        RECT 130.800 505.600 131.600 506.400 ;
        RECT 129.200 499.600 130.000 500.400 ;
        RECT 127.600 495.600 128.400 496.400 ;
        RECT 127.700 494.400 128.300 495.600 ;
        RECT 127.600 493.600 128.400 494.400 ;
        RECT 108.400 491.600 109.200 492.400 ;
        RECT 116.400 491.600 117.200 492.400 ;
        RECT 124.400 491.600 125.200 492.400 ;
        RECT 106.800 489.600 107.600 490.400 ;
        RECT 103.600 485.600 104.400 486.400 ;
        RECT 102.000 481.600 102.800 482.400 ;
        RECT 90.800 477.600 91.600 478.400 ;
        RECT 97.200 477.600 98.000 478.400 ;
        RECT 98.800 477.600 99.600 478.400 ;
        RECT 94.000 469.600 94.800 470.400 ;
        RECT 95.600 469.600 96.400 470.400 ;
        RECT 94.100 468.400 94.700 469.600 ;
        RECT 94.000 467.600 94.800 468.400 ;
        RECT 95.700 466.300 96.300 469.600 ;
        RECT 94.100 465.700 96.300 466.300 ;
        RECT 89.200 457.600 90.000 458.400 ;
        RECT 87.700 451.700 89.900 452.300 ;
        RECT 82.800 449.600 83.600 450.400 ;
        RECT 87.600 449.600 88.400 450.400 ;
        RECT 87.700 448.400 88.300 449.600 ;
        RECT 87.600 447.600 88.400 448.400 ;
        RECT 81.200 433.600 82.000 434.400 ;
        RECT 81.300 428.400 81.900 433.600 ;
        RECT 87.600 431.600 88.400 432.400 ;
        RECT 89.300 430.400 89.900 451.700 ;
        RECT 90.800 451.600 91.600 452.400 ;
        RECT 90.900 430.400 91.500 451.600 ;
        RECT 94.100 446.400 94.700 465.700 ;
        RECT 95.600 457.600 96.400 458.400 ;
        RECT 94.000 445.600 94.800 446.400 ;
        RECT 97.300 432.400 97.900 477.600 ;
        RECT 102.100 470.400 102.700 481.600 ;
        RECT 102.000 469.600 102.800 470.400 ;
        RECT 103.600 469.600 104.400 470.400 ;
        RECT 100.400 459.600 101.200 460.400 ;
        RECT 100.500 454.400 101.100 459.600 ;
        RECT 100.400 453.600 101.200 454.400 ;
        RECT 98.800 451.600 99.600 452.400 ;
        RECT 100.400 451.600 101.200 452.400 ;
        RECT 98.900 444.400 99.500 451.600 ;
        RECT 98.800 443.600 99.600 444.400 ;
        RECT 94.000 431.600 94.800 432.400 ;
        RECT 97.200 431.600 98.000 432.400 ;
        RECT 100.500 432.300 101.100 451.600 ;
        RECT 102.100 450.400 102.700 469.600 ;
        RECT 103.700 468.400 104.300 469.600 ;
        RECT 103.600 467.600 104.400 468.400 ;
        RECT 106.800 463.600 107.600 464.400 ;
        RECT 106.900 462.400 107.500 463.600 ;
        RECT 106.800 461.600 107.600 462.400 ;
        RECT 105.200 455.600 106.000 456.400 ;
        RECT 108.500 452.400 109.100 491.600 ;
        RECT 113.200 489.600 114.000 490.400 ;
        RECT 113.300 488.400 113.900 489.600 ;
        RECT 110.000 487.600 110.800 488.400 ;
        RECT 113.200 487.600 114.000 488.400 ;
        RECT 108.400 451.600 109.200 452.400 ;
        RECT 102.000 449.600 102.800 450.400 ;
        RECT 105.200 449.600 106.000 450.400 ;
        RECT 106.800 449.600 107.600 450.400 ;
        RECT 100.500 431.700 102.700 432.300 ;
        RECT 84.400 429.600 85.200 430.400 ;
        RECT 89.200 429.600 90.000 430.400 ;
        RECT 90.800 429.600 91.600 430.400 ;
        RECT 81.200 427.600 82.000 428.400 ;
        RECT 81.300 414.400 81.900 427.600 ;
        RECT 81.200 413.600 82.000 414.400 ;
        RECT 84.400 413.600 85.200 414.400 ;
        RECT 86.000 411.600 86.800 412.400 ;
        RECT 82.800 409.600 83.600 410.400 ;
        RECT 82.900 408.400 83.500 409.600 ;
        RECT 82.800 407.600 83.600 408.400 ;
        RECT 86.100 406.400 86.700 411.600 ;
        RECT 86.000 405.600 86.800 406.400 ;
        RECT 86.000 403.600 86.800 404.400 ;
        RECT 79.600 401.600 80.400 402.400 ;
        RECT 86.100 392.400 86.700 403.600 ;
        RECT 86.000 391.600 86.800 392.400 ;
        RECT 89.300 390.400 89.900 429.600 ;
        RECT 90.900 422.400 91.500 429.600 ;
        RECT 94.100 428.400 94.700 431.600 ;
        RECT 92.400 427.600 93.200 428.400 ;
        RECT 94.000 427.600 94.800 428.400 ;
        RECT 92.500 424.400 93.100 427.600 ;
        RECT 92.400 423.600 93.200 424.400 ;
        RECT 95.600 423.600 96.400 424.400 ;
        RECT 90.800 421.600 91.600 422.400 ;
        RECT 92.500 416.400 93.100 423.600 ;
        RECT 95.700 420.400 96.300 423.600 ;
        RECT 95.600 419.600 96.400 420.400 ;
        RECT 97.300 418.400 97.900 431.600 ;
        RECT 98.800 429.600 99.600 430.400 ;
        RECT 100.400 429.600 101.200 430.400 ;
        RECT 100.500 428.400 101.100 429.600 ;
        RECT 100.400 427.600 101.200 428.400 ;
        RECT 100.400 425.600 101.200 426.400 ;
        RECT 100.500 418.400 101.100 425.600 ;
        RECT 97.200 417.600 98.000 418.400 ;
        RECT 100.400 417.600 101.200 418.400 ;
        RECT 92.400 415.600 93.200 416.400 ;
        RECT 95.600 415.600 96.400 416.400 ;
        RECT 95.700 414.400 96.300 415.600 ;
        RECT 95.600 413.600 96.400 414.400 ;
        RECT 97.200 413.600 98.000 414.400 ;
        RECT 100.400 414.300 101.200 414.400 ;
        RECT 98.900 413.700 101.200 414.300 ;
        RECT 94.000 411.600 94.800 412.400 ;
        RECT 90.800 409.600 91.600 410.400 ;
        RECT 95.700 410.300 96.300 413.600 ;
        RECT 97.300 410.400 97.900 413.600 ;
        RECT 94.100 409.700 96.300 410.300 ;
        RECT 90.900 404.400 91.500 409.600 ;
        RECT 92.400 405.600 93.200 406.400 ;
        RECT 90.800 403.600 91.600 404.400 ;
        RECT 92.500 398.400 93.100 405.600 ;
        RECT 92.400 397.600 93.200 398.400 ;
        RECT 79.600 389.600 80.400 390.400 ;
        RECT 81.200 389.600 82.000 390.400 ;
        RECT 86.000 389.600 86.800 390.400 ;
        RECT 89.200 389.600 90.000 390.400 ;
        RECT 90.800 389.600 91.600 390.400 ;
        RECT 78.000 387.600 78.800 388.400 ;
        RECT 78.000 379.600 78.800 380.400 ;
        RECT 78.100 376.400 78.700 379.600 ;
        RECT 78.000 375.600 78.800 376.400 ;
        RECT 78.100 374.400 78.700 375.600 ;
        RECT 78.000 373.600 78.800 374.400 ;
        RECT 78.000 369.600 78.800 370.400 ;
        RECT 78.100 368.400 78.700 369.600 ;
        RECT 78.000 367.600 78.800 368.400 ;
        RECT 63.600 363.600 64.400 364.400 ;
        RECT 68.400 363.600 69.200 364.400 ;
        RECT 76.400 363.600 77.200 364.400 ;
        RECT 47.600 357.600 48.400 358.400 ;
        RECT 49.200 357.600 50.000 358.400 ;
        RECT 57.200 357.600 58.000 358.400 ;
        RECT 42.800 353.600 43.600 354.400 ;
        RECT 55.600 353.600 56.400 354.400 ;
        RECT 42.900 352.400 43.500 353.600 ;
        RECT 42.800 351.600 43.600 352.400 ;
        RECT 50.800 351.600 51.600 352.400 ;
        RECT 50.900 348.400 51.500 351.600 ;
        RECT 34.800 347.600 35.600 348.400 ;
        RECT 50.800 347.600 51.600 348.400 ;
        RECT 55.600 347.600 56.400 348.400 ;
        RECT 17.200 335.600 18.000 336.400 ;
        RECT 17.300 324.400 17.900 335.600 ;
        RECT 18.800 326.200 19.600 337.800 ;
        RECT 12.400 323.600 13.200 324.400 ;
        RECT 17.200 323.600 18.000 324.400 ;
        RECT 20.400 324.200 21.200 337.800 ;
        RECT 22.000 324.200 22.800 337.800 ;
        RECT 23.600 324.200 24.400 337.800 ;
        RECT 34.900 336.400 35.500 347.600 ;
        RECT 44.400 345.600 45.200 346.400 ;
        RECT 50.800 345.600 51.600 346.400 ;
        RECT 52.400 345.600 53.200 346.400 ;
        RECT 58.800 345.600 59.600 346.400 ;
        RECT 60.400 346.200 61.200 351.800 ;
        RECT 44.500 336.400 45.100 345.600 ;
        RECT 50.900 336.400 51.500 345.600 ;
        RECT 34.800 335.600 35.600 336.400 ;
        RECT 44.400 335.600 45.200 336.400 ;
        RECT 50.800 335.600 51.600 336.400 ;
        RECT 31.600 323.600 32.400 324.400 ;
        RECT 38.000 323.600 38.800 324.400 ;
        RECT 1.200 319.600 2.000 320.400 ;
        RECT 1.300 308.400 1.900 319.600 ;
        RECT 12.500 318.400 13.100 323.600 ;
        RECT 12.400 317.600 13.200 318.400 ;
        RECT 18.800 309.600 19.600 310.400 ;
        RECT 1.200 307.600 2.000 308.400 ;
        RECT 1.300 294.400 1.900 307.600 ;
        RECT 1.200 293.600 2.000 294.400 ;
        RECT 14.000 293.600 14.800 294.400 ;
        RECT 17.200 293.600 18.000 294.400 ;
        RECT 9.200 264.200 10.000 277.800 ;
        RECT 10.800 264.200 11.600 277.800 ;
        RECT 12.400 264.200 13.200 275.800 ;
        RECT 14.000 267.600 14.800 268.400 ;
        RECT 15.600 264.200 16.400 275.800 ;
        RECT 17.300 266.400 17.900 293.600 ;
        RECT 18.900 292.400 19.500 309.600 ;
        RECT 23.600 304.200 24.400 317.800 ;
        RECT 25.200 304.200 26.000 317.800 ;
        RECT 26.800 304.200 27.600 315.800 ;
        RECT 28.400 307.600 29.200 308.400 ;
        RECT 30.000 304.200 30.800 315.800 ;
        RECT 31.700 306.400 32.300 323.600 ;
        RECT 38.100 320.400 38.700 323.600 ;
        RECT 38.000 319.600 38.800 320.400 ;
        RECT 44.500 318.400 45.100 335.600 ;
        RECT 49.200 323.600 50.000 324.400 ;
        RECT 31.600 305.600 32.400 306.400 ;
        RECT 33.200 304.200 34.000 315.800 ;
        RECT 34.800 304.200 35.600 317.800 ;
        RECT 36.400 304.200 37.200 317.800 ;
        RECT 38.000 304.200 38.800 317.800 ;
        RECT 44.400 317.600 45.200 318.400 ;
        RECT 47.600 317.600 48.400 318.400 ;
        RECT 49.300 308.400 49.900 323.600 ;
        RECT 50.900 318.300 51.500 335.600 ;
        RECT 52.500 332.400 53.100 345.600 ;
        RECT 55.600 335.600 56.400 336.400 ;
        RECT 52.400 331.600 53.200 332.400 ;
        RECT 54.000 331.600 54.800 332.400 ;
        RECT 52.500 322.400 53.100 331.600 ;
        RECT 57.200 323.600 58.000 324.400 ;
        RECT 52.400 321.600 53.200 322.400 ;
        RECT 52.400 318.300 53.200 318.400 ;
        RECT 50.900 317.700 53.200 318.300 ;
        RECT 52.400 317.600 53.200 317.700 ;
        RECT 57.300 310.400 57.900 323.600 ;
        RECT 57.200 309.600 58.000 310.400 ;
        RECT 49.200 307.600 50.000 308.400 ;
        RECT 18.800 291.600 19.600 292.400 ;
        RECT 23.600 284.200 24.400 297.800 ;
        RECT 25.200 284.200 26.000 297.800 ;
        RECT 26.800 286.200 27.600 297.800 ;
        RECT 28.400 295.600 29.200 296.400 ;
        RECT 28.500 294.400 29.100 295.600 ;
        RECT 28.400 293.600 29.200 294.400 ;
        RECT 28.400 291.600 29.200 292.400 ;
        RECT 17.200 265.600 18.000 266.400 ;
        RECT 9.200 244.200 10.000 257.800 ;
        RECT 10.800 244.200 11.600 257.800 ;
        RECT 12.400 246.200 13.200 257.800 ;
        RECT 14.000 253.600 14.800 254.400 ;
        RECT 12.400 233.600 13.200 234.400 ;
        RECT 12.500 232.400 13.100 233.600 ;
        RECT 9.200 231.600 10.000 232.400 ;
        RECT 12.400 231.600 13.200 232.400 ;
        RECT 9.300 230.400 9.900 231.600 ;
        RECT 14.100 230.400 14.700 253.600 ;
        RECT 15.600 246.200 16.400 257.800 ;
        RECT 17.300 256.400 17.900 265.600 ;
        RECT 18.800 264.200 19.600 275.800 ;
        RECT 20.400 264.200 21.200 277.800 ;
        RECT 22.000 264.200 22.800 277.800 ;
        RECT 23.600 264.200 24.400 277.800 ;
        RECT 28.500 270.400 29.100 291.600 ;
        RECT 30.000 286.200 30.800 297.800 ;
        RECT 31.600 295.600 32.400 296.400 ;
        RECT 31.700 294.400 32.300 295.600 ;
        RECT 31.600 293.600 32.400 294.400 ;
        RECT 33.200 286.200 34.000 297.800 ;
        RECT 34.800 284.200 35.600 297.800 ;
        RECT 36.400 284.200 37.200 297.800 ;
        RECT 38.000 284.200 38.800 297.800 ;
        RECT 58.900 296.400 59.500 345.600 ;
        RECT 63.600 344.200 64.400 355.800 ;
        RECT 68.500 350.400 69.100 363.600 ;
        RECT 78.100 358.400 78.700 367.600 ;
        RECT 79.700 358.400 80.300 389.600 ;
        RECT 81.300 378.400 81.900 389.600 ;
        RECT 89.300 384.400 89.900 389.600 ;
        RECT 82.800 383.600 83.600 384.400 ;
        RECT 89.200 383.600 90.000 384.400 ;
        RECT 81.200 377.600 82.000 378.400 ;
        RECT 82.900 376.400 83.500 383.600 ;
        RECT 84.400 377.600 85.200 378.400 ;
        RECT 82.800 375.600 83.600 376.400 ;
        RECT 81.200 371.600 82.000 372.400 ;
        RECT 84.500 370.400 85.100 377.600 ;
        RECT 89.200 375.600 90.000 376.400 ;
        RECT 90.900 376.300 91.500 389.600 ;
        RECT 94.100 380.400 94.700 409.700 ;
        RECT 97.200 409.600 98.000 410.400 ;
        RECT 95.600 403.600 96.400 404.400 ;
        RECT 95.700 390.400 96.300 403.600 ;
        RECT 98.900 398.400 99.500 413.700 ;
        RECT 100.400 413.600 101.200 413.700 ;
        RECT 102.100 412.400 102.700 431.700 ;
        RECT 105.300 426.400 105.900 449.600 ;
        RECT 106.900 448.400 107.500 449.600 ;
        RECT 110.100 448.400 110.700 487.600 ;
        RECT 111.600 483.600 112.400 484.400 ;
        RECT 116.400 483.600 117.200 484.400 ;
        RECT 121.200 483.600 122.000 484.400 ;
        RECT 111.700 476.400 112.300 483.600 ;
        RECT 116.500 480.400 117.100 483.600 ;
        RECT 116.400 479.600 117.200 480.400 ;
        RECT 111.600 475.600 112.400 476.400 ;
        RECT 121.200 475.600 122.000 476.400 ;
        RECT 124.400 475.600 125.200 476.400 ;
        RECT 114.800 473.600 115.600 474.400 ;
        RECT 118.000 473.600 118.800 474.400 ;
        RECT 119.600 473.600 120.400 474.400 ;
        RECT 114.900 472.400 115.500 473.600 ;
        RECT 111.600 471.600 112.400 472.400 ;
        RECT 114.800 471.600 115.600 472.400 ;
        RECT 111.700 470.400 112.300 471.600 ;
        RECT 111.600 469.600 112.400 470.400 ;
        RECT 113.200 469.600 114.000 470.400 ;
        RECT 116.400 469.600 117.200 470.400 ;
        RECT 111.600 465.600 112.400 466.400 ;
        RECT 116.500 462.400 117.100 469.600 ;
        RECT 118.100 464.400 118.700 473.600 ;
        RECT 121.300 472.400 121.900 475.600 ;
        RECT 127.600 473.600 128.400 474.400 ;
        RECT 127.700 472.400 128.300 473.600 ;
        RECT 121.200 471.600 122.000 472.400 ;
        RECT 127.600 471.600 128.400 472.400 ;
        RECT 126.000 469.600 126.800 470.400 ;
        RECT 127.600 469.600 128.400 470.400 ;
        RECT 126.100 468.400 126.700 469.600 ;
        RECT 126.000 467.600 126.800 468.400 ;
        RECT 127.700 466.400 128.300 469.600 ;
        RECT 127.600 465.600 128.400 466.400 ;
        RECT 118.000 463.600 118.800 464.400 ;
        RECT 116.400 462.300 117.200 462.400 ;
        RECT 114.900 461.700 117.200 462.300 ;
        RECT 114.900 452.400 115.500 461.700 ;
        RECT 116.400 461.600 117.200 461.700 ;
        RECT 114.800 451.600 115.600 452.400 ;
        RECT 113.200 449.600 114.000 450.400 ;
        RECT 114.800 449.600 115.600 450.400 ;
        RECT 114.900 448.400 115.500 449.600 ;
        RECT 106.800 447.600 107.600 448.400 ;
        RECT 110.000 447.600 110.800 448.400 ;
        RECT 114.800 447.600 115.600 448.400 ;
        RECT 116.400 448.300 117.200 448.400 ;
        RECT 118.100 448.300 118.700 463.600 ;
        RECT 129.300 458.300 129.900 499.600 ;
        RECT 130.900 498.400 131.500 505.600 ;
        RECT 130.800 497.600 131.600 498.400 ;
        RECT 135.600 473.600 136.400 474.400 ;
        RECT 130.800 472.300 131.600 472.400 ;
        RECT 130.800 471.700 134.700 472.300 ;
        RECT 130.800 471.600 131.600 471.700 ;
        RECT 130.800 469.600 131.600 470.400 ;
        RECT 134.100 468.400 134.700 471.700 ;
        RECT 135.600 469.600 136.400 470.400 ;
        RECT 132.400 468.300 133.200 468.400 ;
        RECT 130.900 467.700 133.200 468.300 ;
        RECT 130.900 458.400 131.500 467.700 ;
        RECT 132.400 467.600 133.200 467.700 ;
        RECT 134.000 467.600 134.800 468.400 ;
        RECT 134.000 465.600 134.800 466.400 ;
        RECT 127.700 457.700 129.900 458.300 ;
        RECT 121.200 453.600 122.000 454.400 ;
        RECT 126.000 453.600 126.800 454.400 ;
        RECT 121.300 452.400 121.900 453.600 ;
        RECT 126.100 452.400 126.700 453.600 ;
        RECT 127.700 452.400 128.300 457.700 ;
        RECT 130.800 457.600 131.600 458.400 ;
        RECT 129.200 455.600 130.000 456.400 ;
        RECT 121.200 451.600 122.000 452.400 ;
        RECT 126.000 451.600 126.800 452.400 ;
        RECT 127.600 451.600 128.400 452.400 ;
        RECT 116.400 447.700 118.700 448.300 ;
        RECT 116.400 447.600 117.200 447.700 ;
        RECT 118.000 443.600 118.800 444.400 ;
        RECT 122.800 443.600 123.600 444.400 ;
        RECT 116.400 441.600 117.200 442.400 ;
        RECT 108.400 433.600 109.200 434.400 ;
        RECT 106.800 429.600 107.600 430.400 ;
        RECT 108.500 428.400 109.100 433.600 ;
        RECT 113.200 431.600 114.000 432.400 ;
        RECT 114.800 431.600 115.600 432.400 ;
        RECT 110.000 429.600 110.800 430.400 ;
        RECT 110.100 428.400 110.700 429.600 ;
        RECT 113.300 428.400 113.900 431.600 ;
        RECT 114.900 430.400 115.500 431.600 ;
        RECT 114.800 429.600 115.600 430.400 ;
        RECT 106.800 427.600 107.600 428.400 ;
        RECT 108.400 427.600 109.200 428.400 ;
        RECT 110.000 427.600 110.800 428.400 ;
        RECT 113.200 427.600 114.000 428.400 ;
        RECT 105.200 425.600 106.000 426.400 ;
        RECT 106.800 419.600 107.600 420.400 ;
        RECT 103.600 417.600 104.400 418.400 ;
        RECT 102.000 411.600 102.800 412.400 ;
        RECT 103.700 410.400 104.300 417.600 ;
        RECT 106.900 410.400 107.500 419.600 ;
        RECT 116.500 418.400 117.100 441.600 ;
        RECT 118.100 434.400 118.700 443.600 ;
        RECT 118.000 433.600 118.800 434.400 ;
        RECT 118.000 429.600 118.800 430.400 ;
        RECT 118.100 422.400 118.700 429.600 ;
        RECT 119.600 427.600 120.400 428.400 ;
        RECT 119.700 424.400 120.300 427.600 ;
        RECT 122.900 426.400 123.500 443.600 ;
        RECT 127.700 436.400 128.300 451.600 ;
        RECT 129.300 440.400 129.900 455.600 ;
        RECT 132.400 453.600 133.200 454.400 ;
        RECT 129.200 439.600 130.000 440.400 ;
        RECT 132.500 438.400 133.100 453.600 ;
        RECT 134.100 452.400 134.700 465.600 ;
        RECT 135.600 459.600 136.400 460.400 ;
        RECT 134.000 451.600 134.800 452.400 ;
        RECT 134.100 442.400 134.700 451.600 ;
        RECT 134.000 441.600 134.800 442.400 ;
        RECT 134.000 439.600 134.800 440.400 ;
        RECT 132.400 437.600 133.200 438.400 ;
        RECT 127.600 435.600 128.400 436.400 ;
        RECT 134.100 434.400 134.700 439.600 ;
        RECT 129.200 433.600 130.000 434.400 ;
        RECT 134.000 433.600 134.800 434.400 ;
        RECT 129.300 432.400 129.900 433.600 ;
        RECT 129.200 431.600 130.000 432.400 ;
        RECT 134.100 430.400 134.700 433.600 ;
        RECT 126.000 429.600 126.800 430.400 ;
        RECT 134.000 429.600 134.800 430.400 ;
        RECT 124.400 427.600 125.200 428.400 ;
        RECT 121.200 425.600 122.000 426.400 ;
        RECT 122.800 425.600 123.600 426.400 ;
        RECT 119.600 423.600 120.400 424.400 ;
        RECT 118.000 421.600 118.800 422.400 ;
        RECT 116.400 417.600 117.200 418.400 ;
        RECT 121.300 416.400 121.900 425.600 ;
        RECT 124.500 422.400 125.100 427.600 ;
        RECT 126.100 424.400 126.700 429.600 ;
        RECT 130.800 425.600 131.600 426.400 ;
        RECT 126.000 423.600 126.800 424.400 ;
        RECT 129.200 423.600 130.000 424.400 ;
        RECT 124.400 421.600 125.200 422.400 ;
        RECT 124.500 418.400 125.100 421.600 ;
        RECT 124.400 417.600 125.200 418.400 ;
        RECT 129.300 418.300 129.900 423.600 ;
        RECT 130.900 422.400 131.500 425.600 ;
        RECT 130.800 421.600 131.600 422.400 ;
        RECT 129.300 417.700 131.500 418.300 ;
        RECT 121.200 415.600 122.000 416.400 ;
        RECT 127.600 415.600 128.400 416.400 ;
        RECT 129.200 415.600 130.000 416.400 ;
        RECT 108.400 413.600 109.200 414.400 ;
        RECT 110.000 413.600 110.800 414.400 ;
        RECT 110.100 412.400 110.700 413.600 ;
        RECT 110.000 411.600 110.800 412.400 ;
        RECT 113.200 412.300 114.000 412.400 ;
        RECT 111.700 411.700 114.000 412.300 ;
        RECT 100.400 409.600 101.200 410.400 ;
        RECT 103.600 409.600 104.400 410.400 ;
        RECT 106.800 409.600 107.600 410.400 ;
        RECT 98.800 397.600 99.600 398.400 ;
        RECT 111.700 392.400 112.300 411.700 ;
        RECT 113.200 411.600 114.000 411.700 ;
        RECT 119.600 411.600 120.400 412.400 ;
        RECT 127.700 404.400 128.300 415.600 ;
        RECT 130.900 414.400 131.500 417.700 ;
        RECT 130.800 413.600 131.600 414.400 ;
        RECT 132.400 413.600 133.200 414.400 ;
        RECT 132.500 412.400 133.100 413.600 ;
        RECT 132.400 411.600 133.200 412.400 ;
        RECT 135.700 410.400 136.300 459.600 ;
        RECT 137.300 446.400 137.900 509.600 ;
        RECT 142.100 506.400 142.700 509.600 ;
        RECT 138.800 505.600 139.600 506.400 ;
        RECT 142.000 505.600 142.800 506.400 ;
        RECT 140.400 503.600 141.200 504.400 ;
        RECT 140.500 500.400 141.100 503.600 ;
        RECT 140.400 499.600 141.200 500.400 ;
        RECT 140.400 484.200 141.200 497.800 ;
        RECT 142.000 484.200 142.800 497.800 ;
        RECT 143.600 484.200 144.400 497.800 ;
        RECT 145.200 486.200 146.000 497.800 ;
        RECT 146.900 496.400 147.500 533.600 ;
        RECT 151.600 524.200 152.400 537.800 ;
        RECT 153.200 524.200 154.000 537.800 ;
        RECT 154.800 524.200 155.600 537.800 ;
        RECT 156.400 526.200 157.200 537.800 ;
        RECT 158.100 536.400 158.700 541.700 ;
        RECT 158.000 535.600 158.800 536.400 ;
        RECT 158.100 534.400 158.700 535.600 ;
        RECT 158.000 533.600 158.800 534.400 ;
        RECT 159.600 526.200 160.400 537.800 ;
        RECT 161.200 533.600 162.000 534.400 ;
        RECT 161.300 532.400 161.900 533.600 ;
        RECT 161.200 531.600 162.000 532.400 ;
        RECT 162.800 526.200 163.600 537.800 ;
        RECT 159.600 523.600 160.400 524.400 ;
        RECT 164.400 524.200 165.200 537.800 ;
        RECT 166.000 524.200 166.800 537.800 ;
        RECT 177.300 532.400 177.900 549.600 ;
        RECT 183.700 548.400 184.300 549.600 ;
        RECT 183.600 547.600 184.400 548.400 ;
        RECT 193.200 547.600 194.000 548.400 ;
        RECT 183.700 546.400 184.300 547.600 ;
        RECT 183.600 545.600 184.400 546.400 ;
        RECT 193.300 542.400 193.900 547.600 ;
        RECT 193.200 541.600 194.000 542.400 ;
        RECT 196.500 540.400 197.100 551.600 ;
        RECT 201.200 549.600 202.000 550.400 ;
        RECT 204.400 549.600 205.200 550.400 ;
        RECT 196.400 539.600 197.200 540.400 ;
        RECT 201.300 538.400 201.900 549.600 ;
        RECT 167.600 531.600 168.400 532.400 ;
        RECT 177.200 531.600 178.000 532.400 ;
        RECT 167.700 524.400 168.300 531.600 ;
        RECT 172.400 529.600 173.200 530.400 ;
        RECT 167.600 523.600 168.400 524.400 ;
        RECT 153.200 513.600 154.000 514.400 ;
        RECT 150.000 503.600 150.800 504.400 ;
        RECT 146.800 495.600 147.600 496.400 ;
        RECT 146.800 491.600 147.600 492.400 ;
        RECT 145.200 477.600 146.000 478.400 ;
        RECT 138.800 471.600 139.600 472.400 ;
        RECT 138.900 460.400 139.500 471.600 ;
        RECT 143.600 469.600 144.400 470.400 ;
        RECT 140.400 465.600 141.200 466.400 ;
        RECT 140.500 462.400 141.100 465.600 ;
        RECT 143.700 464.400 144.300 469.600 ;
        RECT 145.300 468.400 145.900 477.600 ;
        RECT 146.900 470.400 147.500 491.600 ;
        RECT 148.400 486.200 149.200 497.800 ;
        RECT 150.000 493.600 150.800 494.400 ;
        RECT 151.600 486.200 152.400 497.800 ;
        RECT 153.200 484.200 154.000 497.800 ;
        RECT 154.800 484.200 155.600 497.800 ;
        RECT 159.700 492.400 160.300 523.600 ;
        RECT 172.500 510.400 173.100 529.600 ;
        RECT 183.600 524.200 184.400 537.800 ;
        RECT 185.200 524.200 186.000 537.800 ;
        RECT 186.800 526.200 187.600 537.800 ;
        RECT 188.400 535.600 189.200 536.400 ;
        RECT 188.500 534.400 189.100 535.600 ;
        RECT 188.400 533.600 189.200 534.400 ;
        RECT 190.000 526.200 190.800 537.800 ;
        RECT 191.600 535.600 192.400 536.400 ;
        RECT 191.700 534.400 192.300 535.600 ;
        RECT 191.600 533.600 192.400 534.400 ;
        RECT 175.600 511.800 176.400 512.600 ;
        RECT 182.200 511.800 183.000 512.600 ;
        RECT 170.800 509.600 171.600 510.400 ;
        RECT 172.400 509.600 173.200 510.400 ;
        RECT 164.400 507.600 165.200 508.400 ;
        RECT 166.000 505.600 166.800 506.400 ;
        RECT 167.600 505.600 168.400 506.400 ;
        RECT 169.200 505.600 170.000 506.400 ;
        RECT 169.300 504.400 169.900 505.600 ;
        RECT 169.200 503.600 170.000 504.400 ;
        RECT 169.300 492.400 169.900 503.600 ;
        RECT 172.500 502.400 173.100 509.600 ;
        RECT 175.600 508.400 176.200 511.800 ;
        RECT 179.600 508.400 180.400 508.600 ;
        RECT 174.000 507.600 174.800 508.400 ;
        RECT 175.600 507.800 180.400 508.400 ;
        RECT 174.100 506.400 174.700 507.600 ;
        RECT 175.600 507.000 176.200 507.800 ;
        RECT 177.000 507.000 177.800 507.200 ;
        RECT 180.400 507.000 181.200 507.200 ;
        RECT 182.400 507.000 183.000 511.800 ;
        RECT 183.600 509.600 184.400 510.400 ;
        RECT 183.700 508.400 184.300 509.600 ;
        RECT 183.600 507.600 184.400 508.400 ;
        RECT 185.200 507.600 186.000 508.400 ;
        RECT 174.000 505.600 174.800 506.400 ;
        RECT 175.600 506.200 176.400 507.000 ;
        RECT 177.000 506.400 181.200 507.000 ;
        RECT 182.200 506.200 183.000 507.000 ;
        RECT 172.400 501.600 173.200 502.400 ;
        RECT 174.100 496.400 174.700 505.600 ;
        RECT 177.200 503.600 178.000 504.400 ;
        RECT 174.000 495.600 174.800 496.400 ;
        RECT 177.300 494.400 177.900 503.600 ;
        RECT 191.700 500.400 192.300 533.600 ;
        RECT 193.200 526.200 194.000 537.800 ;
        RECT 194.800 524.200 195.600 537.800 ;
        RECT 196.400 524.200 197.200 537.800 ;
        RECT 198.000 524.200 198.800 537.800 ;
        RECT 201.200 537.600 202.000 538.400 ;
        RECT 204.500 532.400 205.100 549.600 ;
        RECT 210.800 544.200 211.600 557.800 ;
        RECT 212.400 544.200 213.200 557.800 ;
        RECT 214.000 544.200 214.800 555.800 ;
        RECT 215.600 549.600 216.400 550.400 ;
        RECT 215.700 548.400 216.300 549.600 ;
        RECT 215.600 547.600 216.400 548.400 ;
        RECT 217.200 544.200 218.000 555.800 ;
        RECT 218.800 545.600 219.600 546.400 ;
        RECT 207.600 537.600 208.400 538.400 ;
        RECT 218.900 536.400 219.500 545.600 ;
        RECT 220.400 544.200 221.200 555.800 ;
        RECT 222.000 544.200 222.800 557.800 ;
        RECT 223.600 544.200 224.400 557.800 ;
        RECT 225.200 544.200 226.000 557.800 ;
        RECT 250.800 551.600 251.600 552.400 ;
        RECT 226.800 549.600 227.600 550.400 ;
        RECT 244.400 549.600 245.200 550.400 ;
        RECT 226.900 548.400 227.500 549.600 ;
        RECT 226.800 547.600 227.600 548.400 ;
        RECT 241.200 547.600 242.000 548.400 ;
        RECT 247.600 547.600 248.400 548.400 ;
        RECT 238.000 545.600 238.800 546.400 ;
        RECT 241.300 542.400 241.900 547.600 ;
        RECT 247.700 542.400 248.300 547.600 ;
        RECT 250.900 544.400 251.500 551.600 ;
        RECT 255.600 549.600 256.400 550.400 ;
        RECT 262.000 549.600 262.800 550.400 ;
        RECT 255.700 546.400 256.300 549.600 ;
        RECT 262.100 548.400 262.700 549.600 ;
        RECT 262.000 547.600 262.800 548.400 ;
        RECT 255.600 545.600 256.400 546.400 ;
        RECT 250.800 543.600 251.600 544.400 ;
        RECT 220.400 541.600 221.200 542.400 ;
        RECT 241.200 541.600 242.000 542.400 ;
        RECT 247.600 541.600 248.400 542.400 ;
        RECT 217.200 535.600 218.000 536.400 ;
        RECT 218.800 535.600 219.600 536.400 ;
        RECT 217.300 534.400 217.900 535.600 ;
        RECT 220.500 534.400 221.100 541.600 ;
        RECT 226.800 539.600 227.600 540.400 ;
        RECT 226.900 538.400 227.500 539.600 ;
        RECT 226.800 537.600 227.600 538.400 ;
        RECT 214.000 533.600 214.800 534.400 ;
        RECT 217.200 533.600 218.000 534.400 ;
        RECT 220.400 533.600 221.200 534.400 ;
        RECT 225.200 533.600 226.000 534.400 ;
        RECT 199.600 531.600 200.400 532.400 ;
        RECT 204.400 531.600 205.200 532.400 ;
        RECT 220.500 530.400 221.100 533.600 ;
        RECT 220.400 529.600 221.200 530.400 ;
        RECT 204.400 509.600 205.200 510.400 ;
        RECT 196.400 503.600 197.200 504.400 ;
        RECT 196.500 500.400 197.100 503.600 ;
        RECT 191.600 499.600 192.400 500.400 ;
        RECT 196.400 499.600 197.200 500.400 ;
        RECT 182.000 497.600 182.800 498.400 ;
        RECT 177.200 493.600 178.000 494.400 ;
        RECT 159.600 491.600 160.400 492.400 ;
        RECT 169.200 491.600 170.000 492.400 ;
        RECT 170.800 483.600 171.600 484.400 ;
        RECT 175.600 483.600 176.400 484.400 ;
        RECT 150.000 471.600 150.800 472.400 ;
        RECT 154.800 471.600 155.600 472.400 ;
        RECT 169.200 471.600 170.000 472.400 ;
        RECT 146.800 469.600 147.600 470.400 ;
        RECT 145.200 467.600 146.000 468.400 ;
        RECT 142.000 463.600 142.800 464.400 ;
        RECT 143.600 463.600 144.400 464.400 ;
        RECT 140.400 461.600 141.200 462.400 ;
        RECT 138.800 459.600 139.600 460.400 ;
        RECT 140.400 455.600 141.200 456.400 ;
        RECT 140.500 452.400 141.100 455.600 ;
        RECT 138.800 451.600 139.600 452.400 ;
        RECT 140.400 451.600 141.200 452.400 ;
        RECT 138.900 450.400 139.500 451.600 ;
        RECT 142.100 450.400 142.700 463.600 ;
        RECT 143.600 459.600 144.400 460.400 ;
        RECT 143.700 450.400 144.300 459.600 ;
        RECT 146.900 458.400 147.500 469.600 ;
        RECT 148.400 467.600 149.200 468.400 ;
        RECT 146.800 457.600 147.600 458.400 ;
        RECT 145.200 453.600 146.000 454.400 ;
        RECT 148.500 452.400 149.100 467.600 ;
        RECT 150.100 458.400 150.700 471.600 ;
        RECT 154.900 470.400 155.500 471.600 ;
        RECT 169.300 470.400 169.900 471.600 ;
        RECT 170.900 470.400 171.500 483.600 ;
        RECT 154.800 469.600 155.600 470.400 ;
        RECT 164.400 469.600 165.200 470.400 ;
        RECT 166.000 469.600 166.800 470.400 ;
        RECT 169.200 469.600 170.000 470.400 ;
        RECT 170.800 469.600 171.600 470.400 ;
        RECT 172.400 469.600 173.200 470.400 ;
        RECT 174.000 469.600 174.800 470.400 ;
        RECT 153.200 465.600 154.000 466.400 ;
        RECT 150.000 457.600 150.800 458.400 ;
        RECT 148.400 451.600 149.200 452.400 ;
        RECT 138.800 449.600 139.600 450.400 ;
        RECT 142.000 449.600 142.800 450.400 ;
        RECT 143.600 449.600 144.400 450.400 ;
        RECT 148.400 449.600 149.200 450.400 ;
        RECT 137.200 445.600 138.000 446.400 ;
        RECT 140.400 443.600 141.200 444.400 ;
        RECT 140.500 436.400 141.100 443.600 ;
        RECT 137.200 435.600 138.000 436.400 ;
        RECT 137.300 412.400 137.900 435.600 ;
        RECT 138.800 424.200 139.600 435.800 ;
        RECT 140.400 435.600 141.200 436.400 ;
        RECT 142.100 418.400 142.700 449.600 ;
        RECT 154.900 444.400 155.500 469.600 ;
        RECT 162.800 467.600 163.600 468.400 ;
        RECT 159.600 457.600 160.400 458.400 ;
        RECT 156.400 451.600 157.200 452.400 ;
        RECT 154.800 443.600 155.600 444.400 ;
        RECT 145.200 431.600 146.000 432.400 ;
        RECT 146.800 431.600 147.600 432.400 ;
        RECT 145.300 430.400 145.900 431.600 ;
        RECT 145.200 429.600 146.000 430.400 ;
        RECT 142.000 417.600 142.800 418.400 ;
        RECT 138.800 413.600 139.600 414.400 ;
        RECT 145.200 413.600 146.000 414.400 ;
        RECT 138.900 412.400 139.500 413.600 ;
        RECT 146.900 412.400 147.500 431.600 ;
        RECT 148.400 424.200 149.200 435.800 ;
        RECT 156.500 432.400 157.100 451.600 ;
        RECT 158.000 443.600 158.800 444.400 ;
        RECT 158.100 432.400 158.700 443.600 ;
        RECT 150.000 427.600 150.800 428.400 ;
        RECT 150.100 420.400 150.700 427.600 ;
        RECT 151.600 426.200 152.400 431.800 ;
        RECT 156.400 431.600 157.200 432.400 ;
        RECT 158.000 431.600 158.800 432.400 ;
        RECT 156.400 429.600 157.200 430.400 ;
        RECT 156.500 428.400 157.100 429.600 ;
        RECT 156.400 427.600 157.200 428.400 ;
        RECT 158.000 427.600 158.800 428.400 ;
        RECT 150.000 419.600 150.800 420.400 ;
        RECT 150.000 417.600 150.800 418.400 ;
        RECT 137.200 411.600 138.000 412.400 ;
        RECT 138.800 411.600 139.600 412.400 ;
        RECT 146.800 411.600 147.600 412.400 ;
        RECT 135.600 409.600 136.400 410.400 ;
        RECT 127.600 403.600 128.400 404.400 ;
        RECT 132.400 403.600 133.200 404.400 ;
        RECT 97.200 391.600 98.000 392.400 ;
        RECT 106.800 391.600 107.600 392.400 ;
        RECT 111.600 391.600 112.400 392.400 ;
        RECT 97.300 390.400 97.900 391.600 ;
        RECT 106.900 390.400 107.500 391.600 ;
        RECT 111.700 390.400 112.300 391.600 ;
        RECT 95.600 389.600 96.400 390.400 ;
        RECT 97.200 389.600 98.000 390.400 ;
        RECT 106.800 389.600 107.600 390.400 ;
        RECT 108.400 389.600 109.200 390.400 ;
        RECT 111.600 389.600 112.400 390.400 ;
        RECT 98.800 387.600 99.600 388.400 ;
        RECT 94.000 379.600 94.800 380.400 ;
        RECT 92.400 377.600 93.200 378.400 ;
        RECT 90.900 375.700 93.100 376.300 ;
        RECT 89.300 372.400 89.900 375.600 ;
        RECT 90.800 373.600 91.600 374.400 ;
        RECT 89.200 371.600 90.000 372.400 ;
        RECT 84.400 369.600 85.200 370.400 ;
        RECT 89.200 369.600 90.000 370.400 ;
        RECT 90.900 366.400 91.500 373.600 ;
        RECT 90.800 365.600 91.600 366.400 ;
        RECT 90.800 363.600 91.600 364.400 ;
        RECT 78.000 357.600 78.800 358.400 ;
        RECT 79.600 357.600 80.400 358.400 ;
        RECT 68.400 349.600 69.200 350.400 ;
        RECT 68.400 347.600 69.200 348.400 ;
        RECT 60.400 341.600 61.200 342.400 ;
        RECT 60.500 338.400 61.100 341.600 ;
        RECT 60.400 337.600 61.200 338.400 ;
        RECT 68.500 336.400 69.100 347.600 ;
        RECT 73.200 344.200 74.000 355.800 ;
        RECT 90.900 352.400 91.500 363.600 ;
        RECT 81.200 351.600 82.000 352.400 ;
        RECT 90.800 351.600 91.600 352.400 ;
        RECT 92.500 350.400 93.100 375.700 ;
        RECT 97.200 366.200 98.000 377.800 ;
        RECT 94.000 353.600 94.800 354.400 ;
        RECT 97.200 353.600 98.000 354.400 ;
        RECT 94.100 352.400 94.700 353.600 ;
        RECT 94.000 351.600 94.800 352.400 ;
        RECT 90.800 349.600 91.600 350.400 ;
        RECT 92.400 349.600 93.200 350.400 ;
        RECT 86.000 347.600 86.800 348.400 ;
        RECT 81.200 345.600 82.000 346.400 ;
        RECT 81.300 342.400 81.900 345.600 ;
        RECT 81.200 341.600 82.000 342.400 ;
        RECT 90.900 340.400 91.500 349.600 ;
        RECT 98.900 348.400 99.500 387.600 ;
        RECT 100.400 385.600 101.200 386.400 ;
        RECT 111.600 385.600 112.400 386.400 ;
        RECT 113.200 386.200 114.000 391.800 ;
        RECT 114.800 387.600 115.600 388.400 ;
        RECT 100.500 368.400 101.100 385.600 ;
        RECT 103.600 383.600 104.400 384.400 ;
        RECT 103.700 372.400 104.300 383.600 ;
        RECT 108.400 381.600 109.200 382.400 ;
        RECT 102.000 371.600 102.800 372.400 ;
        RECT 103.600 371.600 104.400 372.400 ;
        RECT 102.100 370.400 102.700 371.600 ;
        RECT 102.000 369.600 102.800 370.400 ;
        RECT 100.400 367.600 101.200 368.400 ;
        RECT 106.800 366.200 107.600 377.800 ;
        RECT 108.500 374.400 109.100 381.600 ;
        RECT 111.600 379.600 112.400 380.400 ;
        RECT 111.700 376.400 112.300 379.600 ;
        RECT 114.900 378.400 115.500 387.600 ;
        RECT 116.400 384.200 117.200 395.800 ;
        RECT 118.000 389.600 118.800 390.400 ;
        RECT 119.600 389.600 120.400 390.400 ;
        RECT 114.800 377.600 115.600 378.400 ;
        RECT 108.400 373.600 109.200 374.400 ;
        RECT 110.000 370.200 110.800 375.800 ;
        RECT 111.600 375.600 112.400 376.400 ;
        RECT 118.100 372.400 118.700 389.600 ;
        RECT 121.200 387.600 122.000 388.400 ;
        RECT 121.300 386.400 121.900 387.600 ;
        RECT 119.600 385.600 120.400 386.400 ;
        RECT 121.200 385.600 122.000 386.400 ;
        RECT 119.700 374.400 120.300 385.600 ;
        RECT 121.300 382.400 121.900 385.600 ;
        RECT 126.000 384.200 126.800 395.800 ;
        RECT 132.500 394.400 133.100 403.600 ;
        RECT 130.800 393.600 131.600 394.400 ;
        RECT 132.400 393.600 133.200 394.400 ;
        RECT 130.900 392.400 131.500 393.600 ;
        RECT 130.800 391.600 131.600 392.400 ;
        RECT 137.200 392.300 138.000 392.400 ;
        RECT 138.900 392.300 139.500 411.600 ;
        RECT 142.000 403.600 142.800 404.400 ;
        RECT 137.200 391.700 139.500 392.300 ;
        RECT 137.200 391.600 138.000 391.700 ;
        RECT 142.100 390.400 142.700 403.600 ;
        RECT 134.000 389.600 134.800 390.400 ;
        RECT 138.800 389.600 139.600 390.400 ;
        RECT 142.000 389.600 142.800 390.400 ;
        RECT 132.400 387.600 133.200 388.400 ;
        RECT 127.600 383.600 128.400 384.400 ;
        RECT 121.200 381.600 122.000 382.400 ;
        RECT 119.600 373.600 120.400 374.400 ;
        RECT 121.200 373.600 122.000 374.400 ;
        RECT 124.400 373.600 125.200 374.400 ;
        RECT 118.000 371.600 118.800 372.400 ;
        RECT 119.700 358.400 120.300 373.600 ;
        RECT 121.200 371.600 122.000 372.400 ;
        RECT 122.800 371.600 123.600 372.400 ;
        RECT 119.600 357.600 120.400 358.400 ;
        RECT 105.200 351.600 106.000 352.400 ;
        RECT 113.200 351.600 114.000 352.400 ;
        RECT 119.600 351.600 120.400 352.400 ;
        RECT 105.300 350.400 105.900 351.600 ;
        RECT 113.300 350.400 113.900 351.600 ;
        RECT 103.600 349.600 104.400 350.400 ;
        RECT 105.200 349.600 106.000 350.400 ;
        RECT 113.200 349.600 114.000 350.400 ;
        RECT 114.800 349.600 115.600 350.400 ;
        RECT 92.400 347.600 93.200 348.400 ;
        RECT 98.800 347.600 99.600 348.400 ;
        RECT 111.600 347.600 112.400 348.400 ;
        RECT 113.200 347.600 114.000 348.400 ;
        RECT 102.000 345.600 102.800 346.400 ;
        RECT 111.700 346.300 112.300 347.600 ;
        RECT 114.900 346.300 115.500 349.600 ;
        RECT 116.400 347.600 117.200 348.400 ;
        RECT 111.700 345.700 115.500 346.300 ;
        RECT 94.000 341.600 94.800 342.400 ;
        RECT 90.800 339.600 91.600 340.400 ;
        RECT 68.400 335.600 69.200 336.400 ;
        RECT 60.400 321.600 61.200 322.400 ;
        RECT 57.200 295.600 58.000 296.400 ;
        RECT 58.800 295.600 59.600 296.400 ;
        RECT 58.800 293.600 59.600 294.400 ;
        RECT 54.000 291.600 54.800 292.400 ;
        RECT 54.100 290.400 54.700 291.600 ;
        RECT 58.900 290.400 59.500 293.600 ;
        RECT 60.500 292.400 61.100 321.600 ;
        RECT 62.000 304.200 62.800 317.800 ;
        RECT 63.600 304.200 64.400 317.800 ;
        RECT 65.200 304.200 66.000 317.800 ;
        RECT 66.800 304.200 67.600 315.800 ;
        RECT 68.500 306.400 69.100 335.600 ;
        RECT 70.000 324.200 70.800 337.800 ;
        RECT 71.600 324.200 72.400 337.800 ;
        RECT 73.200 324.200 74.000 337.800 ;
        RECT 74.800 326.200 75.600 337.800 ;
        RECT 76.400 335.600 77.200 336.400 ;
        RECT 78.000 326.200 78.800 337.800 ;
        RECT 79.600 333.600 80.400 334.400 ;
        RECT 79.600 331.600 80.400 332.400 ;
        RECT 68.400 305.600 69.200 306.400 ;
        RECT 70.000 304.200 70.800 315.800 ;
        RECT 71.600 307.600 72.400 308.400 ;
        RECT 73.200 304.200 74.000 315.800 ;
        RECT 74.800 304.200 75.600 317.800 ;
        RECT 76.400 304.200 77.200 317.800 ;
        RECT 79.700 312.400 80.300 331.600 ;
        RECT 81.200 326.200 82.000 337.800 ;
        RECT 82.800 324.200 83.600 337.800 ;
        RECT 84.400 324.200 85.200 337.800 ;
        RECT 94.100 336.400 94.700 341.600 ;
        RECT 94.000 335.600 94.800 336.400 ;
        RECT 97.200 333.600 98.000 334.400 ;
        RECT 95.600 331.600 96.400 332.400 ;
        RECT 79.600 311.600 80.400 312.400 ;
        RECT 79.700 310.400 80.300 311.600 ;
        RECT 95.700 310.400 96.300 331.600 ;
        RECT 102.100 318.400 102.700 345.600 ;
        RECT 103.600 331.600 104.400 332.400 ;
        RECT 105.200 331.600 106.000 332.400 ;
        RECT 103.700 322.400 104.300 331.600 ;
        RECT 106.800 330.200 107.600 335.800 ;
        RECT 108.400 335.600 109.200 336.400 ;
        RECT 108.500 334.400 109.100 335.600 ;
        RECT 108.400 333.600 109.200 334.400 ;
        RECT 110.000 326.200 110.800 337.800 ;
        RECT 116.500 332.400 117.100 347.600 ;
        RECT 119.700 342.400 120.300 351.600 ;
        RECT 121.300 350.300 121.900 371.600 ;
        RECT 122.800 363.600 123.600 364.400 ;
        RECT 122.900 352.400 123.500 363.600 ;
        RECT 122.800 351.600 123.600 352.400 ;
        RECT 122.800 350.300 123.600 350.400 ;
        RECT 121.300 349.700 123.600 350.300 ;
        RECT 122.800 349.600 123.600 349.700 ;
        RECT 124.500 348.400 125.100 373.600 ;
        RECT 127.700 372.400 128.300 383.600 ;
        RECT 132.500 380.400 133.100 387.600 ;
        RECT 134.100 384.400 134.700 389.600 ;
        RECT 138.900 388.400 139.500 389.600 ;
        RECT 138.800 387.600 139.600 388.400 ;
        RECT 143.600 387.600 144.400 388.400 ;
        RECT 134.000 383.600 134.800 384.400 ;
        RECT 138.800 383.600 139.600 384.400 ;
        RECT 132.400 379.600 133.200 380.400 ;
        RECT 129.200 375.600 130.000 376.400 ;
        RECT 129.300 372.400 129.900 375.600 ;
        RECT 137.200 373.600 138.000 374.400 ;
        RECT 138.900 372.400 139.500 383.600 ;
        RECT 142.000 377.600 142.800 378.400 ;
        RECT 142.000 375.600 142.800 376.400 ;
        RECT 142.100 372.400 142.700 375.600 ;
        RECT 143.700 374.400 144.300 387.600 ;
        RECT 143.600 373.600 144.400 374.400 ;
        RECT 127.600 371.600 128.400 372.400 ;
        RECT 129.200 371.600 130.000 372.400 ;
        RECT 137.200 371.600 138.000 372.400 ;
        RECT 138.800 371.600 139.600 372.400 ;
        RECT 142.000 371.600 142.800 372.400 ;
        RECT 126.000 369.600 126.800 370.400 ;
        RECT 126.100 364.400 126.700 369.600 ;
        RECT 126.000 363.600 126.800 364.400 ;
        RECT 126.000 351.600 126.800 352.400 ;
        RECT 127.700 350.400 128.300 371.600 ;
        RECT 138.900 370.400 139.500 371.600 ;
        RECT 142.100 370.400 142.700 371.600 ;
        RECT 138.800 369.600 139.600 370.400 ;
        RECT 142.000 369.600 142.800 370.400 ;
        RECT 132.400 367.600 133.200 368.400 ;
        RECT 143.700 366.400 144.300 373.600 ;
        RECT 145.200 371.600 146.000 372.400 ;
        RECT 145.300 368.400 145.900 371.600 ;
        RECT 145.200 367.600 146.000 368.400 ;
        RECT 130.800 365.600 131.600 366.400 ;
        RECT 143.600 365.600 144.400 366.400 ;
        RECT 127.600 349.600 128.400 350.400 ;
        RECT 129.200 349.600 130.000 350.400 ;
        RECT 124.400 347.600 125.200 348.400 ;
        RECT 127.600 347.600 128.400 348.400 ;
        RECT 119.600 341.600 120.400 342.400 ;
        RECT 124.400 341.600 125.200 342.400 ;
        RECT 124.500 338.400 125.100 341.600 ;
        RECT 116.400 331.600 117.200 332.400 ;
        RECT 119.600 326.200 120.400 337.800 ;
        RECT 124.400 337.600 125.200 338.400 ;
        RECT 126.000 330.200 126.800 335.800 ;
        RECT 127.700 332.400 128.300 347.600 ;
        RECT 129.300 344.400 129.900 349.600 ;
        RECT 130.900 348.400 131.500 365.600 ;
        RECT 142.000 363.600 142.800 364.400 ;
        RECT 134.000 353.600 134.800 354.400 ;
        RECT 134.100 350.400 134.700 353.600 ;
        RECT 142.100 350.400 142.700 363.600 ;
        RECT 146.900 354.400 147.500 411.600 ;
        RECT 150.100 410.400 150.700 417.600 ;
        RECT 156.400 415.600 157.200 416.400 ;
        RECT 156.500 414.400 157.100 415.600 ;
        RECT 156.400 413.600 157.200 414.400 ;
        RECT 156.400 411.600 157.200 412.400 ;
        RECT 158.000 412.300 158.800 412.400 ;
        RECT 159.700 412.300 160.300 457.600 ;
        RECT 161.200 451.600 162.000 452.400 ;
        RECT 162.800 451.600 163.600 452.400 ;
        RECT 161.300 450.400 161.900 451.600 ;
        RECT 161.200 449.600 162.000 450.400 ;
        RECT 162.800 449.600 163.600 450.400 ;
        RECT 162.900 432.400 163.500 449.600 ;
        RECT 164.500 446.400 165.100 469.600 ;
        RECT 166.000 463.600 166.800 464.400 ;
        RECT 166.100 448.400 166.700 463.600 ;
        RECT 167.600 461.600 168.400 462.400 ;
        RECT 167.700 456.400 168.300 461.600 ;
        RECT 167.600 455.600 168.400 456.400 ;
        RECT 170.900 456.300 171.500 469.600 ;
        RECT 172.400 467.600 173.200 468.400 ;
        RECT 169.300 455.700 171.500 456.300 ;
        RECT 167.700 452.400 168.300 455.600 ;
        RECT 169.300 452.400 169.900 455.700 ;
        RECT 174.100 454.400 174.700 469.600 ;
        RECT 175.700 456.400 176.300 483.600 ;
        RECT 178.800 475.600 179.600 476.400 ;
        RECT 177.200 471.600 178.000 472.400 ;
        RECT 177.300 470.400 177.900 471.600 ;
        RECT 177.200 469.600 178.000 470.400 ;
        RECT 178.900 468.400 179.500 475.600 ;
        RECT 182.100 470.400 182.700 497.600 ;
        RECT 183.600 491.600 184.400 492.400 ;
        RECT 185.200 484.200 186.000 497.800 ;
        RECT 186.800 484.200 187.600 497.800 ;
        RECT 188.400 484.200 189.200 497.800 ;
        RECT 190.000 486.200 190.800 497.800 ;
        RECT 191.700 496.400 192.300 499.600 ;
        RECT 191.600 495.600 192.400 496.400 ;
        RECT 193.200 486.200 194.000 497.800 ;
        RECT 194.800 493.600 195.600 494.400 ;
        RECT 196.400 486.200 197.200 497.800 ;
        RECT 198.000 484.200 198.800 497.800 ;
        RECT 199.600 484.200 200.400 497.800 ;
        RECT 201.200 495.600 202.000 496.400 ;
        RECT 185.200 473.600 186.000 474.400 ;
        RECT 185.300 472.400 185.900 473.600 ;
        RECT 183.600 471.600 184.400 472.400 ;
        RECT 185.200 471.600 186.000 472.400 ;
        RECT 180.400 469.600 181.200 470.400 ;
        RECT 182.000 469.600 182.800 470.400 ;
        RECT 177.200 467.600 178.000 468.400 ;
        RECT 178.800 467.600 179.600 468.400 ;
        RECT 180.500 466.400 181.100 469.600 ;
        RECT 183.700 466.400 184.300 471.600 ;
        RECT 180.400 465.600 181.200 466.400 ;
        RECT 183.600 465.600 184.400 466.400 ;
        RECT 183.700 460.400 184.300 465.600 ;
        RECT 185.300 460.400 185.900 471.600 ;
        RECT 190.000 464.200 190.800 475.800 ;
        RECT 196.400 469.600 197.200 470.400 ;
        RECT 196.500 468.400 197.100 469.600 ;
        RECT 196.400 467.600 197.200 468.400 ;
        RECT 199.600 464.200 200.400 475.800 ;
        RECT 201.300 468.400 201.900 495.600 ;
        RECT 204.500 492.400 205.100 509.600 ;
        RECT 207.600 504.200 208.400 517.800 ;
        RECT 209.200 504.200 210.000 517.800 ;
        RECT 210.800 504.200 211.600 515.800 ;
        RECT 212.400 507.600 213.200 508.400 ;
        RECT 204.400 491.600 205.200 492.400 ;
        RECT 209.200 487.600 210.000 488.400 ;
        RECT 201.200 467.600 202.000 468.400 ;
        RECT 202.800 466.200 203.600 471.800 ;
        RECT 204.400 469.600 205.200 470.400 ;
        RECT 204.500 468.400 205.100 469.600 ;
        RECT 209.300 468.400 209.900 487.600 ;
        RECT 212.500 484.400 213.100 507.600 ;
        RECT 214.000 504.200 214.800 515.800 ;
        RECT 215.600 505.600 216.400 506.400 ;
        RECT 215.700 500.400 216.300 505.600 ;
        RECT 217.200 504.200 218.000 515.800 ;
        RECT 218.800 504.200 219.600 517.800 ;
        RECT 220.400 504.200 221.200 517.800 ;
        RECT 222.000 504.200 222.800 517.800 ;
        RECT 223.600 509.600 224.400 510.400 ;
        RECT 223.700 502.400 224.300 509.600 ;
        RECT 225.300 504.400 225.900 533.600 ;
        RECT 226.800 523.600 227.600 524.400 ;
        RECT 233.200 523.600 234.000 524.400 ;
        RECT 236.400 524.200 237.200 537.800 ;
        RECT 238.000 524.200 238.800 537.800 ;
        RECT 239.600 524.200 240.400 537.800 ;
        RECT 241.200 526.200 242.000 537.800 ;
        RECT 242.800 535.600 243.600 536.400 ;
        RECT 242.800 533.600 243.600 534.400 ;
        RECT 233.300 514.400 233.900 523.600 ;
        RECT 242.900 518.400 243.500 533.600 ;
        RECT 244.400 526.200 245.200 537.800 ;
        RECT 246.000 533.600 246.800 534.400 ;
        RECT 247.600 526.200 248.400 537.800 ;
        RECT 249.200 524.200 250.000 537.800 ;
        RECT 250.800 524.200 251.600 537.800 ;
        RECT 252.400 531.600 253.200 532.400 ;
        RECT 262.100 532.300 262.700 547.600 ;
        RECT 265.200 544.200 266.000 557.800 ;
        RECT 266.800 544.200 267.600 557.800 ;
        RECT 268.400 544.200 269.200 555.800 ;
        RECT 270.000 547.600 270.800 548.400 ;
        RECT 270.100 540.400 270.700 547.600 ;
        RECT 271.600 544.200 272.400 555.800 ;
        RECT 273.200 545.600 274.000 546.400 ;
        RECT 270.000 539.600 270.800 540.400 ;
        RECT 265.200 535.600 266.000 536.400 ;
        RECT 263.600 532.300 264.400 532.400 ;
        RECT 262.100 531.700 264.400 532.300 ;
        RECT 242.800 517.600 243.600 518.400 ;
        RECT 233.200 513.600 234.000 514.400 ;
        RECT 244.400 511.600 245.200 512.400 ;
        RECT 236.400 509.600 237.200 510.400 ;
        RECT 238.000 509.600 238.800 510.400 ;
        RECT 241.200 509.600 242.000 510.400 ;
        RECT 238.100 506.400 238.700 509.600 ;
        RECT 241.300 508.400 241.900 509.600 ;
        RECT 239.600 507.600 240.400 508.400 ;
        RECT 241.200 507.600 242.000 508.400 ;
        RECT 238.000 505.600 238.800 506.400 ;
        RECT 241.200 505.600 242.000 506.400 ;
        RECT 225.200 503.600 226.000 504.400 ;
        RECT 231.600 503.600 232.400 504.400 ;
        RECT 236.400 503.600 237.200 504.400 ;
        RECT 223.600 501.600 224.400 502.400 ;
        RECT 215.600 499.600 216.400 500.400 ;
        RECT 214.000 493.600 214.800 494.400 ;
        RECT 212.400 483.600 213.200 484.400 ;
        RECT 214.100 478.400 214.700 493.600 ;
        RECT 220.400 484.200 221.200 497.800 ;
        RECT 222.000 484.200 222.800 497.800 ;
        RECT 223.600 484.200 224.400 497.800 ;
        RECT 225.200 486.200 226.000 497.800 ;
        RECT 226.800 495.600 227.600 496.400 ;
        RECT 228.400 486.200 229.200 497.800 ;
        RECT 230.000 493.600 230.800 494.400 ;
        RECT 225.200 483.600 226.000 484.400 ;
        RECT 214.000 477.600 214.800 478.400 ;
        RECT 210.800 471.600 211.600 472.400 ;
        RECT 218.800 471.600 219.600 472.400 ;
        RECT 223.600 471.600 224.400 472.400 ;
        RECT 218.900 470.400 219.500 471.600 ;
        RECT 214.000 469.600 214.800 470.400 ;
        RECT 218.800 469.600 219.600 470.400 ;
        RECT 222.000 469.600 222.800 470.400 ;
        RECT 204.400 467.600 205.200 468.400 ;
        RECT 209.200 467.600 210.000 468.400 ;
        RECT 212.400 467.600 213.200 468.400 ;
        RECT 183.600 459.600 184.400 460.400 ;
        RECT 185.200 459.600 186.000 460.400 ;
        RECT 196.400 459.600 197.200 460.400 ;
        RECT 177.200 457.600 178.000 458.400 ;
        RECT 175.600 455.600 176.400 456.400 ;
        RECT 177.300 454.400 177.900 457.600 ;
        RECT 170.800 453.600 171.600 454.400 ;
        RECT 174.000 453.600 174.800 454.400 ;
        RECT 177.200 453.600 178.000 454.400 ;
        RECT 167.600 451.600 168.400 452.400 ;
        RECT 169.200 451.600 170.000 452.400 ;
        RECT 169.200 449.600 170.000 450.400 ;
        RECT 166.000 447.600 166.800 448.400 ;
        RECT 164.400 445.600 165.200 446.400 ;
        RECT 167.600 443.600 168.400 444.400 ;
        RECT 167.700 438.400 168.300 443.600 ;
        RECT 167.600 437.600 168.400 438.400 ;
        RECT 167.600 433.600 168.400 434.400 ;
        RECT 162.800 431.600 163.600 432.400 ;
        RECT 167.600 431.600 168.400 432.400 ;
        RECT 167.700 430.400 168.300 431.600 ;
        RECT 167.600 429.600 168.400 430.400 ;
        RECT 170.900 428.400 171.500 453.600 ;
        RECT 172.400 451.600 173.200 452.400 ;
        RECT 175.600 451.600 176.400 452.400 ;
        RECT 180.400 451.600 181.200 452.400 ;
        RECT 172.500 430.400 173.100 451.600 ;
        RECT 175.700 450.400 176.300 451.600 ;
        RECT 175.600 449.600 176.400 450.400 ;
        RECT 177.200 443.600 178.000 444.400 ;
        RECT 175.600 432.300 176.400 432.400 ;
        RECT 177.300 432.300 177.900 443.600 ;
        RECT 180.500 438.400 181.100 451.600 ;
        RECT 182.000 446.200 182.800 457.800 ;
        RECT 185.300 454.400 185.900 459.600 ;
        RECT 185.200 453.600 186.000 454.400 ;
        RECT 188.400 451.600 189.200 452.400 ;
        RECT 183.600 449.600 184.400 450.400 ;
        RECT 183.700 438.400 184.300 449.600 ;
        RECT 191.600 446.200 192.400 457.800 ;
        RECT 193.200 453.600 194.000 454.400 ;
        RECT 180.400 437.600 181.200 438.400 ;
        RECT 183.600 437.600 184.400 438.400 ;
        RECT 175.600 431.700 177.900 432.300 ;
        RECT 175.600 431.600 176.400 431.700 ;
        RECT 172.400 429.600 173.200 430.400 ;
        RECT 180.400 429.600 181.200 430.400 ;
        RECT 169.200 427.600 170.000 428.400 ;
        RECT 170.800 427.600 171.600 428.400 ;
        RECT 169.300 426.400 169.900 427.600 ;
        RECT 169.200 425.600 170.000 426.400 ;
        RECT 164.400 421.600 165.200 422.400 ;
        RECT 161.200 415.600 162.000 416.400 ;
        RECT 162.800 413.600 163.600 414.400 ;
        RECT 158.000 411.700 160.300 412.300 ;
        RECT 158.000 411.600 158.800 411.700 ;
        RECT 148.400 409.600 149.200 410.400 ;
        RECT 150.000 409.600 150.800 410.400 ;
        RECT 156.500 390.400 157.100 411.600 ;
        RECT 161.200 409.600 162.000 410.400 ;
        RECT 161.200 407.600 162.000 408.400 ;
        RECT 158.000 405.600 158.800 406.400 ;
        RECT 158.100 398.400 158.700 405.600 ;
        RECT 161.300 398.400 161.900 407.600 ;
        RECT 162.900 406.400 163.500 413.600 ;
        RECT 164.500 412.400 165.100 421.600 ;
        RECT 167.600 413.600 168.400 414.400 ;
        RECT 164.400 411.600 165.200 412.400 ;
        RECT 169.200 411.600 170.000 412.400 ;
        RECT 167.600 409.600 168.400 410.400 ;
        RECT 170.900 408.400 171.500 427.600 ;
        RECT 172.400 425.600 173.200 426.400 ;
        RECT 172.500 418.400 173.100 425.600 ;
        RECT 180.500 424.400 181.100 429.600 ;
        RECT 182.000 427.600 182.800 428.400 ;
        RECT 182.100 426.400 182.700 427.600 ;
        RECT 182.000 425.600 182.800 426.400 ;
        RECT 180.400 423.600 181.200 424.400 ;
        RECT 188.400 424.200 189.200 435.800 ;
        RECT 193.300 428.400 193.900 453.600 ;
        RECT 194.800 450.200 195.600 455.800 ;
        RECT 196.500 450.400 197.100 459.600 ;
        RECT 198.000 455.600 198.800 456.400 ;
        RECT 202.800 456.300 203.600 456.400 ;
        RECT 204.500 456.300 205.100 467.600 ;
        RECT 206.000 463.600 206.800 464.400 ;
        RECT 207.600 463.600 208.400 464.400 ;
        RECT 202.800 455.700 205.100 456.300 ;
        RECT 202.800 455.600 203.600 455.700 ;
        RECT 198.100 452.400 198.700 455.600 ;
        RECT 202.900 452.400 203.500 455.600 ;
        RECT 198.000 451.600 198.800 452.400 ;
        RECT 202.800 451.600 203.600 452.400 ;
        RECT 196.400 449.600 197.200 450.400 ;
        RECT 199.600 447.600 200.400 448.400 ;
        RECT 201.200 443.600 202.000 444.400 ;
        RECT 194.800 433.600 195.600 434.400 ;
        RECT 194.900 430.400 195.500 433.600 ;
        RECT 194.800 429.600 195.600 430.400 ;
        RECT 193.200 427.600 194.000 428.400 ;
        RECT 193.300 420.400 193.900 427.600 ;
        RECT 198.000 424.200 198.800 435.800 ;
        RECT 201.300 434.400 201.900 443.600 ;
        RECT 201.200 433.600 202.000 434.400 ;
        RECT 201.200 426.200 202.000 431.800 ;
        RECT 204.400 430.300 205.200 430.400 ;
        RECT 206.100 430.300 206.700 463.600 ;
        RECT 207.700 458.400 208.300 463.600 ;
        RECT 207.600 457.600 208.400 458.400 ;
        RECT 209.300 454.400 209.900 467.600 ;
        RECT 209.200 453.600 210.000 454.400 ;
        RECT 210.800 453.600 211.600 454.400 ;
        RECT 209.300 448.400 209.900 453.600 ;
        RECT 210.900 450.400 211.500 453.600 ;
        RECT 210.800 449.600 211.600 450.400 ;
        RECT 209.200 447.600 210.000 448.400 ;
        RECT 212.500 434.400 213.100 467.600 ;
        RECT 214.100 464.400 214.700 469.600 ;
        RECT 222.100 468.400 222.700 469.600 ;
        RECT 223.700 468.400 224.300 471.600 ;
        RECT 222.000 467.600 222.800 468.400 ;
        RECT 223.600 467.600 224.400 468.400 ;
        RECT 214.000 463.600 214.800 464.400 ;
        RECT 225.300 458.400 225.900 483.600 ;
        RECT 230.100 478.400 230.700 493.600 ;
        RECT 231.600 486.200 232.400 497.800 ;
        RECT 233.200 484.200 234.000 497.800 ;
        RECT 234.800 484.200 235.600 497.800 ;
        RECT 230.000 477.600 230.800 478.400 ;
        RECT 236.500 474.400 237.100 503.600 ;
        RECT 238.000 491.600 238.800 492.400 ;
        RECT 236.400 473.600 237.200 474.400 ;
        RECT 226.800 471.800 227.600 472.600 ;
        RECT 233.400 471.800 234.200 472.600 ;
        RECT 238.100 472.400 238.700 491.600 ;
        RECT 226.800 468.400 227.400 471.800 ;
        RECT 230.800 468.400 231.600 468.600 ;
        RECT 226.800 467.800 231.600 468.400 ;
        RECT 226.800 467.000 227.400 467.800 ;
        RECT 228.200 467.000 229.000 467.200 ;
        RECT 231.600 467.000 232.400 467.200 ;
        RECT 233.600 467.000 234.200 471.800 ;
        RECT 238.000 471.600 238.800 472.400 ;
        RECT 241.300 470.400 241.900 505.600 ;
        RECT 244.500 498.400 245.100 511.600 ;
        RECT 246.000 507.600 246.800 508.400 ;
        RECT 247.600 507.600 248.400 508.400 ;
        RECT 246.100 506.400 246.700 507.600 ;
        RECT 252.500 506.400 253.100 531.600 ;
        RECT 254.000 509.600 254.800 510.400 ;
        RECT 246.000 505.600 246.800 506.400 ;
        RECT 247.600 505.600 248.400 506.400 ;
        RECT 252.400 505.600 253.200 506.400 ;
        RECT 244.400 497.600 245.200 498.400 ;
        RECT 244.400 491.600 245.200 492.400 ;
        RECT 239.600 469.600 240.400 470.400 ;
        RECT 241.200 469.600 242.000 470.400 ;
        RECT 234.800 467.600 235.600 468.400 ;
        RECT 226.800 466.200 227.600 467.000 ;
        RECT 228.200 466.400 232.400 467.000 ;
        RECT 228.400 465.600 229.200 466.400 ;
        RECT 233.400 466.200 234.200 467.000 ;
        RECT 230.000 463.600 230.800 464.400 ;
        RECT 236.400 463.600 237.200 464.400 ;
        RECT 225.200 457.600 226.000 458.400 ;
        RECT 222.000 455.600 222.800 456.400 ;
        RECT 222.100 454.400 222.700 455.600 ;
        RECT 222.000 453.600 222.800 454.400 ;
        RECT 228.400 453.600 229.200 454.400 ;
        RECT 230.100 452.400 230.700 463.600 ;
        RECT 236.500 454.400 237.100 463.600 ;
        RECT 239.700 454.400 240.300 469.600 ;
        RECT 241.200 467.600 242.000 468.400 ;
        RECT 242.800 467.600 243.600 468.400 ;
        RECT 241.300 466.400 241.900 467.600 ;
        RECT 241.200 465.600 242.000 466.400 ;
        RECT 236.400 453.600 237.200 454.400 ;
        RECT 239.600 453.600 240.400 454.400 ;
        RECT 230.000 451.600 230.800 452.400 ;
        RECT 225.200 449.600 226.000 450.400 ;
        RECT 214.000 437.600 214.800 438.400 ;
        RECT 207.600 433.600 208.400 434.400 ;
        RECT 212.400 433.600 213.200 434.400 ;
        RECT 207.700 432.400 208.300 433.600 ;
        RECT 214.100 432.400 214.700 437.600 ;
        RECT 225.300 436.400 225.900 449.600 ;
        RECT 225.200 435.600 226.000 436.400 ;
        RECT 220.400 433.600 221.200 434.400 ;
        RECT 220.500 432.400 221.100 433.600 ;
        RECT 230.100 432.400 230.700 451.600 ;
        RECT 233.200 443.600 234.000 444.400 ;
        RECT 238.000 443.600 238.800 444.400 ;
        RECT 207.600 431.600 208.400 432.400 ;
        RECT 214.000 431.600 214.800 432.400 ;
        RECT 215.600 431.600 216.400 432.400 ;
        RECT 218.800 431.600 219.600 432.400 ;
        RECT 220.400 431.600 221.200 432.400 ;
        RECT 230.000 431.600 230.800 432.400 ;
        RECT 218.900 430.400 219.500 431.600 ;
        RECT 204.400 429.700 206.700 430.300 ;
        RECT 204.400 429.600 205.200 429.700 ;
        RECT 210.800 429.600 211.600 430.400 ;
        RECT 218.800 429.600 219.600 430.400 ;
        RECT 223.600 429.600 224.400 430.400 ;
        RECT 226.800 429.600 227.600 430.400 ;
        RECT 230.000 429.600 230.800 430.400 ;
        RECT 202.800 427.600 203.600 428.400 ;
        RECT 204.500 422.400 205.100 429.600 ;
        RECT 218.800 427.600 219.600 428.400 ;
        RECT 225.200 425.600 226.000 426.400 ;
        RECT 214.000 423.600 214.800 424.400 ;
        RECT 215.600 423.600 216.400 424.400 ;
        RECT 217.200 423.600 218.000 424.400 ;
        RECT 204.400 421.600 205.200 422.400 ;
        RECT 214.100 420.400 214.700 423.600 ;
        RECT 193.200 419.600 194.000 420.400 ;
        RECT 198.000 419.600 198.800 420.400 ;
        RECT 214.000 419.600 214.800 420.400 ;
        RECT 172.400 417.600 173.200 418.400 ;
        RECT 174.000 415.600 174.800 416.400 ;
        RECT 174.100 412.400 174.700 415.600 ;
        RECT 175.600 413.600 176.400 414.400 ;
        RECT 174.000 411.600 174.800 412.400 ;
        RECT 180.400 411.600 181.200 412.400 ;
        RECT 180.500 410.400 181.100 411.600 ;
        RECT 180.400 409.600 181.200 410.400 ;
        RECT 170.800 407.600 171.600 408.400 ;
        RECT 162.800 405.600 163.600 406.400 ;
        RECT 177.200 403.600 178.000 404.400 ;
        RECT 190.000 404.200 190.800 417.800 ;
        RECT 191.600 404.200 192.400 417.800 ;
        RECT 193.200 406.200 194.000 417.800 ;
        RECT 194.800 413.600 195.600 414.400 ;
        RECT 194.800 411.600 195.600 412.400 ;
        RECT 177.300 400.400 177.900 403.600 ;
        RECT 177.200 399.600 178.000 400.400 ;
        RECT 186.800 399.600 187.600 400.400 ;
        RECT 158.000 397.600 158.800 398.400 ;
        RECT 161.200 397.600 162.000 398.400 ;
        RECT 167.600 397.600 168.400 398.400 ;
        RECT 156.400 389.600 157.200 390.400 ;
        RECT 156.500 388.400 157.100 389.600 ;
        RECT 156.400 387.600 157.200 388.400 ;
        RECT 151.600 385.600 152.400 386.400 ;
        RECT 166.000 385.600 166.800 386.400 ;
        RECT 148.400 377.600 149.200 378.400 ;
        RECT 148.500 370.400 149.100 377.600 ;
        RECT 148.400 369.600 149.200 370.400 ;
        RECT 151.700 364.400 152.300 385.600 ;
        RECT 161.200 383.600 162.000 384.400 ;
        RECT 153.200 371.600 154.000 372.400 ;
        RECT 154.800 370.200 155.600 375.800 ;
        RECT 156.400 373.600 157.200 374.400 ;
        RECT 151.600 363.600 152.400 364.400 ;
        RECT 156.500 358.400 157.100 373.600 ;
        RECT 158.000 366.200 158.800 377.800 ;
        RECT 161.300 374.400 161.900 383.600 ;
        RECT 166.100 374.400 166.700 385.600 ;
        RECT 172.400 383.600 173.200 384.400 ;
        RECT 177.200 384.200 178.000 397.800 ;
        RECT 178.800 384.200 179.600 397.800 ;
        RECT 180.400 384.200 181.200 397.800 ;
        RECT 182.000 384.200 182.800 395.800 ;
        RECT 183.600 385.600 184.400 386.400 ;
        RECT 185.200 384.200 186.000 395.800 ;
        RECT 186.900 388.400 187.500 399.600 ;
        RECT 186.800 387.600 187.600 388.400 ;
        RECT 188.400 384.200 189.200 395.800 ;
        RECT 190.000 384.200 190.800 397.800 ;
        RECT 191.600 384.200 192.400 397.800 ;
        RECT 194.900 390.400 195.500 411.600 ;
        RECT 196.400 406.200 197.200 417.800 ;
        RECT 198.100 416.400 198.700 419.600 ;
        RECT 198.000 415.600 198.800 416.400 ;
        RECT 199.600 406.200 200.400 417.800 ;
        RECT 201.200 404.200 202.000 417.800 ;
        RECT 202.800 404.200 203.600 417.800 ;
        RECT 204.400 404.200 205.200 417.800 ;
        RECT 215.700 414.400 216.300 423.600 ;
        RECT 217.300 416.400 217.900 423.600 ;
        RECT 225.300 416.400 225.900 425.600 ;
        RECT 226.900 418.400 227.500 429.600 ;
        RECT 230.100 424.400 230.700 429.600 ;
        RECT 238.100 428.400 238.700 443.600 ;
        RECT 242.900 438.400 243.500 467.600 ;
        RECT 244.500 464.400 245.100 491.600 ;
        RECT 246.100 488.400 246.700 505.600 ;
        RECT 247.700 502.400 248.300 505.600 ;
        RECT 247.600 501.600 248.400 502.400 ;
        RECT 247.700 498.400 248.300 501.600 ;
        RECT 247.600 497.600 248.400 498.400 ;
        RECT 250.800 495.600 251.600 496.400 ;
        RECT 250.900 494.400 251.500 495.600 ;
        RECT 250.800 493.600 251.600 494.400 ;
        RECT 246.000 487.600 246.800 488.400 ;
        RECT 246.100 466.400 246.700 487.600 ;
        RECT 252.400 483.600 253.200 484.400 ;
        RECT 250.800 471.600 251.600 472.400 ;
        RECT 247.600 469.600 248.400 470.400 ;
        RECT 246.000 465.600 246.800 466.400 ;
        RECT 247.700 464.400 248.300 469.600 ;
        RECT 244.400 463.600 245.200 464.400 ;
        RECT 247.600 463.600 248.400 464.400 ;
        RECT 250.900 460.400 251.500 471.600 ;
        RECT 252.500 466.400 253.100 483.600 ;
        RECT 254.100 470.400 254.700 509.600 ;
        RECT 257.200 504.200 258.000 517.800 ;
        RECT 258.800 504.200 259.600 517.800 ;
        RECT 260.400 504.200 261.200 515.800 ;
        RECT 262.100 510.400 262.700 531.700 ;
        RECT 263.600 531.600 264.400 531.700 ;
        RECT 262.000 509.600 262.800 510.400 ;
        RECT 262.000 507.600 262.800 508.400 ;
        RECT 263.600 504.200 264.400 515.800 ;
        RECT 265.300 506.400 265.900 535.600 ;
        RECT 268.400 524.200 269.200 537.800 ;
        RECT 270.000 524.200 270.800 537.800 ;
        RECT 271.600 526.200 272.400 537.800 ;
        RECT 273.300 536.400 273.900 545.600 ;
        RECT 274.800 544.200 275.600 555.800 ;
        RECT 276.400 544.200 277.200 557.800 ;
        RECT 278.000 544.200 278.800 557.800 ;
        RECT 279.600 544.200 280.400 557.800 ;
        RECT 300.400 545.600 301.200 546.400 ;
        RECT 289.200 543.600 290.000 544.400 ;
        RECT 273.200 535.600 274.000 536.400 ;
        RECT 273.200 533.600 274.000 534.400 ;
        RECT 273.300 522.400 273.900 533.600 ;
        RECT 274.800 526.200 275.600 537.800 ;
        RECT 276.400 535.600 277.200 536.400 ;
        RECT 278.000 526.200 278.800 537.800 ;
        RECT 279.600 524.200 280.400 537.800 ;
        RECT 281.200 524.200 282.000 537.800 ;
        RECT 282.800 524.200 283.600 537.800 ;
        RECT 289.300 536.400 289.900 543.600 ;
        RECT 292.400 541.600 293.200 542.400 ;
        RECT 298.800 541.600 299.600 542.400 ;
        RECT 292.500 538.400 293.100 541.600 ;
        RECT 292.400 537.600 293.200 538.400 ;
        RECT 298.900 536.400 299.500 541.600 ;
        RECT 289.200 535.600 290.000 536.400 ;
        RECT 295.600 535.600 296.400 536.400 ;
        RECT 298.800 535.600 299.600 536.400 ;
        RECT 298.900 534.400 299.500 535.600 ;
        RECT 298.800 533.600 299.600 534.400 ;
        RECT 300.500 522.400 301.100 545.600 ;
        RECT 313.200 544.200 314.000 557.800 ;
        RECT 314.800 544.200 315.600 557.800 ;
        RECT 316.400 544.200 317.200 557.800 ;
        RECT 318.000 544.200 318.800 555.800 ;
        RECT 319.600 545.600 320.400 546.400 ;
        RECT 302.000 537.600 302.800 538.400 ;
        RECT 302.100 534.400 302.700 537.600 ;
        RECT 319.700 536.400 320.300 545.600 ;
        RECT 321.200 544.200 322.000 555.800 ;
        RECT 322.800 547.600 323.600 548.400 ;
        RECT 324.400 544.200 325.200 555.800 ;
        RECT 326.000 544.200 326.800 557.800 ;
        RECT 327.600 544.200 328.400 557.800 ;
        RECT 346.800 551.600 347.600 552.400 ;
        RECT 361.200 551.600 362.000 552.400 ;
        RECT 364.400 551.600 365.200 552.400 ;
        RECT 332.400 549.600 333.200 550.400 ;
        RECT 342.000 549.600 342.800 550.400 ;
        RECT 345.200 549.600 346.000 550.400 ;
        RECT 342.100 540.400 342.700 549.600 ;
        RECT 343.600 547.600 344.400 548.400 ;
        RECT 342.000 539.600 342.800 540.400 ;
        RECT 310.000 535.600 310.800 536.400 ;
        RECT 319.600 535.600 320.400 536.400 ;
        RECT 310.100 534.400 310.700 535.600 ;
        RECT 302.000 533.600 302.800 534.400 ;
        RECT 310.000 533.600 310.800 534.400 ;
        RECT 313.200 529.600 314.000 530.400 ;
        RECT 318.000 529.600 318.800 530.400 ;
        RECT 273.200 521.600 274.000 522.400 ;
        RECT 281.200 521.600 282.000 522.400 ;
        RECT 300.400 521.600 301.200 522.400 ;
        RECT 281.300 518.400 281.900 521.600 ;
        RECT 265.200 505.600 266.000 506.400 ;
        RECT 265.300 494.400 265.900 505.600 ;
        RECT 266.800 504.200 267.600 515.800 ;
        RECT 268.400 504.200 269.200 517.800 ;
        RECT 270.000 504.200 270.800 517.800 ;
        RECT 271.600 504.200 272.400 517.800 ;
        RECT 281.200 517.600 282.000 518.400 ;
        RECT 279.600 509.600 280.400 510.400 ;
        RECT 287.600 509.600 288.400 510.400 ;
        RECT 263.600 493.600 264.400 494.400 ;
        RECT 265.200 493.600 266.000 494.400 ;
        RECT 278.000 493.600 278.800 494.400 ;
        RECT 279.700 490.400 280.300 509.600 ;
        RECT 281.200 503.600 282.000 504.400 ;
        RECT 281.300 498.400 281.900 503.600 ;
        RECT 281.200 497.600 282.000 498.400 ;
        RECT 281.200 493.600 282.000 494.400 ;
        RECT 284.400 493.600 285.200 494.400 ;
        RECT 286.000 493.600 286.800 494.400 ;
        RECT 282.800 491.600 283.600 492.400 ;
        RECT 279.600 489.600 280.400 490.400 ;
        RECT 257.200 471.600 258.000 472.400 ;
        RECT 254.000 469.600 254.800 470.400 ;
        RECT 252.400 465.600 253.200 466.400 ;
        RECT 246.000 459.600 246.800 460.400 ;
        RECT 250.800 459.600 251.600 460.400 ;
        RECT 252.500 460.300 253.100 465.600 ;
        RECT 262.000 464.200 262.800 477.800 ;
        RECT 263.600 464.200 264.400 477.800 ;
        RECT 265.200 464.200 266.000 475.800 ;
        RECT 266.800 467.600 267.600 468.400 ;
        RECT 266.900 462.300 267.500 467.600 ;
        RECT 268.400 464.200 269.200 475.800 ;
        RECT 270.000 465.600 270.800 466.400 ;
        RECT 271.600 464.200 272.400 475.800 ;
        RECT 273.200 464.200 274.000 477.800 ;
        RECT 274.800 464.200 275.600 477.800 ;
        RECT 276.400 464.200 277.200 477.800 ;
        RECT 278.000 463.600 278.800 464.400 ;
        RECT 265.300 461.700 267.500 462.300 ;
        RECT 252.500 459.700 254.700 460.300 ;
        RECT 246.100 452.400 246.700 459.600 ;
        RECT 246.000 451.600 246.800 452.400 ;
        RECT 246.000 447.600 246.800 448.400 ;
        RECT 242.800 437.600 243.600 438.400 ;
        RECT 242.900 432.400 243.500 437.600 ;
        RECT 241.200 431.600 242.000 432.400 ;
        RECT 242.800 431.600 243.600 432.400 ;
        RECT 231.600 427.600 232.400 428.400 ;
        RECT 233.200 427.600 234.000 428.400 ;
        RECT 238.000 427.600 238.800 428.400 ;
        RECT 231.700 426.400 232.300 427.600 ;
        RECT 231.600 425.600 232.400 426.400 ;
        RECT 233.300 424.400 233.900 427.600 ;
        RECT 230.000 423.600 230.800 424.400 ;
        RECT 233.200 423.600 234.000 424.400 ;
        RECT 234.800 423.600 235.600 424.400 ;
        RECT 226.800 417.600 227.600 418.400 ;
        RECT 217.200 415.600 218.000 416.400 ;
        RECT 225.200 415.600 226.000 416.400 ;
        RECT 234.900 414.400 235.500 423.600 ;
        RECT 238.100 416.400 238.700 427.600 ;
        RECT 238.000 415.600 238.800 416.400 ;
        RECT 238.100 414.400 238.700 415.600 ;
        RECT 215.600 413.600 216.400 414.400 ;
        RECT 230.000 413.600 230.800 414.400 ;
        RECT 234.800 413.600 235.600 414.400 ;
        RECT 238.000 413.600 238.800 414.400 ;
        RECT 239.600 413.600 240.400 414.400 ;
        RECT 230.100 412.400 230.700 413.600 ;
        RECT 223.600 411.600 224.400 412.400 ;
        RECT 230.000 411.600 230.800 412.400 ;
        RECT 234.800 411.600 235.600 412.400 ;
        RECT 223.700 410.400 224.300 411.600 ;
        RECT 223.600 409.600 224.400 410.400 ;
        RECT 236.400 410.300 237.200 410.400 ;
        RECT 238.100 410.300 238.700 413.600 ;
        RECT 239.700 412.400 240.300 413.600 ;
        RECT 239.600 412.300 240.400 412.400 ;
        RECT 241.300 412.300 241.900 431.600 ;
        RECT 246.100 430.400 246.700 447.600 ;
        RECT 247.600 444.200 248.400 457.800 ;
        RECT 249.200 444.200 250.000 457.800 ;
        RECT 250.800 444.200 251.600 457.800 ;
        RECT 252.400 446.200 253.200 457.800 ;
        RECT 254.100 456.400 254.700 459.700 ;
        RECT 254.000 455.600 254.800 456.400 ;
        RECT 255.600 446.200 256.400 457.800 ;
        RECT 257.200 453.600 258.000 454.400 ;
        RECT 257.300 452.400 257.900 453.600 ;
        RECT 257.200 451.600 258.000 452.400 ;
        RECT 258.800 446.200 259.600 457.800 ;
        RECT 260.400 444.200 261.200 457.800 ;
        RECT 262.000 444.200 262.800 457.800 ;
        RECT 265.300 448.400 265.900 461.700 ;
        RECT 274.800 455.600 275.600 456.400 ;
        RECT 276.400 455.600 277.200 456.400 ;
        RECT 274.900 454.400 275.500 455.600 ;
        RECT 276.500 454.400 277.100 455.600 ;
        RECT 274.800 453.600 275.600 454.400 ;
        RECT 276.400 453.600 277.200 454.400 ;
        RECT 278.100 452.400 278.700 463.600 ;
        RECT 281.200 455.600 282.000 456.400 ;
        RECT 282.900 454.400 283.500 491.600 ;
        RECT 284.500 488.400 285.100 493.600 ;
        RECT 284.400 487.600 285.200 488.400 ;
        RECT 284.400 485.600 285.200 486.400 ;
        RECT 282.800 453.600 283.600 454.400 ;
        RECT 273.200 451.600 274.000 452.400 ;
        RECT 278.000 451.600 278.800 452.400 ;
        RECT 265.200 447.600 266.000 448.400 ;
        RECT 271.600 443.600 272.400 444.400 ;
        RECT 249.200 441.600 250.000 442.400 ;
        RECT 242.800 429.600 243.600 430.400 ;
        RECT 246.000 429.600 246.800 430.400 ;
        RECT 246.100 418.400 246.700 429.600 ;
        RECT 247.600 423.600 248.400 424.400 ;
        RECT 246.000 417.600 246.800 418.400 ;
        RECT 247.700 416.400 248.300 423.600 ;
        RECT 247.600 415.600 248.400 416.400 ;
        RECT 247.600 413.600 248.400 414.400 ;
        RECT 239.600 411.700 241.900 412.300 ;
        RECT 239.600 411.600 240.400 411.700 ;
        RECT 236.400 409.700 238.700 410.300 ;
        RECT 236.400 409.600 237.200 409.700 ;
        RECT 242.800 409.600 243.600 410.400 ;
        RECT 218.800 407.600 219.600 408.400 ;
        RECT 233.200 407.600 234.000 408.400 ;
        RECT 222.000 403.600 222.800 404.400 ;
        RECT 202.800 401.600 203.600 402.400 ;
        RECT 202.900 398.400 203.500 401.600 ;
        RECT 222.100 400.400 222.700 403.600 ;
        RECT 222.000 399.600 222.800 400.400 ;
        RECT 202.800 397.600 203.600 398.400 ;
        RECT 204.400 397.600 205.200 398.400 ;
        RECT 204.500 392.400 205.100 397.600 ;
        RECT 209.200 393.600 210.000 394.400 ;
        RECT 209.300 392.400 209.900 393.600 ;
        RECT 204.400 391.600 205.200 392.400 ;
        RECT 209.200 391.600 210.000 392.400 ;
        RECT 212.400 391.600 213.200 392.400 ;
        RECT 194.800 389.600 195.600 390.400 ;
        RECT 196.400 390.300 197.200 390.400 ;
        RECT 198.000 390.300 198.800 390.400 ;
        RECT 196.400 389.700 198.800 390.300 ;
        RECT 196.400 389.600 197.200 389.700 ;
        RECT 198.000 389.600 198.800 389.700 ;
        RECT 172.500 378.400 173.100 383.600 ;
        RECT 161.200 373.600 162.000 374.400 ;
        RECT 166.000 373.600 166.800 374.400 ;
        RECT 159.600 371.600 160.400 372.600 ;
        RECT 153.200 357.600 154.000 358.400 ;
        RECT 156.400 357.600 157.200 358.400 ;
        RECT 161.300 354.400 161.900 373.600 ;
        RECT 167.600 366.200 168.400 377.800 ;
        RECT 172.400 377.600 173.200 378.400 ;
        RECT 172.500 376.400 173.100 377.600 ;
        RECT 172.400 375.600 173.200 376.400 ;
        RECT 182.000 364.200 182.800 377.800 ;
        RECT 183.600 364.200 184.400 377.800 ;
        RECT 185.200 366.200 186.000 377.800 ;
        RECT 186.800 373.600 187.600 374.400 ;
        RECT 188.400 366.200 189.200 377.800 ;
        RECT 190.000 375.600 190.800 376.400 ;
        RECT 191.600 366.200 192.400 377.800 ;
        RECT 193.200 364.200 194.000 377.800 ;
        RECT 194.800 364.200 195.600 377.800 ;
        RECT 196.400 364.200 197.200 377.800 ;
        RECT 198.100 372.400 198.700 389.600 ;
        RECT 207.600 387.600 208.400 388.400 ;
        RECT 207.700 386.400 208.300 387.600 ;
        RECT 201.200 385.600 202.000 386.400 ;
        RECT 207.600 385.600 208.400 386.400 ;
        RECT 201.300 384.400 201.900 385.600 ;
        RECT 201.200 383.600 202.000 384.400 ;
        RECT 204.400 383.600 205.200 384.400 ;
        RECT 204.500 374.400 205.100 383.600 ;
        RECT 204.400 373.600 205.200 374.400 ;
        RECT 198.000 371.600 198.800 372.400 ;
        RECT 198.100 362.400 198.700 371.600 ;
        RECT 209.300 370.400 209.900 391.600 ;
        RECT 212.500 388.400 213.100 391.600 ;
        RECT 217.200 389.600 218.000 390.400 ;
        RECT 210.800 387.600 211.600 388.400 ;
        RECT 212.400 387.600 213.200 388.400 ;
        RECT 214.000 385.600 214.800 386.400 ;
        RECT 214.100 378.400 214.700 385.600 ;
        RECT 222.000 384.200 222.800 397.800 ;
        RECT 223.600 384.200 224.400 397.800 ;
        RECT 225.200 384.200 226.000 395.800 ;
        RECT 226.800 387.600 227.600 388.400 ;
        RECT 228.400 384.200 229.200 395.800 ;
        RECT 230.000 385.600 230.800 386.400 ;
        RECT 228.400 381.600 229.200 382.400 ;
        RECT 214.000 377.600 214.800 378.400 ;
        RECT 218.800 377.600 219.600 378.400 ;
        RECT 226.800 377.600 227.600 378.400 ;
        RECT 218.900 374.400 219.500 377.600 ;
        RECT 226.900 374.400 227.500 377.600 ;
        RECT 212.400 373.600 213.200 374.400 ;
        RECT 218.800 373.600 219.600 374.400 ;
        RECT 220.400 373.600 221.200 374.400 ;
        RECT 226.800 373.600 227.600 374.400 ;
        RECT 228.500 372.400 229.100 381.600 ;
        RECT 230.100 376.400 230.700 385.600 ;
        RECT 231.600 384.200 232.400 395.800 ;
        RECT 233.200 384.200 234.000 397.800 ;
        RECT 234.800 384.200 235.600 397.800 ;
        RECT 236.400 384.200 237.200 397.800 ;
        RECT 249.300 394.400 249.900 441.600 ;
        RECT 271.700 434.400 272.300 443.600 ;
        RECT 273.300 438.400 273.900 451.600 ;
        RECT 278.100 438.400 278.700 451.600 ;
        RECT 281.200 443.600 282.000 444.400 ;
        RECT 273.200 437.600 274.000 438.400 ;
        RECT 278.000 437.600 278.800 438.400 ;
        RECT 278.000 435.600 278.800 436.400 ;
        RECT 268.400 433.600 269.200 434.400 ;
        RECT 271.600 433.600 272.400 434.400 ;
        RECT 252.400 431.600 253.200 432.400 ;
        RECT 255.600 431.600 256.400 432.400 ;
        RECT 252.500 424.400 253.100 431.600 ;
        RECT 255.700 430.400 256.300 431.600 ;
        RECT 268.500 430.400 269.100 433.600 ;
        RECT 278.100 432.400 278.700 435.600 ;
        RECT 276.400 431.600 277.200 432.400 ;
        RECT 278.000 431.600 278.800 432.400 ;
        RECT 254.000 429.600 254.800 430.400 ;
        RECT 255.600 429.600 256.400 430.400 ;
        RECT 258.800 429.600 259.600 430.400 ;
        RECT 260.400 429.600 261.200 430.400 ;
        RECT 265.200 429.600 266.000 430.400 ;
        RECT 266.800 429.600 267.600 430.400 ;
        RECT 268.400 429.600 269.200 430.400 ;
        RECT 270.000 429.600 270.800 430.400 ;
        RECT 274.800 429.600 275.600 430.400 ;
        RECT 254.100 424.400 254.700 429.600 ;
        RECT 257.200 427.600 258.000 428.400 ;
        RECT 258.900 426.400 259.500 429.600 ;
        RECT 265.300 428.400 265.900 429.600 ;
        RECT 266.900 428.400 267.500 429.600 ;
        RECT 265.200 427.600 266.000 428.400 ;
        RECT 266.800 427.600 267.600 428.400 ;
        RECT 258.800 426.300 259.600 426.400 ;
        RECT 258.800 425.700 261.100 426.300 ;
        RECT 258.800 425.600 259.600 425.700 ;
        RECT 252.400 423.600 253.200 424.400 ;
        RECT 254.000 423.600 254.800 424.400 ;
        RECT 254.100 418.400 254.700 423.600 ;
        RECT 254.000 417.600 254.800 418.400 ;
        RECT 251.000 415.600 251.800 415.800 ;
        RECT 251.000 415.000 256.600 415.600 ;
        RECT 257.200 415.000 258.000 415.800 ;
        RECT 251.000 410.200 251.600 415.000 ;
        RECT 252.400 414.800 253.200 415.000 ;
        RECT 255.800 414.800 256.600 415.000 ;
        RECT 257.400 414.200 258.000 415.000 ;
        RECT 252.400 413.600 258.000 414.200 ;
        RECT 258.800 413.600 259.600 414.400 ;
        RECT 252.400 412.200 253.000 413.600 ;
        RECT 252.200 411.400 253.000 412.200 ;
        RECT 257.400 410.200 258.000 413.600 ;
        RECT 258.900 412.400 259.500 413.600 ;
        RECT 258.800 411.600 259.600 412.400 ;
        RECT 260.500 410.400 261.100 425.700 ;
        RECT 270.100 424.400 270.700 429.600 ;
        RECT 273.200 427.600 274.000 428.400 ;
        RECT 270.000 423.600 270.800 424.400 ;
        RECT 273.300 418.400 273.900 427.600 ;
        RECT 273.200 417.600 274.000 418.400 ;
        RECT 262.000 415.600 262.800 416.400 ;
        RECT 266.800 415.600 267.600 416.400 ;
        RECT 268.600 415.600 269.400 415.800 ;
        RECT 262.100 414.400 262.700 415.600 ;
        RECT 266.900 414.400 267.500 415.600 ;
        RECT 268.600 415.000 274.200 415.600 ;
        RECT 274.800 415.000 275.600 415.800 ;
        RECT 262.000 413.600 262.800 414.400 ;
        RECT 263.600 413.600 264.400 414.400 ;
        RECT 265.200 413.600 266.000 414.400 ;
        RECT 266.800 413.600 267.600 414.400 ;
        RECT 263.700 412.400 264.300 413.600 ;
        RECT 265.300 412.400 265.900 413.600 ;
        RECT 263.600 411.600 264.400 412.400 ;
        RECT 265.200 411.600 266.000 412.400 ;
        RECT 251.000 409.400 251.800 410.200 ;
        RECT 257.200 409.400 258.000 410.200 ;
        RECT 260.400 409.600 261.200 410.400 ;
        RECT 263.700 404.400 264.300 411.600 ;
        RECT 268.600 410.200 269.200 415.000 ;
        RECT 270.000 414.800 270.800 415.000 ;
        RECT 273.400 414.800 274.200 415.000 ;
        RECT 275.000 414.200 275.600 415.000 ;
        RECT 276.500 414.400 277.100 431.600 ;
        RECT 281.300 430.400 281.900 443.600 ;
        RECT 284.500 438.400 285.100 485.600 ;
        RECT 287.700 472.400 288.300 509.600 ;
        RECT 289.200 507.600 290.000 508.400 ;
        RECT 289.300 498.400 289.900 507.600 ;
        RECT 292.400 504.200 293.200 517.800 ;
        RECT 294.000 504.200 294.800 517.800 ;
        RECT 295.600 504.200 296.400 515.800 ;
        RECT 297.200 507.600 298.000 508.400 ;
        RECT 298.800 504.200 299.600 515.800 ;
        RECT 300.400 505.600 301.200 506.400 ;
        RECT 302.000 504.200 302.800 515.800 ;
        RECT 303.600 504.200 304.400 517.800 ;
        RECT 305.200 504.200 306.000 517.800 ;
        RECT 306.800 504.200 307.600 517.800 ;
        RECT 313.300 510.400 313.900 529.600 ;
        RECT 316.400 524.300 317.200 524.400 ;
        RECT 318.100 524.300 318.700 529.600 ;
        RECT 316.400 523.700 318.700 524.300 ;
        RECT 316.400 523.600 317.200 523.700 ;
        RECT 318.100 514.400 318.700 523.700 ;
        RECT 318.000 513.600 318.800 514.400 ;
        RECT 319.700 512.400 320.300 535.600 ;
        RECT 326.000 524.200 326.800 537.800 ;
        RECT 327.600 524.200 328.400 537.800 ;
        RECT 329.200 524.200 330.000 537.800 ;
        RECT 330.800 526.200 331.600 537.800 ;
        RECT 332.400 535.600 333.200 536.400 ;
        RECT 334.000 526.200 334.800 537.800 ;
        RECT 335.600 535.600 336.400 536.400 ;
        RECT 335.700 534.400 336.300 535.600 ;
        RECT 335.600 533.600 336.400 534.400 ;
        RECT 337.200 526.200 338.000 537.800 ;
        RECT 338.800 524.200 339.600 537.800 ;
        RECT 340.400 524.200 341.200 537.800 ;
        RECT 345.300 532.400 345.900 549.600 ;
        RECT 345.200 531.600 346.000 532.400 ;
        RECT 346.900 522.400 347.500 551.600 ;
        RECT 350.000 549.600 350.800 550.400 ;
        RECT 358.000 549.600 358.800 550.400 ;
        RECT 362.800 549.600 363.600 550.400 ;
        RECT 364.400 549.600 365.200 550.400 ;
        RECT 350.100 548.400 350.700 549.600 ;
        RECT 350.000 547.600 350.800 548.400 ;
        RECT 351.600 547.600 352.400 548.400 ;
        RECT 351.700 546.400 352.300 547.600 ;
        RECT 351.600 545.600 352.400 546.400 ;
        RECT 358.100 540.400 358.700 549.600 ;
        RECT 364.500 548.400 365.100 549.600 ;
        RECT 362.800 547.600 363.600 548.400 ;
        RECT 364.400 547.600 365.200 548.400 ;
        RECT 362.900 546.400 363.500 547.600 ;
        RECT 362.800 545.600 363.600 546.400 ;
        RECT 353.200 539.600 354.000 540.400 ;
        RECT 358.000 539.600 358.800 540.400 ;
        RECT 350.000 535.600 350.800 536.400 ;
        RECT 350.000 533.600 350.800 534.400 ;
        RECT 350.100 530.400 350.700 533.600 ;
        RECT 353.300 532.400 353.900 539.600 ;
        RECT 358.000 533.600 358.800 534.400 ;
        RECT 364.500 532.400 365.100 547.600 ;
        RECT 366.000 545.600 366.800 546.400 ;
        RECT 366.100 534.400 366.700 545.600 ;
        RECT 370.800 543.600 371.600 544.400 ;
        RECT 380.400 544.200 381.200 557.800 ;
        RECT 382.000 544.200 382.800 557.800 ;
        RECT 383.600 544.200 384.400 557.800 ;
        RECT 385.200 544.200 386.000 555.800 ;
        RECT 386.800 545.600 387.600 546.400 ;
        RECT 370.900 538.400 371.500 543.600 ;
        RECT 377.200 539.600 378.000 540.400 ;
        RECT 370.800 537.600 371.600 538.400 ;
        RECT 367.600 535.600 368.400 536.400 ;
        RECT 366.000 533.600 366.800 534.400 ;
        RECT 353.200 531.600 354.000 532.400 ;
        RECT 364.400 531.600 365.200 532.400 ;
        RECT 350.000 529.600 350.800 530.400 ;
        RECT 359.600 529.600 360.400 530.400 ;
        RECT 356.400 527.600 357.200 528.400 ;
        RECT 329.200 521.600 330.000 522.400 ;
        RECT 346.800 521.600 347.600 522.400 ;
        RECT 329.300 514.400 329.900 521.600 ;
        RECT 329.200 513.600 330.000 514.400 ;
        RECT 319.600 511.600 320.400 512.400 ;
        RECT 313.200 509.600 314.000 510.400 ;
        RECT 316.400 509.600 317.400 510.400 ;
        RECT 319.700 506.400 320.300 511.600 ;
        RECT 329.200 509.600 330.000 510.400 ;
        RECT 327.600 507.600 328.400 508.400 ;
        RECT 319.600 505.600 320.400 506.400 ;
        RECT 319.600 503.600 320.400 504.400 ;
        RECT 314.800 501.600 315.600 502.400 ;
        RECT 289.200 497.600 290.000 498.400 ;
        RECT 294.000 497.600 294.800 498.400 ;
        RECT 302.000 497.600 302.800 498.400 ;
        RECT 290.800 493.600 291.600 494.400 ;
        RECT 292.400 491.600 293.200 492.400 ;
        RECT 289.200 489.600 290.000 490.400 ;
        RECT 289.300 474.400 289.900 489.600 ;
        RECT 292.500 486.400 293.100 491.600 ;
        RECT 292.400 485.600 293.200 486.400 ;
        RECT 289.200 473.600 290.000 474.400 ;
        RECT 292.400 473.600 293.200 474.400 ;
        RECT 292.500 472.400 293.100 473.600 ;
        RECT 287.600 471.600 288.400 472.400 ;
        RECT 292.400 471.600 293.200 472.400 ;
        RECT 294.100 470.400 294.700 497.600 ;
        RECT 295.600 495.600 296.400 496.400 ;
        RECT 297.200 493.600 298.000 494.400 ;
        RECT 298.800 491.600 299.600 492.400 ;
        RECT 302.100 490.400 302.700 497.600 ;
        RECT 314.900 496.400 315.500 501.600 ;
        RECT 319.700 498.400 320.300 503.600 ;
        RECT 329.300 498.400 329.900 509.600 ;
        RECT 332.400 507.600 333.200 508.400 ;
        RECT 330.800 503.600 331.600 504.400 ;
        RECT 332.500 504.300 333.100 507.600 ;
        RECT 334.000 506.200 334.800 511.800 ;
        RECT 335.600 511.600 336.400 512.400 ;
        RECT 335.700 508.400 336.300 511.600 ;
        RECT 335.600 507.600 336.400 508.400 ;
        RECT 335.600 505.600 336.400 506.400 ;
        RECT 332.500 503.700 334.700 504.300 ;
        RECT 330.900 498.400 331.500 503.600 ;
        RECT 319.600 497.600 320.400 498.400 ;
        RECT 329.200 497.600 330.000 498.400 ;
        RECT 330.800 497.600 331.600 498.400 ;
        RECT 314.800 495.600 315.600 496.400 ;
        RECT 319.600 495.600 320.400 496.400 ;
        RECT 324.400 495.600 325.200 496.400 ;
        RECT 330.800 495.600 331.600 496.400 ;
        RECT 314.900 492.400 315.500 495.600 ;
        RECT 324.500 494.400 325.100 495.600 ;
        RECT 324.400 493.600 325.200 494.400 ;
        RECT 310.000 491.600 310.800 492.400 ;
        RECT 311.600 491.600 312.400 492.400 ;
        RECT 314.800 491.600 315.600 492.400 ;
        RECT 318.000 491.600 318.800 492.400 ;
        RECT 322.800 491.600 323.600 492.400 ;
        RECT 326.000 491.600 326.800 492.400 ;
        RECT 310.100 490.400 310.700 491.600 ;
        RECT 295.600 489.600 296.400 490.400 ;
        RECT 302.000 489.600 302.800 490.400 ;
        RECT 310.000 489.600 310.800 490.400 ;
        RECT 300.400 487.600 301.200 488.400 ;
        RECT 298.800 483.600 299.600 484.400 ;
        RECT 298.900 482.400 299.500 483.600 ;
        RECT 298.800 481.600 299.600 482.400 ;
        RECT 300.500 478.400 301.100 487.600 ;
        RECT 300.400 477.600 301.200 478.400 ;
        RECT 294.000 469.600 294.800 470.400 ;
        RECT 303.600 469.600 304.400 470.400 ;
        RECT 289.200 467.600 290.000 468.400 ;
        RECT 286.000 463.600 286.800 464.400 ;
        RECT 289.300 458.400 289.900 467.600 ;
        RECT 297.200 465.600 298.000 466.400 ;
        RECT 292.400 463.600 293.200 464.400 ;
        RECT 295.600 463.600 296.400 464.400 ;
        RECT 289.200 457.600 290.000 458.400 ;
        RECT 286.000 455.600 286.800 456.400 ;
        RECT 286.100 454.400 286.700 455.600 ;
        RECT 292.500 454.400 293.100 463.600 ;
        RECT 295.700 456.400 296.300 463.600 ;
        RECT 295.600 455.600 296.400 456.400 ;
        RECT 286.000 453.600 286.800 454.400 ;
        RECT 292.400 453.600 293.200 454.400 ;
        RECT 286.100 452.400 286.700 453.600 ;
        RECT 286.000 451.600 286.800 452.400 ;
        RECT 284.400 437.600 285.200 438.400 ;
        RECT 281.200 429.600 282.000 430.400 ;
        RECT 284.400 429.600 285.200 430.400 ;
        RECT 281.200 427.600 282.000 428.400 ;
        RECT 279.600 423.600 280.400 424.400 ;
        RECT 279.700 418.400 280.300 423.600 ;
        RECT 279.600 417.600 280.400 418.400 ;
        RECT 278.000 415.600 278.800 416.400 ;
        RECT 278.100 414.400 278.700 415.600 ;
        RECT 281.300 414.400 281.900 427.600 ;
        RECT 282.800 425.600 283.600 426.400 ;
        RECT 282.900 422.400 283.500 425.600 ;
        RECT 282.800 421.600 283.600 422.400 ;
        RECT 282.800 417.600 283.600 418.400 ;
        RECT 270.000 413.600 275.600 414.200 ;
        RECT 276.400 413.600 277.200 414.400 ;
        RECT 278.000 413.600 278.800 414.400 ;
        RECT 281.200 413.600 282.000 414.400 ;
        RECT 270.000 412.200 270.600 413.600 ;
        RECT 269.800 411.400 270.600 412.200 ;
        RECT 275.000 410.200 275.600 413.600 ;
        RECT 278.100 412.400 278.700 413.600 ;
        RECT 278.000 411.600 278.800 412.400 ;
        RECT 279.600 411.600 280.400 412.400 ;
        RECT 282.900 410.400 283.500 417.600 ;
        RECT 284.500 416.400 285.100 429.600 ;
        RECT 284.400 415.600 285.200 416.400 ;
        RECT 284.500 414.400 285.100 415.600 ;
        RECT 284.400 413.600 285.200 414.400 ;
        RECT 286.100 412.400 286.700 451.600 ;
        RECT 297.300 446.400 297.900 465.600 ;
        RECT 303.700 464.400 304.300 469.600 ;
        RECT 310.000 466.200 310.800 471.800 ;
        RECT 303.600 463.600 304.400 464.400 ;
        RECT 313.200 464.200 314.000 475.800 ;
        RECT 316.400 475.600 317.200 476.400 ;
        RECT 316.500 470.400 317.100 475.600 ;
        RECT 316.400 469.600 317.200 470.400 ;
        RECT 314.800 465.600 315.600 466.400 ;
        RECT 314.900 462.300 315.500 465.600 ;
        RECT 313.300 461.700 315.500 462.300 ;
        RECT 305.200 451.600 306.000 452.400 ;
        RECT 297.200 445.600 298.000 446.400 ;
        RECT 305.300 444.400 305.900 451.600 ;
        RECT 295.600 443.600 296.400 444.400 ;
        RECT 297.200 443.600 298.000 444.400 ;
        RECT 305.200 443.600 306.000 444.400 ;
        RECT 306.800 444.200 307.600 457.800 ;
        RECT 308.400 444.200 309.200 457.800 ;
        RECT 310.000 444.200 310.800 457.800 ;
        RECT 311.600 446.200 312.400 457.800 ;
        RECT 313.300 456.400 313.900 461.700 ;
        RECT 318.100 460.400 318.700 491.600 ;
        RECT 322.900 486.400 323.500 491.600 ;
        RECT 329.200 489.600 330.000 490.400 ;
        RECT 329.300 488.400 329.900 489.600 ;
        RECT 329.200 487.600 330.000 488.400 ;
        RECT 322.800 485.600 323.600 486.400 ;
        RECT 330.900 484.400 331.500 495.600 ;
        RECT 334.100 494.400 334.700 503.700 ;
        RECT 334.000 493.600 334.800 494.400 ;
        RECT 334.100 492.400 334.700 493.600 ;
        RECT 335.700 492.400 336.300 505.600 ;
        RECT 337.200 504.200 338.000 515.800 ;
        RECT 338.800 509.400 339.600 510.400 ;
        RECT 346.800 504.200 347.600 515.800 ;
        RECT 356.500 514.400 357.100 527.600 ;
        RECT 366.100 522.400 366.700 533.600 ;
        RECT 366.000 521.600 366.800 522.400 ;
        RECT 356.400 513.600 357.200 514.400 ;
        RECT 353.200 507.600 354.000 508.400 ;
        RECT 358.000 506.200 358.800 511.800 ;
        RECT 351.600 503.600 352.400 504.400 ;
        RECT 354.800 503.600 355.600 504.400 ;
        RECT 361.200 504.200 362.000 515.800 ;
        RECT 367.700 510.400 368.300 535.600 ;
        RECT 377.300 532.400 377.900 539.600 ;
        RECT 386.900 536.400 387.500 545.600 ;
        RECT 388.400 544.200 389.200 555.800 ;
        RECT 390.000 549.600 390.800 550.400 ;
        RECT 390.100 548.400 390.700 549.600 ;
        RECT 390.000 547.600 390.800 548.400 ;
        RECT 391.600 544.200 392.400 555.800 ;
        RECT 393.200 544.200 394.000 557.800 ;
        RECT 394.800 544.200 395.600 557.800 ;
        RECT 406.000 553.600 406.800 554.400 ;
        RECT 420.400 551.600 421.200 552.400 ;
        RECT 399.600 549.600 400.400 550.400 ;
        RECT 412.400 549.600 413.200 550.400 ;
        RECT 386.800 535.600 387.600 536.400 ;
        RECT 382.000 533.600 382.800 534.400 ;
        RECT 372.400 531.600 373.200 532.400 ;
        RECT 377.200 531.600 378.000 532.400 ;
        RECT 391.600 531.600 392.400 532.400 ;
        RECT 372.500 530.400 373.100 531.600 ;
        RECT 370.800 529.600 371.600 530.400 ;
        RECT 372.400 529.600 373.200 530.400 ;
        RECT 380.400 529.600 381.200 530.400 ;
        RECT 370.900 528.400 371.500 529.600 ;
        RECT 370.800 527.600 371.600 528.400 ;
        RECT 383.600 527.600 384.400 528.400 ;
        RECT 393.200 524.200 394.000 537.800 ;
        RECT 394.800 524.200 395.600 537.800 ;
        RECT 396.400 524.200 397.200 537.800 ;
        RECT 398.000 526.200 398.800 537.800 ;
        RECT 399.600 535.600 400.400 536.400 ;
        RECT 401.200 526.200 402.000 537.800 ;
        RECT 402.800 533.600 403.600 534.400 ;
        RECT 404.400 526.200 405.200 537.800 ;
        RECT 406.000 524.200 406.800 537.800 ;
        RECT 407.600 524.200 408.400 537.800 ;
        RECT 412.500 532.400 413.100 549.600 ;
        RECT 417.200 547.600 418.000 548.400 ;
        RECT 417.300 546.400 417.900 547.600 ;
        RECT 417.200 545.600 418.000 546.400 ;
        RECT 418.800 544.300 419.600 544.400 ;
        RECT 420.500 544.300 421.100 551.600 ;
        RECT 418.800 543.700 421.100 544.300 ;
        RECT 423.600 544.200 424.400 555.800 ;
        RECT 425.200 553.600 426.000 554.400 ;
        RECT 425.300 550.400 425.900 553.600 ;
        RECT 425.200 549.600 426.000 550.400 ;
        RECT 431.600 549.400 432.400 550.400 ;
        RECT 430.000 545.600 430.800 546.400 ;
        RECT 418.800 543.600 419.600 543.700 ;
        RECT 417.200 535.600 418.000 536.400 ;
        RECT 417.300 534.400 417.900 535.600 ;
        RECT 417.200 533.600 418.000 534.400 ;
        RECT 418.800 533.600 419.600 534.400 ;
        RECT 412.400 531.600 413.200 532.400 ;
        RECT 412.500 524.400 413.100 531.600 ;
        RECT 417.200 527.600 418.000 528.400 ;
        RECT 412.400 523.600 413.200 524.400 ;
        RECT 369.200 521.600 370.000 522.400 ;
        RECT 406.000 521.600 406.800 522.400 ;
        RECT 364.400 509.600 365.200 510.400 ;
        RECT 367.600 509.600 368.400 510.400 ;
        RECT 351.700 500.400 352.300 503.600 ;
        RECT 342.000 499.600 342.800 500.400 ;
        RECT 351.600 499.600 352.400 500.400 ;
        RECT 340.400 493.600 341.200 494.400 ;
        RECT 340.500 492.400 341.100 493.600 ;
        RECT 332.400 491.600 333.200 492.400 ;
        RECT 334.000 491.600 334.800 492.400 ;
        RECT 335.600 491.600 336.400 492.400 ;
        RECT 340.400 491.600 341.200 492.400 ;
        RECT 330.800 483.600 331.600 484.400 ;
        RECT 322.800 464.200 323.600 475.800 ;
        RECT 327.600 473.600 328.400 474.400 ;
        RECT 329.200 471.600 330.000 472.400 ;
        RECT 334.100 470.400 334.700 491.600 ;
        RECT 342.100 490.400 342.700 499.600 ;
        RECT 358.000 495.600 358.800 496.400 ;
        RECT 358.100 494.400 358.700 495.600 ;
        RECT 369.300 494.400 369.900 521.600 ;
        RECT 406.100 518.400 406.700 521.600 ;
        RECT 417.300 518.400 417.900 527.600 ;
        RECT 406.000 517.600 406.800 518.400 ;
        RECT 417.200 517.600 418.000 518.400 ;
        RECT 370.800 504.200 371.600 515.800 ;
        RECT 372.400 513.600 373.200 514.400 ;
        RECT 375.600 513.600 376.400 514.400 ;
        RECT 393.200 513.600 394.000 514.400 ;
        RECT 409.200 513.600 410.000 514.400 ;
        RECT 346.800 493.600 347.600 494.400 ;
        RECT 358.000 493.600 358.800 494.400 ;
        RECT 369.200 493.600 370.000 494.400 ;
        RECT 345.200 492.300 346.000 492.400 ;
        RECT 345.200 491.700 347.500 492.300 ;
        RECT 345.200 491.600 346.000 491.700 ;
        RECT 342.000 489.600 342.800 490.400 ;
        RECT 337.200 485.600 338.000 486.400 ;
        RECT 335.600 483.600 336.400 484.400 ;
        RECT 330.800 469.600 331.600 470.400 ;
        RECT 332.400 469.600 333.200 470.400 ;
        RECT 334.000 469.600 334.800 470.400 ;
        RECT 332.500 468.400 333.100 469.600 ;
        RECT 335.700 468.400 336.300 483.600 ;
        RECT 337.300 478.400 337.900 485.600 ;
        RECT 337.200 477.600 338.000 478.400 ;
        RECT 327.600 467.600 328.400 468.400 ;
        RECT 332.400 467.600 333.200 468.400 ;
        RECT 335.600 467.600 336.400 468.400 ;
        RECT 318.000 459.600 318.800 460.400 ;
        RECT 313.200 455.600 314.000 456.400 ;
        RECT 287.600 433.600 288.400 434.400 ;
        RECT 287.700 432.400 288.300 433.600 ;
        RECT 287.600 431.600 288.400 432.400 ;
        RECT 295.700 430.400 296.300 443.600 ;
        RECT 297.300 440.400 297.900 443.600 ;
        RECT 297.200 439.600 298.000 440.400 ;
        RECT 295.600 429.600 296.400 430.400 ;
        RECT 294.000 419.600 294.800 420.400 ;
        RECT 289.200 415.600 290.000 416.400 ;
        RECT 286.000 411.600 286.800 412.400 ;
        RECT 268.600 409.400 269.400 410.200 ;
        RECT 274.800 409.400 275.600 410.200 ;
        RECT 278.000 409.600 278.800 410.400 ;
        RECT 282.800 409.600 283.600 410.400 ;
        RECT 257.200 403.600 258.000 404.400 ;
        RECT 263.600 403.600 264.400 404.400 ;
        RECT 246.000 393.600 246.800 394.400 ;
        RECT 249.200 393.600 250.000 394.400 ;
        RECT 254.000 393.600 254.800 394.400 ;
        RECT 252.400 391.600 253.200 392.400 ;
        RECT 257.300 390.400 257.900 403.600 ;
        RECT 252.400 389.600 253.200 390.400 ;
        RECT 257.200 389.600 258.000 390.400 ;
        RECT 263.600 389.600 264.400 390.400 ;
        RECT 266.800 389.600 267.600 390.400 ;
        RECT 249.200 387.600 250.000 388.400 ;
        RECT 249.300 380.400 249.900 387.600 ;
        RECT 252.400 383.600 253.200 384.400 ;
        RECT 231.600 379.600 232.400 380.400 ;
        RECT 249.200 379.600 250.000 380.400 ;
        RECT 250.800 379.600 251.600 380.400 ;
        RECT 252.500 380.300 253.100 383.600 ;
        RECT 257.300 382.400 257.900 389.600 ;
        RECT 260.400 383.600 261.200 384.400 ;
        RECT 257.200 381.600 258.000 382.400 ;
        RECT 252.500 379.700 254.700 380.300 ;
        RECT 231.700 378.400 232.300 379.600 ;
        RECT 231.600 377.600 232.400 378.400 ;
        RECT 230.000 375.600 230.800 376.400 ;
        RECT 218.800 371.600 219.600 372.400 ;
        RECT 228.400 371.600 229.200 372.400 ;
        RECT 206.000 369.600 206.800 370.400 ;
        RECT 209.200 369.600 210.000 370.400 ;
        RECT 212.400 369.600 213.200 370.400 ;
        RECT 220.400 367.600 221.200 368.400 ;
        RECT 231.600 367.600 232.400 368.400 ;
        RECT 210.800 363.600 211.600 364.400 ;
        RECT 198.000 361.600 198.800 362.400 ;
        RECT 202.800 361.600 203.600 362.400 ;
        RECT 191.600 359.600 192.400 360.400 ;
        RECT 146.800 353.600 147.600 354.400 ;
        RECT 161.200 353.600 162.000 354.400 ;
        RECT 132.400 349.600 133.200 350.400 ;
        RECT 134.000 349.600 134.800 350.400 ;
        RECT 142.000 350.300 142.800 350.400 ;
        RECT 142.000 349.700 144.300 350.300 ;
        RECT 142.000 349.600 142.800 349.700 ;
        RECT 130.800 347.600 131.600 348.400 ;
        RECT 142.000 347.600 142.800 348.400 ;
        RECT 129.200 343.600 130.000 344.400 ;
        RECT 135.600 343.600 136.400 344.400 ;
        RECT 127.600 331.600 128.400 332.400 ;
        RECT 129.200 326.200 130.000 337.800 ;
        RECT 134.000 335.600 134.800 336.400 ;
        RECT 134.100 334.400 134.700 335.600 ;
        RECT 134.000 333.600 134.800 334.400 ;
        RECT 130.800 331.600 131.600 332.600 ;
        RECT 138.800 326.200 139.600 337.800 ;
        RECT 103.600 321.600 104.400 322.400 ;
        RECT 142.100 320.400 142.700 347.600 ;
        RECT 143.700 338.400 144.300 349.700 ;
        RECT 158.000 349.600 158.800 350.400 ;
        RECT 170.800 349.600 171.600 350.400 ;
        RECT 172.400 349.600 173.200 350.400 ;
        RECT 174.000 349.600 174.800 350.400 ;
        RECT 156.400 346.300 157.200 346.400 ;
        RECT 154.900 345.700 157.200 346.300 ;
        RECT 153.200 343.600 154.000 344.400 ;
        RECT 145.200 339.600 146.000 340.400 ;
        RECT 145.300 338.400 145.900 339.600 ;
        RECT 143.600 337.600 144.400 338.400 ;
        RECT 145.200 337.600 146.000 338.400 ;
        RECT 153.300 336.400 153.900 343.600 ;
        RECT 154.900 338.400 155.500 345.700 ;
        RECT 156.400 345.600 157.200 345.700 ;
        RECT 154.800 337.600 155.600 338.400 ;
        RECT 153.200 335.600 154.000 336.400 ;
        RECT 142.000 319.600 142.800 320.400 ;
        RECT 102.000 317.600 102.800 318.400 ;
        RECT 110.000 317.600 110.800 318.400 ;
        RECT 118.000 311.600 118.800 312.400 ;
        RECT 118.100 310.400 118.700 311.600 ;
        RECT 79.600 309.600 80.400 310.400 ;
        RECT 87.600 309.600 88.400 310.400 ;
        RECT 92.400 309.600 93.200 310.400 ;
        RECT 95.600 309.600 96.400 310.400 ;
        RECT 97.200 309.600 98.000 310.400 ;
        RECT 103.600 309.600 104.400 310.400 ;
        RECT 118.000 309.600 118.800 310.400 ;
        RECT 86.000 307.600 86.800 308.400 ;
        RECT 92.500 306.400 93.100 309.600 ;
        RECT 92.400 305.600 93.200 306.400 ;
        RECT 60.400 291.600 61.200 292.400 ;
        RECT 68.400 291.600 69.200 292.400 ;
        RECT 54.000 289.600 54.800 290.400 ;
        RECT 58.800 289.600 59.600 290.400 ;
        RECT 39.600 283.600 40.400 284.400 ;
        RECT 47.600 283.600 48.400 284.400 ;
        RECT 25.200 269.600 26.000 270.400 ;
        RECT 28.400 269.600 29.200 270.400 ;
        RECT 33.200 263.600 34.000 264.400 ;
        RECT 38.000 263.600 38.800 264.400 ;
        RECT 17.200 255.600 18.000 256.400 ;
        RECT 18.800 246.200 19.600 257.800 ;
        RECT 20.400 244.200 21.200 257.800 ;
        RECT 22.000 244.200 22.800 257.800 ;
        RECT 23.600 244.200 24.400 257.800 ;
        RECT 38.100 256.400 38.700 263.600 ;
        RECT 38.000 255.600 38.800 256.400 ;
        RECT 25.200 251.600 26.000 252.400 ;
        RECT 34.800 247.600 35.600 248.400 ;
        RECT 33.200 243.600 34.000 244.400 ;
        RECT 22.000 239.600 22.800 240.400 ;
        RECT 22.100 238.400 22.700 239.600 ;
        RECT 22.000 237.600 22.800 238.400 ;
        RECT 33.300 236.400 33.900 243.600 ;
        RECT 18.800 235.600 19.600 236.400 ;
        RECT 30.000 235.600 30.800 236.400 ;
        RECT 33.200 235.600 34.000 236.400 ;
        RECT 15.600 233.600 16.400 234.400 ;
        RECT 18.900 232.400 19.500 235.600 ;
        RECT 30.100 234.400 30.700 235.600 ;
        RECT 30.000 233.600 30.800 234.400 ;
        RECT 18.800 231.600 19.600 232.400 ;
        RECT 22.000 231.600 22.800 232.400 ;
        RECT 25.200 231.600 26.000 232.400 ;
        RECT 33.200 231.600 34.000 232.400 ;
        RECT 22.100 230.400 22.700 231.600 ;
        RECT 9.200 229.600 10.000 230.400 ;
        RECT 14.000 229.600 14.800 230.400 ;
        RECT 15.600 229.600 16.400 230.400 ;
        RECT 18.800 229.600 19.600 230.400 ;
        RECT 22.000 229.600 22.800 230.400 ;
        RECT 23.600 229.600 24.400 230.400 ;
        RECT 26.800 229.600 27.600 230.400 ;
        RECT 33.200 229.600 34.000 230.400 ;
        RECT 2.800 227.600 3.600 228.400 ;
        RECT 7.600 227.600 8.400 228.400 ;
        RECT 6.000 225.600 6.800 226.400 ;
        RECT 9.300 212.400 9.900 229.600 ;
        RECT 18.900 228.400 19.500 229.600 ;
        RECT 14.000 227.600 14.800 228.400 ;
        RECT 18.800 227.600 19.600 228.400 ;
        RECT 20.400 227.600 21.200 228.400 ;
        RECT 14.100 216.300 14.700 227.600 ;
        RECT 15.600 216.300 16.400 216.400 ;
        RECT 14.100 215.700 16.400 216.300 ;
        RECT 15.600 215.600 16.400 215.700 ;
        RECT 14.000 213.600 14.800 214.400 ;
        RECT 14.100 212.400 14.700 213.600 ;
        RECT 18.900 212.400 19.500 227.600 ;
        RECT 20.500 226.400 21.100 227.600 ;
        RECT 22.100 226.400 22.700 229.600 ;
        RECT 20.400 225.600 21.200 226.400 ;
        RECT 22.000 225.600 22.800 226.400 ;
        RECT 23.700 214.400 24.300 229.600 ;
        RECT 26.900 228.400 27.500 229.600 ;
        RECT 33.300 228.400 33.900 229.600 ;
        RECT 26.800 227.600 27.600 228.400 ;
        RECT 31.600 227.600 32.400 228.400 ;
        RECT 33.200 227.600 34.000 228.400 ;
        RECT 28.400 223.600 29.200 224.400 ;
        RECT 23.600 213.600 24.400 214.400 ;
        RECT 6.000 211.600 6.800 212.400 ;
        RECT 9.200 211.600 10.000 212.400 ;
        RECT 14.000 211.600 14.800 212.400 ;
        RECT 18.800 211.600 19.600 212.400 ;
        RECT 9.200 209.600 10.000 210.400 ;
        RECT 6.000 203.600 6.800 204.400 ;
        RECT 6.100 188.400 6.700 203.600 ;
        RECT 6.000 187.600 6.800 188.400 ;
        RECT 6.000 185.600 6.800 186.400 ;
        RECT 1.200 170.200 2.000 175.800 ;
        RECT 4.400 166.200 5.200 177.800 ;
        RECT 6.100 176.400 6.700 185.600 ;
        RECT 9.200 184.200 10.000 197.800 ;
        RECT 10.800 184.200 11.600 197.800 ;
        RECT 12.400 184.200 13.200 195.800 ;
        RECT 14.100 190.400 14.700 211.600 ;
        RECT 28.500 210.400 29.100 223.600 ;
        RECT 31.700 216.400 32.300 227.600 ;
        RECT 31.600 215.600 32.400 216.400 ;
        RECT 30.000 211.600 30.800 212.400 ;
        RECT 18.800 209.600 19.600 210.400 ;
        RECT 22.000 209.600 22.800 210.400 ;
        RECT 26.800 209.600 27.600 210.400 ;
        RECT 28.400 209.600 29.200 210.400 ;
        RECT 25.200 207.600 26.000 208.400 ;
        RECT 14.000 189.600 14.800 190.400 ;
        RECT 14.000 187.600 14.800 188.400 ;
        RECT 15.600 184.200 16.400 195.800 ;
        RECT 17.200 185.600 18.000 186.400 ;
        RECT 18.800 184.200 19.600 195.800 ;
        RECT 20.400 184.200 21.200 197.800 ;
        RECT 22.000 184.200 22.800 197.800 ;
        RECT 23.600 184.200 24.400 197.800 ;
        RECT 25.200 191.600 26.000 192.400 ;
        RECT 25.300 190.400 25.900 191.600 ;
        RECT 25.200 189.600 26.000 190.400 ;
        RECT 6.000 175.600 6.800 176.400 ;
        RECT 1.200 146.200 2.000 151.800 ;
        RECT 4.400 144.200 5.200 155.800 ;
        RECT 6.100 148.400 6.700 175.600 ;
        RECT 9.200 171.600 10.000 172.400 ;
        RECT 14.000 166.200 14.800 177.800 ;
        RECT 25.300 176.400 25.900 189.600 ;
        RECT 30.100 178.400 30.700 211.600 ;
        RECT 31.700 182.400 32.300 215.600 ;
        RECT 33.200 213.600 34.000 214.400 ;
        RECT 34.900 212.400 35.500 247.600 ;
        RECT 36.400 241.600 37.200 242.400 ;
        RECT 36.500 232.400 37.100 241.600 ;
        RECT 36.400 231.600 37.200 232.400 ;
        RECT 39.700 226.400 40.300 283.600 ;
        RECT 46.000 269.600 46.800 270.400 ;
        RECT 47.600 264.200 48.400 277.800 ;
        RECT 49.200 264.200 50.000 277.800 ;
        RECT 50.800 264.200 51.600 277.800 ;
        RECT 52.400 264.200 53.200 275.800 ;
        RECT 54.100 270.400 54.700 289.600 ;
        RECT 54.000 269.600 54.800 270.400 ;
        RECT 54.000 265.600 54.800 266.400 ;
        RECT 54.100 260.300 54.700 265.600 ;
        RECT 55.600 264.200 56.400 275.800 ;
        RECT 57.200 267.600 58.000 268.400 ;
        RECT 57.300 266.400 57.900 267.600 ;
        RECT 57.200 265.600 58.000 266.400 ;
        RECT 58.800 264.200 59.600 275.800 ;
        RECT 60.400 264.200 61.200 277.800 ;
        RECT 62.000 264.200 62.800 277.800 ;
        RECT 68.500 272.400 69.100 291.600 ;
        RECT 70.000 284.200 70.800 297.800 ;
        RECT 71.600 284.200 72.400 297.800 ;
        RECT 73.200 286.200 74.000 297.800 ;
        RECT 74.800 293.600 75.600 294.400 ;
        RECT 74.900 292.400 75.500 293.600 ;
        RECT 74.800 291.600 75.600 292.400 ;
        RECT 76.400 286.200 77.200 297.800 ;
        RECT 78.000 295.600 78.800 296.400 ;
        RECT 78.100 294.400 78.700 295.600 ;
        RECT 78.000 293.600 78.800 294.400 ;
        RECT 79.600 286.200 80.400 297.800 ;
        RECT 81.200 284.200 82.000 297.800 ;
        RECT 82.800 284.200 83.600 297.800 ;
        RECT 84.400 284.200 85.200 297.800 ;
        RECT 86.000 295.600 86.800 296.400 ;
        RECT 81.200 279.600 82.000 280.400 ;
        RECT 65.200 271.600 66.000 272.400 ;
        RECT 68.400 271.600 69.200 272.400 ;
        RECT 65.300 270.400 65.900 271.600 ;
        RECT 81.300 270.400 81.900 279.600 ;
        RECT 84.400 278.300 85.200 278.400 ;
        RECT 86.100 278.300 86.700 295.600 ;
        RECT 89.200 283.600 90.000 284.400 ;
        RECT 84.400 277.700 86.700 278.300 ;
        RECT 84.400 277.600 85.200 277.700 ;
        RECT 84.400 273.600 85.200 274.400 ;
        RECT 65.200 269.600 66.000 270.400 ;
        RECT 74.800 269.600 75.600 270.400 ;
        RECT 78.000 269.600 78.800 270.400 ;
        RECT 81.200 269.600 82.000 270.400 ;
        RECT 74.800 267.600 75.600 268.400 ;
        RECT 78.100 268.300 78.700 269.600 ;
        RECT 79.600 268.300 80.400 268.400 ;
        RECT 78.100 267.700 80.400 268.300 ;
        RECT 71.600 265.600 72.400 266.400 ;
        RECT 71.700 264.400 72.300 265.600 ;
        RECT 71.600 263.600 72.400 264.400 ;
        RECT 54.100 259.700 56.300 260.300 ;
        RECT 41.200 251.600 42.000 252.400 ;
        RECT 47.600 244.200 48.400 257.800 ;
        RECT 49.200 244.200 50.000 257.800 ;
        RECT 50.800 246.200 51.600 257.800 ;
        RECT 52.400 253.600 53.200 254.400 ;
        RECT 50.800 243.600 51.600 244.400 ;
        RECT 47.600 229.600 48.400 230.400 ;
        RECT 42.800 227.600 43.600 228.400 ;
        RECT 39.600 225.600 40.400 226.400 ;
        RECT 41.200 225.600 42.000 226.400 ;
        RECT 38.000 223.600 38.800 224.400 ;
        RECT 38.100 212.400 38.700 223.600 ;
        RECT 39.600 213.600 40.400 214.400 ;
        RECT 46.000 213.600 46.800 214.400 ;
        RECT 34.800 211.600 35.600 212.400 ;
        RECT 38.000 211.600 38.800 212.400 ;
        RECT 41.200 211.600 42.000 212.400 ;
        RECT 33.200 209.600 34.000 210.400 ;
        RECT 34.800 209.600 35.600 210.400 ;
        RECT 33.300 198.400 33.900 209.600 ;
        RECT 34.900 208.400 35.500 209.600 ;
        RECT 34.800 207.600 35.600 208.400 ;
        RECT 38.000 203.600 38.800 204.400 ;
        RECT 33.200 197.600 34.000 198.400 ;
        RECT 38.100 194.400 38.700 203.600 ;
        RECT 38.000 193.600 38.800 194.400 ;
        RECT 38.100 188.400 38.700 193.600 ;
        RECT 33.200 187.600 34.000 188.400 ;
        RECT 38.000 187.600 38.800 188.400 ;
        RECT 31.600 181.600 32.400 182.400 ;
        RECT 30.000 177.600 30.800 178.400 ;
        RECT 25.200 175.600 26.000 176.400 ;
        RECT 30.000 175.600 30.800 176.400 ;
        RECT 25.200 173.600 26.000 174.400 ;
        RECT 20.400 171.600 21.200 172.400 ;
        RECT 23.600 171.600 24.400 172.400 ;
        RECT 20.400 169.600 21.200 170.400 ;
        RECT 23.600 169.600 24.400 170.400 ;
        RECT 18.800 167.600 19.600 168.400 ;
        RECT 20.400 167.600 21.200 168.400 ;
        RECT 7.600 149.600 8.400 150.400 ;
        RECT 6.000 147.600 6.800 148.400 ;
        RECT 6.100 136.400 6.700 147.600 ;
        RECT 14.000 144.200 14.800 155.800 ;
        RECT 20.500 152.400 21.100 167.600 ;
        RECT 23.700 158.400 24.300 169.600 ;
        RECT 23.600 157.600 24.400 158.400 ;
        RECT 20.400 151.600 21.200 152.400 ;
        RECT 18.800 147.600 19.600 148.400 ;
        RECT 18.900 144.400 19.500 147.600 ;
        RECT 25.300 144.400 25.900 173.600 ;
        RECT 26.800 171.600 27.600 172.400 ;
        RECT 28.400 171.600 29.200 172.400 ;
        RECT 26.900 160.400 27.500 171.600 ;
        RECT 28.500 168.400 29.100 171.600 ;
        RECT 28.400 167.600 29.200 168.400 ;
        RECT 26.800 159.600 27.600 160.400 ;
        RECT 28.500 158.400 29.100 167.600 ;
        RECT 28.400 157.600 29.200 158.400 ;
        RECT 26.800 153.600 27.600 154.400 ;
        RECT 26.900 148.400 27.500 153.600 ;
        RECT 28.400 149.600 29.200 150.400 ;
        RECT 26.800 147.600 27.600 148.400 ;
        RECT 18.800 143.600 19.600 144.400 ;
        RECT 25.200 143.600 26.000 144.400 ;
        RECT 6.000 135.600 6.800 136.400 ;
        RECT 2.800 129.600 3.600 130.400 ;
        RECT 2.900 124.400 3.500 129.600 ;
        RECT 2.800 123.600 3.600 124.400 ;
        RECT 1.200 106.200 2.000 111.800 ;
        RECT 1.200 87.600 2.000 88.400 ;
        RECT 2.900 64.400 3.500 123.600 ;
        RECT 4.400 104.200 5.200 115.800 ;
        RECT 6.100 108.400 6.700 135.600 ;
        RECT 10.800 131.600 11.600 132.400 ;
        RECT 9.200 109.600 10.000 110.400 ;
        RECT 6.000 107.600 6.800 108.400 ;
        RECT 6.000 86.200 6.800 97.800 ;
        RECT 10.900 74.400 11.500 131.600 ;
        RECT 12.400 124.200 13.200 137.800 ;
        RECT 14.000 124.200 14.800 137.800 ;
        RECT 15.600 124.200 16.400 137.800 ;
        RECT 17.200 126.200 18.000 137.800 ;
        RECT 18.800 135.600 19.600 136.400 ;
        RECT 20.400 126.200 21.200 137.800 ;
        RECT 22.000 135.600 22.800 136.400 ;
        RECT 22.100 134.400 22.700 135.600 ;
        RECT 22.000 133.600 22.800 134.400 ;
        RECT 23.600 126.200 24.400 137.800 ;
        RECT 25.200 124.200 26.000 137.800 ;
        RECT 26.800 124.200 27.600 137.800 ;
        RECT 14.000 104.200 14.800 115.800 ;
        RECT 23.600 115.600 24.400 116.400 ;
        RECT 18.800 113.600 19.600 114.400 ;
        RECT 20.400 111.600 21.200 112.400 ;
        RECT 20.500 108.400 21.100 111.600 ;
        RECT 23.700 110.400 24.300 115.600 ;
        RECT 26.800 113.600 27.600 114.400 ;
        RECT 26.900 112.400 27.500 113.600 ;
        RECT 26.800 111.600 27.600 112.400 ;
        RECT 28.500 112.300 29.100 149.600 ;
        RECT 30.100 132.400 30.700 175.600 ;
        RECT 33.300 172.400 33.900 187.600 ;
        RECT 38.000 185.600 38.800 186.400 ;
        RECT 39.600 186.200 40.400 191.800 ;
        RECT 41.300 188.400 41.900 211.600 ;
        RECT 41.200 187.600 42.000 188.400 ;
        RECT 41.300 186.400 41.900 187.600 ;
        RECT 41.200 185.600 42.000 186.400 ;
        RECT 38.100 184.400 38.700 185.600 ;
        RECT 36.400 183.600 37.200 184.400 ;
        RECT 38.000 183.600 38.800 184.400 ;
        RECT 42.800 184.200 43.600 195.800 ;
        RECT 31.600 171.600 32.400 172.400 ;
        RECT 33.200 171.600 34.000 172.400 ;
        RECT 36.500 152.400 37.100 183.600 ;
        RECT 38.000 181.600 38.800 182.400 ;
        RECT 38.100 178.400 38.700 181.600 ;
        RECT 38.000 177.600 38.800 178.400 ;
        RECT 39.600 177.600 40.400 178.400 ;
        RECT 38.000 163.600 38.800 164.400 ;
        RECT 38.100 154.400 38.700 163.600 ;
        RECT 38.000 153.600 38.800 154.400 ;
        RECT 31.600 151.600 32.400 152.400 ;
        RECT 36.400 151.600 37.200 152.400 ;
        RECT 31.700 148.400 32.300 151.600 ;
        RECT 39.700 150.400 40.300 177.600 ;
        RECT 46.100 176.300 46.700 213.600 ;
        RECT 47.700 192.400 48.300 229.600 ;
        RECT 47.600 191.600 48.400 192.400 ;
        RECT 47.600 189.600 48.400 190.400 ;
        RECT 49.200 185.600 50.000 186.400 ;
        RECT 46.100 175.700 48.300 176.300 ;
        RECT 41.200 171.600 42.000 172.400 ;
        RECT 41.300 168.400 41.900 171.600 ;
        RECT 42.800 169.600 43.600 170.400 ;
        RECT 41.200 167.600 42.000 168.400 ;
        RECT 33.200 149.600 34.000 150.400 ;
        RECT 36.400 149.600 37.200 150.400 ;
        RECT 39.600 149.600 40.400 150.400 ;
        RECT 33.300 148.400 33.900 149.600 ;
        RECT 31.600 147.600 32.400 148.400 ;
        RECT 33.200 147.600 34.000 148.400 ;
        RECT 36.500 146.400 37.100 149.600 ;
        RECT 38.000 147.600 38.800 148.400 ;
        RECT 39.600 147.600 40.400 148.400 ;
        RECT 36.400 145.600 37.200 146.400 ;
        RECT 38.100 144.400 38.700 147.600 ;
        RECT 39.700 146.400 40.300 147.600 ;
        RECT 39.600 145.600 40.400 146.400 ;
        RECT 38.000 143.600 38.800 144.400 ;
        RECT 41.300 142.400 41.900 167.600 ;
        RECT 38.000 141.600 38.800 142.400 ;
        RECT 41.200 141.600 42.000 142.400 ;
        RECT 36.400 134.300 37.200 134.400 ;
        RECT 34.900 133.700 37.200 134.300 ;
        RECT 30.000 131.600 30.800 132.400 ;
        RECT 33.200 131.600 34.000 132.400 ;
        RECT 30.000 112.300 30.800 112.400 ;
        RECT 28.500 111.700 30.800 112.300 ;
        RECT 30.000 111.600 30.800 111.700 ;
        RECT 30.100 110.400 30.700 111.600 ;
        RECT 22.000 109.600 22.800 110.400 ;
        RECT 23.600 109.600 24.400 110.400 ;
        RECT 30.000 109.600 30.800 110.400 ;
        RECT 20.400 107.600 21.200 108.400 ;
        RECT 25.200 107.600 26.000 108.400 ;
        RECT 26.800 107.600 27.600 108.400 ;
        RECT 25.300 106.400 25.900 107.600 ;
        RECT 25.200 105.600 26.000 106.400 ;
        RECT 26.800 105.600 27.600 106.400 ;
        RECT 20.400 103.600 21.200 104.400 ;
        RECT 20.500 98.400 21.100 103.600 ;
        RECT 12.400 93.600 13.200 94.400 ;
        RECT 7.600 73.600 8.400 74.400 ;
        RECT 10.800 73.600 11.600 74.400 ;
        RECT 6.000 69.600 6.800 70.400 ;
        RECT 2.800 63.600 3.600 64.400 ;
        RECT 6.100 30.400 6.700 69.600 ;
        RECT 7.700 52.400 8.300 73.600 ;
        RECT 10.800 71.600 11.600 72.400 ;
        RECT 9.200 63.600 10.000 64.400 ;
        RECT 9.300 62.400 9.900 63.600 ;
        RECT 9.200 61.600 10.000 62.400 ;
        RECT 12.500 60.400 13.100 93.600 ;
        RECT 14.000 91.800 14.800 92.600 ;
        RECT 14.100 90.400 14.700 91.800 ;
        RECT 14.000 89.600 14.800 90.400 ;
        RECT 15.600 86.200 16.400 97.800 ;
        RECT 20.400 97.600 21.200 98.400 ;
        RECT 18.800 90.200 19.600 95.800 ;
        RECT 23.600 95.600 24.400 96.400 ;
        RECT 22.000 93.600 22.800 94.400 ;
        RECT 20.400 89.600 21.200 90.400 ;
        RECT 20.500 74.400 21.100 89.600 ;
        RECT 20.400 73.600 21.200 74.400 ;
        RECT 17.200 71.600 18.000 72.400 ;
        RECT 14.000 69.600 14.800 70.400 ;
        RECT 14.100 64.400 14.700 69.600 ;
        RECT 15.600 67.600 16.400 68.400 ;
        RECT 14.000 63.600 14.800 64.400 ;
        RECT 15.700 62.400 16.300 67.600 ;
        RECT 17.300 66.400 17.900 71.600 ;
        RECT 22.100 68.400 22.700 93.600 ;
        RECT 23.700 92.400 24.300 95.600 ;
        RECT 26.900 94.400 27.500 105.600 ;
        RECT 31.600 97.600 32.400 98.400 ;
        RECT 25.200 93.600 26.000 94.400 ;
        RECT 26.800 93.600 27.600 94.400 ;
        RECT 23.600 91.600 24.400 92.400 ;
        RECT 23.600 83.600 24.400 84.400 ;
        RECT 23.700 70.400 24.300 83.600 ;
        RECT 26.900 72.400 27.500 93.600 ;
        RECT 28.400 91.600 29.200 92.400 ;
        RECT 31.700 90.400 32.300 97.600 ;
        RECT 33.300 94.400 33.900 131.600 ;
        RECT 34.900 118.400 35.500 133.700 ;
        RECT 36.400 133.600 37.200 133.700 ;
        RECT 34.800 117.600 35.600 118.400 ;
        RECT 38.100 110.400 38.700 141.600 ;
        RECT 41.200 135.600 42.000 136.400 ;
        RECT 39.600 129.600 40.400 130.400 ;
        RECT 42.900 130.300 43.500 169.600 ;
        RECT 46.100 166.300 46.700 175.700 ;
        RECT 47.700 174.400 48.300 175.700 ;
        RECT 47.600 173.600 48.400 174.400 ;
        RECT 44.500 165.700 46.700 166.300 ;
        RECT 44.500 132.400 45.100 165.700 ;
        RECT 46.000 163.600 46.800 164.400 ;
        RECT 46.100 152.400 46.700 163.600 ;
        RECT 46.000 151.600 46.800 152.400 ;
        RECT 49.300 152.300 49.900 185.600 ;
        RECT 50.900 176.400 51.500 243.600 ;
        RECT 52.500 240.400 53.100 253.600 ;
        RECT 54.000 246.200 54.800 257.800 ;
        RECT 55.700 256.400 56.300 259.700 ;
        RECT 55.600 255.600 56.400 256.400 ;
        RECT 57.200 246.200 58.000 257.800 ;
        RECT 58.800 244.200 59.600 257.800 ;
        RECT 60.400 244.200 61.200 257.800 ;
        RECT 62.000 244.200 62.800 257.800 ;
        RECT 74.800 255.600 75.600 256.400 ;
        RECT 78.100 252.400 78.700 267.700 ;
        RECT 79.600 267.600 80.400 267.700 ;
        RECT 82.800 267.600 83.600 268.400 ;
        RECT 81.200 265.600 82.000 266.400 ;
        RECT 81.300 258.400 81.900 265.600 ;
        RECT 81.200 257.600 82.000 258.400 ;
        RECT 82.900 254.400 83.500 267.600 ;
        RECT 82.800 253.600 83.600 254.400 ;
        RECT 84.500 252.400 85.100 273.600 ;
        RECT 87.600 267.600 88.400 268.400 ;
        RECT 87.700 252.400 88.300 267.600 ;
        RECT 89.300 256.400 89.900 283.600 ;
        RECT 92.500 274.400 93.100 305.600 ;
        RECT 95.700 290.400 96.300 309.600 ;
        RECT 97.300 308.400 97.900 309.600 ;
        RECT 103.700 308.400 104.300 309.600 ;
        RECT 97.200 307.600 98.000 308.400 ;
        RECT 103.600 307.600 104.400 308.400 ;
        RECT 95.600 289.600 96.400 290.400 ;
        RECT 94.000 283.600 94.800 284.400 ;
        RECT 97.300 280.400 97.900 307.600 ;
        RECT 119.600 304.200 120.400 317.800 ;
        RECT 121.200 304.200 122.000 317.800 ;
        RECT 122.800 304.200 123.600 317.800 ;
        RECT 124.400 304.200 125.200 315.800 ;
        RECT 126.000 305.600 126.800 306.400 ;
        RECT 122.800 301.600 123.600 302.400 ;
        RECT 122.900 298.400 123.500 301.600 ;
        RECT 122.800 297.600 123.600 298.400 ;
        RECT 126.100 296.400 126.700 305.600 ;
        RECT 127.600 304.200 128.400 315.800 ;
        RECT 129.200 309.600 130.000 310.400 ;
        RECT 129.300 308.400 129.900 309.600 ;
        RECT 129.200 307.600 130.000 308.400 ;
        RECT 130.800 304.200 131.600 315.800 ;
        RECT 132.400 304.200 133.200 317.800 ;
        RECT 134.000 304.200 134.800 317.800 ;
        RECT 137.200 311.600 138.000 312.400 ;
        RECT 137.300 310.400 137.900 311.600 ;
        RECT 158.100 310.400 158.700 349.600 ;
        RECT 169.200 343.600 170.000 344.400 ;
        RECT 169.300 342.400 169.900 343.600 ;
        RECT 169.200 341.600 170.000 342.400 ;
        RECT 172.500 340.400 173.100 349.600 ;
        RECT 174.100 344.400 174.700 349.600 ;
        RECT 174.000 343.600 174.800 344.400 ;
        RECT 186.800 344.200 187.600 357.800 ;
        RECT 188.400 344.200 189.200 357.800 ;
        RECT 190.000 344.200 190.800 355.800 ;
        RECT 191.700 348.400 192.300 359.600 ;
        RECT 191.600 347.600 192.400 348.400 ;
        RECT 193.200 344.200 194.000 355.800 ;
        RECT 194.800 345.600 195.600 346.400 ;
        RECT 194.900 342.400 195.500 345.600 ;
        RECT 196.400 344.200 197.200 355.800 ;
        RECT 198.000 344.200 198.800 357.800 ;
        RECT 199.600 344.200 200.400 357.800 ;
        RECT 201.200 344.200 202.000 357.800 ;
        RECT 202.900 350.400 203.500 361.600 ;
        RECT 210.900 360.400 211.500 363.600 ;
        RECT 218.800 361.600 219.600 362.400 ;
        RECT 210.800 359.600 211.600 360.400 ;
        RECT 210.800 357.600 211.600 358.400 ;
        RECT 218.900 350.400 219.500 361.600 ;
        RECT 220.500 358.400 221.100 367.600 ;
        RECT 222.000 361.600 222.800 362.400 ;
        RECT 222.100 358.400 222.700 361.600 ;
        RECT 220.400 357.600 221.200 358.400 ;
        RECT 222.000 357.600 222.800 358.400 ;
        RECT 202.800 349.600 203.600 350.400 ;
        RECT 212.400 349.600 213.200 350.400 ;
        RECT 218.800 349.600 219.600 350.400 ;
        RECT 212.500 348.400 213.100 349.600 ;
        RECT 212.400 347.600 213.200 348.400 ;
        RECT 174.000 341.600 174.800 342.400 ;
        RECT 194.800 341.600 195.600 342.400 ;
        RECT 210.800 341.600 211.600 342.400 ;
        RECT 172.400 339.600 173.200 340.400 ;
        RECT 164.400 324.200 165.200 337.800 ;
        RECT 166.000 324.200 166.800 337.800 ;
        RECT 167.600 324.200 168.400 337.800 ;
        RECT 169.200 326.200 170.000 337.800 ;
        RECT 170.800 335.600 171.600 336.400 ;
        RECT 172.400 326.200 173.200 337.800 ;
        RECT 174.100 334.400 174.700 341.600 ;
        RECT 196.400 339.600 197.200 340.400 ;
        RECT 174.000 333.600 174.800 334.400 ;
        RECT 175.600 326.200 176.400 337.800 ;
        RECT 177.200 324.200 178.000 337.800 ;
        RECT 178.800 324.200 179.600 337.800 ;
        RECT 191.600 333.600 192.400 334.400 ;
        RECT 191.700 332.400 192.300 333.600 ;
        RECT 180.400 331.600 181.200 332.400 ;
        RECT 183.600 331.600 184.400 332.400 ;
        RECT 188.400 331.600 189.200 332.400 ;
        RECT 191.600 331.600 192.400 332.400 ;
        RECT 161.200 317.600 162.000 318.400 ;
        RECT 169.200 311.600 170.000 312.400 ;
        RECT 169.300 310.400 169.900 311.600 ;
        RECT 137.200 309.600 138.000 310.400 ;
        RECT 146.800 309.600 147.600 310.400 ;
        RECT 156.400 309.600 157.200 310.400 ;
        RECT 158.000 309.600 158.800 310.400 ;
        RECT 169.200 309.600 170.000 310.400 ;
        RECT 156.500 308.400 157.100 309.600 ;
        RECT 156.400 307.600 157.200 308.400 ;
        RECT 143.600 305.600 144.400 306.400 ;
        RECT 143.700 302.400 144.300 305.600 ;
        RECT 154.800 303.600 155.600 304.400 ;
        RECT 143.600 301.600 144.400 302.400 ;
        RECT 108.400 295.600 109.200 296.400 ;
        RECT 126.000 295.600 126.800 296.400 ;
        RECT 100.400 293.600 101.200 294.400 ;
        RECT 105.200 293.600 106.000 294.400 ;
        RECT 100.500 292.400 101.100 293.600 ;
        RECT 100.400 291.600 101.200 292.400 ;
        RECT 102.000 291.600 102.800 292.400 ;
        RECT 106.800 291.600 107.600 292.400 ;
        RECT 110.000 291.600 110.800 292.400 ;
        RECT 111.600 291.600 112.400 292.400 ;
        RECT 113.200 291.600 114.000 292.400 ;
        RECT 118.000 291.600 118.800 292.400 ;
        RECT 121.200 291.600 122.000 292.400 ;
        RECT 97.200 279.600 98.000 280.400 ;
        RECT 92.400 273.600 93.200 274.400 ;
        RECT 92.400 271.600 93.200 272.400 ;
        RECT 92.500 270.400 93.100 271.600 ;
        RECT 92.400 269.600 93.200 270.400 ;
        RECT 90.800 265.600 91.600 266.400 ;
        RECT 90.900 258.400 91.500 265.600 ;
        RECT 94.000 264.200 94.800 277.800 ;
        RECT 95.600 264.200 96.400 277.800 ;
        RECT 97.200 264.200 98.000 277.800 ;
        RECT 98.800 264.200 99.600 275.800 ;
        RECT 100.500 268.400 101.100 291.600 ;
        RECT 106.900 286.400 107.500 291.600 ;
        RECT 111.700 290.400 112.300 291.600 ;
        RECT 111.600 289.600 112.400 290.400 ;
        RECT 113.300 286.400 113.900 291.600 ;
        RECT 106.800 285.600 107.600 286.400 ;
        RECT 113.200 285.600 114.000 286.400 ;
        RECT 114.800 283.600 115.600 284.400 ;
        RECT 100.400 267.600 101.200 268.400 ;
        RECT 100.400 265.600 101.200 266.400 ;
        RECT 90.800 257.600 91.600 258.400 ;
        RECT 100.500 256.400 101.100 265.600 ;
        RECT 102.000 264.200 102.800 275.800 ;
        RECT 103.600 269.600 104.400 270.400 ;
        RECT 103.700 268.400 104.300 269.600 ;
        RECT 103.600 267.600 104.400 268.400 ;
        RECT 105.200 264.200 106.000 275.800 ;
        RECT 106.800 264.200 107.600 277.800 ;
        RECT 108.400 264.200 109.200 277.800 ;
        RECT 114.900 270.400 115.500 283.600 ;
        RECT 113.200 269.600 114.000 270.400 ;
        RECT 114.800 269.600 115.600 270.400 ;
        RECT 113.300 268.400 113.900 269.600 ;
        RECT 121.300 268.400 121.900 291.600 ;
        RECT 122.800 283.600 123.600 284.400 ;
        RECT 122.900 276.400 123.500 283.600 ;
        RECT 126.100 278.400 126.700 295.600 ;
        RECT 132.400 284.200 133.200 297.800 ;
        RECT 134.000 284.200 134.800 297.800 ;
        RECT 135.600 284.200 136.400 297.800 ;
        RECT 137.200 286.200 138.000 297.800 ;
        RECT 138.800 295.600 139.600 296.400 ;
        RECT 140.400 286.200 141.200 297.800 ;
        RECT 142.000 293.600 142.800 294.400 ;
        RECT 143.600 286.200 144.400 297.800 ;
        RECT 143.600 283.600 144.400 284.400 ;
        RECT 145.200 284.200 146.000 297.800 ;
        RECT 146.800 284.200 147.600 297.800 ;
        RECT 154.900 294.400 155.500 303.600 ;
        RECT 154.800 293.600 155.600 294.400 ;
        RECT 156.500 292.400 157.100 307.600 ;
        RECT 158.100 302.400 158.700 309.600 ;
        RECT 161.200 303.600 162.000 304.400 ;
        RECT 169.200 303.600 170.000 304.400 ;
        RECT 170.800 304.200 171.600 317.800 ;
        RECT 172.400 304.200 173.200 317.800 ;
        RECT 174.000 304.200 174.800 317.800 ;
        RECT 175.600 304.200 176.400 315.800 ;
        RECT 177.200 305.600 178.000 306.400 ;
        RECT 158.000 301.600 158.800 302.400 ;
        RECT 161.300 296.400 161.900 303.600 ;
        RECT 169.300 298.400 169.900 303.600 ;
        RECT 169.200 297.600 170.000 298.400 ;
        RECT 177.300 296.400 177.900 305.600 ;
        RECT 178.800 304.200 179.600 315.800 ;
        RECT 180.500 310.400 181.100 331.600 ;
        RECT 188.500 330.400 189.100 331.600 ;
        RECT 188.400 329.600 189.200 330.400 ;
        RECT 196.500 318.400 197.100 339.600 ;
        RECT 202.800 324.200 203.600 337.800 ;
        RECT 204.400 324.200 205.200 337.800 ;
        RECT 206.000 326.200 206.800 337.800 ;
        RECT 207.600 333.600 208.400 334.400 ;
        RECT 207.700 324.400 208.300 333.600 ;
        RECT 209.200 326.200 210.000 337.800 ;
        RECT 210.900 336.400 211.500 341.600 ;
        RECT 210.800 335.600 211.600 336.400 ;
        RECT 207.600 323.600 208.400 324.400 ;
        RECT 210.900 322.400 211.500 335.600 ;
        RECT 212.400 326.200 213.200 337.800 ;
        RECT 214.000 324.200 214.800 337.800 ;
        RECT 215.600 324.200 216.400 337.800 ;
        RECT 217.200 324.200 218.000 337.800 ;
        RECT 220.500 332.400 221.100 357.600 ;
        RECT 228.400 349.600 229.200 350.400 ;
        RECT 226.800 341.600 227.600 342.400 ;
        RECT 226.900 338.400 227.500 341.600 ;
        RECT 226.800 337.600 227.600 338.400 ;
        RECT 218.800 331.600 219.600 332.400 ;
        RECT 220.400 331.600 221.200 332.400 ;
        RECT 218.900 326.400 219.500 331.600 ;
        RECT 231.700 330.400 232.300 367.600 ;
        RECT 244.400 364.200 245.200 377.800 ;
        RECT 246.000 364.200 246.800 377.800 ;
        RECT 247.600 364.200 248.400 377.800 ;
        RECT 249.200 366.200 250.000 377.800 ;
        RECT 250.900 376.400 251.500 379.600 ;
        RECT 250.800 375.600 251.600 376.400 ;
        RECT 234.800 359.600 235.600 360.400 ;
        RECT 233.200 349.600 234.000 350.400 ;
        RECT 233.300 348.400 233.900 349.600 ;
        RECT 233.200 347.600 234.000 348.400 ;
        RECT 234.900 338.400 235.500 359.600 ;
        RECT 238.000 349.600 238.800 350.400 ;
        RECT 236.400 345.600 237.200 346.400 ;
        RECT 234.800 337.600 235.600 338.400 ;
        RECT 231.600 329.600 232.400 330.400 ;
        RECT 218.800 325.600 219.600 326.400 ;
        RECT 210.800 321.600 211.600 322.400 ;
        RECT 217.200 321.600 218.000 322.400 ;
        RECT 180.400 309.600 181.200 310.400 ;
        RECT 180.400 307.600 181.200 308.400 ;
        RECT 180.500 304.400 181.100 307.600 ;
        RECT 180.400 303.600 181.200 304.400 ;
        RECT 182.000 304.200 182.800 315.800 ;
        RECT 183.600 304.200 184.400 317.800 ;
        RECT 185.200 304.200 186.000 317.800 ;
        RECT 196.400 317.600 197.200 318.400 ;
        RECT 191.600 311.600 192.400 312.400 ;
        RECT 194.800 311.600 195.600 312.400 ;
        RECT 204.400 311.600 205.200 312.400 ;
        RECT 191.700 310.400 192.300 311.600 ;
        RECT 191.600 309.600 192.400 310.400 ;
        RECT 186.800 303.600 187.600 304.400 ;
        RECT 161.200 295.600 162.000 296.400 ;
        RECT 177.200 295.600 178.000 296.400 ;
        RECT 151.600 291.600 152.400 292.400 ;
        RECT 156.400 291.600 157.200 292.400 ;
        RECT 164.400 291.600 165.200 292.400 ;
        RECT 166.000 291.600 166.800 292.400 ;
        RECT 175.600 291.600 176.400 292.400 ;
        RECT 151.700 288.400 152.300 291.600 ;
        RECT 151.600 287.600 152.400 288.400 ;
        RECT 126.000 277.600 126.800 278.400 ;
        RECT 122.800 275.600 123.600 276.400 ;
        RECT 130.800 275.600 131.600 276.400 ;
        RECT 122.800 273.600 123.600 274.400 ;
        RECT 122.900 270.400 123.500 273.600 ;
        RECT 122.800 269.600 123.600 270.400 ;
        RECT 113.200 267.600 114.000 268.400 ;
        RECT 121.200 267.600 122.000 268.400 ;
        RECT 124.400 267.600 125.200 268.400 ;
        RECT 118.000 265.600 118.800 266.400 ;
        RECT 119.600 263.600 120.400 264.400 ;
        RECT 119.700 260.400 120.300 263.600 ;
        RECT 114.800 259.600 115.600 260.400 ;
        RECT 119.600 259.600 120.400 260.400 ;
        RECT 89.200 255.600 90.000 256.400 ;
        RECT 100.400 255.600 101.200 256.400 ;
        RECT 63.600 251.600 64.400 252.400 ;
        RECT 68.400 251.600 69.200 252.400 ;
        RECT 78.000 251.600 78.800 252.400 ;
        RECT 84.400 251.600 85.200 252.400 ;
        RECT 87.600 251.600 88.400 252.400 ;
        RECT 52.400 239.600 53.200 240.400 ;
        RECT 52.400 224.200 53.200 237.800 ;
        RECT 54.000 224.200 54.800 237.800 ;
        RECT 55.600 224.200 56.400 235.800 ;
        RECT 57.200 227.600 58.000 228.400 ;
        RECT 58.800 224.200 59.600 235.800 ;
        RECT 60.400 225.600 61.200 226.400 ;
        RECT 55.600 221.600 56.400 222.400 ;
        RECT 55.700 214.400 56.300 221.600 ;
        RECT 60.500 220.400 61.100 225.600 ;
        RECT 62.000 224.200 62.800 235.800 ;
        RECT 63.600 224.200 64.400 237.800 ;
        RECT 65.200 224.200 66.000 237.800 ;
        RECT 66.800 224.200 67.600 237.800 ;
        RECT 68.500 230.400 69.100 251.600 ;
        RECT 71.600 243.600 72.400 244.400 ;
        RECT 86.000 243.600 86.800 244.400 ;
        RECT 95.600 243.600 96.400 244.400 ;
        RECT 105.200 244.200 106.000 257.800 ;
        RECT 106.800 244.200 107.600 257.800 ;
        RECT 108.400 244.200 109.200 257.800 ;
        RECT 110.000 246.200 110.800 257.800 ;
        RECT 111.600 255.600 112.400 256.400 ;
        RECT 113.200 246.200 114.000 257.800 ;
        RECT 114.900 254.400 115.500 259.600 ;
        RECT 114.800 253.600 115.600 254.400 ;
        RECT 116.400 246.200 117.200 257.800 ;
        RECT 118.000 244.200 118.800 257.800 ;
        RECT 119.600 244.200 120.400 257.800 ;
        RECT 124.500 252.400 125.100 267.600 ;
        RECT 126.000 263.600 126.800 264.400 ;
        RECT 126.100 256.400 126.700 263.600 ;
        RECT 130.900 256.400 131.500 275.600 ;
        RECT 138.800 267.600 139.600 268.400 ;
        RECT 126.000 255.600 126.800 256.400 ;
        RECT 130.800 255.600 131.600 256.400 ;
        RECT 130.800 253.600 131.600 254.400 ;
        RECT 130.900 252.400 131.500 253.600 ;
        RECT 124.400 251.600 125.200 252.400 ;
        RECT 130.800 251.600 131.600 252.400 ;
        RECT 137.200 251.600 138.000 252.400 ;
        RECT 129.200 243.600 130.000 244.400 ;
        RECT 135.600 243.600 136.400 244.400 ;
        RECT 71.700 242.400 72.300 243.600 ;
        RECT 71.600 241.600 72.400 242.400 ;
        RECT 78.000 241.600 78.800 242.400 ;
        RECT 78.100 234.400 78.700 241.600 ;
        RECT 78.000 233.600 78.800 234.400 ;
        RECT 82.800 233.600 83.600 234.400 ;
        RECT 68.400 229.600 69.200 230.400 ;
        RECT 76.400 229.600 77.400 230.400 ;
        RECT 82.800 229.600 83.600 230.400 ;
        RECT 68.500 226.400 69.100 229.600 ;
        RECT 82.900 228.400 83.500 229.600 ;
        RECT 82.800 227.600 83.600 228.400 ;
        RECT 84.400 227.600 85.200 228.400 ;
        RECT 68.400 225.600 69.200 226.400 ;
        RECT 84.500 222.400 85.100 227.600 ;
        RECT 84.400 221.600 85.200 222.400 ;
        RECT 60.400 219.600 61.200 220.400 ;
        RECT 66.800 219.600 67.600 220.400 ;
        RECT 66.900 218.400 67.500 219.600 ;
        RECT 66.800 217.600 67.600 218.400 ;
        RECT 74.800 215.600 75.600 216.400 ;
        RECT 55.600 213.600 56.400 214.400 ;
        RECT 68.400 211.600 69.200 212.400 ;
        RECT 71.600 211.600 72.400 212.400 ;
        RECT 76.400 211.600 77.200 212.400 ;
        RECT 78.000 211.600 78.800 212.400 ;
        RECT 82.800 211.600 83.600 212.400 ;
        RECT 52.400 184.200 53.200 195.800 ;
        RECT 57.200 195.600 58.000 196.400 ;
        RECT 58.800 191.600 59.600 192.400 ;
        RECT 66.800 191.600 67.600 192.400 ;
        RECT 58.800 189.600 59.600 190.400 ;
        RECT 62.000 189.600 62.800 190.400 ;
        RECT 66.800 189.600 67.600 190.400 ;
        RECT 63.600 187.600 64.400 188.400 ;
        RECT 65.200 187.600 66.000 188.400 ;
        RECT 52.400 177.600 53.200 178.400 ;
        RECT 50.800 175.600 51.600 176.400 ;
        RECT 57.200 166.200 58.000 177.800 ;
        RECT 63.700 176.400 64.300 187.600 ;
        RECT 65.300 182.400 65.900 187.600 ;
        RECT 66.900 182.400 67.500 189.600 ;
        RECT 68.500 188.400 69.100 211.600 ;
        RECT 70.000 195.600 70.800 196.400 ;
        RECT 70.100 192.400 70.700 195.600 ;
        RECT 71.700 194.400 72.300 211.600 ;
        RECT 76.500 208.400 77.100 211.600 ;
        RECT 76.400 207.600 77.200 208.400 ;
        RECT 78.100 202.400 78.700 211.600 ;
        RECT 79.600 207.600 80.400 208.400 ;
        RECT 78.000 201.600 78.800 202.400 ;
        RECT 82.900 198.400 83.500 211.600 ;
        RECT 84.400 206.200 85.200 217.800 ;
        RECT 84.400 201.600 85.200 202.400 ;
        RECT 82.800 197.600 83.600 198.400 ;
        RECT 71.600 193.600 72.400 194.400 ;
        RECT 73.200 193.600 74.000 194.400 ;
        RECT 70.000 191.600 70.800 192.400 ;
        RECT 73.300 190.400 73.900 193.600 ;
        RECT 78.000 191.600 78.800 192.400 ;
        RECT 78.100 190.400 78.700 191.600 ;
        RECT 71.600 189.600 72.400 190.400 ;
        RECT 73.200 189.600 74.000 190.400 ;
        RECT 78.000 189.600 78.800 190.400 ;
        RECT 79.600 189.600 80.400 190.400 ;
        RECT 71.700 188.400 72.300 189.600 ;
        RECT 68.400 187.600 69.200 188.400 ;
        RECT 71.600 187.600 72.400 188.400 ;
        RECT 65.200 181.600 66.000 182.400 ;
        RECT 66.800 181.600 67.600 182.400 ;
        RECT 63.600 175.600 64.400 176.400 ;
        RECT 65.200 171.800 66.000 172.600 ;
        RECT 65.300 170.400 65.900 171.800 ;
        RECT 65.200 169.600 66.000 170.400 ;
        RECT 66.800 166.200 67.600 177.800 ;
        RECT 68.500 174.400 69.100 187.600 ;
        RECT 78.100 180.400 78.700 189.600 ;
        RECT 79.700 186.400 80.300 189.600 ;
        RECT 79.600 185.600 80.400 186.400 ;
        RECT 82.800 183.600 83.600 184.400 ;
        RECT 82.900 182.400 83.500 183.600 ;
        RECT 82.800 181.600 83.600 182.400 ;
        RECT 78.000 179.600 78.800 180.400 ;
        RECT 73.200 177.600 74.000 178.400 ;
        RECT 68.400 173.600 69.200 174.400 ;
        RECT 57.200 159.600 58.000 160.400 ;
        RECT 55.600 153.600 56.400 154.400 ;
        RECT 47.700 151.700 49.900 152.300 ;
        RECT 47.700 150.400 48.300 151.700 ;
        RECT 50.800 151.600 51.600 152.400 ;
        RECT 50.900 150.400 51.500 151.600 ;
        RECT 55.700 150.400 56.300 153.600 ;
        RECT 57.300 150.400 57.900 159.600 ;
        RECT 68.500 156.400 69.100 173.600 ;
        RECT 70.000 170.200 70.800 175.800 ;
        RECT 73.300 172.400 73.900 177.600 ;
        RECT 82.900 176.400 83.500 181.600 ;
        RECT 76.400 175.600 77.200 176.400 ;
        RECT 81.200 175.600 82.000 176.400 ;
        RECT 82.800 175.600 83.600 176.400 ;
        RECT 76.500 174.400 77.100 175.600 ;
        RECT 81.300 174.400 81.900 175.600 ;
        RECT 84.500 174.400 85.100 201.600 ;
        RECT 86.100 198.400 86.700 243.600 ;
        RECT 102.000 227.600 102.800 228.400 ;
        RECT 105.200 226.200 106.000 231.800 ;
        RECT 106.800 227.600 107.600 228.400 ;
        RECT 87.600 223.600 88.400 224.400 ;
        RECT 95.600 223.600 96.400 224.400 ;
        RECT 86.000 197.600 86.800 198.400 ;
        RECT 87.700 196.300 88.300 223.600 ;
        RECT 95.700 218.400 96.300 223.600 ;
        RECT 106.900 218.400 107.500 227.600 ;
        RECT 108.400 224.200 109.200 235.800 ;
        RECT 114.800 230.300 115.600 230.400 ;
        RECT 114.800 229.700 117.100 230.300 ;
        RECT 114.800 229.600 115.600 229.700 ;
        RECT 116.500 218.400 117.100 229.700 ;
        RECT 118.000 224.200 118.800 235.800 ;
        RECT 124.400 233.600 125.200 234.400 ;
        RECT 124.500 232.400 125.100 233.600 ;
        RECT 124.400 231.600 125.200 232.400 ;
        RECT 127.600 231.600 128.400 232.400 ;
        RECT 122.800 223.600 123.600 224.400 ;
        RECT 92.400 217.600 93.200 218.400 ;
        RECT 92.500 216.400 93.100 217.600 ;
        RECT 92.400 215.600 93.200 216.400 ;
        RECT 92.400 213.600 93.200 214.400 ;
        RECT 92.500 212.600 93.100 213.600 ;
        RECT 92.400 211.800 93.200 212.600 ;
        RECT 94.000 206.200 94.800 217.800 ;
        RECT 95.600 217.600 96.400 218.400 ;
        RECT 106.800 217.600 107.600 218.400 ;
        RECT 116.400 217.600 117.200 218.400 ;
        RECT 122.900 216.400 123.500 223.600 ;
        RECT 97.200 210.200 98.000 215.800 ;
        RECT 100.400 215.600 101.200 216.400 ;
        RECT 118.000 215.600 118.800 216.400 ;
        RECT 122.800 215.600 123.600 216.400 ;
        RECT 98.800 213.600 99.600 214.400 ;
        RECT 98.900 198.400 99.500 213.600 ;
        RECT 100.500 212.400 101.100 215.600 ;
        RECT 102.000 213.600 102.800 214.400 ;
        RECT 110.000 213.600 110.800 214.400 ;
        RECT 111.600 213.600 112.400 214.400 ;
        RECT 100.400 211.600 101.200 212.400 ;
        RECT 108.400 211.600 109.200 212.400 ;
        RECT 105.200 209.600 106.000 210.400 ;
        RECT 105.300 208.400 105.900 209.600 ;
        RECT 105.200 207.600 106.000 208.400 ;
        RECT 98.800 197.600 99.600 198.400 ;
        RECT 86.100 195.700 88.300 196.300 ;
        RECT 86.100 190.400 86.700 195.700 ;
        RECT 86.000 189.600 86.800 190.400 ;
        RECT 76.400 173.600 77.200 174.400 ;
        RECT 81.200 173.600 82.000 174.400 ;
        RECT 82.800 173.600 83.600 174.400 ;
        RECT 84.400 173.600 85.200 174.400 ;
        RECT 73.200 171.600 74.000 172.400 ;
        RECT 78.000 171.600 78.800 172.400 ;
        RECT 79.600 171.600 80.400 172.400 ;
        RECT 78.100 166.400 78.700 171.600 ;
        RECT 78.000 165.600 78.800 166.400 ;
        RECT 68.400 155.600 69.200 156.400 ;
        RECT 73.200 155.600 74.000 156.400 ;
        RECT 63.600 153.600 64.400 154.400 ;
        RECT 63.700 152.400 64.300 153.600 ;
        RECT 63.600 151.600 64.400 152.400 ;
        RECT 46.000 149.600 46.800 150.400 ;
        RECT 47.600 149.600 48.400 150.400 ;
        RECT 50.800 150.300 51.600 150.400 ;
        RECT 49.300 149.700 51.600 150.300 ;
        RECT 46.100 148.400 46.700 149.600 ;
        RECT 46.000 147.600 46.800 148.400 ;
        RECT 46.100 140.400 46.700 147.600 ;
        RECT 46.000 139.600 46.800 140.400 ;
        RECT 46.000 133.600 46.800 134.400 ;
        RECT 47.700 132.400 48.300 149.600 ;
        RECT 49.300 132.400 49.900 149.700 ;
        RECT 50.800 149.600 51.600 149.700 ;
        RECT 55.600 149.600 56.400 150.400 ;
        RECT 57.200 149.600 58.000 150.400 ;
        RECT 60.400 149.600 61.200 150.400 ;
        RECT 63.600 149.600 64.400 150.400 ;
        RECT 66.800 149.600 67.600 150.400 ;
        RECT 68.400 149.600 69.200 150.400 ;
        RECT 54.000 147.600 54.800 148.400 ;
        RECT 58.800 147.600 59.600 148.400 ;
        RECT 54.100 146.400 54.700 147.600 ;
        RECT 54.000 145.600 54.800 146.400 ;
        RECT 57.200 134.300 58.000 134.400 ;
        RECT 58.900 134.300 59.500 147.600 ;
        RECT 57.200 133.700 59.500 134.300 ;
        RECT 57.200 133.600 58.000 133.700 ;
        RECT 44.400 131.600 45.200 132.400 ;
        RECT 47.600 131.600 48.400 132.400 ;
        RECT 49.200 131.600 50.000 132.400 ;
        RECT 54.000 131.600 54.800 132.400 ;
        RECT 55.600 131.600 56.400 132.400 ;
        RECT 58.800 132.300 59.600 132.400 ;
        RECT 60.500 132.300 61.100 149.600 ;
        RECT 58.800 131.700 61.100 132.300 ;
        RECT 58.800 131.600 59.600 131.700 ;
        RECT 42.900 129.700 45.100 130.300 ;
        RECT 42.800 127.600 43.600 128.400 ;
        RECT 41.200 123.600 42.000 124.400 ;
        RECT 38.000 109.600 38.800 110.400 ;
        RECT 39.600 109.600 40.400 110.400 ;
        RECT 34.800 107.600 35.600 108.400 ;
        RECT 33.200 93.600 34.000 94.400 ;
        RECT 34.800 93.600 35.600 94.400 ;
        RECT 34.900 92.400 35.500 93.600 ;
        RECT 34.800 91.600 35.600 92.400 ;
        RECT 36.400 91.600 37.200 92.400 ;
        RECT 28.400 89.600 29.200 90.400 ;
        RECT 31.600 89.600 32.400 90.400 ;
        RECT 38.100 82.400 38.700 109.600 ;
        RECT 39.700 104.400 40.300 109.600 ;
        RECT 39.600 103.600 40.400 104.400 ;
        RECT 39.600 101.600 40.400 102.400 ;
        RECT 39.700 92.400 40.300 101.600 ;
        RECT 41.300 92.400 41.900 123.600 ;
        RECT 42.900 118.400 43.500 127.600 ;
        RECT 42.800 117.600 43.600 118.400 ;
        RECT 44.500 104.400 45.100 129.700 ;
        RECT 46.000 123.600 46.800 124.400 ;
        RECT 46.100 110.400 46.700 123.600 ;
        RECT 47.700 110.400 48.300 131.600 ;
        RECT 54.100 126.400 54.700 131.600 ;
        RECT 57.200 129.600 58.000 130.400 ;
        RECT 54.000 125.600 54.800 126.400 ;
        RECT 50.800 123.600 51.600 124.400 ;
        RECT 50.900 116.400 51.500 123.600 ;
        RECT 50.800 115.600 51.600 116.400 ;
        RECT 54.100 114.400 54.700 125.600 ;
        RECT 54.000 113.600 54.800 114.400 ;
        RECT 50.800 111.600 51.600 112.400 ;
        RECT 54.000 111.600 54.800 112.400 ;
        RECT 50.900 110.400 51.500 111.600 ;
        RECT 54.100 110.400 54.700 111.600 ;
        RECT 57.300 110.400 57.900 129.600 ;
        RECT 58.900 112.400 59.500 131.600 ;
        RECT 62.000 129.600 62.800 130.400 ;
        RECT 62.100 124.400 62.700 129.600 ;
        RECT 62.000 123.600 62.800 124.400 ;
        RECT 58.800 111.600 59.600 112.400 ;
        RECT 63.700 110.400 64.300 149.600 ;
        RECT 68.500 148.400 69.100 149.600 ;
        RECT 68.400 147.600 69.200 148.400 ;
        RECT 70.000 147.600 70.800 148.400 ;
        RECT 70.100 146.300 70.700 147.600 ;
        RECT 68.500 145.700 70.700 146.300 ;
        RECT 71.600 146.200 72.400 151.800 ;
        RECT 73.300 148.400 73.900 155.600 ;
        RECT 73.200 147.600 74.000 148.400 ;
        RECT 68.500 144.400 69.100 145.700 ;
        RECT 68.400 143.600 69.200 144.400 ;
        RECT 74.800 144.200 75.600 155.800 ;
        RECT 78.100 152.400 78.700 165.600 ;
        RECT 78.000 151.600 78.800 152.400 ;
        RECT 76.400 149.400 77.200 150.400 ;
        RECT 76.400 145.600 77.200 146.400 ;
        RECT 68.500 136.400 69.100 143.600 ;
        RECT 71.600 141.600 72.400 142.400 ;
        RECT 68.400 135.600 69.200 136.400 ;
        RECT 68.500 134.400 69.100 135.600 ;
        RECT 68.400 133.600 69.200 134.400 ;
        RECT 65.200 131.600 66.000 132.400 ;
        RECT 66.800 131.600 67.600 132.400 ;
        RECT 66.900 128.400 67.500 131.600 ;
        RECT 70.000 130.200 70.800 135.800 ;
        RECT 66.800 127.600 67.600 128.400 ;
        RECT 68.400 123.600 69.200 124.400 ;
        RECT 68.500 110.400 69.100 123.600 ;
        RECT 46.000 109.600 46.800 110.400 ;
        RECT 47.600 109.600 48.400 110.400 ;
        RECT 50.800 109.600 51.600 110.400 ;
        RECT 54.000 109.600 54.800 110.400 ;
        RECT 57.200 109.600 58.000 110.400 ;
        RECT 63.600 109.600 64.400 110.400 ;
        RECT 68.400 109.600 69.200 110.400 ;
        RECT 70.000 110.300 70.800 110.400 ;
        RECT 71.700 110.300 72.300 141.600 ;
        RECT 73.200 126.200 74.000 137.800 ;
        RECT 76.500 134.400 77.100 145.600 ;
        RECT 78.000 137.600 78.800 138.400 ;
        RECT 76.400 133.600 77.200 134.400 ;
        RECT 74.800 131.600 75.600 132.600 ;
        RECT 73.200 111.600 74.000 112.400 ;
        RECT 78.100 110.400 78.700 137.600 ;
        RECT 81.300 136.400 81.900 173.600 ;
        RECT 82.900 172.400 83.500 173.600 ;
        RECT 82.800 171.600 83.600 172.400 ;
        RECT 82.800 169.600 83.600 170.400 ;
        RECT 84.500 158.300 85.100 173.600 ;
        RECT 82.900 157.700 85.100 158.300 ;
        RECT 82.900 142.400 83.500 157.700 ;
        RECT 84.400 144.200 85.200 155.800 ;
        RECT 82.800 141.600 83.600 142.400 ;
        RECT 86.100 138.400 86.700 189.600 ;
        RECT 87.600 186.200 88.400 191.800 ;
        RECT 89.200 187.600 90.000 188.400 ;
        RECT 90.800 184.200 91.600 195.800 ;
        RECT 94.000 191.600 94.800 192.400 ;
        RECT 94.100 190.400 94.700 191.600 ;
        RECT 94.000 189.600 94.800 190.400 ;
        RECT 92.400 187.600 93.200 188.400 ;
        RECT 87.600 177.600 88.400 178.400 ;
        RECT 87.700 170.400 88.300 177.600 ;
        RECT 90.800 175.600 91.600 176.400 ;
        RECT 90.900 172.400 91.500 175.600 ;
        RECT 92.500 174.400 93.100 187.600 ;
        RECT 100.400 184.200 101.200 195.800 ;
        RECT 102.000 189.600 102.800 190.400 ;
        RECT 102.100 178.400 102.700 189.600 ;
        RECT 105.300 186.300 105.900 207.600 ;
        RECT 111.700 198.400 112.300 213.600 ;
        RECT 113.200 211.600 114.000 212.400 ;
        RECT 116.400 211.600 117.200 212.400 ;
        RECT 116.500 198.400 117.100 211.600 ;
        RECT 118.100 210.400 118.700 215.600 ;
        RECT 124.400 213.600 125.200 214.400 ;
        RECT 121.200 211.600 122.000 212.400 ;
        RECT 121.300 210.400 121.900 211.600 ;
        RECT 118.000 209.600 118.800 210.400 ;
        RECT 121.200 209.600 122.000 210.400 ;
        RECT 106.800 197.600 107.600 198.400 ;
        RECT 111.600 197.600 112.400 198.400 ;
        RECT 116.400 197.600 117.200 198.400 ;
        RECT 106.900 188.400 107.500 197.600 ;
        RECT 114.800 193.600 115.600 194.400 ;
        RECT 108.400 191.600 109.200 192.400 ;
        RECT 111.600 191.600 112.400 192.400 ;
        RECT 114.900 190.400 115.500 193.600 ;
        RECT 108.400 189.600 109.200 190.400 ;
        RECT 113.200 189.600 114.000 190.400 ;
        RECT 114.800 189.600 115.600 190.400 ;
        RECT 106.800 187.600 107.600 188.400 ;
        RECT 105.300 185.700 107.500 186.300 ;
        RECT 105.200 184.300 106.000 184.400 ;
        RECT 103.700 183.700 106.000 184.300 ;
        RECT 103.700 178.400 104.300 183.700 ;
        RECT 105.200 183.600 106.000 183.700 ;
        RECT 94.000 177.600 94.800 178.400 ;
        RECT 102.000 177.600 102.800 178.400 ;
        RECT 103.600 177.600 104.400 178.400 ;
        RECT 94.100 176.400 94.700 177.600 ;
        RECT 94.000 175.600 94.800 176.400 ;
        RECT 92.400 173.600 93.200 174.400 ;
        RECT 103.700 172.400 104.300 177.600 ;
        RECT 106.900 176.400 107.500 185.700 ;
        RECT 113.300 184.400 113.900 189.600 ;
        RECT 113.200 183.600 114.000 184.400 ;
        RECT 110.000 179.600 110.800 180.400 ;
        RECT 106.800 175.600 107.600 176.400 ;
        RECT 110.100 174.400 110.700 179.600 ;
        RECT 105.200 173.600 106.000 174.400 ;
        RECT 110.000 173.600 110.800 174.400 ;
        RECT 105.300 172.400 105.900 173.600 ;
        RECT 113.300 172.400 113.900 183.600 ;
        RECT 114.800 177.600 115.600 178.400 ;
        RECT 114.900 176.400 115.500 177.600 ;
        RECT 118.100 176.400 118.700 209.600 ;
        RECT 121.200 191.600 122.000 192.400 ;
        RECT 122.800 191.600 123.600 192.400 ;
        RECT 121.300 190.400 121.900 191.600 ;
        RECT 119.600 189.600 120.400 190.400 ;
        RECT 121.200 189.600 122.000 190.400 ;
        RECT 114.800 175.600 115.600 176.400 ;
        RECT 118.000 176.300 118.800 176.400 ;
        RECT 119.700 176.300 120.300 189.600 ;
        RECT 121.200 183.600 122.000 184.400 ;
        RECT 121.300 178.400 121.900 183.600 ;
        RECT 122.900 178.400 123.500 191.600 ;
        RECT 124.500 188.400 125.100 213.600 ;
        RECT 126.000 211.600 126.800 212.400 ;
        RECT 126.100 190.400 126.700 211.600 ;
        RECT 127.700 190.400 128.300 231.600 ;
        RECT 129.300 230.400 129.900 243.600 ;
        RECT 129.200 229.600 130.000 230.400 ;
        RECT 130.800 229.600 131.600 230.400 ;
        RECT 134.000 229.600 134.800 230.400 ;
        RECT 135.700 228.400 136.300 243.600 ;
        RECT 135.600 227.600 136.400 228.400 ;
        RECT 138.800 227.600 139.600 228.400 ;
        RECT 132.400 223.600 133.200 224.400 ;
        RECT 135.600 213.600 136.400 214.400 ;
        RECT 134.000 212.300 134.800 212.400 ;
        RECT 132.500 211.700 134.800 212.300 ;
        RECT 129.200 209.600 130.000 210.400 ;
        RECT 129.300 208.300 129.900 209.600 ;
        RECT 130.800 208.300 131.600 208.400 ;
        RECT 129.300 207.700 131.600 208.300 ;
        RECT 130.800 207.600 131.600 207.700 ;
        RECT 130.900 190.400 131.500 207.600 ;
        RECT 132.500 198.400 133.100 211.700 ;
        RECT 134.000 211.600 134.800 211.700 ;
        RECT 134.000 209.600 134.800 210.400 ;
        RECT 135.700 198.400 136.300 213.600 ;
        RECT 137.200 207.600 138.000 208.400 ;
        RECT 132.400 197.600 133.200 198.400 ;
        RECT 135.600 197.600 136.400 198.400 ;
        RECT 126.000 189.600 126.800 190.400 ;
        RECT 127.600 189.600 128.400 190.400 ;
        RECT 129.200 189.600 130.000 190.400 ;
        RECT 130.800 189.600 131.600 190.400 ;
        RECT 135.600 189.600 136.400 190.400 ;
        RECT 124.400 187.600 125.200 188.400 ;
        RECT 127.600 187.600 128.400 188.400 ;
        RECT 121.200 177.600 122.000 178.400 ;
        RECT 122.800 177.600 123.600 178.400 ;
        RECT 129.300 176.400 129.900 189.600 ;
        RECT 132.400 187.600 133.200 188.400 ;
        RECT 132.500 178.400 133.100 187.600 ;
        RECT 134.000 185.600 134.800 186.400 ;
        RECT 132.400 177.600 133.200 178.400 ;
        RECT 118.000 175.700 120.300 176.300 ;
        RECT 118.000 175.600 118.800 175.700 ;
        RECT 126.000 175.600 126.800 176.400 ;
        RECT 129.200 175.600 130.000 176.400 ;
        RECT 129.300 174.400 129.900 175.600 ;
        RECT 129.200 173.600 130.000 174.400 ;
        RECT 90.800 171.600 91.600 172.400 ;
        RECT 97.200 171.600 98.000 172.400 ;
        RECT 98.800 171.600 99.600 172.400 ;
        RECT 103.600 171.600 104.400 172.400 ;
        RECT 105.200 171.600 106.000 172.400 ;
        RECT 113.200 171.600 114.000 172.400 ;
        RECT 121.200 171.600 122.000 172.400 ;
        RECT 129.200 171.600 130.000 172.400 ;
        RECT 87.600 169.600 88.400 170.400 ;
        RECT 94.000 155.600 94.800 156.400 ;
        RECT 94.100 154.400 94.700 155.600 ;
        RECT 89.200 153.600 90.000 154.400 ;
        RECT 94.000 153.600 94.800 154.400 ;
        RECT 92.400 149.600 93.200 150.400 ;
        RECT 92.500 142.300 93.100 149.600 ;
        RECT 90.900 141.700 93.100 142.300 ;
        RECT 81.200 135.600 82.000 136.400 ;
        RECT 82.800 126.200 83.600 137.800 ;
        RECT 86.000 137.600 86.800 138.400 ;
        RECT 89.200 135.600 90.000 136.400 ;
        RECT 89.300 134.400 89.900 135.600 ;
        RECT 89.200 133.600 90.000 134.400 ;
        RECT 87.600 123.600 88.400 124.400 ;
        RECT 87.700 122.400 88.300 123.600 ;
        RECT 84.400 121.600 85.200 122.400 ;
        RECT 87.600 121.600 88.400 122.400 ;
        RECT 82.800 111.600 83.600 112.400 ;
        RECT 82.900 110.400 83.500 111.600 ;
        RECT 70.000 109.700 72.300 110.300 ;
        RECT 70.000 109.600 70.800 109.700 ;
        RECT 78.000 109.600 78.800 110.400 ;
        RECT 82.800 109.600 83.600 110.400 ;
        RECT 47.600 107.600 48.400 108.400 ;
        RECT 49.200 107.600 50.000 108.400 ;
        RECT 60.400 107.600 61.200 108.400 ;
        RECT 44.400 103.600 45.200 104.400 ;
        RECT 42.800 97.600 43.600 98.400 ;
        RECT 47.700 94.400 48.300 107.600 ;
        RECT 60.500 106.400 61.100 107.600 ;
        RECT 60.400 105.600 61.200 106.400 ;
        RECT 60.500 98.400 61.100 105.600 ;
        RECT 47.600 93.600 48.400 94.400 ;
        RECT 39.600 91.600 40.400 92.400 ;
        RECT 41.200 91.600 42.000 92.400 ;
        RECT 46.000 91.600 46.800 92.400 ;
        RECT 39.700 90.400 40.300 91.600 ;
        RECT 39.600 89.600 40.400 90.400 ;
        RECT 38.000 81.600 38.800 82.400 ;
        RECT 41.300 76.400 41.900 91.600 ;
        RECT 42.800 89.600 43.600 90.400 ;
        RECT 30.000 75.600 30.800 76.400 ;
        RECT 41.200 75.600 42.000 76.400 ;
        RECT 28.400 73.600 29.200 74.400 ;
        RECT 26.800 71.600 27.600 72.400 ;
        RECT 28.500 70.400 29.100 73.600 ;
        RECT 30.100 70.400 30.700 75.600 ;
        RECT 38.000 73.600 38.800 74.400 ;
        RECT 38.100 72.400 38.700 73.600 ;
        RECT 31.600 71.600 32.400 72.400 ;
        RECT 36.400 71.600 37.200 72.400 ;
        RECT 38.000 71.600 38.800 72.400 ;
        RECT 23.600 69.600 24.400 70.400 ;
        RECT 25.200 69.600 26.000 70.400 ;
        RECT 28.400 69.600 29.200 70.400 ;
        RECT 30.000 69.600 30.800 70.400 ;
        RECT 22.000 67.600 22.800 68.400 ;
        RECT 17.200 65.600 18.000 66.400 ;
        RECT 14.000 61.600 14.800 62.400 ;
        RECT 15.600 61.600 16.400 62.400 ;
        RECT 12.400 59.600 13.200 60.400 ;
        RECT 7.600 51.600 8.400 52.400 ;
        RECT 4.400 29.600 5.200 30.400 ;
        RECT 6.000 29.600 6.800 30.400 ;
        RECT 7.700 30.300 8.300 51.600 ;
        RECT 9.200 44.200 10.000 57.800 ;
        RECT 10.800 44.200 11.600 57.800 ;
        RECT 12.400 46.200 13.200 57.800 ;
        RECT 14.100 54.400 14.700 61.600 ;
        RECT 23.700 60.400 24.300 69.600 ;
        RECT 31.700 68.400 32.300 71.600 ;
        RECT 33.200 69.600 34.000 70.400 ;
        RECT 36.500 68.400 37.100 71.600 ;
        RECT 41.200 69.600 42.000 70.400 ;
        RECT 31.600 67.600 32.400 68.400 ;
        RECT 36.400 67.600 37.200 68.400 ;
        RECT 42.800 67.600 43.600 68.400 ;
        RECT 42.900 66.400 43.500 67.600 ;
        RECT 33.200 65.600 34.000 66.400 ;
        RECT 36.400 65.600 37.200 66.400 ;
        RECT 42.800 65.600 43.600 66.400 ;
        RECT 44.400 66.200 45.200 71.800 ;
        RECT 46.100 70.400 46.700 91.600 ;
        RECT 49.200 90.200 50.000 95.800 ;
        RECT 52.400 86.200 53.200 97.800 ;
        RECT 60.400 97.600 61.200 98.400 ;
        RECT 58.800 95.600 59.600 96.400 ;
        RECT 55.600 93.600 56.400 94.400 ;
        RECT 46.000 69.600 46.800 70.400 ;
        RECT 46.000 67.600 46.800 68.400 ;
        RECT 17.200 59.600 18.000 60.400 ;
        RECT 23.600 59.600 24.400 60.400 ;
        RECT 14.000 53.600 14.800 54.400 ;
        RECT 15.600 46.200 16.400 57.800 ;
        RECT 17.300 56.400 17.900 59.600 ;
        RECT 33.300 58.400 33.900 65.600 ;
        RECT 34.800 63.600 35.600 64.400 ;
        RECT 17.200 55.600 18.000 56.400 ;
        RECT 17.300 38.400 17.900 55.600 ;
        RECT 18.800 46.200 19.600 57.800 ;
        RECT 20.400 44.200 21.200 57.800 ;
        RECT 22.000 44.200 22.800 57.800 ;
        RECT 23.600 44.200 24.400 57.800 ;
        RECT 33.200 57.600 34.000 58.400 ;
        RECT 34.900 52.400 35.500 63.600 ;
        RECT 36.500 62.400 37.100 65.600 ;
        RECT 44.400 63.600 45.200 64.400 ;
        RECT 36.400 61.600 37.200 62.400 ;
        RECT 36.500 54.400 37.100 61.600 ;
        RECT 44.500 58.400 45.100 63.600 ;
        RECT 44.400 57.600 45.200 58.400 ;
        RECT 46.100 54.400 46.700 67.600 ;
        RECT 47.600 64.200 48.400 75.800 ;
        RECT 49.200 71.600 50.000 72.400 ;
        RECT 49.300 70.200 49.900 71.600 ;
        RECT 55.700 70.400 56.300 93.600 ;
        RECT 58.900 92.400 59.500 95.600 ;
        RECT 58.800 91.600 59.600 92.400 ;
        RECT 62.000 86.200 62.800 97.800 ;
        RECT 63.700 94.400 64.300 109.600 ;
        RECT 68.400 95.600 69.200 96.400 ;
        RECT 63.600 93.600 64.400 94.400 ;
        RECT 62.000 83.600 62.800 84.400 ;
        RECT 49.200 69.400 50.000 70.200 ;
        RECT 52.400 69.600 53.200 70.400 ;
        RECT 55.600 69.600 56.400 70.400 ;
        RECT 49.200 65.600 50.000 66.400 ;
        RECT 49.300 58.400 49.900 65.600 ;
        RECT 49.200 57.600 50.000 58.400 ;
        RECT 49.300 56.400 49.900 57.600 ;
        RECT 49.200 55.600 50.000 56.400 ;
        RECT 36.400 53.600 37.200 54.400 ;
        RECT 46.000 53.600 46.800 54.400 ;
        RECT 34.800 51.600 35.600 52.400 ;
        RECT 9.200 30.300 10.000 30.400 ;
        RECT 7.700 29.700 10.000 30.300 ;
        RECT 4.500 12.400 5.100 29.600 ;
        RECT 7.700 12.400 8.300 29.700 ;
        RECT 9.200 29.600 10.000 29.700 ;
        RECT 14.000 24.200 14.800 37.800 ;
        RECT 15.600 24.200 16.400 37.800 ;
        RECT 17.200 37.600 18.000 38.400 ;
        RECT 22.000 37.600 22.800 38.400 ;
        RECT 17.200 24.200 18.000 35.800 ;
        RECT 18.800 27.600 19.600 28.400 ;
        RECT 20.400 24.200 21.200 35.800 ;
        RECT 22.100 26.400 22.700 37.600 ;
        RECT 22.000 25.600 22.800 26.400 ;
        RECT 22.100 20.400 22.700 25.600 ;
        RECT 23.600 24.200 24.400 35.800 ;
        RECT 25.200 24.200 26.000 37.800 ;
        RECT 26.800 24.200 27.600 37.800 ;
        RECT 28.400 24.200 29.200 37.800 ;
        RECT 30.000 29.600 30.800 30.400 ;
        RECT 30.100 22.400 30.700 29.600 ;
        RECT 30.000 21.600 30.800 22.400 ;
        RECT 17.200 19.600 18.000 20.400 ;
        RECT 22.000 19.600 22.800 20.400 ;
        RECT 4.400 11.600 5.200 12.400 ;
        RECT 7.600 11.600 8.400 12.400 ;
        RECT 9.200 4.200 10.000 17.800 ;
        RECT 10.800 4.200 11.600 17.800 ;
        RECT 12.400 6.200 13.200 17.800 ;
        RECT 14.000 13.600 14.800 14.400 ;
        RECT 15.600 6.200 16.400 17.800 ;
        RECT 17.300 16.400 17.900 19.600 ;
        RECT 17.200 15.600 18.000 16.400 ;
        RECT 18.800 6.200 19.600 17.800 ;
        RECT 20.400 4.200 21.200 17.800 ;
        RECT 22.000 4.200 22.800 17.800 ;
        RECT 23.600 4.200 24.400 17.800 ;
        RECT 33.200 15.600 34.000 16.400 ;
        RECT 34.900 12.400 35.500 51.600 ;
        RECT 36.500 18.400 37.100 53.600 ;
        RECT 41.200 50.300 42.000 50.400 ;
        RECT 39.700 49.700 42.000 50.300 ;
        RECT 38.000 43.600 38.800 44.400 ;
        RECT 38.100 40.400 38.700 43.600 ;
        RECT 38.000 39.600 38.800 40.400 ;
        RECT 38.000 38.300 38.800 38.400 ;
        RECT 39.700 38.300 40.300 49.700 ;
        RECT 41.200 49.600 42.000 49.700 ;
        RECT 42.800 47.600 43.600 48.400 ;
        RECT 41.200 39.600 42.000 40.400 ;
        RECT 38.000 37.700 40.300 38.300 ;
        RECT 38.000 37.600 38.800 37.700 ;
        RECT 41.300 32.400 41.900 39.600 ;
        RECT 41.200 31.600 42.000 32.400 ;
        RECT 39.600 27.600 40.400 28.400 ;
        RECT 36.400 17.600 37.200 18.400 ;
        RECT 36.500 14.400 37.100 17.600 ;
        RECT 41.200 16.300 42.000 16.400 ;
        RECT 42.900 16.300 43.500 47.600 ;
        RECT 52.500 30.400 53.100 69.600 ;
        RECT 57.200 64.200 58.000 75.800 ;
        RECT 62.100 74.400 62.700 83.600 ;
        RECT 63.700 74.400 64.300 93.600 ;
        RECT 66.800 89.600 67.600 90.400 ;
        RECT 68.400 89.600 69.200 90.400 ;
        RECT 66.900 88.400 67.500 89.600 ;
        RECT 68.500 88.400 69.100 89.600 ;
        RECT 65.200 87.600 66.000 88.400 ;
        RECT 66.800 87.600 67.600 88.400 ;
        RECT 68.400 87.600 69.200 88.400 ;
        RECT 65.300 78.400 65.900 87.600 ;
        RECT 65.200 77.600 66.000 78.400 ;
        RECT 62.000 73.600 62.800 74.400 ;
        RECT 63.600 73.600 64.400 74.400 ;
        RECT 66.900 72.300 67.500 87.600 ;
        RECT 70.100 72.400 70.700 109.600 ;
        RECT 73.200 97.600 74.000 98.400 ;
        RECT 71.600 95.600 72.400 96.400 ;
        RECT 71.700 92.400 72.300 95.600 ;
        RECT 73.300 94.400 73.900 97.600 ;
        RECT 73.200 93.600 74.000 94.400 ;
        RECT 71.600 91.600 72.400 92.400 ;
        RECT 74.800 91.600 75.600 92.400 ;
        RECT 76.400 91.600 77.200 92.400 ;
        RECT 76.500 90.400 77.100 91.600 ;
        RECT 76.400 89.600 77.200 90.400 ;
        RECT 73.200 85.600 74.000 86.400 ;
        RECT 68.400 72.300 69.200 72.400 ;
        RECT 66.900 71.700 69.200 72.300 ;
        RECT 68.400 71.600 69.200 71.700 ;
        RECT 70.000 71.600 70.800 72.400 ;
        RECT 65.200 69.600 66.000 70.400 ;
        RECT 71.600 69.600 72.400 70.400 ;
        RECT 63.600 67.600 64.400 68.400 ;
        RECT 70.000 67.600 70.800 68.400 ;
        RECT 71.600 67.600 72.400 68.400 ;
        RECT 63.700 66.400 64.300 67.600 ;
        RECT 70.100 66.400 70.700 67.600 ;
        RECT 63.600 65.600 64.400 66.400 ;
        RECT 70.000 65.600 70.800 66.400 ;
        RECT 68.400 63.600 69.200 64.400 ;
        RECT 63.600 59.600 64.400 60.400 ;
        RECT 60.400 55.600 61.200 56.400 ;
        RECT 60.500 54.400 61.100 55.600 ;
        RECT 60.400 53.600 61.200 54.400 ;
        RECT 63.700 52.400 64.300 59.600 ;
        RECT 68.500 52.400 69.100 63.600 ;
        RECT 71.700 52.400 72.300 67.600 ;
        RECT 73.300 58.400 73.900 85.600 ;
        RECT 78.100 82.400 78.700 109.600 ;
        RECT 84.500 108.400 85.100 121.600 ;
        RECT 87.600 115.600 88.400 116.400 ;
        RECT 86.000 113.600 86.800 114.400 ;
        RECT 87.700 112.400 88.300 115.600 ;
        RECT 87.600 111.600 88.400 112.400 ;
        RECT 89.200 111.600 90.000 112.400 ;
        RECT 84.400 107.600 85.200 108.400 ;
        RECT 79.600 103.600 80.400 104.400 ;
        RECT 79.700 98.400 80.300 103.600 ;
        RECT 89.300 102.400 89.900 111.600 ;
        RECT 90.900 110.400 91.500 141.700 ;
        RECT 94.100 134.300 94.700 153.600 ;
        RECT 95.600 151.600 96.400 152.400 ;
        RECT 97.300 148.400 97.900 171.600 ;
        RECT 98.900 166.400 99.500 171.600 ;
        RECT 121.300 170.400 121.900 171.600 ;
        RECT 113.200 169.600 114.000 170.400 ;
        RECT 121.200 169.600 122.000 170.400 ;
        RECT 110.000 167.600 110.800 168.400 ;
        RECT 98.800 165.600 99.600 166.400 ;
        RECT 106.800 165.600 107.600 166.400 ;
        RECT 103.600 157.600 104.400 158.400 ;
        RECT 103.700 152.400 104.300 157.600 ;
        RECT 106.900 156.400 107.500 165.600 ;
        RECT 106.800 155.600 107.600 156.400 ;
        RECT 106.900 154.400 107.500 155.600 ;
        RECT 106.800 153.600 107.600 154.400 ;
        RECT 102.000 151.600 102.800 152.400 ;
        RECT 103.600 151.600 104.400 152.400 ;
        RECT 108.400 151.600 109.200 152.400 ;
        RECT 98.800 149.600 99.600 150.400 ;
        RECT 105.200 149.600 106.000 150.400 ;
        RECT 97.200 147.600 98.000 148.400 ;
        RECT 98.900 146.400 99.500 149.600 ;
        RECT 110.100 148.400 110.700 167.600 ;
        RECT 111.600 163.600 112.400 164.400 ;
        RECT 111.700 156.400 112.300 163.600 ;
        RECT 111.600 155.600 112.400 156.400 ;
        RECT 111.600 153.600 112.400 154.400 ;
        RECT 111.600 149.600 112.400 150.400 ;
        RECT 111.700 148.400 112.300 149.600 ;
        RECT 110.000 147.600 110.800 148.400 ;
        RECT 111.600 147.600 112.400 148.400 ;
        RECT 98.800 145.600 99.600 146.400 ;
        RECT 95.600 137.600 96.400 138.400 ;
        RECT 92.500 133.700 94.700 134.300 ;
        RECT 92.500 114.400 93.100 133.700 ;
        RECT 98.900 132.400 99.500 145.600 ;
        RECT 102.000 143.600 102.800 144.400 ;
        RECT 100.400 133.600 101.200 134.400 ;
        RECT 100.500 132.400 101.100 133.600 ;
        RECT 94.000 131.600 94.800 132.400 ;
        RECT 98.800 131.600 99.600 132.400 ;
        RECT 100.400 131.600 101.200 132.400 ;
        RECT 95.600 130.300 96.400 130.400 ;
        RECT 94.100 129.700 96.400 130.300 ;
        RECT 94.100 118.400 94.700 129.700 ;
        RECT 95.600 129.600 96.400 129.700 ;
        RECT 98.900 122.400 99.500 131.600 ;
        RECT 102.000 130.200 102.800 135.800 ;
        RECT 103.600 133.600 104.400 134.400 ;
        RECT 105.200 126.200 106.000 137.800 ;
        RECT 106.800 131.800 107.600 132.600 ;
        RECT 106.900 130.400 107.500 131.800 ;
        RECT 110.000 131.600 110.800 132.400 ;
        RECT 106.800 129.600 107.600 130.400 ;
        RECT 98.800 121.600 99.600 122.400 ;
        RECT 103.600 121.600 104.400 122.400 ;
        RECT 103.700 118.400 104.300 121.600 ;
        RECT 94.000 117.600 94.800 118.400 ;
        RECT 103.600 117.600 104.400 118.400 ;
        RECT 92.400 114.300 93.200 114.400 ;
        RECT 92.400 113.700 94.700 114.300 ;
        RECT 92.400 113.600 93.200 113.700 ;
        RECT 90.800 109.600 91.600 110.400 ;
        RECT 89.200 101.600 90.000 102.400 ;
        RECT 79.600 98.300 80.400 98.400 ;
        RECT 79.600 97.700 81.900 98.300 ;
        RECT 79.600 97.600 80.400 97.700 ;
        RECT 79.600 95.600 80.400 96.400 ;
        RECT 78.000 81.600 78.800 82.400 ;
        RECT 78.000 73.600 78.800 74.400 ;
        RECT 79.600 73.600 80.400 74.400 ;
        RECT 74.800 71.600 75.600 72.400 ;
        RECT 74.900 68.400 75.500 71.600 ;
        RECT 74.800 67.600 75.600 68.400 ;
        RECT 74.800 61.600 75.600 62.400 ;
        RECT 73.200 57.600 74.000 58.400 ;
        RECT 74.900 54.400 75.500 61.600 ;
        RECT 74.800 53.600 75.600 54.400 ;
        RECT 76.400 53.600 77.200 54.400 ;
        RECT 76.500 52.400 77.100 53.600 ;
        RECT 78.100 52.400 78.700 73.600 ;
        RECT 79.600 69.600 80.400 70.400 ;
        RECT 79.700 66.400 80.300 69.600 ;
        RECT 81.300 68.400 81.900 97.700 ;
        RECT 90.900 96.300 91.500 109.600 ;
        RECT 92.400 96.300 93.200 96.400 ;
        RECT 90.900 95.700 93.200 96.300 ;
        RECT 92.400 95.600 93.200 95.700 ;
        RECT 82.800 93.600 83.600 94.400 ;
        RECT 89.200 93.600 90.000 94.400 ;
        RECT 82.900 72.400 83.500 93.600 ;
        RECT 87.600 91.600 88.400 92.400 ;
        RECT 84.400 89.600 85.200 90.400 ;
        RECT 84.500 86.400 85.100 89.600 ;
        RECT 84.400 85.600 85.200 86.400 ;
        RECT 87.600 83.600 88.400 84.400 ;
        RECT 82.800 71.600 83.600 72.400 ;
        RECT 82.900 70.400 83.500 71.600 ;
        RECT 82.800 69.600 83.600 70.400 ;
        RECT 84.400 69.600 85.200 70.400 ;
        RECT 81.200 67.600 82.000 68.400 ;
        RECT 79.600 65.600 80.400 66.400 ;
        RECT 82.900 54.400 83.500 69.600 ;
        RECT 84.500 60.400 85.100 69.600 ;
        RECT 86.000 65.600 86.800 66.400 ;
        RECT 84.400 59.600 85.200 60.400 ;
        RECT 82.800 53.600 83.600 54.400 ;
        RECT 86.000 53.600 86.800 54.400 ;
        RECT 86.100 52.400 86.700 53.600 ;
        RECT 87.700 52.400 88.300 83.600 ;
        RECT 89.300 62.400 89.900 93.600 ;
        RECT 92.500 92.400 93.100 95.600 ;
        RECT 92.400 91.600 93.200 92.400 ;
        RECT 94.100 90.400 94.700 113.700 ;
        RECT 95.600 113.600 96.400 114.400 ;
        RECT 106.800 113.600 107.600 114.400 ;
        RECT 95.700 112.400 96.300 113.600 ;
        RECT 106.900 112.400 107.500 113.600 ;
        RECT 95.600 111.600 96.400 112.400 ;
        RECT 98.800 112.300 99.600 112.400 ;
        RECT 98.800 111.700 101.100 112.300 ;
        RECT 98.800 111.600 99.600 111.700 ;
        RECT 100.500 110.400 101.100 111.700 ;
        RECT 106.800 111.600 107.600 112.400 ;
        RECT 110.100 110.400 110.700 131.600 ;
        RECT 113.300 130.400 113.900 169.600 ;
        RECT 116.400 163.600 117.200 164.400 ;
        RECT 119.600 163.600 120.400 164.400 ;
        RECT 116.500 156.400 117.100 163.600 ;
        RECT 114.800 155.600 115.600 156.400 ;
        RECT 116.400 155.600 117.200 156.400 ;
        RECT 114.900 152.400 115.500 155.600 ;
        RECT 114.800 151.600 115.600 152.400 ;
        RECT 116.400 151.600 117.200 152.400 ;
        RECT 119.700 152.300 120.300 163.600 ;
        RECT 134.100 156.400 134.700 185.600 ;
        RECT 137.300 176.400 137.900 207.600 ;
        RECT 138.900 190.400 139.500 227.600 ;
        RECT 143.700 226.400 144.300 283.600 ;
        RECT 164.500 278.400 165.100 291.600 ;
        RECT 164.400 277.600 165.200 278.400 ;
        RECT 164.400 271.600 165.200 272.400 ;
        RECT 164.500 270.400 165.100 271.600 ;
        RECT 153.200 269.600 154.000 270.400 ;
        RECT 162.800 269.600 163.600 270.400 ;
        RECT 164.400 269.600 165.200 270.400 ;
        RECT 150.000 263.600 150.800 264.400 ;
        RECT 153.300 252.400 153.900 269.600 ;
        RECT 162.900 268.400 163.500 269.600 ;
        RECT 162.800 267.600 163.600 268.400 ;
        RECT 166.100 260.400 166.700 291.600 ;
        RECT 169.200 289.600 170.000 290.400 ;
        RECT 175.700 288.400 176.300 291.600 ;
        RECT 175.600 287.600 176.400 288.400 ;
        RECT 174.000 275.600 174.800 276.400 ;
        RECT 169.200 271.600 170.000 272.400 ;
        RECT 167.600 265.600 168.400 266.400 ;
        RECT 169.300 262.400 169.900 271.600 ;
        RECT 174.100 266.400 174.700 275.600 ;
        RECT 175.700 270.400 176.300 287.600 ;
        RECT 178.800 284.200 179.600 297.800 ;
        RECT 180.400 284.200 181.200 297.800 ;
        RECT 182.000 286.200 182.800 297.800 ;
        RECT 183.600 293.600 184.400 294.400 ;
        RECT 185.200 286.200 186.000 297.800 ;
        RECT 186.900 296.400 187.500 303.600 ;
        RECT 186.800 295.600 187.600 296.400 ;
        RECT 186.900 282.400 187.500 295.600 ;
        RECT 188.400 286.200 189.200 297.800 ;
        RECT 190.000 284.200 190.800 297.800 ;
        RECT 191.600 284.200 192.400 297.800 ;
        RECT 193.200 284.200 194.000 297.800 ;
        RECT 186.800 281.600 187.600 282.400 ;
        RECT 191.600 281.600 192.400 282.400 ;
        RECT 175.600 269.600 176.400 270.400 ;
        RECT 178.800 269.600 179.600 270.400 ;
        RECT 174.000 265.600 174.800 266.400 ;
        RECT 169.200 261.600 170.000 262.400 ;
        RECT 166.000 259.600 166.800 260.400 ;
        RECT 153.200 251.600 154.000 252.400 ;
        RECT 145.200 243.600 146.000 244.400 ;
        RECT 154.800 244.200 155.600 257.800 ;
        RECT 156.400 244.200 157.200 257.800 ;
        RECT 158.000 244.200 158.800 257.800 ;
        RECT 159.600 246.200 160.400 257.800 ;
        RECT 161.200 255.600 162.000 256.400 ;
        RECT 162.800 246.200 163.600 257.800 ;
        RECT 164.400 253.600 165.200 254.400 ;
        RECT 166.000 246.200 166.800 257.800 ;
        RECT 167.600 244.200 168.400 257.800 ;
        RECT 169.200 244.200 170.000 257.800 ;
        RECT 174.000 252.300 174.800 252.400 ;
        RECT 175.700 252.300 176.300 269.600 ;
        RECT 183.600 264.200 184.400 277.800 ;
        RECT 185.200 264.200 186.000 277.800 ;
        RECT 186.800 264.200 187.600 275.800 ;
        RECT 188.400 267.600 189.200 268.400 ;
        RECT 188.400 265.600 189.200 266.400 ;
        RECT 188.500 262.400 189.100 265.600 ;
        RECT 190.000 264.200 190.800 275.800 ;
        RECT 191.700 266.400 192.300 281.600 ;
        RECT 194.900 280.400 195.500 311.600 ;
        RECT 204.500 310.400 205.100 311.600 ;
        RECT 196.400 309.600 197.200 310.400 ;
        RECT 204.400 309.600 205.200 310.400 ;
        RECT 207.600 305.600 208.400 306.400 ;
        RECT 196.400 303.600 197.200 304.400 ;
        RECT 196.500 290.400 197.100 303.600 ;
        RECT 207.700 298.400 208.300 305.600 ;
        RECT 209.200 304.200 210.000 317.800 ;
        RECT 210.800 304.200 211.600 317.800 ;
        RECT 212.400 304.200 213.200 315.800 ;
        RECT 214.000 307.600 214.800 308.400 ;
        RECT 214.100 306.400 214.700 307.600 ;
        RECT 214.000 305.600 214.800 306.400 ;
        RECT 215.600 304.200 216.400 315.800 ;
        RECT 217.300 306.400 217.900 321.600 ;
        RECT 236.500 318.400 237.100 345.600 ;
        RECT 242.800 344.200 243.600 357.800 ;
        RECT 244.400 344.200 245.200 357.800 ;
        RECT 246.000 344.200 246.800 355.800 ;
        RECT 247.600 347.600 248.400 348.400 ;
        RECT 249.200 344.200 250.000 355.800 ;
        RECT 250.900 346.400 251.500 375.600 ;
        RECT 252.400 366.200 253.200 377.800 ;
        RECT 254.100 374.400 254.700 379.700 ;
        RECT 254.000 373.600 254.800 374.400 ;
        RECT 255.600 366.200 256.400 377.800 ;
        RECT 257.200 364.200 258.000 377.800 ;
        RECT 258.800 364.200 259.600 377.800 ;
        RECT 260.500 374.400 261.100 383.600 ;
        RECT 260.400 373.600 261.200 374.400 ;
        RECT 266.900 372.400 267.500 389.600 ;
        RECT 273.200 384.200 274.000 397.800 ;
        RECT 274.800 384.200 275.600 397.800 ;
        RECT 276.400 384.200 277.200 395.800 ;
        RECT 278.100 388.400 278.700 409.600 ;
        RECT 282.800 407.600 283.600 408.400 ;
        RECT 282.900 398.400 283.500 407.600 ;
        RECT 282.800 397.600 283.600 398.400 ;
        RECT 278.000 387.600 278.800 388.400 ;
        RECT 279.600 384.200 280.400 395.800 ;
        RECT 281.200 385.600 282.000 386.400 ;
        RECT 281.300 380.400 281.900 385.600 ;
        RECT 282.800 384.200 283.600 395.800 ;
        RECT 284.400 384.200 285.200 397.800 ;
        RECT 286.000 384.200 286.800 397.800 ;
        RECT 287.600 384.200 288.400 397.800 ;
        RECT 289.300 390.400 289.900 415.600 ;
        RECT 294.100 410.400 294.700 419.600 ;
        RECT 295.700 416.400 296.300 429.600 ;
        RECT 297.200 424.200 298.000 437.800 ;
        RECT 298.800 424.200 299.600 437.800 ;
        RECT 300.400 424.200 301.200 437.800 ;
        RECT 302.000 424.200 302.800 435.800 ;
        RECT 303.600 425.600 304.400 426.400 ;
        RECT 305.200 424.200 306.000 435.800 ;
        RECT 306.800 427.600 307.600 428.400 ;
        RECT 308.400 424.200 309.200 435.800 ;
        RECT 310.000 424.200 310.800 437.800 ;
        RECT 311.600 424.200 312.400 437.800 ;
        RECT 313.300 426.400 313.900 455.600 ;
        RECT 314.800 446.200 315.600 457.800 ;
        RECT 316.400 453.600 317.200 454.400 ;
        RECT 318.000 446.200 318.800 457.800 ;
        RECT 319.600 444.200 320.400 457.800 ;
        RECT 321.200 444.200 322.000 457.800 ;
        RECT 327.700 438.400 328.300 467.600 ;
        RECT 335.700 464.400 336.300 467.600 ;
        RECT 335.600 463.600 336.400 464.400 ;
        RECT 340.400 463.600 341.200 464.400 ;
        RECT 340.500 462.400 341.100 463.600 ;
        RECT 340.400 461.600 341.200 462.400 ;
        RECT 330.800 449.600 331.600 450.400 ;
        RECT 330.900 448.400 331.500 449.600 ;
        RECT 330.800 447.600 331.600 448.400 ;
        RECT 335.600 446.200 336.400 457.800 ;
        RECT 342.100 456.400 342.700 489.600 ;
        RECT 345.200 487.600 346.000 488.400 ;
        RECT 343.600 483.600 344.400 484.400 ;
        RECT 343.700 456.400 344.300 483.600 ;
        RECT 346.900 470.400 347.500 491.700 ;
        RECT 348.400 491.600 349.200 492.400 ;
        RECT 351.600 491.600 352.400 492.400 ;
        RECT 354.800 491.600 355.600 492.400 ;
        RECT 356.400 491.600 357.200 492.400 ;
        RECT 346.800 469.600 347.600 470.400 ;
        RECT 345.200 467.600 346.000 468.400 ;
        RECT 342.000 455.600 342.800 456.400 ;
        RECT 343.600 455.600 344.400 456.400 ;
        RECT 343.600 451.600 344.400 452.600 ;
        RECT 345.200 446.200 346.000 457.800 ;
        RECT 327.600 437.600 328.400 438.400 ;
        RECT 346.900 436.400 347.500 469.600 ;
        RECT 348.500 464.400 349.100 491.600 ;
        RECT 354.900 488.400 355.500 491.600 ;
        RECT 356.500 490.400 357.100 491.600 ;
        RECT 356.400 489.600 357.200 490.400 ;
        RECT 354.800 487.600 355.600 488.400 ;
        RECT 356.400 479.600 357.200 480.400 ;
        RECT 354.800 475.600 355.600 476.400 ;
        RECT 354.800 473.600 355.600 474.400 ;
        RECT 350.000 471.600 350.800 472.400 ;
        RECT 354.900 470.400 355.500 473.600 ;
        RECT 356.500 470.400 357.100 479.600 ;
        RECT 354.800 469.600 355.600 470.400 ;
        RECT 356.400 469.600 357.200 470.400 ;
        RECT 348.400 463.600 349.200 464.400 ;
        RECT 353.200 461.600 354.000 462.400 ;
        RECT 348.400 450.200 349.200 455.800 ;
        RECT 350.000 455.600 350.800 456.400 ;
        RECT 353.300 452.400 353.900 461.600 ;
        RECT 353.200 451.600 354.000 452.400 ;
        RECT 351.600 447.600 352.400 448.400 ;
        RECT 348.400 443.600 349.200 444.400 ;
        RECT 313.200 425.600 314.000 426.400 ;
        RECT 316.400 425.600 317.200 426.400 ;
        RECT 326.000 425.600 326.800 426.400 ;
        RECT 329.200 426.200 330.000 431.800 ;
        RECT 295.600 415.600 296.400 416.400 ;
        RECT 303.600 415.600 304.400 416.400 ;
        RECT 298.800 413.600 299.600 414.400 ;
        RECT 303.700 412.400 304.300 415.600 ;
        RECT 300.400 411.600 301.200 412.400 ;
        RECT 303.600 411.600 304.400 412.400 ;
        RECT 294.000 409.600 294.800 410.400 ;
        RECT 290.800 407.600 291.600 408.400 ;
        RECT 297.200 397.600 298.000 398.400 ;
        RECT 289.200 389.600 290.000 390.400 ;
        RECT 284.400 381.600 285.200 382.400 ;
        RECT 281.200 379.600 282.000 380.400 ;
        RECT 281.200 377.600 282.000 378.400 ;
        RECT 270.000 373.600 270.800 374.400 ;
        RECT 274.800 373.600 275.600 374.400 ;
        RECT 263.600 371.600 264.400 372.400 ;
        RECT 266.800 371.600 267.600 372.400 ;
        RECT 270.000 369.600 270.800 370.400 ;
        RECT 250.800 345.600 251.600 346.400 ;
        RECT 238.000 341.600 238.800 342.400 ;
        RECT 238.100 336.400 238.700 341.600 ;
        RECT 250.900 340.400 251.500 345.600 ;
        RECT 252.400 344.200 253.200 355.800 ;
        RECT 254.000 344.200 254.800 357.800 ;
        RECT 255.600 344.200 256.400 357.800 ;
        RECT 257.200 344.200 258.000 357.800 ;
        RECT 266.800 357.600 267.600 358.400 ;
        RECT 258.800 351.600 259.600 352.400 ;
        RECT 258.900 350.400 259.500 351.600 ;
        RECT 270.100 350.400 270.700 369.600 ;
        RECT 281.300 358.400 281.900 377.600 ;
        RECT 284.500 358.400 285.100 381.600 ;
        RECT 286.000 379.600 286.800 380.400 ;
        RECT 286.100 378.400 286.700 379.600 ;
        RECT 300.500 378.400 301.100 411.600 ;
        RECT 308.400 404.200 309.200 417.800 ;
        RECT 310.000 404.200 310.800 417.800 ;
        RECT 311.600 406.200 312.400 417.800 ;
        RECT 313.200 413.600 314.000 414.400 ;
        RECT 314.800 406.200 315.600 417.800 ;
        RECT 316.500 416.400 317.100 425.600 ;
        RECT 316.400 415.600 317.200 416.400 ;
        RECT 316.500 412.400 317.100 415.600 ;
        RECT 316.400 411.600 317.200 412.400 ;
        RECT 318.000 406.200 318.800 417.800 ;
        RECT 319.600 404.200 320.400 417.800 ;
        RECT 321.200 404.200 322.000 417.800 ;
        RECT 322.800 404.200 323.600 417.800 ;
        RECT 326.100 400.400 326.700 425.600 ;
        RECT 332.400 424.200 333.200 435.800 ;
        RECT 335.600 429.600 336.400 430.400 ;
        RECT 337.200 427.600 338.000 428.400 ;
        RECT 335.600 410.200 336.400 415.800 ;
        RECT 337.300 414.400 337.900 427.600 ;
        RECT 342.000 424.200 342.800 435.800 ;
        RECT 346.800 435.600 347.600 436.400 ;
        RECT 346.800 433.600 347.600 434.400 ;
        RECT 346.900 432.400 347.500 433.600 ;
        RECT 346.800 431.600 347.600 432.400 ;
        RECT 348.500 430.400 349.100 443.600 ;
        RECT 356.500 438.400 357.100 469.600 ;
        RECT 358.100 468.400 358.700 493.600 ;
        RECT 359.600 491.600 360.400 492.400 ;
        RECT 367.600 491.600 368.400 492.400 ;
        RECT 370.800 491.600 371.600 492.400 ;
        RECT 364.400 489.600 365.200 490.400 ;
        RECT 364.500 488.400 365.100 489.600 ;
        RECT 364.400 487.600 365.200 488.400 ;
        RECT 359.600 483.600 360.400 484.400 ;
        RECT 359.700 470.400 360.300 483.600 ;
        RECT 364.500 476.400 365.100 487.600 ;
        RECT 366.000 477.600 366.800 478.400 ;
        RECT 364.400 475.600 365.200 476.400 ;
        RECT 361.200 473.600 362.000 474.400 ;
        RECT 364.400 471.600 365.200 472.400 ;
        RECT 364.500 470.400 365.100 471.600 ;
        RECT 366.100 470.400 366.700 477.600 ;
        RECT 367.700 474.400 368.300 491.600 ;
        RECT 370.900 480.400 371.500 491.600 ;
        RECT 372.500 484.400 373.100 513.600 ;
        RECT 375.700 512.400 376.300 513.600 ;
        RECT 375.600 511.600 376.400 512.400 ;
        RECT 378.800 511.600 379.600 512.400 ;
        RECT 391.600 511.600 392.400 512.400 ;
        RECT 398.000 511.600 398.800 512.400 ;
        RECT 378.900 510.400 379.500 511.600 ;
        RECT 391.700 510.400 392.300 511.600 ;
        RECT 409.300 510.400 409.900 513.600 ;
        RECT 410.800 511.600 411.600 512.400 ;
        RECT 377.200 510.300 378.000 510.400 ;
        RECT 375.700 509.700 378.000 510.300 ;
        RECT 374.000 491.600 374.800 492.400 ;
        RECT 372.400 483.600 373.200 484.400 ;
        RECT 370.800 479.600 371.600 480.400 ;
        RECT 367.600 473.600 368.400 474.400 ;
        RECT 359.600 469.600 360.400 470.400 ;
        RECT 364.400 469.600 365.200 470.400 ;
        RECT 366.000 469.600 366.800 470.400 ;
        RECT 358.000 467.600 358.800 468.400 ;
        RECT 364.500 466.400 365.100 469.600 ;
        RECT 364.400 465.600 365.200 466.400 ;
        RECT 364.400 455.600 365.200 456.400 ;
        RECT 358.000 453.600 358.800 454.400 ;
        RECT 361.200 453.600 362.000 454.400 ;
        RECT 350.000 437.600 350.800 438.400 ;
        RECT 356.400 437.600 357.200 438.400 ;
        RECT 350.100 430.400 350.700 437.600 ;
        RECT 356.400 435.600 357.200 436.400 ;
        RECT 354.800 431.600 355.600 432.400 ;
        RECT 354.900 430.400 355.500 431.600 ;
        RECT 348.400 429.600 349.200 430.400 ;
        RECT 350.000 429.600 350.800 430.400 ;
        RECT 354.800 429.600 355.600 430.400 ;
        RECT 354.800 427.600 355.600 428.400 ;
        RECT 337.200 413.600 338.000 414.400 ;
        RECT 337.300 412.400 337.900 413.600 ;
        RECT 337.200 411.600 338.000 412.400 ;
        RECT 332.400 407.600 333.200 408.400 ;
        RECT 338.800 406.200 339.600 417.800 ;
        RECT 342.000 415.600 342.800 416.400 ;
        RECT 342.100 412.400 342.700 415.600 ;
        RECT 342.000 411.600 342.800 412.400 ;
        RECT 348.400 406.200 349.200 417.800 ;
        RECT 353.200 417.600 354.000 418.400 ;
        RECT 353.300 410.400 353.900 417.600 ;
        RECT 354.900 414.400 355.500 427.600 ;
        RECT 354.800 413.600 355.600 414.400 ;
        RECT 356.500 412.400 357.100 435.600 ;
        RECT 358.100 428.400 358.700 453.600 ;
        RECT 361.300 452.400 361.900 453.600 ;
        RECT 361.200 451.600 362.000 452.400 ;
        RECT 362.800 451.600 363.600 452.400 ;
        RECT 364.500 450.400 365.100 455.600 ;
        RECT 366.100 452.400 366.700 469.600 ;
        RECT 367.600 466.200 368.400 471.800 ;
        RECT 370.800 464.200 371.600 475.800 ;
        RECT 372.500 472.400 373.100 483.600 ;
        RECT 375.700 478.400 376.300 509.700 ;
        RECT 377.200 509.600 378.000 509.700 ;
        RECT 378.800 509.600 379.600 510.400 ;
        RECT 383.600 509.600 384.400 510.400 ;
        RECT 390.000 509.600 390.800 510.400 ;
        RECT 391.600 509.600 392.400 510.400 ;
        RECT 396.400 509.600 397.200 510.400 ;
        RECT 402.800 509.600 403.600 510.400 ;
        RECT 409.200 509.600 410.000 510.400 ;
        RECT 378.800 503.600 379.600 504.400 ;
        RECT 378.900 492.400 379.500 503.600 ;
        RECT 383.700 502.400 384.300 509.600 ;
        RECT 386.800 507.600 387.600 508.400 ;
        RECT 396.400 507.600 397.200 508.400 ;
        RECT 383.600 501.600 384.400 502.400 ;
        RECT 383.700 498.400 384.300 501.600 ;
        RECT 383.600 497.600 384.400 498.400 ;
        RECT 377.200 491.600 378.000 492.400 ;
        RECT 378.800 491.600 379.600 492.400 ;
        RECT 377.300 488.400 377.900 491.600 ;
        RECT 378.800 489.600 379.600 490.400 ;
        RECT 377.200 487.600 378.000 488.400 ;
        RECT 375.600 477.600 376.400 478.400 ;
        RECT 372.400 471.600 373.200 472.400 ;
        RECT 372.500 468.400 373.100 471.600 ;
        RECT 378.900 470.400 379.500 489.600 ;
        RECT 380.400 487.600 381.200 488.400 ;
        RECT 385.200 486.200 386.000 497.800 ;
        RECT 386.900 496.400 387.500 507.600 ;
        RECT 393.200 503.600 394.000 504.400 ;
        RECT 391.600 501.600 392.400 502.400 ;
        RECT 386.800 495.600 387.600 496.400 ;
        RECT 386.900 490.400 387.500 495.600 ;
        RECT 391.700 492.400 392.300 501.600 ;
        RECT 393.300 500.400 393.900 503.600 ;
        RECT 393.200 499.600 394.000 500.400 ;
        RECT 393.200 495.600 394.000 496.400 ;
        RECT 391.600 491.600 392.400 492.400 ;
        RECT 386.800 489.600 387.600 490.400 ;
        RECT 394.800 486.200 395.600 497.800 ;
        RECT 396.500 494.400 397.100 507.600 ;
        RECT 396.400 493.600 397.200 494.400 ;
        RECT 391.600 479.600 392.400 480.400 ;
        RECT 374.000 469.600 374.800 470.400 ;
        RECT 378.800 469.600 379.600 470.400 ;
        RECT 372.400 467.600 373.200 468.400 ;
        RECT 375.600 459.600 376.400 460.400 ;
        RECT 372.400 457.600 373.200 458.400 ;
        RECT 369.200 455.600 370.000 456.400 ;
        RECT 369.300 454.400 369.900 455.600 ;
        RECT 369.200 453.600 370.000 454.400 ;
        RECT 372.500 452.400 373.100 457.600 ;
        RECT 375.700 452.400 376.300 459.600 ;
        RECT 377.200 457.600 378.000 458.400 ;
        RECT 377.300 452.400 377.900 457.600 ;
        RECT 366.000 451.600 366.800 452.400 ;
        RECT 367.600 451.600 368.400 452.400 ;
        RECT 372.400 451.600 373.200 452.400 ;
        RECT 375.600 451.600 376.400 452.400 ;
        RECT 377.200 451.600 378.000 452.400 ;
        RECT 367.700 450.400 368.300 451.600 ;
        RECT 364.400 449.600 365.200 450.400 ;
        RECT 367.600 449.600 368.400 450.400 ;
        RECT 375.700 444.400 376.300 451.600 ;
        RECT 375.600 443.600 376.400 444.400 ;
        RECT 372.400 437.600 373.200 438.400 ;
        RECT 367.600 435.600 368.400 436.400 ;
        RECT 364.400 431.600 365.200 432.400 ;
        RECT 361.200 429.600 362.000 430.400 ;
        RECT 358.000 427.600 358.800 428.400 ;
        RECT 358.100 418.400 358.700 427.600 ;
        RECT 364.500 420.400 365.100 431.600 ;
        RECT 367.700 430.400 368.300 435.600 ;
        RECT 372.500 430.400 373.100 437.600 ;
        RECT 378.900 430.400 379.500 469.600 ;
        RECT 380.400 464.200 381.200 475.800 ;
        RECT 385.200 475.600 386.000 476.400 ;
        RECT 391.700 470.400 392.300 479.600 ;
        RECT 393.200 475.600 394.000 476.400 ;
        RECT 393.300 472.400 393.900 475.600 ;
        RECT 393.200 471.600 394.000 472.400 ;
        RECT 396.500 472.300 397.100 493.600 ;
        RECT 398.000 490.200 398.800 495.800 ;
        RECT 399.600 493.600 400.400 494.400 ;
        RECT 399.700 490.400 400.300 493.600 ;
        RECT 401.200 491.600 402.000 492.400 ;
        RECT 399.600 489.600 400.400 490.400 ;
        RECT 402.900 474.400 403.500 509.600 ;
        RECT 410.900 506.400 411.500 511.600 ;
        RECT 415.600 509.600 416.400 510.400 ;
        RECT 414.000 507.600 414.800 508.400 ;
        RECT 410.800 505.600 411.600 506.400 ;
        RECT 404.400 501.600 405.200 502.400 ;
        RECT 404.500 498.400 405.100 501.600 ;
        RECT 404.400 497.600 405.200 498.400 ;
        RECT 410.800 493.600 411.600 494.400 ;
        RECT 409.200 491.600 410.000 492.400 ;
        RECT 406.000 489.600 406.800 490.400 ;
        RECT 406.100 488.400 406.700 489.600 ;
        RECT 406.000 487.600 406.800 488.400 ;
        RECT 406.100 484.400 406.700 487.600 ;
        RECT 406.000 483.600 406.800 484.400 ;
        RECT 407.600 477.600 408.400 478.400 ;
        RECT 402.800 473.600 403.600 474.400 ;
        RECT 396.500 471.700 398.700 472.300 ;
        RECT 391.600 469.600 392.400 470.400 ;
        RECT 396.400 469.600 397.200 470.400 ;
        RECT 388.400 467.600 389.200 468.400 ;
        RECT 388.500 464.400 389.100 467.600 ;
        RECT 388.400 463.600 389.200 464.400 ;
        RECT 393.200 463.600 394.000 464.400 ;
        RECT 382.000 453.600 382.800 454.400 ;
        RECT 383.600 453.600 384.400 454.400 ;
        RECT 386.800 453.600 387.600 454.400 ;
        RECT 382.000 449.600 382.800 450.400 ;
        RECT 382.100 438.400 382.700 449.600 ;
        RECT 382.000 437.600 382.800 438.400 ;
        RECT 382.000 435.600 382.800 436.400 ;
        RECT 382.100 430.400 382.700 435.600 ;
        RECT 367.600 429.600 368.400 430.400 ;
        RECT 372.400 429.600 373.200 430.400 ;
        RECT 377.200 429.600 378.000 430.400 ;
        RECT 378.800 429.600 379.600 430.400 ;
        RECT 382.000 429.600 382.800 430.400 ;
        RECT 369.200 427.600 370.000 428.400 ;
        RECT 374.000 423.600 374.800 424.400 ;
        RECT 364.400 419.600 365.200 420.400 ;
        RECT 367.600 419.600 368.400 420.400 ;
        RECT 358.000 417.600 358.800 418.400 ;
        RECT 366.000 417.600 366.800 418.400 ;
        RECT 361.200 415.600 362.000 416.400 ;
        RECT 364.400 415.600 365.200 416.400 ;
        RECT 364.500 412.400 365.100 415.600 ;
        RECT 366.100 414.400 366.700 417.600 ;
        RECT 367.700 416.400 368.300 419.600 ;
        RECT 374.100 416.400 374.700 423.600 ;
        RECT 377.300 420.400 377.900 429.600 ;
        RECT 380.400 427.600 381.200 428.400 ;
        RECT 377.200 419.600 378.000 420.400 ;
        RECT 367.600 415.600 368.400 416.400 ;
        RECT 369.200 416.300 370.000 416.400 ;
        RECT 369.200 415.700 373.100 416.300 ;
        RECT 369.200 415.600 370.000 415.700 ;
        RECT 372.500 414.400 373.100 415.700 ;
        RECT 374.000 415.600 374.800 416.400 ;
        RECT 366.000 413.600 366.800 414.400 ;
        RECT 370.800 413.600 371.600 414.400 ;
        RECT 372.400 413.600 373.200 414.400 ;
        RECT 356.400 411.600 357.200 412.400 ;
        RECT 364.400 411.600 365.200 412.400 ;
        RECT 353.200 409.600 354.000 410.400 ;
        RECT 359.600 409.600 360.400 410.400 ;
        RECT 350.000 407.600 350.800 408.400 ;
        RECT 326.000 399.600 326.800 400.400 ;
        RECT 337.200 399.600 338.000 400.400 ;
        RECT 337.300 398.400 337.900 399.600 ;
        RECT 311.600 389.600 312.400 390.400 ;
        RECT 286.000 377.600 286.800 378.400 ;
        RECT 300.400 377.600 301.200 378.400 ;
        RECT 289.200 373.600 290.000 374.400 ;
        RECT 311.700 372.400 312.300 389.600 ;
        RECT 313.200 384.200 314.000 397.800 ;
        RECT 314.800 384.200 315.600 397.800 ;
        RECT 316.400 384.200 317.200 395.800 ;
        RECT 318.000 387.600 318.800 388.400 ;
        RECT 318.100 382.400 318.700 387.600 ;
        RECT 319.600 384.200 320.400 395.800 ;
        RECT 321.200 385.600 322.000 386.400 ;
        RECT 321.200 383.600 322.000 384.400 ;
        RECT 322.800 384.200 323.600 395.800 ;
        RECT 324.400 384.200 325.200 397.800 ;
        RECT 326.000 384.200 326.800 397.800 ;
        RECT 327.600 384.200 328.400 397.800 ;
        RECT 329.200 397.600 330.000 398.400 ;
        RECT 337.200 397.600 338.000 398.400 ;
        RECT 342.000 397.600 342.800 398.400 ;
        RECT 313.200 381.600 314.000 382.400 ;
        RECT 318.000 381.600 318.800 382.400 ;
        RECT 313.300 378.400 313.900 381.600 ;
        RECT 321.300 378.400 321.900 383.600 ;
        RECT 313.200 377.600 314.000 378.400 ;
        RECT 321.200 377.600 322.000 378.400 ;
        RECT 329.300 376.400 329.900 397.600 ;
        RECT 350.100 386.400 350.700 407.600 ;
        RECT 370.900 400.400 371.500 413.600 ;
        RECT 372.400 411.600 373.200 412.400 ;
        RECT 375.600 411.600 376.400 412.400 ;
        RECT 375.700 410.400 376.300 411.600 ;
        RECT 377.300 410.400 377.900 419.600 ;
        RECT 382.000 418.300 382.800 418.400 ;
        RECT 383.700 418.300 384.300 453.600 ;
        RECT 386.900 452.400 387.500 453.600 ;
        RECT 385.200 451.600 386.000 452.400 ;
        RECT 386.800 451.600 387.600 452.400 ;
        RECT 385.300 444.400 385.900 451.600 ;
        RECT 385.200 443.600 386.000 444.400 ;
        RECT 385.300 432.400 385.900 443.600 ;
        RECT 385.200 431.600 386.000 432.400 ;
        RECT 385.200 429.600 386.000 430.400 ;
        RECT 382.000 417.700 384.300 418.300 ;
        RECT 382.000 417.600 382.800 417.700 ;
        RECT 380.400 415.600 381.200 416.400 ;
        RECT 380.500 412.400 381.100 415.600 ;
        RECT 382.100 414.400 382.700 417.600 ;
        RECT 383.600 416.300 384.400 416.400 ;
        RECT 385.300 416.300 385.900 429.600 ;
        RECT 388.500 428.400 389.100 463.600 ;
        RECT 390.000 453.600 390.800 454.400 ;
        RECT 390.000 449.600 390.800 450.400 ;
        RECT 391.600 450.200 392.400 455.800 ;
        RECT 393.300 430.400 393.900 463.600 ;
        RECT 396.500 462.400 397.100 469.600 ;
        RECT 398.100 468.400 398.700 471.700 ;
        RECT 398.000 467.600 398.800 468.400 ;
        RECT 399.600 467.600 400.400 468.400 ;
        RECT 399.700 466.400 400.300 467.600 ;
        RECT 398.000 465.600 398.800 466.400 ;
        RECT 399.600 465.600 400.400 466.400 ;
        RECT 402.800 466.200 403.600 471.800 ;
        RECT 404.400 471.600 405.200 472.400 ;
        RECT 404.500 468.400 405.100 471.600 ;
        RECT 404.400 467.600 405.200 468.400 ;
        RECT 404.500 466.400 405.100 467.600 ;
        RECT 404.400 465.600 405.200 466.400 ;
        RECT 396.400 461.600 397.200 462.400 ;
        RECT 396.400 459.600 397.200 460.400 ;
        RECT 394.800 446.200 395.600 457.800 ;
        RECT 396.500 430.400 397.100 459.600 ;
        RECT 398.100 454.400 398.700 465.600 ;
        RECT 401.200 463.600 402.000 464.400 ;
        RECT 406.000 464.200 406.800 475.800 ;
        RECT 398.000 453.600 398.800 454.400 ;
        RECT 399.600 453.600 400.400 454.400 ;
        RECT 399.700 452.400 400.300 453.600 ;
        RECT 399.600 451.600 400.400 452.400 ;
        RECT 401.300 450.400 401.900 463.600 ;
        RECT 401.200 449.600 402.000 450.400 ;
        RECT 404.400 446.200 405.200 457.800 ;
        RECT 406.000 433.600 406.800 434.400 ;
        RECT 398.000 431.600 398.800 432.400 ;
        RECT 406.100 430.400 406.700 433.600 ;
        RECT 407.700 430.400 408.300 477.600 ;
        RECT 409.200 475.600 410.000 476.400 ;
        RECT 409.300 470.400 409.900 475.600 ;
        RECT 410.900 472.400 411.500 493.600 ;
        RECT 412.400 490.200 413.200 495.800 ;
        RECT 415.600 486.200 416.400 497.800 ;
        RECT 418.900 496.400 419.500 533.600 ;
        RECT 420.500 510.400 421.100 543.700 ;
        RECT 430.100 534.400 430.700 545.600 ;
        RECT 433.200 544.200 434.000 555.800 ;
        RECT 434.800 547.600 435.600 548.400 ;
        RECT 434.900 544.400 435.500 547.600 ;
        RECT 436.400 546.200 437.200 551.800 ;
        RECT 444.400 551.600 445.200 552.400 ;
        RECT 463.600 551.600 464.400 552.400 ;
        RECT 439.600 549.600 440.400 550.400 ;
        RECT 441.200 549.600 442.000 550.400 ;
        RECT 447.600 549.600 448.400 550.400 ;
        RECT 438.000 547.600 438.800 548.400 ;
        RECT 434.800 543.600 435.600 544.400 ;
        RECT 434.900 534.400 435.500 543.600 ;
        RECT 438.100 538.400 438.700 547.600 ;
        RECT 430.000 533.600 430.800 534.400 ;
        RECT 434.800 533.600 435.600 534.400 ;
        RECT 430.100 522.400 430.700 533.600 ;
        RECT 433.200 531.600 434.000 532.400 ;
        RECT 431.600 523.600 432.400 524.400 ;
        RECT 430.000 521.600 430.800 522.400 ;
        RECT 431.700 520.400 432.300 523.600 ;
        RECT 431.600 519.600 432.400 520.400 ;
        RECT 428.400 511.600 429.200 512.400 ;
        RECT 420.400 509.600 421.200 510.400 ;
        RECT 422.000 509.600 422.800 510.400 ;
        RECT 425.200 510.300 426.000 510.400 ;
        RECT 425.200 509.700 427.500 510.300 ;
        RECT 425.200 509.600 426.000 509.700 ;
        RECT 420.500 498.300 421.100 509.600 ;
        RECT 422.100 504.400 422.700 509.600 ;
        RECT 423.600 507.600 424.400 508.400 ;
        RECT 422.000 503.600 422.800 504.400 ;
        RECT 422.100 502.400 422.700 503.600 ;
        RECT 422.000 501.600 422.800 502.400 ;
        RECT 420.500 497.700 422.700 498.300 ;
        RECT 418.800 495.600 419.600 496.400 ;
        RECT 420.400 495.600 421.200 496.400 ;
        RECT 418.900 494.400 419.500 495.600 ;
        RECT 418.800 493.600 419.600 494.400 ;
        RECT 420.500 492.400 421.100 495.600 ;
        RECT 420.400 491.600 421.200 492.400 ;
        RECT 414.000 473.600 414.800 474.400 ;
        RECT 410.800 471.600 411.600 472.400 ;
        RECT 409.200 469.600 410.000 470.400 ;
        RECT 410.900 462.400 411.500 471.600 ;
        RECT 410.800 461.600 411.600 462.400 ;
        RECT 410.800 455.600 411.600 456.400 ;
        RECT 412.400 455.600 413.200 456.400 ;
        RECT 410.800 452.300 411.600 452.400 ;
        RECT 412.500 452.300 413.100 455.600 ;
        RECT 414.100 452.400 414.700 473.600 ;
        RECT 415.600 464.200 416.400 475.800 ;
        RECT 422.100 468.400 422.700 497.700 ;
        RECT 425.200 486.200 426.000 497.800 ;
        RECT 426.900 484.400 427.500 509.700 ;
        RECT 428.500 508.400 429.100 511.600 ;
        RECT 428.400 507.600 429.200 508.400 ;
        RECT 428.400 503.600 429.200 504.400 ;
        RECT 431.600 503.600 432.400 504.400 ;
        RECT 433.300 504.300 433.900 531.600 ;
        RECT 436.400 526.200 437.200 537.800 ;
        RECT 438.000 537.600 438.800 538.400 ;
        RECT 438.000 533.600 438.800 534.400 ;
        RECT 438.100 532.400 438.700 533.600 ;
        RECT 438.000 531.600 438.800 532.400 ;
        RECT 438.000 529.600 438.800 530.400 ;
        RECT 438.100 520.400 438.700 529.600 ;
        RECT 439.700 528.400 440.300 549.600 ;
        RECT 444.400 531.800 445.200 532.600 ;
        RECT 444.500 528.400 445.100 531.800 ;
        RECT 439.600 527.600 440.400 528.400 ;
        RECT 444.400 527.600 445.200 528.400 ;
        RECT 446.000 526.200 446.800 537.800 ;
        RECT 447.700 534.400 448.300 549.600 ;
        RECT 449.200 547.600 450.000 548.400 ;
        RECT 457.200 547.600 458.000 548.400 ;
        RECT 449.300 546.400 449.900 547.600 ;
        RECT 449.200 545.600 450.000 546.400 ;
        RECT 455.600 545.600 456.400 546.400 ;
        RECT 450.800 543.600 451.600 544.400 ;
        RECT 450.900 540.400 451.500 543.600 ;
        RECT 450.800 539.600 451.600 540.400 ;
        RECT 450.800 537.600 451.600 538.400 ;
        RECT 447.600 533.600 448.400 534.400 ;
        RECT 449.200 530.200 450.000 535.800 ;
        RECT 450.900 534.400 451.500 537.600 ;
        RECT 455.700 536.400 456.300 545.600 ;
        RECT 455.600 535.600 456.400 536.400 ;
        RECT 450.800 533.600 451.600 534.400 ;
        RECT 452.400 531.600 453.200 532.400 ;
        RECT 454.000 531.600 454.800 532.400 ;
        RECT 452.400 527.600 453.200 528.400 ;
        RECT 452.400 525.600 453.200 526.400 ;
        RECT 438.000 519.600 438.800 520.400 ;
        RECT 436.400 511.600 437.200 512.400 ;
        RECT 434.800 509.600 435.600 510.400 ;
        RECT 434.900 506.400 435.500 509.600 ;
        RECT 436.400 507.600 437.200 508.400 ;
        RECT 434.800 505.600 435.600 506.400 ;
        RECT 433.300 503.700 435.500 504.300 ;
        RECT 425.200 483.600 426.000 484.400 ;
        RECT 426.800 483.600 427.600 484.400 ;
        RECT 425.300 468.400 425.900 483.600 ;
        RECT 426.800 479.600 427.600 480.400 ;
        RECT 426.900 472.400 427.500 479.600 ;
        RECT 426.800 471.600 427.600 472.400 ;
        RECT 422.000 467.600 422.800 468.400 ;
        RECT 425.200 467.600 426.000 468.400 ;
        RECT 420.400 465.600 421.200 466.400 ;
        RECT 420.500 464.400 421.100 465.600 ;
        RECT 420.400 463.600 421.200 464.400 ;
        RECT 423.600 463.600 424.400 464.400 ;
        RECT 415.600 461.600 416.400 462.400 ;
        RECT 415.700 454.400 416.300 461.600 ;
        RECT 415.600 453.600 416.400 454.400 ;
        RECT 422.000 453.600 422.800 454.400 ;
        RECT 410.800 451.700 413.100 452.300 ;
        RECT 410.800 451.600 411.600 451.700 ;
        RECT 414.000 451.600 414.800 452.400 ;
        RECT 420.400 451.600 421.200 452.400 ;
        RECT 423.700 452.300 424.300 463.600 ;
        RECT 428.500 456.300 429.100 503.600 ;
        RECT 430.000 487.600 430.800 488.400 ;
        RECT 430.000 485.600 430.800 486.400 ;
        RECT 430.100 480.400 430.700 485.600 ;
        RECT 430.000 479.600 430.800 480.400 ;
        RECT 430.100 472.400 430.700 479.600 ;
        RECT 431.700 474.400 432.300 503.600 ;
        RECT 434.900 498.400 435.500 503.700 ;
        RECT 433.200 497.600 434.000 498.400 ;
        RECT 434.800 497.600 435.600 498.400 ;
        RECT 433.300 492.400 433.900 497.600 ;
        RECT 438.100 492.400 438.700 519.600 ;
        RECT 452.500 518.400 453.100 525.600 ;
        RECT 452.400 517.600 453.200 518.400 ;
        RECT 454.100 510.400 454.700 531.600 ;
        RECT 457.300 528.400 457.900 547.600 ;
        RECT 458.800 543.600 459.600 544.400 ;
        RECT 458.900 532.400 459.500 543.600 ;
        RECT 458.800 531.600 459.600 532.400 ;
        RECT 462.000 529.600 462.800 530.400 ;
        RECT 457.200 527.600 458.000 528.400 ;
        RECT 441.200 509.600 442.000 510.400 ;
        RECT 447.600 509.600 448.400 510.400 ;
        RECT 454.000 509.600 454.800 510.400 ;
        RECT 455.600 509.600 456.400 510.400 ;
        RECT 439.600 507.600 440.400 508.400 ;
        RECT 444.400 503.600 445.200 504.400 ;
        RECT 441.200 493.600 442.000 494.400 ;
        RECT 433.200 491.600 434.000 492.400 ;
        RECT 438.000 491.600 438.800 492.400 ;
        RECT 439.600 491.600 440.400 492.400 ;
        RECT 433.200 479.600 434.000 480.400 ;
        RECT 431.600 473.600 432.400 474.400 ;
        RECT 430.000 471.600 430.800 472.400 ;
        RECT 433.300 470.400 433.900 479.600 ;
        RECT 438.100 476.400 438.700 491.600 ;
        RECT 434.800 475.600 435.600 476.400 ;
        RECT 438.000 475.600 438.800 476.400 ;
        RECT 434.900 470.400 435.500 475.600 ;
        RECT 438.000 471.600 438.800 472.400 ;
        RECT 433.200 469.600 434.000 470.400 ;
        RECT 434.800 469.600 435.600 470.400 ;
        RECT 438.100 468.400 438.700 471.600 ;
        RECT 439.700 470.400 440.300 491.600 ;
        RECT 441.300 490.300 441.900 493.600 ;
        RECT 444.500 492.400 445.100 503.600 ;
        RECT 447.700 498.400 448.300 509.600 ;
        RECT 454.100 508.400 454.700 509.600 ;
        RECT 454.000 507.600 454.800 508.400 ;
        RECT 449.200 503.600 450.000 504.400 ;
        RECT 447.600 497.600 448.400 498.400 ;
        RECT 447.600 495.600 448.400 496.400 ;
        RECT 442.800 492.300 443.600 492.400 ;
        RECT 444.400 492.300 445.200 492.400 ;
        RECT 442.800 491.700 445.200 492.300 ;
        RECT 442.800 491.600 443.600 491.700 ;
        RECT 444.400 491.600 445.200 491.700 ;
        RECT 441.300 489.700 443.500 490.300 ;
        RECT 441.200 473.600 442.000 474.400 ;
        RECT 441.300 470.400 441.900 473.600 ;
        RECT 442.900 472.400 443.500 489.700 ;
        RECT 446.000 489.600 446.800 490.400 ;
        RECT 446.100 488.400 446.700 489.600 ;
        RECT 446.000 487.600 446.800 488.400 ;
        RECT 446.100 474.400 446.700 487.600 ;
        RECT 447.600 479.600 448.400 480.400 ;
        RECT 447.700 478.400 448.300 479.600 ;
        RECT 449.300 478.400 449.900 503.600 ;
        RECT 455.700 502.400 456.300 509.600 ;
        RECT 463.700 506.400 464.300 551.600 ;
        RECT 466.800 544.200 467.600 555.800 ;
        RECT 468.400 549.600 469.200 550.400 ;
        RECT 468.500 544.400 469.100 549.600 ;
        RECT 474.800 549.400 475.600 550.400 ;
        RECT 468.400 543.600 469.200 544.400 ;
        RECT 476.400 544.200 477.200 555.800 ;
        RECT 494.000 553.600 494.800 554.400 ;
        RECT 494.100 552.400 494.700 553.600 ;
        RECT 478.000 549.600 478.800 550.400 ;
        RECT 474.800 537.600 475.600 538.400 ;
        RECT 466.800 535.600 467.600 536.400 ;
        RECT 466.900 534.400 467.500 535.600 ;
        RECT 474.900 534.400 475.500 537.600 ;
        RECT 478.100 534.400 478.700 549.600 ;
        RECT 479.600 546.200 480.400 551.800 ;
        RECT 487.600 551.600 488.400 552.400 ;
        RECT 494.000 551.600 494.800 552.400 ;
        RECT 482.800 549.600 483.600 550.400 ;
        RECT 486.000 549.600 486.800 550.400 ;
        RECT 490.800 549.600 491.600 550.400 ;
        RECT 481.200 547.600 482.000 548.400 ;
        RECT 481.300 538.400 481.900 547.600 ;
        RECT 481.200 537.600 482.000 538.400 ;
        RECT 465.200 533.600 466.000 534.400 ;
        RECT 466.800 533.600 467.600 534.400 ;
        RECT 471.600 533.600 472.400 534.400 ;
        RECT 474.800 533.600 475.600 534.400 ;
        RECT 478.000 533.600 478.800 534.400 ;
        RECT 465.300 532.400 465.900 533.600 ;
        RECT 482.900 532.400 483.500 549.600 ;
        RECT 486.100 548.400 486.700 549.600 ;
        RECT 486.000 547.600 486.800 548.400 ;
        RECT 486.000 543.600 486.800 544.400 ;
        RECT 486.100 534.400 486.700 543.600 ;
        RECT 487.600 537.600 488.400 538.400 ;
        RECT 487.700 534.400 488.300 537.600 ;
        RECT 490.900 534.400 491.500 549.600 ;
        RECT 492.400 547.600 493.200 548.400 ;
        RECT 492.500 544.400 493.100 547.600 ;
        RECT 492.400 543.600 493.200 544.400 ;
        RECT 498.800 544.200 499.600 555.800 ;
        RECT 505.200 549.600 506.000 550.400 ;
        RECT 508.400 544.200 509.200 555.800 ;
        RECT 510.000 547.600 510.800 548.400 ;
        RECT 492.500 536.400 493.100 543.600 ;
        RECT 510.100 542.400 510.700 547.600 ;
        RECT 511.600 546.200 512.400 551.800 ;
        RECT 518.000 551.600 518.800 552.400 ;
        RECT 521.200 552.300 522.000 552.400 ;
        RECT 521.200 551.700 523.500 552.300 ;
        RECT 521.200 551.600 522.000 551.700 ;
        RECT 521.300 550.400 521.900 551.600 ;
        RECT 514.800 549.600 515.600 550.400 ;
        RECT 519.600 549.600 520.400 550.400 ;
        RECT 521.200 549.600 522.000 550.400 ;
        RECT 513.200 547.600 514.000 548.400 ;
        RECT 513.300 544.400 513.900 547.600 ;
        RECT 513.200 543.600 514.000 544.400 ;
        RECT 502.000 541.600 502.800 542.400 ;
        RECT 510.000 541.600 510.800 542.400 ;
        RECT 492.400 535.600 493.200 536.400 ;
        RECT 498.800 535.600 499.600 536.400 ;
        RECT 498.900 534.400 499.500 535.600 ;
        RECT 484.400 533.600 485.200 534.400 ;
        RECT 486.000 533.600 486.800 534.400 ;
        RECT 487.600 533.600 488.400 534.400 ;
        RECT 490.800 533.600 491.600 534.400 ;
        RECT 492.400 533.600 493.200 534.400 ;
        RECT 497.200 533.600 498.000 534.400 ;
        RECT 498.800 533.600 499.600 534.400 ;
        RECT 484.500 532.400 485.100 533.600 ;
        RECT 492.500 532.400 493.100 533.600 ;
        RECT 497.300 532.400 497.900 533.600 ;
        RECT 465.200 531.600 466.000 532.400 ;
        RECT 466.800 531.600 467.600 532.400 ;
        RECT 473.200 531.600 474.000 532.400 ;
        RECT 474.800 531.600 475.600 532.400 ;
        RECT 482.800 531.600 483.600 532.400 ;
        RECT 484.400 531.600 485.200 532.400 ;
        RECT 489.200 531.600 490.000 532.400 ;
        RECT 492.400 531.600 493.200 532.400 ;
        RECT 497.200 531.600 498.000 532.400 ;
        RECT 465.200 521.600 466.000 522.400 ;
        RECT 465.300 512.400 465.900 521.600 ;
        RECT 465.200 511.600 466.000 512.400 ;
        RECT 466.900 510.400 467.500 531.600 ;
        RECT 473.300 526.400 473.900 531.600 ;
        RECT 473.200 525.600 474.000 526.400 ;
        RECT 474.900 518.400 475.500 531.600 ;
        RECT 481.200 529.600 482.000 530.400 ;
        RECT 487.600 527.600 488.400 528.400 ;
        RECT 474.800 517.600 475.600 518.400 ;
        RECT 482.800 515.600 483.600 516.400 ;
        RECT 482.900 514.400 483.500 515.600 ;
        RECT 482.800 513.600 483.600 514.400 ;
        RECT 484.400 513.600 485.200 514.400 ;
        RECT 468.400 511.600 469.200 512.400 ;
        RECT 466.800 509.600 467.600 510.400 ;
        RECT 468.500 508.400 469.100 511.600 ;
        RECT 470.000 509.600 470.800 510.400 ;
        RECT 471.600 509.600 472.400 510.400 ;
        RECT 476.400 509.600 477.200 510.400 ;
        RECT 468.400 507.600 469.200 508.400 ;
        RECT 463.600 505.600 464.400 506.400 ;
        RECT 470.100 504.400 470.700 509.600 ;
        RECT 471.700 506.400 472.300 509.600 ;
        RECT 479.600 507.600 480.400 508.400 ;
        RECT 479.700 506.400 480.300 507.600 ;
        RECT 471.600 505.600 472.400 506.400 ;
        RECT 479.600 505.600 480.400 506.400 ;
        RECT 457.200 503.600 458.000 504.400 ;
        RECT 465.200 503.600 466.000 504.400 ;
        RECT 470.000 503.600 470.800 504.400 ;
        RECT 455.600 501.600 456.400 502.400 ;
        RECT 452.400 497.600 453.200 498.400 ;
        RECT 452.500 494.400 453.100 497.600 ;
        RECT 454.000 495.600 454.800 496.400 ;
        RECT 454.100 494.400 454.700 495.600 ;
        RECT 452.400 493.600 453.200 494.400 ;
        RECT 454.000 493.600 454.800 494.400 ;
        RECT 452.400 491.600 453.200 492.400 ;
        RECT 454.000 491.600 454.800 492.400 ;
        RECT 447.600 477.600 448.400 478.400 ;
        RECT 449.200 477.600 450.000 478.400 ;
        RECT 447.600 475.600 448.400 476.400 ;
        RECT 446.000 473.600 446.800 474.400 ;
        RECT 442.800 471.600 443.600 472.400 ;
        RECT 439.600 469.600 440.400 470.400 ;
        RECT 441.200 469.600 442.000 470.400 ;
        RECT 431.600 467.600 432.400 468.400 ;
        RECT 438.000 467.600 438.800 468.400 ;
        RECT 430.000 463.600 430.800 464.400 ;
        RECT 430.100 462.400 430.700 463.600 ;
        RECT 441.300 462.400 441.900 469.600 ;
        RECT 442.900 468.400 443.500 471.600 ;
        RECT 444.400 469.600 445.200 470.400 ;
        RECT 446.000 469.600 446.800 470.400 ;
        RECT 446.100 468.400 446.700 469.600 ;
        RECT 442.800 467.600 443.600 468.400 ;
        RECT 446.000 467.600 446.800 468.400 ;
        RECT 430.000 461.600 430.800 462.400 ;
        RECT 434.800 461.600 435.600 462.400 ;
        RECT 441.200 461.600 442.000 462.400 ;
        RECT 426.900 455.700 429.100 456.300 ;
        RECT 426.900 452.400 427.500 455.700 ;
        RECT 428.400 453.600 429.200 454.400 ;
        RECT 430.000 453.600 430.800 454.400 ;
        RECT 422.100 451.700 424.300 452.300 ;
        RECT 410.900 450.400 411.500 451.600 ;
        RECT 410.800 449.600 411.600 450.400 ;
        RECT 417.200 449.600 418.000 450.400 ;
        RECT 409.200 443.600 410.000 444.400 ;
        RECT 414.000 437.600 414.800 438.400 ;
        RECT 412.400 433.600 413.200 434.400 ;
        RECT 393.200 429.600 394.000 430.400 ;
        RECT 396.400 429.600 397.200 430.400 ;
        RECT 401.200 429.600 402.000 430.400 ;
        RECT 402.800 429.600 403.600 430.400 ;
        RECT 406.000 429.600 406.800 430.400 ;
        RECT 407.600 429.600 408.400 430.400 ;
        RECT 410.800 429.600 411.600 430.400 ;
        RECT 388.400 427.600 389.200 428.400 ;
        RECT 398.000 427.600 398.800 428.400 ;
        RECT 409.200 427.600 410.000 428.400 ;
        RECT 396.400 425.600 397.200 426.400 ;
        RECT 388.400 423.600 389.200 424.400 ;
        RECT 390.000 423.600 390.800 424.400 ;
        RECT 383.600 415.700 385.900 416.300 ;
        RECT 383.600 415.600 384.400 415.700 ;
        RECT 382.000 413.600 382.800 414.400 ;
        RECT 383.700 412.400 384.300 415.600 ;
        RECT 388.500 412.400 389.100 423.600 ;
        RECT 390.100 416.400 390.700 423.600 ;
        RECT 396.500 422.400 397.100 425.600 ;
        RECT 396.400 421.600 397.200 422.400 ;
        RECT 390.000 415.600 390.800 416.400 ;
        RECT 391.600 415.600 392.400 416.400 ;
        RECT 380.400 411.600 381.200 412.400 ;
        RECT 383.600 411.600 384.400 412.400 ;
        RECT 388.400 411.600 389.200 412.400 ;
        RECT 394.800 411.600 395.600 412.400 ;
        RECT 396.400 411.600 397.200 412.400 ;
        RECT 375.600 409.600 376.400 410.400 ;
        RECT 377.200 409.600 378.000 410.400 ;
        RECT 380.400 403.600 381.200 404.400 ;
        RECT 370.800 399.600 371.600 400.400 ;
        RECT 350.000 385.600 350.800 386.400 ;
        RECT 337.200 383.600 338.000 384.400 ;
        RECT 351.600 384.200 352.400 397.800 ;
        RECT 353.200 384.200 354.000 397.800 ;
        RECT 354.800 384.200 355.600 397.800 ;
        RECT 356.400 384.200 357.200 395.800 ;
        RECT 358.000 385.600 358.800 386.400 ;
        RECT 359.600 384.200 360.400 395.800 ;
        RECT 361.200 387.600 362.000 388.400 ;
        RECT 361.300 384.400 361.900 387.600 ;
        RECT 361.200 383.600 362.000 384.400 ;
        RECT 362.800 384.200 363.600 395.800 ;
        RECT 364.400 384.200 365.200 397.800 ;
        RECT 366.000 384.200 366.800 397.800 ;
        RECT 367.600 389.600 368.400 390.400 ;
        RECT 337.300 376.400 337.900 383.600 ;
        RECT 359.600 381.600 360.400 382.400 ;
        RECT 342.000 379.600 342.800 380.400 ;
        RECT 342.100 376.400 342.700 379.600 ;
        RECT 319.600 375.600 320.400 376.400 ;
        RECT 329.200 375.600 330.000 376.400 ;
        RECT 337.200 375.600 338.000 376.400 ;
        RECT 342.000 375.600 342.800 376.400 ;
        RECT 338.800 373.600 339.600 374.400 ;
        RECT 308.400 371.600 309.200 372.400 ;
        RECT 310.000 371.600 310.800 372.400 ;
        RECT 311.600 371.600 312.400 372.400 ;
        RECT 326.000 371.600 326.800 372.400 ;
        RECT 330.800 371.600 331.600 372.400 ;
        RECT 332.400 371.600 333.200 372.400 ;
        RECT 343.600 371.600 344.400 372.400 ;
        RECT 346.800 371.600 347.600 372.400 ;
        RECT 308.500 370.400 309.100 371.600 ;
        RECT 308.400 369.600 309.200 370.400 ;
        RECT 310.100 366.400 310.700 371.600 ;
        RECT 310.000 365.600 310.800 366.400 ;
        RECT 286.000 363.600 286.800 364.400 ;
        RECT 311.700 364.300 312.300 371.600 ;
        RECT 321.200 369.600 322.000 370.400 ;
        RECT 310.100 363.700 312.300 364.300 ;
        RECT 281.200 357.600 282.000 358.400 ;
        RECT 284.400 357.600 285.200 358.400 ;
        RECT 258.800 349.600 259.600 350.400 ;
        RECT 270.000 349.600 270.800 350.400 ;
        RECT 271.600 349.600 272.400 350.400 ;
        RECT 250.800 339.600 251.600 340.400 ;
        RECT 257.200 339.600 258.000 340.400 ;
        RECT 238.000 335.600 238.800 336.400 ;
        RECT 239.600 323.600 240.400 324.400 ;
        RECT 249.200 324.200 250.000 337.800 ;
        RECT 250.800 324.200 251.600 337.800 ;
        RECT 252.400 326.200 253.200 337.800 ;
        RECT 254.000 333.600 254.800 334.400 ;
        RECT 254.000 331.600 254.800 332.400 ;
        RECT 254.100 326.400 254.700 331.600 ;
        RECT 254.000 325.600 254.800 326.400 ;
        RECT 255.600 326.200 256.400 337.800 ;
        RECT 257.300 336.400 257.900 339.600 ;
        RECT 257.200 335.600 258.000 336.400 ;
        RECT 258.800 326.200 259.600 337.800 ;
        RECT 217.200 305.600 218.000 306.400 ;
        RECT 217.300 304.400 217.900 305.600 ;
        RECT 217.200 303.600 218.000 304.400 ;
        RECT 218.800 304.200 219.600 315.800 ;
        RECT 220.400 304.200 221.200 317.800 ;
        RECT 222.000 304.200 222.800 317.800 ;
        RECT 223.600 304.200 224.400 317.800 ;
        RECT 236.400 317.600 237.200 318.400 ;
        RECT 239.700 312.400 240.300 323.600 ;
        RECT 239.600 311.600 240.400 312.400 ;
        RECT 242.800 311.600 243.600 312.400 ;
        RECT 247.600 311.600 248.400 312.400 ;
        RECT 233.200 309.600 234.200 310.400 ;
        RECT 238.000 309.600 238.800 310.400 ;
        RECT 238.100 308.400 238.700 309.600 ;
        RECT 238.000 307.600 238.800 308.400 ;
        RECT 234.800 303.600 235.600 304.400 ;
        RECT 207.600 297.600 208.400 298.400 ;
        RECT 204.400 293.600 205.200 294.400 ;
        RECT 206.000 293.600 206.800 294.400 ;
        RECT 209.200 293.600 210.000 294.400 ;
        RECT 199.600 291.600 200.400 292.400 ;
        RECT 204.500 292.300 205.100 293.600 ;
        RECT 212.400 292.300 213.200 292.400 ;
        RECT 204.500 291.700 213.200 292.300 ;
        RECT 212.400 291.600 213.200 291.700 ;
        RECT 222.000 291.600 222.800 292.400 ;
        RECT 196.400 289.600 197.200 290.400 ;
        RECT 194.800 279.600 195.600 280.400 ;
        RECT 191.600 265.600 192.400 266.400 ;
        RECT 191.700 264.400 192.300 265.600 ;
        RECT 191.600 263.600 192.400 264.400 ;
        RECT 193.200 264.200 194.000 275.800 ;
        RECT 194.800 264.200 195.600 277.800 ;
        RECT 196.400 264.200 197.200 277.800 ;
        RECT 198.000 264.200 198.800 277.800 ;
        RECT 199.700 270.400 200.300 291.600 ;
        RECT 214.000 289.600 214.800 290.400 ;
        RECT 217.200 289.600 218.000 290.400 ;
        RECT 207.600 283.600 208.400 284.400 ;
        RECT 212.400 273.600 213.200 274.400 ;
        RECT 212.500 270.400 213.100 273.600 ;
        RECT 199.600 269.600 200.400 270.400 ;
        RECT 212.400 269.600 213.200 270.400 ;
        RECT 186.800 261.600 187.600 262.400 ;
        RECT 188.400 261.600 189.200 262.400 ;
        RECT 185.200 259.600 186.000 260.400 ;
        RECT 178.800 253.600 179.600 254.400 ;
        RECT 182.000 253.600 182.800 254.400 ;
        RECT 174.000 251.700 176.300 252.300 ;
        RECT 174.000 251.600 174.800 251.700 ;
        RECT 162.800 241.600 163.600 242.400 ;
        RECT 143.600 225.600 144.400 226.400 ;
        RECT 142.000 206.200 142.800 217.800 ;
        RECT 143.700 214.400 144.300 225.600 ;
        RECT 158.000 224.200 158.800 237.800 ;
        RECT 159.600 224.200 160.400 237.800 ;
        RECT 161.200 224.200 162.000 235.800 ;
        RECT 162.900 228.400 163.500 241.600 ;
        RECT 162.800 227.600 163.600 228.400 ;
        RECT 164.400 224.200 165.200 235.800 ;
        RECT 166.000 225.600 166.800 226.400 ;
        RECT 166.100 218.400 166.700 225.600 ;
        RECT 167.600 224.200 168.400 235.800 ;
        RECT 169.200 224.200 170.000 237.800 ;
        RECT 170.800 224.200 171.600 237.800 ;
        RECT 172.400 224.200 173.200 237.800 ;
        RECT 174.100 230.400 174.700 251.600 ;
        RECT 178.900 244.400 179.500 253.600 ;
        RECT 182.000 249.600 182.800 250.400 ;
        RECT 178.800 243.600 179.600 244.400 ;
        RECT 182.100 242.400 182.700 249.600 ;
        RECT 182.000 241.600 182.800 242.400 ;
        RECT 182.000 237.600 182.800 238.400 ;
        RECT 174.000 229.600 174.800 230.400 ;
        RECT 185.300 228.400 185.900 259.600 ;
        RECT 186.900 252.400 187.500 261.600 ;
        RECT 188.500 254.400 189.100 261.600 ;
        RECT 193.200 259.600 194.000 260.400 ;
        RECT 193.300 254.400 193.900 259.600 ;
        RECT 188.400 253.600 189.200 254.400 ;
        RECT 193.200 253.600 194.000 254.400 ;
        RECT 186.800 251.600 187.600 252.400 ;
        RECT 186.800 241.600 187.600 242.400 ;
        RECT 186.900 238.400 187.500 241.600 ;
        RECT 193.300 238.400 193.900 253.600 ;
        RECT 199.700 252.400 200.300 269.600 ;
        RECT 207.600 267.600 208.600 268.400 ;
        RECT 212.400 267.600 213.200 268.400 ;
        RECT 210.800 263.600 211.600 264.400 ;
        RECT 199.600 251.600 200.400 252.400 ;
        RECT 202.800 244.200 203.600 257.800 ;
        RECT 204.400 244.200 205.200 257.800 ;
        RECT 206.000 246.200 206.800 257.800 ;
        RECT 207.600 253.600 208.400 254.400 ;
        RECT 209.200 246.200 210.000 257.800 ;
        RECT 210.900 256.400 211.500 263.600 ;
        RECT 214.100 262.400 214.700 289.600 ;
        RECT 217.300 274.400 217.900 289.600 ;
        RECT 226.800 284.200 227.600 297.800 ;
        RECT 228.400 284.200 229.200 297.800 ;
        RECT 230.000 286.200 230.800 297.800 ;
        RECT 231.600 293.600 232.400 294.400 ;
        RECT 233.200 286.200 234.000 297.800 ;
        RECT 234.900 296.400 235.500 303.600 ;
        RECT 234.800 295.600 235.600 296.400 ;
        RECT 236.400 286.200 237.200 297.800 ;
        RECT 236.400 283.600 237.200 284.400 ;
        RECT 238.000 284.200 238.800 297.800 ;
        RECT 239.600 284.200 240.400 297.800 ;
        RECT 241.200 284.200 242.000 297.800 ;
        RECT 242.900 290.400 243.500 311.600 ;
        RECT 247.700 310.400 248.300 311.600 ;
        RECT 247.600 309.600 248.400 310.400 ;
        RECT 249.200 309.600 250.000 310.400 ;
        RECT 246.000 305.600 246.800 306.400 ;
        RECT 247.600 295.600 248.400 296.400 ;
        RECT 242.800 289.600 243.600 290.400 ;
        RECT 228.400 281.600 229.200 282.400 ;
        RECT 228.500 278.400 229.100 281.600 ;
        RECT 228.400 277.600 229.200 278.400 ;
        RECT 217.200 273.600 218.000 274.400 ;
        RECT 217.200 271.600 218.000 272.400 ;
        RECT 222.000 271.600 222.800 272.400 ;
        RECT 217.300 262.400 217.900 271.600 ;
        RECT 220.400 265.600 221.200 266.400 ;
        RECT 225.200 263.600 226.000 264.400 ;
        RECT 214.000 261.600 214.800 262.400 ;
        RECT 217.200 261.600 218.000 262.400 ;
        RECT 210.800 255.600 211.600 256.400 ;
        RECT 212.400 246.200 213.200 257.800 ;
        RECT 214.000 244.200 214.800 257.800 ;
        RECT 215.600 244.200 216.400 257.800 ;
        RECT 217.200 244.200 218.000 257.800 ;
        RECT 225.300 252.400 225.900 263.600 ;
        RECT 236.500 254.400 237.100 283.600 ;
        RECT 239.600 264.200 240.400 277.800 ;
        RECT 241.200 264.200 242.000 277.800 ;
        RECT 242.800 264.200 243.600 275.800 ;
        RECT 244.400 267.600 245.200 268.400 ;
        RECT 246.000 264.200 246.800 275.800 ;
        RECT 247.700 266.400 248.300 295.600 ;
        RECT 249.300 282.400 249.900 309.600 ;
        RECT 254.100 308.400 254.700 325.600 ;
        RECT 258.800 323.600 259.600 324.400 ;
        RECT 260.400 324.200 261.200 337.800 ;
        RECT 262.000 324.200 262.800 337.800 ;
        RECT 263.600 324.200 264.400 337.800 ;
        RECT 268.400 333.600 269.200 334.400 ;
        RECT 258.900 318.400 259.500 323.600 ;
        RECT 268.500 318.400 269.100 333.600 ;
        RECT 258.800 317.600 259.600 318.400 ;
        RECT 268.400 317.600 269.200 318.400 ;
        RECT 270.100 314.400 270.700 349.600 ;
        RECT 271.700 340.400 272.300 349.600 ;
        RECT 273.200 347.600 274.000 348.400 ;
        RECT 273.300 346.400 273.900 347.600 ;
        RECT 281.300 346.400 281.900 357.600 ;
        RECT 286.100 350.400 286.700 363.600 ;
        RECT 289.200 351.600 290.000 352.400 ;
        RECT 289.300 350.400 289.900 351.600 ;
        RECT 286.000 349.600 286.800 350.400 ;
        RECT 289.200 349.600 290.000 350.400 ;
        RECT 273.200 345.600 274.000 346.400 ;
        RECT 281.200 345.600 282.000 346.400 ;
        RECT 282.800 345.600 283.600 346.400 ;
        RECT 271.600 339.600 272.400 340.400 ;
        RECT 282.900 336.400 283.500 345.600 ;
        RECT 294.000 344.200 294.800 357.800 ;
        RECT 295.600 344.200 296.400 357.800 ;
        RECT 297.200 344.200 298.000 355.800 ;
        RECT 298.800 347.600 299.600 348.400 ;
        RECT 300.400 344.200 301.200 355.800 ;
        RECT 302.000 349.600 302.800 350.400 ;
        RECT 302.100 346.400 302.700 349.600 ;
        RECT 302.000 345.600 302.800 346.400 ;
        RECT 303.600 344.200 304.400 355.800 ;
        RECT 305.200 344.200 306.000 357.800 ;
        RECT 306.800 344.200 307.600 357.800 ;
        RECT 308.400 344.200 309.200 357.800 ;
        RECT 310.100 350.400 310.700 363.700 ;
        RECT 321.300 350.400 321.900 369.600 ;
        RECT 310.000 349.600 310.800 350.400 ;
        RECT 318.000 349.600 319.000 350.400 ;
        RECT 321.200 349.600 322.000 350.400 ;
        RECT 324.400 349.600 325.200 350.400 ;
        RECT 321.200 343.600 322.000 344.400 ;
        RECT 294.000 339.600 294.800 340.400 ;
        RECT 292.400 337.600 293.200 338.400 ;
        RECT 273.200 335.600 274.000 336.400 ;
        RECT 278.000 335.600 278.800 336.400 ;
        RECT 282.800 335.600 283.600 336.400 ;
        RECT 287.600 331.600 288.400 332.400 ;
        RECT 290.800 331.600 291.600 332.400 ;
        RECT 281.200 329.600 282.000 330.400 ;
        RECT 284.400 329.600 285.200 330.400 ;
        RECT 281.300 328.400 281.900 329.600 ;
        RECT 287.700 328.400 288.300 331.600 ;
        RECT 290.900 330.400 291.500 331.600 ;
        RECT 290.800 329.600 291.600 330.400 ;
        RECT 281.200 327.600 282.000 328.400 ;
        RECT 287.600 327.600 288.400 328.400 ;
        RECT 276.400 323.600 277.200 324.400 ;
        RECT 279.600 323.600 280.400 324.400 ;
        RECT 289.200 323.600 290.000 324.400 ;
        RECT 265.200 313.600 266.000 314.400 ;
        RECT 270.000 313.600 270.800 314.400 ;
        RECT 257.200 311.600 258.000 312.400 ;
        RECT 257.300 310.400 257.900 311.600 ;
        RECT 265.300 310.400 265.900 313.600 ;
        RECT 271.600 312.300 272.400 312.400 ;
        RECT 271.600 311.700 273.900 312.300 ;
        RECT 271.600 311.600 272.400 311.700 ;
        RECT 257.200 309.600 258.000 310.400 ;
        RECT 262.000 309.600 262.800 310.400 ;
        RECT 265.200 309.600 266.000 310.400 ;
        RECT 266.800 309.600 267.600 310.400 ;
        RECT 254.000 308.300 254.800 308.400 ;
        RECT 254.000 307.700 256.300 308.300 ;
        RECT 254.000 307.600 254.800 307.700 ;
        RECT 255.700 292.400 256.300 307.700 ;
        RECT 263.600 303.600 264.400 304.400 ;
        RECT 263.700 302.400 264.300 303.600 ;
        RECT 263.600 301.600 264.400 302.400 ;
        RECT 257.200 293.600 258.000 294.400 ;
        RECT 263.700 292.400 264.300 301.600 ;
        RECT 255.600 291.600 256.400 292.400 ;
        RECT 263.600 291.600 264.400 292.400 ;
        RECT 265.200 291.600 266.000 292.400 ;
        RECT 250.800 283.600 251.600 284.400 ;
        RECT 249.200 281.600 250.000 282.400 ;
        RECT 247.600 265.600 248.400 266.400 ;
        RECT 242.800 257.600 243.600 258.400 ;
        RECT 233.200 253.600 234.000 254.400 ;
        RECT 236.400 253.600 237.200 254.400 ;
        RECT 239.600 253.600 240.400 254.400 ;
        RECT 239.700 252.400 240.300 253.600 ;
        RECT 242.900 252.400 243.500 257.600 ;
        RECT 247.700 256.400 248.300 265.600 ;
        RECT 249.200 264.200 250.000 275.800 ;
        RECT 250.800 264.200 251.600 277.800 ;
        RECT 252.400 264.200 253.200 277.800 ;
        RECT 254.000 264.200 254.800 277.800 ;
        RECT 255.700 270.400 256.300 291.600 ;
        RECT 255.600 269.600 256.400 270.400 ;
        RECT 265.300 270.300 265.900 291.600 ;
        RECT 266.900 286.400 267.500 309.600 ;
        RECT 273.300 308.400 273.900 311.700 ;
        RECT 274.800 311.600 275.600 312.400 ;
        RECT 274.800 310.300 275.600 310.400 ;
        RECT 276.500 310.300 277.100 323.600 ;
        RECT 279.700 310.400 280.300 323.600 ;
        RECT 289.300 314.400 289.900 323.600 ;
        RECT 289.200 313.600 290.000 314.400 ;
        RECT 284.400 311.600 285.200 312.400 ;
        RECT 292.500 310.400 293.100 337.600 ;
        RECT 294.100 328.400 294.700 339.600 ;
        RECT 321.300 334.400 321.900 343.600 ;
        RECT 324.500 342.400 325.100 349.600 ;
        RECT 326.100 344.400 326.700 371.600 ;
        RECT 330.900 370.400 331.500 371.600 ;
        RECT 330.800 369.600 331.600 370.400 ;
        RECT 327.600 349.600 328.400 350.400 ;
        RECT 327.700 346.400 328.300 349.600 ;
        RECT 329.200 347.600 330.000 348.400 ;
        RECT 329.300 346.400 329.900 347.600 ;
        RECT 327.600 345.600 328.400 346.400 ;
        RECT 329.200 345.600 330.000 346.400 ;
        RECT 326.000 343.600 326.800 344.400 ;
        RECT 324.400 341.600 325.200 342.400 ;
        RECT 332.500 338.400 333.100 371.600 ;
        RECT 343.700 350.400 344.300 371.600 ;
        RECT 351.600 364.200 352.400 377.800 ;
        RECT 353.200 364.200 354.000 377.800 ;
        RECT 354.800 366.200 355.600 377.800 ;
        RECT 356.400 373.600 357.200 374.400 ;
        RECT 358.000 366.200 358.800 377.800 ;
        RECT 359.700 376.400 360.300 381.600 ;
        RECT 359.600 375.600 360.400 376.400 ;
        RECT 361.200 366.200 362.000 377.800 ;
        RECT 362.800 364.200 363.600 377.800 ;
        RECT 364.400 364.200 365.200 377.800 ;
        RECT 366.000 364.200 366.800 377.800 ;
        RECT 367.700 372.400 368.300 389.600 ;
        RECT 375.600 386.200 376.400 391.800 ;
        RECT 378.800 384.200 379.600 395.800 ;
        RECT 380.500 390.200 381.100 403.600 ;
        RECT 382.000 399.600 382.800 400.400 ;
        RECT 380.400 389.400 381.200 390.200 ;
        RECT 375.600 379.600 376.400 380.400 ;
        RECT 375.700 378.400 376.300 379.600 ;
        RECT 375.600 377.600 376.400 378.400 ;
        RECT 367.600 371.600 368.400 372.400 ;
        RECT 380.400 369.600 381.200 370.400 ;
        RECT 367.600 359.600 368.400 360.400 ;
        RECT 343.600 349.600 344.400 350.400 ;
        RECT 337.200 347.600 338.000 348.400 ;
        RECT 337.300 346.400 337.900 347.600 ;
        RECT 337.200 345.600 338.000 346.400 ;
        RECT 345.200 345.600 346.000 346.400 ;
        RECT 335.600 341.600 336.400 342.400 ;
        RECT 332.400 337.600 333.200 338.400 ;
        RECT 326.000 335.600 326.800 336.400 ;
        RECT 326.100 334.400 326.700 335.600 ;
        RECT 305.200 333.600 306.000 334.400 ;
        RECT 316.400 333.600 317.200 334.400 ;
        RECT 321.200 333.600 322.000 334.400 ;
        RECT 326.000 333.600 326.800 334.400 ;
        RECT 327.600 333.600 328.400 334.400 ;
        RECT 329.200 333.600 330.000 334.400 ;
        RECT 334.000 333.600 334.800 334.400 ;
        RECT 305.300 332.400 305.900 333.600 ;
        RECT 316.500 332.400 317.100 333.600 ;
        RECT 297.200 331.600 298.000 332.400 ;
        RECT 305.200 331.600 306.000 332.400 ;
        RECT 314.800 331.600 315.600 332.400 ;
        RECT 316.400 331.600 317.200 332.400 ;
        RECT 297.300 330.400 297.900 331.600 ;
        RECT 305.300 330.400 305.900 331.600 ;
        RECT 297.200 329.600 298.000 330.400 ;
        RECT 305.200 329.600 306.000 330.400 ;
        RECT 294.000 327.600 294.800 328.400 ;
        RECT 300.400 327.600 301.200 328.400 ;
        RECT 295.600 323.600 296.400 324.400 ;
        RECT 302.000 323.600 302.800 324.400 ;
        RECT 274.800 309.700 277.100 310.300 ;
        RECT 274.800 309.600 275.600 309.700 ;
        RECT 278.000 309.600 278.800 310.400 ;
        RECT 279.600 309.600 280.400 310.400 ;
        RECT 284.400 309.600 285.200 310.400 ;
        RECT 292.400 309.600 293.200 310.400 ;
        RECT 268.400 307.600 269.200 308.400 ;
        RECT 273.200 307.600 274.000 308.400 ;
        RECT 266.800 285.600 267.600 286.400 ;
        RECT 266.900 282.400 267.500 285.600 ;
        RECT 266.800 281.600 267.600 282.400 ;
        RECT 268.500 270.400 269.100 307.600 ;
        RECT 278.100 302.400 278.700 309.600 ;
        RECT 279.600 307.600 280.400 308.400 ;
        RECT 282.800 307.600 283.600 308.400 ;
        RECT 287.600 307.600 288.400 308.400 ;
        RECT 294.000 307.600 294.800 308.400 ;
        RECT 290.800 305.600 291.600 306.400 ;
        RECT 289.200 303.600 290.000 304.400 ;
        RECT 278.000 301.600 278.800 302.400 ;
        RECT 270.000 291.600 270.800 292.400 ;
        RECT 274.800 284.200 275.600 297.800 ;
        RECT 276.400 284.200 277.200 297.800 ;
        RECT 278.000 286.200 278.800 297.800 ;
        RECT 279.600 293.600 280.400 294.400 ;
        RECT 279.700 292.400 280.300 293.600 ;
        RECT 279.600 291.600 280.400 292.400 ;
        RECT 281.200 286.200 282.000 297.800 ;
        RECT 282.800 295.600 283.600 296.400 ;
        RECT 284.400 286.200 285.200 297.800 ;
        RECT 286.000 284.200 286.800 297.800 ;
        RECT 287.600 284.200 288.400 297.800 ;
        RECT 289.200 284.200 290.000 297.800 ;
        RECT 290.900 292.400 291.500 305.600 ;
        RECT 294.100 298.400 294.700 307.600 ;
        RECT 294.000 297.600 294.800 298.400 ;
        RECT 294.000 293.600 294.800 294.400 ;
        RECT 290.800 291.600 291.600 292.400 ;
        RECT 292.400 289.600 293.200 290.400 ;
        RECT 290.800 287.600 291.600 288.400 ;
        RECT 276.400 281.600 277.200 282.400 ;
        RECT 276.500 270.400 277.100 281.600 ;
        RECT 279.600 279.600 280.400 280.400 ;
        RECT 289.200 279.600 290.000 280.400 ;
        RECT 279.700 272.400 280.300 279.600 ;
        RECT 278.000 271.600 278.800 272.400 ;
        RECT 279.600 271.600 280.400 272.400 ;
        RECT 287.600 272.300 288.400 272.400 ;
        RECT 286.100 271.700 288.400 272.300 ;
        RECT 278.100 270.400 278.700 271.600 ;
        RECT 286.100 270.400 286.700 271.700 ;
        RECT 287.600 271.600 288.400 271.700 ;
        RECT 266.800 270.300 267.600 270.400 ;
        RECT 265.300 269.700 267.600 270.300 ;
        RECT 266.800 269.600 267.600 269.700 ;
        RECT 268.400 269.600 269.200 270.400 ;
        RECT 276.400 269.600 277.200 270.400 ;
        RECT 278.000 269.600 278.800 270.400 ;
        RECT 286.000 269.600 286.800 270.400 ;
        RECT 287.600 269.600 288.400 270.400 ;
        RECT 263.600 265.600 264.400 266.400 ;
        RECT 266.900 264.400 267.500 269.600 ;
        RECT 270.000 267.600 270.800 268.400 ;
        RECT 270.100 266.400 270.700 267.600 ;
        RECT 270.000 265.600 270.800 266.400 ;
        RECT 266.800 263.600 267.600 264.400 ;
        RECT 266.900 258.400 267.500 263.600 ;
        RECT 247.600 255.600 248.400 256.400 ;
        RECT 225.200 251.600 226.000 252.400 ;
        RECT 239.600 251.600 240.400 252.400 ;
        RECT 242.800 251.600 243.600 252.400 ;
        RECT 247.600 251.600 248.400 252.400 ;
        RECT 258.800 251.600 259.600 252.400 ;
        RECT 258.900 248.400 259.500 251.600 ;
        RECT 244.400 247.600 245.200 248.400 ;
        RECT 258.800 247.600 259.600 248.400 ;
        RECT 244.500 244.400 245.100 247.600 ;
        RECT 226.800 243.600 227.600 244.400 ;
        RECT 244.400 243.600 245.200 244.400 ;
        RECT 250.800 243.600 251.600 244.400 ;
        RECT 260.400 244.200 261.200 257.800 ;
        RECT 262.000 244.200 262.800 257.800 ;
        RECT 263.600 244.200 264.400 257.800 ;
        RECT 265.200 246.200 266.000 257.800 ;
        RECT 266.800 257.600 267.600 258.400 ;
        RECT 266.800 255.600 267.600 256.400 ;
        RECT 268.400 246.200 269.200 257.800 ;
        RECT 270.000 257.600 270.800 258.400 ;
        RECT 270.100 254.400 270.700 257.600 ;
        RECT 270.000 253.600 270.800 254.400 ;
        RECT 271.600 246.200 272.400 257.800 ;
        RECT 273.200 244.200 274.000 257.800 ;
        RECT 274.800 244.200 275.600 257.800 ;
        RECT 220.400 241.600 221.200 242.400 ;
        RECT 220.500 238.400 221.100 241.600 ;
        RECT 226.900 238.400 227.500 243.600 ;
        RECT 186.800 237.600 187.600 238.400 ;
        RECT 193.200 237.600 194.000 238.400 ;
        RECT 185.200 227.600 186.000 228.400 ;
        RECT 185.300 226.400 185.900 227.600 ;
        RECT 185.200 225.600 186.000 226.400 ;
        RECT 196.400 224.200 197.200 237.800 ;
        RECT 198.000 224.200 198.800 237.800 ;
        RECT 199.600 224.200 200.400 235.800 ;
        RECT 201.200 227.600 202.000 228.400 ;
        RECT 201.300 222.400 201.900 227.600 ;
        RECT 202.800 224.200 203.600 235.800 ;
        RECT 204.400 225.600 205.200 226.400 ;
        RECT 201.200 221.600 202.000 222.400 ;
        RECT 150.000 217.600 150.800 218.400 ;
        RECT 150.100 216.400 150.700 217.600 ;
        RECT 150.000 215.600 150.800 216.400 ;
        RECT 143.600 213.600 144.400 214.400 ;
        RECT 148.400 211.600 149.200 212.400 ;
        RECT 148.500 210.400 149.100 211.600 ;
        RECT 148.400 209.600 149.200 210.400 ;
        RECT 145.200 207.600 146.000 208.400 ;
        RECT 145.300 198.400 145.900 207.600 ;
        RECT 151.600 206.200 152.400 217.800 ;
        RECT 166.000 217.600 166.800 218.400 ;
        RECT 172.400 217.600 173.200 218.400 ;
        RECT 154.800 210.200 155.600 215.800 ;
        RECT 158.000 215.600 158.800 216.400 ;
        RECT 158.100 198.400 158.700 215.600 ;
        RECT 167.600 215.000 168.400 215.800 ;
        RECT 169.000 215.000 173.200 215.600 ;
        RECT 174.200 215.000 175.000 215.800 ;
        RECT 164.400 213.600 165.200 214.400 ;
        RECT 166.000 213.600 166.800 214.400 ;
        RECT 167.600 214.200 168.200 215.000 ;
        RECT 169.000 214.800 169.800 215.000 ;
        RECT 172.400 214.800 173.200 215.000 ;
        RECT 167.600 213.600 172.400 214.200 ;
        RECT 164.400 211.600 165.200 212.400 ;
        RECT 164.500 198.400 165.100 211.600 ;
        RECT 166.100 208.400 166.700 213.600 ;
        RECT 167.600 210.200 168.200 213.600 ;
        RECT 171.600 213.400 172.400 213.600 ;
        RECT 174.400 210.200 175.000 215.000 ;
        RECT 175.600 213.600 176.400 214.400 ;
        RECT 167.600 209.400 168.400 210.200 ;
        RECT 174.200 209.400 175.000 210.200 ;
        RECT 166.000 207.600 166.800 208.400 ;
        RECT 178.800 203.600 179.600 204.400 ;
        RECT 188.400 204.200 189.200 217.800 ;
        RECT 190.000 204.200 190.800 217.800 ;
        RECT 191.600 204.200 192.400 217.800 ;
        RECT 193.200 206.200 194.000 217.800 ;
        RECT 194.800 215.600 195.600 216.400 ;
        RECT 196.400 206.200 197.200 217.800 ;
        RECT 198.000 217.600 198.800 218.400 ;
        RECT 198.100 214.400 198.700 217.600 ;
        RECT 198.000 213.600 198.800 214.400 ;
        RECT 199.600 206.200 200.400 217.800 ;
        RECT 201.200 204.200 202.000 217.800 ;
        RECT 202.800 204.200 203.600 217.800 ;
        RECT 204.500 216.400 205.100 225.600 ;
        RECT 206.000 224.200 206.800 235.800 ;
        RECT 207.600 224.200 208.400 237.800 ;
        RECT 209.200 224.200 210.000 237.800 ;
        RECT 210.800 224.200 211.600 237.800 ;
        RECT 220.400 237.600 221.200 238.400 ;
        RECT 226.800 237.600 227.600 238.400 ;
        RECT 212.400 229.600 213.200 230.400 ;
        RECT 209.200 221.600 210.000 222.400 ;
        RECT 204.400 215.600 205.200 216.400 ;
        RECT 204.400 211.600 205.200 212.400 ;
        RECT 142.000 197.600 142.800 198.400 ;
        RECT 145.200 197.600 146.000 198.400 ;
        RECT 158.000 197.600 158.800 198.400 ;
        RECT 161.200 197.600 162.000 198.400 ;
        RECT 164.400 197.600 165.200 198.400 ;
        RECT 138.800 189.600 139.600 190.400 ;
        RECT 151.600 189.600 152.400 190.400 ;
        RECT 159.600 189.600 160.400 190.400 ;
        RECT 138.900 180.400 139.500 189.600 ;
        RECT 159.700 186.400 160.300 189.600 ;
        RECT 161.300 188.400 161.900 197.600 ;
        RECT 162.600 191.800 163.400 192.600 ;
        RECT 169.200 191.800 170.000 192.600 ;
        RECT 161.200 187.600 162.000 188.400 ;
        RECT 162.600 187.000 163.200 191.800 ;
        RECT 165.200 188.400 166.000 188.600 ;
        RECT 169.400 188.400 170.000 191.800 ;
        RECT 170.800 189.600 171.600 190.400 ;
        RECT 172.400 189.600 173.200 190.400 ;
        RECT 170.900 188.400 171.500 189.600 ;
        RECT 172.500 188.400 173.100 189.600 ;
        RECT 165.200 187.800 170.000 188.400 ;
        RECT 164.400 187.000 165.200 187.200 ;
        RECT 167.800 187.000 168.600 187.200 ;
        RECT 169.400 187.000 170.000 187.800 ;
        RECT 170.800 187.600 171.600 188.400 ;
        RECT 172.400 187.600 173.200 188.400 ;
        RECT 146.800 185.600 147.600 186.400 ;
        RECT 150.000 185.600 150.800 186.400 ;
        RECT 159.600 185.600 160.400 186.400 ;
        RECT 162.600 186.200 163.400 187.000 ;
        RECT 164.400 186.400 168.600 187.000 ;
        RECT 169.200 186.200 170.000 187.000 ;
        RECT 177.200 185.600 178.000 186.400 ;
        RECT 145.200 183.600 146.000 184.400 ;
        RECT 138.800 179.600 139.600 180.400 ;
        RECT 145.300 176.400 145.900 183.600 ;
        RECT 146.900 176.400 147.500 185.600 ;
        RECT 156.400 183.600 157.200 184.400 ;
        RECT 137.200 175.600 138.000 176.400 ;
        RECT 145.200 175.600 146.000 176.400 ;
        RECT 146.800 175.600 147.600 176.400 ;
        RECT 156.500 172.400 157.100 183.600 ;
        RECT 135.600 171.600 136.400 172.400 ;
        RECT 140.400 171.600 141.200 172.400 ;
        RECT 156.400 171.600 157.200 172.400 ;
        RECT 135.700 168.400 136.300 171.600 ;
        RECT 137.200 169.600 138.000 170.400 ;
        RECT 135.600 167.600 136.400 168.400 ;
        RECT 137.300 158.400 137.900 169.600 ;
        RECT 142.000 165.600 142.800 166.400 ;
        RECT 151.600 165.600 152.400 166.400 ;
        RECT 138.800 163.600 139.600 164.400 ;
        RECT 140.400 163.600 141.200 164.400 ;
        RECT 137.200 157.600 138.000 158.400 ;
        RECT 122.800 155.600 123.600 156.400 ;
        RECT 134.000 155.600 134.800 156.400 ;
        RECT 119.700 151.700 121.900 152.300 ;
        RECT 118.000 149.600 118.800 150.400 ;
        RECT 119.600 149.600 120.400 150.400 ;
        RECT 119.700 146.400 120.300 149.600 ;
        RECT 121.300 148.400 121.900 151.700 ;
        RECT 122.900 148.400 123.500 155.600 ;
        RECT 129.200 153.600 130.000 154.400 ;
        RECT 127.600 152.300 128.400 152.400 ;
        RECT 126.100 151.700 128.400 152.300 ;
        RECT 124.400 149.600 125.200 150.400 ;
        RECT 124.500 148.400 125.100 149.600 ;
        RECT 121.200 147.600 122.000 148.400 ;
        RECT 122.800 147.600 123.600 148.400 ;
        RECT 124.400 147.600 125.200 148.400 ;
        RECT 119.600 145.600 120.400 146.400 ;
        RECT 122.800 145.600 123.600 146.400 ;
        RECT 122.900 138.400 123.500 145.600 ;
        RECT 113.200 129.600 114.000 130.400 ;
        RECT 113.300 116.400 113.900 129.600 ;
        RECT 114.800 126.200 115.600 137.800 ;
        RECT 122.800 137.600 123.600 138.400 ;
        RECT 121.200 133.600 122.000 134.400 ;
        RECT 121.300 126.400 121.900 133.600 ;
        RECT 124.500 132.400 125.100 147.600 ;
        RECT 126.100 146.400 126.700 151.700 ;
        RECT 127.600 151.600 128.400 151.700 ;
        RECT 127.600 149.600 128.400 150.400 ;
        RECT 129.300 150.300 129.900 153.600 ;
        RECT 130.800 151.600 131.600 152.400 ;
        RECT 134.000 151.600 134.800 152.400 ;
        RECT 130.800 150.300 131.600 150.400 ;
        RECT 129.300 149.700 131.600 150.300 ;
        RECT 130.800 149.600 131.600 149.700 ;
        RECT 127.600 147.600 128.400 148.400 ;
        RECT 134.100 146.400 134.700 151.600 ;
        RECT 137.200 149.600 138.000 150.400 ;
        RECT 137.300 148.400 137.900 149.600 ;
        RECT 135.600 147.600 136.400 148.400 ;
        RECT 137.200 147.600 138.000 148.400 ;
        RECT 126.000 145.600 126.800 146.400 ;
        RECT 134.000 145.600 134.800 146.400 ;
        RECT 135.700 144.400 136.300 147.600 ;
        RECT 135.600 143.600 136.400 144.400 ;
        RECT 129.200 139.600 130.000 140.400 ;
        RECT 126.000 135.600 126.800 136.400 ;
        RECT 124.400 131.600 125.200 132.400 ;
        RECT 124.400 129.600 125.200 130.400 ;
        RECT 121.200 125.600 122.000 126.400 ;
        RECT 126.100 124.400 126.700 135.600 ;
        RECT 129.300 134.400 129.900 139.600 ;
        RECT 138.900 138.300 139.500 163.600 ;
        RECT 140.500 160.400 141.100 163.600 ;
        RECT 140.400 159.600 141.200 160.400 ;
        RECT 140.500 156.400 141.100 159.600 ;
        RECT 140.400 155.600 141.200 156.400 ;
        RECT 140.400 151.600 141.200 152.400 ;
        RECT 140.500 146.400 141.100 151.600 ;
        RECT 142.100 148.400 142.700 165.600 ;
        RECT 161.200 164.200 162.000 177.800 ;
        RECT 162.800 164.200 163.600 177.800 ;
        RECT 164.400 164.200 165.200 177.800 ;
        RECT 166.000 166.200 166.800 177.800 ;
        RECT 167.600 175.600 168.400 176.400 ;
        RECT 167.700 168.400 168.300 175.600 ;
        RECT 167.600 167.600 168.400 168.400 ;
        RECT 169.200 166.200 170.000 177.800 ;
        RECT 170.800 173.600 171.600 174.400 ;
        RECT 161.200 161.600 162.000 162.400 ;
        RECT 151.600 157.600 152.400 158.400 ;
        RECT 146.800 151.800 147.600 152.600 ;
        RECT 153.400 151.800 154.200 152.600 ;
        RECT 146.800 148.400 147.400 151.800 ;
        RECT 150.800 148.400 151.600 148.600 ;
        RECT 142.000 147.600 142.800 148.400 ;
        RECT 146.800 147.800 151.600 148.400 ;
        RECT 140.400 145.600 141.200 146.400 ;
        RECT 138.900 137.700 141.100 138.300 ;
        RECT 138.800 135.600 139.600 136.400 ;
        RECT 140.500 134.400 141.100 137.700 ;
        RECT 142.100 134.400 142.700 147.600 ;
        RECT 146.800 147.000 147.400 147.800 ;
        RECT 148.200 147.000 149.000 147.200 ;
        RECT 151.600 147.000 152.400 147.200 ;
        RECT 153.600 147.000 154.200 151.800 ;
        RECT 154.800 147.600 155.600 148.400 ;
        RECT 146.800 146.200 147.600 147.000 ;
        RECT 148.200 146.400 152.400 147.000 ;
        RECT 148.400 145.600 149.200 146.400 ;
        RECT 153.400 146.200 154.200 147.000 ;
        RECT 143.600 143.600 144.400 144.400 ;
        RECT 143.700 140.400 144.300 143.600 ;
        RECT 143.600 139.600 144.400 140.400 ;
        RECT 127.600 133.600 128.400 134.400 ;
        RECT 129.200 133.600 130.000 134.400 ;
        RECT 134.000 133.600 134.800 134.400 ;
        RECT 140.400 133.600 141.200 134.400 ;
        RECT 142.000 133.600 142.800 134.400 ;
        RECT 150.000 133.600 150.800 134.400 ;
        RECT 135.600 131.600 136.400 132.400 ;
        RECT 142.000 131.600 142.800 132.400 ;
        RECT 145.200 131.600 146.000 132.400 ;
        RECT 132.400 129.600 133.200 130.400 ;
        RECT 134.000 129.600 134.800 130.400 ;
        RECT 138.800 129.600 139.600 130.400 ;
        RECT 145.200 130.300 146.000 130.400 ;
        RECT 143.700 129.700 146.000 130.300 ;
        RECT 130.800 127.600 131.600 128.400 ;
        RECT 119.600 123.600 120.400 124.400 ;
        RECT 126.000 123.600 126.800 124.400 ;
        RECT 132.500 124.300 133.100 129.600 ;
        RECT 130.900 123.700 133.100 124.300 ;
        RECT 113.200 115.600 114.000 116.400 ;
        RECT 118.000 115.600 118.800 116.400 ;
        RECT 113.200 111.600 114.000 112.400 ;
        RECT 98.800 109.600 99.600 110.400 ;
        RECT 100.400 109.600 101.200 110.400 ;
        RECT 110.000 109.600 110.800 110.400 ;
        RECT 113.300 108.400 113.900 111.600 ;
        RECT 118.100 110.400 118.700 115.600 ;
        RECT 119.600 113.600 120.400 114.400 ;
        RECT 119.700 112.400 120.300 113.600 ;
        RECT 119.600 111.600 120.400 112.400 ;
        RECT 121.200 111.600 122.000 112.400 ;
        RECT 127.600 111.600 128.400 112.400 ;
        RECT 121.300 110.400 121.900 111.600 ;
        RECT 118.000 109.600 118.800 110.400 ;
        RECT 121.200 110.300 122.000 110.400 ;
        RECT 121.200 109.700 123.500 110.300 ;
        RECT 121.200 109.600 122.000 109.700 ;
        RECT 97.200 107.600 98.000 108.400 ;
        RECT 100.400 108.300 101.200 108.400 ;
        RECT 98.900 107.700 101.200 108.300 ;
        RECT 97.300 98.400 97.900 107.600 ;
        RECT 97.200 97.600 98.000 98.400 ;
        RECT 97.200 93.600 98.000 94.400 ;
        RECT 90.800 89.600 91.600 90.400 ;
        RECT 94.000 89.600 94.800 90.400 ;
        RECT 90.900 84.400 91.500 89.600 ;
        RECT 94.100 88.400 94.700 89.600 ;
        RECT 94.000 87.600 94.800 88.400 ;
        RECT 90.800 83.600 91.600 84.400 ;
        RECT 90.800 69.600 91.600 70.400 ;
        RECT 92.400 69.600 93.200 70.400 ;
        RECT 90.900 68.400 91.500 69.600 ;
        RECT 92.500 68.400 93.100 69.600 ;
        RECT 90.800 67.600 91.600 68.400 ;
        RECT 92.400 67.600 93.200 68.400 ;
        RECT 89.200 61.600 90.000 62.400 ;
        RECT 63.600 51.600 64.400 52.400 ;
        RECT 68.400 51.600 69.200 52.400 ;
        RECT 71.600 51.600 72.400 52.400 ;
        RECT 76.400 51.600 77.200 52.400 ;
        RECT 78.000 51.600 78.800 52.400 ;
        RECT 86.000 51.600 86.800 52.400 ;
        RECT 87.600 51.600 88.400 52.400 ;
        RECT 65.200 43.600 66.000 44.400 ;
        RECT 63.600 35.600 64.400 36.400 ;
        RECT 62.000 33.600 62.800 34.400 ;
        RECT 55.600 31.600 56.400 32.400 ;
        RECT 44.400 30.300 45.200 30.400 ;
        RECT 44.400 29.700 46.700 30.300 ;
        RECT 44.400 29.600 45.200 29.700 ;
        RECT 41.200 15.700 43.500 16.300 ;
        RECT 41.200 15.600 42.000 15.700 ;
        RECT 36.400 13.600 37.200 14.400 ;
        RECT 34.800 11.600 35.600 12.400 ;
        RECT 38.000 11.600 38.800 12.400 ;
        RECT 41.300 10.400 41.900 15.600 ;
        RECT 42.800 13.600 43.600 14.400 ;
        RECT 46.100 12.400 46.700 29.700 ;
        RECT 52.400 29.600 53.200 30.400 ;
        RECT 60.400 29.600 61.200 30.400 ;
        RECT 62.100 28.400 62.700 33.600 ;
        RECT 65.300 30.400 65.900 43.600 ;
        RECT 68.500 38.300 69.100 51.600 ;
        RECT 71.600 49.600 72.400 50.400 ;
        RECT 79.600 43.600 80.400 44.400 ;
        RECT 68.500 37.700 70.700 38.300 ;
        RECT 65.200 29.600 66.000 30.400 ;
        RECT 50.800 27.600 51.600 28.400 ;
        RECT 62.000 27.600 62.800 28.400 ;
        RECT 50.900 18.400 51.500 27.600 ;
        RECT 57.200 23.600 58.000 24.400 ;
        RECT 68.400 24.200 69.200 35.800 ;
        RECT 70.100 32.400 70.700 37.700 ;
        RECT 70.000 31.600 70.800 32.400 ;
        RECT 76.400 31.600 77.200 32.400 ;
        RECT 54.000 19.600 54.800 20.400 ;
        RECT 50.800 17.600 51.600 18.400 ;
        RECT 46.000 11.600 46.800 12.400 ;
        RECT 41.200 9.600 42.000 10.400 ;
        RECT 52.400 10.200 53.200 15.800 ;
        RECT 54.100 14.400 54.700 19.600 ;
        RECT 54.000 13.600 54.800 14.400 ;
        RECT 55.600 6.200 56.400 17.800 ;
        RECT 57.300 12.600 57.900 23.600 ;
        RECT 70.100 18.400 70.700 31.600 ;
        RECT 76.500 30.200 77.100 31.600 ;
        RECT 76.400 29.400 77.200 30.200 ;
        RECT 76.400 25.600 77.200 26.400 ;
        RECT 76.500 20.400 77.100 25.600 ;
        RECT 78.000 24.200 78.800 35.800 ;
        RECT 76.400 19.600 77.200 20.400 ;
        RECT 57.200 11.800 58.000 12.600 ;
        RECT 65.200 6.200 66.000 17.800 ;
        RECT 70.000 17.600 70.800 18.400 ;
        RECT 73.200 17.600 74.000 18.400 ;
        RECT 78.000 15.600 78.800 16.400 ;
        RECT 78.100 14.400 78.700 15.600 ;
        RECT 78.000 13.600 78.800 14.400 ;
        RECT 79.700 12.400 80.300 43.600 ;
        RECT 82.800 33.600 83.600 34.400 ;
        RECT 81.200 26.200 82.000 31.800 ;
        RECT 82.900 28.400 83.500 33.600 ;
        RECT 84.400 31.600 85.200 32.400 ;
        RECT 84.400 29.600 85.200 30.400 ;
        RECT 82.800 27.600 83.600 28.400 ;
        RECT 82.900 16.400 83.500 27.600 ;
        RECT 86.100 24.400 86.700 51.600 ;
        RECT 87.700 50.400 88.300 51.600 ;
        RECT 87.600 49.600 88.400 50.400 ;
        RECT 90.900 46.400 91.500 67.600 ;
        RECT 92.500 66.400 93.100 67.600 ;
        RECT 92.400 65.600 93.200 66.400 ;
        RECT 97.300 58.400 97.900 93.600 ;
        RECT 98.900 90.300 99.500 107.700 ;
        RECT 100.400 107.600 101.200 107.700 ;
        RECT 102.000 107.600 102.800 108.400 ;
        RECT 108.400 107.600 109.200 108.400 ;
        RECT 113.200 107.600 114.000 108.400 ;
        RECT 114.800 107.600 115.600 108.400 ;
        RECT 121.200 107.600 122.000 108.400 ;
        RECT 108.500 106.400 109.100 107.600 ;
        RECT 108.400 105.600 109.200 106.400 ;
        RECT 114.900 98.400 115.500 107.600 ;
        RECT 121.300 98.400 121.900 107.600 ;
        RECT 114.800 97.600 115.600 98.400 ;
        RECT 121.200 97.600 122.000 98.400 ;
        RECT 105.200 95.600 106.000 96.400 ;
        RECT 113.200 95.600 114.000 96.400 ;
        RECT 102.000 93.600 102.800 94.400 ;
        RECT 100.400 91.600 101.200 92.400 ;
        RECT 98.900 89.700 101.100 90.300 ;
        RECT 98.800 81.600 99.600 82.400 ;
        RECT 98.900 70.400 99.500 81.600 ;
        RECT 100.500 78.400 101.100 89.700 ;
        RECT 102.100 86.300 102.700 93.600 ;
        RECT 105.300 92.400 105.900 95.600 ;
        RECT 119.600 93.600 120.400 94.400 ;
        RECT 105.200 91.600 106.000 92.400 ;
        RECT 110.000 91.600 110.800 92.400 ;
        RECT 118.000 91.600 118.800 92.400 ;
        RECT 110.100 90.400 110.700 91.600 ;
        RECT 103.600 89.600 104.400 90.400 ;
        RECT 106.800 89.600 107.600 90.400 ;
        RECT 110.000 89.600 110.800 90.400 ;
        RECT 111.600 89.600 112.400 90.400 ;
        RECT 114.800 89.600 115.600 90.400 ;
        RECT 121.200 89.600 122.000 90.400 ;
        RECT 103.700 88.400 104.300 89.600 ;
        RECT 106.900 88.400 107.500 89.600 ;
        RECT 114.900 88.400 115.500 89.600 ;
        RECT 103.600 87.600 104.400 88.400 ;
        RECT 106.800 87.600 107.600 88.400 ;
        RECT 108.400 87.600 109.200 88.400 ;
        RECT 114.800 87.600 115.600 88.400 ;
        RECT 102.100 85.700 104.300 86.300 ;
        RECT 103.700 78.400 104.300 85.700 ;
        RECT 106.800 85.600 107.600 86.400 ;
        RECT 106.900 78.400 107.500 85.600 ;
        RECT 122.900 82.400 123.500 109.700 ;
        RECT 127.700 108.400 128.300 111.600 ;
        RECT 127.600 107.600 128.400 108.400 ;
        RECT 124.400 105.600 125.200 106.400 ;
        RECT 129.200 103.600 130.000 104.400 ;
        RECT 124.400 93.600 125.200 94.400 ;
        RECT 127.600 93.600 128.400 94.400 ;
        RECT 124.500 88.400 125.100 93.600 ;
        RECT 126.000 91.600 126.800 92.400 ;
        RECT 124.400 87.600 125.200 88.400 ;
        RECT 126.100 84.300 126.700 91.600 ;
        RECT 124.500 83.700 126.700 84.300 ;
        RECT 122.800 81.600 123.600 82.400 ;
        RECT 100.400 77.600 101.200 78.400 ;
        RECT 103.600 77.600 104.400 78.400 ;
        RECT 106.800 77.600 107.600 78.400 ;
        RECT 98.800 69.600 99.600 70.400 ;
        RECT 100.400 67.600 101.200 68.400 ;
        RECT 98.800 65.600 99.600 66.400 ;
        RECT 98.900 64.400 99.500 65.600 ;
        RECT 98.800 63.600 99.600 64.400 ;
        RECT 100.500 58.400 101.100 67.600 ;
        RECT 102.000 65.600 102.800 66.400 ;
        RECT 105.200 65.600 106.000 66.400 ;
        RECT 108.400 65.600 109.200 66.400 ;
        RECT 105.300 58.400 105.900 65.600 ;
        RECT 108.500 64.400 109.100 65.600 ;
        RECT 108.400 63.600 109.200 64.400 ;
        RECT 113.200 64.200 114.000 75.800 ;
        RECT 119.600 73.600 120.400 74.400 ;
        RECT 119.700 70.400 120.300 73.600 ;
        RECT 121.200 71.600 122.000 72.400 ;
        RECT 119.600 69.600 120.400 70.400 ;
        RECT 118.000 67.600 118.800 68.400 ;
        RECT 92.400 57.600 93.200 58.400 ;
        RECT 97.200 57.600 98.000 58.400 ;
        RECT 100.400 57.600 101.200 58.400 ;
        RECT 105.200 57.600 106.000 58.400 ;
        RECT 92.500 52.400 93.100 57.600 ;
        RECT 95.600 55.600 96.400 56.400 ;
        RECT 111.600 55.600 112.400 56.400 ;
        RECT 119.600 55.600 120.400 56.400 ;
        RECT 95.700 54.400 96.300 55.600 ;
        RECT 111.700 54.400 112.300 55.600 ;
        RECT 95.600 53.600 96.400 54.400 ;
        RECT 111.600 53.600 112.400 54.400 ;
        RECT 119.700 52.400 120.300 55.600 ;
        RECT 121.300 52.400 121.900 71.600 ;
        RECT 122.800 64.200 123.600 75.800 ;
        RECT 124.500 52.400 125.100 83.700 ;
        RECT 127.700 78.400 128.300 93.600 ;
        RECT 129.300 92.400 129.900 103.600 ;
        RECT 129.200 91.600 130.000 92.400 ;
        RECT 130.900 90.400 131.500 123.700 ;
        RECT 134.100 118.400 134.700 129.600 ;
        RECT 138.900 128.400 139.500 129.600 ;
        RECT 138.800 127.600 139.600 128.400 ;
        RECT 135.600 125.600 136.400 126.400 ;
        RECT 134.000 117.600 134.800 118.400 ;
        RECT 135.700 114.400 136.300 125.600 ;
        RECT 142.000 123.600 142.800 124.400 ;
        RECT 135.600 113.600 136.400 114.400 ;
        RECT 142.100 114.300 142.700 123.600 ;
        RECT 140.500 113.700 142.700 114.300 ;
        RECT 135.700 112.400 136.300 113.600 ;
        RECT 132.400 111.600 133.200 112.400 ;
        RECT 135.600 111.600 136.400 112.400 ;
        RECT 132.500 108.400 133.100 111.600 ;
        RECT 140.500 110.400 141.100 113.700 ;
        RECT 142.000 111.600 142.800 112.400 ;
        RECT 140.400 109.600 141.200 110.400 ;
        RECT 142.000 109.600 142.800 110.400 ;
        RECT 132.400 107.600 133.200 108.400 ;
        RECT 137.200 107.600 138.000 108.400 ;
        RECT 140.400 107.600 141.200 108.400 ;
        RECT 132.500 96.400 133.100 107.600 ;
        RECT 137.300 100.400 137.900 107.600 ;
        RECT 137.200 99.600 138.000 100.400 ;
        RECT 140.500 98.400 141.100 107.600 ;
        RECT 143.700 98.400 144.300 129.700 ;
        RECT 145.200 129.600 146.000 129.700 ;
        RECT 146.800 129.600 147.600 130.400 ;
        RECT 150.100 124.400 150.700 133.600 ;
        RECT 154.900 128.400 155.500 147.600 ;
        RECT 161.300 138.400 161.900 161.600 ;
        RECT 170.900 160.400 171.500 173.600 ;
        RECT 172.400 166.200 173.200 177.800 ;
        RECT 174.000 164.200 174.800 177.800 ;
        RECT 175.600 164.200 176.400 177.800 ;
        RECT 177.300 168.400 177.900 185.600 ;
        RECT 178.900 176.400 179.500 203.600 ;
        RECT 182.000 189.600 182.800 190.400 ;
        RECT 178.800 175.600 179.600 176.400 ;
        RECT 182.100 172.400 182.700 189.600 ;
        RECT 183.600 184.200 184.400 197.800 ;
        RECT 185.200 184.200 186.000 197.800 ;
        RECT 186.800 184.200 187.600 197.800 ;
        RECT 188.400 184.200 189.200 195.800 ;
        RECT 190.000 185.600 190.800 186.400 ;
        RECT 191.600 184.200 192.400 195.800 ;
        RECT 193.200 187.600 194.000 188.400 ;
        RECT 194.800 184.200 195.600 195.800 ;
        RECT 196.400 184.200 197.200 197.800 ;
        RECT 198.000 184.200 198.800 197.800 ;
        RECT 199.600 191.600 200.400 192.400 ;
        RECT 190.000 181.600 190.800 182.400 ;
        RECT 185.200 173.600 186.000 174.400 ;
        RECT 185.300 172.400 185.900 173.600 ;
        RECT 190.100 172.400 190.700 181.600 ;
        RECT 193.200 177.600 194.000 178.400 ;
        RECT 194.800 175.600 195.600 176.400 ;
        RECT 194.900 174.400 195.500 175.600 ;
        RECT 193.200 173.600 194.000 174.400 ;
        RECT 194.800 173.600 195.600 174.400 ;
        RECT 180.400 171.600 181.200 172.400 ;
        RECT 182.000 171.600 182.800 172.400 ;
        RECT 185.200 171.600 186.000 172.400 ;
        RECT 190.000 171.600 190.800 172.400 ;
        RECT 177.200 167.600 178.000 168.400 ;
        RECT 170.800 159.600 171.600 160.400 ;
        RECT 169.200 144.200 170.000 157.800 ;
        RECT 170.800 144.200 171.600 157.800 ;
        RECT 172.400 144.200 173.200 155.800 ;
        RECT 174.000 147.600 174.800 148.400 ;
        RECT 175.600 144.200 176.400 155.800 ;
        RECT 177.300 146.400 177.900 167.600 ;
        RECT 177.200 145.600 178.000 146.400 ;
        RECT 177.300 142.400 177.900 145.600 ;
        RECT 178.800 144.200 179.600 155.800 ;
        RECT 180.400 144.200 181.200 157.800 ;
        RECT 182.000 144.200 182.800 157.800 ;
        RECT 183.600 144.200 184.400 157.800 ;
        RECT 185.200 149.600 186.000 150.400 ;
        RECT 177.200 141.600 178.000 142.400 ;
        RECT 180.400 141.600 181.200 142.400 ;
        RECT 156.400 137.600 157.200 138.400 ;
        RECT 161.200 137.600 162.000 138.400 ;
        RECT 156.500 134.400 157.100 137.600 ;
        RECT 158.000 135.600 158.800 136.400 ;
        RECT 156.400 133.600 157.200 134.400 ;
        RECT 158.100 132.400 158.700 135.600 ;
        RECT 156.400 131.600 157.200 132.400 ;
        RECT 158.000 131.600 158.800 132.400 ;
        RECT 153.200 127.600 154.000 128.400 ;
        RECT 154.800 127.600 155.600 128.400 ;
        RECT 153.300 124.400 153.900 127.600 ;
        RECT 146.800 123.600 147.600 124.400 ;
        RECT 150.000 123.600 150.800 124.400 ;
        RECT 153.200 123.600 154.000 124.400 ;
        RECT 145.200 109.600 146.000 110.400 ;
        RECT 146.900 110.300 147.500 123.600 ;
        RECT 156.500 118.400 157.100 131.600 ;
        RECT 161.200 129.600 162.000 130.400 ;
        RECT 161.300 128.400 161.900 129.600 ;
        RECT 161.200 127.600 162.000 128.400 ;
        RECT 158.000 123.600 158.800 124.400 ;
        RECT 164.400 123.600 165.200 124.400 ;
        RECT 174.000 124.200 174.800 137.800 ;
        RECT 175.600 124.200 176.400 137.800 ;
        RECT 177.200 124.200 178.000 137.800 ;
        RECT 178.800 126.200 179.600 137.800 ;
        RECT 180.500 136.400 181.100 141.600 ;
        RECT 185.300 140.400 185.900 149.600 ;
        RECT 185.200 139.600 186.000 140.400 ;
        RECT 180.400 135.600 181.200 136.400 ;
        RECT 156.400 117.600 157.200 118.400 ;
        RECT 150.000 111.600 150.800 112.400 ;
        RECT 153.200 111.600 154.000 112.400 ;
        RECT 146.900 109.700 149.100 110.300 ;
        RECT 145.300 104.400 145.900 109.600 ;
        RECT 146.800 107.600 147.600 108.400 ;
        RECT 145.200 103.600 146.000 104.400 ;
        RECT 140.400 97.600 141.200 98.400 ;
        RECT 143.600 97.600 144.400 98.400 ;
        RECT 132.400 95.600 133.200 96.400 ;
        RECT 135.600 94.300 136.400 94.400 ;
        RECT 134.100 93.700 136.400 94.300 ;
        RECT 132.400 91.600 133.200 92.400 ;
        RECT 130.800 89.600 131.600 90.400 ;
        RECT 132.500 88.400 133.100 91.600 ;
        RECT 132.400 87.600 133.200 88.400 ;
        RECT 130.800 83.600 131.600 84.400 ;
        RECT 134.100 84.300 134.700 93.700 ;
        RECT 135.600 93.600 136.400 93.700 ;
        RECT 145.200 93.600 146.000 94.400 ;
        RECT 135.600 91.600 136.400 92.400 ;
        RECT 137.200 91.600 138.000 92.400 ;
        RECT 135.700 88.400 136.300 91.600 ;
        RECT 140.400 89.600 141.200 90.400 ;
        RECT 142.000 89.600 142.800 90.400 ;
        RECT 140.500 88.400 141.100 89.600 ;
        RECT 135.600 87.600 136.400 88.400 ;
        RECT 140.400 87.600 141.200 88.400 ;
        RECT 132.500 83.700 134.700 84.300 ;
        RECT 127.600 77.600 128.400 78.400 ;
        RECT 130.900 76.400 131.500 83.600 ;
        RECT 132.500 78.400 133.100 83.700 ;
        RECT 132.400 77.600 133.200 78.400 ;
        RECT 130.800 75.600 131.600 76.400 ;
        RECT 126.000 66.200 126.800 71.800 ;
        RECT 134.000 69.600 134.800 70.400 ;
        RECT 129.200 65.600 130.000 66.400 ;
        RECT 130.800 65.600 131.600 66.400 ;
        RECT 129.300 52.400 129.900 65.600 ;
        RECT 92.400 51.600 93.200 52.400 ;
        RECT 94.000 51.600 94.800 52.400 ;
        RECT 113.200 51.600 114.000 52.400 ;
        RECT 119.600 51.600 120.400 52.400 ;
        RECT 121.200 51.600 122.000 52.400 ;
        RECT 124.400 51.600 125.200 52.400 ;
        RECT 129.200 51.600 130.000 52.400 ;
        RECT 87.600 45.600 88.400 46.400 ;
        RECT 90.800 45.600 91.600 46.400 ;
        RECT 86.000 24.300 86.800 24.400 ;
        RECT 84.500 23.700 86.800 24.300 ;
        RECT 82.800 15.600 83.600 16.400 ;
        RECT 82.800 13.600 83.600 14.400 ;
        RECT 78.000 11.600 78.800 12.400 ;
        RECT 79.600 11.600 80.400 12.400 ;
        RECT 84.500 10.400 85.100 23.700 ;
        RECT 86.000 23.600 86.800 23.700 ;
        RECT 87.700 12.400 88.300 45.600 ;
        RECT 90.800 43.600 91.600 44.400 ;
        RECT 89.200 35.600 90.000 36.400 ;
        RECT 89.300 32.400 89.900 35.600 ;
        RECT 89.200 31.600 90.000 32.400 ;
        RECT 90.900 30.400 91.500 43.600 ;
        RECT 92.500 32.400 93.100 51.600 ;
        RECT 100.400 43.600 101.200 44.400 ;
        RECT 92.400 31.600 93.200 32.400 ;
        RECT 90.800 29.600 91.600 30.400 ;
        RECT 92.400 29.600 93.200 30.400 ;
        RECT 89.200 27.600 90.000 28.400 ;
        RECT 94.000 27.600 94.800 28.400 ;
        RECT 89.300 14.400 89.900 27.600 ;
        RECT 95.600 26.200 96.400 31.800 ;
        RECT 90.800 23.600 91.600 24.400 ;
        RECT 98.800 24.200 99.600 35.800 ;
        RECT 100.500 28.400 101.100 43.600 ;
        RECT 113.300 38.400 113.900 51.600 ;
        RECT 124.500 50.400 125.100 51.600 ;
        RECT 124.400 49.600 125.200 50.400 ;
        RECT 118.000 43.600 118.800 44.400 ;
        RECT 126.000 43.600 126.800 44.400 ;
        RECT 113.200 37.600 114.000 38.400 ;
        RECT 113.300 36.400 113.900 37.600 ;
        RECT 102.000 31.600 102.800 32.400 ;
        RECT 102.100 30.400 102.700 31.600 ;
        RECT 102.000 29.600 102.800 30.400 ;
        RECT 100.400 27.600 101.200 28.400 ;
        RECT 90.900 18.400 91.500 23.600 ;
        RECT 100.500 20.400 101.100 27.600 ;
        RECT 108.400 24.200 109.200 35.800 ;
        RECT 113.200 35.600 114.000 36.400 ;
        RECT 114.800 33.600 115.600 34.400 ;
        RECT 114.900 28.400 115.500 33.600 ;
        RECT 116.400 31.600 117.200 32.400 ;
        RECT 116.400 30.300 117.200 30.400 ;
        RECT 118.100 30.300 118.700 43.600 ;
        RECT 121.200 35.600 122.000 36.400 ;
        RECT 121.300 32.400 121.900 35.600 ;
        RECT 121.200 31.600 122.000 32.400 ;
        RECT 126.100 30.400 126.700 43.600 ;
        RECT 127.600 33.600 128.400 34.400 ;
        RECT 116.400 29.700 118.700 30.300 ;
        RECT 116.400 29.600 117.200 29.700 ;
        RECT 124.400 29.600 125.200 30.400 ;
        RECT 126.000 29.600 126.800 30.400 ;
        RECT 127.700 28.400 128.300 33.600 ;
        RECT 129.300 32.400 129.900 51.600 ;
        RECT 130.900 36.400 131.500 65.600 ;
        RECT 135.700 52.400 136.300 87.600 ;
        RECT 143.600 85.600 144.400 86.400 ;
        RECT 138.800 81.600 139.600 82.400 ;
        RECT 137.200 63.600 138.000 64.400 ;
        RECT 135.600 51.600 136.400 52.400 ;
        RECT 137.300 50.400 137.900 63.600 ;
        RECT 138.900 52.400 139.500 81.600 ;
        RECT 143.700 72.300 144.300 85.600 ;
        RECT 145.300 74.400 145.900 93.600 ;
        RECT 148.500 88.400 149.100 109.700 ;
        RECT 150.100 92.400 150.700 111.600 ;
        RECT 153.300 110.400 153.900 111.600 ;
        RECT 158.100 110.400 158.700 123.600 ;
        RECT 164.500 112.400 165.100 123.600 ;
        RECT 180.500 120.400 181.100 135.600 ;
        RECT 182.000 126.200 182.800 137.800 ;
        RECT 183.600 133.600 184.400 134.400 ;
        RECT 183.600 131.600 184.400 132.400 ;
        RECT 170.800 119.600 171.600 120.400 ;
        RECT 180.400 119.600 181.200 120.400 ;
        RECT 170.900 118.400 171.500 119.600 ;
        RECT 170.800 117.600 171.600 118.400 ;
        RECT 183.700 114.300 184.300 131.600 ;
        RECT 185.200 126.200 186.000 137.800 ;
        RECT 186.800 124.200 187.600 137.800 ;
        RECT 188.400 124.200 189.200 137.800 ;
        RECT 190.100 136.400 190.700 171.600 ;
        RECT 191.600 169.600 192.400 170.400 ;
        RECT 191.700 162.400 192.300 169.600 ;
        RECT 191.600 161.600 192.400 162.400 ;
        RECT 193.300 158.400 193.900 173.600 ;
        RECT 199.700 170.400 200.300 191.600 ;
        RECT 204.500 190.400 205.100 211.600 ;
        RECT 209.300 198.400 209.900 221.600 ;
        RECT 212.500 212.400 213.100 229.600 ;
        RECT 225.200 225.600 226.000 226.400 ;
        RECT 217.200 223.600 218.000 224.400 ;
        RECT 220.400 223.600 221.200 224.400 ;
        RECT 239.600 224.200 240.400 237.800 ;
        RECT 241.200 224.200 242.000 237.800 ;
        RECT 242.800 224.200 243.600 235.800 ;
        RECT 244.500 230.400 245.100 243.600 ;
        RECT 244.400 229.600 245.200 230.400 ;
        RECT 244.400 227.600 245.200 228.400 ;
        RECT 244.400 223.600 245.200 224.400 ;
        RECT 246.000 224.200 246.800 235.800 ;
        RECT 247.600 225.600 248.400 226.400 ;
        RECT 212.400 211.600 213.200 212.400 ;
        RECT 215.600 211.600 216.400 212.400 ;
        RECT 209.200 197.600 210.000 198.400 ;
        RECT 217.300 194.400 217.900 223.600 ;
        RECT 244.500 218.400 245.100 223.600 ;
        RECT 247.700 218.400 248.300 225.600 ;
        RECT 249.200 224.200 250.000 235.800 ;
        RECT 250.800 224.200 251.600 237.800 ;
        RECT 252.400 224.200 253.200 237.800 ;
        RECT 254.000 224.200 254.800 237.800 ;
        RECT 266.800 231.600 267.600 232.400 ;
        RECT 271.600 231.600 272.400 232.400 ;
        RECT 266.900 230.400 267.500 231.600 ;
        RECT 276.500 230.400 277.100 269.600 ;
        RECT 284.400 267.600 285.200 268.400 ;
        RECT 286.000 267.600 286.800 268.400 ;
        RECT 284.500 266.400 285.100 267.600 ;
        RECT 278.000 265.600 278.800 266.400 ;
        RECT 284.400 265.600 285.200 266.400 ;
        RECT 278.100 240.400 278.700 265.600 ;
        RECT 281.200 263.600 282.000 264.400 ;
        RECT 281.300 242.300 281.900 263.600 ;
        RECT 286.000 257.600 286.800 258.400 ;
        RECT 287.700 256.400 288.300 269.600 ;
        RECT 284.400 255.600 285.200 256.400 ;
        RECT 287.600 255.600 288.400 256.400 ;
        RECT 284.500 254.400 285.100 255.600 ;
        RECT 284.400 253.600 285.200 254.400 ;
        RECT 286.000 252.300 286.800 252.400 ;
        RECT 279.700 241.700 281.900 242.300 ;
        RECT 284.500 251.700 286.800 252.300 ;
        RECT 278.000 239.600 278.800 240.400 ;
        RECT 279.700 232.400 280.300 241.700 ;
        RECT 279.600 231.600 280.400 232.400 ;
        RECT 255.600 229.600 256.400 230.400 ;
        RECT 265.200 229.600 266.000 230.400 ;
        RECT 266.800 229.600 267.600 230.400 ;
        RECT 276.400 229.600 277.200 230.400 ;
        RECT 282.800 230.300 283.600 230.400 ;
        RECT 284.500 230.300 285.100 251.700 ;
        RECT 286.000 251.600 286.800 251.700 ;
        RECT 286.000 249.600 286.800 250.400 ;
        RECT 286.100 238.400 286.700 249.600 ;
        RECT 286.000 237.600 286.800 238.400 ;
        RECT 289.300 232.400 289.900 279.600 ;
        RECT 290.900 272.400 291.500 287.600 ;
        RECT 290.800 271.600 291.600 272.400 ;
        RECT 292.500 268.300 293.100 289.600 ;
        RECT 294.100 278.400 294.700 293.600 ;
        RECT 294.000 277.600 294.800 278.400 ;
        RECT 295.700 274.400 296.300 323.600 ;
        RECT 297.200 309.600 298.000 310.400 ;
        RECT 295.600 273.600 296.400 274.400 ;
        RECT 297.300 270.400 297.900 309.600 ;
        RECT 298.600 307.600 299.600 308.400 ;
        RECT 302.100 304.300 302.700 323.600 ;
        RECT 314.900 322.400 315.500 331.600 ;
        RECT 321.300 326.400 321.900 333.600 ;
        RECT 326.000 331.600 326.800 332.400 ;
        RECT 327.700 328.400 328.300 333.600 ;
        RECT 329.300 332.400 329.900 333.600 ;
        RECT 329.200 331.600 330.000 332.400 ;
        RECT 332.400 331.600 333.200 332.400 ;
        RECT 329.200 329.600 330.000 330.400 ;
        RECT 327.600 327.600 328.400 328.400 ;
        RECT 321.200 325.600 322.000 326.400 ;
        RECT 314.800 321.600 315.600 322.400 ;
        RECT 306.800 309.600 307.600 310.400 ;
        RECT 306.900 306.400 307.500 309.600 ;
        RECT 306.800 305.600 307.600 306.400 ;
        RECT 300.500 303.700 302.700 304.300 ;
        RECT 308.400 304.200 309.200 317.800 ;
        RECT 310.000 304.200 310.800 317.800 ;
        RECT 311.600 304.200 312.400 317.800 ;
        RECT 313.200 304.200 314.000 315.800 ;
        RECT 314.800 305.600 315.600 306.400 ;
        RECT 314.900 304.400 315.500 305.600 ;
        RECT 298.800 297.600 299.600 298.400 ;
        RECT 298.800 273.600 299.600 274.400 ;
        RECT 295.600 269.600 296.400 270.400 ;
        RECT 297.200 269.600 298.000 270.400 ;
        RECT 290.900 267.700 293.100 268.300 ;
        RECT 290.900 258.400 291.500 267.700 ;
        RECT 292.400 265.600 293.200 266.400 ;
        RECT 290.800 257.600 291.600 258.400 ;
        RECT 290.900 254.400 291.500 257.600 ;
        RECT 290.800 253.600 291.600 254.400 ;
        RECT 292.500 252.300 293.100 265.600 ;
        RECT 295.700 264.400 296.300 269.600 ;
        RECT 295.600 263.600 296.400 264.400 ;
        RECT 298.900 254.400 299.500 273.600 ;
        RECT 300.500 268.400 301.100 303.700 ;
        RECT 314.800 303.600 315.600 304.400 ;
        RECT 316.400 304.200 317.200 315.800 ;
        RECT 318.000 307.600 318.800 308.400 ;
        RECT 318.100 304.400 318.700 307.600 ;
        RECT 318.000 303.600 318.800 304.400 ;
        RECT 319.600 304.200 320.400 315.800 ;
        RECT 321.200 304.200 322.000 317.800 ;
        RECT 322.800 304.200 323.600 317.800 ;
        RECT 334.100 314.400 334.700 333.600 ;
        RECT 334.000 313.600 334.800 314.400 ;
        RECT 332.400 307.600 333.200 308.400 ;
        RECT 324.400 305.600 325.200 306.400 ;
        RECT 316.400 297.600 317.200 298.400 ;
        RECT 316.500 294.400 317.100 297.600 ;
        RECT 316.400 293.600 317.200 294.400 ;
        RECT 305.200 291.600 306.000 292.400 ;
        RECT 322.800 291.600 323.600 292.400 ;
        RECT 305.200 289.600 306.000 290.400 ;
        RECT 314.800 289.600 315.600 290.400 ;
        RECT 319.600 289.600 320.400 290.400 ;
        RECT 322.800 289.600 323.600 290.400 ;
        RECT 313.200 285.600 314.000 286.400 ;
        RECT 302.000 273.600 302.800 274.400 ;
        RECT 302.100 270.400 302.700 273.600 ;
        RECT 302.000 269.600 302.800 270.400 ;
        RECT 300.400 267.600 301.200 268.400 ;
        RECT 308.400 267.600 309.200 268.400 ;
        RECT 300.400 265.600 301.200 266.400 ;
        RECT 300.500 258.400 301.100 265.600 ;
        RECT 300.400 257.600 301.200 258.400 ;
        RECT 313.300 256.400 313.900 285.600 ;
        RECT 319.700 284.400 320.300 289.600 ;
        RECT 314.800 283.600 315.600 284.400 ;
        RECT 319.600 283.600 320.400 284.400 ;
        RECT 314.900 268.300 315.500 283.600 ;
        RECT 324.500 278.300 325.100 305.600 ;
        RECT 335.700 298.400 336.300 341.600 ;
        RECT 337.200 329.600 338.000 330.400 ;
        RECT 337.200 327.600 338.000 328.400 ;
        RECT 337.300 324.400 337.900 327.600 ;
        RECT 340.400 325.600 341.200 326.400 ;
        RECT 337.200 323.600 338.000 324.400 ;
        RECT 337.300 312.400 337.900 323.600 ;
        RECT 340.500 322.400 341.100 325.600 ;
        RECT 340.400 321.600 341.200 322.400 ;
        RECT 337.200 311.600 338.000 312.400 ;
        RECT 332.400 297.600 333.200 298.400 ;
        RECT 335.600 297.600 336.400 298.400 ;
        RECT 327.600 293.600 328.400 294.400 ;
        RECT 329.200 293.600 330.000 294.400 ;
        RECT 329.300 292.400 329.900 293.600 ;
        RECT 329.200 291.600 330.000 292.400 ;
        RECT 330.800 291.600 331.600 292.400 ;
        RECT 326.000 289.600 326.800 290.400 ;
        RECT 326.100 280.400 326.700 289.600 ;
        RECT 329.300 286.400 329.900 291.600 ;
        RECT 332.500 290.400 333.100 297.600 ;
        RECT 334.000 293.600 334.800 294.400 ;
        RECT 334.100 290.400 334.700 293.600 ;
        RECT 332.400 289.600 333.200 290.400 ;
        RECT 334.000 289.600 334.800 290.400 ;
        RECT 334.100 286.400 334.700 289.600 ;
        RECT 329.200 285.600 330.000 286.400 ;
        RECT 334.000 285.600 334.800 286.400 ;
        RECT 335.600 281.600 336.400 282.400 ;
        RECT 326.000 279.600 326.800 280.400 ;
        RECT 334.000 279.600 334.800 280.400 ;
        RECT 314.900 267.700 317.100 268.300 ;
        RECT 308.400 255.600 309.200 256.400 ;
        RECT 313.200 255.600 314.000 256.400 ;
        RECT 308.500 254.400 309.100 255.600 ;
        RECT 297.200 253.600 298.000 254.400 ;
        RECT 298.800 253.600 299.600 254.400 ;
        RECT 303.600 253.600 304.400 254.400 ;
        RECT 308.400 253.600 309.200 254.400 ;
        RECT 314.800 253.600 315.600 254.400 ;
        RECT 297.300 252.400 297.900 253.600 ;
        RECT 290.900 251.700 293.100 252.300 ;
        RECT 289.200 231.600 290.000 232.400 ;
        RECT 282.800 229.700 285.100 230.300 ;
        RECT 282.800 229.600 283.600 229.700 ;
        RECT 287.600 229.600 288.400 230.400 ;
        RECT 249.200 221.600 250.000 222.400 ;
        RECT 249.300 218.400 249.900 221.600 ;
        RECT 220.400 204.200 221.200 217.800 ;
        RECT 222.000 204.200 222.800 217.800 ;
        RECT 223.600 206.200 224.400 217.800 ;
        RECT 225.200 213.600 226.000 214.400 ;
        RECT 226.800 206.200 227.600 217.800 ;
        RECT 228.400 217.600 229.200 218.400 ;
        RECT 228.500 216.400 229.100 217.600 ;
        RECT 228.400 215.600 229.200 216.400 ;
        RECT 217.200 193.600 218.000 194.400 ;
        RECT 207.600 191.600 208.400 192.400 ;
        RECT 207.700 190.400 208.300 191.600 ;
        RECT 204.400 189.600 205.200 190.400 ;
        RECT 207.600 189.600 208.400 190.400 ;
        RECT 214.000 189.600 214.800 190.400 ;
        RECT 218.800 189.600 219.600 190.400 ;
        RECT 210.800 187.600 211.600 188.400 ;
        RECT 212.400 187.600 213.200 188.400 ;
        RECT 212.500 186.400 213.100 187.600 ;
        RECT 206.000 185.600 206.800 186.400 ;
        RECT 212.400 185.600 213.200 186.400 ;
        RECT 204.400 183.600 205.200 184.400 ;
        RECT 204.500 172.400 205.100 183.600 ;
        RECT 206.100 174.400 206.700 185.600 ;
        RECT 214.100 184.400 214.700 189.600 ;
        RECT 215.600 187.600 216.400 188.400 ;
        RECT 214.000 183.600 214.800 184.400 ;
        RECT 218.900 180.400 219.500 189.600 ;
        RECT 223.600 187.600 224.400 188.400 ;
        RECT 225.200 183.600 226.000 184.400 ;
        RECT 225.300 182.400 225.900 183.600 ;
        RECT 225.200 181.600 226.000 182.400 ;
        RECT 207.600 179.600 208.400 180.400 ;
        RECT 218.800 179.600 219.600 180.400 ;
        RECT 206.000 173.600 206.800 174.400 ;
        RECT 201.200 171.600 202.000 172.400 ;
        RECT 204.400 171.600 205.200 172.400 ;
        RECT 196.400 169.600 197.200 170.400 ;
        RECT 199.600 169.600 200.400 170.400 ;
        RECT 201.200 169.600 202.000 170.400 ;
        RECT 193.200 157.600 194.000 158.400 ;
        RECT 204.500 150.400 205.100 171.600 ;
        RECT 207.700 150.400 208.300 179.600 ;
        RECT 228.500 178.400 229.100 215.600 ;
        RECT 230.000 206.200 230.800 217.800 ;
        RECT 231.600 204.200 232.400 217.800 ;
        RECT 233.200 204.200 234.000 217.800 ;
        RECT 234.800 204.200 235.600 217.800 ;
        RECT 244.400 217.600 245.200 218.400 ;
        RECT 247.600 217.600 248.400 218.400 ;
        RECT 249.200 217.600 250.000 218.400 ;
        RECT 246.000 215.600 246.800 216.400 ;
        RECT 236.400 203.600 237.200 204.400 ;
        RECT 244.400 203.600 245.200 204.400 ;
        RECT 236.500 194.400 237.100 203.600 ;
        RECT 236.400 193.600 237.200 194.400 ;
        RECT 244.400 193.600 245.200 194.400 ;
        RECT 233.200 189.600 234.000 190.400 ;
        RECT 234.800 189.600 235.600 190.400 ;
        RECT 239.600 189.600 240.400 190.400 ;
        RECT 231.600 187.600 232.400 188.400 ;
        RECT 233.300 184.400 233.900 189.600 ;
        RECT 238.000 187.600 238.800 188.400 ;
        RECT 239.700 184.400 240.300 189.600 ;
        RECT 233.200 183.600 234.000 184.400 ;
        RECT 239.600 183.600 240.400 184.400 ;
        RECT 212.400 175.600 213.200 176.400 ;
        RECT 209.200 169.600 210.000 170.400 ;
        RECT 201.200 149.600 202.000 150.400 ;
        RECT 204.400 149.600 205.200 150.400 ;
        RECT 207.600 149.600 208.400 150.400 ;
        RECT 209.200 149.600 210.000 150.400 ;
        RECT 198.000 147.600 198.800 148.400 ;
        RECT 196.400 143.600 197.200 144.400 ;
        RECT 193.200 139.600 194.000 140.400 ;
        RECT 190.000 135.600 190.800 136.400 ;
        RECT 193.300 132.400 193.900 139.600 ;
        RECT 196.500 134.400 197.100 143.600 ;
        RECT 198.100 138.400 198.700 147.600 ;
        RECT 204.400 145.600 205.200 146.400 ;
        RECT 198.000 137.600 198.800 138.400 ;
        RECT 207.600 135.600 208.400 136.400 ;
        RECT 196.400 133.600 197.200 134.400 ;
        RECT 201.200 133.600 202.000 134.400 ;
        RECT 202.800 133.600 203.600 134.400 ;
        RECT 202.900 132.400 203.500 133.600 ;
        RECT 207.700 132.400 208.300 135.600 ;
        RECT 209.300 132.400 209.900 149.600 ;
        RECT 212.500 146.400 213.100 175.600 ;
        RECT 218.800 164.200 219.600 177.800 ;
        RECT 220.400 164.200 221.200 177.800 ;
        RECT 222.000 164.200 222.800 177.800 ;
        RECT 223.600 166.200 224.400 177.800 ;
        RECT 225.200 177.600 226.000 178.400 ;
        RECT 225.300 176.400 225.900 177.600 ;
        RECT 225.200 175.600 226.000 176.400 ;
        RECT 225.300 168.400 225.900 175.600 ;
        RECT 225.200 167.600 226.000 168.400 ;
        RECT 226.800 166.200 227.600 177.800 ;
        RECT 228.400 177.600 229.200 178.400 ;
        RECT 228.400 173.600 229.200 174.400 ;
        RECT 228.500 172.400 229.100 173.600 ;
        RECT 228.400 171.600 229.200 172.400 ;
        RECT 230.000 166.200 230.800 177.800 ;
        RECT 231.600 164.200 232.400 177.800 ;
        RECT 233.200 164.200 234.000 177.800 ;
        RECT 246.100 174.400 246.700 215.600 ;
        RECT 255.700 212.400 256.300 229.600 ;
        RECT 263.600 227.600 264.600 228.400 ;
        RECT 274.800 227.600 275.600 228.400 ;
        RECT 282.900 226.400 283.500 229.600 ;
        RECT 284.400 227.600 285.200 228.400 ;
        RECT 290.900 228.300 291.500 251.700 ;
        RECT 297.200 251.600 298.000 252.400 ;
        RECT 292.400 249.600 293.200 250.400 ;
        RECT 302.000 249.600 302.800 250.400 ;
        RECT 292.500 244.400 293.100 249.600 ;
        RECT 300.400 245.600 301.200 246.400 ;
        RECT 292.400 243.600 293.200 244.400 ;
        RECT 300.500 232.400 301.100 245.600 ;
        RECT 302.100 236.400 302.700 249.600 ;
        RECT 302.000 235.600 302.800 236.400 ;
        RECT 303.700 232.400 304.300 253.600 ;
        RECT 314.800 249.600 315.600 250.400 ;
        RECT 310.000 243.600 310.800 244.400 ;
        RECT 313.200 243.600 314.000 244.400 ;
        RECT 297.200 232.300 298.000 232.400 ;
        RECT 295.700 231.700 298.000 232.300 ;
        RECT 295.700 230.400 296.300 231.700 ;
        RECT 297.200 231.600 298.000 231.700 ;
        RECT 300.400 231.600 301.200 232.400 ;
        RECT 302.000 231.600 302.800 232.400 ;
        RECT 303.600 231.600 304.400 232.400 ;
        RECT 305.200 231.600 306.000 232.400 ;
        RECT 295.600 229.600 296.400 230.400 ;
        RECT 297.200 229.600 298.000 230.400 ;
        RECT 302.100 228.400 302.700 231.600 ;
        RECT 305.300 228.400 305.900 231.600 ;
        RECT 289.300 227.700 291.500 228.300 ;
        RECT 282.800 225.600 283.600 226.400 ;
        RECT 279.600 223.600 280.400 224.400 ;
        RECT 255.600 211.600 256.400 212.400 ;
        RECT 258.800 204.200 259.600 217.800 ;
        RECT 260.400 204.200 261.200 217.800 ;
        RECT 262.000 206.200 262.800 217.800 ;
        RECT 263.600 213.600 264.400 214.400 ;
        RECT 265.200 206.200 266.000 217.800 ;
        RECT 266.800 215.600 267.600 216.400 ;
        RECT 268.400 206.200 269.200 217.800 ;
        RECT 270.000 204.200 270.800 217.800 ;
        RECT 271.600 204.200 272.400 217.800 ;
        RECT 273.200 204.200 274.000 217.800 ;
        RECT 274.800 215.600 275.600 216.400 ;
        RECT 274.900 212.400 275.500 215.600 ;
        RECT 279.700 214.400 280.300 223.600 ;
        RECT 284.500 216.400 285.100 227.600 ;
        RECT 287.600 226.300 288.400 226.400 ;
        RECT 286.100 225.700 288.400 226.300 ;
        RECT 284.400 215.600 285.200 216.400 ;
        RECT 279.600 213.600 280.400 214.400 ;
        RECT 274.800 211.600 275.600 212.400 ;
        RECT 282.800 205.600 283.600 206.400 ;
        RECT 247.600 191.600 248.400 192.400 ;
        RECT 249.200 189.600 250.000 190.400 ;
        RECT 254.000 189.600 254.800 190.400 ;
        RECT 258.800 189.600 259.600 190.400 ;
        RECT 249.300 188.400 249.900 189.600 ;
        RECT 247.600 187.600 248.400 188.400 ;
        RECT 249.200 187.600 250.000 188.400 ;
        RECT 246.000 173.600 246.800 174.400 ;
        RECT 249.300 172.400 249.900 187.600 ;
        RECT 254.100 182.400 254.700 189.600 ;
        RECT 263.600 184.200 264.400 197.800 ;
        RECT 265.200 184.200 266.000 197.800 ;
        RECT 266.800 184.200 267.600 195.800 ;
        RECT 268.400 187.600 269.200 188.400 ;
        RECT 270.000 184.200 270.800 195.800 ;
        RECT 271.600 195.600 272.400 196.400 ;
        RECT 271.700 186.400 272.300 195.600 ;
        RECT 271.600 185.600 272.400 186.400 ;
        RECT 273.200 184.200 274.000 195.800 ;
        RECT 274.800 184.200 275.600 197.800 ;
        RECT 276.400 184.200 277.200 197.800 ;
        RECT 278.000 184.200 278.800 197.800 ;
        RECT 286.100 194.400 286.700 225.700 ;
        RECT 287.600 225.600 288.400 225.700 ;
        RECT 287.600 215.600 288.400 216.400 ;
        RECT 287.700 206.400 288.300 215.600 ;
        RECT 287.600 205.600 288.400 206.400 ;
        RECT 286.000 193.600 286.800 194.400 ;
        RECT 287.600 193.600 288.400 194.400 ;
        RECT 289.300 192.400 289.900 227.700 ;
        RECT 294.000 227.600 294.800 228.400 ;
        RECT 295.600 227.600 296.400 228.400 ;
        RECT 302.000 227.600 302.800 228.400 ;
        RECT 303.600 227.600 304.400 228.400 ;
        RECT 305.200 227.600 306.000 228.400 ;
        RECT 295.700 222.400 296.300 227.600 ;
        RECT 295.600 221.600 296.400 222.400 ;
        RECT 310.100 218.400 310.700 243.600 ;
        RECT 313.300 234.300 313.900 243.600 ;
        RECT 311.700 233.700 313.900 234.300 ;
        RECT 311.700 230.400 312.300 233.700 ;
        RECT 313.200 231.600 314.000 232.400 ;
        RECT 314.900 232.300 315.500 249.600 ;
        RECT 316.500 248.400 317.100 267.700 ;
        RECT 318.000 264.200 318.800 277.800 ;
        RECT 319.600 264.200 320.400 277.800 ;
        RECT 322.900 277.700 325.100 278.300 ;
        RECT 321.200 264.200 322.000 275.800 ;
        RECT 322.900 270.400 323.500 277.700 ;
        RECT 322.800 269.600 323.600 270.400 ;
        RECT 322.800 267.600 323.600 268.400 ;
        RECT 324.400 264.200 325.200 275.800 ;
        RECT 326.000 265.600 326.800 266.400 ;
        RECT 327.600 264.200 328.400 275.800 ;
        RECT 329.200 264.200 330.000 277.800 ;
        RECT 330.800 264.200 331.600 277.800 ;
        RECT 332.400 264.200 333.200 277.800 ;
        RECT 318.000 257.600 318.800 258.400 ;
        RECT 318.100 250.400 318.700 257.600 ;
        RECT 327.600 255.600 328.400 256.400 ;
        RECT 327.700 254.400 328.300 255.600 ;
        RECT 334.100 254.400 334.700 279.600 ;
        RECT 327.600 253.600 328.400 254.400 ;
        RECT 334.000 253.600 334.800 254.400 ;
        RECT 319.600 251.600 320.400 252.400 ;
        RECT 324.400 251.600 325.200 252.400 ;
        RECT 329.200 251.600 330.000 252.400 ;
        RECT 324.500 250.400 325.100 251.600 ;
        RECT 318.000 249.600 318.800 250.400 ;
        RECT 321.200 249.600 322.000 250.400 ;
        RECT 324.400 249.600 325.200 250.400 ;
        RECT 316.400 247.600 317.200 248.400 ;
        RECT 319.600 247.600 320.400 248.400 ;
        RECT 316.400 245.600 317.200 246.400 ;
        RECT 316.500 244.400 317.100 245.600 ;
        RECT 316.400 243.600 317.200 244.400 ;
        RECT 316.500 234.300 317.100 243.600 ;
        RECT 319.700 238.400 320.300 247.600 ;
        RECT 321.300 244.400 321.900 249.600 ;
        RECT 329.300 248.400 329.900 251.600 ;
        RECT 324.400 247.600 325.200 248.400 ;
        RECT 329.200 247.600 330.000 248.400 ;
        RECT 321.200 243.600 322.000 244.400 ;
        RECT 326.000 243.600 326.800 244.400 ;
        RECT 329.200 243.600 330.000 244.400 ;
        RECT 326.100 238.400 326.700 243.600 ;
        RECT 319.600 237.600 320.400 238.400 ;
        RECT 326.000 237.600 326.800 238.400 ;
        RECT 316.500 233.700 318.700 234.300 ;
        RECT 318.100 232.400 318.700 233.700 ;
        RECT 321.200 233.600 322.000 234.400 ;
        RECT 316.400 232.300 317.200 232.400 ;
        RECT 314.900 231.700 317.200 232.300 ;
        RECT 316.400 231.600 317.200 231.700 ;
        RECT 318.000 231.600 318.800 232.400 ;
        RECT 311.600 229.600 312.400 230.400 ;
        RECT 319.600 229.600 320.400 230.400 ;
        RECT 311.600 227.600 312.400 228.400 ;
        RECT 311.700 222.400 312.300 227.600 ;
        RECT 326.000 223.600 326.800 224.400 ;
        RECT 311.600 221.600 312.400 222.400 ;
        RECT 300.400 217.600 301.200 218.400 ;
        RECT 310.000 217.600 310.800 218.400 ;
        RECT 297.200 213.600 298.000 214.400 ;
        RECT 290.800 203.600 291.600 204.400 ;
        RECT 290.900 196.400 291.500 203.600 ;
        RECT 290.800 195.600 291.600 196.400 ;
        RECT 289.200 191.600 290.000 192.400 ;
        RECT 254.000 181.600 254.800 182.400 ;
        RECT 289.300 178.400 289.900 191.600 ;
        RECT 294.000 189.600 294.800 190.400 ;
        RECT 295.600 189.600 296.400 190.400 ;
        RECT 292.400 185.600 293.200 186.400 ;
        RECT 290.800 183.600 291.600 184.400 ;
        RECT 238.000 171.600 238.800 172.400 ;
        RECT 249.200 171.600 250.000 172.400 ;
        RECT 223.600 155.600 224.400 156.400 ;
        RECT 223.700 154.400 224.300 155.600 ;
        RECT 223.600 153.600 224.400 154.400 ;
        RECT 214.000 151.600 214.800 152.400 ;
        RECT 214.000 149.600 214.800 150.400 ;
        RECT 220.400 149.600 221.200 150.400 ;
        RECT 217.200 147.600 218.000 148.400 ;
        RECT 218.800 147.600 219.600 148.400 ;
        RECT 222.000 147.600 222.800 148.400 ;
        RECT 218.900 146.400 219.500 147.600 ;
        RECT 212.400 145.600 213.200 146.400 ;
        RECT 218.800 145.600 219.600 146.400 ;
        RECT 210.800 143.600 211.600 144.400 ;
        RECT 215.600 143.600 216.400 144.400 ;
        RECT 233.200 144.200 234.000 157.800 ;
        RECT 234.800 144.200 235.600 157.800 ;
        RECT 236.400 144.200 237.200 155.800 ;
        RECT 238.100 150.400 238.700 171.600 ;
        RECT 241.200 159.600 242.000 160.400 ;
        RECT 238.000 149.600 238.800 150.400 ;
        RECT 238.000 147.600 238.800 148.400 ;
        RECT 238.100 144.400 238.700 147.600 ;
        RECT 238.000 143.600 238.800 144.400 ;
        RECT 239.600 144.200 240.400 155.800 ;
        RECT 241.300 146.400 241.900 159.600 ;
        RECT 241.200 145.600 242.000 146.400 ;
        RECT 242.800 144.200 243.600 155.800 ;
        RECT 244.400 144.200 245.200 157.800 ;
        RECT 246.000 144.200 246.800 157.800 ;
        RECT 247.600 144.200 248.400 157.800 ;
        RECT 249.300 150.400 249.900 171.600 ;
        RECT 250.800 164.200 251.600 177.800 ;
        RECT 252.400 164.200 253.200 177.800 ;
        RECT 254.000 166.200 254.800 177.800 ;
        RECT 255.600 173.600 256.400 174.400 ;
        RECT 257.200 166.200 258.000 177.800 ;
        RECT 258.800 175.600 259.600 176.400 ;
        RECT 258.900 160.400 259.500 175.600 ;
        RECT 260.400 166.200 261.200 177.800 ;
        RECT 262.000 164.200 262.800 177.800 ;
        RECT 263.600 164.200 264.400 177.800 ;
        RECT 265.200 164.200 266.000 177.800 ;
        RECT 274.800 177.600 275.600 178.400 ;
        RECT 289.200 177.600 290.000 178.400 ;
        RECT 290.900 174.400 291.500 183.600 ;
        RECT 276.400 173.600 277.200 174.400 ;
        RECT 281.200 173.600 282.000 174.400 ;
        RECT 290.800 173.600 291.600 174.400 ;
        RECT 278.000 169.600 278.800 170.400 ;
        RECT 258.800 159.600 259.600 160.400 ;
        RECT 257.200 155.600 258.000 156.400 ;
        RECT 271.600 153.600 272.400 154.400 ;
        RECT 260.400 151.600 261.200 152.400 ;
        RECT 249.200 149.600 250.000 150.400 ;
        RECT 252.400 149.600 253.200 150.400 ;
        RECT 266.800 149.600 267.600 150.400 ;
        RECT 249.200 145.600 250.000 146.400 ;
        RECT 193.200 131.600 194.000 132.400 ;
        RECT 202.800 131.600 203.600 132.400 ;
        RECT 207.600 131.600 208.400 132.400 ;
        RECT 209.200 131.600 210.000 132.400 ;
        RECT 198.000 129.600 198.800 130.400 ;
        RECT 209.200 129.600 210.000 130.400 ;
        RECT 193.200 117.600 194.000 118.400 ;
        RECT 182.100 113.700 184.300 114.300 ;
        RECT 164.400 111.600 165.200 112.400 ;
        RECT 153.200 109.600 154.000 110.400 ;
        RECT 158.000 109.600 158.800 110.400 ;
        RECT 174.000 109.600 174.800 110.400 ;
        RECT 175.600 109.600 176.400 110.400 ;
        RECT 180.400 109.600 181.200 110.400 ;
        RECT 158.000 107.600 158.800 108.400 ;
        RECT 159.600 107.600 160.400 108.400 ;
        RECT 156.400 105.600 157.200 106.400 ;
        RECT 150.000 91.600 150.800 92.400 ;
        RECT 146.800 87.600 147.600 88.400 ;
        RECT 148.400 87.600 149.200 88.400 ;
        RECT 150.000 75.600 150.800 76.400 ;
        RECT 145.200 73.600 146.000 74.400 ;
        RECT 148.400 73.600 149.200 74.400 ;
        RECT 145.200 72.300 146.000 72.400 ;
        RECT 143.700 71.700 146.000 72.300 ;
        RECT 145.200 71.600 146.000 71.700 ;
        RECT 146.800 69.600 147.600 70.400 ;
        RECT 146.900 68.400 147.500 69.600 ;
        RECT 140.400 67.600 141.200 68.400 ;
        RECT 146.800 67.600 147.600 68.400 ;
        RECT 140.400 55.600 141.200 56.400 ;
        RECT 143.600 56.300 144.400 56.400 ;
        RECT 146.800 56.300 147.600 56.400 ;
        RECT 143.600 55.700 147.600 56.300 ;
        RECT 143.600 55.600 144.400 55.700 ;
        RECT 146.800 55.600 147.600 55.700 ;
        RECT 140.500 52.400 141.100 55.600 ;
        RECT 138.800 51.600 139.600 52.400 ;
        RECT 140.400 51.600 141.200 52.400 ;
        RECT 145.200 51.600 146.000 52.400 ;
        RECT 146.800 51.600 147.600 52.400 ;
        RECT 137.200 49.600 138.000 50.400 ;
        RECT 134.000 45.600 134.800 46.400 ;
        RECT 134.100 44.400 134.700 45.600 ;
        RECT 134.000 43.600 134.800 44.400 ;
        RECT 130.800 35.600 131.600 36.400 ;
        RECT 134.100 34.400 134.700 43.600 ;
        RECT 134.000 33.600 134.800 34.400 ;
        RECT 129.200 31.600 130.000 32.400 ;
        RECT 134.000 31.600 134.800 32.400 ;
        RECT 114.800 27.600 115.600 28.400 ;
        RECT 126.000 27.600 126.800 28.400 ;
        RECT 127.600 27.600 128.400 28.400 ;
        RECT 126.100 20.400 126.700 27.600 ;
        RECT 129.200 25.600 130.000 26.400 ;
        RECT 100.400 19.600 101.200 20.400 ;
        RECT 126.000 19.600 126.800 20.400 ;
        RECT 90.800 17.600 91.600 18.400 ;
        RECT 89.200 13.600 90.000 14.400 ;
        RECT 87.600 11.600 88.400 12.400 ;
        RECT 84.400 9.600 85.200 10.400 ;
        RECT 95.600 6.200 96.400 17.800 ;
        RECT 100.500 14.400 101.100 19.600 ;
        RECT 100.400 13.600 101.200 14.400 ;
        RECT 102.000 13.600 102.800 14.400 ;
        RECT 100.500 12.400 101.100 13.600 ;
        RECT 102.100 12.400 102.700 13.600 ;
        RECT 100.400 11.600 101.200 12.400 ;
        RECT 102.000 11.600 102.800 12.400 ;
        RECT 105.200 6.200 106.000 17.800 ;
        RECT 110.000 17.600 110.800 18.400 ;
        RECT 108.400 10.200 109.200 15.800 ;
        RECT 114.800 6.200 115.600 17.800 ;
        RECT 116.400 11.600 117.200 12.400 ;
        RECT 122.800 11.600 123.600 12.600 ;
        RECT 124.400 6.200 125.200 17.800 ;
        RECT 127.600 10.200 128.400 15.800 ;
        RECT 129.300 14.400 129.900 25.600 ;
        RECT 132.400 23.600 133.200 24.400 ;
        RECT 130.800 19.600 131.600 20.400 ;
        RECT 130.900 18.400 131.500 19.600 ;
        RECT 130.800 17.600 131.600 18.400 ;
        RECT 129.200 13.600 130.000 14.400 ;
        RECT 132.500 12.400 133.100 23.600 ;
        RECT 134.100 18.400 134.700 31.600 ;
        RECT 137.300 30.400 137.900 49.600 ;
        RECT 145.300 48.400 145.900 51.600 ;
        RECT 148.500 48.400 149.100 73.600 ;
        RECT 150.100 70.400 150.700 75.600 ;
        RECT 156.500 74.400 157.100 105.600 ;
        RECT 158.100 104.400 158.700 107.600 ;
        RECT 158.000 103.600 158.800 104.400 ;
        RECT 158.000 83.600 158.800 84.400 ;
        RECT 158.100 78.400 158.700 83.600 ;
        RECT 158.000 77.600 158.800 78.400 ;
        RECT 156.400 73.600 157.200 74.400 ;
        RECT 150.000 69.600 150.800 70.400 ;
        RECT 156.500 68.400 157.100 73.600 ;
        RECT 156.400 67.600 157.200 68.400 ;
        RECT 158.000 66.200 158.800 71.800 ;
        RECT 154.800 55.600 155.600 56.400 ;
        RECT 153.200 53.600 154.000 54.400 ;
        RECT 145.200 47.600 146.000 48.400 ;
        RECT 148.400 47.600 149.200 48.400 ;
        RECT 145.300 38.400 145.900 47.600 ;
        RECT 153.300 46.400 153.900 53.600 ;
        RECT 154.900 52.400 155.500 55.600 ;
        RECT 159.700 54.400 160.300 107.600 ;
        RECT 174.100 104.400 174.700 109.600 ;
        RECT 180.500 108.400 181.100 109.600 ;
        RECT 180.400 107.600 181.200 108.400 ;
        RECT 174.000 103.600 174.800 104.400 ;
        RECT 178.800 103.600 179.600 104.400 ;
        RECT 162.800 86.200 163.600 97.800 ;
        RECT 169.200 93.600 170.000 94.400 ;
        RECT 161.200 64.200 162.000 75.800 ;
        RECT 162.800 69.400 163.600 70.400 ;
        RECT 164.400 67.600 165.200 68.400 ;
        RECT 162.800 65.600 163.600 66.400 ;
        RECT 162.900 62.300 163.500 65.600 ;
        RECT 161.300 61.700 163.500 62.300 ;
        RECT 159.600 53.600 160.400 54.400 ;
        RECT 154.800 51.600 155.600 52.400 ;
        RECT 156.400 51.600 157.200 52.400 ;
        RECT 153.200 45.600 154.000 46.400 ;
        RECT 140.400 37.600 141.200 38.400 ;
        RECT 145.200 37.600 146.000 38.400 ;
        RECT 137.200 29.600 138.000 30.400 ;
        RECT 138.800 27.600 139.600 28.400 ;
        RECT 138.900 20.400 139.500 27.600 ;
        RECT 145.200 24.200 146.000 35.800 ;
        RECT 146.800 29.600 147.600 30.400 ;
        RECT 146.900 26.400 147.500 29.600 ;
        RECT 153.200 29.400 154.000 30.400 ;
        RECT 146.800 25.600 147.600 26.400 ;
        RECT 146.800 23.600 147.600 24.400 ;
        RECT 154.800 24.200 155.600 35.800 ;
        RECT 156.500 30.400 157.100 51.600 ;
        RECT 159.600 49.600 160.400 50.400 ;
        RECT 159.700 48.400 160.300 49.600 ;
        RECT 159.600 47.600 160.400 48.400 ;
        RECT 156.400 29.600 157.200 30.400 ;
        RECT 158.000 26.200 158.800 31.800 ;
        RECT 161.300 28.400 161.900 61.700 ;
        RECT 162.800 59.600 163.600 60.400 ;
        RECT 162.900 52.400 163.500 59.600 ;
        RECT 164.500 54.400 165.100 67.600 ;
        RECT 169.300 54.400 169.900 93.600 ;
        RECT 170.800 91.800 171.600 92.600 ;
        RECT 170.900 82.400 171.500 91.800 ;
        RECT 172.400 86.200 173.200 97.800 ;
        RECT 175.600 90.200 176.400 95.800 ;
        RECT 178.900 94.400 179.500 103.600 ;
        RECT 178.800 93.600 179.600 94.400 ;
        RECT 182.100 92.400 182.700 113.700 ;
        RECT 183.600 109.600 184.400 110.400 ;
        RECT 185.200 109.600 186.000 110.400 ;
        RECT 183.700 106.400 184.300 109.600 ;
        RECT 186.800 107.600 187.600 108.400 ;
        RECT 191.600 107.600 192.400 108.400 ;
        RECT 186.900 106.400 187.500 107.600 ;
        RECT 183.600 105.600 184.400 106.400 ;
        RECT 186.800 105.600 187.600 106.400 ;
        RECT 182.000 91.600 182.800 92.400 ;
        RECT 175.600 85.600 176.400 86.400 ;
        RECT 170.800 81.600 171.600 82.400 ;
        RECT 175.700 78.400 176.300 85.600 ;
        RECT 185.200 84.200 186.000 97.800 ;
        RECT 186.800 84.200 187.600 97.800 ;
        RECT 188.400 86.200 189.200 97.800 ;
        RECT 190.000 93.600 190.800 94.400 ;
        RECT 191.600 86.200 192.400 97.800 ;
        RECT 193.300 96.400 193.900 117.600 ;
        RECT 198.100 116.400 198.700 129.600 ;
        RECT 198.000 115.600 198.800 116.400 ;
        RECT 195.000 111.800 195.800 112.600 ;
        RECT 201.200 111.800 202.000 112.600 ;
        RECT 195.000 107.000 195.600 111.800 ;
        RECT 196.200 109.800 197.000 110.600 ;
        RECT 196.400 108.400 197.000 109.800 ;
        RECT 198.000 109.600 198.800 110.400 ;
        RECT 201.400 108.400 202.000 111.800 ;
        RECT 202.800 109.600 203.600 110.400 ;
        RECT 202.900 108.400 203.500 109.600 ;
        RECT 210.900 108.400 211.500 143.600 ;
        RECT 218.800 133.600 219.600 134.400 ;
        RECT 218.900 132.400 219.500 133.600 ;
        RECT 218.800 131.600 219.600 132.400 ;
        RECT 220.400 124.200 221.200 137.800 ;
        RECT 222.000 124.200 222.800 137.800 ;
        RECT 223.600 124.200 224.400 137.800 ;
        RECT 225.200 126.200 226.000 137.800 ;
        RECT 226.800 135.600 227.600 136.400 ;
        RECT 223.600 119.600 224.400 120.400 ;
        RECT 218.800 115.600 219.600 116.400 ;
        RECT 218.900 112.400 219.500 115.600 ;
        RECT 223.700 114.400 224.300 119.600 ;
        RECT 226.900 118.400 227.500 135.600 ;
        RECT 228.400 126.200 229.200 137.800 ;
        RECT 230.000 133.600 230.800 134.400 ;
        RECT 231.600 126.200 232.400 137.800 ;
        RECT 233.200 124.200 234.000 137.800 ;
        RECT 234.800 124.200 235.600 137.800 ;
        RECT 249.300 136.400 249.900 145.600 ;
        RECT 247.600 135.600 248.400 136.400 ;
        RECT 249.200 135.600 250.000 136.400 ;
        RECT 244.400 133.600 245.200 134.400 ;
        RECT 244.400 131.600 245.200 132.400 ;
        RECT 238.000 127.600 238.800 128.400 ;
        RECT 228.400 121.600 229.200 122.400 ;
        RECT 226.800 117.600 227.600 118.400 ;
        RECT 226.900 114.400 227.500 117.600 ;
        RECT 220.400 113.600 221.200 114.400 ;
        RECT 223.600 113.600 224.400 114.400 ;
        RECT 226.800 113.600 227.600 114.400 ;
        RECT 214.000 111.600 214.800 112.400 ;
        RECT 217.200 111.600 218.000 112.400 ;
        RECT 218.800 111.600 219.600 112.400 ;
        RECT 214.100 108.400 214.700 111.600 ;
        RECT 215.600 109.600 216.400 110.400 ;
        RECT 196.400 107.800 202.000 108.400 ;
        RECT 196.400 107.000 197.200 107.200 ;
        RECT 199.800 107.000 200.600 107.200 ;
        RECT 201.400 107.000 202.000 107.800 ;
        RECT 202.800 107.600 203.600 108.400 ;
        RECT 207.600 107.600 208.400 108.400 ;
        RECT 209.200 107.600 210.000 108.400 ;
        RECT 210.800 107.600 211.600 108.400 ;
        RECT 214.000 107.600 214.800 108.400 ;
        RECT 195.000 106.400 200.600 107.000 ;
        RECT 195.000 106.200 195.800 106.400 ;
        RECT 201.200 106.200 202.000 107.000 ;
        RECT 204.400 103.600 205.200 104.400 ;
        RECT 193.200 95.600 194.000 96.400 ;
        RECT 194.800 86.200 195.600 97.800 ;
        RECT 196.400 84.200 197.200 97.800 ;
        RECT 198.000 84.200 198.800 97.800 ;
        RECT 199.600 84.200 200.400 97.800 ;
        RECT 201.200 91.600 202.000 92.400 ;
        RECT 186.800 81.600 187.600 82.400 ;
        RECT 186.900 78.400 187.500 81.600 ;
        RECT 190.000 79.600 190.800 80.400 ;
        RECT 175.600 77.600 176.400 78.400 ;
        RECT 182.000 77.600 182.800 78.400 ;
        RECT 186.800 77.600 187.600 78.400 ;
        RECT 170.800 64.200 171.600 75.800 ;
        RECT 182.100 72.400 182.700 77.600 ;
        RECT 188.400 73.600 189.200 74.400 ;
        RECT 182.000 71.600 182.800 72.400 ;
        RECT 182.100 70.400 182.700 71.600 ;
        RECT 178.800 69.600 179.600 70.400 ;
        RECT 182.000 69.600 182.800 70.400 ;
        RECT 186.800 69.600 187.600 70.400 ;
        RECT 177.200 67.600 178.000 68.400 ;
        RECT 174.000 61.600 174.800 62.400 ;
        RECT 164.400 53.600 165.200 54.400 ;
        RECT 166.000 53.600 166.800 54.400 ;
        RECT 169.200 53.600 170.000 54.400 ;
        RECT 162.800 51.600 163.600 52.400 ;
        RECT 162.900 50.400 163.500 51.600 ;
        RECT 162.800 49.600 163.600 50.400 ;
        RECT 161.200 27.600 162.000 28.400 ;
        RECT 162.800 25.600 163.600 26.400 ;
        RECT 162.900 24.400 163.500 25.600 ;
        RECT 162.800 23.600 163.600 24.400 ;
        RECT 138.800 19.600 139.600 20.400 ;
        RECT 146.900 18.400 147.500 23.600 ;
        RECT 154.800 21.600 155.600 22.400 ;
        RECT 134.000 17.600 134.800 18.400 ;
        RECT 146.800 17.600 147.600 18.400 ;
        RECT 134.000 15.600 134.800 16.400 ;
        RECT 134.100 12.400 134.700 15.600 ;
        RECT 154.900 12.400 155.500 21.600 ;
        RECT 164.500 20.400 165.100 53.600 ;
        RECT 174.100 32.400 174.700 61.600 ;
        RECT 178.900 60.400 179.500 69.600 ;
        RECT 186.900 68.400 187.500 69.600 ;
        RECT 188.500 68.400 189.100 73.600 ;
        RECT 190.100 70.400 190.700 79.600 ;
        RECT 199.600 73.600 200.400 74.400 ;
        RECT 199.700 72.400 200.300 73.600 ;
        RECT 196.400 71.600 197.200 72.400 ;
        RECT 199.600 71.600 200.400 72.400 ;
        RECT 196.500 70.400 197.100 71.600 ;
        RECT 201.300 70.400 201.900 91.600 ;
        RECT 204.500 90.400 205.100 103.600 ;
        RECT 204.400 89.600 205.200 90.400 ;
        RECT 207.700 80.400 208.300 107.600 ;
        RECT 209.300 98.400 209.900 107.600 ;
        RECT 210.800 105.600 211.600 106.400 ;
        RECT 215.700 104.400 216.300 109.600 ;
        RECT 217.300 108.400 217.900 111.600 ;
        RECT 218.800 109.600 219.600 110.400 ;
        RECT 222.000 109.600 222.800 110.400 ;
        RECT 225.200 109.600 226.000 110.400 ;
        RECT 217.200 107.600 218.000 108.400 ;
        RECT 218.800 107.600 219.600 108.400 ;
        RECT 212.400 103.600 213.200 104.400 ;
        RECT 215.600 103.600 216.400 104.400 ;
        RECT 209.200 97.600 210.000 98.400 ;
        RECT 212.500 92.400 213.100 103.600 ;
        RECT 218.900 94.400 219.500 107.600 ;
        RECT 222.100 94.400 222.700 109.600 ;
        RECT 225.300 108.400 225.900 109.600 ;
        RECT 225.200 107.600 226.000 108.400 ;
        RECT 226.800 107.600 227.600 108.400 ;
        RECT 226.900 106.400 227.500 107.600 ;
        RECT 225.200 105.600 226.000 106.400 ;
        RECT 226.800 105.600 227.600 106.400 ;
        RECT 223.600 103.600 224.400 104.400 ;
        RECT 223.700 98.400 224.300 103.600 ;
        RECT 223.600 97.600 224.400 98.400 ;
        RECT 225.300 96.300 225.900 105.600 ;
        RECT 226.900 98.400 227.500 105.600 ;
        RECT 226.800 97.600 227.600 98.400 ;
        RECT 226.800 96.300 227.600 96.400 ;
        RECT 225.300 95.700 227.600 96.300 ;
        RECT 226.800 95.600 227.600 95.700 ;
        RECT 226.900 94.400 227.500 95.600 ;
        RECT 217.200 93.600 218.000 94.400 ;
        RECT 218.800 93.600 219.600 94.400 ;
        RECT 222.000 93.600 222.800 94.400 ;
        RECT 226.800 93.600 227.600 94.400 ;
        RECT 217.300 92.400 217.900 93.600 ;
        RECT 212.400 91.600 213.200 92.400 ;
        RECT 215.600 91.600 216.400 92.400 ;
        RECT 217.200 91.600 218.000 92.400 ;
        RECT 222.100 90.400 222.700 93.600 ;
        RECT 226.800 91.600 227.600 92.400 ;
        RECT 212.400 89.600 213.200 90.400 ;
        RECT 215.600 89.600 216.400 90.400 ;
        RECT 222.000 89.600 222.800 90.400 ;
        RECT 207.600 79.600 208.400 80.400 ;
        RECT 202.800 71.600 203.600 72.400 ;
        RECT 190.000 69.600 190.800 70.400 ;
        RECT 191.600 69.600 192.400 70.400 ;
        RECT 196.400 69.600 197.200 70.400 ;
        RECT 201.200 69.600 202.000 70.400 ;
        RECT 202.900 68.400 203.500 71.600 ;
        RECT 207.600 69.600 208.400 70.400 ;
        RECT 186.800 67.600 187.600 68.400 ;
        RECT 188.400 67.600 189.200 68.400 ;
        RECT 193.200 67.600 194.000 68.400 ;
        RECT 201.200 67.600 202.000 68.400 ;
        RECT 202.800 67.600 203.600 68.400 ;
        RECT 193.300 66.400 193.900 67.600 ;
        RECT 193.200 65.600 194.000 66.400 ;
        RECT 196.400 65.600 197.200 66.400 ;
        RECT 178.800 59.600 179.600 60.400 ;
        RECT 178.800 53.600 179.600 54.400 ;
        RECT 185.200 51.600 186.000 52.400 ;
        RECT 167.600 31.600 168.400 32.400 ;
        RECT 174.000 31.600 174.800 32.400 ;
        RECT 180.200 31.600 181.000 32.400 ;
        RECT 167.700 28.400 168.300 31.600 ;
        RECT 180.300 30.400 180.900 31.600 ;
        RECT 180.200 29.600 181.000 30.400 ;
        RECT 167.600 27.600 168.400 28.400 ;
        RECT 172.400 23.600 173.200 24.400 ;
        RECT 164.400 19.600 165.200 20.400 ;
        RECT 132.400 11.600 133.200 12.400 ;
        RECT 134.000 11.600 134.800 12.400 ;
        RECT 154.800 11.600 155.600 12.400 ;
        RECT 156.400 4.200 157.200 17.800 ;
        RECT 158.000 4.200 158.800 17.800 ;
        RECT 159.600 4.200 160.400 17.800 ;
        RECT 161.200 6.200 162.000 17.800 ;
        RECT 162.800 15.600 163.600 16.400 ;
        RECT 164.400 6.200 165.200 17.800 ;
        RECT 166.000 13.600 166.800 14.400 ;
        RECT 167.600 6.200 168.400 17.800 ;
        RECT 169.200 4.200 170.000 17.800 ;
        RECT 170.800 4.200 171.600 17.800 ;
        RECT 172.500 14.400 173.100 23.600 ;
        RECT 185.300 20.400 185.900 51.600 ;
        RECT 188.400 44.200 189.200 57.800 ;
        RECT 190.000 44.200 190.800 57.800 ;
        RECT 191.600 46.200 192.400 57.800 ;
        RECT 193.200 55.600 194.000 56.400 ;
        RECT 193.300 54.400 193.900 55.600 ;
        RECT 193.200 53.600 194.000 54.400 ;
        RECT 194.800 46.200 195.600 57.800 ;
        RECT 196.500 56.400 197.100 65.600 ;
        RECT 212.400 64.200 213.200 77.800 ;
        RECT 214.000 64.200 214.800 77.800 ;
        RECT 215.600 64.200 216.400 75.800 ;
        RECT 217.200 67.600 218.000 68.400 ;
        RECT 218.800 64.200 219.600 75.800 ;
        RECT 220.400 65.600 221.200 66.400 ;
        RECT 222.000 64.200 222.800 75.800 ;
        RECT 223.600 64.200 224.400 77.800 ;
        RECT 225.200 64.200 226.000 77.800 ;
        RECT 226.800 64.200 227.600 77.800 ;
        RECT 196.400 55.600 197.200 56.400 ;
        RECT 196.500 54.400 197.100 55.600 ;
        RECT 196.400 53.600 197.200 54.400 ;
        RECT 188.400 29.600 189.200 30.400 ;
        RECT 188.500 20.400 189.100 29.600 ;
        RECT 190.000 24.200 190.800 37.800 ;
        RECT 191.600 24.200 192.400 37.800 ;
        RECT 193.200 24.200 194.000 37.800 ;
        RECT 194.800 24.200 195.600 35.800 ;
        RECT 196.500 26.400 197.100 53.600 ;
        RECT 198.000 46.200 198.800 57.800 ;
        RECT 199.600 44.200 200.400 57.800 ;
        RECT 201.200 44.200 202.000 57.800 ;
        RECT 202.800 44.200 203.600 57.800 ;
        RECT 212.400 57.600 213.200 58.400 ;
        RECT 222.000 57.600 222.800 58.400 ;
        RECT 222.100 56.400 222.700 57.600 ;
        RECT 220.400 55.600 221.200 56.400 ;
        RECT 222.000 55.600 222.800 56.400 ;
        RECT 228.500 56.300 229.100 121.600 ;
        RECT 238.100 116.400 238.700 127.600 ;
        RECT 238.000 115.600 238.800 116.400 ;
        RECT 238.100 112.400 238.700 115.600 ;
        RECT 238.000 111.600 238.800 112.400 ;
        RECT 244.500 110.400 245.100 131.600 ;
        RECT 247.700 120.400 248.300 135.600 ;
        RECT 249.300 134.400 249.900 135.600 ;
        RECT 249.200 133.600 250.000 134.400 ;
        RECT 252.500 132.400 253.100 149.600 ;
        RECT 263.600 147.600 264.400 148.400 ;
        RECT 262.000 143.600 262.800 144.400 ;
        RECT 254.000 135.600 254.800 136.400 ;
        RECT 254.100 132.400 254.700 135.600 ;
        RECT 262.100 134.400 262.700 143.600 ;
        RECT 263.700 134.400 264.300 147.600 ;
        RECT 260.400 133.600 261.200 134.400 ;
        RECT 262.000 133.600 262.800 134.400 ;
        RECT 263.600 133.600 264.400 134.400 ;
        RECT 252.400 131.600 253.200 132.400 ;
        RECT 254.000 131.600 254.800 132.400 ;
        RECT 262.000 131.600 262.800 132.400 ;
        RECT 257.200 129.600 258.000 130.400 ;
        RECT 257.300 124.400 257.900 129.600 ;
        RECT 250.800 123.600 251.600 124.400 ;
        RECT 257.200 123.600 258.000 124.400 ;
        RECT 247.600 119.600 248.400 120.400 ;
        RECT 249.200 117.600 250.000 118.400 ;
        RECT 233.200 109.600 234.000 110.400 ;
        RECT 236.400 109.600 237.200 110.400 ;
        RECT 241.200 109.600 242.000 110.400 ;
        RECT 244.400 109.600 245.200 110.400 ;
        RECT 241.300 106.400 241.900 109.600 ;
        RECT 242.800 107.600 243.600 108.400 ;
        RECT 233.200 105.600 234.000 106.400 ;
        RECT 234.800 105.600 235.600 106.400 ;
        RECT 236.400 105.600 237.200 106.400 ;
        RECT 241.200 105.600 242.000 106.400 ;
        RECT 231.600 95.600 232.400 96.400 ;
        RECT 231.700 94.300 232.300 95.600 ;
        RECT 233.300 94.300 233.900 105.600 ;
        RECT 234.900 94.400 235.500 105.600 ;
        RECT 242.900 104.400 243.500 107.600 ;
        RECT 238.000 103.600 238.800 104.400 ;
        RECT 242.800 103.600 243.600 104.400 ;
        RECT 247.600 103.600 248.400 104.400 ;
        RECT 238.100 94.400 238.700 103.600 ;
        RECT 247.700 98.400 248.300 103.600 ;
        RECT 239.600 97.600 240.400 98.400 ;
        RECT 247.600 97.600 248.400 98.400 ;
        RECT 239.700 94.400 240.300 97.600 ;
        RECT 244.400 95.600 245.200 96.400 ;
        RECT 231.700 94.000 233.900 94.300 ;
        RECT 231.600 93.700 233.900 94.000 ;
        RECT 231.600 93.200 232.400 93.700 ;
        RECT 234.800 93.600 235.600 94.400 ;
        RECT 238.000 93.600 238.800 94.400 ;
        RECT 239.600 93.600 240.400 94.400 ;
        RECT 241.200 93.600 242.000 94.400 ;
        RECT 241.300 92.400 241.900 93.600 ;
        RECT 239.600 91.600 240.400 92.400 ;
        RECT 241.200 91.600 242.000 92.400 ;
        RECT 244.500 90.400 245.100 95.600 ;
        RECT 234.800 89.600 235.600 90.400 ;
        RECT 244.400 89.600 245.200 90.400 ;
        RECT 246.000 79.600 246.800 80.400 ;
        RECT 238.000 71.600 238.800 72.400 ;
        RECT 238.100 70.400 238.700 71.600 ;
        RECT 238.000 69.600 238.800 70.400 ;
        RECT 246.100 68.400 246.700 79.600 ;
        RECT 247.600 70.300 248.400 70.400 ;
        RECT 249.300 70.300 249.900 117.600 ;
        RECT 250.900 116.400 251.500 123.600 ;
        RECT 250.800 115.600 251.600 116.400 ;
        RECT 250.800 111.200 251.600 112.400 ;
        RECT 252.400 104.200 253.200 117.800 ;
        RECT 254.000 104.200 254.800 117.800 ;
        RECT 255.600 104.200 256.400 115.800 ;
        RECT 257.300 112.400 257.900 123.600 ;
        RECT 262.100 118.400 262.700 131.600 ;
        RECT 265.200 127.600 266.000 128.400 ;
        RECT 265.300 122.400 265.900 127.600 ;
        RECT 265.200 121.600 266.000 122.400 ;
        RECT 266.900 120.400 267.500 149.600 ;
        RECT 266.800 119.600 267.600 120.400 ;
        RECT 262.000 117.600 262.800 118.400 ;
        RECT 257.200 111.600 258.000 112.400 ;
        RECT 257.200 107.600 258.000 108.400 ;
        RECT 257.300 106.400 257.900 107.600 ;
        RECT 257.200 105.600 258.000 106.400 ;
        RECT 258.800 104.200 259.600 115.800 ;
        RECT 260.400 113.600 261.200 114.400 ;
        RECT 260.500 110.400 261.100 113.600 ;
        RECT 260.400 109.600 261.200 110.400 ;
        RECT 260.500 106.400 261.100 109.600 ;
        RECT 260.400 105.600 261.200 106.400 ;
        RECT 260.500 100.400 261.100 105.600 ;
        RECT 262.000 104.200 262.800 115.800 ;
        RECT 263.600 104.200 264.400 117.800 ;
        RECT 265.200 104.200 266.000 117.800 ;
        RECT 266.800 104.200 267.600 117.800 ;
        RECT 271.700 102.400 272.300 153.600 ;
        RECT 273.200 144.200 274.000 157.800 ;
        RECT 274.800 144.200 275.600 157.800 ;
        RECT 276.400 144.200 277.200 155.800 ;
        RECT 278.100 154.400 278.700 169.600 ;
        RECT 284.400 163.600 285.200 164.400 ;
        RECT 284.500 160.400 285.100 163.600 ;
        RECT 281.200 159.600 282.000 160.400 ;
        RECT 284.400 159.600 285.200 160.400 ;
        RECT 278.000 153.600 278.800 154.400 ;
        RECT 278.000 147.600 278.800 148.400 ;
        RECT 279.600 144.200 280.400 155.800 ;
        RECT 281.300 146.400 281.900 159.600 ;
        RECT 281.200 145.600 282.000 146.400 ;
        RECT 281.300 140.400 281.900 145.600 ;
        RECT 282.800 144.200 283.600 155.800 ;
        RECT 284.400 144.200 285.200 157.800 ;
        RECT 286.000 144.200 286.800 157.800 ;
        RECT 287.600 144.200 288.400 157.800 ;
        RECT 292.500 156.400 293.100 185.600 ;
        RECT 294.100 184.400 294.700 189.600 ;
        RECT 295.600 187.600 296.400 188.400 ;
        RECT 294.000 183.600 294.800 184.400 ;
        RECT 297.300 174.400 297.900 213.600 ;
        RECT 300.500 198.400 301.100 217.600 ;
        RECT 318.000 215.600 318.800 216.400 ;
        RECT 302.000 213.600 302.800 214.400 ;
        RECT 318.100 212.400 318.700 215.600 ;
        RECT 318.000 211.600 318.800 212.400 ;
        RECT 310.000 204.300 310.800 204.400 ;
        RECT 310.000 203.700 312.300 204.300 ;
        RECT 319.600 204.200 320.400 217.800 ;
        RECT 321.200 204.200 322.000 217.800 ;
        RECT 322.800 204.200 323.600 217.800 ;
        RECT 324.400 206.200 325.200 217.800 ;
        RECT 326.100 216.400 326.700 223.600 ;
        RECT 326.000 215.600 326.800 216.400 ;
        RECT 327.600 206.200 328.400 217.800 ;
        RECT 329.300 214.400 329.900 243.600 ;
        RECT 334.100 226.400 334.700 253.600 ;
        RECT 335.700 250.400 336.300 281.600 ;
        RECT 337.300 256.400 337.900 311.600 ;
        RECT 338.800 303.600 339.600 304.400 ;
        RECT 338.800 295.600 339.600 296.400 ;
        RECT 338.900 276.400 339.500 295.600 ;
        RECT 340.500 280.400 341.100 321.600 ;
        RECT 342.000 311.600 342.800 312.400 ;
        RECT 342.100 286.400 342.700 311.600 ;
        RECT 345.300 292.400 345.900 345.600 ;
        RECT 346.800 344.200 347.600 357.800 ;
        RECT 348.400 344.200 349.200 357.800 ;
        RECT 350.000 344.200 350.800 355.800 ;
        RECT 351.600 347.600 352.400 348.400 ;
        RECT 351.700 346.400 352.300 347.600 ;
        RECT 351.600 345.600 352.400 346.400 ;
        RECT 353.200 344.200 354.000 355.800 ;
        RECT 354.800 345.600 355.600 346.400 ;
        RECT 354.900 342.300 355.500 345.600 ;
        RECT 356.400 344.200 357.200 355.800 ;
        RECT 358.000 344.200 358.800 357.800 ;
        RECT 359.600 344.200 360.400 357.800 ;
        RECT 361.200 344.200 362.000 357.800 ;
        RECT 362.800 349.600 363.600 350.400 ;
        RECT 353.300 341.700 355.500 342.300 ;
        RECT 353.300 338.400 353.900 341.700 ;
        RECT 346.800 324.200 347.600 337.800 ;
        RECT 348.400 324.200 349.200 337.800 ;
        RECT 350.000 324.200 350.800 337.800 ;
        RECT 351.600 326.200 352.400 337.800 ;
        RECT 353.200 337.600 354.000 338.400 ;
        RECT 353.300 336.400 353.900 337.600 ;
        RECT 353.200 335.600 354.000 336.400 ;
        RECT 354.800 326.200 355.600 337.800 ;
        RECT 356.400 333.600 357.200 334.400 ;
        RECT 358.000 326.200 358.800 337.800 ;
        RECT 359.600 324.200 360.400 337.800 ;
        RECT 361.200 324.200 362.000 337.800 ;
        RECT 362.900 332.400 363.500 349.600 ;
        RECT 362.800 331.600 363.600 332.400 ;
        RECT 364.400 331.600 365.200 332.400 ;
        RECT 359.600 317.600 360.400 318.400 ;
        RECT 358.000 313.600 358.800 314.400 ;
        RECT 348.400 311.600 349.200 312.400 ;
        RECT 351.600 309.600 352.400 310.400 ;
        RECT 346.800 307.600 347.600 308.400 ;
        RECT 348.400 295.600 349.200 296.400 ;
        RECT 348.500 292.400 349.100 295.600 ;
        RECT 351.700 294.400 352.300 309.600 ;
        RECT 356.400 305.600 357.200 306.400 ;
        RECT 358.100 304.300 358.700 313.600 ;
        RECT 359.700 310.400 360.300 317.600 ;
        RECT 364.500 310.400 365.100 331.600 ;
        RECT 359.600 309.600 360.400 310.400 ;
        RECT 364.400 309.600 365.200 310.400 ;
        RECT 356.500 303.700 358.700 304.300 ;
        RECT 351.600 294.300 352.400 294.400 ;
        RECT 351.600 293.700 353.900 294.300 ;
        RECT 351.600 293.600 352.400 293.700 ;
        RECT 345.200 291.600 346.000 292.400 ;
        RECT 348.400 291.600 349.200 292.400 ;
        RECT 346.800 289.600 347.600 290.400 ;
        RECT 351.600 289.600 352.400 290.400 ;
        RECT 346.900 286.400 347.500 289.600 ;
        RECT 342.000 285.600 342.800 286.400 ;
        RECT 346.800 285.600 347.600 286.400 ;
        RECT 340.400 279.600 341.200 280.400 ;
        RECT 338.800 275.600 339.600 276.400 ;
        RECT 343.600 273.600 344.400 274.400 ;
        RECT 345.200 273.600 346.000 274.400 ;
        RECT 340.400 267.600 341.200 268.400 ;
        RECT 343.600 267.600 344.400 268.400 ;
        RECT 337.200 255.600 338.000 256.400 ;
        RECT 338.800 255.600 339.600 256.400 ;
        RECT 335.600 249.600 336.400 250.400 ;
        RECT 335.700 234.400 336.300 249.600 ;
        RECT 337.300 248.400 337.900 255.600 ;
        RECT 338.900 254.400 339.500 255.600 ;
        RECT 338.800 253.600 339.600 254.400 ;
        RECT 337.200 247.600 338.000 248.400 ;
        RECT 335.600 233.600 336.400 234.400 ;
        RECT 338.900 232.400 339.500 253.600 ;
        RECT 340.500 238.400 341.100 267.600 ;
        RECT 342.000 263.600 342.800 264.400 ;
        RECT 342.100 254.400 342.700 263.600 ;
        RECT 342.000 253.600 342.800 254.400 ;
        RECT 342.000 252.300 342.800 252.400 ;
        RECT 343.700 252.300 344.300 267.600 ;
        RECT 342.000 251.700 344.300 252.300 ;
        RECT 342.000 251.600 342.800 251.700 ;
        RECT 343.600 250.300 344.400 250.400 ;
        RECT 345.300 250.300 345.900 273.600 ;
        RECT 346.900 272.400 347.500 285.600 ;
        RECT 346.800 271.600 347.600 272.400 ;
        RECT 348.400 271.600 349.200 272.400 ;
        RECT 351.600 271.600 352.400 272.400 ;
        RECT 348.500 270.400 349.100 271.600 ;
        RECT 351.700 270.400 352.300 271.600 ;
        RECT 353.300 270.400 353.900 293.700 ;
        RECT 354.800 293.600 355.600 294.400 ;
        RECT 354.900 292.400 355.500 293.600 ;
        RECT 354.800 291.600 355.600 292.400 ;
        RECT 356.500 288.400 357.100 303.700 ;
        RECT 359.600 303.600 360.400 304.400 ;
        RECT 359.700 298.400 360.300 303.600 ;
        RECT 359.600 297.600 360.400 298.400 ;
        RECT 359.600 291.600 360.400 292.400 ;
        RECT 361.200 291.600 362.000 292.400 ;
        RECT 359.700 290.400 360.300 291.600 ;
        RECT 359.600 289.600 360.400 290.400 ;
        RECT 354.800 287.600 355.600 288.400 ;
        RECT 356.400 287.600 357.200 288.400 ;
        RECT 354.900 286.400 355.500 287.600 ;
        RECT 354.800 285.600 355.600 286.400 ;
        RECT 356.500 274.400 357.100 287.600 ;
        RECT 359.700 276.400 360.300 289.600 ;
        RECT 362.800 283.600 363.600 284.400 ;
        RECT 361.200 277.600 362.000 278.400 ;
        RECT 359.600 275.600 360.400 276.400 ;
        RECT 356.400 273.600 357.200 274.400 ;
        RECT 356.400 271.600 357.200 272.400 ;
        RECT 359.600 272.300 360.400 272.400 ;
        RECT 361.300 272.300 361.900 277.600 ;
        RECT 359.600 271.700 361.900 272.300 ;
        RECT 359.600 271.600 360.400 271.700 ;
        RECT 348.400 269.600 349.200 270.400 ;
        RECT 350.000 269.600 350.800 270.400 ;
        RECT 351.600 269.600 352.400 270.400 ;
        RECT 353.200 269.600 354.000 270.400 ;
        RECT 354.800 269.600 355.600 270.400 ;
        RECT 359.600 269.600 360.400 270.400 ;
        RECT 346.800 265.600 347.600 266.400 ;
        RECT 346.900 254.400 347.500 265.600 ;
        RECT 350.100 258.300 350.700 269.600 ;
        RECT 354.900 268.400 355.500 269.600 ;
        RECT 353.200 267.600 354.000 268.400 ;
        RECT 354.800 267.600 355.600 268.400 ;
        RECT 362.900 268.300 363.500 283.600 ;
        RECT 364.500 282.400 365.100 309.600 ;
        RECT 367.700 294.400 368.300 359.600 ;
        RECT 380.400 351.600 381.200 352.400 ;
        RECT 380.500 348.400 381.100 351.600 ;
        RECT 382.100 350.400 382.700 399.600 ;
        RECT 383.700 398.400 384.300 411.600 ;
        RECT 394.900 410.400 395.500 411.600 ;
        RECT 391.600 409.600 392.400 410.400 ;
        RECT 393.200 409.600 394.000 410.400 ;
        RECT 394.800 409.600 395.600 410.400 ;
        RECT 391.700 408.400 392.300 409.600 ;
        RECT 396.500 408.400 397.100 411.600 ;
        RECT 391.600 407.600 392.400 408.400 ;
        RECT 394.800 407.600 395.600 408.400 ;
        RECT 396.400 407.600 397.200 408.400 ;
        RECT 394.900 406.400 395.500 407.600 ;
        RECT 394.800 405.600 395.600 406.400 ;
        RECT 398.100 406.300 398.700 427.600 ;
        RECT 407.600 421.600 408.400 422.400 ;
        RECT 399.600 419.600 400.400 420.400 ;
        RECT 399.700 410.400 400.300 419.600 ;
        RECT 401.300 415.700 405.100 416.300 ;
        RECT 401.300 414.400 401.900 415.700 ;
        RECT 401.200 413.600 402.000 414.400 ;
        RECT 402.800 413.600 403.600 414.400 ;
        RECT 404.500 414.300 405.100 415.700 ;
        RECT 406.000 414.300 406.800 414.400 ;
        RECT 404.500 413.700 406.800 414.300 ;
        RECT 406.000 413.600 406.800 413.700 ;
        RECT 402.900 412.400 403.500 413.600 ;
        RECT 407.700 412.400 408.300 421.600 ;
        RECT 409.300 418.400 409.900 427.600 ;
        RECT 409.200 417.600 410.000 418.400 ;
        RECT 410.800 417.600 411.600 418.400 ;
        RECT 412.500 416.400 413.100 433.600 ;
        RECT 414.100 432.400 414.700 437.600 ;
        RECT 415.600 434.300 416.400 434.400 ;
        RECT 417.300 434.300 417.900 449.600 ;
        RECT 420.400 443.600 421.200 444.400 ;
        RECT 420.500 438.400 421.100 443.600 ;
        RECT 420.400 437.600 421.200 438.400 ;
        RECT 415.600 433.700 417.900 434.300 ;
        RECT 415.600 433.600 416.400 433.700 ;
        RECT 414.000 431.600 414.800 432.400 ;
        RECT 414.000 429.600 414.800 430.400 ;
        RECT 420.400 424.200 421.200 435.800 ;
        RECT 412.400 415.600 413.200 416.400 ;
        RECT 415.600 415.600 416.400 416.400 ;
        RECT 417.200 415.600 418.000 416.400 ;
        RECT 422.100 416.300 422.700 451.700 ;
        RECT 426.800 451.600 427.600 452.400 ;
        RECT 430.100 450.400 430.700 453.600 ;
        RECT 431.600 451.600 432.400 452.400 ;
        RECT 423.600 449.600 424.400 450.400 ;
        RECT 430.000 449.600 430.800 450.400 ;
        RECT 420.500 415.700 422.700 416.300 ;
        RECT 415.700 412.400 416.300 415.600 ;
        RECT 417.300 412.400 417.900 415.600 ;
        RECT 401.200 411.600 402.000 412.400 ;
        RECT 402.800 411.600 403.600 412.400 ;
        RECT 406.000 411.600 406.800 412.400 ;
        RECT 407.600 411.600 408.400 412.400 ;
        RECT 410.800 411.600 411.600 412.400 ;
        RECT 415.600 411.600 416.400 412.400 ;
        RECT 417.200 411.600 418.000 412.400 ;
        RECT 401.300 410.400 401.900 411.600 ;
        RECT 399.600 409.600 400.400 410.400 ;
        RECT 401.200 409.600 402.000 410.400 ;
        RECT 402.900 408.400 403.500 411.600 ;
        RECT 410.900 410.400 411.500 411.600 ;
        RECT 420.500 410.400 421.100 415.700 ;
        RECT 422.000 413.600 422.800 414.400 ;
        RECT 422.100 412.400 422.700 413.600 ;
        RECT 422.000 411.600 422.800 412.400 ;
        RECT 410.800 409.600 411.600 410.400 ;
        RECT 420.400 409.600 421.200 410.400 ;
        RECT 423.700 408.400 424.300 449.600 ;
        RECT 431.700 446.400 432.300 451.600 ;
        RECT 434.900 450.400 435.500 461.600 ;
        RECT 436.400 453.600 437.200 454.400 ;
        RECT 439.600 453.600 440.400 454.400 ;
        RECT 434.800 449.600 435.600 450.400 ;
        RECT 436.500 448.400 437.100 453.600 ;
        RECT 438.000 451.600 438.800 452.400 ;
        RECT 444.400 451.600 445.200 452.400 ;
        RECT 436.400 447.600 437.200 448.400 ;
        RECT 431.600 445.600 432.400 446.400 ;
        RECT 426.800 443.600 427.600 444.400 ;
        RECT 431.600 443.600 432.400 444.400 ;
        RECT 434.800 443.600 435.600 444.400 ;
        RECT 425.200 429.600 426.000 430.400 ;
        RECT 425.200 427.600 426.000 428.400 ;
        RECT 402.800 407.600 403.600 408.400 ;
        RECT 423.600 407.600 424.400 408.400 ;
        RECT 396.500 405.700 398.700 406.300 ;
        RECT 396.500 398.400 397.100 405.700 ;
        RECT 399.600 405.600 400.400 406.400 ;
        RECT 399.700 398.400 400.300 405.600 ;
        RECT 423.600 403.600 424.400 404.400 ;
        RECT 383.600 397.600 384.400 398.400 ;
        RECT 393.200 397.600 394.000 398.400 ;
        RECT 396.400 397.600 397.200 398.400 ;
        RECT 399.600 397.600 400.400 398.400 ;
        RECT 386.800 389.600 387.600 390.400 ;
        RECT 386.900 382.400 387.500 389.600 ;
        RECT 388.400 384.200 389.200 395.800 ;
        RECT 409.200 393.600 410.000 394.400 ;
        RECT 401.200 389.600 402.000 390.400 ;
        RECT 394.800 385.600 395.600 386.400 ;
        RECT 398.000 385.600 398.800 386.400 ;
        RECT 386.800 381.600 387.600 382.400 ;
        RECT 394.900 380.400 395.500 385.600 ;
        RECT 396.400 381.600 397.200 382.400 ;
        RECT 394.800 379.600 395.600 380.400 ;
        RECT 390.000 364.200 390.800 377.800 ;
        RECT 391.600 364.200 392.400 377.800 ;
        RECT 393.200 364.200 394.000 377.800 ;
        RECT 394.800 366.200 395.600 377.800 ;
        RECT 396.500 376.400 397.100 381.600 ;
        RECT 398.100 380.400 398.700 385.600 ;
        RECT 404.400 383.600 405.200 384.400 ;
        RECT 409.200 383.600 410.000 384.400 ;
        RECT 418.800 384.200 419.600 397.800 ;
        RECT 420.400 384.200 421.200 397.800 ;
        RECT 422.000 384.200 422.800 397.800 ;
        RECT 423.600 384.200 424.400 395.800 ;
        RECT 425.300 386.400 425.900 427.600 ;
        RECT 426.900 420.400 427.500 443.600 ;
        RECT 430.000 424.200 430.800 435.800 ;
        RECT 426.800 419.600 427.600 420.400 ;
        RECT 428.400 417.600 429.200 418.400 ;
        RECT 428.500 414.400 429.100 417.600 ;
        RECT 428.400 413.600 429.200 414.400 ;
        RECT 430.000 412.300 430.800 412.400 ;
        RECT 431.700 412.300 432.300 443.600 ;
        RECT 433.200 426.200 434.000 431.800 ;
        RECT 434.900 426.400 435.500 443.600 ;
        RECT 438.100 430.300 438.700 451.600 ;
        RECT 441.200 449.600 442.000 450.400 ;
        RECT 444.400 450.300 445.200 450.400 ;
        RECT 446.100 450.300 446.700 467.600 ;
        RECT 444.400 449.700 446.700 450.300 ;
        RECT 447.700 450.300 448.300 475.600 ;
        RECT 452.500 468.400 453.100 491.600 ;
        RECT 454.100 484.400 454.700 491.600 ;
        RECT 455.700 490.400 456.300 501.600 ;
        RECT 457.300 496.400 457.900 503.600 ;
        RECT 457.200 495.600 458.000 496.400 ;
        RECT 465.300 496.300 465.900 503.600 ;
        RECT 476.400 497.600 477.200 498.400 ;
        RECT 463.700 495.700 465.900 496.300 ;
        RECT 463.700 490.400 464.300 495.700 ;
        RECT 471.600 495.600 472.400 496.400 ;
        RECT 476.500 494.400 477.100 497.600 ;
        RECT 479.700 494.400 480.300 505.600 ;
        RECT 481.200 503.600 482.000 504.400 ;
        RECT 465.200 493.600 466.000 494.400 ;
        RECT 473.200 493.600 474.000 494.400 ;
        RECT 476.400 493.600 477.200 494.400 ;
        RECT 479.600 493.600 480.400 494.400 ;
        RECT 455.600 489.600 456.400 490.400 ;
        RECT 463.600 489.600 464.400 490.400 ;
        RECT 454.000 483.600 454.800 484.400 ;
        RECT 455.600 483.600 456.400 484.400 ;
        RECT 452.400 467.600 453.200 468.400 ;
        RECT 450.800 451.600 451.600 452.400 ;
        RECT 449.200 450.300 450.000 450.400 ;
        RECT 447.700 449.700 450.000 450.300 ;
        RECT 444.400 449.600 445.200 449.700 ;
        RECT 449.200 449.600 450.000 449.700 ;
        RECT 441.300 444.400 441.900 449.600 ;
        RECT 446.000 447.600 446.800 448.400 ;
        RECT 450.900 448.300 451.500 451.600 ;
        RECT 449.300 447.700 451.500 448.300 ;
        RECT 441.200 443.600 442.000 444.400 ;
        RECT 444.400 443.600 445.200 444.400 ;
        RECT 444.500 434.300 445.100 443.600 ;
        RECT 442.900 433.700 445.100 434.300 ;
        RECT 442.900 432.400 443.500 433.700 ;
        RECT 442.800 431.600 443.600 432.400 ;
        RECT 439.600 430.300 440.400 430.400 ;
        RECT 438.100 429.700 440.400 430.300 ;
        RECT 434.800 425.600 435.600 426.400 ;
        RECT 438.100 422.400 438.700 429.700 ;
        RECT 439.600 429.600 440.400 429.700 ;
        RECT 444.400 426.200 445.200 431.800 ;
        RECT 446.000 427.600 446.800 428.400 ;
        RECT 442.800 423.600 443.600 424.400 ;
        RECT 447.600 424.200 448.400 435.800 ;
        RECT 438.000 421.600 438.800 422.400 ;
        RECT 436.400 415.600 437.200 416.400 ;
        RECT 441.200 415.600 442.000 416.400 ;
        RECT 434.800 413.600 435.600 414.400 ;
        RECT 436.500 412.400 437.100 415.600 ;
        RECT 430.000 411.700 432.300 412.300 ;
        RECT 430.000 411.600 430.800 411.700 ;
        RECT 436.400 411.600 437.200 412.400 ;
        RECT 441.300 410.400 441.900 415.600 ;
        RECT 442.900 414.400 443.500 423.600 ;
        RECT 444.400 417.600 445.200 418.400 ;
        RECT 442.800 413.600 443.600 414.400 ;
        RECT 444.500 412.400 445.100 417.600 ;
        RECT 449.300 416.400 449.900 447.700 ;
        RECT 452.400 447.600 453.200 448.400 ;
        RECT 450.800 443.600 451.600 444.400 ;
        RECT 452.500 436.400 453.100 447.600 ;
        RECT 454.100 446.400 454.700 483.600 ;
        RECT 465.300 472.400 465.900 493.600 ;
        RECT 466.800 491.600 467.600 492.400 ;
        RECT 466.800 489.600 467.600 490.400 ;
        RECT 470.000 489.600 470.800 490.400 ;
        RECT 466.900 478.400 467.500 489.600 ;
        RECT 470.100 488.400 470.700 489.600 ;
        RECT 470.000 487.600 470.800 488.400 ;
        RECT 471.600 481.600 472.400 482.400 ;
        RECT 466.800 477.600 467.600 478.400 ;
        RECT 465.200 471.600 466.000 472.400 ;
        RECT 466.900 470.400 467.500 477.600 ;
        RECT 468.400 473.600 469.200 474.400 ;
        RECT 460.400 469.600 461.200 470.400 ;
        RECT 465.200 469.600 466.000 470.400 ;
        RECT 466.800 469.600 467.600 470.400 ;
        RECT 460.500 464.400 461.100 469.600 ;
        RECT 465.300 468.400 465.900 469.600 ;
        RECT 468.500 468.400 469.100 473.600 ;
        RECT 471.700 472.400 472.300 481.600 ;
        RECT 471.600 471.600 472.400 472.400 ;
        RECT 465.200 467.600 466.000 468.400 ;
        RECT 468.400 467.600 469.200 468.400 ;
        RECT 471.700 466.400 472.300 471.600 ;
        RECT 473.300 468.400 473.900 493.600 ;
        RECT 474.800 491.600 475.600 492.400 ;
        RECT 474.900 490.400 475.500 491.600 ;
        RECT 474.800 489.600 475.600 490.400 ;
        RECT 474.800 469.600 475.600 470.400 ;
        RECT 473.200 467.600 474.000 468.400 ;
        RECT 471.600 465.600 472.400 466.400 ;
        RECT 460.400 463.600 461.200 464.400 ;
        RECT 470.000 463.600 470.800 464.400 ;
        RECT 460.500 458.400 461.100 463.600 ;
        RECT 460.400 457.600 461.200 458.400 ;
        RECT 455.600 455.600 456.400 456.400 ;
        RECT 470.100 456.300 470.700 463.600 ;
        RECT 471.600 461.600 472.400 462.400 ;
        RECT 468.500 455.700 470.700 456.300 ;
        RECT 463.600 451.600 464.400 452.400 ;
        RECT 463.700 446.400 464.300 451.600 ;
        RECT 468.500 450.400 469.100 455.700 ;
        RECT 470.000 453.600 470.800 454.400 ;
        RECT 471.700 452.400 472.300 461.600 ;
        RECT 474.900 454.400 475.500 469.600 ;
        RECT 476.500 456.400 477.100 493.600 ;
        RECT 478.000 487.600 478.800 488.400 ;
        RECT 478.100 484.400 478.700 487.600 ;
        RECT 478.000 483.600 478.800 484.400 ;
        RECT 478.100 482.400 478.700 483.600 ;
        RECT 478.000 481.600 478.800 482.400 ;
        RECT 481.300 474.400 481.900 503.600 ;
        RECT 482.800 486.200 483.600 497.800 ;
        RECT 478.000 473.600 478.800 474.400 ;
        RECT 481.200 473.600 482.000 474.400 ;
        RECT 478.100 472.400 478.700 473.600 ;
        RECT 478.000 471.600 478.800 472.400 ;
        RECT 481.200 471.600 482.000 472.400 ;
        RECT 484.500 470.400 485.100 513.600 ;
        RECT 487.700 510.400 488.300 527.600 ;
        RECT 489.300 518.400 489.900 531.600 ;
        RECT 494.000 529.600 494.800 530.400 ;
        RECT 498.800 529.600 499.600 530.400 ;
        RECT 500.400 530.200 501.200 535.800 ;
        RECT 502.100 534.400 502.700 541.600 ;
        RECT 502.000 533.600 502.800 534.400 ;
        RECT 494.100 528.400 494.700 529.600 ;
        RECT 490.800 527.600 491.600 528.400 ;
        RECT 494.000 527.600 494.800 528.400 ;
        RECT 489.200 517.600 490.000 518.400 ;
        RECT 490.900 512.400 491.500 527.600 ;
        RECT 498.900 518.400 499.500 529.600 ;
        RECT 503.600 526.200 504.400 537.800 ;
        RECT 505.200 531.600 506.000 532.600 ;
        RECT 513.200 526.200 514.000 537.800 ;
        RECT 514.900 534.400 515.500 549.600 ;
        RECT 518.000 547.600 518.800 548.400 ;
        RECT 514.800 533.600 515.600 534.400 ;
        RECT 519.700 532.400 520.300 549.600 ;
        RECT 522.900 546.400 523.500 551.700 ;
        RECT 529.200 551.600 530.000 552.400 ;
        RECT 532.400 551.600 533.200 552.400 ;
        RECT 526.000 549.600 526.800 550.400 ;
        RECT 527.600 549.600 528.400 550.400 ;
        RECT 522.800 545.600 523.600 546.400 ;
        RECT 522.900 534.400 523.500 545.600 ;
        RECT 526.100 536.400 526.700 549.600 ;
        RECT 527.700 548.400 528.300 549.600 ;
        RECT 529.300 548.400 529.900 551.600 ;
        RECT 532.400 549.600 533.200 550.400 ;
        RECT 527.600 547.600 528.400 548.400 ;
        RECT 529.200 547.600 530.000 548.400 ;
        RECT 534.000 547.600 534.800 548.400 ;
        RECT 527.600 543.600 528.400 544.400 ;
        RECT 527.700 538.400 528.300 543.600 ;
        RECT 532.400 541.600 533.200 542.400 ;
        RECT 527.600 537.600 528.400 538.400 ;
        RECT 526.000 535.600 526.800 536.400 ;
        RECT 522.800 533.600 523.600 534.400 ;
        RECT 519.600 531.600 520.400 532.400 ;
        RECT 522.800 531.600 523.600 532.400 ;
        RECT 530.800 531.600 531.600 532.400 ;
        RECT 519.600 529.600 520.400 530.400 ;
        RECT 518.000 527.600 518.800 528.400 ;
        RECT 519.700 522.400 520.300 529.600 ;
        RECT 521.200 523.600 522.000 524.400 ;
        RECT 519.600 521.600 520.400 522.400 ;
        RECT 521.300 520.400 521.900 523.600 ;
        RECT 516.400 519.600 517.200 520.400 ;
        RECT 521.200 519.600 522.000 520.400 ;
        RECT 498.800 517.600 499.600 518.400 ;
        RECT 503.600 517.600 504.400 518.400 ;
        RECT 490.800 511.600 491.600 512.400 ;
        RECT 490.900 510.400 491.500 511.600 ;
        RECT 498.900 510.400 499.500 517.600 ;
        RECT 503.700 514.400 504.300 517.600 ;
        RECT 503.600 513.600 504.400 514.400 ;
        RECT 505.200 513.600 506.000 514.400 ;
        RECT 505.300 510.400 505.900 513.600 ;
        RECT 516.500 512.400 517.100 519.600 ;
        RECT 522.900 514.400 523.500 531.600 ;
        RECT 530.900 530.400 531.500 531.600 ;
        RECT 530.800 529.600 531.600 530.400 ;
        RECT 522.800 513.600 523.600 514.400 ;
        RECT 511.600 511.600 512.400 512.400 ;
        RECT 516.400 511.600 517.200 512.400 ;
        RECT 518.000 511.600 518.800 512.400 ;
        RECT 522.800 511.600 523.600 512.400 ;
        RECT 526.000 512.300 526.800 512.400 ;
        RECT 526.000 511.700 529.900 512.300 ;
        RECT 526.000 511.600 526.800 511.700 ;
        RECT 486.000 509.600 486.800 510.400 ;
        RECT 487.600 509.600 488.400 510.400 ;
        RECT 490.800 509.600 491.600 510.400 ;
        RECT 494.000 509.600 494.800 510.400 ;
        RECT 498.800 509.600 499.600 510.400 ;
        RECT 505.200 509.600 506.000 510.400 ;
        RECT 510.000 509.600 510.800 510.400 ;
        RECT 486.100 476.400 486.700 509.600 ;
        RECT 490.800 501.600 491.600 502.400 ;
        RECT 490.900 496.400 491.500 501.600 ;
        RECT 489.200 495.600 490.000 496.400 ;
        RECT 490.800 495.600 491.600 496.400 ;
        RECT 489.300 492.400 489.900 495.600 ;
        RECT 489.200 491.600 490.000 492.400 ;
        RECT 489.200 489.600 490.000 490.400 ;
        RECT 489.300 478.400 489.900 489.600 ;
        RECT 492.400 486.200 493.200 497.800 ;
        RECT 494.100 484.400 494.700 509.600 ;
        RECT 500.400 507.600 501.200 508.400 ;
        RECT 500.500 506.400 501.100 507.600 ;
        RECT 500.400 505.600 501.200 506.400 ;
        RECT 495.600 503.600 496.400 504.400 ;
        RECT 495.700 498.400 496.300 503.600 ;
        RECT 495.600 497.600 496.400 498.400 ;
        RECT 495.600 490.200 496.400 495.800 ;
        RECT 500.500 494.400 501.100 505.600 ;
        RECT 503.600 503.600 504.400 504.400 ;
        RECT 506.800 503.600 507.600 504.400 ;
        RECT 508.400 503.600 509.200 504.400 ;
        RECT 503.700 496.400 504.300 503.600 ;
        RECT 506.900 498.400 507.500 503.600 ;
        RECT 508.500 500.400 509.100 503.600 ;
        RECT 508.400 499.600 509.200 500.400 ;
        RECT 506.800 497.600 507.600 498.400 ;
        RECT 503.600 495.600 504.400 496.400 ;
        RECT 506.900 494.400 507.500 497.600 ;
        RECT 500.400 493.600 501.200 494.400 ;
        RECT 506.800 493.600 507.600 494.400 ;
        RECT 497.200 491.600 498.000 492.400 ;
        RECT 498.800 491.600 499.600 492.400 ;
        RECT 497.300 490.400 497.900 491.600 ;
        RECT 497.200 489.600 498.000 490.400 ;
        RECT 492.400 483.600 493.200 484.400 ;
        RECT 494.000 483.600 494.800 484.400 ;
        RECT 489.200 477.600 490.000 478.400 ;
        RECT 486.000 475.600 486.800 476.400 ;
        RECT 487.600 476.300 488.400 476.400 ;
        RECT 487.600 475.700 489.900 476.300 ;
        RECT 487.600 475.600 488.400 475.700 ;
        RECT 486.000 471.600 486.800 472.400 ;
        RECT 486.100 470.400 486.700 471.600 ;
        RECT 487.700 470.400 488.300 475.600 ;
        RECT 482.800 469.600 483.600 470.400 ;
        RECT 484.400 469.600 485.200 470.400 ;
        RECT 486.000 469.600 486.800 470.400 ;
        RECT 487.600 469.600 488.400 470.400 ;
        RECT 478.000 463.600 478.800 464.400 ;
        RECT 476.400 455.600 477.200 456.400 ;
        RECT 481.200 455.600 482.000 456.400 ;
        RECT 481.300 454.400 481.900 455.600 ;
        RECT 474.800 453.600 475.600 454.400 ;
        RECT 476.400 453.600 477.200 454.400 ;
        RECT 479.600 453.600 480.400 454.400 ;
        RECT 481.200 453.600 482.000 454.400 ;
        RECT 471.600 451.600 472.400 452.400 ;
        RECT 474.800 451.600 475.600 452.400 ;
        RECT 474.900 450.400 475.500 451.600 ;
        RECT 468.400 449.600 469.200 450.400 ;
        RECT 471.600 449.600 472.400 450.400 ;
        RECT 474.800 449.600 475.600 450.400 ;
        RECT 454.000 445.600 454.800 446.400 ;
        RECT 463.600 445.600 464.400 446.400 ;
        RECT 454.000 437.600 454.800 438.400 ;
        RECT 452.400 435.600 453.200 436.400 ;
        RECT 450.800 429.600 451.600 430.400 ;
        RECT 450.900 418.400 451.500 429.600 ;
        RECT 450.800 417.600 451.600 418.400 ;
        RECT 449.200 415.600 450.000 416.400 ;
        RECT 449.300 414.400 449.900 415.600 ;
        RECT 452.500 414.400 453.100 435.600 ;
        RECT 454.100 430.400 454.700 437.600 ;
        RECT 454.000 429.600 454.800 430.400 ;
        RECT 457.200 424.200 458.000 435.800 ;
        RECT 462.000 433.600 462.800 434.400 ;
        RECT 457.200 415.600 458.000 416.400 ;
        RECT 449.200 413.600 450.000 414.400 ;
        RECT 452.400 413.600 453.200 414.400 ;
        RECT 444.400 411.600 445.200 412.400 ;
        RECT 457.300 410.400 457.900 415.600 ;
        RECT 460.400 413.600 461.200 414.400 ;
        RECT 463.700 412.400 464.300 445.600 ;
        RECT 465.200 443.600 466.000 444.400 ;
        RECT 465.300 418.400 465.900 443.600 ;
        RECT 471.700 438.400 472.300 449.600 ;
        RECT 471.600 437.600 472.400 438.400 ;
        RECT 470.000 435.600 470.800 436.400 ;
        RECT 470.100 434.400 470.700 435.600 ;
        RECT 474.900 434.400 475.500 449.600 ;
        RECT 476.500 438.400 477.100 453.600 ;
        RECT 479.700 452.400 480.300 453.600 ;
        RECT 482.900 452.400 483.500 469.600 ;
        RECT 484.500 456.400 485.100 469.600 ;
        RECT 486.100 460.400 486.700 469.600 ;
        RECT 486.000 459.600 486.800 460.400 ;
        RECT 484.400 455.600 485.200 456.400 ;
        RECT 486.000 455.600 486.800 456.400 ;
        RECT 486.100 454.400 486.700 455.600 ;
        RECT 486.000 453.600 486.800 454.400 ;
        RECT 489.300 452.400 489.900 475.700 ;
        RECT 492.500 452.400 493.100 483.600 ;
        RECT 494.100 478.400 494.700 483.600 ;
        RECT 495.600 481.600 496.400 482.400 ;
        RECT 494.000 477.600 494.800 478.400 ;
        RECT 495.700 470.400 496.300 481.600 ;
        RECT 497.300 472.400 497.900 489.600 ;
        RECT 498.900 488.400 499.500 491.600 ;
        RECT 498.800 487.600 499.600 488.400 ;
        RECT 497.200 471.600 498.000 472.400 ;
        RECT 500.500 472.300 501.100 493.600 ;
        RECT 503.600 491.600 504.400 492.400 ;
        RECT 503.700 488.400 504.300 491.600 ;
        RECT 506.800 489.600 507.600 490.400 ;
        RECT 502.000 487.600 502.800 488.400 ;
        RECT 503.600 487.600 504.400 488.400 ;
        RECT 498.900 471.700 501.100 472.300 ;
        RECT 495.600 469.600 496.400 470.400 ;
        RECT 495.700 466.400 496.300 469.600 ;
        RECT 498.900 468.400 499.500 471.700 ;
        RECT 502.100 470.400 502.700 487.600 ;
        RECT 506.900 478.400 507.500 489.600 ;
        RECT 506.800 477.600 507.600 478.400 ;
        RECT 503.600 471.600 504.400 472.400 ;
        RECT 508.400 471.600 509.200 472.400 ;
        RECT 500.400 469.600 501.200 470.400 ;
        RECT 502.000 469.600 502.800 470.400 ;
        RECT 500.500 468.400 501.100 469.600 ;
        RECT 502.100 468.400 502.700 469.600 ;
        RECT 498.800 467.600 499.600 468.400 ;
        RECT 500.400 467.600 501.200 468.400 ;
        RECT 502.000 467.600 502.800 468.400 ;
        RECT 505.200 467.600 506.000 468.400 ;
        RECT 495.600 465.600 496.400 466.400 ;
        RECT 497.200 463.600 498.000 464.400 ;
        RECT 497.300 454.400 497.900 463.600 ;
        RECT 505.300 458.400 505.900 467.600 ;
        RECT 506.800 465.600 507.600 466.400 ;
        RECT 506.900 458.400 507.500 465.600 ;
        RECT 505.200 457.600 506.000 458.400 ;
        RECT 506.800 457.600 507.600 458.400 ;
        RECT 508.400 455.600 509.200 456.400 ;
        RECT 494.000 453.600 494.800 454.400 ;
        RECT 497.200 453.600 498.000 454.400 ;
        RECT 498.800 453.600 499.600 454.400 ;
        RECT 505.200 453.600 506.000 454.400 ;
        RECT 508.500 452.400 509.100 455.600 ;
        RECT 479.600 451.600 480.400 452.400 ;
        RECT 482.800 451.600 483.600 452.400 ;
        RECT 484.400 451.600 485.200 452.400 ;
        RECT 489.200 451.600 490.000 452.400 ;
        RECT 492.400 451.600 493.200 452.400 ;
        RECT 495.600 451.600 496.400 452.400 ;
        RECT 500.400 451.600 501.200 452.400 ;
        RECT 505.200 451.600 506.000 452.400 ;
        RECT 508.400 451.600 509.200 452.400 ;
        RECT 492.400 449.600 493.200 450.400 ;
        RECT 495.700 444.400 496.300 451.600 ;
        RECT 503.600 449.600 504.400 450.400 ;
        RECT 495.600 443.600 496.400 444.400 ;
        RECT 476.400 437.600 477.200 438.400 ;
        RECT 470.000 433.600 470.800 434.400 ;
        RECT 474.800 433.600 475.600 434.400 ;
        RECT 474.900 432.400 475.500 433.600 ;
        RECT 474.800 431.600 475.600 432.400 ;
        RECT 471.600 429.600 472.400 430.400 ;
        RECT 465.200 417.600 466.000 418.400 ;
        RECT 471.700 416.400 472.300 429.600 ;
        RECT 481.200 427.600 482.000 428.400 ;
        RECT 481.300 418.400 481.900 427.600 ;
        RECT 486.000 424.200 486.800 437.800 ;
        RECT 487.600 424.200 488.400 437.800 ;
        RECT 489.200 424.200 490.000 437.800 ;
        RECT 490.800 424.200 491.600 435.800 ;
        RECT 492.400 425.600 493.200 426.400 ;
        RECT 494.000 424.200 494.800 435.800 ;
        RECT 495.700 430.400 496.300 443.600 ;
        RECT 495.600 429.600 496.400 430.400 ;
        RECT 495.600 427.600 496.400 428.400 ;
        RECT 497.200 424.200 498.000 435.800 ;
        RECT 498.800 424.200 499.600 437.800 ;
        RECT 500.400 424.200 501.200 437.800 ;
        RECT 498.800 419.600 499.600 420.400 ;
        RECT 481.200 417.600 482.000 418.400 ;
        RECT 498.900 416.400 499.500 419.600 ;
        RECT 471.600 415.600 472.400 416.400 ;
        RECT 476.400 415.000 477.200 415.800 ;
        RECT 477.800 415.000 482.000 415.600 ;
        RECT 483.000 415.000 483.800 415.800 ;
        RECT 490.800 415.600 491.600 416.400 ;
        RECT 498.800 415.600 499.600 416.400 ;
        RECT 466.800 413.600 467.600 414.400 ;
        RECT 473.200 413.600 474.000 414.400 ;
        RECT 474.800 413.600 475.600 414.400 ;
        RECT 476.400 414.200 477.000 415.000 ;
        RECT 477.800 414.800 478.600 415.000 ;
        RECT 481.200 414.800 482.000 415.000 ;
        RECT 476.400 413.600 481.200 414.200 ;
        RECT 463.600 411.600 464.400 412.400 ;
        RECT 465.200 411.600 466.000 412.400 ;
        RECT 471.600 411.600 472.400 412.400 ;
        RECT 426.800 409.600 427.600 410.400 ;
        RECT 433.200 409.600 434.000 410.400 ;
        RECT 441.200 409.600 442.000 410.400 ;
        RECT 447.600 409.600 448.400 410.400 ;
        RECT 457.200 409.600 458.000 410.400 ;
        RECT 426.900 408.400 427.500 409.600 ;
        RECT 433.300 408.400 433.900 409.600 ;
        RECT 465.300 408.400 465.900 411.600 ;
        RECT 468.400 409.600 469.200 410.400 ;
        RECT 426.800 407.600 427.600 408.400 ;
        RECT 433.200 407.600 434.000 408.400 ;
        RECT 465.200 407.600 466.000 408.400 ;
        RECT 465.200 406.300 466.000 406.400 ;
        RECT 468.500 406.300 469.100 409.600 ;
        RECT 473.300 408.400 473.900 413.600 ;
        RECT 476.400 410.200 477.000 413.600 ;
        RECT 480.400 413.400 481.200 413.600 ;
        RECT 483.200 410.200 483.800 415.000 ;
        RECT 484.400 413.600 485.200 414.400 ;
        RECT 484.500 410.400 485.100 413.600 ;
        RECT 489.200 411.600 490.000 412.400 ;
        RECT 476.400 409.400 477.200 410.200 ;
        RECT 483.000 409.400 483.800 410.200 ;
        RECT 484.400 409.600 485.200 410.400 ;
        RECT 486.000 409.600 486.800 410.400 ;
        RECT 473.200 407.600 474.000 408.400 ;
        RECT 465.200 405.700 469.100 406.300 ;
        RECT 465.200 405.600 466.000 405.700 ;
        RECT 430.000 403.600 430.800 404.400 ;
        RECT 444.400 403.600 445.200 404.400 ;
        RECT 471.600 403.600 472.400 404.400 ;
        RECT 430.100 398.400 430.700 403.600 ;
        RECT 430.000 397.600 430.800 398.400 ;
        RECT 425.200 385.600 426.000 386.400 ;
        RECT 425.300 384.400 425.900 385.600 ;
        RECT 425.200 383.600 426.000 384.400 ;
        RECT 426.800 384.200 427.600 395.800 ;
        RECT 428.400 387.600 429.200 388.400 ;
        RECT 430.000 384.200 430.800 395.800 ;
        RECT 431.600 384.200 432.400 397.800 ;
        RECT 433.200 384.200 434.000 397.800 ;
        RECT 442.800 397.600 443.600 398.400 ;
        RECT 442.900 392.400 443.500 397.600 ;
        RECT 442.800 391.600 443.600 392.400 ;
        RECT 438.000 389.600 438.800 390.400 ;
        RECT 404.500 380.400 405.100 383.600 ;
        RECT 398.000 379.600 398.800 380.400 ;
        RECT 404.400 379.600 405.200 380.400 ;
        RECT 396.400 375.600 397.200 376.400 ;
        RECT 398.000 366.200 398.800 377.800 ;
        RECT 399.600 373.600 400.400 374.400 ;
        RECT 401.200 366.200 402.000 377.800 ;
        RECT 402.800 364.200 403.600 377.800 ;
        RECT 404.400 364.200 405.200 377.800 ;
        RECT 407.600 377.600 408.400 378.400 ;
        RECT 407.700 372.400 408.300 377.600 ;
        RECT 407.600 371.600 408.400 372.400 ;
        RECT 393.200 353.600 394.000 354.400 ;
        RECT 393.300 350.400 393.900 353.600 ;
        RECT 394.800 351.600 395.600 352.400 ;
        RECT 401.200 351.600 402.000 352.400 ;
        RECT 407.600 351.600 408.400 352.400 ;
        RECT 409.300 350.400 409.900 383.600 ;
        RECT 431.600 381.600 432.400 382.400 ;
        RECT 417.200 375.600 418.000 376.400 ;
        RECT 431.700 374.400 432.300 381.600 ;
        RECT 438.100 378.400 438.700 389.600 ;
        RECT 442.800 387.600 443.600 388.400 ;
        RECT 444.500 386.400 445.100 403.600 ;
        RECT 446.000 393.600 446.800 394.400 ;
        RECT 450.800 389.600 451.600 390.400 ;
        RECT 444.400 385.600 445.200 386.400 ;
        RECT 438.000 377.600 438.800 378.400 ;
        RECT 418.800 373.600 419.600 374.400 ;
        RECT 431.600 373.600 432.400 374.400 ;
        RECT 420.400 371.600 421.200 372.400 ;
        RECT 433.200 371.600 434.000 372.400 ;
        RECT 420.500 370.400 421.100 371.600 ;
        RECT 444.500 370.400 445.100 385.600 ;
        RECT 447.600 373.600 448.400 374.400 ;
        RECT 450.900 372.400 451.500 389.600 ;
        RECT 452.400 387.600 453.200 388.400 ;
        RECT 452.500 382.400 453.100 387.600 ;
        RECT 466.800 384.200 467.600 397.800 ;
        RECT 468.400 384.200 469.200 397.800 ;
        RECT 470.000 384.200 470.800 395.800 ;
        RECT 471.700 388.400 472.300 403.600 ;
        RECT 484.500 400.400 485.100 409.600 ;
        RECT 486.100 408.400 486.700 409.600 ;
        RECT 486.000 407.600 486.800 408.400 ;
        RECT 489.200 403.600 490.000 404.400 ;
        RECT 484.400 399.600 485.200 400.400 ;
        RECT 471.600 387.600 472.400 388.400 ;
        RECT 473.200 384.200 474.000 395.800 ;
        RECT 474.800 387.600 475.600 388.400 ;
        RECT 474.900 386.400 475.500 387.600 ;
        RECT 474.800 385.600 475.600 386.400 ;
        RECT 474.900 384.400 475.500 385.600 ;
        RECT 474.800 383.600 475.600 384.400 ;
        RECT 476.400 384.200 477.200 395.800 ;
        RECT 478.000 384.200 478.800 397.800 ;
        RECT 479.600 384.200 480.400 397.800 ;
        RECT 481.200 384.200 482.000 397.800 ;
        RECT 489.300 392.400 489.900 403.600 ;
        RECT 490.900 398.400 491.500 415.600 ;
        RECT 495.600 413.200 496.400 414.400 ;
        RECT 502.000 413.600 502.800 414.400 ;
        RECT 498.800 411.600 499.600 412.400 ;
        RECT 502.100 410.400 502.700 413.600 ;
        RECT 502.000 409.600 502.800 410.400 ;
        RECT 503.700 400.400 504.300 449.600 ;
        RECT 505.300 448.400 505.900 451.600 ;
        RECT 505.200 447.600 506.000 448.400 ;
        RECT 505.300 436.400 505.900 447.600 ;
        RECT 505.200 435.600 506.000 436.400 ;
        RECT 505.200 429.600 506.000 430.400 ;
        RECT 508.500 416.400 509.100 451.600 ;
        RECT 510.100 446.400 510.700 509.600 ;
        RECT 511.700 508.400 512.300 511.600 ;
        RECT 522.900 510.400 523.500 511.600 ;
        RECT 529.300 510.400 529.900 511.700 ;
        RECT 521.200 509.600 522.000 510.400 ;
        RECT 522.800 509.600 523.600 510.400 ;
        RECT 527.600 509.600 528.400 510.400 ;
        RECT 529.200 509.600 530.000 510.400 ;
        RECT 521.300 508.400 521.900 509.600 ;
        RECT 511.600 507.600 512.400 508.400 ;
        RECT 521.200 507.600 522.000 508.400 ;
        RECT 519.600 505.600 520.400 506.400 ;
        RECT 516.400 503.600 517.200 504.400 ;
        RECT 516.500 498.400 517.100 503.600 ;
        RECT 518.000 499.600 518.800 500.400 ;
        RECT 516.400 497.600 517.200 498.400 ;
        RECT 511.600 495.600 512.400 496.400 ;
        RECT 518.100 494.400 518.700 499.600 ;
        RECT 518.000 493.600 518.800 494.400 ;
        RECT 516.400 491.600 517.200 492.400 ;
        RECT 521.300 490.400 521.900 507.600 ;
        RECT 522.900 506.400 523.500 509.600 ;
        RECT 527.700 508.400 528.300 509.600 ;
        RECT 527.600 507.600 528.400 508.400 ;
        RECT 529.200 507.600 530.000 508.400 ;
        RECT 522.800 505.600 523.600 506.400 ;
        RECT 527.700 502.300 528.300 507.600 ;
        RECT 529.300 504.400 529.900 507.600 ;
        RECT 529.200 503.600 530.000 504.400 ;
        RECT 526.100 501.700 528.300 502.300 ;
        RECT 511.600 489.600 512.400 490.400 ;
        RECT 513.200 489.600 514.000 490.400 ;
        RECT 521.200 489.600 522.000 490.400 ;
        RECT 522.800 489.600 523.600 490.400 ;
        RECT 511.700 478.400 512.300 489.600 ;
        RECT 513.300 488.400 513.900 489.600 ;
        RECT 513.200 487.600 514.000 488.400 ;
        RECT 519.600 487.600 520.400 488.400 ;
        RECT 516.400 483.600 517.200 484.400 ;
        RECT 516.500 478.400 517.100 483.600 ;
        RECT 511.600 477.600 512.400 478.400 ;
        RECT 516.400 477.600 517.200 478.400 ;
        RECT 518.000 473.600 518.800 474.400 ;
        RECT 518.100 470.400 518.700 473.600 ;
        RECT 518.000 469.600 518.800 470.400 ;
        RECT 519.600 469.600 520.400 470.400 ;
        RECT 521.200 469.600 522.000 470.400 ;
        RECT 514.800 465.600 515.600 466.400 ;
        RECT 514.900 458.400 515.500 465.600 ;
        RECT 521.300 460.400 521.900 469.600 ;
        RECT 521.200 459.600 522.000 460.400 ;
        RECT 514.800 457.600 515.600 458.400 ;
        RECT 522.900 456.400 523.500 489.600 ;
        RECT 524.400 486.200 525.200 497.800 ;
        RECT 524.400 483.600 525.200 484.400 ;
        RECT 524.500 478.400 525.100 483.600 ;
        RECT 524.400 477.600 525.200 478.400 ;
        RECT 526.100 470.400 526.700 501.700 ;
        RECT 527.600 497.600 528.400 498.400 ;
        RECT 526.000 469.600 526.800 470.400 ;
        RECT 526.100 468.400 526.700 469.600 ;
        RECT 526.000 467.600 526.800 468.400 ;
        RECT 522.800 455.600 523.600 456.400 ;
        RECT 513.200 451.600 514.000 452.400 ;
        RECT 514.800 451.600 515.600 452.400 ;
        RECT 518.000 451.600 518.800 452.400 ;
        RECT 519.600 451.600 520.400 452.400 ;
        RECT 527.700 452.300 528.300 497.600 ;
        RECT 529.200 495.600 530.000 496.400 ;
        RECT 529.300 492.400 529.900 495.600 ;
        RECT 529.200 491.600 530.000 492.400 ;
        RECT 529.200 471.600 530.000 472.400 ;
        RECT 530.900 472.300 531.500 529.600 ;
        RECT 532.500 502.400 533.100 541.600 ;
        RECT 534.100 538.400 534.700 547.600 ;
        RECT 538.800 545.600 539.600 546.400 ;
        RECT 538.900 544.400 539.500 545.600 ;
        RECT 537.200 543.600 538.000 544.400 ;
        RECT 538.800 543.600 539.600 544.400 ;
        RECT 543.600 544.200 544.400 555.800 ;
        RECT 550.000 551.600 550.800 552.400 ;
        RECT 550.100 550.400 550.700 551.600 ;
        RECT 550.000 549.600 550.800 550.400 ;
        RECT 545.200 547.600 546.000 548.400 ;
        RECT 534.000 537.600 534.800 538.400 ;
        RECT 537.300 534.400 537.900 543.600 ;
        RECT 545.300 542.400 545.900 547.600 ;
        RECT 553.200 544.200 554.000 555.800 ;
        RECT 554.800 547.600 555.600 548.400 ;
        RECT 554.900 546.400 555.500 547.600 ;
        RECT 554.800 545.600 555.600 546.400 ;
        RECT 556.400 546.200 557.200 551.800 ;
        RECT 561.200 545.600 562.000 546.400 ;
        RECT 559.600 543.600 560.400 544.400 ;
        RECT 545.200 541.600 546.000 542.400 ;
        RECT 538.800 539.600 539.600 540.400 ;
        RECT 537.200 533.600 538.000 534.400 ;
        RECT 538.900 532.400 539.500 539.600 ;
        RECT 543.600 535.600 544.400 536.400 ;
        RECT 538.800 531.600 539.600 532.400 ;
        RECT 543.600 529.600 544.400 530.400 ;
        RECT 542.000 515.600 542.800 516.400 ;
        RECT 535.600 513.600 536.400 514.400 ;
        RECT 535.700 512.400 536.300 513.600 ;
        RECT 542.100 512.400 542.700 515.600 ;
        RECT 535.600 511.600 536.400 512.400 ;
        RECT 542.000 511.600 542.800 512.400 ;
        RECT 543.700 510.400 544.300 529.600 ;
        RECT 545.200 523.600 546.000 524.400 ;
        RECT 554.800 524.200 555.600 537.800 ;
        RECT 556.400 524.200 557.200 537.800 ;
        RECT 558.000 524.200 558.800 537.800 ;
        RECT 559.600 526.200 560.400 537.800 ;
        RECT 561.300 536.400 561.900 545.600 ;
        RECT 569.200 544.200 570.000 557.800 ;
        RECT 570.800 544.200 571.600 557.800 ;
        RECT 572.400 544.200 573.200 557.800 ;
        RECT 574.000 544.200 574.800 555.800 ;
        RECT 575.600 545.600 576.400 546.400 ;
        RECT 577.200 544.200 578.000 555.800 ;
        RECT 578.800 547.600 579.600 548.400 ;
        RECT 580.400 544.200 581.200 555.800 ;
        RECT 582.000 544.200 582.800 557.800 ;
        RECT 583.600 544.200 584.400 557.800 ;
        RECT 591.600 555.600 592.400 556.400 ;
        RECT 607.600 555.600 608.400 556.400 ;
        RECT 588.400 549.600 589.200 550.400 ;
        RECT 586.800 545.600 587.600 546.400 ;
        RECT 586.900 538.400 587.500 545.600 ;
        RECT 561.200 535.600 562.000 536.400 ;
        RECT 562.800 526.200 563.600 537.800 ;
        RECT 564.400 535.600 565.200 536.400 ;
        RECT 564.500 534.400 565.100 535.600 ;
        RECT 564.400 533.600 565.200 534.400 ;
        RECT 566.000 526.200 566.800 537.800 ;
        RECT 567.600 524.200 568.400 537.800 ;
        RECT 569.200 524.200 570.000 537.800 ;
        RECT 586.800 537.600 587.600 538.400 ;
        RECT 578.800 533.600 579.600 534.400 ;
        RECT 572.400 531.600 573.200 532.400 ;
        RECT 580.400 531.600 581.200 532.400 ;
        RECT 582.000 531.600 582.800 532.400 ;
        RECT 572.500 524.400 573.100 531.600 ;
        RECT 572.400 523.600 573.200 524.400 ;
        RECT 545.300 516.400 545.900 523.600 ;
        RECT 575.600 517.600 576.400 518.400 ;
        RECT 545.200 515.600 546.000 516.400 ;
        RECT 545.200 513.600 546.000 514.400 ;
        RECT 548.400 511.600 549.200 512.400 ;
        RECT 538.800 509.600 539.600 510.400 ;
        RECT 543.600 509.600 544.400 510.400 ;
        RECT 545.200 510.300 546.000 510.400 ;
        RECT 545.200 509.700 547.500 510.300 ;
        RECT 545.200 509.600 546.000 509.700 ;
        RECT 537.200 507.600 538.000 508.400 ;
        RECT 543.600 507.600 544.400 508.400 ;
        RECT 535.600 505.600 536.400 506.400 ;
        RECT 532.400 501.600 533.200 502.400 ;
        RECT 532.500 496.400 533.100 501.600 ;
        RECT 537.300 500.400 537.900 507.600 ;
        RECT 538.800 503.600 539.600 504.400 ;
        RECT 537.200 499.600 538.000 500.400 ;
        RECT 532.400 495.600 533.200 496.400 ;
        RECT 534.000 486.200 534.800 497.800 ;
        RECT 537.200 490.200 538.000 495.800 ;
        RECT 538.900 494.400 539.500 503.600 ;
        RECT 543.700 500.400 544.300 507.600 ;
        RECT 543.600 500.300 544.400 500.400 ;
        RECT 543.600 499.700 545.900 500.300 ;
        RECT 543.600 499.600 544.400 499.700 ;
        RECT 543.600 495.600 544.400 496.400 ;
        RECT 545.300 494.400 545.900 499.700 ;
        RECT 538.800 493.600 539.600 494.400 ;
        RECT 545.200 493.600 546.000 494.400 ;
        RECT 540.400 491.600 541.200 492.400 ;
        RECT 540.500 484.400 541.100 491.600 ;
        RECT 543.600 489.600 544.400 490.400 ;
        RECT 540.400 483.600 541.200 484.400 ;
        RECT 545.300 476.400 545.900 493.600 ;
        RECT 546.900 492.400 547.500 509.700 ;
        RECT 554.800 504.200 555.600 515.800 ;
        RECT 561.200 509.600 562.000 510.400 ;
        RECT 561.300 506.400 561.900 509.600 ;
        RECT 561.200 505.600 562.000 506.400 ;
        RECT 564.400 504.200 565.200 515.800 ;
        RECT 566.000 507.600 566.800 508.400 ;
        RECT 566.100 500.300 566.700 507.600 ;
        RECT 567.600 506.200 568.400 511.800 ;
        RECT 569.200 511.600 570.000 512.400 ;
        RECT 578.800 511.600 579.600 512.400 ;
        RECT 572.400 507.600 573.200 508.400 ;
        RECT 575.600 507.600 576.400 508.400 ;
        RECT 570.800 503.600 571.600 504.400 ;
        RECT 567.600 500.300 568.400 500.400 ;
        RECT 566.100 499.700 568.400 500.300 ;
        RECT 567.600 499.600 568.400 499.700 ;
        RECT 546.800 491.600 547.600 492.400 ;
        RECT 546.800 489.600 547.600 490.400 ;
        RECT 556.400 486.200 557.200 497.800 ;
        RECT 562.800 495.600 563.600 496.400 ;
        RECT 562.900 492.400 563.500 495.600 ;
        RECT 562.800 491.600 563.600 492.400 ;
        RECT 566.000 486.200 566.800 497.800 ;
        RECT 567.700 494.400 568.300 499.600 ;
        RECT 567.600 493.600 568.400 494.400 ;
        RECT 569.200 490.200 570.000 495.800 ;
        RECT 570.900 490.400 571.500 503.600 ;
        RECT 575.700 494.400 576.300 507.600 ;
        RECT 578.900 498.400 579.500 511.600 ;
        RECT 578.800 497.600 579.600 498.400 ;
        RECT 574.000 493.600 574.800 494.400 ;
        RECT 575.600 493.600 576.400 494.400 ;
        RECT 574.100 492.400 574.700 493.600 ;
        RECT 572.400 491.600 573.200 492.400 ;
        RECT 574.000 491.600 574.800 492.400 ;
        RECT 570.800 489.600 571.600 490.400 ;
        RECT 551.600 483.600 552.400 484.400 ;
        RECT 578.800 483.600 579.600 484.400 ;
        RECT 545.200 475.600 546.000 476.400 ;
        RECT 530.900 471.700 533.100 472.300 ;
        RECT 529.300 470.400 529.900 471.600 ;
        RECT 529.200 469.600 530.000 470.400 ;
        RECT 530.800 469.600 531.600 470.400 ;
        RECT 530.800 453.600 531.600 454.400 ;
        RECT 530.900 452.400 531.500 453.600 ;
        RECT 532.500 452.400 533.100 471.700 ;
        RECT 538.800 471.800 539.600 472.600 ;
        RECT 545.400 471.800 546.200 472.600 ;
        RECT 538.800 468.400 539.400 471.800 ;
        RECT 542.800 468.400 543.600 468.600 ;
        RECT 538.800 467.800 543.600 468.400 ;
        RECT 538.800 467.000 539.400 467.800 ;
        RECT 540.200 467.000 541.000 467.200 ;
        RECT 543.600 467.000 544.400 467.200 ;
        RECT 545.600 467.000 546.200 471.800 ;
        RECT 548.400 469.600 549.200 470.400 ;
        RECT 548.500 468.400 549.100 469.600 ;
        RECT 548.400 467.600 549.200 468.400 ;
        RECT 535.600 465.600 536.400 466.400 ;
        RECT 538.800 466.200 539.600 467.000 ;
        RECT 540.200 466.400 544.400 467.000 ;
        RECT 545.400 466.200 546.200 467.000 ;
        RECT 535.700 458.400 536.300 465.600 ;
        RECT 543.600 463.600 544.400 464.400 ;
        RECT 543.700 458.400 544.300 463.600 ;
        RECT 535.600 457.600 536.400 458.400 ;
        RECT 540.400 457.600 541.200 458.400 ;
        RECT 543.600 457.600 544.400 458.400 ;
        RECT 529.200 452.300 530.000 452.400 ;
        RECT 527.700 451.700 530.000 452.300 ;
        RECT 529.200 451.600 530.000 451.700 ;
        RECT 530.800 451.600 531.600 452.400 ;
        RECT 532.400 451.600 533.200 452.400 ;
        RECT 542.000 451.600 542.800 452.400 ;
        RECT 514.900 450.400 515.500 451.600 ;
        RECT 514.800 449.600 515.600 450.400 ;
        RECT 516.400 449.600 517.200 450.400 ;
        RECT 516.500 448.400 517.100 449.600 ;
        RECT 511.600 447.600 512.400 448.400 ;
        RECT 513.200 447.600 514.000 448.400 ;
        RECT 516.400 447.600 517.200 448.400 ;
        RECT 513.300 446.400 513.900 447.600 ;
        RECT 510.000 445.600 510.800 446.400 ;
        RECT 513.200 445.600 514.000 446.400 ;
        RECT 519.700 444.400 520.300 451.600 ;
        RECT 526.000 449.600 526.800 450.400 ;
        RECT 519.600 443.600 520.400 444.400 ;
        RECT 529.200 443.600 530.000 444.400 ;
        RECT 535.600 443.600 536.400 444.400 ;
        RECT 529.300 438.400 529.900 443.600 ;
        RECT 535.700 440.400 536.300 443.600 ;
        RECT 535.600 439.600 536.400 440.400 ;
        RECT 511.600 437.600 512.400 438.400 ;
        RECT 519.600 429.600 520.400 430.400 ;
        RECT 508.400 415.600 509.200 416.400 ;
        RECT 505.200 413.600 506.000 414.400 ;
        RECT 510.000 413.600 510.800 414.400 ;
        RECT 514.800 413.600 515.600 414.400 ;
        RECT 505.300 412.400 505.900 413.600 ;
        RECT 505.200 411.600 506.000 412.400 ;
        RECT 513.200 411.600 514.000 412.400 ;
        RECT 513.300 410.400 513.900 411.600 ;
        RECT 514.900 410.400 515.500 413.600 ;
        RECT 516.400 411.600 517.200 412.400 ;
        RECT 513.200 409.600 514.000 410.400 ;
        RECT 514.800 409.600 515.600 410.400 ;
        RECT 516.400 409.600 517.200 410.400 ;
        RECT 518.000 409.600 518.800 410.400 ;
        RECT 516.500 406.400 517.100 409.600 ;
        RECT 518.100 408.400 518.700 409.600 ;
        RECT 518.000 407.600 518.800 408.400 ;
        RECT 516.400 405.600 517.200 406.400 ;
        RECT 508.400 401.600 509.200 402.400 ;
        RECT 503.600 399.600 504.400 400.400 ;
        RECT 490.800 397.600 491.600 398.400 ;
        RECT 506.800 395.600 507.600 396.400 ;
        RECT 489.200 391.600 490.000 392.400 ;
        RECT 482.800 389.600 483.600 390.400 ;
        RECT 452.400 381.600 453.200 382.400 ;
        RECT 457.200 377.600 458.000 378.400 ;
        RECT 457.300 372.400 457.900 377.600 ;
        RECT 450.800 371.600 451.600 372.400 ;
        RECT 457.200 371.600 458.000 372.400 ;
        RECT 420.400 369.600 421.200 370.400 ;
        RECT 423.600 369.600 424.400 370.400 ;
        RECT 438.000 369.600 438.800 370.400 ;
        RECT 444.400 369.600 445.200 370.400 ;
        RECT 449.200 369.600 450.000 370.400 ;
        RECT 438.100 360.400 438.700 369.600 ;
        RECT 438.000 359.600 438.800 360.400 ;
        RECT 450.900 358.400 451.500 371.600 ;
        RECT 458.800 364.200 459.600 377.800 ;
        RECT 460.400 364.200 461.200 377.800 ;
        RECT 462.000 364.200 462.800 377.800 ;
        RECT 463.600 366.200 464.400 377.800 ;
        RECT 465.200 375.600 466.000 376.400 ;
        RECT 465.300 372.400 465.900 375.600 ;
        RECT 465.200 371.600 466.000 372.400 ;
        RECT 466.800 366.200 467.600 377.800 ;
        RECT 468.400 373.600 469.200 374.400 ;
        RECT 470.000 366.200 470.800 377.800 ;
        RECT 471.600 364.200 472.400 377.800 ;
        RECT 473.200 364.200 474.000 377.800 ;
        RECT 482.900 374.400 483.500 389.600 ;
        RECT 506.900 388.400 507.500 395.600 ;
        RECT 508.500 390.400 509.100 401.600 ;
        RECT 510.000 399.600 510.800 400.400 ;
        RECT 510.100 398.400 510.700 399.600 ;
        RECT 510.000 397.600 510.800 398.400 ;
        RECT 516.400 393.600 517.200 394.400 ;
        RECT 513.200 391.600 514.000 392.400 ;
        RECT 508.400 389.600 509.200 390.400 ;
        RECT 516.500 388.400 517.100 393.600 ;
        RECT 519.700 390.400 520.300 429.600 ;
        RECT 521.200 424.200 522.000 437.800 ;
        RECT 522.800 424.200 523.600 437.800 ;
        RECT 524.400 424.200 525.200 437.800 ;
        RECT 529.200 437.600 530.000 438.400 ;
        RECT 526.000 424.200 526.800 435.800 ;
        RECT 527.600 425.600 528.400 426.400 ;
        RECT 529.200 424.200 530.000 435.800 ;
        RECT 530.800 427.600 531.600 428.400 ;
        RECT 530.900 422.400 531.500 427.600 ;
        RECT 532.400 424.200 533.200 435.800 ;
        RECT 534.000 424.200 534.800 437.800 ;
        RECT 535.600 424.200 536.400 437.800 ;
        RECT 542.100 430.400 542.700 451.600 ;
        RECT 548.500 440.400 549.100 467.600 ;
        RECT 551.700 460.400 552.300 483.600 ;
        RECT 554.800 473.600 555.600 474.400 ;
        RECT 553.200 471.600 554.000 472.400 ;
        RECT 554.900 470.400 555.500 473.600 ;
        RECT 557.800 471.800 558.600 472.600 ;
        RECT 564.400 471.800 565.200 472.600 ;
        RECT 554.800 469.600 555.600 470.400 ;
        RECT 554.900 466.400 555.500 469.600 ;
        RECT 556.400 467.600 557.200 468.400 ;
        RECT 556.500 466.400 557.100 467.600 ;
        RECT 557.800 467.000 558.400 471.800 ;
        RECT 560.400 468.400 561.200 468.600 ;
        RECT 564.600 468.400 565.200 471.800 ;
        RECT 569.000 471.800 569.800 472.600 ;
        RECT 575.600 471.800 576.400 472.600 ;
        RECT 560.400 467.800 565.200 468.400 ;
        RECT 559.600 467.000 560.400 467.200 ;
        RECT 563.000 467.000 563.800 467.200 ;
        RECT 564.600 467.000 565.200 467.800 ;
        RECT 566.000 467.600 566.800 468.400 ;
        RECT 567.600 467.600 568.400 468.400 ;
        RECT 554.800 465.600 555.600 466.400 ;
        RECT 556.400 465.600 557.200 466.400 ;
        RECT 557.800 466.200 558.600 467.000 ;
        RECT 559.600 466.400 563.800 467.000 ;
        RECT 564.400 466.200 565.200 467.000 ;
        RECT 562.800 463.600 563.600 464.400 ;
        RECT 562.900 460.400 563.500 463.600 ;
        RECT 551.600 459.600 552.400 460.400 ;
        RECT 562.800 459.600 563.600 460.400 ;
        RECT 550.000 444.200 550.800 457.800 ;
        RECT 551.600 444.200 552.400 457.800 ;
        RECT 553.200 444.200 554.000 457.800 ;
        RECT 554.800 446.200 555.600 457.800 ;
        RECT 556.400 455.600 557.200 456.400 ;
        RECT 558.000 446.200 558.800 457.800 ;
        RECT 559.600 457.600 560.400 458.400 ;
        RECT 559.700 454.400 560.300 457.600 ;
        RECT 559.600 453.600 560.400 454.400 ;
        RECT 559.600 451.600 560.400 452.400 ;
        RECT 559.600 449.600 560.400 450.400 ;
        RECT 545.200 439.600 546.000 440.400 ;
        RECT 548.400 439.600 549.200 440.400 ;
        RECT 551.600 439.600 552.400 440.400 ;
        RECT 545.300 430.400 545.900 439.600 ;
        RECT 551.700 430.400 552.300 439.600 ;
        RECT 559.700 438.400 560.300 449.600 ;
        RECT 561.200 446.200 562.000 457.800 ;
        RECT 562.800 444.200 563.600 457.800 ;
        RECT 564.400 444.200 565.200 457.800 ;
        RECT 566.100 442.400 566.700 467.600 ;
        RECT 569.000 467.000 569.600 471.800 ;
        RECT 571.600 468.400 572.400 468.600 ;
        RECT 575.800 468.400 576.400 471.800 ;
        RECT 577.200 469.600 578.000 470.400 ;
        RECT 578.800 469.600 579.600 470.400 ;
        RECT 577.300 468.400 577.900 469.600 ;
        RECT 578.900 468.400 579.500 469.600 ;
        RECT 571.600 467.800 576.400 468.400 ;
        RECT 570.800 467.000 571.600 467.200 ;
        RECT 574.200 467.000 575.000 467.200 ;
        RECT 575.800 467.000 576.400 467.800 ;
        RECT 577.200 467.600 578.000 468.400 ;
        RECT 578.800 467.600 579.600 468.400 ;
        RECT 569.000 466.200 569.800 467.000 ;
        RECT 570.800 466.400 575.000 467.000 ;
        RECT 575.600 466.200 576.400 467.000 ;
        RECT 572.400 453.600 573.200 454.400 ;
        RECT 566.000 441.600 566.800 442.400 ;
        RECT 559.600 437.600 560.400 438.400 ;
        RECT 542.000 429.600 542.800 430.400 ;
        RECT 545.200 429.600 546.000 430.400 ;
        RECT 546.800 429.600 547.600 430.400 ;
        RECT 551.600 429.600 552.400 430.400 ;
        RECT 554.800 429.600 555.600 430.400 ;
        RECT 556.400 429.600 557.200 430.400 ;
        RECT 561.200 429.600 562.000 430.400 ;
        RECT 526.000 421.600 526.800 422.400 ;
        RECT 530.800 421.600 531.600 422.400 ;
        RECT 526.100 418.400 526.700 421.600 ;
        RECT 545.300 420.400 545.900 429.600 ;
        RECT 545.200 419.600 546.000 420.400 ;
        RECT 546.900 418.400 547.500 429.600 ;
        RECT 526.000 417.600 526.800 418.400 ;
        RECT 542.000 417.600 542.800 418.400 ;
        RECT 546.800 417.600 547.600 418.400 ;
        RECT 521.200 415.600 522.000 416.400 ;
        RECT 537.400 415.600 538.200 415.800 ;
        RECT 537.400 415.000 543.000 415.600 ;
        RECT 543.600 415.000 544.400 415.800 ;
        RECT 550.000 415.600 550.800 416.400 ;
        RECT 532.400 413.600 533.200 414.400 ;
        RECT 535.600 413.600 536.400 414.400 ;
        RECT 532.500 412.400 533.100 413.600 ;
        RECT 532.400 411.600 533.200 412.400 ;
        RECT 521.200 409.600 522.000 410.400 ;
        RECT 537.400 410.200 538.000 415.000 ;
        RECT 538.800 414.800 539.600 415.000 ;
        RECT 542.200 414.800 543.000 415.000 ;
        RECT 543.800 414.200 544.400 415.000 ;
        RECT 538.800 413.600 544.400 414.200 ;
        RECT 545.200 413.600 546.000 414.400 ;
        RECT 546.800 413.600 547.600 414.400 ;
        RECT 538.800 412.200 539.400 413.600 ;
        RECT 538.600 411.400 539.400 412.200 ;
        RECT 543.800 410.200 544.400 413.600 ;
        RECT 545.300 412.400 545.900 413.600 ;
        RECT 545.200 411.600 546.000 412.400 ;
        RECT 537.400 409.400 538.200 410.200 ;
        RECT 543.600 409.400 544.400 410.200 ;
        RECT 550.100 410.300 550.700 415.600 ;
        RECT 551.700 414.400 552.300 429.600 ;
        RECT 553.200 427.600 554.000 428.400 ;
        RECT 553.200 423.600 554.000 424.400 ;
        RECT 553.300 414.400 553.900 423.600 ;
        RECT 554.900 418.300 555.500 429.600 ;
        RECT 561.300 428.400 561.900 429.600 ;
        RECT 561.200 427.600 562.000 428.400 ;
        RECT 570.800 427.600 571.600 428.400 ;
        RECT 566.000 423.600 566.800 424.400 ;
        RECT 569.200 423.600 570.000 424.400 ;
        RECT 566.000 421.600 566.800 422.400 ;
        RECT 558.000 419.600 558.800 420.400 ;
        RECT 554.900 417.700 557.100 418.300 ;
        RECT 551.600 413.600 552.400 414.400 ;
        RECT 553.200 413.600 554.000 414.400 ;
        RECT 551.600 410.300 552.400 410.400 ;
        RECT 550.100 409.700 552.400 410.300 ;
        RECT 529.200 403.600 530.000 404.400 ;
        RECT 548.400 403.600 549.200 404.400 ;
        RECT 529.300 398.400 529.900 403.600 ;
        RECT 519.600 389.600 520.400 390.400 ;
        RECT 521.200 389.600 522.000 390.400 ;
        RECT 494.000 387.600 494.800 388.400 ;
        RECT 506.800 387.600 507.600 388.400 ;
        RECT 514.800 387.600 515.600 388.400 ;
        RECT 516.400 387.600 517.200 388.400 ;
        RECT 484.400 383.600 485.200 384.400 ;
        RECT 484.500 382.400 485.100 383.600 ;
        RECT 484.400 381.600 485.200 382.400 ;
        RECT 484.500 376.400 485.100 381.600 ;
        RECT 506.900 376.400 507.500 387.600 ;
        RECT 511.600 385.600 512.400 386.400 ;
        RECT 511.700 384.400 512.300 385.600 ;
        RECT 511.600 383.600 512.400 384.400 ;
        RECT 514.800 383.600 515.600 384.400 ;
        RECT 508.400 381.600 509.200 382.400 ;
        RECT 508.500 378.400 509.100 381.600 ;
        RECT 514.900 378.400 515.500 383.600 ;
        RECT 521.300 382.400 521.900 389.600 ;
        RECT 526.000 384.200 526.800 397.800 ;
        RECT 527.600 384.200 528.400 397.800 ;
        RECT 529.200 397.600 530.000 398.400 ;
        RECT 529.200 384.200 530.000 395.800 ;
        RECT 530.800 387.600 531.600 388.400 ;
        RECT 532.400 384.200 533.200 395.800 ;
        RECT 534.000 385.600 534.800 386.400 ;
        RECT 534.100 382.400 534.700 385.600 ;
        RECT 535.600 384.200 536.400 395.800 ;
        RECT 537.200 384.200 538.000 397.800 ;
        RECT 538.800 384.200 539.600 397.800 ;
        RECT 540.400 384.200 541.200 397.800 ;
        RECT 548.500 392.400 549.100 403.600 ;
        RECT 548.400 391.600 549.200 392.400 ;
        RECT 550.100 390.400 550.700 409.700 ;
        RECT 551.600 409.600 552.400 409.700 ;
        RECT 551.600 397.600 552.400 398.400 ;
        RECT 551.700 390.400 552.300 397.600 ;
        RECT 542.000 389.600 542.800 390.400 ;
        RECT 550.000 389.600 551.000 390.400 ;
        RECT 551.600 389.600 552.400 390.400 ;
        RECT 521.200 381.600 522.000 382.400 ;
        RECT 534.000 381.600 534.800 382.400 ;
        RECT 537.200 381.600 538.000 382.400 ;
        RECT 508.400 377.600 509.200 378.400 ;
        RECT 514.800 377.600 515.600 378.400 ;
        RECT 484.400 375.600 485.200 376.400 ;
        RECT 498.800 375.600 499.600 376.400 ;
        RECT 506.800 375.600 507.600 376.400 ;
        RECT 498.900 374.400 499.500 375.600 ;
        RECT 478.000 373.600 478.800 374.400 ;
        RECT 482.800 373.600 483.600 374.400 ;
        RECT 498.800 373.600 499.600 374.400 ;
        RECT 500.400 373.600 501.200 374.400 ;
        RECT 478.100 372.400 478.700 373.600 ;
        RECT 476.400 371.600 477.200 372.400 ;
        RECT 478.000 371.600 478.800 372.400 ;
        RECT 486.000 371.600 486.800 372.400 ;
        RECT 505.200 371.600 506.000 372.400 ;
        RECT 511.600 371.600 512.400 372.400 ;
        RECT 412.400 351.600 413.200 352.400 ;
        RECT 382.000 349.600 382.800 350.400 ;
        RECT 388.400 349.600 389.200 350.400 ;
        RECT 390.000 349.600 390.800 350.400 ;
        RECT 393.200 349.600 394.000 350.400 ;
        RECT 398.000 349.600 398.800 350.400 ;
        RECT 399.600 349.600 400.400 350.400 ;
        RECT 409.200 349.600 410.000 350.400 ;
        RECT 423.600 349.600 424.400 350.400 ;
        RECT 374.000 347.600 374.800 348.400 ;
        RECT 380.400 347.600 381.200 348.400 ;
        RECT 374.100 346.400 374.700 347.600 ;
        RECT 374.000 345.600 374.800 346.400 ;
        RECT 378.800 345.600 379.600 346.400 ;
        RECT 370.800 343.600 371.600 344.400 ;
        RECT 370.900 330.400 371.500 343.600 ;
        RECT 378.900 338.400 379.500 345.600 ;
        RECT 380.400 343.600 381.200 344.400 ;
        RECT 378.800 337.600 379.600 338.400 ;
        RECT 380.500 336.400 381.100 343.600 ;
        RECT 382.000 339.600 382.800 340.400 ;
        RECT 380.400 335.600 381.200 336.400 ;
        RECT 375.600 333.600 376.400 334.400 ;
        RECT 377.200 333.600 378.000 334.400 ;
        RECT 374.000 331.600 374.800 332.400 ;
        RECT 370.800 329.600 371.600 330.400 ;
        RECT 372.400 329.600 373.200 330.400 ;
        RECT 370.800 315.600 371.600 316.400 ;
        RECT 370.900 312.400 371.500 315.600 ;
        RECT 372.500 314.400 373.100 329.600 ;
        RECT 374.000 327.600 374.800 328.400 ;
        RECT 375.700 320.300 376.300 333.600 ;
        RECT 377.300 324.400 377.900 333.600 ;
        RECT 378.800 331.600 379.600 332.400 ;
        RECT 378.900 328.400 379.500 331.600 ;
        RECT 378.800 327.600 379.600 328.400 ;
        RECT 377.200 323.600 378.000 324.400 ;
        RECT 374.100 319.700 376.300 320.300 ;
        RECT 372.400 313.600 373.200 314.400 ;
        RECT 370.800 311.600 371.600 312.400 ;
        RECT 370.800 309.600 371.600 310.400 ;
        RECT 369.200 307.600 370.000 308.400 ;
        RECT 369.300 298.400 369.900 307.600 ;
        RECT 369.200 297.600 370.000 298.400 ;
        RECT 367.600 293.600 368.400 294.400 ;
        RECT 370.900 292.400 371.500 309.600 ;
        RECT 374.100 294.400 374.700 319.700 ;
        RECT 375.600 317.600 376.400 318.400 ;
        RECT 375.700 314.400 376.300 317.600 ;
        RECT 375.600 313.600 376.400 314.400 ;
        RECT 382.100 310.400 382.700 339.600 ;
        RECT 383.600 333.600 384.400 334.400 ;
        RECT 391.600 333.600 392.400 334.400 ;
        RECT 383.700 322.400 384.300 333.600 ;
        RECT 391.700 330.400 392.300 333.600 ;
        RECT 398.100 332.400 398.700 349.600 ;
        RECT 398.000 331.600 398.800 332.400 ;
        RECT 385.200 329.600 386.000 330.400 ;
        RECT 391.600 329.600 392.400 330.400 ;
        RECT 399.700 328.400 400.300 349.600 ;
        RECT 404.400 347.600 405.200 348.400 ;
        RECT 409.200 347.600 410.000 348.400 ;
        RECT 401.200 345.600 402.000 346.400 ;
        RECT 401.300 334.400 401.900 345.600 ;
        RECT 402.800 343.600 403.600 344.400 ;
        RECT 402.900 340.400 403.500 343.600 ;
        RECT 402.800 339.600 403.600 340.400 ;
        RECT 401.200 333.600 402.000 334.400 ;
        RECT 399.600 327.600 400.400 328.400 ;
        RECT 398.000 323.600 398.800 324.400 ;
        RECT 383.600 321.600 384.400 322.400 ;
        RECT 398.100 320.400 398.700 323.600 ;
        RECT 398.000 319.600 398.800 320.400 ;
        RECT 399.600 317.600 400.400 318.400 ;
        RECT 388.400 315.600 389.200 316.400 ;
        RECT 385.200 311.600 386.000 312.400 ;
        RECT 386.800 311.600 387.600 312.400 ;
        RECT 375.600 309.600 376.400 310.400 ;
        RECT 378.800 309.600 379.600 310.400 ;
        RECT 382.000 309.600 382.800 310.400 ;
        RECT 383.600 309.600 384.400 310.400 ;
        RECT 372.400 293.600 373.200 294.400 ;
        RECT 374.000 293.600 374.800 294.400 ;
        RECT 366.000 291.600 366.800 292.400 ;
        RECT 370.800 291.600 371.600 292.400 ;
        RECT 364.400 281.600 365.200 282.400 ;
        RECT 364.400 271.600 365.200 272.400 ;
        RECT 362.900 267.700 365.100 268.300 ;
        RECT 353.300 262.400 353.900 267.600 ;
        RECT 362.800 265.600 363.600 266.400 ;
        RECT 353.200 261.600 354.000 262.400 ;
        RECT 362.900 260.400 363.500 265.600 ;
        RECT 362.800 259.600 363.600 260.400 ;
        RECT 350.100 257.700 352.300 258.300 ;
        RECT 350.000 255.600 350.800 256.400 ;
        RECT 346.800 253.600 347.600 254.400 ;
        RECT 346.800 251.600 347.600 252.400 ;
        RECT 343.600 249.700 345.900 250.300 ;
        RECT 343.600 249.600 344.400 249.700 ;
        RECT 343.700 248.400 344.300 249.600 ;
        RECT 343.600 247.600 344.400 248.400 ;
        RECT 345.200 247.600 346.000 248.400 ;
        RECT 345.300 244.400 345.900 247.600 ;
        RECT 346.800 245.600 347.600 246.400 ;
        RECT 342.000 243.600 342.800 244.400 ;
        RECT 345.200 243.600 346.000 244.400 ;
        RECT 340.400 237.600 341.200 238.400 ;
        RECT 342.100 236.300 342.700 243.600 ;
        RECT 340.500 235.700 342.700 236.300 ;
        RECT 340.500 232.400 341.100 235.700 ;
        RECT 342.000 233.600 342.800 234.400 ;
        RECT 346.900 232.400 347.500 245.600 ;
        RECT 351.700 238.400 352.300 257.700 ;
        RECT 356.400 251.600 357.200 252.400 ;
        RECT 351.600 237.600 352.400 238.400 ;
        RECT 353.200 235.600 354.000 236.400 ;
        RECT 348.400 233.600 349.200 234.400 ;
        RECT 351.600 233.600 352.400 234.400 ;
        RECT 338.800 231.600 339.600 232.400 ;
        RECT 340.400 231.600 341.200 232.400 ;
        RECT 346.800 231.600 347.600 232.400 ;
        RECT 351.600 231.600 352.400 232.400 ;
        RECT 354.800 231.600 355.600 232.400 ;
        RECT 340.400 229.600 341.200 230.400 ;
        RECT 346.800 229.600 347.600 230.400 ;
        RECT 353.200 229.600 354.000 230.400 ;
        RECT 337.200 227.600 338.000 228.400 ;
        RECT 334.000 225.600 334.800 226.400 ;
        RECT 337.300 222.400 337.900 227.600 ;
        RECT 337.200 221.600 338.000 222.400 ;
        RECT 329.200 213.600 330.000 214.400 ;
        RECT 330.800 206.200 331.600 217.800 ;
        RECT 310.000 203.600 310.800 203.700 ;
        RECT 310.000 201.600 310.800 202.400 ;
        RECT 310.100 198.400 310.700 201.600 ;
        RECT 300.400 197.600 301.200 198.400 ;
        RECT 310.000 197.600 310.800 198.400 ;
        RECT 300.400 187.600 301.200 188.400 ;
        RECT 311.700 186.400 312.300 203.700 ;
        RECT 324.400 203.600 325.200 204.400 ;
        RECT 332.400 204.200 333.200 217.800 ;
        RECT 334.000 204.200 334.800 217.800 ;
        RECT 337.300 214.400 337.900 221.600 ;
        RECT 346.900 220.400 347.500 229.600 ;
        RECT 348.400 227.600 349.200 228.400 ;
        RECT 346.800 219.600 347.600 220.400 ;
        RECT 351.600 219.600 352.400 220.400 ;
        RECT 351.700 218.400 352.300 219.600 ;
        RECT 351.600 217.600 352.400 218.400 ;
        RECT 340.400 215.600 341.200 216.400 ;
        RECT 337.200 213.600 338.000 214.400 ;
        RECT 340.500 212.400 341.100 215.600 ;
        RECT 343.600 213.600 344.400 214.400 ;
        RECT 350.000 213.600 350.800 214.400 ;
        RECT 340.400 211.600 341.200 212.400 ;
        RECT 324.500 198.400 325.100 203.600 ;
        RECT 324.400 197.600 325.200 198.400 ;
        RECT 313.200 189.600 314.000 190.400 ;
        RECT 314.800 189.600 315.600 190.400 ;
        RECT 318.000 189.600 318.800 190.400 ;
        RECT 332.400 189.600 333.200 190.400 ;
        RECT 308.400 185.600 309.200 186.400 ;
        RECT 311.600 185.600 312.400 186.400 ;
        RECT 298.800 175.600 299.600 176.400 ;
        RECT 297.200 173.600 298.000 174.400 ;
        RECT 297.300 160.400 297.900 173.600 ;
        RECT 297.200 159.600 298.000 160.400 ;
        RECT 292.400 155.600 293.200 156.400 ;
        RECT 298.900 154.400 299.500 175.600 ;
        RECT 310.000 164.200 310.800 177.800 ;
        RECT 311.600 164.200 312.400 177.800 ;
        RECT 313.200 166.200 314.000 177.800 ;
        RECT 314.900 176.400 315.500 189.600 ;
        RECT 316.400 187.600 317.200 188.400 ;
        RECT 316.500 182.400 317.100 187.600 ;
        RECT 321.200 183.600 322.000 184.400 ;
        RECT 316.400 181.600 317.200 182.400 ;
        RECT 321.300 180.400 321.900 183.600 ;
        RECT 321.200 179.600 322.000 180.400 ;
        RECT 314.800 175.600 315.600 176.400 ;
        RECT 314.800 173.600 315.600 174.400 ;
        RECT 316.400 166.200 317.200 177.800 ;
        RECT 318.000 175.600 318.800 176.400 ;
        RECT 318.000 165.600 318.800 166.400 ;
        RECT 319.600 166.200 320.400 177.800 ;
        RECT 298.800 153.600 299.600 154.400 ;
        RECT 318.100 152.400 318.700 165.600 ;
        RECT 321.200 164.200 322.000 177.800 ;
        RECT 322.800 164.200 323.600 177.800 ;
        RECT 324.400 164.200 325.200 177.800 ;
        RECT 332.500 172.400 333.100 189.600 ;
        RECT 334.000 184.200 334.800 197.800 ;
        RECT 335.600 184.200 336.400 197.800 ;
        RECT 337.200 184.200 338.000 197.800 ;
        RECT 338.800 184.200 339.600 195.800 ;
        RECT 340.400 195.600 341.200 196.400 ;
        RECT 340.500 186.400 341.100 195.600 ;
        RECT 340.400 185.600 341.200 186.400 ;
        RECT 340.400 183.600 341.200 184.400 ;
        RECT 342.000 184.200 342.800 195.800 ;
        RECT 343.700 194.400 344.300 213.600 ;
        RECT 345.200 211.600 346.000 212.400 ;
        RECT 345.300 204.400 345.900 211.600 ;
        RECT 345.200 203.600 346.000 204.400 ;
        RECT 343.600 193.600 344.400 194.400 ;
        RECT 343.600 187.600 344.400 188.400 ;
        RECT 343.700 184.400 344.300 187.600 ;
        RECT 343.600 183.600 344.400 184.400 ;
        RECT 345.200 184.200 346.000 195.800 ;
        RECT 346.800 184.200 347.600 197.800 ;
        RECT 348.400 184.200 349.200 197.800 ;
        RECT 353.300 194.400 353.900 229.600 ;
        RECT 354.900 226.400 355.500 231.600 ;
        RECT 356.500 228.400 357.100 251.600 ;
        RECT 359.600 244.200 360.400 257.800 ;
        RECT 361.200 244.200 362.000 257.800 ;
        RECT 362.800 246.200 363.600 257.800 ;
        RECT 364.500 254.400 365.100 267.700 ;
        RECT 366.100 266.300 366.700 291.600 ;
        RECT 369.200 289.600 370.000 290.400 ;
        RECT 369.300 284.400 369.900 289.600 ;
        RECT 372.500 288.400 373.100 293.600 ;
        RECT 374.100 290.400 374.700 293.600 ;
        RECT 374.000 289.600 374.800 290.400 ;
        RECT 372.400 287.600 373.200 288.400 ;
        RECT 375.700 286.300 376.300 309.600 ;
        RECT 377.200 307.600 378.000 308.400 ;
        RECT 380.400 307.600 381.200 308.400 ;
        RECT 377.200 297.600 378.000 298.400 ;
        RECT 377.300 288.400 377.900 297.600 ;
        RECT 380.400 293.600 381.200 294.400 ;
        RECT 382.100 288.400 382.700 309.600 ;
        RECT 383.700 308.400 384.300 309.600 ;
        RECT 383.600 307.600 384.400 308.400 ;
        RECT 386.900 298.400 387.500 311.600 ;
        RECT 388.500 310.400 389.100 315.600 ;
        RECT 396.400 311.600 397.200 312.400 ;
        RECT 388.400 309.600 389.200 310.400 ;
        RECT 391.600 309.600 392.400 310.400 ;
        RECT 394.800 309.600 395.600 310.400 ;
        RECT 388.500 298.400 389.100 309.600 ;
        RECT 390.000 307.600 390.800 308.400 ;
        RECT 390.100 302.400 390.700 307.600 ;
        RECT 390.000 301.600 390.800 302.400 ;
        RECT 386.800 297.600 387.600 298.400 ;
        RECT 388.400 297.600 389.200 298.400 ;
        RECT 386.800 293.600 387.600 294.400 ;
        RECT 390.000 293.600 390.800 294.400 ;
        RECT 385.200 291.600 386.000 292.400 ;
        RECT 377.200 287.600 378.000 288.400 ;
        RECT 380.400 287.600 381.200 288.400 ;
        RECT 382.000 287.600 382.800 288.400 ;
        RECT 375.700 285.700 377.900 286.300 ;
        RECT 369.200 283.600 370.000 284.400 ;
        RECT 372.400 275.600 373.200 276.400 ;
        RECT 372.500 274.400 373.100 275.600 ;
        RECT 372.400 273.600 373.200 274.400 ;
        RECT 377.300 272.400 377.900 285.700 ;
        RECT 378.800 281.600 379.600 282.400 ;
        RECT 378.900 274.400 379.500 281.600 ;
        RECT 380.500 278.400 381.100 287.600 ;
        RECT 385.300 286.400 385.900 291.600 ;
        RECT 385.200 285.600 386.000 286.400 ;
        RECT 382.000 283.600 382.800 284.400 ;
        RECT 383.600 283.600 384.400 284.400 ;
        RECT 380.400 277.600 381.200 278.400 ;
        RECT 382.100 274.400 382.700 283.600 ;
        RECT 383.700 278.400 384.300 283.600 ;
        RECT 385.200 281.600 386.000 282.400 ;
        RECT 383.600 277.600 384.400 278.400 ;
        RECT 385.300 274.400 385.900 281.600 ;
        RECT 378.800 273.600 379.600 274.400 ;
        RECT 382.000 273.600 382.800 274.400 ;
        RECT 385.200 273.600 386.000 274.400 ;
        RECT 369.200 271.600 370.000 272.400 ;
        RECT 375.600 271.600 376.400 272.400 ;
        RECT 377.200 271.600 378.000 272.400 ;
        RECT 382.000 271.600 382.800 272.400 ;
        RECT 375.700 270.400 376.300 271.600 ;
        RECT 377.300 270.400 377.900 271.600 ;
        RECT 382.100 270.400 382.700 271.600 ;
        RECT 367.600 269.600 368.400 270.400 ;
        RECT 372.400 269.600 373.200 270.400 ;
        RECT 375.600 269.600 376.400 270.400 ;
        RECT 377.200 269.600 378.000 270.400 ;
        RECT 382.000 269.600 382.800 270.400 ;
        RECT 383.600 269.600 384.400 270.400 ;
        RECT 367.700 268.400 368.300 269.600 ;
        RECT 372.500 268.400 373.100 269.600 ;
        RECT 367.600 267.600 368.400 268.400 ;
        RECT 372.400 267.600 373.200 268.400 ;
        RECT 366.100 265.700 368.300 266.300 ;
        RECT 366.000 263.600 366.800 264.400 ;
        RECT 366.100 262.400 366.700 263.600 ;
        RECT 367.700 262.400 368.300 265.700 ;
        RECT 366.000 261.600 366.800 262.400 ;
        RECT 367.600 261.600 368.400 262.400 ;
        RECT 367.600 259.600 368.400 260.400 ;
        RECT 364.400 253.600 365.200 254.400 ;
        RECT 366.000 246.200 366.800 257.800 ;
        RECT 367.700 256.400 368.300 259.600 ;
        RECT 367.600 255.600 368.400 256.400 ;
        RECT 369.200 246.200 370.000 257.800 ;
        RECT 370.800 244.200 371.600 257.800 ;
        RECT 372.400 244.200 373.200 257.800 ;
        RECT 374.000 244.200 374.800 257.800 ;
        RECT 375.700 256.400 376.300 269.600 ;
        RECT 377.300 264.400 377.900 269.600 ;
        RECT 386.900 266.400 387.500 293.600 ;
        RECT 390.100 286.400 390.700 293.600 ;
        RECT 391.700 292.400 392.300 309.600 ;
        RECT 393.200 307.600 394.000 308.400 ;
        RECT 394.900 306.400 395.500 309.600 ;
        RECT 396.500 308.400 397.100 311.600 ;
        RECT 398.000 309.600 398.800 310.400 ;
        RECT 398.100 308.400 398.700 309.600 ;
        RECT 396.400 307.600 397.200 308.400 ;
        RECT 398.000 307.600 398.800 308.400 ;
        RECT 394.800 305.600 395.600 306.400 ;
        RECT 396.400 305.600 397.200 306.400 ;
        RECT 393.200 303.600 394.000 304.400 ;
        RECT 393.300 294.400 393.900 303.600 ;
        RECT 396.500 298.400 397.100 305.600 ;
        RECT 399.700 298.400 400.300 317.600 ;
        RECT 401.300 312.400 401.900 333.600 ;
        RECT 404.500 318.400 405.100 347.600 ;
        RECT 407.600 345.600 408.400 346.400 ;
        RECT 415.600 345.600 416.400 346.400 ;
        RECT 410.800 343.600 411.600 344.400 ;
        RECT 410.900 342.400 411.500 343.600 ;
        RECT 410.800 341.600 411.600 342.400 ;
        RECT 414.000 341.600 414.800 342.400 ;
        RECT 414.100 338.400 414.700 341.600 ;
        RECT 406.000 331.600 406.800 332.400 ;
        RECT 404.400 317.600 405.200 318.400 ;
        RECT 402.800 315.600 403.600 316.400 ;
        RECT 401.200 311.600 402.000 312.400 ;
        RECT 402.900 310.400 403.500 315.600 ;
        RECT 402.800 309.600 403.600 310.400 ;
        RECT 404.400 309.600 405.200 310.400 ;
        RECT 404.500 308.400 405.100 309.600 ;
        RECT 402.800 307.600 403.600 308.400 ;
        RECT 404.400 307.600 405.200 308.400 ;
        RECT 402.900 306.400 403.500 307.600 ;
        RECT 402.800 305.600 403.600 306.400 ;
        RECT 396.400 297.600 397.200 298.400 ;
        RECT 399.600 297.600 400.400 298.400 ;
        RECT 401.200 297.600 402.000 298.400 ;
        RECT 399.700 296.400 400.300 297.600 ;
        RECT 399.600 295.600 400.400 296.400 ;
        RECT 393.200 293.600 394.000 294.400 ;
        RECT 391.600 291.600 392.400 292.400 ;
        RECT 390.000 285.600 390.800 286.400 ;
        RECT 390.000 277.600 390.800 278.400 ;
        RECT 391.700 276.300 392.300 291.600 ;
        RECT 398.000 289.600 398.800 290.400 ;
        RECT 396.400 285.600 397.200 286.400 ;
        RECT 390.100 275.700 392.300 276.300 ;
        RECT 390.100 270.400 390.700 275.700 ;
        RECT 391.600 274.300 392.400 274.400 ;
        RECT 391.600 273.700 393.900 274.300 ;
        RECT 391.600 273.600 392.400 273.700 ;
        RECT 390.000 269.600 390.800 270.400 ;
        RECT 386.800 265.600 387.600 266.400 ;
        RECT 377.200 263.600 378.000 264.400 ;
        RECT 386.800 261.600 387.600 262.400 ;
        RECT 386.900 258.400 387.500 261.600 ;
        RECT 386.800 257.600 387.600 258.400 ;
        RECT 390.000 257.600 390.800 258.400 ;
        RECT 391.600 257.600 392.400 258.400 ;
        RECT 375.600 255.600 376.400 256.400 ;
        RECT 388.400 255.600 389.200 256.400 ;
        RECT 383.600 243.600 384.400 244.400 ;
        RECT 383.700 240.400 384.300 243.600 ;
        RECT 388.500 240.400 389.100 255.600 ;
        RECT 390.100 250.300 390.700 257.600 ;
        RECT 391.700 252.400 392.300 257.600 ;
        RECT 391.600 251.600 392.400 252.400 ;
        RECT 390.100 249.700 392.300 250.300 ;
        RECT 391.700 246.400 392.300 249.700 ;
        RECT 393.300 248.400 393.900 273.700 ;
        RECT 394.800 269.600 395.600 270.400 ;
        RECT 394.900 252.300 395.500 269.600 ;
        RECT 396.500 268.400 397.100 285.600 ;
        RECT 396.400 267.600 397.200 268.400 ;
        RECT 398.100 258.400 398.700 289.600 ;
        RECT 399.600 283.600 400.400 284.400 ;
        RECT 399.600 275.600 400.400 276.400 ;
        RECT 401.300 270.400 401.900 297.600 ;
        RECT 402.800 291.600 403.600 292.400 ;
        RECT 401.200 270.300 402.000 270.400 ;
        RECT 399.700 269.700 402.000 270.300 ;
        RECT 398.000 257.600 398.800 258.400 ;
        RECT 398.000 255.600 398.800 256.400 ;
        RECT 398.100 254.400 398.700 255.600 ;
        RECT 398.000 253.600 398.800 254.400 ;
        RECT 399.700 252.400 400.300 269.700 ;
        RECT 401.200 269.600 402.000 269.700 ;
        RECT 401.200 267.600 402.000 268.400 ;
        RECT 401.300 266.400 401.900 267.600 ;
        RECT 401.200 265.600 402.000 266.400 ;
        RECT 402.900 260.400 403.500 291.600 ;
        RECT 406.100 286.400 406.700 331.600 ;
        RECT 407.600 324.200 408.400 337.800 ;
        RECT 409.200 324.200 410.000 337.800 ;
        RECT 410.800 324.200 411.600 337.800 ;
        RECT 412.400 326.200 413.200 337.800 ;
        RECT 414.000 337.600 414.800 338.400 ;
        RECT 414.100 336.400 414.700 337.600 ;
        RECT 414.000 335.600 414.800 336.400 ;
        RECT 407.600 311.600 408.400 312.400 ;
        RECT 412.400 311.600 413.200 312.400 ;
        RECT 407.600 309.600 408.400 310.400 ;
        RECT 409.200 307.600 410.000 308.400 ;
        RECT 410.800 307.600 411.600 308.400 ;
        RECT 410.900 306.400 411.500 307.600 ;
        RECT 414.100 306.400 414.700 335.600 ;
        RECT 415.600 326.200 416.400 337.800 ;
        RECT 417.200 333.600 418.000 334.400 ;
        RECT 417.300 332.400 417.900 333.600 ;
        RECT 417.200 331.600 418.000 332.400 ;
        RECT 418.800 326.200 419.600 337.800 ;
        RECT 420.400 324.200 421.200 337.800 ;
        RECT 422.000 324.200 422.800 337.800 ;
        RECT 423.700 332.400 424.300 349.600 ;
        RECT 425.200 344.200 426.000 357.800 ;
        RECT 426.800 344.200 427.600 357.800 ;
        RECT 428.400 344.200 429.200 357.800 ;
        RECT 430.000 344.200 430.800 355.800 ;
        RECT 431.600 345.600 432.400 346.400 ;
        RECT 431.700 342.400 432.300 345.600 ;
        RECT 433.200 344.200 434.000 355.800 ;
        RECT 434.800 351.600 435.600 352.400 ;
        RECT 434.900 348.400 435.500 351.600 ;
        RECT 434.800 347.600 435.600 348.400 ;
        RECT 431.600 341.600 432.400 342.400 ;
        RECT 434.900 338.400 435.500 347.600 ;
        RECT 436.400 344.200 437.200 355.800 ;
        RECT 438.000 344.200 438.800 357.800 ;
        RECT 439.600 344.200 440.400 357.800 ;
        RECT 450.800 357.600 451.600 358.400 ;
        RECT 446.000 351.600 446.800 352.400 ;
        RECT 442.800 349.600 443.600 350.400 ;
        RECT 431.600 337.600 432.400 338.400 ;
        RECT 434.800 337.600 435.600 338.400 ;
        RECT 423.600 331.600 424.400 332.400 ;
        RECT 431.700 330.400 432.300 337.600 ;
        RECT 436.400 335.600 437.200 336.400 ;
        RECT 434.800 333.600 435.600 334.400 ;
        RECT 431.600 329.600 432.400 330.400 ;
        RECT 434.900 328.400 435.500 333.600 ;
        RECT 436.500 330.400 437.100 335.600 ;
        RECT 439.600 333.600 440.400 334.400 ;
        RECT 436.400 329.600 437.200 330.400 ;
        RECT 441.200 329.600 442.000 330.400 ;
        RECT 434.800 327.600 435.600 328.400 ;
        RECT 433.200 323.600 434.000 324.400 ;
        RECT 433.300 320.400 433.900 323.600 ;
        RECT 423.600 319.600 424.400 320.400 ;
        RECT 433.200 319.600 434.000 320.400 ;
        RECT 418.800 315.600 419.600 316.400 ;
        RECT 415.600 309.600 416.400 310.400 ;
        RECT 417.200 309.600 418.000 310.400 ;
        RECT 410.800 305.600 411.600 306.400 ;
        RECT 414.000 305.600 414.800 306.400 ;
        RECT 412.400 303.600 413.200 304.400 ;
        RECT 412.500 302.400 413.100 303.600 ;
        RECT 412.400 301.600 413.200 302.400 ;
        RECT 415.700 300.400 416.300 309.600 ;
        RECT 417.300 308.400 417.900 309.600 ;
        RECT 418.900 308.400 419.500 315.600 ;
        RECT 423.700 312.400 424.300 319.600 ;
        RECT 436.500 318.400 437.100 329.600 ;
        RECT 442.900 324.400 443.500 349.600 ;
        RECT 446.100 334.400 446.700 351.600 ;
        RECT 460.200 347.600 461.200 348.400 ;
        RECT 449.200 345.600 450.000 346.400 ;
        RECT 449.300 344.400 449.900 345.600 ;
        RECT 449.200 343.600 450.000 344.400 ;
        RECT 470.000 344.200 470.800 357.800 ;
        RECT 471.600 344.200 472.400 357.800 ;
        RECT 473.200 344.200 474.000 357.800 ;
        RECT 474.800 344.200 475.600 355.800 ;
        RECT 476.500 346.400 477.100 371.600 ;
        RECT 505.300 366.400 505.900 371.600 ;
        RECT 511.700 366.400 512.300 371.600 ;
        RECT 505.200 365.600 506.000 366.400 ;
        RECT 511.600 365.600 512.400 366.400 ;
        RECT 482.800 363.600 483.600 364.400 ;
        RECT 521.200 363.600 522.000 364.400 ;
        RECT 530.800 364.200 531.600 377.800 ;
        RECT 532.400 364.200 533.200 377.800 ;
        RECT 534.000 364.200 534.800 377.800 ;
        RECT 535.600 366.200 536.400 377.800 ;
        RECT 537.300 376.400 537.900 381.600 ;
        RECT 542.100 380.400 542.700 389.600 ;
        RECT 553.300 384.400 553.900 413.600 ;
        RECT 554.800 411.600 555.600 412.400 ;
        RECT 554.900 402.400 555.500 411.600 ;
        RECT 556.500 408.400 557.100 417.700 ;
        RECT 558.100 410.400 558.700 419.600 ;
        RECT 566.100 418.400 566.700 421.600 ;
        RECT 566.000 417.600 566.800 418.400 ;
        RECT 561.400 415.600 562.200 415.800 ;
        RECT 561.400 415.000 567.000 415.600 ;
        RECT 567.600 415.000 568.400 415.800 ;
        RECT 558.000 409.600 558.800 410.400 ;
        RECT 561.400 410.200 562.000 415.000 ;
        RECT 562.800 414.800 563.600 415.000 ;
        RECT 566.200 414.800 567.000 415.000 ;
        RECT 567.800 414.200 568.400 415.000 ;
        RECT 569.300 414.400 569.900 423.600 ;
        RECT 570.900 414.400 571.500 427.600 ;
        RECT 562.800 413.600 568.400 414.200 ;
        RECT 569.200 413.600 570.000 414.400 ;
        RECT 570.800 413.600 571.600 414.400 ;
        RECT 562.800 412.200 563.400 413.600 ;
        RECT 562.600 411.400 563.400 412.200 ;
        RECT 567.800 410.200 568.400 413.600 ;
        RECT 569.300 412.400 569.900 413.600 ;
        RECT 569.200 411.600 570.000 412.400 ;
        RECT 572.500 412.300 573.100 453.600 ;
        RECT 575.600 443.600 576.400 444.400 ;
        RECT 575.700 440.400 576.300 443.600 ;
        RECT 580.500 442.400 581.100 531.600 ;
        RECT 580.400 441.600 581.200 442.400 ;
        RECT 575.600 439.600 576.400 440.400 ;
        RECT 574.000 429.600 574.800 430.400 ;
        RECT 574.100 416.300 574.700 429.600 ;
        RECT 575.600 424.200 576.400 437.800 ;
        RECT 577.200 424.200 578.000 437.800 ;
        RECT 578.800 424.200 579.600 437.800 ;
        RECT 580.400 424.200 581.200 435.800 ;
        RECT 582.100 428.400 582.700 531.600 ;
        RECT 583.600 527.600 584.400 528.400 ;
        RECT 583.700 526.400 584.300 527.600 ;
        RECT 583.600 525.600 584.400 526.400 ;
        RECT 588.500 524.400 589.100 549.600 ;
        RECT 583.600 523.600 584.400 524.400 ;
        RECT 588.400 523.600 589.200 524.400 ;
        RECT 583.700 510.400 584.300 523.600 ;
        RECT 583.600 509.600 584.400 510.400 ;
        RECT 585.200 504.200 586.000 517.800 ;
        RECT 586.800 504.200 587.600 517.800 ;
        RECT 588.400 504.200 589.200 517.800 ;
        RECT 590.000 504.200 590.800 515.800 ;
        RECT 591.700 506.400 592.300 555.600 ;
        RECT 593.200 547.600 594.000 548.400 ;
        RECT 596.400 547.600 597.200 548.400 ;
        RECT 594.800 545.600 595.600 546.400 ;
        RECT 594.900 540.400 595.500 545.600 ;
        RECT 594.800 539.600 595.600 540.400 ;
        RECT 596.500 534.300 597.100 547.600 ;
        RECT 602.800 539.600 603.600 540.400 ;
        RECT 598.000 534.300 598.800 534.400 ;
        RECT 596.500 533.700 598.800 534.300 ;
        RECT 598.000 533.600 598.800 533.700 ;
        RECT 602.900 532.400 603.500 539.600 ;
        RECT 612.400 533.600 613.200 534.400 ;
        RECT 598.000 531.600 598.800 532.400 ;
        RECT 602.800 531.600 603.600 532.400 ;
        RECT 598.100 520.400 598.700 531.600 ;
        RECT 599.600 529.600 600.400 530.400 ;
        RECT 594.800 519.600 595.600 520.400 ;
        RECT 598.000 519.600 598.800 520.400 ;
        RECT 591.600 505.600 592.400 506.400 ;
        RECT 591.700 500.400 592.300 505.600 ;
        RECT 593.200 504.200 594.000 515.800 ;
        RECT 594.900 508.400 595.500 519.600 ;
        RECT 594.800 507.600 595.600 508.400 ;
        RECT 596.400 504.200 597.200 515.800 ;
        RECT 598.000 504.200 598.800 517.800 ;
        RECT 599.600 504.200 600.400 517.800 ;
        RECT 604.400 510.300 605.200 510.400 ;
        RECT 604.400 509.700 606.700 510.300 ;
        RECT 604.400 509.600 605.200 509.700 ;
        RECT 591.600 499.600 592.400 500.400 ;
        RECT 594.800 499.600 595.600 500.400 ;
        RECT 588.400 484.200 589.200 497.800 ;
        RECT 590.000 484.200 590.800 497.800 ;
        RECT 591.600 484.200 592.400 497.800 ;
        RECT 593.200 486.200 594.000 497.800 ;
        RECT 594.900 496.400 595.500 499.600 ;
        RECT 594.800 495.600 595.600 496.400 ;
        RECT 594.900 478.300 595.500 495.600 ;
        RECT 596.400 486.200 597.200 497.800 ;
        RECT 598.000 493.600 598.800 494.400 ;
        RECT 598.100 492.400 598.700 493.600 ;
        RECT 598.000 491.600 598.800 492.400 ;
        RECT 599.600 486.200 600.400 497.800 ;
        RECT 601.200 484.200 602.000 497.800 ;
        RECT 602.800 484.200 603.600 497.800 ;
        RECT 606.100 492.400 606.700 509.700 ;
        RECT 606.000 491.600 606.800 492.400 ;
        RECT 588.400 469.600 589.200 470.400 ;
        RECT 588.500 466.400 589.100 469.600 ;
        RECT 583.600 465.600 584.400 466.400 ;
        RECT 588.400 465.600 589.200 466.400 ;
        RECT 583.700 452.400 584.300 465.600 ;
        RECT 590.000 464.200 590.800 477.800 ;
        RECT 591.600 464.200 592.400 477.800 ;
        RECT 593.200 464.200 594.000 477.800 ;
        RECT 594.900 477.700 597.100 478.300 ;
        RECT 594.800 464.200 595.600 475.800 ;
        RECT 596.500 466.400 597.100 477.700 ;
        RECT 596.400 465.600 597.200 466.400 ;
        RECT 596.500 460.400 597.100 465.600 ;
        RECT 598.000 464.200 598.800 475.800 ;
        RECT 599.600 467.600 600.400 468.400 ;
        RECT 601.200 464.200 602.000 475.800 ;
        RECT 602.800 464.200 603.600 477.800 ;
        RECT 604.400 464.200 605.200 477.800 ;
        RECT 591.600 459.600 592.400 460.400 ;
        RECT 596.400 459.600 597.200 460.400 ;
        RECT 583.600 451.600 584.400 452.400 ;
        RECT 583.700 442.300 584.300 451.600 ;
        RECT 585.200 444.200 586.000 457.800 ;
        RECT 586.800 444.200 587.600 457.800 ;
        RECT 588.400 444.200 589.200 457.800 ;
        RECT 590.000 446.200 590.800 457.800 ;
        RECT 591.700 456.400 592.300 459.600 ;
        RECT 591.600 455.600 592.400 456.400 ;
        RECT 593.200 446.200 594.000 457.800 ;
        RECT 594.800 453.600 595.600 454.400 ;
        RECT 594.900 450.400 595.500 453.600 ;
        RECT 594.800 449.600 595.600 450.400 ;
        RECT 596.400 446.200 597.200 457.800 ;
        RECT 598.000 444.200 598.800 457.800 ;
        RECT 599.600 444.200 600.400 457.800 ;
        RECT 606.100 442.400 606.700 491.600 ;
        RECT 583.700 441.700 585.900 442.300 ;
        RECT 582.000 427.600 582.800 428.400 ;
        RECT 582.000 425.600 582.800 426.400 ;
        RECT 582.100 416.400 582.700 425.600 ;
        RECT 583.600 424.200 584.400 435.800 ;
        RECT 585.300 430.400 585.900 441.700 ;
        RECT 599.600 441.600 600.400 442.400 ;
        RECT 606.000 441.600 606.800 442.400 ;
        RECT 585.200 429.600 586.000 430.400 ;
        RECT 585.200 427.600 586.000 428.400 ;
        RECT 585.300 422.400 585.900 427.600 ;
        RECT 586.800 424.200 587.600 435.800 ;
        RECT 588.400 424.200 589.200 437.800 ;
        RECT 590.000 424.200 590.800 437.800 ;
        RECT 585.200 421.600 586.000 422.400 ;
        RECT 574.100 415.700 576.300 416.300 ;
        RECT 572.500 411.700 574.700 412.300 ;
        RECT 574.100 410.400 574.700 411.700 ;
        RECT 561.400 409.400 562.200 410.200 ;
        RECT 567.600 409.400 568.400 410.200 ;
        RECT 574.000 409.600 574.800 410.400 ;
        RECT 556.400 407.600 557.200 408.400 ;
        RECT 567.600 407.600 568.400 408.400 ;
        RECT 554.800 401.600 555.600 402.400 ;
        RECT 554.900 388.400 555.500 401.600 ;
        RECT 558.000 399.600 558.800 400.400 ;
        RECT 558.100 392.400 558.700 399.600 ;
        RECT 567.700 398.400 568.300 407.600 ;
        RECT 572.400 403.600 573.200 404.400 ;
        RECT 567.600 397.600 568.400 398.400 ;
        RECT 561.200 393.600 562.000 394.400 ;
        RECT 558.000 391.600 558.800 392.400 ;
        RECT 566.000 391.600 566.800 392.400 ;
        RECT 556.400 389.600 557.200 390.400 ;
        RECT 558.000 389.600 558.800 390.400 ;
        RECT 561.200 389.600 562.000 390.400 ;
        RECT 554.800 387.600 555.600 388.400 ;
        RECT 556.500 386.400 557.100 389.600 ;
        RECT 559.600 387.600 560.400 388.400 ;
        RECT 556.400 385.600 557.200 386.400 ;
        RECT 553.200 383.600 554.000 384.400 ;
        RECT 554.800 383.600 555.600 384.400 ;
        RECT 542.000 379.600 542.800 380.400 ;
        RECT 546.800 379.600 547.600 380.400 ;
        RECT 537.200 375.600 538.000 376.400 ;
        RECT 482.900 360.400 483.500 363.600 ;
        RECT 479.600 359.600 480.400 360.400 ;
        RECT 482.800 359.600 483.600 360.400 ;
        RECT 476.400 345.600 477.200 346.400 ;
        RECT 478.000 344.200 478.800 355.800 ;
        RECT 479.700 348.400 480.300 359.600 ;
        RECT 479.600 347.600 480.400 348.400 ;
        RECT 481.200 344.200 482.000 355.800 ;
        RECT 482.800 344.200 483.600 357.800 ;
        RECT 484.400 344.200 485.200 357.800 ;
        RECT 489.200 349.600 490.000 350.400 ;
        RECT 495.600 349.600 496.400 350.400 ;
        RECT 502.000 344.200 502.800 357.800 ;
        RECT 503.600 344.200 504.400 357.800 ;
        RECT 505.200 344.200 506.000 355.800 ;
        RECT 506.800 347.600 507.600 348.400 ;
        RECT 508.400 344.200 509.200 355.800 ;
        RECT 510.000 345.600 510.800 346.400 ;
        RECT 511.600 344.200 512.400 355.800 ;
        RECT 513.200 344.200 514.000 357.800 ;
        RECT 514.800 344.200 515.600 357.800 ;
        RECT 516.400 344.200 517.200 357.800 ;
        RECT 521.300 352.400 521.900 363.600 ;
        RECT 532.400 359.600 533.200 360.400 ;
        RECT 532.500 354.400 533.100 359.600 ;
        RECT 532.400 353.600 533.200 354.400 ;
        RECT 534.000 353.600 534.800 354.400 ;
        RECT 532.500 352.400 533.100 353.600 ;
        RECT 521.200 351.600 522.000 352.400 ;
        RECT 532.400 351.600 533.200 352.400 ;
        RECT 518.000 349.600 518.800 350.400 ;
        RECT 529.200 347.600 530.000 348.400 ;
        RECT 529.300 346.400 529.900 347.600 ;
        RECT 522.800 345.600 523.600 346.400 ;
        RECT 529.200 345.600 530.000 346.400 ;
        RECT 452.400 339.600 453.200 340.400 ;
        RECT 462.000 339.600 462.800 340.400 ;
        RECT 452.500 334.400 453.100 339.600 ;
        RECT 455.600 335.600 456.400 336.400 ;
        RECT 455.700 334.400 456.300 335.600 ;
        RECT 446.000 333.600 446.800 334.400 ;
        RECT 450.800 333.600 451.600 334.400 ;
        RECT 452.400 333.600 453.200 334.400 ;
        RECT 455.600 333.600 456.400 334.400 ;
        RECT 447.600 331.600 448.400 332.400 ;
        RECT 447.700 330.400 448.300 331.600 ;
        RECT 455.700 330.400 456.300 333.600 ;
        RECT 462.100 332.400 462.700 339.600 ;
        RECT 466.800 335.600 467.600 336.400 ;
        RECT 468.400 335.600 469.200 336.400 ;
        RECT 490.800 335.600 491.600 336.400 ;
        RECT 505.200 335.600 506.000 336.400 ;
        RECT 468.500 334.400 469.100 335.600 ;
        RECT 465.200 333.600 466.000 334.400 ;
        RECT 468.400 333.600 469.200 334.400 ;
        RECT 482.800 333.600 483.600 334.400 ;
        RECT 484.400 333.600 485.200 334.400 ;
        RECT 489.200 333.600 490.000 334.400 ;
        RECT 460.400 331.600 461.200 332.400 ;
        RECT 462.000 331.600 462.800 332.400 ;
        RECT 444.400 329.600 445.200 330.400 ;
        RECT 447.600 329.600 448.400 330.400 ;
        RECT 450.800 329.600 451.600 330.400 ;
        RECT 455.600 329.600 456.400 330.400 ;
        RECT 442.800 323.600 443.600 324.400 ;
        RECT 444.500 320.400 445.100 329.600 ;
        RECT 454.000 327.600 454.800 328.400 ;
        RECT 449.200 323.600 450.000 324.400 ;
        RECT 444.400 319.600 445.200 320.400 ;
        RECT 423.600 311.600 424.400 312.400 ;
        RECT 420.400 309.600 421.200 310.400 ;
        RECT 423.600 309.600 424.400 310.400 ;
        RECT 428.400 309.600 429.200 310.400 ;
        RECT 417.200 307.600 418.000 308.400 ;
        RECT 418.800 307.600 419.600 308.400 ;
        RECT 420.500 302.400 421.100 309.600 ;
        RECT 418.800 301.600 419.600 302.400 ;
        RECT 420.400 301.600 421.200 302.400 ;
        RECT 415.600 299.600 416.400 300.400 ;
        RECT 406.000 285.600 406.800 286.400 ;
        RECT 409.200 284.200 410.000 297.800 ;
        RECT 410.800 284.200 411.600 297.800 ;
        RECT 412.400 284.200 413.200 297.800 ;
        RECT 414.000 286.200 414.800 297.800 ;
        RECT 415.600 295.600 416.400 296.400 ;
        RECT 417.200 286.200 418.000 297.800 ;
        RECT 418.900 294.400 419.500 301.600 ;
        RECT 418.800 293.600 419.600 294.400 ;
        RECT 420.400 286.200 421.200 297.800 ;
        RECT 422.000 284.200 422.800 297.800 ;
        RECT 423.600 284.200 424.400 297.800 ;
        RECT 428.500 292.400 429.100 309.600 ;
        RECT 433.200 304.200 434.000 317.800 ;
        RECT 434.800 304.200 435.600 317.800 ;
        RECT 436.400 317.600 437.200 318.400 ;
        RECT 436.400 304.200 437.200 315.800 ;
        RECT 438.000 309.600 438.800 310.400 ;
        RECT 438.100 308.400 438.700 309.600 ;
        RECT 438.000 307.600 438.800 308.400 ;
        RECT 439.600 304.200 440.400 315.800 ;
        RECT 441.200 305.600 442.000 306.400 ;
        RECT 442.800 304.200 443.600 315.800 ;
        RECT 444.400 304.200 445.200 317.800 ;
        RECT 446.000 304.200 446.800 317.800 ;
        RECT 447.600 304.200 448.400 317.800 ;
        RECT 449.300 310.400 449.900 323.600 ;
        RECT 450.800 319.600 451.600 320.400 ;
        RECT 449.200 309.600 450.000 310.400 ;
        RECT 450.900 304.400 451.500 319.600 ;
        RECT 454.100 316.400 454.700 327.600 ;
        RECT 460.500 326.400 461.100 331.600 ;
        RECT 460.400 325.600 461.200 326.400 ;
        RECT 460.400 317.600 461.200 318.400 ;
        RECT 454.000 315.600 454.800 316.400 ;
        RECT 457.200 315.600 458.000 316.400 ;
        RECT 458.800 315.600 459.600 316.400 ;
        RECT 449.200 303.600 450.000 304.400 ;
        RECT 450.800 303.600 451.600 304.400 ;
        RECT 457.200 303.600 458.000 304.400 ;
        RECT 442.800 301.600 443.600 302.400 ;
        RECT 434.800 299.600 435.600 300.400 ;
        RECT 434.900 298.400 435.500 299.600 ;
        RECT 442.900 298.400 443.500 301.600 ;
        RECT 434.800 297.600 435.600 298.400 ;
        RECT 442.800 297.600 443.600 298.400 ;
        RECT 434.800 293.600 435.600 294.400 ;
        RECT 438.000 293.600 438.800 294.400 ;
        RECT 442.800 293.600 443.600 294.400 ;
        RECT 447.600 293.600 448.400 294.400 ;
        RECT 428.400 291.600 429.200 292.400 ;
        RECT 433.200 291.600 434.000 292.400 ;
        RECT 433.300 278.400 433.900 291.600 ;
        RECT 434.900 288.400 435.500 293.600 ;
        RECT 439.600 291.600 440.400 292.400 ;
        RECT 441.200 291.600 442.000 292.400 ;
        RECT 434.800 287.600 435.600 288.400 ;
        RECT 439.600 285.600 440.400 286.400 ;
        RECT 420.400 277.600 421.200 278.400 ;
        RECT 433.200 277.600 434.000 278.400 ;
        RECT 407.600 273.600 408.400 274.400 ;
        RECT 410.800 273.600 411.600 274.400 ;
        RECT 414.000 273.600 414.800 274.400 ;
        RECT 417.200 273.600 418.000 274.400 ;
        RECT 409.200 269.600 410.000 270.400 ;
        RECT 410.900 268.400 411.500 273.600 ;
        RECT 414.100 272.400 414.700 273.600 ;
        RECT 414.000 271.600 414.800 272.400 ;
        RECT 412.400 269.600 413.200 270.400 ;
        RECT 414.000 269.600 414.800 270.400 ;
        RECT 404.400 267.600 405.200 268.400 ;
        RECT 407.600 267.600 408.400 268.400 ;
        RECT 410.800 267.600 411.600 268.400 ;
        RECT 402.800 259.600 403.600 260.400 ;
        RECT 401.200 253.600 402.000 254.400 ;
        RECT 396.400 252.300 397.200 252.400 ;
        RECT 394.900 251.700 397.200 252.300 ;
        RECT 396.400 251.600 397.200 251.700 ;
        RECT 399.600 251.600 400.400 252.400 ;
        RECT 393.200 247.600 394.000 248.400 ;
        RECT 401.300 246.400 401.900 253.600 ;
        RECT 402.900 252.400 403.500 259.600 ;
        RECT 404.500 254.400 405.100 267.600 ;
        RECT 407.700 266.400 408.300 267.600 ;
        RECT 407.600 265.600 408.400 266.400 ;
        RECT 406.000 263.600 406.800 264.400 ;
        RECT 406.100 256.400 406.700 263.600 ;
        RECT 406.000 255.600 406.800 256.400 ;
        RECT 406.100 254.400 406.700 255.600 ;
        RECT 412.500 254.400 413.100 269.600 ;
        RECT 414.100 260.400 414.700 269.600 ;
        RECT 420.500 268.400 421.100 277.600 ;
        RECT 433.200 275.600 434.000 276.400 ;
        RECT 431.600 271.600 432.400 272.400 ;
        RECT 431.700 270.400 432.300 271.600 ;
        RECT 433.300 270.400 433.900 275.600 ;
        RECT 439.700 274.400 440.300 285.600 ;
        RECT 441.300 278.400 441.900 291.600 ;
        RECT 442.900 278.400 443.500 293.600 ;
        RECT 447.600 291.600 448.400 292.400 ;
        RECT 441.200 277.600 442.000 278.400 ;
        RECT 442.800 277.600 443.600 278.400 ;
        RECT 434.800 273.600 435.600 274.400 ;
        RECT 439.600 273.600 440.400 274.400 ;
        RECT 442.800 271.600 443.600 272.400 ;
        RECT 444.400 271.600 445.200 272.400 ;
        RECT 446.000 271.600 446.800 272.400 ;
        RECT 442.900 270.400 443.500 271.600 ;
        RECT 444.500 270.400 445.100 271.600 ;
        RECT 446.100 270.400 446.700 271.600 ;
        RECT 422.000 269.600 422.800 270.400 ;
        RECT 426.800 269.600 427.600 270.400 ;
        RECT 430.000 269.600 430.800 270.400 ;
        RECT 431.600 269.600 432.400 270.400 ;
        RECT 433.200 269.600 434.000 270.400 ;
        RECT 441.200 269.600 442.000 270.400 ;
        RECT 442.800 269.600 443.600 270.400 ;
        RECT 444.400 269.600 445.200 270.400 ;
        RECT 446.000 269.600 446.800 270.400 ;
        RECT 415.600 267.600 416.400 268.400 ;
        RECT 417.200 267.600 418.000 268.400 ;
        RECT 420.400 267.600 421.200 268.400 ;
        RECT 417.300 264.400 417.900 267.600 ;
        RECT 417.200 263.600 418.000 264.400 ;
        RECT 420.500 260.400 421.100 267.600 ;
        RECT 414.000 259.600 414.800 260.400 ;
        RECT 415.600 259.600 416.400 260.400 ;
        RECT 420.400 259.600 421.200 260.400 ;
        RECT 414.100 254.400 414.700 259.600 ;
        RECT 404.400 253.600 405.200 254.400 ;
        RECT 406.000 253.600 406.800 254.400 ;
        RECT 409.200 253.600 410.000 254.400 ;
        RECT 412.400 253.600 413.200 254.400 ;
        RECT 414.000 253.600 414.800 254.400 ;
        RECT 402.800 251.600 403.600 252.400 ;
        RECT 404.400 251.600 405.200 252.400 ;
        RECT 407.600 251.600 408.400 252.400 ;
        RECT 409.300 246.400 409.900 253.600 ;
        RECT 410.800 251.600 411.600 252.400 ;
        RECT 391.600 245.600 392.400 246.400 ;
        RECT 401.200 245.600 402.000 246.400 ;
        RECT 409.200 245.600 410.000 246.400 ;
        RECT 410.900 244.400 411.500 251.600 ;
        RECT 406.000 243.600 406.800 244.400 ;
        RECT 410.800 243.600 411.600 244.400 ;
        RECT 383.600 239.600 384.400 240.400 ;
        RECT 388.400 239.600 389.200 240.400 ;
        RECT 359.600 237.600 360.400 238.400 ;
        RECT 359.700 230.400 360.300 237.600 ;
        RECT 358.000 229.600 358.800 230.400 ;
        RECT 359.600 229.600 360.400 230.400 ;
        RECT 364.400 229.600 365.200 230.400 ;
        RECT 370.800 229.600 371.600 230.400 ;
        RECT 370.900 228.400 371.500 229.600 ;
        RECT 356.400 227.600 357.200 228.400 ;
        RECT 366.000 227.600 366.800 228.400 ;
        RECT 370.800 227.600 371.600 228.400 ;
        RECT 372.400 227.600 373.200 228.400 ;
        RECT 354.800 225.600 355.600 226.400 ;
        RECT 356.500 216.400 357.100 227.600 ;
        RECT 366.100 226.300 366.700 227.600 ;
        RECT 372.500 226.300 373.100 227.600 ;
        RECT 366.100 225.700 373.100 226.300 ;
        RECT 375.600 224.200 376.400 237.800 ;
        RECT 377.200 224.200 378.000 237.800 ;
        RECT 378.800 224.200 379.600 235.800 ;
        RECT 380.400 227.600 381.200 228.400 ;
        RECT 382.000 224.200 382.800 235.800 ;
        RECT 383.600 225.600 384.400 226.400 ;
        RECT 383.700 220.400 384.300 225.600 ;
        RECT 385.200 224.200 386.000 235.800 ;
        RECT 386.800 224.200 387.600 237.800 ;
        RECT 388.400 224.200 389.200 237.800 ;
        RECT 390.000 224.200 390.800 237.800 ;
        RECT 399.600 233.600 400.400 234.400 ;
        RECT 404.400 233.600 405.200 234.400 ;
        RECT 401.200 229.600 402.000 230.400 ;
        RECT 404.500 226.400 405.100 233.600 ;
        RECT 406.100 232.400 406.700 243.600 ;
        RECT 410.900 242.400 411.500 243.600 ;
        RECT 410.800 241.600 411.600 242.400 ;
        RECT 409.200 235.600 410.000 236.400 ;
        RECT 406.000 231.600 406.800 232.400 ;
        RECT 407.600 231.600 408.400 232.400 ;
        RECT 409.300 228.400 409.900 235.600 ;
        RECT 409.200 227.600 410.000 228.400 ;
        RECT 404.400 225.600 405.200 226.400 ;
        RECT 410.800 225.600 411.600 226.400 ;
        RECT 401.200 221.600 402.000 222.400 ;
        RECT 367.600 219.600 368.400 220.400 ;
        RECT 383.600 219.600 384.400 220.400 ;
        RECT 356.400 215.600 357.200 216.400 ;
        RECT 361.200 204.200 362.000 217.800 ;
        RECT 362.800 204.200 363.600 217.800 ;
        RECT 364.400 204.200 365.200 217.800 ;
        RECT 366.000 206.200 366.800 217.800 ;
        RECT 367.700 216.400 368.300 219.600 ;
        RECT 401.300 218.400 401.900 221.600 ;
        RECT 367.600 215.600 368.400 216.400 ;
        RECT 367.700 196.400 368.300 215.600 ;
        RECT 369.200 206.200 370.000 217.800 ;
        RECT 370.800 215.600 371.600 216.400 ;
        RECT 370.900 214.400 371.500 215.600 ;
        RECT 370.800 213.600 371.600 214.400 ;
        RECT 372.400 206.200 373.200 217.800 ;
        RECT 374.000 204.200 374.800 217.800 ;
        RECT 375.600 204.200 376.400 217.800 ;
        RECT 401.200 217.600 402.000 218.400 ;
        RECT 410.900 216.400 411.500 225.600 ;
        RECT 386.800 215.600 387.600 216.400 ;
        RECT 410.800 215.600 411.600 216.400 ;
        RECT 385.200 213.600 386.000 214.400 ;
        RECT 410.800 213.600 411.600 214.400 ;
        RECT 378.800 211.600 379.600 212.400 ;
        RECT 398.000 211.600 398.800 212.400 ;
        RECT 402.800 211.600 403.600 212.400 ;
        RECT 378.900 202.400 379.500 211.600 ;
        RECT 388.400 209.600 389.200 210.400 ;
        RECT 391.600 203.600 392.400 204.400 ;
        RECT 374.000 201.600 374.800 202.400 ;
        RECT 378.800 201.600 379.600 202.400 ;
        RECT 367.600 195.600 368.400 196.400 ;
        RECT 353.200 193.600 354.000 194.400 ;
        RECT 358.000 193.600 358.800 194.400 ;
        RECT 366.000 193.600 366.800 194.400 ;
        RECT 374.100 190.400 374.700 201.600 ;
        RECT 361.200 189.600 362.000 190.400 ;
        RECT 366.000 189.600 366.800 190.400 ;
        RECT 374.000 189.600 374.800 190.400 ;
        RECT 362.800 187.600 363.600 188.400 ;
        RECT 364.400 187.600 365.200 188.400 ;
        RECT 358.000 183.600 358.800 184.400 ;
        RECT 337.200 179.600 338.000 180.400 ;
        RECT 337.300 174.400 337.900 179.600 ;
        RECT 340.500 178.400 341.100 183.600 ;
        RECT 346.800 181.600 347.600 182.400 ;
        RECT 346.900 178.400 347.500 181.600 ;
        RECT 353.200 179.600 354.000 180.400 ;
        RECT 340.400 177.600 341.200 178.400 ;
        RECT 346.800 177.600 347.600 178.400 ;
        RECT 346.900 174.400 347.500 177.600 ;
        RECT 350.000 175.600 350.800 176.400 ;
        RECT 337.200 173.600 338.000 174.400 ;
        RECT 343.600 173.600 344.400 174.400 ;
        RECT 346.800 173.600 347.600 174.400 ;
        RECT 348.400 173.600 349.200 174.400 ;
        RECT 353.300 172.400 353.900 179.600 ;
        RECT 356.400 177.600 357.200 178.400 ;
        RECT 356.500 174.400 357.100 177.600 ;
        RECT 358.100 174.400 358.700 183.600 ;
        RECT 362.900 178.400 363.500 187.600 ;
        RECT 362.800 177.600 363.600 178.400 ;
        RECT 364.500 174.400 365.100 187.600 ;
        RECT 356.400 173.600 357.200 174.400 ;
        RECT 358.000 173.600 358.800 174.400 ;
        RECT 364.400 173.600 365.200 174.400 ;
        RECT 366.100 172.400 366.700 189.600 ;
        RECT 374.100 178.400 374.700 189.600 ;
        RECT 375.600 184.200 376.400 197.800 ;
        RECT 377.200 184.200 378.000 197.800 ;
        RECT 378.800 184.200 379.600 197.800 ;
        RECT 380.400 184.200 381.200 195.800 ;
        RECT 382.000 195.600 382.800 196.400 ;
        RECT 382.100 186.400 382.700 195.600 ;
        RECT 382.000 185.600 382.800 186.400 ;
        RECT 383.600 184.200 384.400 195.800 ;
        RECT 385.200 187.600 386.000 188.400 ;
        RECT 386.800 184.200 387.600 195.800 ;
        RECT 388.400 184.200 389.200 197.800 ;
        RECT 390.000 184.200 390.800 197.800 ;
        RECT 380.400 181.600 381.200 182.400 ;
        RECT 380.500 178.400 381.100 181.600 ;
        RECT 391.700 178.400 392.300 203.600 ;
        RECT 396.400 189.600 397.200 190.400 ;
        RECT 396.500 188.400 397.100 189.600 ;
        RECT 396.400 187.600 397.200 188.400 ;
        RECT 398.100 180.400 398.700 211.600 ;
        RECT 402.900 190.400 403.500 211.600 ;
        RECT 412.500 210.400 413.100 253.600 ;
        RECT 415.700 250.400 416.300 259.600 ;
        RECT 418.800 255.600 419.600 256.400 ;
        RECT 418.900 252.400 419.500 255.600 ;
        RECT 418.800 251.600 419.600 252.400 ;
        RECT 420.400 251.600 421.200 252.400 ;
        RECT 414.000 249.600 414.800 250.400 ;
        RECT 415.600 249.600 416.400 250.400 ;
        RECT 417.200 249.600 418.000 250.400 ;
        RECT 420.500 248.400 421.100 251.600 ;
        RECT 420.400 247.600 421.200 248.400 ;
        RECT 422.100 244.400 422.700 269.600 ;
        RECT 425.200 267.600 426.000 268.400 ;
        RECT 428.400 267.600 429.200 268.400 ;
        RECT 425.300 264.400 425.900 267.600 ;
        RECT 425.200 263.600 426.000 264.400 ;
        RECT 426.800 261.600 427.600 262.400 ;
        RECT 423.600 255.600 424.400 256.400 ;
        RECT 426.900 254.400 427.500 261.600 ;
        RECT 428.500 260.400 429.100 267.600 ;
        RECT 430.100 262.400 430.700 269.600 ;
        RECT 441.300 268.400 441.900 269.600 ;
        RECT 433.200 267.600 434.000 268.400 ;
        RECT 441.200 267.600 442.000 268.400 ;
        RECT 431.600 263.600 432.400 264.400 ;
        RECT 430.000 261.600 430.800 262.400 ;
        RECT 428.400 259.600 429.200 260.400 ;
        RECT 430.000 255.600 430.800 256.400 ;
        RECT 430.100 254.400 430.700 255.600 ;
        RECT 426.800 253.600 427.600 254.400 ;
        RECT 430.000 253.600 430.800 254.400 ;
        RECT 423.600 251.600 424.400 252.400 ;
        RECT 428.400 251.600 429.200 252.400 ;
        RECT 428.500 250.400 429.100 251.600 ;
        RECT 423.600 249.600 424.400 250.400 ;
        RECT 428.400 249.600 429.200 250.400 ;
        RECT 431.700 250.300 432.300 263.600 ;
        RECT 433.300 258.400 433.900 267.600 ;
        RECT 441.200 259.600 442.000 260.400 ;
        RECT 433.200 257.600 434.000 258.400 ;
        RECT 441.300 256.400 441.900 259.600 ;
        RECT 436.400 255.600 437.200 256.400 ;
        RECT 441.200 255.600 442.000 256.400 ;
        RECT 436.500 254.400 437.100 255.600 ;
        RECT 433.200 253.600 434.000 254.400 ;
        RECT 436.400 253.600 437.200 254.400 ;
        RECT 439.600 253.600 440.400 254.400 ;
        RECT 433.300 250.400 433.900 253.600 ;
        RECT 434.800 251.600 435.600 252.400 ;
        RECT 433.200 250.300 434.000 250.400 ;
        RECT 431.700 249.700 434.000 250.300 ;
        RECT 433.200 249.600 434.000 249.700 ;
        RECT 422.000 243.600 422.800 244.400 ;
        RECT 418.800 241.600 419.600 242.400 ;
        RECT 418.900 238.400 419.500 241.600 ;
        RECT 418.800 237.600 419.600 238.400 ;
        RECT 428.500 232.400 429.100 249.600 ;
        RECT 428.400 231.600 429.200 232.400 ;
        RECT 415.600 227.600 416.400 228.400 ;
        RECT 428.400 227.600 429.200 228.400 ;
        RECT 430.000 227.600 430.800 228.400 ;
        RECT 420.400 213.600 421.200 214.400 ;
        RECT 425.200 213.600 426.000 214.400 ;
        RECT 410.800 209.600 411.600 210.400 ;
        RECT 412.400 209.600 413.200 210.400 ;
        RECT 423.600 209.600 424.400 210.400 ;
        RECT 426.800 209.600 427.600 210.400 ;
        RECT 412.400 203.600 413.200 204.400 ;
        RECT 417.200 203.600 418.000 204.400 ;
        RECT 402.800 189.600 403.600 190.400 ;
        RECT 404.400 189.600 405.200 190.400 ;
        RECT 404.500 188.400 405.100 189.600 ;
        RECT 404.400 187.600 405.200 188.400 ;
        RECT 404.400 183.600 405.200 184.400 ;
        RECT 407.600 184.200 408.400 197.800 ;
        RECT 409.200 184.200 410.000 197.800 ;
        RECT 410.800 184.200 411.600 195.800 ;
        RECT 412.500 194.400 413.100 203.600 ;
        RECT 417.300 198.400 417.900 203.600 ;
        RECT 417.200 197.600 418.000 198.400 ;
        RECT 412.400 193.600 413.200 194.400 ;
        RECT 412.400 187.600 413.200 188.400 ;
        RECT 398.000 179.600 398.800 180.400 ;
        RECT 370.800 177.600 371.600 178.400 ;
        RECT 374.000 177.600 374.800 178.400 ;
        RECT 380.400 177.600 381.200 178.400 ;
        RECT 385.200 177.600 386.000 178.400 ;
        RECT 369.200 173.600 370.000 174.400 ;
        RECT 370.900 172.400 371.500 177.600 ;
        RECT 377.200 173.600 378.000 174.400 ;
        RECT 326.000 171.600 326.800 172.400 ;
        RECT 332.400 171.600 333.200 172.400 ;
        RECT 345.200 171.600 346.000 172.400 ;
        RECT 353.200 171.600 354.000 172.400 ;
        RECT 364.400 172.300 365.200 172.400 ;
        RECT 366.000 172.300 366.800 172.400 ;
        RECT 364.400 171.700 366.800 172.300 ;
        RECT 364.400 171.600 365.200 171.700 ;
        RECT 366.000 171.600 366.800 171.700 ;
        RECT 369.200 171.600 370.000 172.400 ;
        RECT 370.800 171.600 371.600 172.400 ;
        RECT 319.600 159.600 320.400 160.400 ;
        RECT 314.800 151.600 315.600 152.400 ;
        RECT 318.000 151.600 318.800 152.400 ;
        RECT 289.200 149.600 290.000 150.400 ;
        RECT 310.000 149.600 310.800 150.400 ;
        RECT 289.300 146.400 289.900 149.600 ;
        RECT 298.800 147.600 299.600 148.400 ;
        RECT 308.400 147.600 309.200 148.400 ;
        RECT 289.200 145.600 290.000 146.400 ;
        RECT 308.500 144.400 309.100 147.600 ;
        RECT 297.200 143.600 298.000 144.400 ;
        RECT 308.400 143.600 309.200 144.400 ;
        RECT 281.200 139.600 282.000 140.400 ;
        RECT 276.400 131.600 277.200 132.400 ;
        RECT 276.500 130.400 277.100 131.600 ;
        RECT 276.400 129.600 277.200 130.400 ;
        RECT 278.000 124.200 278.800 137.800 ;
        RECT 279.600 124.200 280.400 137.800 ;
        RECT 281.200 124.200 282.000 137.800 ;
        RECT 282.800 126.200 283.600 137.800 ;
        RECT 284.400 135.600 285.200 136.400 ;
        RECT 284.500 132.400 285.100 135.600 ;
        RECT 284.400 131.600 285.200 132.400 ;
        RECT 282.800 117.600 283.600 118.400 ;
        RECT 276.400 113.600 277.200 114.400 ;
        RECT 279.600 111.600 280.400 112.400 ;
        RECT 279.700 108.400 280.300 111.600 ;
        RECT 282.900 110.400 283.500 117.600 ;
        RECT 284.500 110.400 285.100 131.600 ;
        RECT 286.000 126.200 286.800 137.800 ;
        RECT 287.600 133.600 288.400 134.400 ;
        RECT 287.600 131.600 288.400 132.400 ;
        RECT 282.800 109.600 283.600 110.400 ;
        RECT 284.400 109.600 285.200 110.400 ;
        RECT 279.600 107.600 280.400 108.400 ;
        RECT 281.200 107.600 282.000 108.400 ;
        RECT 284.400 107.600 285.200 108.400 ;
        RECT 271.600 101.600 272.400 102.400 ;
        RECT 255.600 99.600 256.400 100.400 ;
        RECT 260.400 99.600 261.200 100.400 ;
        RECT 266.800 99.600 267.600 100.400 ;
        RECT 250.800 95.600 251.600 96.400 ;
        RECT 252.400 73.600 253.200 74.400 ;
        RECT 247.600 69.700 249.900 70.300 ;
        RECT 247.600 69.600 248.400 69.700 ;
        RECT 246.000 67.600 246.800 68.400 ;
        RECT 236.400 63.600 237.200 64.400 ;
        RECT 236.500 56.400 237.100 63.600 ;
        RECT 246.100 58.400 246.700 67.600 ;
        RECT 252.500 62.400 253.100 73.600 ;
        RECT 255.700 72.400 256.300 99.600 ;
        RECT 260.400 84.200 261.200 97.800 ;
        RECT 262.000 84.200 262.800 97.800 ;
        RECT 263.600 84.200 264.400 97.800 ;
        RECT 265.200 86.200 266.000 97.800 ;
        RECT 266.900 96.400 267.500 99.600 ;
        RECT 266.800 95.600 267.600 96.400 ;
        RECT 258.800 73.600 259.600 74.400 ;
        RECT 255.600 71.600 256.400 72.400 ;
        RECT 257.200 67.600 258.000 68.400 ;
        RECT 266.900 66.400 267.500 95.600 ;
        RECT 268.400 86.200 269.200 97.800 ;
        RECT 270.000 93.600 270.800 94.400 ;
        RECT 270.100 92.400 270.700 93.600 ;
        RECT 270.000 91.600 270.800 92.400 ;
        RECT 271.600 86.200 272.400 97.800 ;
        RECT 273.200 84.200 274.000 97.800 ;
        RECT 274.800 84.200 275.600 97.800 ;
        RECT 279.600 91.600 280.400 92.400 ;
        RECT 284.500 80.400 285.100 107.600 ;
        RECT 287.700 92.400 288.300 131.600 ;
        RECT 289.200 126.200 290.000 137.800 ;
        RECT 290.800 124.200 291.600 137.800 ;
        RECT 292.400 124.200 293.200 137.800 ;
        RECT 297.300 134.400 297.900 143.600 ;
        RECT 297.200 133.600 298.000 134.400 ;
        RECT 306.800 131.600 307.600 132.400 ;
        RECT 314.900 118.400 315.500 151.600 ;
        RECT 318.000 143.600 318.800 144.400 ;
        RECT 314.800 117.600 315.600 118.400 ;
        RECT 290.800 113.600 291.600 114.400 ;
        RECT 290.900 110.400 291.500 113.600 ;
        RECT 294.200 111.800 295.000 112.600 ;
        RECT 300.400 111.800 301.200 112.600 ;
        RECT 290.800 109.600 291.600 110.400 ;
        RECT 292.400 107.600 293.200 108.400 ;
        RECT 294.200 107.000 294.800 111.800 ;
        RECT 295.400 109.800 296.200 110.600 ;
        RECT 295.600 108.400 296.200 109.800 ;
        RECT 300.600 108.400 301.200 111.800 ;
        RECT 318.100 108.400 318.700 143.600 ;
        RECT 319.700 134.400 320.300 159.600 ;
        RECT 322.800 145.600 323.600 146.400 ;
        RECT 319.600 133.600 320.400 134.400 ;
        RECT 322.900 132.400 323.500 145.600 ;
        RECT 327.600 144.200 328.400 157.800 ;
        RECT 329.200 144.200 330.000 157.800 ;
        RECT 330.800 144.200 331.600 155.800 ;
        RECT 332.500 150.400 333.100 171.600 ;
        RECT 334.000 169.600 334.800 170.400 ;
        RECT 340.400 169.600 341.200 170.400 ;
        RECT 342.000 169.600 342.800 170.400 ;
        RECT 351.600 169.600 352.400 170.400 ;
        RECT 340.500 166.400 341.100 169.600 ;
        RECT 351.700 168.400 352.300 169.600 ;
        RECT 351.600 167.600 352.400 168.400 ;
        RECT 340.400 165.600 341.200 166.400 ;
        RECT 332.400 149.600 333.200 150.400 ;
        RECT 332.400 147.600 333.200 148.400 ;
        RECT 334.000 144.200 334.800 155.800 ;
        RECT 335.600 145.600 336.400 146.400 ;
        RECT 337.200 144.200 338.000 155.800 ;
        RECT 338.800 144.200 339.600 157.800 ;
        RECT 340.400 144.200 341.200 157.800 ;
        RECT 342.000 144.200 342.800 157.800 ;
        RECT 351.600 153.600 352.400 154.400 ;
        RECT 343.600 149.600 344.400 150.400 ;
        RECT 348.400 145.600 349.200 146.400 ;
        RECT 322.800 131.600 323.600 132.400 ;
        RECT 329.200 124.200 330.000 137.800 ;
        RECT 330.800 124.200 331.600 137.800 ;
        RECT 332.400 126.200 333.200 137.800 ;
        RECT 334.000 133.600 334.800 134.400 ;
        RECT 335.600 126.200 336.400 137.800 ;
        RECT 337.200 137.600 338.000 138.400 ;
        RECT 337.300 136.400 337.900 137.600 ;
        RECT 337.200 135.600 338.000 136.400 ;
        RECT 337.300 120.400 337.900 135.600 ;
        RECT 338.800 126.200 339.600 137.800 ;
        RECT 340.400 124.200 341.200 137.800 ;
        RECT 342.000 124.200 342.800 137.800 ;
        RECT 343.600 124.200 344.400 137.800 ;
        RECT 345.200 131.600 346.000 132.400 ;
        RECT 345.300 124.400 345.900 131.600 ;
        RECT 345.200 123.600 346.000 124.400 ;
        RECT 330.800 119.600 331.600 120.400 ;
        RECT 337.200 119.600 338.000 120.400 ;
        RECT 322.800 109.600 323.600 110.400 ;
        RECT 295.600 107.800 301.200 108.400 ;
        RECT 295.600 107.000 296.400 107.200 ;
        RECT 299.000 107.000 299.800 107.200 ;
        RECT 300.600 107.000 301.200 107.800 ;
        RECT 302.000 107.600 302.800 108.400 ;
        RECT 308.400 107.600 309.200 108.400 ;
        RECT 318.000 107.600 318.800 108.400 ;
        RECT 294.200 106.400 299.800 107.000 ;
        RECT 289.200 105.600 290.000 106.400 ;
        RECT 294.200 106.200 295.000 106.400 ;
        RECT 300.400 106.200 301.200 107.000 ;
        RECT 308.500 106.400 309.100 107.600 ;
        RECT 308.400 105.600 309.200 106.400 ;
        RECT 286.000 91.600 286.800 92.400 ;
        RECT 287.600 91.600 288.400 92.400 ;
        RECT 284.400 79.600 285.200 80.400 ;
        RECT 266.800 65.600 267.600 66.400 ;
        RECT 268.400 64.200 269.200 77.800 ;
        RECT 270.000 64.200 270.800 77.800 ;
        RECT 271.600 64.200 272.400 77.800 ;
        RECT 273.200 64.200 274.000 75.800 ;
        RECT 274.800 65.600 275.600 66.400 ;
        RECT 276.400 64.200 277.200 75.800 ;
        RECT 278.000 67.600 278.800 68.400 ;
        RECT 279.600 64.200 280.400 75.800 ;
        RECT 281.200 64.200 282.000 77.800 ;
        RECT 282.800 64.200 283.600 77.800 ;
        RECT 286.100 70.400 286.700 91.600 ;
        RECT 286.000 69.600 286.800 70.400 ;
        RECT 289.300 68.400 289.900 105.600 ;
        RECT 297.200 103.600 298.000 104.400 ;
        RECT 310.000 103.600 310.800 104.400 ;
        RECT 292.400 84.200 293.200 97.800 ;
        RECT 294.000 84.200 294.800 97.800 ;
        RECT 295.600 86.200 296.400 97.800 ;
        RECT 297.300 94.400 297.900 103.600 ;
        RECT 297.200 93.600 298.000 94.400 ;
        RECT 298.800 86.200 299.600 97.800 ;
        RECT 300.400 95.600 301.200 96.400 ;
        RECT 302.000 86.200 302.800 97.800 ;
        RECT 303.600 84.200 304.400 97.800 ;
        RECT 305.200 84.200 306.000 97.800 ;
        RECT 306.800 84.200 307.600 97.800 ;
        RECT 303.600 73.600 304.400 74.400 ;
        RECT 289.200 67.600 290.000 68.400 ;
        RECT 292.400 67.600 293.200 68.400 ;
        RECT 284.400 63.600 285.200 64.400 ;
        RECT 252.400 61.600 253.200 62.400 ;
        RECT 246.000 57.600 246.800 58.400 ;
        RECT 226.900 55.700 229.100 56.300 ;
        RECT 215.600 53.600 216.400 54.400 ;
        RECT 218.800 53.600 219.600 54.400 ;
        RECT 223.600 53.600 224.400 54.400 ;
        RECT 204.400 51.600 205.200 52.400 ;
        RECT 218.900 50.400 219.500 53.600 ;
        RECT 226.900 50.400 227.500 55.700 ;
        RECT 231.600 55.600 232.400 56.400 ;
        RECT 236.400 55.600 237.200 56.400 ;
        RECT 241.200 55.600 242.000 56.400 ;
        RECT 228.400 53.600 229.200 54.400 ;
        RECT 218.800 49.600 219.600 50.400 ;
        RECT 226.800 49.600 227.600 50.400 ;
        RECT 223.600 47.600 224.400 48.400 ;
        RECT 217.200 43.600 218.000 44.400 ;
        RECT 196.400 25.600 197.200 26.400 ;
        RECT 183.600 19.600 184.400 20.400 ;
        RECT 185.200 19.600 186.000 20.400 ;
        RECT 188.400 19.600 189.200 20.400 ;
        RECT 172.400 13.600 173.200 14.400 ;
        RECT 183.700 12.400 184.300 19.600 ;
        RECT 177.200 11.600 178.000 12.400 ;
        RECT 183.600 11.600 184.400 12.400 ;
        RECT 188.400 4.200 189.200 17.800 ;
        RECT 190.000 4.200 190.800 17.800 ;
        RECT 191.600 6.200 192.400 17.800 ;
        RECT 193.200 13.600 194.000 14.400 ;
        RECT 194.800 6.200 195.600 17.800 ;
        RECT 196.500 16.400 197.100 25.600 ;
        RECT 198.000 24.200 198.800 35.800 ;
        RECT 199.600 27.600 200.400 28.400 ;
        RECT 201.200 24.200 202.000 35.800 ;
        RECT 202.800 24.200 203.600 37.800 ;
        RECT 204.400 24.200 205.200 37.800 ;
        RECT 217.300 32.400 217.900 43.600 ;
        RECT 223.700 32.400 224.300 47.600 ;
        RECT 217.200 31.600 218.000 32.400 ;
        RECT 222.000 31.600 222.800 32.400 ;
        RECT 223.600 31.600 224.400 32.400 ;
        RECT 217.200 29.600 218.000 30.400 ;
        RECT 220.400 29.600 221.200 30.400 ;
        RECT 222.100 28.400 222.700 31.600 ;
        RECT 228.500 28.400 229.100 53.600 ;
        RECT 231.700 50.400 232.300 55.600 ;
        RECT 238.000 53.600 238.800 54.400 ;
        RECT 246.000 51.600 246.800 52.400 ;
        RECT 231.600 49.600 232.400 50.400 ;
        RECT 236.400 49.600 237.200 50.400 ;
        RECT 250.800 44.200 251.600 57.800 ;
        RECT 252.400 44.200 253.200 57.800 ;
        RECT 254.000 46.200 254.800 57.800 ;
        RECT 255.600 53.600 256.400 54.400 ;
        RECT 255.700 50.400 256.300 53.600 ;
        RECT 255.600 49.600 256.400 50.400 ;
        RECT 257.200 46.200 258.000 57.800 ;
        RECT 258.800 55.600 259.600 56.400 ;
        RECT 246.000 39.600 246.800 40.400 ;
        RECT 222.000 27.600 222.800 28.400 ;
        RECT 228.400 27.600 229.200 28.400 ;
        RECT 215.600 25.600 216.400 26.400 ;
        RECT 231.600 25.600 232.400 26.400 ;
        RECT 196.400 15.600 197.200 16.400 ;
        RECT 198.000 6.200 198.800 17.800 ;
        RECT 199.600 4.200 200.400 17.800 ;
        RECT 201.200 4.200 202.000 17.800 ;
        RECT 202.800 4.200 203.600 17.800 ;
        RECT 215.700 12.400 216.300 25.600 ;
        RECT 217.200 23.600 218.000 24.400 ;
        RECT 223.600 23.600 224.400 24.400 ;
        RECT 217.300 14.400 217.900 23.600 ;
        RECT 223.700 14.400 224.300 23.600 ;
        RECT 231.700 22.400 232.300 25.600 ;
        RECT 241.200 24.200 242.000 37.800 ;
        RECT 242.800 24.200 243.600 37.800 ;
        RECT 244.400 24.200 245.200 35.800 ;
        RECT 246.100 28.400 246.700 39.600 ;
        RECT 246.000 27.600 246.800 28.400 ;
        RECT 247.600 24.200 248.400 35.800 ;
        RECT 249.200 25.600 250.000 26.400 ;
        RECT 231.600 21.600 232.400 22.400 ;
        RECT 249.300 18.400 249.900 25.600 ;
        RECT 250.800 24.200 251.600 35.800 ;
        RECT 252.400 24.200 253.200 37.800 ;
        RECT 254.000 24.200 254.800 37.800 ;
        RECT 255.600 24.200 256.400 37.800 ;
        RECT 257.200 29.600 258.000 30.400 ;
        RECT 252.400 21.600 253.200 22.400 ;
        RECT 252.500 18.400 253.100 21.600 ;
        RECT 258.900 18.400 259.500 55.600 ;
        RECT 260.400 46.200 261.200 57.800 ;
        RECT 262.000 44.200 262.800 57.800 ;
        RECT 263.600 44.200 264.400 57.800 ;
        RECT 265.200 44.200 266.000 57.800 ;
        RECT 274.800 55.600 275.600 56.400 ;
        RECT 278.000 53.600 278.800 54.400 ;
        RECT 270.000 51.600 270.800 52.400 ;
        RECT 279.600 51.600 280.400 52.400 ;
        RECT 270.100 38.400 270.700 51.600 ;
        RECT 284.500 50.400 285.100 63.600 ;
        RECT 289.300 54.400 289.900 67.600 ;
        RECT 310.100 64.400 310.700 103.600 ;
        RECT 316.400 93.600 317.400 94.400 ;
        RECT 311.600 69.600 312.400 70.400 ;
        RECT 294.000 63.600 294.800 64.400 ;
        RECT 310.000 63.600 310.800 64.400 ;
        RECT 289.200 53.600 290.000 54.400 ;
        RECT 289.200 51.600 290.000 52.400 ;
        RECT 282.800 49.600 283.600 50.400 ;
        RECT 284.400 49.600 285.200 50.400 ;
        RECT 289.300 44.400 289.900 51.600 ;
        RECT 294.100 50.400 294.700 63.600 ;
        RECT 311.700 58.400 312.300 69.600 ;
        RECT 313.200 64.200 314.000 77.800 ;
        RECT 314.800 64.200 315.600 77.800 ;
        RECT 316.400 64.200 317.200 77.800 ;
        RECT 318.000 64.200 318.800 75.800 ;
        RECT 319.600 65.600 320.400 66.400 ;
        RECT 321.200 64.200 322.000 75.800 ;
        RECT 322.900 70.400 323.500 109.600 ;
        RECT 324.400 104.200 325.200 117.800 ;
        RECT 326.000 104.200 326.800 117.800 ;
        RECT 327.600 104.200 328.400 117.800 ;
        RECT 329.200 104.200 330.000 115.800 ;
        RECT 330.900 106.400 331.500 119.600 ;
        RECT 330.800 105.600 331.600 106.400 ;
        RECT 330.900 96.400 331.500 105.600 ;
        RECT 332.400 104.200 333.200 115.800 ;
        RECT 334.000 107.600 334.800 108.400 ;
        RECT 335.600 104.200 336.400 115.800 ;
        RECT 337.200 104.200 338.000 117.800 ;
        RECT 338.800 104.200 339.600 117.800 ;
        RECT 343.600 109.600 344.400 110.400 ;
        RECT 348.500 100.400 349.100 145.600 ;
        RECT 353.300 132.400 353.900 171.600 ;
        RECT 354.800 169.600 355.600 170.400 ;
        RECT 362.800 169.600 363.600 170.400 ;
        RECT 354.900 152.400 355.500 169.600 ;
        RECT 361.200 167.600 362.000 168.400 ;
        RECT 356.400 155.600 357.200 156.400 ;
        RECT 354.800 151.600 355.600 152.400 ;
        RECT 354.800 147.600 355.600 148.400 ;
        RECT 354.800 145.600 355.600 146.400 ;
        RECT 354.900 136.400 355.500 145.600 ;
        RECT 354.800 135.600 355.600 136.400 ;
        RECT 356.500 132.400 357.100 155.600 ;
        RECT 358.000 153.600 358.800 154.400 ;
        RECT 359.600 149.600 360.400 150.400 ;
        RECT 359.700 136.400 360.300 149.600 ;
        RECT 359.600 135.600 360.400 136.400 ;
        RECT 353.200 131.600 354.000 132.400 ;
        RECT 356.400 132.300 357.200 132.400 ;
        RECT 354.900 131.700 357.200 132.300 ;
        RECT 353.200 123.600 354.000 124.400 ;
        RECT 350.000 109.600 350.800 110.400 ;
        RECT 350.100 108.400 350.700 109.600 ;
        RECT 353.300 108.400 353.900 123.600 ;
        RECT 354.900 110.400 355.500 131.700 ;
        RECT 356.400 131.600 357.200 131.700 ;
        RECT 354.800 109.600 355.600 110.400 ;
        RECT 350.000 107.600 350.800 108.400 ;
        RECT 353.200 107.600 354.000 108.400 ;
        RECT 358.000 103.600 358.800 104.400 ;
        RECT 348.400 99.600 349.200 100.400 ;
        RECT 332.400 97.600 333.200 98.400 ;
        RECT 330.800 95.600 331.600 96.400 ;
        RECT 326.000 83.600 326.800 84.400 ;
        RECT 342.000 84.200 342.800 97.800 ;
        RECT 343.600 84.200 344.400 97.800 ;
        RECT 345.200 84.200 346.000 97.800 ;
        RECT 346.800 86.200 347.600 97.800 ;
        RECT 348.500 96.400 349.100 99.600 ;
        RECT 348.400 95.600 349.200 96.400 ;
        RECT 350.000 86.200 350.800 97.800 ;
        RECT 351.600 93.600 352.400 94.400 ;
        RECT 353.200 86.200 354.000 97.800 ;
        RECT 354.800 84.200 355.600 97.800 ;
        RECT 356.400 84.200 357.200 97.800 ;
        RECT 358.100 92.400 358.700 103.600 ;
        RECT 358.000 91.600 358.800 92.400 ;
        RECT 358.100 90.800 358.700 91.600 ;
        RECT 358.000 90.000 358.800 90.800 ;
        RECT 326.100 80.400 326.700 83.600 ;
        RECT 326.000 79.600 326.800 80.400 ;
        RECT 337.200 79.600 338.000 80.400 ;
        RECT 359.600 79.600 360.400 80.400 ;
        RECT 322.800 69.600 323.600 70.400 ;
        RECT 322.800 67.600 323.600 68.400 ;
        RECT 322.900 66.400 323.500 67.600 ;
        RECT 322.800 65.600 323.600 66.400 ;
        RECT 324.400 64.200 325.200 75.800 ;
        RECT 326.000 64.200 326.800 77.800 ;
        RECT 327.600 64.200 328.400 77.800 ;
        RECT 337.300 68.400 337.900 79.600 ;
        RECT 354.800 73.600 355.600 74.400 ;
        RECT 342.000 71.600 342.800 72.400 ;
        RECT 345.400 71.800 346.200 72.600 ;
        RECT 351.600 71.800 352.400 72.600 ;
        RECT 338.800 69.600 339.600 70.400 ;
        RECT 337.200 67.600 338.000 68.400 ;
        RECT 338.800 63.600 339.600 64.400 ;
        RECT 297.200 51.600 298.000 52.400 ;
        RECT 294.000 49.600 294.800 50.400 ;
        RECT 274.800 43.600 275.600 44.400 ;
        RECT 279.600 43.600 280.400 44.400 ;
        RECT 287.600 43.600 288.400 44.400 ;
        RECT 289.200 43.600 290.000 44.400 ;
        RECT 270.000 37.600 270.800 38.400 ;
        RECT 273.200 29.600 274.000 30.400 ;
        RECT 265.200 23.600 266.000 24.400 ;
        RECT 260.400 19.600 261.200 20.400 ;
        RECT 217.200 13.600 218.000 14.400 ;
        RECT 223.600 13.600 224.400 14.400 ;
        RECT 204.400 11.600 205.200 12.400 ;
        RECT 215.600 11.600 216.400 12.400 ;
        RECT 223.600 11.600 224.400 12.400 ;
        RECT 228.400 4.200 229.200 17.800 ;
        RECT 230.000 4.200 230.800 17.800 ;
        RECT 231.600 6.200 232.400 17.800 ;
        RECT 233.200 13.600 234.000 14.400 ;
        RECT 234.800 6.200 235.600 17.800 ;
        RECT 236.400 17.600 237.200 18.400 ;
        RECT 236.500 16.400 237.100 17.600 ;
        RECT 236.400 15.600 237.200 16.400 ;
        RECT 238.000 6.200 238.800 17.800 ;
        RECT 239.600 4.200 240.400 17.800 ;
        RECT 241.200 4.200 242.000 17.800 ;
        RECT 242.800 4.200 243.600 17.800 ;
        RECT 249.200 17.600 250.000 18.400 ;
        RECT 252.400 17.600 253.200 18.400 ;
        RECT 258.800 17.600 259.600 18.400 ;
        RECT 260.500 12.400 261.100 19.600 ;
        RECT 265.300 12.400 265.900 23.600 ;
        RECT 273.300 12.400 273.900 29.600 ;
        RECT 274.900 20.400 275.500 43.600 ;
        RECT 279.700 40.400 280.300 43.600 ;
        RECT 279.600 39.600 280.400 40.400 ;
        RECT 279.600 24.200 280.400 37.800 ;
        RECT 281.200 24.200 282.000 37.800 ;
        RECT 282.800 24.200 283.600 35.800 ;
        RECT 284.400 29.600 285.200 30.400 ;
        RECT 284.500 28.400 285.100 29.600 ;
        RECT 284.400 27.600 285.200 28.400 ;
        RECT 286.000 24.200 286.800 35.800 ;
        RECT 287.700 28.400 288.300 43.600 ;
        RECT 287.600 27.600 288.400 28.400 ;
        RECT 287.600 25.600 288.400 26.400 ;
        RECT 287.700 22.300 288.300 25.600 ;
        RECT 289.200 24.200 290.000 35.800 ;
        RECT 290.800 24.200 291.600 37.800 ;
        RECT 292.400 24.200 293.200 37.800 ;
        RECT 294.000 24.200 294.800 37.800 ;
        RECT 295.600 30.300 296.400 30.400 ;
        RECT 297.300 30.300 297.900 51.600 ;
        RECT 303.600 44.200 304.400 57.800 ;
        RECT 305.200 44.200 306.000 57.800 ;
        RECT 306.800 46.200 307.600 57.800 ;
        RECT 308.400 53.600 309.200 54.400 ;
        RECT 310.000 46.200 310.800 57.800 ;
        RECT 311.600 57.600 312.400 58.400 ;
        RECT 311.600 55.600 312.400 56.400 ;
        RECT 295.600 29.700 297.900 30.300 ;
        RECT 295.600 29.600 296.400 29.700 ;
        RECT 286.100 21.700 288.300 22.300 ;
        RECT 274.800 19.600 275.600 20.400 ;
        RECT 286.100 18.400 286.700 21.700 ;
        RECT 260.400 11.600 261.200 12.400 ;
        RECT 265.200 11.600 266.000 12.400 ;
        RECT 273.200 11.600 274.000 12.400 ;
        RECT 278.000 4.200 278.800 17.800 ;
        RECT 279.600 4.200 280.400 17.800 ;
        RECT 281.200 6.200 282.000 17.800 ;
        RECT 282.800 13.600 283.600 14.400 ;
        RECT 284.400 6.200 285.200 17.800 ;
        RECT 286.000 17.600 286.800 18.400 ;
        RECT 286.100 16.400 286.700 17.600 ;
        RECT 286.000 15.600 286.800 16.400 ;
        RECT 287.600 6.200 288.400 17.800 ;
        RECT 289.200 4.200 290.000 17.800 ;
        RECT 290.800 4.200 291.600 17.800 ;
        RECT 292.400 4.200 293.200 17.800 ;
        RECT 297.300 12.400 297.900 29.700 ;
        RECT 303.600 27.600 304.600 28.400 ;
        RECT 310.000 25.600 310.800 26.400 ;
        RECT 310.100 12.400 310.700 25.600 ;
        RECT 311.700 18.400 312.300 55.600 ;
        RECT 313.200 46.200 314.000 57.800 ;
        RECT 313.200 43.600 314.000 44.400 ;
        RECT 314.800 44.200 315.600 57.800 ;
        RECT 316.400 44.200 317.200 57.800 ;
        RECT 318.000 44.200 318.800 57.800 ;
        RECT 319.600 57.600 320.400 58.400 ;
        RECT 326.000 57.600 326.800 58.400 ;
        RECT 319.700 52.400 320.300 57.600 ;
        RECT 319.600 51.600 320.400 52.400 ;
        RECT 313.300 38.400 313.900 43.600 ;
        RECT 313.200 37.600 314.000 38.400 ;
        RECT 316.400 31.800 317.200 32.600 ;
        RECT 323.000 31.800 323.800 32.600 ;
        RECT 314.800 29.600 315.600 30.400 ;
        RECT 316.400 28.400 317.000 31.800 ;
        RECT 320.400 28.400 321.200 28.600 ;
        RECT 314.800 27.600 315.600 28.400 ;
        RECT 316.400 27.800 321.200 28.400 ;
        RECT 316.400 27.000 317.000 27.800 ;
        RECT 317.800 27.000 318.600 27.200 ;
        RECT 321.200 27.000 322.000 27.200 ;
        RECT 323.200 27.000 323.800 31.800 ;
        RECT 326.100 30.400 326.700 57.600 ;
        RECT 338.900 52.400 339.500 63.600 ;
        RECT 342.100 58.400 342.700 71.600 ;
        RECT 343.600 67.600 344.400 68.400 ;
        RECT 342.000 57.600 342.800 58.400 ;
        RECT 340.400 53.600 341.200 54.400 ;
        RECT 330.800 51.600 331.600 52.400 ;
        RECT 337.200 51.600 338.000 52.400 ;
        RECT 338.800 51.600 339.600 52.400 ;
        RECT 327.600 49.600 328.400 50.400 ;
        RECT 330.900 38.400 331.500 51.600 ;
        RECT 337.300 50.300 337.900 51.600 ;
        RECT 337.300 49.700 339.500 50.300 ;
        RECT 334.000 43.600 334.800 44.400 ;
        RECT 330.800 37.600 331.600 38.400 ;
        RECT 327.600 31.600 328.400 32.400 ;
        RECT 327.700 30.400 328.300 31.600 ;
        RECT 326.000 29.600 326.800 30.400 ;
        RECT 327.600 29.600 328.400 30.400 ;
        RECT 316.400 26.200 317.200 27.000 ;
        RECT 317.800 26.400 322.000 27.000 ;
        RECT 323.000 26.200 323.800 27.000 ;
        RECT 334.100 20.400 334.700 43.600 ;
        RECT 338.900 38.400 339.500 49.700 ;
        RECT 340.500 46.400 341.100 53.600 ;
        RECT 343.700 50.400 344.300 67.600 ;
        RECT 345.400 67.000 346.000 71.800 ;
        RECT 346.600 69.800 347.400 70.600 ;
        RECT 346.800 68.400 347.400 69.800 ;
        RECT 351.800 68.400 352.400 71.800 ;
        RECT 358.000 69.600 358.800 70.400 ;
        RECT 359.700 68.400 360.300 79.600 ;
        RECT 361.300 78.400 361.900 167.600 ;
        RECT 362.800 150.300 363.600 150.400 ;
        RECT 364.500 150.300 365.100 171.600 ;
        RECT 369.300 170.400 369.900 171.600 ;
        RECT 369.200 169.600 370.000 170.400 ;
        RECT 370.900 156.400 371.500 171.600 ;
        RECT 385.300 170.400 385.900 177.600 ;
        RECT 374.000 169.600 374.800 170.400 ;
        RECT 380.400 169.600 381.200 170.400 ;
        RECT 385.200 169.600 386.000 170.400 ;
        RECT 374.100 158.400 374.700 169.600 ;
        RECT 383.600 167.600 384.400 168.400 ;
        RECT 380.400 165.600 381.200 166.400 ;
        RECT 380.500 158.400 381.100 165.600 ;
        RECT 374.000 157.600 374.800 158.400 ;
        RECT 380.400 157.600 381.200 158.400 ;
        RECT 370.800 155.600 371.600 156.400 ;
        RECT 366.000 153.600 366.800 154.400 ;
        RECT 362.800 149.700 365.100 150.300 ;
        RECT 362.800 149.600 363.600 149.700 ;
        RECT 362.900 138.400 363.500 149.600 ;
        RECT 366.100 148.400 366.700 153.600 ;
        RECT 369.200 151.600 370.000 152.400 ;
        RECT 370.800 151.600 371.600 152.400 ;
        RECT 377.200 151.600 378.000 152.400 ;
        RECT 364.400 147.600 365.200 148.400 ;
        RECT 366.000 147.600 366.800 148.400 ;
        RECT 364.500 144.400 365.100 147.600 ;
        RECT 369.300 146.400 369.900 151.600 ;
        RECT 369.200 145.600 370.000 146.400 ;
        RECT 364.400 143.600 365.200 144.400 ;
        RECT 369.200 143.600 370.000 144.400 ;
        RECT 362.800 137.600 363.600 138.400 ;
        RECT 364.500 134.400 365.100 143.600 ;
        RECT 369.300 140.400 369.900 143.600 ;
        RECT 369.200 139.600 370.000 140.400 ;
        RECT 369.200 137.600 370.000 138.400 ;
        RECT 362.800 133.600 363.600 134.400 ;
        RECT 364.400 133.600 365.200 134.400 ;
        RECT 367.600 133.600 368.400 134.400 ;
        RECT 369.300 132.400 369.900 137.600 ;
        RECT 366.000 131.600 366.800 132.400 ;
        RECT 369.200 131.600 370.000 132.400 ;
        RECT 369.300 116.400 369.900 131.600 ;
        RECT 366.000 115.600 366.800 116.400 ;
        RECT 369.200 115.600 370.000 116.400 ;
        RECT 364.400 107.600 365.200 108.400 ;
        RECT 362.800 105.600 363.600 106.400 ;
        RECT 362.900 102.400 363.500 105.600 ;
        RECT 362.800 101.600 363.600 102.400 ;
        RECT 361.200 77.600 362.000 78.400 ;
        RECT 364.400 77.600 365.200 78.400 ;
        RECT 364.500 72.400 365.100 77.600 ;
        RECT 364.400 71.600 365.200 72.400 ;
        RECT 366.100 70.400 366.700 115.600 ;
        RECT 369.200 113.600 370.000 114.400 ;
        RECT 369.300 112.400 369.900 113.600 ;
        RECT 369.200 111.600 370.000 112.400 ;
        RECT 369.200 107.600 370.000 108.400 ;
        RECT 369.200 91.600 370.000 92.400 ;
        RECT 367.600 79.600 368.400 80.400 ;
        RECT 366.000 69.600 366.800 70.400 ;
        RECT 346.800 67.800 352.400 68.400 ;
        RECT 346.800 67.000 347.600 67.200 ;
        RECT 350.200 67.000 351.000 67.200 ;
        RECT 351.800 67.000 352.400 67.800 ;
        RECT 353.200 67.600 354.000 68.400 ;
        RECT 356.400 67.600 357.200 68.400 ;
        RECT 359.600 67.600 360.400 68.400 ;
        RECT 361.200 67.600 362.000 68.400 ;
        RECT 345.400 66.400 351.000 67.000 ;
        RECT 345.400 66.200 346.200 66.400 ;
        RECT 351.600 66.200 352.400 67.000 ;
        RECT 366.100 66.400 366.700 69.600 ;
        RECT 367.700 68.400 368.300 79.600 ;
        RECT 370.900 72.400 371.500 151.600 ;
        RECT 374.000 149.600 374.800 150.400 ;
        RECT 375.600 149.600 376.400 150.400 ;
        RECT 380.400 149.600 381.200 150.400 ;
        RECT 374.100 144.400 374.700 149.600 ;
        RECT 375.700 148.400 376.300 149.600 ;
        RECT 375.600 147.600 376.400 148.400 ;
        RECT 374.000 143.600 374.800 144.400 ;
        RECT 380.500 142.400 381.100 149.600 ;
        RECT 383.700 148.400 384.300 167.600 ;
        RECT 390.000 166.200 390.800 177.800 ;
        RECT 391.600 177.600 392.400 178.400 ;
        RECT 398.000 175.600 398.800 176.400 ;
        RECT 398.100 172.600 398.700 175.600 ;
        RECT 398.000 171.800 398.800 172.600 ;
        RECT 399.600 166.200 400.400 177.800 ;
        RECT 401.200 173.600 402.000 174.400 ;
        RECT 402.800 170.200 403.600 175.800 ;
        RECT 404.500 174.400 405.100 183.600 ;
        RECT 412.500 182.400 413.100 187.600 ;
        RECT 414.000 184.200 414.800 195.800 ;
        RECT 415.600 185.600 416.400 186.400 ;
        RECT 417.200 184.200 418.000 195.800 ;
        RECT 418.800 184.200 419.600 197.800 ;
        RECT 420.400 184.200 421.200 197.800 ;
        RECT 422.000 184.200 422.800 197.800 ;
        RECT 412.400 181.600 413.200 182.400 ;
        RECT 423.700 182.300 424.300 209.600 ;
        RECT 422.100 181.700 424.300 182.300 ;
        RECT 410.800 175.600 411.600 176.400 ;
        RECT 414.000 175.600 414.800 176.400 ;
        RECT 417.200 175.600 418.000 176.400 ;
        RECT 404.400 173.600 405.200 174.400 ;
        RECT 404.500 158.400 405.100 173.600 ;
        RECT 414.100 172.400 414.700 175.600 ;
        RECT 417.300 174.400 417.900 175.600 ;
        RECT 415.600 173.600 416.400 174.400 ;
        RECT 417.200 173.600 418.000 174.400 ;
        RECT 406.000 171.600 406.800 172.400 ;
        RECT 414.000 171.600 414.800 172.400 ;
        RECT 406.100 162.400 406.700 171.600 ;
        RECT 409.200 169.600 410.000 170.400 ;
        RECT 415.700 168.400 416.300 173.600 ;
        RECT 417.200 171.600 418.000 172.400 ;
        RECT 417.300 170.400 417.900 171.600 ;
        RECT 417.200 169.600 418.000 170.400 ;
        RECT 415.600 167.600 416.400 168.400 ;
        RECT 420.400 167.600 421.200 168.400 ;
        RECT 407.600 163.600 408.400 164.400 ;
        RECT 406.000 161.600 406.800 162.400 ;
        RECT 404.400 157.600 405.200 158.400 ;
        RECT 390.000 155.600 390.800 156.400 ;
        RECT 402.800 155.600 403.600 156.400 ;
        RECT 390.100 152.400 390.700 155.600 ;
        RECT 398.000 153.600 398.800 154.400 ;
        RECT 404.400 153.600 405.200 154.400 ;
        RECT 385.200 151.600 386.000 152.400 ;
        RECT 388.400 151.600 389.200 152.400 ;
        RECT 390.000 151.600 390.800 152.400 ;
        RECT 396.400 151.600 397.200 152.400 ;
        RECT 401.200 151.600 402.000 152.400 ;
        RECT 385.200 149.600 386.000 150.400 ;
        RECT 393.200 149.600 394.000 150.400 ;
        RECT 399.600 149.600 400.400 150.400 ;
        RECT 382.000 147.600 382.800 148.400 ;
        RECT 383.600 147.600 384.400 148.400 ;
        RECT 390.000 147.600 390.800 148.400 ;
        RECT 380.400 141.600 381.200 142.400 ;
        RECT 393.300 140.400 393.900 149.600 ;
        RECT 394.800 147.600 395.600 148.400 ;
        RECT 393.200 139.600 394.000 140.400 ;
        RECT 382.000 135.600 382.800 136.400 ;
        RECT 377.200 133.600 378.000 134.400 ;
        RECT 382.100 132.400 382.700 135.600 ;
        RECT 382.000 131.600 382.800 132.400 ;
        RECT 377.200 129.600 378.000 130.400 ;
        RECT 374.000 127.600 374.800 128.400 ;
        RECT 377.300 122.400 377.900 129.600 ;
        RECT 386.800 124.200 387.600 137.800 ;
        RECT 388.400 124.200 389.200 137.800 ;
        RECT 390.000 126.200 390.800 137.800 ;
        RECT 391.600 133.600 392.400 134.400 ;
        RECT 393.200 126.200 394.000 137.800 ;
        RECT 394.800 135.600 395.600 136.400 ;
        RECT 396.400 126.200 397.200 137.800 ;
        RECT 394.800 123.600 395.600 124.400 ;
        RECT 398.000 124.200 398.800 137.800 ;
        RECT 399.600 124.200 400.400 137.800 ;
        RECT 401.200 124.200 402.000 137.800 ;
        RECT 377.200 121.600 378.000 122.400 ;
        RECT 378.800 104.200 379.600 117.800 ;
        RECT 380.400 104.200 381.200 117.800 ;
        RECT 382.000 104.200 382.800 115.800 ;
        RECT 383.600 107.600 384.400 108.400 ;
        RECT 385.200 104.200 386.000 115.800 ;
        RECT 386.800 109.600 387.600 110.400 ;
        RECT 386.900 106.400 387.500 109.600 ;
        RECT 386.800 105.600 387.600 106.400 ;
        RECT 386.900 100.400 387.500 105.600 ;
        RECT 388.400 104.200 389.200 115.800 ;
        RECT 390.000 104.200 390.800 117.800 ;
        RECT 391.600 104.200 392.400 117.800 ;
        RECT 393.200 104.200 394.000 117.800 ;
        RECT 394.900 110.400 395.500 123.600 ;
        RECT 401.200 121.600 402.000 122.400 ;
        RECT 394.800 109.600 395.600 110.400 ;
        RECT 382.000 99.600 382.800 100.400 ;
        RECT 386.800 99.600 387.600 100.400 ;
        RECT 374.000 84.200 374.800 97.800 ;
        RECT 375.600 84.200 376.400 97.800 ;
        RECT 377.200 86.200 378.000 97.800 ;
        RECT 378.800 93.600 379.600 94.400 ;
        RECT 378.900 82.400 379.500 93.600 ;
        RECT 380.400 86.200 381.200 97.800 ;
        RECT 382.100 96.400 382.700 99.600 ;
        RECT 401.300 98.400 401.900 121.600 ;
        RECT 404.500 110.300 405.100 153.600 ;
        RECT 407.700 152.400 408.300 163.600 ;
        RECT 410.800 161.600 411.600 162.400 ;
        RECT 409.200 157.600 410.000 158.400 ;
        RECT 407.600 151.600 408.400 152.400 ;
        RECT 406.000 149.600 406.800 150.400 ;
        RECT 406.100 132.400 406.700 149.600 ;
        RECT 409.300 148.400 409.900 157.600 ;
        RECT 410.900 150.400 411.500 161.600 ;
        RECT 412.400 157.600 413.200 158.400 ;
        RECT 410.800 149.600 411.600 150.400 ;
        RECT 409.200 147.600 410.000 148.400 ;
        RECT 409.300 134.400 409.900 147.600 ;
        RECT 410.900 138.400 411.500 149.600 ;
        RECT 412.500 148.400 413.100 157.600 ;
        RECT 414.000 151.600 414.800 152.400 ;
        RECT 420.500 148.400 421.100 167.600 ;
        RECT 412.400 147.600 413.200 148.400 ;
        RECT 417.200 147.600 418.000 148.400 ;
        RECT 420.400 147.600 421.200 148.400 ;
        RECT 412.400 139.600 413.200 140.400 ;
        RECT 410.800 137.600 411.600 138.400 ;
        RECT 409.200 133.600 410.000 134.400 ;
        RECT 406.000 131.600 406.800 132.400 ;
        RECT 410.800 127.600 411.600 128.400 ;
        RECT 406.000 121.600 406.800 122.400 ;
        RECT 406.100 118.400 406.700 121.600 ;
        RECT 406.000 117.600 406.800 118.400 ;
        RECT 404.500 109.700 406.700 110.300 ;
        RECT 402.800 103.600 403.600 104.400 ;
        RECT 404.400 103.600 405.200 104.400 ;
        RECT 402.900 102.400 403.500 103.600 ;
        RECT 402.800 101.600 403.600 102.400 ;
        RECT 382.000 95.600 382.800 96.400 ;
        RECT 383.600 86.200 384.400 97.800 ;
        RECT 385.200 84.200 386.000 97.800 ;
        RECT 386.800 84.200 387.600 97.800 ;
        RECT 388.400 84.200 389.200 97.800 ;
        RECT 401.200 97.600 402.000 98.400 ;
        RECT 404.500 92.400 405.100 103.600 ;
        RECT 404.400 91.600 405.200 92.400 ;
        RECT 401.200 89.600 402.000 90.400 ;
        RECT 398.000 83.600 398.800 84.400 ;
        RECT 378.800 81.600 379.600 82.400 ;
        RECT 398.000 81.600 398.800 82.400 ;
        RECT 398.100 78.400 398.700 81.600 ;
        RECT 398.000 77.600 398.800 78.400 ;
        RECT 386.800 73.600 387.600 74.400 ;
        RECT 390.000 73.600 390.800 74.400 ;
        RECT 386.900 72.400 387.500 73.600 ;
        RECT 370.800 71.600 371.600 72.400 ;
        RECT 374.000 71.600 374.800 72.400 ;
        RECT 382.000 71.600 382.800 72.400 ;
        RECT 386.800 71.600 387.600 72.400 ;
        RECT 393.200 71.600 394.000 72.400 ;
        RECT 394.800 71.600 395.600 72.400 ;
        RECT 396.200 71.800 397.000 72.600 ;
        RECT 401.300 72.400 401.900 89.600 ;
        RECT 406.100 84.400 406.700 109.700 ;
        RECT 407.600 107.600 408.400 108.400 ;
        RECT 407.700 96.400 408.300 107.600 ;
        RECT 410.800 104.200 411.600 115.800 ;
        RECT 407.600 95.600 408.400 96.400 ;
        RECT 407.600 93.600 408.400 94.400 ;
        RECT 412.500 92.400 413.100 139.600 ;
        RECT 414.000 135.600 414.800 136.400 ;
        RECT 414.100 134.400 414.700 135.600 ;
        RECT 414.000 133.600 414.800 134.400 ;
        RECT 415.600 123.600 416.400 124.400 ;
        RECT 415.700 110.400 416.300 123.600 ;
        RECT 422.100 118.400 422.700 181.700 ;
        RECT 423.600 177.600 424.400 178.400 ;
        RECT 423.700 172.400 424.300 177.600 ;
        RECT 423.600 171.600 424.400 172.400 ;
        RECT 425.200 171.600 426.000 172.400 ;
        RECT 423.700 150.400 424.300 171.600 ;
        RECT 423.600 149.600 424.400 150.400 ;
        RECT 425.300 120.400 425.900 171.600 ;
        RECT 426.800 170.200 427.600 175.800 ;
        RECT 428.500 158.300 429.100 227.600 ;
        RECT 434.900 224.400 435.500 251.600 ;
        RECT 436.500 240.400 437.100 253.600 ;
        RECT 441.300 250.400 441.900 255.600 ;
        RECT 444.500 254.400 445.100 269.600 ;
        RECT 449.300 268.400 449.900 303.600 ;
        RECT 450.800 299.600 451.600 300.400 ;
        RECT 450.900 296.400 451.500 299.600 ;
        RECT 457.300 296.400 457.900 303.600 ;
        RECT 458.900 296.400 459.500 315.600 ;
        RECT 450.800 295.600 451.600 296.400 ;
        RECT 457.200 295.600 458.000 296.400 ;
        RECT 458.800 295.600 459.600 296.400 ;
        RECT 450.800 293.600 451.600 294.400 ;
        RECT 460.500 290.400 461.100 317.600 ;
        RECT 465.300 316.400 465.900 333.600 ;
        RECT 468.500 330.400 469.100 333.600 ;
        RECT 471.600 331.600 472.400 332.400 ;
        RECT 478.000 331.600 478.800 332.400 ;
        RECT 481.200 331.600 482.000 332.400 ;
        RECT 468.400 329.600 469.200 330.400 ;
        RECT 470.000 329.600 470.800 330.400 ;
        RECT 466.800 327.600 467.600 328.400 ;
        RECT 465.200 315.600 466.000 316.400 ;
        RECT 466.800 309.600 467.600 310.400 ;
        RECT 465.200 307.600 466.000 308.400 ;
        RECT 463.600 293.600 464.400 294.400 ;
        RECT 462.000 291.600 462.800 292.400 ;
        RECT 460.400 289.600 461.200 290.400 ;
        RECT 452.400 287.600 453.200 288.400 ;
        RECT 463.600 287.600 464.400 288.400 ;
        RECT 452.500 278.400 453.100 287.600 ;
        RECT 465.300 284.400 465.900 307.600 ;
        RECT 470.100 300.400 470.700 329.600 ;
        RECT 471.700 326.400 472.300 331.600 ;
        RECT 478.100 330.400 478.700 331.600 ;
        RECT 478.000 329.600 478.800 330.400 ;
        RECT 471.600 325.600 472.400 326.400 ;
        RECT 471.700 312.400 472.300 325.600 ;
        RECT 474.800 323.600 475.600 324.400 ;
        RECT 474.900 312.400 475.500 323.600 ;
        RECT 478.100 314.400 478.700 329.600 ;
        RECT 481.300 318.400 481.900 331.600 ;
        RECT 482.900 330.400 483.500 333.600 ;
        RECT 484.500 332.400 485.100 333.600 ;
        RECT 484.400 331.600 485.200 332.400 ;
        RECT 482.800 329.600 483.600 330.400 ;
        RECT 487.600 329.600 488.400 330.400 ;
        RECT 487.700 326.400 488.300 329.600 ;
        RECT 487.600 325.600 488.400 326.400 ;
        RECT 486.000 323.600 486.800 324.400 ;
        RECT 481.200 317.600 482.000 318.400 ;
        RECT 478.000 313.600 478.800 314.400 ;
        RECT 481.200 313.600 482.000 314.400 ;
        RECT 484.400 313.600 485.200 314.400 ;
        RECT 481.300 312.400 481.900 313.600 ;
        RECT 471.600 311.600 472.400 312.400 ;
        RECT 474.800 311.600 475.600 312.400 ;
        RECT 479.600 311.600 480.400 312.400 ;
        RECT 481.200 311.600 482.000 312.400 ;
        RECT 484.500 310.400 485.100 313.600 ;
        RECT 486.100 312.400 486.700 323.600 ;
        RECT 487.600 315.600 488.400 316.400 ;
        RECT 487.700 312.400 488.300 315.600 ;
        RECT 486.000 311.600 486.800 312.400 ;
        RECT 487.600 311.600 488.400 312.400 ;
        RECT 471.600 309.600 472.400 310.400 ;
        RECT 476.400 309.600 477.200 310.400 ;
        RECT 484.400 309.600 485.200 310.400 ;
        RECT 486.000 307.600 486.800 308.400 ;
        RECT 471.600 305.600 472.400 306.400 ;
        RECT 479.600 305.600 480.400 306.400 ;
        RECT 471.700 300.400 472.300 305.600 ;
        RECT 481.200 303.600 482.000 304.400 ;
        RECT 486.100 302.400 486.700 307.600 ;
        RECT 487.600 303.600 488.400 304.400 ;
        RECT 476.400 301.600 477.200 302.400 ;
        RECT 486.000 301.600 486.800 302.400 ;
        RECT 470.000 299.600 470.800 300.400 ;
        RECT 471.600 299.600 472.400 300.400 ;
        RECT 466.800 295.600 467.600 296.400 ;
        RECT 466.900 290.400 467.500 295.600 ;
        RECT 468.400 291.600 469.200 292.400 ;
        RECT 466.800 289.600 467.600 290.400 ;
        RECT 466.800 287.600 467.600 288.400 ;
        RECT 463.600 283.600 464.400 284.400 ;
        RECT 465.200 283.600 466.000 284.400 ;
        RECT 452.400 277.600 453.200 278.400 ;
        RECT 450.800 273.600 451.600 274.400 ;
        RECT 455.600 273.600 456.400 274.400 ;
        RECT 450.900 270.400 451.500 273.600 ;
        RECT 454.000 271.600 454.800 272.400 ;
        RECT 454.100 270.400 454.700 271.600 ;
        RECT 450.800 269.600 451.600 270.400 ;
        RECT 454.000 269.600 454.800 270.400 ;
        RECT 446.000 267.600 446.800 268.400 ;
        RECT 449.200 267.600 450.000 268.400 ;
        RECT 444.400 253.600 445.200 254.400 ;
        RECT 439.600 249.600 440.400 250.400 ;
        RECT 441.200 249.600 442.000 250.400 ;
        RECT 436.400 239.600 437.200 240.400 ;
        RECT 434.800 223.600 435.600 224.400 ;
        RECT 441.300 220.400 441.900 249.600 ;
        RECT 444.500 226.400 445.100 253.600 ;
        RECT 446.100 250.300 446.700 267.600 ;
        RECT 447.600 253.600 448.400 254.400 ;
        RECT 447.700 252.400 448.300 253.600 ;
        RECT 447.600 251.600 448.400 252.400 ;
        RECT 449.300 250.300 449.900 267.600 ;
        RECT 450.900 256.400 451.500 269.600 ;
        RECT 454.000 259.600 454.800 260.400 ;
        RECT 450.800 255.600 451.600 256.400 ;
        RECT 454.100 254.400 454.700 259.600 ;
        RECT 455.700 258.400 456.300 273.600 ;
        RECT 463.700 272.400 464.300 283.600 ;
        RECT 465.200 277.600 466.000 278.400 ;
        RECT 463.600 271.600 464.400 272.400 ;
        RECT 465.300 270.400 465.900 277.600 ;
        RECT 466.900 276.400 467.500 287.600 ;
        RECT 468.500 278.400 469.100 291.600 ;
        RECT 471.700 286.400 472.300 299.600 ;
        RECT 476.500 298.400 477.100 301.600 ;
        RECT 476.400 297.600 477.200 298.400 ;
        RECT 478.000 295.600 478.800 296.400 ;
        RECT 473.200 293.600 474.000 294.400 ;
        RECT 474.800 293.600 475.600 294.400 ;
        RECT 473.300 292.400 473.900 293.600 ;
        RECT 478.100 292.400 478.700 295.600 ;
        RECT 479.600 293.600 480.400 294.400 ;
        RECT 482.800 293.600 483.600 294.400 ;
        RECT 486.000 293.600 486.800 294.400 ;
        RECT 473.200 291.600 474.000 292.400 ;
        RECT 478.000 291.600 478.800 292.400 ;
        RECT 484.400 291.600 485.200 292.400 ;
        RECT 479.600 289.600 480.400 290.400 ;
        RECT 471.600 285.600 472.400 286.400 ;
        RECT 471.600 283.600 472.400 284.400 ;
        RECT 468.400 277.600 469.200 278.400 ;
        RECT 466.800 275.600 467.600 276.400 ;
        RECT 466.900 274.400 467.500 275.600 ;
        RECT 466.800 273.600 467.600 274.400 ;
        RECT 470.000 274.300 470.800 274.400 ;
        RECT 468.500 273.700 470.800 274.300 ;
        RECT 465.200 269.600 466.000 270.400 ;
        RECT 463.600 261.600 464.400 262.400 ;
        RECT 455.600 257.600 456.400 258.400 ;
        RECT 452.400 253.600 453.200 254.400 ;
        RECT 454.000 253.600 454.800 254.400 ;
        RECT 455.600 253.600 456.400 254.400 ;
        RECT 457.200 253.600 458.000 254.400 ;
        RECT 452.400 251.600 453.200 252.400 ;
        RECT 455.700 250.400 456.300 253.600 ;
        RECT 458.800 251.600 459.600 252.400 ;
        RECT 446.100 249.700 448.300 250.300 ;
        RECT 449.300 249.700 451.500 250.300 ;
        RECT 447.700 246.400 448.300 249.700 ;
        RECT 449.200 247.600 450.000 248.400 ;
        RECT 447.600 245.600 448.400 246.400 ;
        RECT 446.000 229.600 446.800 230.400 ;
        RECT 444.400 225.600 445.200 226.400 ;
        RECT 446.100 224.400 446.700 229.600 ;
        RECT 447.700 228.400 448.300 245.600 ;
        RECT 449.300 230.400 449.900 247.600 ;
        RECT 450.900 234.300 451.500 249.700 ;
        RECT 452.400 249.600 453.200 250.400 ;
        RECT 455.600 249.600 456.400 250.400 ;
        RECT 452.500 246.400 453.100 249.600 ;
        RECT 452.400 245.600 453.200 246.400 ;
        RECT 463.700 242.400 464.300 261.600 ;
        RECT 465.200 259.600 466.000 260.400 ;
        RECT 465.300 254.400 465.900 259.600 ;
        RECT 468.500 258.400 469.100 273.700 ;
        RECT 470.000 273.600 470.800 273.700 ;
        RECT 471.700 272.400 472.300 283.600 ;
        RECT 479.700 282.400 480.300 289.600 ;
        RECT 481.200 283.600 482.000 284.400 ;
        RECT 479.600 281.600 480.400 282.400 ;
        RECT 474.800 279.600 475.600 280.400 ;
        RECT 474.900 278.400 475.500 279.600 ;
        RECT 474.800 277.600 475.600 278.400 ;
        RECT 474.800 275.600 475.600 276.400 ;
        RECT 478.000 275.600 478.800 276.400 ;
        RECT 471.600 271.600 472.400 272.400 ;
        RECT 474.900 270.400 475.500 275.600 ;
        RECT 478.100 272.400 478.700 275.600 ;
        RECT 479.600 273.600 480.400 274.400 ;
        RECT 476.400 271.600 477.200 272.400 ;
        RECT 478.000 271.600 478.800 272.400 ;
        RECT 471.600 269.600 472.400 270.400 ;
        RECT 474.800 269.600 475.600 270.400 ;
        RECT 471.700 262.400 472.300 269.600 ;
        RECT 471.600 261.600 472.400 262.400 ;
        RECT 466.800 257.600 467.600 258.400 ;
        RECT 468.400 257.600 469.200 258.400 ;
        RECT 471.600 257.600 472.400 258.400 ;
        RECT 465.200 253.600 466.000 254.400 ;
        RECT 465.200 251.600 466.000 252.400 ;
        RECT 465.300 250.400 465.900 251.600 ;
        RECT 465.200 249.600 466.000 250.400 ;
        RECT 466.900 248.400 467.500 257.600 ;
        RECT 470.000 253.600 470.800 254.400 ;
        RECT 471.700 252.400 472.300 257.600 ;
        RECT 474.900 252.400 475.500 269.600 ;
        RECT 476.500 268.400 477.100 271.600 ;
        RECT 478.000 269.600 478.800 270.400 ;
        RECT 476.400 267.600 477.200 268.400 ;
        RECT 479.700 266.400 480.300 273.600 ;
        RECT 476.400 265.600 477.200 266.400 ;
        RECT 479.600 265.600 480.400 266.400 ;
        RECT 471.600 251.600 472.400 252.400 ;
        RECT 474.800 251.600 475.600 252.400 ;
        RECT 473.200 249.600 474.000 250.400 ;
        RECT 465.200 247.600 466.000 248.400 ;
        RECT 466.800 247.600 467.600 248.400 ;
        RECT 463.600 241.600 464.400 242.400 ;
        RECT 454.000 239.600 454.800 240.400 ;
        RECT 450.900 233.700 453.100 234.300 ;
        RECT 450.800 231.600 451.600 232.400 ;
        RECT 449.200 229.600 450.000 230.400 ;
        RECT 450.900 228.400 451.500 231.600 ;
        RECT 452.500 230.400 453.100 233.700 ;
        RECT 454.100 230.400 454.700 239.600 ;
        RECT 463.600 237.600 464.400 238.400 ;
        RECT 462.000 234.300 462.800 234.400 ;
        RECT 457.300 233.700 462.800 234.300 ;
        RECT 457.300 230.400 457.900 233.700 ;
        RECT 462.000 233.600 462.800 233.700 ;
        RECT 452.400 229.600 453.200 230.400 ;
        RECT 454.000 229.600 454.800 230.400 ;
        RECT 457.200 229.600 458.000 230.400 ;
        RECT 460.400 229.600 461.200 230.400 ;
        RECT 447.600 227.600 448.400 228.400 ;
        RECT 450.800 227.600 451.600 228.400 ;
        RECT 455.600 227.600 456.400 228.400 ;
        RECT 458.800 227.600 459.600 228.400 ;
        RECT 442.800 223.600 443.600 224.400 ;
        RECT 446.000 223.600 446.800 224.400 ;
        RECT 441.200 219.600 442.000 220.400 ;
        RECT 434.800 211.600 435.600 212.400 ;
        RECT 433.200 199.600 434.000 200.400 ;
        RECT 431.600 183.600 432.400 184.400 ;
        RECT 430.000 166.200 430.800 177.800 ;
        RECT 431.700 172.400 432.300 183.600 ;
        RECT 433.300 174.400 433.900 199.600 ;
        RECT 434.900 188.400 435.500 211.600 ;
        RECT 436.400 204.200 437.200 217.800 ;
        RECT 438.000 204.200 438.800 217.800 ;
        RECT 439.600 204.200 440.400 217.800 ;
        RECT 441.200 206.200 442.000 217.800 ;
        RECT 442.900 216.400 443.500 223.600 ;
        RECT 442.800 215.600 443.600 216.400 ;
        RECT 442.900 200.400 443.500 215.600 ;
        RECT 444.400 206.200 445.200 217.800 ;
        RECT 446.000 213.600 446.800 214.400 ;
        RECT 447.600 206.200 448.400 217.800 ;
        RECT 449.200 204.200 450.000 217.800 ;
        RECT 450.800 204.200 451.600 217.800 ;
        RECT 455.700 216.400 456.300 227.600 ;
        RECT 458.900 224.400 459.500 227.600 ;
        RECT 458.800 223.600 459.600 224.400 ;
        RECT 460.500 220.400 461.100 229.600 ;
        RECT 463.700 220.400 464.300 237.600 ;
        RECT 460.400 219.600 461.200 220.400 ;
        RECT 463.600 219.600 464.400 220.400 ;
        RECT 465.300 216.400 465.900 247.600 ;
        RECT 473.300 238.400 473.900 249.600 ;
        RECT 474.900 240.400 475.500 251.600 ;
        RECT 476.500 248.400 477.100 265.600 ;
        RECT 478.000 261.600 478.800 262.400 ;
        RECT 478.100 258.400 478.700 261.600 ;
        RECT 481.300 258.400 481.900 283.600 ;
        RECT 482.800 273.600 483.600 274.400 ;
        RECT 482.800 271.600 483.600 272.400 ;
        RECT 482.900 270.400 483.500 271.600 ;
        RECT 482.800 269.600 483.600 270.400 ;
        RECT 478.000 257.600 478.800 258.400 ;
        RECT 481.200 257.600 482.000 258.400 ;
        RECT 482.900 256.400 483.500 269.600 ;
        RECT 484.500 266.400 485.100 291.600 ;
        RECT 486.100 270.400 486.700 293.600 ;
        RECT 487.700 282.400 488.300 303.600 ;
        RECT 489.300 300.400 489.900 333.600 ;
        RECT 495.600 331.600 496.400 332.400 ;
        RECT 500.400 331.600 501.200 332.400 ;
        RECT 494.000 329.600 494.800 330.400 ;
        RECT 494.100 328.400 494.700 329.600 ;
        RECT 494.000 327.600 494.800 328.400 ;
        RECT 495.600 327.600 496.400 328.400 ;
        RECT 490.800 323.600 491.600 324.400 ;
        RECT 490.900 322.400 491.500 323.600 ;
        RECT 490.800 321.600 491.600 322.400 ;
        RECT 490.800 317.600 491.600 318.400 ;
        RECT 490.900 308.400 491.500 317.600 ;
        RECT 495.700 310.400 496.300 327.600 ;
        RECT 498.800 323.600 499.600 324.400 ;
        RECT 498.900 312.300 499.500 323.600 ;
        RECT 500.500 316.400 501.100 331.600 ;
        RECT 505.300 330.400 505.900 335.600 ;
        RECT 510.000 331.600 510.800 332.400 ;
        RECT 505.200 329.600 506.000 330.400 ;
        RECT 502.000 323.600 502.800 324.400 ;
        RECT 502.100 318.400 502.700 323.600 ;
        RECT 502.000 317.600 502.800 318.400 ;
        RECT 505.300 318.300 505.900 329.600 ;
        RECT 506.800 323.600 507.600 324.400 ;
        RECT 506.900 320.400 507.500 323.600 ;
        RECT 506.800 319.600 507.600 320.400 ;
        RECT 505.300 317.700 507.500 318.300 ;
        RECT 500.400 315.600 501.200 316.400 ;
        RECT 502.000 313.600 502.800 314.400 ;
        RECT 497.300 311.700 499.500 312.300 ;
        RECT 495.600 309.600 496.400 310.400 ;
        RECT 497.300 308.400 497.900 311.700 ;
        RECT 505.200 311.600 506.000 312.400 ;
        RECT 505.300 310.400 505.900 311.600 ;
        RECT 498.800 309.600 499.600 310.400 ;
        RECT 500.400 309.600 501.200 310.400 ;
        RECT 502.000 309.600 502.800 310.400 ;
        RECT 505.200 309.600 506.000 310.400 ;
        RECT 490.800 307.600 491.600 308.400 ;
        RECT 492.400 307.600 493.200 308.400 ;
        RECT 497.200 307.600 498.000 308.400 ;
        RECT 492.500 306.400 493.100 307.600 ;
        RECT 492.400 305.600 493.200 306.400 ;
        RECT 494.000 305.600 494.800 306.400 ;
        RECT 489.200 299.600 490.000 300.400 ;
        RECT 494.100 298.400 494.700 305.600 ;
        RECT 497.200 301.600 498.000 302.400 ;
        RECT 497.300 298.400 497.900 301.600 ;
        RECT 489.200 297.600 490.000 298.400 ;
        RECT 494.000 297.600 494.800 298.400 ;
        RECT 497.200 297.600 498.000 298.400 ;
        RECT 489.300 296.400 489.900 297.600 ;
        RECT 489.200 295.600 490.000 296.400 ;
        RECT 490.800 296.300 491.600 296.400 ;
        RECT 490.800 295.700 493.100 296.300 ;
        RECT 490.800 295.600 491.600 295.700 ;
        RECT 489.200 293.600 490.000 294.400 ;
        RECT 490.800 293.600 491.600 294.400 ;
        RECT 489.300 292.400 489.900 293.600 ;
        RECT 489.200 291.600 490.000 292.400 ;
        RECT 487.600 281.600 488.400 282.400 ;
        RECT 490.900 280.400 491.500 293.600 ;
        RECT 492.500 292.400 493.100 295.700 ;
        RECT 495.600 293.600 496.400 294.400 ;
        RECT 498.900 292.400 499.500 309.600 ;
        RECT 500.400 307.600 501.200 308.400 ;
        RECT 502.100 306.300 502.700 309.600 ;
        RECT 506.900 308.400 507.500 317.700 ;
        RECT 508.400 313.600 509.200 314.400 ;
        RECT 508.400 309.600 509.200 310.400 ;
        RECT 506.800 307.600 507.600 308.400 ;
        RECT 508.500 308.300 509.100 309.600 ;
        RECT 510.100 308.300 510.700 331.600 ;
        RECT 516.400 324.200 517.200 337.800 ;
        RECT 518.000 324.200 518.800 337.800 ;
        RECT 519.600 324.200 520.400 337.800 ;
        RECT 521.200 326.200 522.000 337.800 ;
        RECT 522.900 336.400 523.500 345.600 ;
        RECT 526.000 343.600 526.800 344.400 ;
        RECT 530.800 343.600 531.600 344.400 ;
        RECT 526.100 342.400 526.700 343.600 ;
        RECT 526.000 341.600 526.800 342.400 ;
        RECT 530.900 340.400 531.500 343.600 ;
        RECT 526.000 339.600 526.800 340.400 ;
        RECT 530.800 339.600 531.600 340.400 ;
        RECT 522.800 335.600 523.600 336.400 ;
        RECT 524.400 326.200 525.200 337.800 ;
        RECT 526.100 334.400 526.700 339.600 ;
        RECT 526.000 333.600 526.800 334.400 ;
        RECT 526.000 331.600 526.800 332.400 ;
        RECT 518.000 321.600 518.800 322.400 ;
        RECT 524.400 321.600 525.200 322.400 ;
        RECT 513.200 317.600 514.000 318.400 ;
        RECT 513.300 312.400 513.900 317.600 ;
        RECT 518.100 312.400 518.700 321.600 ;
        RECT 521.200 319.600 522.000 320.400 ;
        RECT 521.300 314.400 521.900 319.600 ;
        RECT 522.800 317.600 523.600 318.400 ;
        RECT 521.200 313.600 522.000 314.400 ;
        RECT 511.600 311.600 512.400 312.400 ;
        RECT 513.200 311.600 514.000 312.400 ;
        RECT 518.000 311.600 518.800 312.400 ;
        RECT 521.200 311.600 522.000 312.400 ;
        RECT 511.600 309.600 512.400 310.400 ;
        RECT 521.300 308.400 521.900 311.600 ;
        RECT 508.500 307.700 510.700 308.300 ;
        RECT 500.500 305.700 502.700 306.300 ;
        RECT 500.500 296.400 501.100 305.700 ;
        RECT 502.000 299.600 502.800 300.400 ;
        RECT 500.400 295.600 501.200 296.400 ;
        RECT 492.400 291.600 493.200 292.400 ;
        RECT 494.000 291.600 494.800 292.400 ;
        RECT 498.800 291.600 499.600 292.400 ;
        RECT 490.800 279.600 491.600 280.400 ;
        RECT 492.500 278.400 493.100 291.600 ;
        RECT 495.600 289.600 496.400 290.400 ;
        RECT 498.800 289.600 499.600 290.400 ;
        RECT 500.400 289.600 501.200 290.400 ;
        RECT 495.700 288.400 496.300 289.600 ;
        RECT 495.600 287.600 496.400 288.400 ;
        RECT 497.200 281.600 498.000 282.400 ;
        RECT 492.400 277.600 493.200 278.400 ;
        RECT 487.600 275.600 488.400 276.400 ;
        RECT 486.000 269.600 486.800 270.400 ;
        RECT 487.700 268.400 488.300 275.600 ;
        RECT 489.200 273.600 490.000 274.400 ;
        RECT 489.300 270.400 489.900 273.600 ;
        RECT 489.200 269.600 490.000 270.400 ;
        RECT 492.400 270.300 493.200 270.400 ;
        RECT 490.900 269.700 493.200 270.300 ;
        RECT 486.000 267.600 486.800 268.400 ;
        RECT 487.600 267.600 488.400 268.400 ;
        RECT 486.100 266.400 486.700 267.600 ;
        RECT 484.400 265.600 485.200 266.400 ;
        RECT 486.000 265.600 486.800 266.400 ;
        RECT 484.400 263.600 485.200 264.400 ;
        RECT 484.500 262.400 485.100 263.600 ;
        RECT 484.400 261.600 485.200 262.400 ;
        RECT 479.600 255.600 480.400 256.400 ;
        RECT 482.800 255.600 483.600 256.400 ;
        RECT 486.100 256.300 486.700 265.600 ;
        RECT 490.900 256.400 491.500 269.700 ;
        RECT 492.400 269.600 493.200 269.700 ;
        RECT 495.600 269.600 496.400 270.400 ;
        RECT 497.300 270.300 497.900 281.600 ;
        RECT 498.900 276.300 499.500 289.600 ;
        RECT 500.500 286.400 501.100 289.600 ;
        RECT 500.400 285.600 501.200 286.400 ;
        RECT 500.500 278.400 501.100 285.600 ;
        RECT 500.400 277.600 501.200 278.400 ;
        RECT 500.400 276.300 501.200 276.400 ;
        RECT 498.900 275.700 501.200 276.300 ;
        RECT 500.400 275.600 501.200 275.700 ;
        RECT 502.100 272.400 502.700 299.600 ;
        RECT 506.900 296.400 507.500 307.600 ;
        RECT 506.800 295.600 507.600 296.400 ;
        RECT 506.800 293.600 507.600 294.400 ;
        RECT 506.900 282.400 507.500 293.600 ;
        RECT 508.400 291.600 509.200 292.400 ;
        RECT 506.800 281.600 507.600 282.400 ;
        RECT 505.200 279.600 506.000 280.400 ;
        RECT 505.300 278.400 505.900 279.600 ;
        RECT 505.200 277.600 506.000 278.400 ;
        RECT 502.000 271.600 502.800 272.400 ;
        RECT 506.800 271.600 507.600 272.400 ;
        RECT 497.300 269.700 499.500 270.300 ;
        RECT 494.000 267.600 494.800 268.400 ;
        RECT 494.100 264.400 494.700 267.600 ;
        RECT 495.700 266.400 496.300 269.600 ;
        RECT 497.200 267.600 498.000 268.400 ;
        RECT 495.600 265.600 496.400 266.400 ;
        RECT 494.000 263.600 494.800 264.400 ;
        RECT 492.400 257.600 493.200 258.400 ;
        RECT 494.100 256.400 494.700 263.600 ;
        RECT 495.600 261.600 496.400 262.400 ;
        RECT 487.600 256.300 488.400 256.400 ;
        RECT 486.100 255.700 488.400 256.300 ;
        RECT 482.800 251.600 483.600 252.400 ;
        RECT 484.400 251.600 485.200 252.400 ;
        RECT 482.900 250.400 483.500 251.600 ;
        RECT 482.800 249.600 483.600 250.400 ;
        RECT 476.400 247.600 477.200 248.400 ;
        RECT 481.200 243.600 482.000 244.400 ;
        RECT 481.300 242.400 481.900 243.600 ;
        RECT 482.900 242.400 483.500 249.600 ;
        RECT 484.400 245.600 485.200 246.400 ;
        RECT 484.500 244.400 485.100 245.600 ;
        RECT 484.400 243.600 485.200 244.400 ;
        RECT 481.200 241.600 482.000 242.400 ;
        RECT 482.800 241.600 483.600 242.400 ;
        RECT 474.800 239.600 475.600 240.400 ;
        RECT 473.200 237.600 474.000 238.400 ;
        RECT 466.800 234.300 467.600 234.400 ;
        RECT 466.800 233.700 472.300 234.300 ;
        RECT 466.800 233.600 467.600 233.700 ;
        RECT 471.700 232.400 472.300 233.700 ;
        RECT 474.800 233.600 475.600 234.400 ;
        RECT 476.400 233.600 477.200 234.400 ;
        RECT 474.900 232.400 475.500 233.600 ;
        RECT 470.000 231.600 470.800 232.400 ;
        RECT 471.600 231.600 472.400 232.400 ;
        RECT 474.800 231.600 475.600 232.400 ;
        RECT 470.000 230.300 470.800 230.400 ;
        RECT 473.200 230.300 474.000 230.400 ;
        RECT 470.000 229.700 474.000 230.300 ;
        RECT 470.000 229.600 470.800 229.700 ;
        RECT 473.200 229.600 474.000 229.700 ;
        RECT 466.800 227.600 467.600 228.400 ;
        RECT 471.600 227.600 472.400 228.400 ;
        RECT 466.900 226.400 467.500 227.600 ;
        RECT 466.800 225.600 467.600 226.400 ;
        RECT 468.400 223.600 469.200 224.400 ;
        RECT 468.500 216.400 469.100 223.600 ;
        RECT 471.700 216.400 472.300 227.600 ;
        RECT 476.500 226.300 477.100 233.600 ;
        RECT 484.500 232.400 485.100 243.600 ;
        RECT 478.000 231.600 478.800 232.400 ;
        RECT 481.200 231.600 482.000 232.400 ;
        RECT 484.400 231.600 485.200 232.400 ;
        RECT 478.000 229.600 478.800 230.400 ;
        RECT 482.800 229.600 483.600 230.400 ;
        RECT 478.100 228.400 478.700 229.600 ;
        RECT 482.900 228.400 483.500 229.600 ;
        RECT 478.000 227.600 478.800 228.400 ;
        RECT 481.200 227.600 482.000 228.400 ;
        RECT 482.800 227.600 483.600 228.400 ;
        RECT 476.500 225.700 478.700 226.300 ;
        RECT 474.800 219.600 475.600 220.400 ;
        RECT 474.900 216.400 475.500 219.600 ;
        RECT 478.100 216.400 478.700 225.700 ;
        RECT 481.300 218.400 481.900 227.600 ;
        RECT 482.900 218.400 483.500 227.600 ;
        RECT 481.200 217.600 482.000 218.400 ;
        RECT 482.800 217.600 483.600 218.400 ;
        RECT 481.300 216.400 481.900 217.600 ;
        RECT 455.600 215.600 456.400 216.400 ;
        RECT 465.200 215.600 466.000 216.400 ;
        RECT 468.400 215.600 469.200 216.400 ;
        RECT 471.600 215.600 472.400 216.400 ;
        RECT 474.800 215.600 475.600 216.400 ;
        RECT 478.000 215.600 478.800 216.400 ;
        RECT 481.200 215.600 482.000 216.400 ;
        RECT 486.100 214.400 486.700 255.700 ;
        RECT 487.600 255.600 488.400 255.700 ;
        RECT 489.200 255.600 490.000 256.400 ;
        RECT 490.800 255.600 491.600 256.400 ;
        RECT 494.000 255.600 494.800 256.400 ;
        RECT 489.200 253.600 490.000 254.400 ;
        RECT 487.600 233.600 488.400 234.400 ;
        RECT 487.600 231.600 488.400 232.400 ;
        RECT 487.700 228.400 488.300 231.600 ;
        RECT 489.300 230.400 489.900 253.600 ;
        RECT 490.900 244.400 491.500 255.600 ;
        RECT 495.700 252.400 496.300 261.600 ;
        RECT 497.200 253.600 498.000 254.400 ;
        RECT 495.600 251.600 496.400 252.400 ;
        RECT 495.700 250.400 496.300 251.600 ;
        RECT 495.600 249.600 496.400 250.400 ;
        RECT 490.800 243.600 491.600 244.400 ;
        RECT 490.800 239.600 491.600 240.400 ;
        RECT 490.900 238.400 491.500 239.600 ;
        RECT 490.800 237.600 491.600 238.400 ;
        RECT 495.600 237.600 496.400 238.400 ;
        RECT 492.400 233.600 493.200 234.400 ;
        RECT 495.700 232.400 496.300 237.600 ;
        RECT 495.600 231.600 496.400 232.400 ;
        RECT 489.200 229.600 490.000 230.400 ;
        RECT 494.000 229.600 494.800 230.400 ;
        RECT 497.200 229.600 498.000 230.400 ;
        RECT 487.600 227.600 488.400 228.400 ;
        RECT 497.200 225.600 498.000 226.400 ;
        RECT 497.300 220.400 497.900 225.600 ;
        RECT 497.200 219.600 498.000 220.400 ;
        RECT 498.900 220.300 499.500 269.700 ;
        RECT 503.600 269.600 504.400 270.400 ;
        RECT 505.200 269.600 506.000 270.400 ;
        RECT 500.400 265.600 501.200 266.400 ;
        RECT 502.000 265.600 502.800 266.400 ;
        RECT 500.500 260.400 501.100 265.600 ;
        RECT 502.100 264.400 502.700 265.600 ;
        RECT 502.000 263.600 502.800 264.400 ;
        RECT 502.100 262.400 502.700 263.600 ;
        RECT 502.000 261.600 502.800 262.400 ;
        RECT 503.700 260.400 504.300 269.600 ;
        RECT 505.300 264.400 505.900 269.600 ;
        RECT 505.200 263.600 506.000 264.400 ;
        RECT 500.400 259.600 501.200 260.400 ;
        RECT 503.600 259.600 504.400 260.400 ;
        RECT 506.900 258.400 507.500 271.600 ;
        RECT 508.500 270.400 509.100 291.600 ;
        RECT 510.100 274.400 510.700 307.700 ;
        RECT 516.400 307.600 517.200 308.400 ;
        RECT 521.200 307.600 522.000 308.400 ;
        RECT 511.600 305.600 512.400 306.400 ;
        RECT 511.700 298.400 512.300 305.600 ;
        RECT 518.000 303.600 518.800 304.400 ;
        RECT 511.600 297.600 512.400 298.400 ;
        RECT 518.100 294.400 518.700 303.600 ;
        RECT 521.300 302.400 521.900 307.600 ;
        RECT 521.200 301.600 522.000 302.400 ;
        RECT 521.200 297.600 522.000 298.400 ;
        RECT 521.300 296.400 521.900 297.600 ;
        RECT 522.900 296.400 523.500 317.600 ;
        RECT 521.200 295.600 522.000 296.400 ;
        RECT 522.800 295.600 523.600 296.400 ;
        RECT 513.200 294.300 514.000 294.400 ;
        RECT 511.700 293.700 514.000 294.300 ;
        RECT 510.000 273.600 510.800 274.400 ;
        RECT 511.700 270.400 512.300 293.700 ;
        RECT 513.200 293.600 514.000 293.700 ;
        RECT 518.000 293.600 518.800 294.400 ;
        RECT 521.300 292.400 521.900 295.600 ;
        RECT 518.000 291.600 518.800 292.400 ;
        RECT 521.200 291.600 522.000 292.400 ;
        RECT 518.100 290.400 518.700 291.600 ;
        RECT 516.400 289.600 517.200 290.400 ;
        RECT 518.000 289.600 518.800 290.400 ;
        RECT 513.200 281.600 514.000 282.400 ;
        RECT 508.400 269.600 509.200 270.400 ;
        RECT 511.600 269.600 512.400 270.400 ;
        RECT 511.600 267.600 512.400 268.400 ;
        RECT 508.400 263.600 509.200 264.400 ;
        RECT 502.000 257.600 502.800 258.400 ;
        RECT 506.800 257.600 507.600 258.400 ;
        RECT 500.400 255.600 501.200 256.400 ;
        RECT 500.500 246.400 501.100 255.600 ;
        RECT 502.100 254.400 502.700 257.600 ;
        RECT 505.200 255.600 506.000 256.400 ;
        RECT 505.300 254.400 505.900 255.600 ;
        RECT 502.000 253.600 502.800 254.400 ;
        RECT 505.200 253.600 506.000 254.400 ;
        RECT 508.500 252.400 509.100 263.600 ;
        RECT 511.700 258.400 512.300 267.600 ;
        RECT 513.300 266.400 513.900 281.600 ;
        RECT 516.500 274.400 517.100 289.600 ;
        RECT 521.200 285.600 522.000 286.400 ;
        RECT 519.600 283.600 520.400 284.400 ;
        RECT 519.700 278.400 520.300 283.600 ;
        RECT 519.600 277.600 520.400 278.400 ;
        RECT 516.400 273.600 517.200 274.400 ;
        RECT 516.400 269.600 517.200 270.400 ;
        RECT 516.500 266.400 517.100 269.600 ;
        RECT 521.300 266.400 521.900 285.600 ;
        RECT 522.800 279.600 523.600 280.400 ;
        RECT 522.900 268.400 523.500 279.600 ;
        RECT 524.500 278.400 525.100 321.600 ;
        RECT 526.100 318.400 526.700 331.600 ;
        RECT 527.600 326.200 528.400 337.800 ;
        RECT 529.200 324.200 530.000 337.800 ;
        RECT 530.800 324.200 531.600 337.800 ;
        RECT 526.000 317.600 526.800 318.400 ;
        RECT 527.600 313.600 528.400 314.400 ;
        RECT 532.400 313.600 533.200 314.400 ;
        RECT 526.000 309.600 526.800 310.400 ;
        RECT 526.100 304.400 526.700 309.600 ;
        RECT 527.700 308.400 528.300 313.600 ;
        RECT 529.200 311.600 530.000 312.400 ;
        RECT 529.300 310.400 529.900 311.600 ;
        RECT 534.100 310.400 534.700 353.600 ;
        RECT 535.600 343.600 536.400 344.400 ;
        RECT 535.700 332.400 536.300 343.600 ;
        RECT 537.300 336.400 537.900 375.600 ;
        RECT 538.800 366.200 539.600 377.800 ;
        RECT 540.400 373.600 541.200 374.400 ;
        RECT 542.000 366.200 542.800 377.800 ;
        RECT 543.600 364.200 544.400 377.800 ;
        RECT 545.200 364.200 546.000 377.800 ;
        RECT 546.900 370.800 547.500 379.600 ;
        RECT 554.900 374.400 555.500 383.600 ;
        RECT 554.800 373.600 555.600 374.400 ;
        RECT 558.000 373.600 558.800 374.400 ;
        RECT 558.100 372.400 558.700 373.600 ;
        RECT 554.800 371.600 555.600 372.400 ;
        RECT 558.000 371.600 558.800 372.400 ;
        RECT 546.800 370.000 547.600 370.800 ;
        RECT 554.900 366.400 555.500 371.600 ;
        RECT 551.600 365.600 552.400 366.400 ;
        RECT 554.800 365.600 555.600 366.400 ;
        RECT 551.700 358.400 552.300 365.600 ;
        RECT 554.800 359.600 555.600 360.400 ;
        RECT 542.000 357.600 542.800 358.400 ;
        RECT 551.600 357.600 552.400 358.400 ;
        RECT 538.800 355.600 539.600 356.400 ;
        RECT 538.900 350.400 539.500 355.600 ;
        RECT 540.400 351.600 541.200 352.400 ;
        RECT 540.500 350.400 541.100 351.600 ;
        RECT 538.800 349.600 539.600 350.400 ;
        RECT 540.400 349.600 541.200 350.400 ;
        RECT 537.200 335.600 538.000 336.400 ;
        RECT 537.200 333.600 538.000 334.400 ;
        RECT 535.600 331.600 536.400 332.400 ;
        RECT 537.300 312.400 537.900 333.600 ;
        RECT 537.200 311.600 538.000 312.400 ;
        RECT 538.800 312.300 539.600 312.400 ;
        RECT 540.500 312.300 541.100 349.600 ;
        RECT 538.800 311.700 541.100 312.300 ;
        RECT 538.800 311.600 539.600 311.700 ;
        RECT 538.900 310.400 539.500 311.600 ;
        RECT 529.200 309.600 530.000 310.400 ;
        RECT 534.000 309.600 534.800 310.400 ;
        RECT 538.800 309.600 539.600 310.400 ;
        RECT 527.600 307.600 528.400 308.400 ;
        RECT 529.200 307.600 530.000 308.400 ;
        RECT 534.000 308.300 534.800 308.400 ;
        RECT 532.500 307.700 534.800 308.300 ;
        RECT 526.000 303.600 526.800 304.400 ;
        RECT 526.000 301.600 526.800 302.400 ;
        RECT 526.100 294.400 526.700 301.600 ;
        RECT 526.000 293.600 526.800 294.400 ;
        RECT 526.000 291.600 526.800 292.400 ;
        RECT 526.000 283.600 526.800 284.400 ;
        RECT 524.400 277.600 525.200 278.400 ;
        RECT 526.100 272.300 526.700 283.600 ;
        RECT 527.700 276.400 528.300 307.600 ;
        RECT 529.300 298.400 529.900 307.600 ;
        RECT 529.200 297.600 530.000 298.400 ;
        RECT 532.500 294.400 533.100 307.700 ;
        RECT 534.000 307.600 534.800 307.700 ;
        RECT 542.100 306.400 542.700 357.600 ;
        RECT 551.700 356.400 552.300 357.600 ;
        RECT 551.600 355.600 552.400 356.400 ;
        RECT 554.900 352.400 555.500 359.600 ;
        RECT 559.700 354.400 560.300 387.600 ;
        RECT 566.100 386.400 566.700 391.600 ;
        RECT 572.500 390.400 573.100 403.600 ;
        RECT 572.400 389.600 573.200 390.400 ;
        RECT 567.600 387.600 568.400 388.400 ;
        RECT 570.800 387.600 571.600 388.400 ;
        RECT 572.400 387.600 573.200 388.400 ;
        RECT 561.200 385.600 562.000 386.400 ;
        RECT 566.000 385.600 566.800 386.400 ;
        RECT 561.300 370.400 561.900 385.600 ;
        RECT 566.000 383.600 566.800 384.400 ;
        RECT 562.800 375.600 563.600 376.400 ;
        RECT 566.100 374.400 566.700 383.600 ;
        RECT 564.400 373.600 565.200 374.400 ;
        RECT 566.000 373.600 566.800 374.400 ;
        RECT 561.200 369.600 562.000 370.400 ;
        RECT 559.600 353.600 560.400 354.400 ;
        RECT 554.800 351.600 555.600 352.400 ;
        RECT 558.000 351.600 558.800 352.400 ;
        RECT 558.100 348.400 558.700 351.600 ;
        RECT 559.700 350.400 560.300 353.600 ;
        RECT 561.200 351.600 562.000 352.400 ;
        RECT 564.400 351.600 565.200 352.400 ;
        RECT 559.600 349.600 560.400 350.400 ;
        RECT 543.600 347.600 544.400 348.400 ;
        RECT 558.000 347.600 558.800 348.400 ;
        RECT 559.600 347.600 560.400 348.400 ;
        RECT 554.800 343.600 555.600 344.400 ;
        RECT 554.900 340.300 555.500 343.600 ;
        RECT 553.300 339.700 555.500 340.300 ;
        RECT 543.600 331.600 544.400 332.400 ;
        RECT 546.800 323.600 547.600 324.400 ;
        RECT 548.400 324.200 549.200 337.800 ;
        RECT 550.000 324.200 550.800 337.800 ;
        RECT 551.600 326.200 552.400 337.800 ;
        RECT 553.300 334.400 553.900 339.700 ;
        RECT 564.500 338.400 565.100 351.600 ;
        RECT 566.100 348.400 566.700 373.600 ;
        RECT 567.700 372.400 568.300 387.600 ;
        RECT 570.900 384.400 571.500 387.600 ;
        RECT 572.500 386.400 573.100 387.600 ;
        RECT 572.400 385.600 573.200 386.400 ;
        RECT 570.800 383.600 571.600 384.400 ;
        RECT 569.200 373.600 570.000 374.400 ;
        RECT 567.600 371.600 568.400 372.400 ;
        RECT 570.800 367.600 571.600 368.400 ;
        RECT 567.600 349.600 568.400 350.400 ;
        RECT 566.000 347.600 566.800 348.400 ;
        RECT 553.200 333.600 554.000 334.400 ;
        RECT 554.800 326.200 555.600 337.800 ;
        RECT 556.400 335.600 557.200 336.400 ;
        RECT 558.000 326.200 558.800 337.800 ;
        RECT 559.600 324.200 560.400 337.800 ;
        RECT 561.200 324.200 562.000 337.800 ;
        RECT 562.800 324.200 563.600 337.800 ;
        RECT 564.400 337.600 565.200 338.400 ;
        RECT 570.900 334.400 571.500 367.600 ;
        RECT 574.100 362.400 574.700 409.600 ;
        RECT 575.700 390.400 576.300 415.700 ;
        RECT 582.000 415.600 582.800 416.400 ;
        RECT 578.800 411.600 579.600 412.400 ;
        RECT 575.600 389.600 576.400 390.400 ;
        RECT 577.200 389.600 578.000 390.400 ;
        RECT 577.300 372.400 577.900 389.600 ;
        RECT 577.200 371.600 578.000 372.400 ;
        RECT 574.000 361.600 574.800 362.400 ;
        RECT 574.000 344.200 574.800 357.800 ;
        RECT 575.600 344.200 576.400 357.800 ;
        RECT 577.200 344.200 578.000 355.800 ;
        RECT 578.900 350.400 579.500 411.600 ;
        RECT 583.600 404.200 584.400 417.800 ;
        RECT 585.200 404.200 586.000 417.800 ;
        RECT 586.800 406.200 587.600 417.800 ;
        RECT 588.400 413.600 589.200 414.400 ;
        RECT 590.000 406.200 590.800 417.800 ;
        RECT 591.600 415.600 592.400 416.400 ;
        RECT 591.700 398.300 592.300 415.600 ;
        RECT 593.200 406.200 594.000 417.800 ;
        RECT 594.800 404.200 595.600 417.800 ;
        RECT 596.400 404.200 597.200 417.800 ;
        RECT 598.000 404.200 598.800 417.800 ;
        RECT 599.700 412.400 600.300 441.600 ;
        RECT 612.500 428.400 613.100 533.600 ;
        RECT 612.400 427.600 613.200 428.400 ;
        RECT 601.200 423.600 602.000 424.400 ;
        RECT 601.300 416.400 601.900 423.600 ;
        RECT 601.200 415.600 602.000 416.400 ;
        RECT 599.600 411.600 600.400 412.400 ;
        RECT 607.600 403.600 608.400 404.400 ;
        RECT 604.400 399.600 605.200 400.400 ;
        RECT 606.000 399.600 606.800 400.400 ;
        RECT 582.000 384.200 582.800 397.800 ;
        RECT 583.600 384.200 584.400 397.800 ;
        RECT 590.100 397.700 592.300 398.300 ;
        RECT 585.200 384.200 586.000 395.800 ;
        RECT 586.800 389.600 587.600 390.400 ;
        RECT 586.900 388.400 587.500 389.600 ;
        RECT 586.800 387.600 587.600 388.400 ;
        RECT 588.400 384.200 589.200 395.800 ;
        RECT 590.100 386.400 590.700 397.700 ;
        RECT 590.000 385.600 590.800 386.400 ;
        RECT 582.000 371.600 582.800 372.400 ;
        RECT 583.600 364.200 584.400 377.800 ;
        RECT 585.200 364.200 586.000 377.800 ;
        RECT 586.800 364.200 587.600 377.800 ;
        RECT 588.400 366.200 589.200 377.800 ;
        RECT 590.100 376.400 590.700 385.600 ;
        RECT 591.600 384.200 592.400 395.800 ;
        RECT 593.200 384.200 594.000 397.800 ;
        RECT 594.800 384.200 595.600 397.800 ;
        RECT 596.400 384.200 597.200 397.800 ;
        RECT 590.000 375.600 590.800 376.400 ;
        RECT 591.600 366.200 592.400 377.800 ;
        RECT 593.200 375.600 594.000 376.400 ;
        RECT 593.300 374.400 593.900 375.600 ;
        RECT 593.200 373.600 594.000 374.400 ;
        RECT 593.200 371.600 594.000 372.400 ;
        RECT 578.800 349.600 579.600 350.400 ;
        RECT 578.800 347.600 579.600 348.400 ;
        RECT 578.900 342.300 579.500 347.600 ;
        RECT 580.400 344.200 581.200 355.800 ;
        RECT 582.000 345.600 582.800 346.400 ;
        RECT 578.900 341.700 581.100 342.300 ;
        RECT 580.500 338.400 581.100 341.700 ;
        RECT 572.400 337.600 573.200 338.400 ;
        RECT 580.400 337.600 581.200 338.400 ;
        RECT 570.800 333.600 571.600 334.400 ;
        RECT 578.800 333.600 579.600 334.400 ;
        RECT 578.900 332.400 579.500 333.600 ;
        RECT 578.800 331.600 579.600 332.400 ;
        RECT 582.100 330.300 582.700 345.600 ;
        RECT 583.600 344.200 584.400 355.800 ;
        RECT 585.200 344.200 586.000 357.800 ;
        RECT 586.800 344.200 587.600 357.800 ;
        RECT 588.400 344.200 589.200 357.800 ;
        RECT 590.000 349.600 590.800 350.400 ;
        RECT 590.100 348.400 590.700 349.600 ;
        RECT 590.000 347.600 590.800 348.400 ;
        RECT 585.200 341.600 586.000 342.400 ;
        RECT 585.300 334.400 585.900 341.600 ;
        RECT 588.400 335.600 589.200 336.400 ;
        RECT 593.300 334.400 593.900 371.600 ;
        RECT 594.800 366.200 595.600 377.800 ;
        RECT 596.400 364.200 597.200 377.800 ;
        RECT 598.000 364.200 598.800 377.800 ;
        RECT 604.500 352.400 605.100 399.600 ;
        RECT 606.100 398.400 606.700 399.600 ;
        RECT 606.000 397.600 606.800 398.400 ;
        RECT 607.700 372.400 608.300 403.600 ;
        RECT 612.500 396.400 613.100 427.600 ;
        RECT 612.400 395.600 613.200 396.400 ;
        RECT 607.600 371.600 608.400 372.400 ;
        RECT 604.400 351.600 605.200 352.400 ;
        RECT 598.000 349.600 599.000 350.400 ;
        RECT 604.400 349.600 605.200 350.400 ;
        RECT 594.800 337.600 595.600 338.400 ;
        RECT 585.200 333.600 586.000 334.400 ;
        RECT 590.000 333.600 590.800 334.400 ;
        RECT 593.200 333.600 594.000 334.400 ;
        RECT 585.300 332.400 585.900 333.600 ;
        RECT 585.200 331.600 586.000 332.400 ;
        RECT 593.200 331.600 594.000 332.400 ;
        RECT 593.300 330.400 593.900 331.600 ;
        RECT 594.900 330.400 595.500 337.600 ;
        RECT 598.100 336.400 598.700 349.600 ;
        RECT 599.600 347.600 600.400 348.400 ;
        RECT 601.200 347.600 602.000 348.400 ;
        RECT 606.000 347.600 606.800 348.400 ;
        RECT 598.000 335.600 598.800 336.400 ;
        RECT 599.700 334.400 600.300 347.600 ;
        RECT 599.600 333.600 600.400 334.400 ;
        RECT 599.700 332.400 600.300 333.600 ;
        RECT 599.600 331.600 600.400 332.400 ;
        RECT 580.500 329.700 582.700 330.300 ;
        RECT 546.900 318.400 547.500 323.600 ;
        RECT 546.800 317.600 547.600 318.400 ;
        RECT 542.000 305.600 542.800 306.400 ;
        RECT 534.000 303.600 534.800 304.400 ;
        RECT 537.200 303.600 538.000 304.400 ;
        RECT 542.000 303.600 542.800 304.400 ;
        RECT 546.800 303.600 547.600 304.400 ;
        RECT 554.800 303.600 555.600 304.400 ;
        RECT 558.000 304.200 558.800 317.800 ;
        RECT 559.600 304.200 560.400 317.800 ;
        RECT 561.200 304.200 562.000 315.800 ;
        RECT 562.800 307.600 563.600 308.400 ;
        RECT 564.400 304.200 565.200 315.800 ;
        RECT 566.000 305.600 566.800 306.400 ;
        RECT 566.100 304.400 566.700 305.600 ;
        RECT 566.000 303.600 566.800 304.400 ;
        RECT 567.600 304.200 568.400 315.800 ;
        RECT 569.200 304.200 570.000 317.800 ;
        RECT 570.800 304.200 571.600 317.800 ;
        RECT 572.400 304.200 573.200 317.800 ;
        RECT 575.600 311.600 576.400 312.400 ;
        RECT 574.000 309.600 574.800 310.400 ;
        RECT 574.100 306.400 574.700 309.600 ;
        RECT 574.000 305.600 574.800 306.400 ;
        RECT 532.400 293.600 533.200 294.400 ;
        RECT 534.100 292.400 534.700 303.600 ;
        RECT 537.300 296.400 537.900 303.600 ;
        RECT 537.200 295.600 538.000 296.400 ;
        RECT 542.100 294.400 542.700 303.600 ;
        RECT 535.600 293.600 536.400 294.400 ;
        RECT 542.000 293.600 542.800 294.400 ;
        RECT 534.000 291.600 534.800 292.400 ;
        RECT 530.800 289.600 531.600 290.400 ;
        RECT 529.200 283.600 530.000 284.400 ;
        RECT 529.300 280.400 529.900 283.600 ;
        RECT 530.800 281.600 531.600 282.400 ;
        RECT 529.200 279.600 530.000 280.400 ;
        RECT 530.900 278.400 531.500 281.600 ;
        RECT 530.800 277.600 531.600 278.400 ;
        RECT 532.400 277.600 533.200 278.400 ;
        RECT 527.600 275.600 528.400 276.400 ;
        RECT 527.600 272.300 528.400 272.400 ;
        RECT 526.100 271.700 528.400 272.300 ;
        RECT 527.600 271.600 528.400 271.700 ;
        RECT 527.600 269.600 528.400 270.400 ;
        RECT 530.800 269.600 531.600 270.400 ;
        RECT 522.800 267.600 523.600 268.400 ;
        RECT 513.200 265.600 514.000 266.400 ;
        RECT 514.800 265.600 515.600 266.400 ;
        RECT 516.400 265.600 517.200 266.400 ;
        RECT 521.200 265.600 522.000 266.400 ;
        RECT 524.400 265.600 525.200 266.400 ;
        RECT 521.300 264.400 521.900 265.600 ;
        RECT 521.200 263.600 522.000 264.400 ;
        RECT 519.600 261.600 520.400 262.400 ;
        RECT 514.800 259.600 515.600 260.400 ;
        RECT 514.900 258.400 515.500 259.600 ;
        RECT 519.700 258.400 520.300 261.600 ;
        RECT 522.800 259.600 523.600 260.400 ;
        RECT 511.600 257.600 512.400 258.400 ;
        RECT 514.800 257.600 515.600 258.400 ;
        RECT 518.000 257.600 518.800 258.400 ;
        RECT 519.600 257.600 520.400 258.400 ;
        RECT 510.000 255.600 510.800 256.400 ;
        RECT 516.400 255.600 517.200 256.400 ;
        RECT 510.100 252.400 510.700 255.600 ;
        RECT 508.400 251.600 509.200 252.400 ;
        RECT 510.000 251.600 510.800 252.400 ;
        RECT 511.600 251.600 512.400 252.400 ;
        RECT 513.200 251.600 514.000 252.400 ;
        RECT 502.000 249.600 502.800 250.400 ;
        RECT 500.400 245.600 501.200 246.400 ;
        RECT 500.400 241.600 501.200 242.400 ;
        RECT 500.500 230.400 501.100 241.600 ;
        RECT 502.100 230.400 502.700 249.600 ;
        RECT 508.500 248.400 509.100 251.600 ;
        RECT 511.700 250.400 512.300 251.600 ;
        RECT 511.600 249.600 512.400 250.400 ;
        RECT 508.400 247.600 509.200 248.400 ;
        RECT 505.200 245.600 506.000 246.400 ;
        RECT 503.600 243.600 504.400 244.400 ;
        RECT 503.700 242.400 504.300 243.600 ;
        RECT 503.600 241.600 504.400 242.400 ;
        RECT 505.300 236.400 505.900 245.600 ;
        RECT 506.800 243.600 507.600 244.400 ;
        RECT 506.900 238.400 507.500 243.600 ;
        RECT 506.800 237.600 507.600 238.400 ;
        RECT 505.200 235.600 506.000 236.400 ;
        RECT 506.800 235.600 507.600 236.400 ;
        RECT 500.400 229.600 501.200 230.400 ;
        RECT 502.000 229.600 502.800 230.400 ;
        RECT 500.400 227.600 501.200 228.400 ;
        RECT 500.500 222.400 501.100 227.600 ;
        RECT 500.400 221.600 501.200 222.400 ;
        RECT 505.300 220.400 505.900 235.600 ;
        RECT 508.500 234.400 509.100 247.600 ;
        RECT 510.000 245.600 510.800 246.400 ;
        RECT 508.400 233.600 509.200 234.400 ;
        RECT 508.400 231.600 509.200 232.400 ;
        RECT 506.800 229.600 507.600 230.400 ;
        RECT 508.500 228.400 509.100 231.600 ;
        RECT 508.400 228.300 509.200 228.400 ;
        RECT 510.100 228.300 510.700 245.600 ;
        RECT 513.300 238.400 513.900 251.600 ;
        RECT 516.500 250.400 517.100 255.600 ;
        RECT 518.100 254.400 518.700 257.600 ;
        RECT 518.000 253.600 518.800 254.400 ;
        RECT 522.900 252.400 523.500 259.600 ;
        RECT 518.000 251.600 518.800 252.400 ;
        RECT 519.600 251.600 520.400 252.400 ;
        RECT 522.800 251.600 523.600 252.400 ;
        RECT 516.400 249.600 517.200 250.400 ;
        RECT 514.800 239.600 515.600 240.400 ;
        RECT 513.200 237.600 514.000 238.400 ;
        RECT 511.600 235.600 512.400 236.400 ;
        RECT 511.700 234.400 512.300 235.600 ;
        RECT 511.600 233.600 512.400 234.400 ;
        RECT 514.900 232.400 515.500 239.600 ;
        RECT 518.100 232.400 518.700 251.600 ;
        RECT 522.800 239.600 523.600 240.400 ;
        RECT 519.600 233.600 520.400 234.400 ;
        RECT 522.900 232.400 523.500 239.600 ;
        RECT 524.500 238.400 525.100 265.600 ;
        RECT 527.700 258.400 528.300 269.600 ;
        RECT 529.200 267.600 530.000 268.400 ;
        RECT 529.300 258.400 529.900 267.600 ;
        RECT 530.900 260.400 531.500 269.600 ;
        RECT 530.800 259.600 531.600 260.400 ;
        RECT 527.600 257.600 528.400 258.400 ;
        RECT 529.200 257.600 530.000 258.400 ;
        RECT 526.000 253.600 526.800 254.400 ;
        RECT 526.100 250.300 526.700 253.600 ;
        RECT 530.900 252.400 531.500 259.600 ;
        RECT 527.600 251.600 528.400 252.400 ;
        RECT 530.800 251.600 531.600 252.400 ;
        RECT 526.100 249.700 528.300 250.300 ;
        RECT 524.400 237.600 525.200 238.400 ;
        RECT 526.000 235.600 526.800 236.400 ;
        RECT 526.100 234.400 526.700 235.600 ;
        RECT 526.000 233.600 526.800 234.400 ;
        RECT 514.800 231.600 515.600 232.400 ;
        RECT 518.000 231.600 518.800 232.400 ;
        RECT 522.800 231.600 523.600 232.400 ;
        RECT 524.400 231.600 525.200 232.400 ;
        RECT 524.500 230.400 525.100 231.600 ;
        RECT 513.200 229.600 514.000 230.400 ;
        RECT 516.400 229.600 517.200 230.400 ;
        RECT 518.000 229.600 518.800 230.400 ;
        RECT 524.400 229.600 525.200 230.400 ;
        RECT 513.300 228.400 513.900 229.600 ;
        RECT 508.400 227.700 510.700 228.300 ;
        RECT 508.400 227.600 509.200 227.700 ;
        RECT 513.200 227.600 514.000 228.400 ;
        RECT 498.900 219.700 501.100 220.300 ;
        RECT 486.000 213.600 486.800 214.400 ;
        RECT 484.400 211.600 485.200 212.400 ;
        RECT 489.200 209.600 490.000 210.400 ;
        RECT 466.800 203.600 467.600 204.400 ;
        RECT 470.000 203.600 470.800 204.400 ;
        RECT 473.200 203.600 474.000 204.400 ;
        RECT 476.400 203.600 477.200 204.400 ;
        RECT 479.600 203.600 480.400 204.400 ;
        RECT 442.800 199.600 443.600 200.400 ;
        RECT 450.800 199.600 451.600 200.400 ;
        RECT 438.000 189.600 438.800 190.400 ;
        RECT 438.100 188.400 438.700 189.600 ;
        RECT 434.800 187.600 435.600 188.400 ;
        RECT 438.000 187.600 438.800 188.400 ;
        RECT 438.000 185.600 438.800 186.400 ;
        RECT 433.200 173.600 434.000 174.400 ;
        RECT 431.600 171.600 432.400 172.400 ;
        RECT 433.200 171.600 434.000 172.400 ;
        RECT 426.900 157.700 429.100 158.300 ;
        RECT 426.900 134.400 427.500 157.700 ;
        RECT 428.400 155.600 429.200 156.400 ;
        RECT 428.500 152.400 429.100 155.600 ;
        RECT 428.400 151.600 429.200 152.400 ;
        RECT 431.600 151.600 432.400 152.400 ;
        RECT 428.500 150.400 429.100 151.600 ;
        RECT 428.400 149.600 429.200 150.400 ;
        RECT 430.000 149.600 430.800 150.400 ;
        RECT 434.800 149.600 435.600 150.400 ;
        RECT 431.600 143.600 432.400 144.400 ;
        RECT 431.600 137.600 432.400 138.400 ;
        RECT 426.800 133.600 427.600 134.400 ;
        RECT 431.700 132.400 432.300 137.600 ;
        RECT 433.200 133.600 434.000 134.400 ;
        RECT 431.600 131.600 432.400 132.400 ;
        RECT 433.200 131.600 434.000 132.400 ;
        RECT 433.300 130.400 433.900 131.600 ;
        RECT 428.400 129.600 429.200 130.400 ;
        RECT 433.200 129.600 434.000 130.400 ;
        RECT 426.800 125.600 427.600 126.400 ;
        RECT 425.200 119.600 426.000 120.400 ;
        RECT 426.900 118.400 427.500 125.600 ;
        RECT 428.500 122.400 429.100 129.600 ;
        RECT 433.200 127.600 434.000 128.400 ;
        RECT 431.600 123.600 432.400 124.400 ;
        RECT 428.400 121.600 429.200 122.400 ;
        RECT 422.000 117.600 422.800 118.400 ;
        RECT 426.800 117.600 427.600 118.400 ;
        RECT 431.700 116.400 432.300 123.600 ;
        RECT 415.600 109.600 416.400 110.400 ;
        RECT 415.700 108.400 416.300 109.600 ;
        RECT 418.800 109.400 419.600 110.400 ;
        RECT 415.600 107.600 416.400 108.400 ;
        RECT 420.400 104.200 421.200 115.800 ;
        RECT 428.400 115.600 429.200 116.400 ;
        RECT 431.600 115.600 432.400 116.400 ;
        RECT 428.500 112.400 429.100 115.600 ;
        RECT 422.000 111.600 422.800 112.400 ;
        RECT 418.800 99.600 419.600 100.400 ;
        RECT 414.000 93.600 414.800 94.400 ;
        RECT 418.900 92.400 419.500 99.600 ;
        RECT 422.100 98.400 422.700 111.600 ;
        RECT 423.600 106.200 424.400 111.800 ;
        RECT 428.400 111.600 429.200 112.400 ;
        RECT 428.400 109.600 429.200 110.400 ;
        RECT 428.500 108.400 429.100 109.600 ;
        RECT 433.300 108.400 433.900 127.600 ;
        RECT 428.400 107.600 429.200 108.400 ;
        RECT 433.200 107.600 434.000 108.400 ;
        RECT 425.200 105.600 426.000 106.400 ;
        RECT 422.000 97.600 422.800 98.400 ;
        RECT 420.400 95.600 421.200 96.400 ;
        RECT 412.400 91.600 413.200 92.400 ;
        RECT 418.800 91.600 419.600 92.400 ;
        RECT 406.000 83.600 406.800 84.400 ;
        RECT 375.600 69.600 376.400 70.400 ;
        RECT 378.800 69.600 379.600 70.400 ;
        RECT 390.000 69.600 390.800 70.400 ;
        RECT 367.600 67.600 368.400 68.400 ;
        RECT 377.200 67.600 378.000 68.400 ;
        RECT 367.700 66.400 368.300 67.600 ;
        RECT 362.800 65.600 363.600 66.400 ;
        RECT 366.000 65.600 366.800 66.400 ;
        RECT 367.600 65.600 368.400 66.400 ;
        RECT 372.400 65.600 373.200 66.400 ;
        RECT 346.800 63.600 347.600 64.400 ;
        RECT 370.800 63.600 371.600 64.400 ;
        RECT 346.900 54.400 347.500 63.600 ;
        RECT 377.300 62.400 377.900 67.600 ;
        RECT 370.800 61.600 371.600 62.400 ;
        RECT 377.200 61.600 378.000 62.400 ;
        RECT 353.200 59.600 354.000 60.400 ;
        RECT 353.300 58.400 353.900 59.600 ;
        RECT 370.900 58.400 371.500 61.600 ;
        RECT 353.200 57.600 354.000 58.400 ;
        RECT 354.800 57.600 355.600 58.400 ;
        RECT 362.800 57.600 363.600 58.400 ;
        RECT 367.600 57.600 368.400 58.400 ;
        RECT 370.800 57.600 371.600 58.400 ;
        RECT 354.900 56.400 355.500 57.600 ;
        RECT 354.800 55.600 355.600 56.400 ;
        RECT 361.200 55.600 362.000 56.400 ;
        RECT 362.900 54.400 363.500 57.600 ;
        RECT 369.200 55.600 370.000 56.400 ;
        RECT 378.900 54.400 379.500 69.600 ;
        RECT 388.400 67.600 389.200 68.400 ;
        RECT 385.200 63.600 386.000 64.400 ;
        RECT 346.800 53.600 347.600 54.400 ;
        RECT 348.400 53.600 349.200 54.400 ;
        RECT 351.600 53.600 352.400 54.400 ;
        RECT 354.800 53.600 355.600 54.400 ;
        RECT 356.400 53.600 357.200 54.400 ;
        RECT 362.800 53.600 363.600 54.400 ;
        RECT 378.800 53.600 379.600 54.400 ;
        RECT 348.500 52.400 349.100 53.600 ;
        RECT 348.400 51.600 349.200 52.400 ;
        RECT 343.600 50.300 344.400 50.400 ;
        RECT 345.200 50.300 346.000 50.400 ;
        RECT 343.600 49.700 346.000 50.300 ;
        RECT 343.600 49.600 344.400 49.700 ;
        RECT 345.200 49.600 346.000 49.700 ;
        RECT 340.400 45.600 341.200 46.400 ;
        RECT 338.800 37.600 339.600 38.400 ;
        RECT 337.400 31.800 338.200 32.600 ;
        RECT 338.900 32.400 339.500 37.600 ;
        RECT 335.600 27.600 336.400 28.400 ;
        RECT 335.700 26.400 336.300 27.600 ;
        RECT 337.400 27.000 338.000 31.800 ;
        RECT 338.800 31.600 339.600 32.400 ;
        RECT 343.600 31.800 344.400 32.600 ;
        RECT 338.600 29.800 339.400 30.600 ;
        RECT 338.800 28.400 339.400 29.800 ;
        RECT 343.800 28.400 344.400 31.800 ;
        RECT 345.300 28.400 345.900 49.600 ;
        RECT 346.800 45.600 347.600 46.400 ;
        RECT 346.900 32.400 347.500 45.600 ;
        RECT 351.700 38.400 352.300 53.600 ;
        RECT 354.900 46.400 355.500 53.600 ;
        RECT 354.800 45.600 355.600 46.400 ;
        RECT 356.500 38.400 357.100 53.600 ;
        RECT 358.000 51.600 358.800 52.400 ;
        RECT 361.200 51.600 362.000 52.400 ;
        RECT 358.100 50.400 358.700 51.600 ;
        RECT 361.300 50.400 361.900 51.600 ;
        RECT 362.900 50.400 363.500 53.600 ;
        RECT 364.400 51.600 365.200 52.400 ;
        RECT 375.600 51.600 376.400 52.400 ;
        RECT 358.000 49.600 358.800 50.400 ;
        RECT 361.200 49.600 362.000 50.400 ;
        RECT 362.800 49.600 363.600 50.400 ;
        RECT 351.600 37.600 352.400 38.400 ;
        RECT 356.400 37.600 357.200 38.400 ;
        RECT 350.000 33.600 350.800 34.400 ;
        RECT 346.800 31.600 347.600 32.400 ;
        RECT 338.800 27.800 344.400 28.400 ;
        RECT 338.800 27.000 339.600 27.200 ;
        RECT 342.200 27.000 343.000 27.200 ;
        RECT 343.800 27.000 344.400 27.800 ;
        RECT 345.200 27.600 346.000 28.400 ;
        RECT 337.400 26.400 343.000 27.000 ;
        RECT 335.600 25.600 336.400 26.400 ;
        RECT 337.400 26.200 338.200 26.400 ;
        RECT 343.600 26.200 344.400 27.000 ;
        RECT 346.900 26.400 347.500 31.600 ;
        RECT 348.400 29.600 349.200 30.400 ;
        RECT 348.500 28.400 349.100 29.600 ;
        RECT 348.400 27.600 349.200 28.400 ;
        RECT 346.800 25.600 347.600 26.400 ;
        RECT 327.600 19.600 328.400 20.400 ;
        RECT 334.000 19.600 334.800 20.400 ;
        RECT 311.600 17.600 312.400 18.400 ;
        RECT 297.200 11.600 298.000 12.400 ;
        RECT 310.000 11.600 310.800 12.400 ;
        RECT 318.000 11.600 318.800 12.400 ;
        RECT 322.800 4.200 323.600 17.800 ;
        RECT 324.400 4.200 325.200 17.800 ;
        RECT 326.000 6.200 326.800 17.800 ;
        RECT 327.700 14.400 328.300 19.600 ;
        RECT 346.900 18.400 347.500 25.600 ;
        RECT 327.600 13.600 328.400 14.400 ;
        RECT 329.200 6.200 330.000 17.800 ;
        RECT 330.800 17.600 331.600 18.400 ;
        RECT 330.900 16.400 331.500 17.600 ;
        RECT 330.800 15.600 331.600 16.400 ;
        RECT 332.400 6.200 333.200 17.800 ;
        RECT 334.000 4.200 334.800 17.800 ;
        RECT 335.600 4.200 336.400 17.800 ;
        RECT 337.200 4.200 338.000 17.800 ;
        RECT 346.800 17.600 347.600 18.400 ;
        RECT 348.500 14.400 349.100 27.600 ;
        RECT 350.100 16.400 350.700 33.600 ;
        RECT 356.400 29.600 357.200 30.400 ;
        RECT 353.200 25.600 354.000 26.400 ;
        RECT 356.500 16.400 357.100 29.600 ;
        RECT 361.300 26.400 361.900 49.600 ;
        RECT 380.400 44.200 381.200 57.800 ;
        RECT 382.000 44.200 382.800 57.800 ;
        RECT 383.600 46.200 384.400 57.800 ;
        RECT 385.300 56.400 385.900 63.600 ;
        RECT 388.500 58.400 389.100 67.600 ;
        RECT 390.100 60.400 390.700 69.600 ;
        RECT 393.300 64.400 393.900 71.600 ;
        RECT 394.900 68.400 395.500 71.600 ;
        RECT 394.800 67.600 395.600 68.400 ;
        RECT 396.200 67.000 396.800 71.800 ;
        RECT 401.200 71.600 402.000 72.400 ;
        RECT 402.800 71.800 403.600 72.600 ;
        RECT 398.800 68.400 399.600 68.600 ;
        RECT 403.000 68.400 403.600 71.800 ;
        RECT 406.100 68.400 406.700 83.600 ;
        RECT 410.800 73.600 411.600 74.400 ;
        RECT 410.800 69.600 411.600 70.400 ;
        RECT 398.800 67.800 403.600 68.400 ;
        RECT 398.000 67.000 398.800 67.200 ;
        RECT 401.400 67.000 402.200 67.200 ;
        RECT 403.000 67.000 403.600 67.800 ;
        RECT 406.000 67.600 406.800 68.400 ;
        RECT 407.600 67.600 408.400 68.400 ;
        RECT 409.200 67.600 410.000 68.400 ;
        RECT 396.200 66.200 397.000 67.000 ;
        RECT 398.000 66.400 402.200 67.000 ;
        RECT 402.800 66.200 403.600 67.000 ;
        RECT 409.300 64.400 409.900 67.600 ;
        RECT 412.500 66.400 413.100 91.600 ;
        RECT 415.600 89.600 416.400 90.400 ;
        RECT 415.700 88.400 416.300 89.600 ;
        RECT 415.600 87.600 416.400 88.400 ;
        RECT 420.500 72.400 421.100 95.600 ;
        RECT 425.300 94.300 425.900 105.600 ;
        RECT 433.300 98.400 433.900 107.600 ;
        RECT 434.900 102.400 435.500 149.600 ;
        RECT 438.100 146.400 438.700 185.600 ;
        RECT 442.800 184.200 443.600 197.800 ;
        RECT 444.400 184.200 445.200 197.800 ;
        RECT 446.000 184.200 446.800 195.800 ;
        RECT 447.600 187.600 448.400 188.400 ;
        RECT 447.700 182.400 448.300 187.600 ;
        RECT 449.200 184.200 450.000 195.800 ;
        RECT 450.900 188.400 451.500 199.600 ;
        RECT 450.800 187.600 451.600 188.400 ;
        RECT 450.900 186.400 451.500 187.600 ;
        RECT 450.800 185.600 451.600 186.400 ;
        RECT 452.400 184.200 453.200 195.800 ;
        RECT 454.000 184.200 454.800 197.800 ;
        RECT 455.600 184.200 456.400 197.800 ;
        RECT 457.200 184.200 458.000 197.800 ;
        RECT 466.900 190.400 467.500 203.600 ;
        RECT 466.800 189.600 467.600 190.400 ;
        RECT 466.800 183.600 467.600 184.400 ;
        RECT 447.600 181.600 448.400 182.400 ;
        RECT 450.800 181.600 451.600 182.400 ;
        RECT 439.600 166.200 440.400 177.800 ;
        RECT 446.000 173.600 446.800 174.400 ;
        RECT 444.400 169.600 445.200 170.400 ;
        RECT 444.500 164.400 445.100 169.600 ;
        RECT 446.100 168.400 446.700 173.600 ;
        RECT 447.600 171.600 448.400 172.400 ;
        RECT 449.200 171.600 450.000 172.400 ;
        RECT 446.000 167.600 446.800 168.400 ;
        RECT 447.700 166.300 448.300 171.600 ;
        RECT 446.100 165.700 448.300 166.300 ;
        RECT 444.400 164.300 445.200 164.400 ;
        RECT 442.900 163.700 445.200 164.300 ;
        RECT 442.900 150.400 443.500 163.700 ;
        RECT 444.400 163.600 445.200 163.700 ;
        RECT 446.100 158.400 446.700 165.700 ;
        RECT 446.000 157.600 446.800 158.400 ;
        RECT 450.900 154.400 451.500 181.600 ;
        RECT 457.200 173.600 458.000 174.400 ;
        RECT 452.400 169.600 453.200 170.400 ;
        RECT 457.300 168.400 457.900 173.600 ;
        RECT 463.600 171.600 464.400 172.400 ;
        RECT 452.400 167.600 453.200 168.400 ;
        RECT 457.200 167.600 458.000 168.400 ;
        RECT 450.800 153.600 451.600 154.400 ;
        RECT 447.600 152.300 448.400 152.400 ;
        RECT 447.600 151.700 449.900 152.300 ;
        RECT 447.600 151.600 448.400 151.700 ;
        RECT 449.300 150.400 449.900 151.700 ;
        RECT 450.800 151.600 451.600 152.400 ;
        RECT 441.200 149.600 442.000 150.400 ;
        RECT 442.800 149.600 443.600 150.400 ;
        RECT 447.600 149.600 448.400 150.400 ;
        RECT 449.200 149.600 450.000 150.400 ;
        RECT 438.000 145.600 438.800 146.400 ;
        RECT 439.600 145.600 440.400 146.400 ;
        RECT 439.700 140.400 440.300 145.600 ;
        RECT 439.600 139.600 440.400 140.400 ;
        RECT 441.300 136.400 441.900 149.600 ;
        RECT 441.200 135.600 442.000 136.400 ;
        RECT 438.000 133.600 438.800 134.400 ;
        RECT 436.400 121.600 437.200 122.400 ;
        RECT 436.500 110.400 437.100 121.600 ;
        RECT 441.300 114.400 441.900 135.600 ;
        RECT 442.900 130.300 443.500 149.600 ;
        RECT 447.600 135.600 448.400 136.400 ;
        RECT 444.400 131.600 445.200 132.400 ;
        RECT 444.400 130.300 445.200 130.400 ;
        RECT 442.900 129.700 445.200 130.300 ;
        RECT 444.400 129.600 445.200 129.700 ;
        RECT 442.800 127.600 443.600 128.400 ;
        RECT 441.200 113.600 442.000 114.400 ;
        RECT 439.600 111.600 440.400 112.400 ;
        RECT 436.400 109.600 437.200 110.400 ;
        RECT 434.800 101.600 435.600 102.400 ;
        RECT 428.400 97.600 429.200 98.400 ;
        RECT 433.200 97.600 434.000 98.400 ;
        RECT 430.000 95.600 430.800 96.400 ;
        RECT 425.300 93.700 427.500 94.300 ;
        RECT 426.900 92.400 427.500 93.700 ;
        RECT 423.600 91.600 424.400 92.400 ;
        RECT 425.200 91.600 426.000 92.400 ;
        RECT 426.800 91.600 427.600 92.400 ;
        RECT 423.700 80.400 424.300 91.600 ;
        RECT 425.200 89.600 426.000 90.400 ;
        RECT 425.300 84.400 425.900 89.600 ;
        RECT 425.200 83.600 426.000 84.400 ;
        RECT 423.600 79.600 424.400 80.400 ;
        RECT 414.000 71.600 414.800 72.400 ;
        RECT 417.200 71.600 418.000 72.400 ;
        RECT 420.400 71.600 421.200 72.400 ;
        RECT 422.000 71.600 422.800 72.400 ;
        RECT 417.200 69.600 418.000 70.400 ;
        RECT 415.600 67.600 416.400 68.400 ;
        RECT 412.400 65.600 413.200 66.400 ;
        RECT 417.300 64.400 417.900 69.600 ;
        RECT 393.200 63.600 394.000 64.400 ;
        RECT 409.200 63.600 410.000 64.400 ;
        RECT 417.200 63.600 418.000 64.400 ;
        RECT 399.600 61.600 400.400 62.400 ;
        RECT 418.800 61.600 419.600 62.400 ;
        RECT 390.000 59.600 390.800 60.400 ;
        RECT 385.200 55.600 386.000 56.400 ;
        RECT 385.200 53.600 386.000 54.400 ;
        RECT 385.200 51.600 386.000 52.400 ;
        RECT 367.600 29.600 368.400 30.400 ;
        RECT 359.600 25.600 360.400 26.400 ;
        RECT 361.200 25.600 362.000 26.400 ;
        RECT 362.800 25.600 363.600 26.400 ;
        RECT 362.900 16.400 363.500 25.600 ;
        RECT 350.000 15.600 350.800 16.400 ;
        RECT 356.400 15.600 357.200 16.400 ;
        RECT 359.600 15.600 360.400 16.400 ;
        RECT 362.800 15.600 363.600 16.400 ;
        RECT 348.400 13.600 349.200 14.400 ;
        RECT 359.600 13.600 360.400 14.400 ;
        RECT 367.700 12.400 368.300 29.600 ;
        RECT 369.200 24.200 370.000 37.800 ;
        RECT 370.800 24.200 371.600 37.800 ;
        RECT 372.400 24.200 373.200 37.800 ;
        RECT 374.000 24.200 374.800 35.800 ;
        RECT 375.600 25.600 376.400 26.400 ;
        RECT 375.700 22.400 376.300 25.600 ;
        RECT 377.200 24.200 378.000 35.800 ;
        RECT 378.800 27.600 379.600 28.400 ;
        RECT 380.400 24.200 381.200 35.800 ;
        RECT 382.000 24.200 382.800 37.800 ;
        RECT 383.600 24.200 384.400 37.800 ;
        RECT 385.300 30.400 385.900 51.600 ;
        RECT 386.800 46.200 387.600 57.800 ;
        RECT 388.400 57.600 389.200 58.400 ;
        RECT 388.400 55.600 389.200 56.400 ;
        RECT 390.000 46.200 390.800 57.800 ;
        RECT 391.600 44.200 392.400 57.800 ;
        RECT 393.200 44.200 394.000 57.800 ;
        RECT 394.800 44.200 395.600 57.800 ;
        RECT 385.200 29.600 386.000 30.400 ;
        RECT 394.800 23.600 395.600 24.400 ;
        RECT 375.600 21.600 376.400 22.400 ;
        RECT 380.400 21.600 381.200 22.400 ;
        RECT 367.600 11.600 368.400 12.400 ;
        RECT 372.400 4.200 373.200 17.800 ;
        RECT 374.000 4.200 374.800 17.800 ;
        RECT 375.600 6.200 376.400 17.800 ;
        RECT 377.200 13.600 378.000 14.400 ;
        RECT 378.800 6.200 379.600 17.800 ;
        RECT 380.500 16.400 381.100 21.600 ;
        RECT 394.900 18.400 395.500 23.600 ;
        RECT 380.400 15.600 381.200 16.400 ;
        RECT 382.000 6.200 382.800 17.800 ;
        RECT 383.600 4.200 384.400 17.800 ;
        RECT 385.200 4.200 386.000 17.800 ;
        RECT 386.800 4.200 387.600 17.800 ;
        RECT 394.800 17.600 395.600 18.400 ;
        RECT 396.400 17.600 397.200 18.400 ;
        RECT 399.700 12.400 400.300 61.600 ;
        RECT 404.400 59.600 405.200 60.400 ;
        RECT 404.500 58.400 405.100 59.600 ;
        RECT 404.400 57.600 405.200 58.400 ;
        RECT 407.600 50.200 408.400 55.800 ;
        RECT 409.200 55.600 410.000 56.400 ;
        RECT 409.300 54.400 409.900 55.600 ;
        RECT 409.200 53.600 410.000 54.400 ;
        RECT 407.600 27.600 408.400 28.400 ;
        RECT 399.600 11.600 400.400 12.400 ;
        RECT 404.400 10.200 405.200 15.800 ;
        RECT 407.600 6.200 408.400 17.800 ;
        RECT 409.300 16.400 409.900 53.600 ;
        RECT 410.800 46.200 411.600 57.800 ;
        RECT 414.000 53.600 414.800 54.400 ;
        RECT 414.100 52.400 414.700 53.600 ;
        RECT 418.900 52.400 419.500 61.600 ;
        RECT 420.500 60.400 421.100 71.600 ;
        RECT 422.100 68.400 422.700 71.600 ;
        RECT 423.700 70.400 424.300 79.600 ;
        RECT 425.300 74.400 425.900 83.600 ;
        RECT 426.900 76.400 427.500 91.600 ;
        RECT 428.400 87.600 429.200 88.400 ;
        RECT 428.500 78.400 429.100 87.600 ;
        RECT 430.100 84.400 430.700 95.600 ;
        RECT 433.300 94.400 433.900 97.600 ;
        RECT 433.200 93.600 434.000 94.400 ;
        RECT 438.000 93.600 438.800 94.400 ;
        RECT 439.700 92.400 440.300 111.600 ;
        RECT 441.200 109.600 442.000 110.400 ;
        RECT 441.300 100.400 441.900 109.600 ;
        RECT 442.900 108.400 443.500 127.600 ;
        RECT 447.700 126.400 448.300 135.600 ;
        RECT 452.500 134.400 453.100 167.600 ;
        RECT 454.000 165.600 454.800 166.400 ;
        RECT 454.100 148.400 454.700 165.600 ;
        RECT 460.400 155.600 461.200 156.400 ;
        RECT 455.600 153.600 456.400 154.400 ;
        RECT 454.000 147.600 454.800 148.400 ;
        RECT 455.700 138.400 456.300 153.600 ;
        RECT 463.700 144.400 464.300 171.600 ;
        RECT 465.200 169.600 466.000 170.400 ;
        RECT 466.900 156.400 467.500 183.600 ;
        RECT 470.100 176.400 470.700 203.600 ;
        RECT 470.000 175.600 470.800 176.400 ;
        RECT 470.000 173.600 470.800 174.400 ;
        RECT 468.400 169.600 469.200 170.400 ;
        RECT 468.500 166.400 469.100 169.600 ;
        RECT 468.400 165.600 469.200 166.400 ;
        RECT 470.100 160.400 470.700 173.600 ;
        RECT 471.600 171.600 472.400 172.400 ;
        RECT 470.000 159.600 470.800 160.400 ;
        RECT 463.600 143.600 464.400 144.400 ;
        RECT 465.200 144.200 466.000 155.800 ;
        RECT 466.800 155.600 467.600 156.400 ;
        RECT 470.000 155.600 470.800 156.400 ;
        RECT 466.800 149.600 467.600 150.400 ;
        RECT 463.700 138.400 464.300 143.600 ;
        RECT 455.600 137.600 456.400 138.400 ;
        RECT 463.600 137.600 464.400 138.400 ;
        RECT 453.800 135.000 454.600 135.800 ;
        RECT 455.600 135.000 459.800 135.600 ;
        RECT 460.400 135.000 461.200 135.800 ;
        RECT 452.400 133.600 453.200 134.400 ;
        RECT 449.200 131.600 450.000 132.400 ;
        RECT 450.800 131.600 451.600 132.400 ;
        RECT 447.600 125.600 448.400 126.400 ;
        RECT 444.400 123.600 445.200 124.400 ;
        RECT 444.500 116.400 445.100 123.600 ;
        RECT 446.000 119.600 446.800 120.400 ;
        RECT 444.400 115.600 445.200 116.400 ;
        RECT 446.100 114.400 446.700 119.600 ;
        RECT 446.000 113.600 446.800 114.400 ;
        RECT 444.400 111.600 445.200 112.400 ;
        RECT 444.400 110.300 445.200 110.400 ;
        RECT 446.100 110.300 446.700 113.600 ;
        RECT 444.400 109.700 446.700 110.300 ;
        RECT 444.400 109.600 445.200 109.700 ;
        RECT 442.800 107.600 443.600 108.400 ;
        RECT 441.200 99.600 442.000 100.400 ;
        RECT 433.200 91.600 434.000 92.400 ;
        RECT 436.400 91.600 437.200 92.400 ;
        RECT 439.600 91.600 440.400 92.400 ;
        RECT 441.200 91.600 442.000 92.400 ;
        RECT 442.900 92.300 443.500 107.600 ;
        RECT 449.300 106.400 449.900 131.600 ;
        RECT 450.900 128.400 451.500 131.600 ;
        RECT 452.400 129.600 453.200 130.400 ;
        RECT 453.800 130.200 454.400 135.000 ;
        RECT 455.600 134.800 456.400 135.000 ;
        RECT 459.000 134.800 459.800 135.000 ;
        RECT 460.600 134.200 461.200 135.000 ;
        RECT 456.400 133.600 461.200 134.200 ;
        RECT 456.400 133.400 457.200 133.600 ;
        RECT 460.600 130.200 461.200 133.600 ;
        RECT 450.800 127.600 451.600 128.400 ;
        RECT 450.800 115.600 451.600 116.400 ;
        RECT 450.900 112.400 451.500 115.600 ;
        RECT 450.800 111.600 451.600 112.400 ;
        RECT 450.800 109.600 451.600 110.400 ;
        RECT 444.400 105.600 445.200 106.400 ;
        RECT 447.600 105.600 448.400 106.400 ;
        RECT 449.200 105.600 450.000 106.400 ;
        RECT 447.700 96.400 448.300 105.600 ;
        RECT 449.200 103.600 450.000 104.400 ;
        RECT 449.300 98.400 449.900 103.600 ;
        RECT 450.900 100.400 451.500 109.600 ;
        RECT 452.500 104.400 453.100 129.600 ;
        RECT 453.800 129.400 454.600 130.200 ;
        RECT 460.400 129.400 461.200 130.200 ;
        RECT 454.000 109.600 454.800 110.400 ;
        RECT 455.600 109.600 456.400 110.400 ;
        RECT 452.400 103.600 453.200 104.400 ;
        RECT 450.800 99.600 451.600 100.400 ;
        RECT 449.200 97.600 450.000 98.400 ;
        RECT 447.600 95.600 448.400 96.400 ;
        RECT 452.400 95.600 453.200 96.400 ;
        RECT 447.600 93.600 448.400 94.400 ;
        RECT 444.400 92.300 445.200 92.400 ;
        RECT 442.900 91.700 445.200 92.300 ;
        RECT 444.400 91.600 445.200 91.700 ;
        RECT 430.000 83.600 430.800 84.400 ;
        RECT 428.400 77.600 429.200 78.400 ;
        RECT 426.800 75.600 427.600 76.400 ;
        RECT 425.200 73.600 426.000 74.400 ;
        RECT 425.200 71.600 426.000 72.400 ;
        RECT 426.800 71.600 427.600 72.400 ;
        RECT 430.000 71.600 430.800 72.400 ;
        RECT 423.600 69.600 424.400 70.400 ;
        RECT 425.300 68.400 425.900 71.600 ;
        RECT 426.900 70.400 427.500 71.600 ;
        RECT 426.800 69.600 427.600 70.400 ;
        RECT 428.400 69.600 429.200 70.400 ;
        RECT 428.500 68.400 429.100 69.600 ;
        RECT 422.000 67.600 422.800 68.400 ;
        RECT 425.200 67.600 426.000 68.400 ;
        RECT 428.400 67.600 429.200 68.400 ;
        RECT 423.600 65.600 424.400 66.400 ;
        RECT 423.700 64.400 424.300 65.600 ;
        RECT 423.600 63.600 424.400 64.400 ;
        RECT 420.400 59.600 421.200 60.400 ;
        RECT 422.000 59.600 422.800 60.400 ;
        RECT 414.000 51.600 414.800 52.400 ;
        RECT 418.800 51.600 419.600 52.400 ;
        RECT 418.900 38.400 419.500 51.600 ;
        RECT 420.400 46.200 421.200 57.800 ;
        RECT 422.100 50.400 422.700 59.600 ;
        RECT 423.700 52.400 424.300 63.600 ;
        RECT 425.200 57.600 426.000 58.400 ;
        RECT 425.300 56.300 425.900 57.600 ;
        RECT 426.800 56.300 427.600 56.400 ;
        RECT 425.300 55.700 427.600 56.300 ;
        RECT 426.800 55.600 427.600 55.700 ;
        RECT 423.600 51.600 424.400 52.400 ;
        RECT 422.000 49.600 422.800 50.400 ;
        RECT 418.800 37.600 419.600 38.400 ;
        RECT 422.100 28.400 422.700 49.600 ;
        RECT 426.800 31.600 427.600 32.400 ;
        RECT 428.500 30.400 429.100 67.600 ;
        RECT 430.100 34.400 430.700 71.600 ;
        RECT 431.600 51.600 432.400 52.400 ;
        RECT 431.600 49.600 432.400 50.400 ;
        RECT 431.700 38.400 432.300 49.600 ;
        RECT 431.600 37.600 432.400 38.400 ;
        RECT 430.000 33.600 430.800 34.400 ;
        RECT 423.600 29.600 424.400 30.400 ;
        RECT 426.800 29.600 427.600 30.400 ;
        RECT 428.400 29.600 429.200 30.400 ;
        RECT 431.600 29.600 432.400 30.400 ;
        RECT 422.000 27.600 422.800 28.400 ;
        RECT 425.200 27.600 426.000 28.400 ;
        RECT 423.600 21.600 424.400 22.400 ;
        RECT 409.200 15.600 410.000 16.400 ;
        RECT 410.800 13.600 411.600 14.400 ;
        RECT 410.900 12.400 411.500 13.600 ;
        RECT 410.800 11.600 411.600 12.400 ;
        RECT 417.200 6.200 418.000 17.800 ;
        RECT 423.700 12.400 424.300 21.600 ;
        RECT 425.300 14.400 425.900 27.600 ;
        RECT 426.900 18.400 427.500 29.600 ;
        RECT 433.300 22.400 433.900 91.600 ;
        RECT 439.600 83.600 440.400 84.400 ;
        RECT 438.000 77.600 438.800 78.400 ;
        RECT 438.100 70.400 438.700 77.600 ;
        RECT 439.700 70.400 440.300 83.600 ;
        RECT 441.300 78.400 441.900 91.600 ;
        RECT 444.500 90.400 445.100 91.600 ;
        RECT 442.800 89.600 443.600 90.400 ;
        RECT 444.400 89.600 445.200 90.400 ;
        RECT 441.200 77.600 442.000 78.400 ;
        RECT 438.000 69.600 438.800 70.400 ;
        RECT 439.600 69.600 440.400 70.400 ;
        RECT 441.200 69.600 442.000 70.400 ;
        RECT 442.900 70.300 443.500 89.600 ;
        RECT 446.000 79.600 446.800 80.400 ;
        RECT 446.100 74.400 446.700 79.600 ;
        RECT 444.400 73.600 445.200 74.400 ;
        RECT 446.000 73.600 446.800 74.400 ;
        RECT 444.500 72.400 445.100 73.600 ;
        RECT 446.100 72.400 446.700 73.600 ;
        RECT 444.400 71.600 445.200 72.400 ;
        RECT 446.000 71.600 446.800 72.400 ;
        RECT 444.400 70.300 445.200 70.400 ;
        RECT 442.900 69.700 445.200 70.300 ;
        RECT 444.400 69.600 445.200 69.700 ;
        RECT 439.600 67.600 440.400 68.400 ;
        RECT 434.800 63.600 435.600 64.400 ;
        RECT 434.900 60.400 435.500 63.600 ;
        RECT 434.800 59.600 435.600 60.400 ;
        RECT 439.700 58.400 440.300 67.600 ;
        RECT 441.300 64.400 441.900 69.600 ;
        RECT 447.700 68.400 448.300 93.600 ;
        RECT 452.500 92.400 453.100 95.600 ;
        RECT 449.200 91.600 450.000 92.400 ;
        RECT 452.400 91.600 453.200 92.400 ;
        RECT 449.200 89.600 450.000 90.400 ;
        RECT 452.400 71.600 453.200 72.400 ;
        RECT 449.200 69.600 450.000 70.400 ;
        RECT 447.600 67.600 448.400 68.400 ;
        RECT 441.200 63.600 442.000 64.400 ;
        RECT 434.800 57.600 435.600 58.400 ;
        RECT 439.600 57.600 440.400 58.400 ;
        RECT 436.400 55.600 437.200 56.400 ;
        RECT 442.800 56.300 443.600 56.400 ;
        RECT 439.700 55.700 443.600 56.300 ;
        RECT 436.500 50.400 437.100 55.600 ;
        RECT 439.700 54.400 440.300 55.700 ;
        RECT 442.800 55.600 443.600 55.700 ;
        RECT 444.400 55.600 445.200 56.400 ;
        RECT 446.000 55.600 446.800 56.400 ;
        RECT 439.600 53.600 440.400 54.400 ;
        RECT 441.200 53.600 442.000 54.400 ;
        RECT 439.600 52.300 440.400 52.400 ;
        RECT 438.100 51.700 440.400 52.300 ;
        RECT 434.800 49.600 435.600 50.400 ;
        RECT 436.400 49.600 437.200 50.400 ;
        RECT 434.800 31.600 435.600 32.400 ;
        RECT 436.400 31.600 437.200 32.400 ;
        RECT 433.200 21.600 434.000 22.400 ;
        RECT 433.200 19.600 434.000 20.400 ;
        RECT 433.300 18.400 433.900 19.600 ;
        RECT 426.800 17.600 427.600 18.400 ;
        RECT 433.200 17.600 434.000 18.400 ;
        RECT 425.200 13.600 426.000 14.400 ;
        RECT 423.600 11.600 424.400 12.400 ;
        RECT 425.200 11.600 426.000 12.400 ;
        RECT 430.000 11.600 430.800 12.400 ;
        RECT 425.300 8.400 425.900 11.600 ;
        RECT 434.900 8.400 435.500 31.600 ;
        RECT 436.500 30.400 437.100 31.600 ;
        RECT 438.100 30.400 438.700 51.700 ;
        RECT 439.600 51.600 440.400 51.700 ;
        RECT 439.600 49.600 440.400 50.400 ;
        RECT 436.400 29.600 437.200 30.400 ;
        RECT 438.000 29.600 438.800 30.400 ;
        RECT 439.600 28.300 440.400 28.400 ;
        RECT 441.300 28.300 441.900 53.600 ;
        RECT 444.500 50.400 445.100 55.600 ;
        RECT 446.100 52.400 446.700 55.600 ;
        RECT 447.700 54.400 448.300 67.600 ;
        RECT 449.300 60.400 449.900 69.600 ;
        RECT 450.800 67.600 451.600 68.400 ;
        RECT 449.200 59.600 450.000 60.400 ;
        RECT 447.600 53.600 448.400 54.400 ;
        RECT 449.300 52.400 449.900 59.600 ;
        RECT 450.900 54.400 451.500 67.600 ;
        RECT 454.100 66.400 454.700 109.600 ;
        RECT 455.700 108.400 456.300 109.600 ;
        RECT 455.600 107.600 456.400 108.400 ;
        RECT 462.000 107.600 462.800 108.400 ;
        RECT 463.600 103.600 464.400 104.400 ;
        RECT 463.700 102.400 464.300 103.600 ;
        RECT 463.600 101.600 464.400 102.400 ;
        RECT 463.700 96.400 464.300 101.600 ;
        RECT 466.900 96.400 467.500 149.600 ;
        RECT 470.100 136.400 470.700 155.600 ;
        RECT 471.600 149.600 472.400 150.400 ;
        RECT 471.700 148.400 472.300 149.600 ;
        RECT 471.600 147.600 472.400 148.400 ;
        RECT 471.600 145.600 472.400 146.400 ;
        RECT 470.000 135.600 470.800 136.400 ;
        RECT 468.400 109.600 469.200 110.400 ;
        RECT 470.100 108.300 470.700 135.600 ;
        RECT 471.700 114.400 472.300 145.600 ;
        RECT 473.300 138.400 473.900 203.600 ;
        RECT 476.500 192.400 477.100 203.600 ;
        RECT 479.700 196.400 480.300 203.600 ;
        RECT 474.800 186.200 475.600 191.800 ;
        RECT 476.400 191.600 477.200 192.400 ;
        RECT 476.400 189.600 477.200 190.400 ;
        RECT 474.800 177.600 475.600 178.400 ;
        RECT 474.900 172.400 475.500 177.600 ;
        RECT 476.500 174.400 477.100 189.600 ;
        RECT 478.000 184.200 478.800 195.800 ;
        RECT 479.600 195.600 480.400 196.400 ;
        RECT 479.600 189.400 480.400 190.400 ;
        RECT 481.200 187.600 482.000 188.400 ;
        RECT 487.600 184.200 488.400 195.800 ;
        RECT 489.300 194.400 489.900 209.600 ;
        RECT 495.600 204.200 496.400 217.800 ;
        RECT 497.200 204.200 498.000 217.800 ;
        RECT 498.800 206.200 499.600 217.800 ;
        RECT 500.500 214.400 501.100 219.700 ;
        RECT 505.200 219.600 506.000 220.400 ;
        RECT 500.400 213.600 501.200 214.400 ;
        RECT 502.000 206.200 502.800 217.800 ;
        RECT 503.600 215.600 504.400 216.400 ;
        RECT 503.700 210.400 504.300 215.600 ;
        RECT 503.600 209.600 504.400 210.400 ;
        RECT 505.200 206.200 506.000 217.800 ;
        RECT 506.800 204.200 507.600 217.800 ;
        RECT 508.400 204.200 509.200 217.800 ;
        RECT 510.000 204.200 510.800 217.800 ;
        RECT 511.600 215.600 512.400 216.400 ;
        RECT 511.700 212.400 512.300 215.600 ;
        RECT 516.500 214.400 517.100 229.600 ;
        RECT 518.100 222.400 518.700 229.600 ;
        RECT 519.600 227.600 520.400 228.400 ;
        RECT 519.600 225.600 520.400 226.400 ;
        RECT 526.000 225.600 526.800 226.400 ;
        RECT 518.000 221.600 518.800 222.400 ;
        RECT 519.700 218.400 520.300 225.600 ;
        RECT 522.800 221.600 523.600 222.400 ;
        RECT 519.600 217.600 520.400 218.400 ;
        RECT 516.400 213.600 517.200 214.400 ;
        RECT 519.700 212.400 520.300 217.600 ;
        RECT 522.900 216.400 523.500 221.600 ;
        RECT 522.800 215.600 523.600 216.400 ;
        RECT 526.100 214.400 526.700 225.600 ;
        RECT 526.000 213.600 526.800 214.400 ;
        RECT 527.700 212.400 528.300 249.700 ;
        RECT 530.800 235.600 531.600 236.400 ;
        RECT 530.800 233.600 531.600 234.400 ;
        RECT 529.200 231.600 530.000 232.400 ;
        RECT 530.800 231.600 531.600 232.400 ;
        RECT 529.300 222.400 529.900 231.600 ;
        RECT 530.900 230.400 531.500 231.600 ;
        RECT 530.800 229.600 531.600 230.400 ;
        RECT 530.800 223.600 531.600 224.400 ;
        RECT 529.200 221.600 530.000 222.400 ;
        RECT 511.600 211.600 512.400 212.400 ;
        RECT 519.600 211.600 520.400 212.400 ;
        RECT 527.600 211.600 528.400 212.400 ;
        RECT 530.900 210.400 531.500 223.600 ;
        RECT 532.500 218.400 533.100 277.600 ;
        RECT 534.100 276.400 534.700 291.600 ;
        RECT 538.800 289.600 539.600 290.400 ;
        RECT 537.200 279.600 538.000 280.400 ;
        RECT 534.000 275.600 534.800 276.400 ;
        RECT 534.000 273.600 534.800 274.400 ;
        RECT 534.100 270.400 534.700 273.600 ;
        RECT 537.300 272.400 537.900 279.600 ;
        RECT 537.200 271.600 538.000 272.400 ;
        RECT 540.400 271.600 541.200 272.400 ;
        RECT 545.200 271.600 546.000 272.400 ;
        RECT 534.000 269.600 534.800 270.400 ;
        RECT 535.600 267.600 536.400 268.400 ;
        RECT 535.700 262.400 536.300 267.600 ;
        RECT 535.600 261.600 536.400 262.400 ;
        RECT 534.000 255.600 534.800 256.400 ;
        RECT 535.600 255.600 536.400 256.400 ;
        RECT 534.000 252.300 534.800 252.400 ;
        RECT 535.700 252.300 536.300 255.600 ;
        RECT 537.300 254.400 537.900 271.600 ;
        RECT 538.800 269.600 539.600 270.400 ;
        RECT 538.900 264.400 539.500 269.600 ;
        RECT 540.500 268.400 541.100 271.600 ;
        RECT 540.400 267.600 541.200 268.400 ;
        RECT 543.600 265.600 544.400 266.400 ;
        RECT 538.800 263.600 539.600 264.400 ;
        RECT 542.000 263.600 542.800 264.400 ;
        RECT 545.200 263.600 546.000 264.400 ;
        RECT 537.200 253.600 538.000 254.400 ;
        RECT 538.900 252.400 539.500 263.600 ;
        RECT 542.100 262.400 542.700 263.600 ;
        RECT 542.000 261.600 542.800 262.400 ;
        RECT 542.100 258.300 542.700 261.600 ;
        RECT 542.100 257.700 544.300 258.300 ;
        RECT 542.000 255.600 542.800 256.400 ;
        RECT 542.100 252.400 542.700 255.600 ;
        RECT 543.700 254.400 544.300 257.700 ;
        RECT 545.300 256.400 545.900 263.600 ;
        RECT 546.900 260.400 547.500 303.600 ;
        RECT 548.400 284.200 549.200 297.800 ;
        RECT 550.000 284.200 550.800 297.800 ;
        RECT 551.600 284.200 552.400 297.800 ;
        RECT 553.200 286.200 554.000 297.800 ;
        RECT 554.900 296.400 555.500 303.600 ;
        RECT 572.400 301.600 573.200 302.400 ;
        RECT 554.800 295.600 555.600 296.400 ;
        RECT 554.800 293.600 555.600 294.400 ;
        RECT 550.000 271.600 550.800 272.400 ;
        RECT 548.400 267.600 549.200 268.400 ;
        RECT 546.800 259.600 547.600 260.400 ;
        RECT 546.800 257.600 547.600 258.400 ;
        RECT 545.200 255.600 546.000 256.400 ;
        RECT 543.600 253.600 544.400 254.400 ;
        RECT 545.200 253.600 546.000 254.400 ;
        RECT 548.400 254.300 549.200 254.400 ;
        RECT 550.100 254.300 550.700 271.600 ;
        RECT 554.900 268.400 555.500 293.600 ;
        RECT 556.400 286.200 557.200 297.800 ;
        RECT 558.000 295.600 558.800 296.400 ;
        RECT 558.100 294.400 558.700 295.600 ;
        RECT 558.000 293.600 558.800 294.400 ;
        RECT 558.000 291.600 558.800 292.400 ;
        RECT 559.600 286.200 560.400 297.800 ;
        RECT 561.200 284.200 562.000 297.800 ;
        RECT 562.800 284.200 563.600 297.800 ;
        RECT 572.500 294.400 573.100 301.600 ;
        RECT 575.700 298.400 576.300 311.600 ;
        RECT 578.800 305.600 579.600 306.400 ;
        RECT 575.600 297.600 576.400 298.400 ;
        RECT 572.400 293.600 573.200 294.400 ;
        RECT 578.900 292.400 579.500 305.600 ;
        RECT 580.500 304.400 581.100 329.700 ;
        RECT 593.200 329.600 594.000 330.400 ;
        RECT 594.800 329.600 595.600 330.400 ;
        RECT 591.600 323.600 592.400 324.400 ;
        RECT 585.200 311.600 586.000 312.400 ;
        RECT 591.700 312.300 592.300 323.600 ;
        RECT 593.200 312.300 594.000 312.400 ;
        RECT 591.700 311.700 594.000 312.300 ;
        RECT 593.200 311.600 594.000 311.700 ;
        RECT 599.700 308.400 600.300 331.600 ;
        RECT 585.200 307.600 586.000 308.400 ;
        RECT 590.000 307.600 590.800 308.400 ;
        RECT 599.600 307.600 600.400 308.400 ;
        RECT 582.000 305.600 582.800 306.400 ;
        RECT 580.400 303.600 581.200 304.400 ;
        RECT 590.100 302.400 590.700 307.600 ;
        RECT 593.200 305.600 594.000 306.400 ;
        RECT 593.200 303.600 594.000 304.400 ;
        RECT 594.800 303.600 595.600 304.400 ;
        RECT 590.000 301.600 590.800 302.400 ;
        RECT 590.000 299.600 590.800 300.400 ;
        RECT 569.200 291.600 570.000 292.400 ;
        RECT 578.800 291.600 579.600 292.400 ;
        RECT 556.400 275.600 557.200 276.400 ;
        RECT 567.600 275.600 568.400 276.400 ;
        RECT 556.500 270.400 557.100 275.600 ;
        RECT 564.400 273.600 565.200 274.400 ;
        RECT 564.500 272.400 565.100 273.600 ;
        RECT 561.200 271.600 562.000 272.400 ;
        RECT 564.400 271.600 565.200 272.400 ;
        RECT 556.400 269.600 557.200 270.400 ;
        RECT 554.800 267.600 555.600 268.400 ;
        RECT 551.600 263.600 552.400 264.400 ;
        RECT 558.000 263.600 558.800 264.400 ;
        RECT 548.400 253.700 550.700 254.300 ;
        RECT 548.400 253.600 549.200 253.700 ;
        RECT 534.000 251.700 536.300 252.300 ;
        RECT 534.000 251.600 534.800 251.700 ;
        RECT 538.800 251.600 539.600 252.400 ;
        RECT 542.000 251.600 542.800 252.400 ;
        RECT 538.800 249.600 539.600 250.400 ;
        RECT 545.300 246.400 545.900 253.600 ;
        RECT 545.200 245.600 546.000 246.400 ;
        RECT 550.100 246.300 550.700 253.700 ;
        RECT 551.700 250.300 552.300 263.600 ;
        RECT 554.800 254.300 555.600 254.400 ;
        RECT 554.800 253.700 557.100 254.300 ;
        RECT 554.800 253.600 555.600 253.700 ;
        RECT 553.200 250.300 554.000 250.400 ;
        RECT 551.700 249.700 554.000 250.300 ;
        RECT 553.200 249.600 554.000 249.700 ;
        RECT 550.100 245.700 552.300 246.300 ;
        RECT 535.600 243.600 536.400 244.400 ;
        RECT 550.000 243.600 550.800 244.400 ;
        RECT 535.700 238.400 536.300 243.600 ;
        RECT 537.200 241.600 538.000 242.400 ;
        RECT 535.600 237.600 536.400 238.400 ;
        RECT 537.300 234.400 537.900 241.600 ;
        RECT 540.400 237.600 541.200 238.400 ;
        RECT 537.200 233.600 538.000 234.400 ;
        RECT 540.500 232.400 541.100 237.600 ;
        RECT 543.600 233.600 544.400 234.400 ;
        RECT 550.100 232.400 550.700 243.600 ;
        RECT 540.400 231.600 541.200 232.400 ;
        RECT 545.200 231.600 546.000 232.400 ;
        RECT 546.800 231.600 547.600 232.400 ;
        RECT 548.400 231.600 549.200 232.400 ;
        RECT 550.000 231.600 550.800 232.400 ;
        RECT 545.300 230.400 545.900 231.600 ;
        RECT 538.800 229.600 539.600 230.400 ;
        RECT 542.000 229.600 542.800 230.400 ;
        RECT 545.200 229.600 546.000 230.400 ;
        RECT 534.000 227.600 534.800 228.400 ;
        RECT 534.100 218.400 534.700 227.600 ;
        RECT 546.900 222.400 547.500 231.600 ;
        RECT 551.700 228.400 552.300 245.700 ;
        RECT 554.800 237.600 555.600 238.400 ;
        RECT 551.600 227.600 552.400 228.400 ;
        RECT 553.200 227.600 554.000 228.400 ;
        RECT 551.700 226.400 552.300 227.600 ;
        RECT 551.600 225.600 552.400 226.400 ;
        RECT 548.400 223.600 549.200 224.400 ;
        RECT 546.800 221.600 547.600 222.400 ;
        RECT 538.800 219.600 539.600 220.400 ;
        RECT 538.900 218.400 539.500 219.600 ;
        RECT 532.400 217.600 533.200 218.400 ;
        RECT 534.000 217.600 534.800 218.400 ;
        RECT 538.800 217.600 539.600 218.400 ;
        RECT 546.900 214.400 547.500 221.600 ;
        RECT 553.300 220.400 553.900 227.600 ;
        RECT 556.500 220.400 557.100 253.700 ;
        RECT 558.100 238.400 558.700 263.600 ;
        RECT 561.300 258.400 561.900 271.600 ;
        RECT 567.700 270.400 568.300 275.600 ;
        RECT 569.300 270.400 569.900 291.600 ;
        RECT 575.600 289.600 576.400 290.400 ;
        RECT 575.700 276.400 576.300 289.600 ;
        RECT 585.200 284.200 586.000 297.800 ;
        RECT 586.800 284.200 587.600 297.800 ;
        RECT 588.400 286.200 589.200 297.800 ;
        RECT 590.100 294.400 590.700 299.600 ;
        RECT 590.000 293.600 590.800 294.400 ;
        RECT 591.600 286.200 592.400 297.800 ;
        RECT 593.300 296.400 593.900 303.600 ;
        RECT 594.900 300.400 595.500 303.600 ;
        RECT 594.800 299.600 595.600 300.400 ;
        RECT 593.200 295.600 594.000 296.400 ;
        RECT 593.300 284.300 593.900 295.600 ;
        RECT 594.800 286.200 595.600 297.800 ;
        RECT 593.300 283.700 595.500 284.300 ;
        RECT 596.400 284.200 597.200 297.800 ;
        RECT 598.000 284.200 598.800 297.800 ;
        RECT 599.600 284.200 600.400 297.800 ;
        RECT 601.300 292.400 601.900 347.600 ;
        RECT 602.800 343.600 603.600 344.400 ;
        RECT 602.900 338.400 603.500 343.600 ;
        RECT 606.100 338.400 606.700 347.600 ;
        RECT 602.800 337.600 603.600 338.400 ;
        RECT 606.000 337.600 606.800 338.400 ;
        RECT 607.700 336.400 608.300 371.600 ;
        RECT 602.800 335.600 603.600 336.400 ;
        RECT 607.600 335.600 608.400 336.400 ;
        RECT 604.400 309.600 605.200 310.400 ;
        RECT 604.500 306.400 605.100 309.600 ;
        RECT 602.800 305.600 603.600 306.400 ;
        RECT 604.400 305.600 605.200 306.400 ;
        RECT 601.200 291.600 602.000 292.400 ;
        RECT 572.400 275.600 573.200 276.400 ;
        RECT 575.600 275.600 576.400 276.400 ;
        RECT 578.800 275.600 579.600 276.400 ;
        RECT 572.500 274.400 573.100 275.600 ;
        RECT 572.400 273.600 573.200 274.400 ;
        RECT 575.600 273.600 576.400 274.400 ;
        RECT 575.700 272.400 576.300 273.600 ;
        RECT 575.600 271.600 576.400 272.400 ;
        RECT 567.600 269.600 568.400 270.400 ;
        RECT 569.200 269.600 570.000 270.400 ;
        RECT 578.800 269.600 579.600 270.400 ;
        RECT 586.800 269.600 587.600 270.400 ;
        RECT 564.400 267.600 565.200 268.400 ;
        RECT 577.200 267.600 578.000 268.400 ;
        RECT 564.400 263.600 565.200 264.400 ;
        RECT 561.200 257.600 562.000 258.400 ;
        RECT 561.300 248.400 561.900 257.600 ;
        RECT 564.500 254.400 565.100 263.600 ;
        RECT 577.200 259.600 578.000 260.400 ;
        RECT 570.800 257.600 571.600 258.400 ;
        RECT 564.400 253.600 565.200 254.400 ;
        RECT 561.200 247.600 562.000 248.400 ;
        RECT 566.000 243.600 566.800 244.400 ;
        RECT 566.100 238.400 566.700 243.600 ;
        RECT 558.000 237.600 558.800 238.400 ;
        RECT 566.000 237.600 566.800 238.400 ;
        RECT 566.000 235.600 566.800 236.400 ;
        RECT 559.600 233.600 560.400 234.400 ;
        RECT 558.000 229.600 558.800 230.400 ;
        RECT 559.700 228.400 560.300 233.600 ;
        RECT 562.800 231.600 563.600 232.400 ;
        RECT 562.800 229.600 563.600 230.400 ;
        RECT 566.100 228.400 566.700 235.600 ;
        RECT 577.300 230.400 577.900 259.600 ;
        RECT 578.900 252.400 579.500 269.600 ;
        RECT 586.800 265.600 587.600 266.400 ;
        RECT 578.800 251.600 579.600 252.400 ;
        RECT 580.400 244.200 581.200 257.800 ;
        RECT 582.000 244.200 582.800 257.800 ;
        RECT 583.600 244.200 584.400 257.800 ;
        RECT 585.200 246.200 586.000 257.800 ;
        RECT 586.900 256.400 587.500 265.600 ;
        RECT 588.400 264.200 589.200 277.800 ;
        RECT 590.000 264.200 590.800 277.800 ;
        RECT 591.600 264.200 592.400 277.800 ;
        RECT 593.200 264.200 594.000 275.800 ;
        RECT 594.900 266.400 595.500 283.700 ;
        RECT 602.900 282.400 603.500 305.600 ;
        RECT 609.200 283.600 610.000 284.400 ;
        RECT 609.300 282.400 609.900 283.600 ;
        RECT 602.800 281.600 603.600 282.400 ;
        RECT 606.000 281.600 606.800 282.400 ;
        RECT 609.200 281.600 610.000 282.400 ;
        RECT 594.800 265.600 595.600 266.400 ;
        RECT 596.400 264.200 597.200 275.800 ;
        RECT 598.000 267.600 598.800 268.400 ;
        RECT 599.600 264.200 600.400 275.800 ;
        RECT 601.200 264.200 602.000 277.800 ;
        RECT 602.800 264.200 603.600 277.800 ;
        RECT 604.400 267.600 605.200 268.400 ;
        RECT 586.800 255.600 587.600 256.400 ;
        RECT 586.900 244.300 587.500 255.600 ;
        RECT 588.400 246.200 589.200 257.800 ;
        RECT 590.000 253.600 590.800 254.400 ;
        RECT 591.600 246.200 592.400 257.800 ;
        RECT 585.300 243.700 587.500 244.300 ;
        RECT 593.200 244.200 594.000 257.800 ;
        RECT 594.800 244.200 595.600 257.800 ;
        RECT 604.500 252.400 605.100 267.600 ;
        RECT 604.400 251.600 605.200 252.400 ;
        RECT 577.200 229.600 578.000 230.400 ;
        RECT 559.600 227.600 560.400 228.400 ;
        RECT 566.000 227.600 566.800 228.400 ;
        RECT 572.400 227.600 573.200 228.400 ;
        RECT 569.200 223.600 570.000 224.400 ;
        RECT 569.300 222.400 569.900 223.600 ;
        RECT 569.200 221.600 570.000 222.400 ;
        RECT 553.200 219.600 554.000 220.400 ;
        RECT 556.400 219.600 557.200 220.400 ;
        RECT 535.600 213.600 536.400 214.400 ;
        RECT 546.800 213.600 547.600 214.400 ;
        RECT 530.800 209.600 531.600 210.400 ;
        RECT 516.400 205.600 517.200 206.400 ;
        RECT 489.200 193.600 490.000 194.400 ;
        RECT 503.600 193.600 504.400 194.400 ;
        RECT 495.600 191.600 496.400 192.400 ;
        RECT 498.800 191.600 499.600 192.400 ;
        RECT 500.400 191.600 501.200 192.400 ;
        RECT 502.000 191.600 502.800 192.400 ;
        RECT 510.000 191.600 510.800 192.400 ;
        RECT 495.700 190.400 496.300 191.600 ;
        RECT 494.000 189.600 494.800 190.400 ;
        RECT 495.600 189.600 496.400 190.400 ;
        RECT 494.100 188.400 494.700 189.600 ;
        RECT 494.000 187.600 494.800 188.400 ;
        RECT 500.500 184.400 501.100 191.600 ;
        RECT 492.400 183.600 493.200 184.400 ;
        RECT 498.800 183.600 499.600 184.400 ;
        RECT 500.400 183.600 501.200 184.400 ;
        RECT 476.400 173.600 477.200 174.400 ;
        RECT 478.000 173.600 478.800 174.400 ;
        RECT 482.800 173.600 483.600 174.400 ;
        RECT 478.100 172.400 478.700 173.600 ;
        RECT 482.900 172.400 483.500 173.600 ;
        RECT 474.800 171.600 475.600 172.400 ;
        RECT 478.000 171.600 478.800 172.400 ;
        RECT 482.800 171.600 483.600 172.400 ;
        RECT 484.400 171.600 485.200 172.400 ;
        RECT 474.800 169.600 475.600 170.400 ;
        RECT 476.400 169.600 477.200 170.400 ;
        RECT 474.800 144.200 475.600 155.800 ;
        RECT 476.500 148.400 477.100 169.600 ;
        RECT 482.900 166.400 483.500 171.600 ;
        RECT 484.500 168.400 485.100 171.600 ;
        RECT 489.200 169.600 490.000 170.400 ;
        RECT 489.300 168.400 489.900 169.600 ;
        RECT 484.400 167.600 485.200 168.400 ;
        RECT 486.000 167.600 486.800 168.400 ;
        RECT 489.200 167.600 490.000 168.400 ;
        RECT 482.800 165.600 483.600 166.400 ;
        RECT 490.800 166.200 491.600 177.800 ;
        RECT 492.500 174.400 493.100 183.600 ;
        RECT 497.200 179.600 498.000 180.400 ;
        RECT 492.400 173.600 493.200 174.400 ;
        RECT 497.300 172.400 497.900 179.600 ;
        RECT 498.900 178.400 499.500 183.600 ;
        RECT 502.100 178.400 502.700 191.600 ;
        RECT 513.200 189.600 514.000 190.400 ;
        RECT 503.600 187.600 504.400 188.400 ;
        RECT 503.700 186.400 504.300 187.600 ;
        RECT 516.500 186.400 517.100 205.600 ;
        RECT 548.400 204.200 549.200 217.800 ;
        RECT 550.000 204.200 550.800 217.800 ;
        RECT 551.600 204.200 552.400 217.800 ;
        RECT 553.200 206.200 554.000 217.800 ;
        RECT 554.800 215.600 555.600 216.400 ;
        RECT 554.900 214.400 555.500 215.600 ;
        RECT 554.800 213.600 555.600 214.400 ;
        RECT 518.000 193.600 518.800 194.400 ;
        RECT 526.000 193.600 526.800 194.400 ;
        RECT 518.100 192.400 518.700 193.600 ;
        RECT 518.000 191.600 518.800 192.400 ;
        RECT 519.600 187.600 520.400 188.400 ;
        RECT 522.800 187.600 523.600 188.400 ;
        RECT 522.900 186.400 523.500 187.600 ;
        RECT 526.100 186.400 526.700 193.600 ;
        RECT 537.200 191.600 538.000 192.400 ;
        RECT 537.300 190.400 537.900 191.600 ;
        RECT 529.200 189.600 530.000 190.400 ;
        RECT 537.200 189.600 538.000 190.400 ;
        RECT 503.600 185.600 504.400 186.400 ;
        RECT 516.400 185.600 517.200 186.400 ;
        RECT 522.800 185.600 523.600 186.400 ;
        RECT 526.000 185.600 526.800 186.400 ;
        RECT 516.500 184.400 517.100 185.600 ;
        RECT 529.300 184.400 529.900 189.600 ;
        RECT 514.800 183.600 515.600 184.400 ;
        RECT 516.400 183.600 517.200 184.400 ;
        RECT 529.200 183.600 530.000 184.400 ;
        RECT 538.800 184.200 539.600 197.800 ;
        RECT 540.400 184.200 541.200 197.800 ;
        RECT 542.000 184.200 542.800 197.800 ;
        RECT 543.600 184.200 544.400 195.800 ;
        RECT 545.200 185.600 546.000 186.400 ;
        RECT 546.800 184.200 547.600 195.800 ;
        RECT 548.400 187.600 549.200 188.400 ;
        RECT 514.900 182.400 515.500 183.600 ;
        RECT 514.800 181.600 515.600 182.400 ;
        RECT 510.000 179.600 510.800 180.400 ;
        RECT 510.100 178.400 510.700 179.600 ;
        RECT 498.800 177.600 499.600 178.400 ;
        RECT 497.200 171.600 498.000 172.400 ;
        RECT 492.400 167.600 493.200 168.400 ;
        RECT 479.600 157.600 480.400 158.400 ;
        RECT 484.400 155.600 485.200 156.400 ;
        RECT 476.400 147.600 477.200 148.400 ;
        RECT 478.000 146.200 478.800 151.800 ;
        RECT 484.500 150.400 485.100 155.600 ;
        RECT 487.600 153.600 488.400 154.400 ;
        RECT 489.200 151.600 490.000 152.400 ;
        RECT 489.300 150.400 489.900 151.600 ;
        RECT 482.800 149.600 483.600 150.400 ;
        RECT 484.400 149.600 485.200 150.400 ;
        RECT 489.200 149.600 490.000 150.400 ;
        RECT 490.800 149.600 491.600 150.400 ;
        RECT 481.200 147.600 482.000 148.400 ;
        RECT 481.300 146.400 481.900 147.600 ;
        RECT 482.900 146.400 483.500 149.600 ;
        RECT 489.300 148.400 489.900 149.600 ;
        RECT 489.200 147.600 490.000 148.400 ;
        RECT 481.200 145.600 482.000 146.400 ;
        RECT 482.800 145.600 483.600 146.400 ;
        RECT 486.000 145.600 486.800 146.400 ;
        RECT 478.000 143.600 478.800 144.400 ;
        RECT 473.200 137.600 474.000 138.400 ;
        RECT 473.200 135.600 474.000 136.400 ;
        RECT 478.100 134.400 478.700 143.600 ;
        RECT 479.600 137.600 480.400 138.400 ;
        RECT 481.200 137.600 482.000 138.400 ;
        RECT 476.400 133.600 477.200 134.400 ;
        RECT 478.000 133.600 478.800 134.400 ;
        RECT 478.100 132.400 478.700 133.600 ;
        RECT 474.800 131.600 475.600 132.400 ;
        RECT 478.000 131.600 478.800 132.400 ;
        RECT 474.900 128.400 475.500 131.600 ;
        RECT 474.800 128.300 475.600 128.400 ;
        RECT 474.800 127.700 477.100 128.300 ;
        RECT 474.800 127.600 475.600 127.700 ;
        RECT 471.600 113.600 472.400 114.400 ;
        RECT 476.500 112.400 477.100 127.700 ;
        RECT 476.400 111.600 477.200 112.400 ;
        RECT 476.500 110.400 477.100 111.600 ;
        RECT 476.400 109.600 477.200 110.400 ;
        RECT 471.600 108.300 472.400 108.400 ;
        RECT 470.100 107.700 472.400 108.300 ;
        RECT 471.600 107.600 472.400 107.700 ;
        RECT 478.000 107.600 478.800 108.400 ;
        RECT 478.100 106.400 478.700 107.600 ;
        RECT 468.400 105.600 469.200 106.400 ;
        RECT 471.600 105.600 472.400 106.400 ;
        RECT 478.000 105.600 478.800 106.400 ;
        RECT 463.600 95.600 464.400 96.400 ;
        RECT 466.800 95.600 467.600 96.400 ;
        RECT 455.600 93.600 456.400 94.400 ;
        RECT 458.800 93.600 459.600 94.400 ;
        RECT 455.600 91.600 456.400 92.400 ;
        RECT 455.700 90.400 456.300 91.600 ;
        RECT 455.600 89.600 456.400 90.400 ;
        RECT 457.200 89.600 458.000 90.400 ;
        RECT 458.900 86.400 459.500 93.600 ;
        RECT 466.900 92.400 467.500 95.600 ;
        RECT 471.700 92.400 472.300 105.600 ;
        RECT 474.800 103.600 475.600 104.400 ;
        RECT 473.200 93.600 474.000 94.400 ;
        RECT 474.900 92.400 475.500 103.600 ;
        RECT 476.400 95.600 477.200 96.400 ;
        RECT 465.200 91.600 466.000 92.400 ;
        RECT 466.800 91.600 467.600 92.400 ;
        RECT 471.600 91.600 472.400 92.400 ;
        RECT 474.800 91.600 475.600 92.400 ;
        RECT 458.800 85.600 459.600 86.400 ;
        RECT 455.600 75.600 456.400 76.400 ;
        RECT 457.200 75.600 458.000 76.400 ;
        RECT 457.300 70.400 457.900 75.600 ;
        RECT 463.600 73.600 464.400 74.400 ;
        RECT 457.200 69.600 458.000 70.400 ;
        RECT 458.800 67.600 459.600 68.400 ;
        RECT 454.000 65.600 454.800 66.400 ;
        RECT 458.900 58.400 459.500 67.600 ;
        RECT 458.800 57.600 459.600 58.400 ;
        RECT 452.400 55.600 453.200 56.400 ;
        RECT 455.600 55.600 456.400 56.400 ;
        RECT 450.800 53.600 451.600 54.400 ;
        RECT 455.700 52.400 456.300 55.600 ;
        RECT 465.300 52.400 465.900 91.600 ;
        RECT 470.000 83.600 470.800 84.400 ;
        RECT 466.800 65.600 467.600 66.400 ;
        RECT 466.900 52.400 467.500 65.600 ;
        RECT 468.400 64.200 469.200 75.800 ;
        RECT 470.100 72.400 470.700 83.600 ;
        RECT 471.700 74.400 472.300 91.600 ;
        RECT 476.500 90.400 477.100 95.600 ;
        RECT 476.400 89.600 477.200 90.400 ;
        RECT 478.100 84.400 478.700 105.600 ;
        RECT 479.700 92.400 480.300 137.600 ;
        RECT 481.300 130.400 481.900 137.600 ;
        RECT 482.800 133.600 483.600 134.400 ;
        RECT 484.400 133.600 485.200 134.400 ;
        RECT 482.800 132.300 483.600 132.400 ;
        RECT 484.500 132.300 485.100 133.600 ;
        RECT 482.800 131.700 485.100 132.300 ;
        RECT 482.800 131.600 483.600 131.700 ;
        RECT 481.200 129.600 482.000 130.400 ;
        RECT 484.400 129.600 485.200 130.400 ;
        RECT 481.200 121.600 482.000 122.400 ;
        RECT 481.300 118.400 481.900 121.600 ;
        RECT 481.200 117.600 482.000 118.400 ;
        RECT 482.800 111.600 483.600 112.400 ;
        RECT 482.900 110.400 483.500 111.600 ;
        RECT 481.200 109.600 482.000 110.400 ;
        RECT 482.800 109.600 483.600 110.400 ;
        RECT 482.800 103.600 483.600 104.400 ;
        RECT 482.900 100.400 483.500 103.600 ;
        RECT 482.800 99.600 483.600 100.400 ;
        RECT 484.500 92.400 485.100 129.600 ;
        RECT 486.100 110.400 486.700 145.600 ;
        RECT 489.200 133.600 490.000 134.400 ;
        RECT 487.600 131.600 488.400 132.400 ;
        RECT 487.700 130.400 488.300 131.600 ;
        RECT 489.300 130.400 489.900 133.600 ;
        RECT 487.600 129.600 488.400 130.400 ;
        RECT 489.200 129.600 490.000 130.400 ;
        RECT 487.600 119.600 488.400 120.400 ;
        RECT 486.000 109.600 486.800 110.400 ;
        RECT 486.100 102.400 486.700 109.600 ;
        RECT 487.700 108.400 488.300 119.600 ;
        RECT 489.200 117.600 490.000 118.400 ;
        RECT 489.300 112.400 489.900 117.600 ;
        RECT 489.200 111.600 490.000 112.400 ;
        RECT 489.200 109.600 490.000 110.400 ;
        RECT 490.900 110.300 491.500 149.600 ;
        RECT 492.500 148.400 493.100 167.600 ;
        RECT 495.600 151.600 496.400 152.400 ;
        RECT 492.400 147.600 493.200 148.400 ;
        RECT 494.000 133.600 494.800 134.400 ;
        RECT 494.100 132.400 494.700 133.600 ;
        RECT 494.000 131.600 494.800 132.400 ;
        RECT 492.400 129.600 493.200 130.400 ;
        RECT 495.700 118.400 496.300 151.600 ;
        RECT 497.200 143.600 498.000 144.400 ;
        RECT 497.300 142.400 497.900 143.600 ;
        RECT 497.200 141.600 498.000 142.400 ;
        RECT 497.200 132.300 498.000 132.400 ;
        RECT 498.900 132.300 499.500 177.600 ;
        RECT 500.400 166.200 501.200 177.800 ;
        RECT 502.000 177.600 502.800 178.400 ;
        RECT 510.000 177.600 510.800 178.400 ;
        RECT 502.000 173.600 502.800 174.400 ;
        RECT 502.100 166.400 502.700 173.600 ;
        RECT 503.600 170.200 504.400 175.800 ;
        RECT 521.200 175.600 522.000 176.400 ;
        RECT 521.300 174.400 521.900 175.600 ;
        RECT 529.300 174.400 529.900 183.600 ;
        RECT 548.500 182.300 549.100 187.600 ;
        RECT 550.000 184.200 550.800 195.800 ;
        RECT 551.600 184.200 552.400 197.800 ;
        RECT 553.200 184.200 554.000 197.800 ;
        RECT 554.900 186.400 555.500 213.600 ;
        RECT 556.400 206.200 557.200 217.800 ;
        RECT 558.000 217.600 558.800 218.400 ;
        RECT 558.100 214.400 558.700 217.600 ;
        RECT 558.000 213.600 558.800 214.400 ;
        RECT 559.600 206.200 560.400 217.800 ;
        RECT 561.200 204.200 562.000 217.800 ;
        RECT 562.800 204.200 563.600 217.800 ;
        RECT 567.600 215.600 568.400 216.400 ;
        RECT 567.700 212.400 568.300 215.600 ;
        RECT 572.500 214.400 573.100 227.600 ;
        RECT 572.400 213.600 573.200 214.400 ;
        RECT 567.600 211.600 568.400 212.400 ;
        RECT 572.500 204.400 573.100 213.600 ;
        RECT 577.300 212.400 577.900 229.600 ;
        RECT 578.800 224.200 579.600 237.800 ;
        RECT 580.400 224.200 581.200 237.800 ;
        RECT 582.000 224.200 582.800 237.800 ;
        RECT 583.600 224.200 584.400 235.800 ;
        RECT 585.300 226.400 585.900 243.700 ;
        RECT 588.400 237.600 589.200 238.400 ;
        RECT 585.200 225.600 586.000 226.400 ;
        RECT 586.800 224.200 587.600 235.800 ;
        RECT 588.500 228.400 589.100 237.600 ;
        RECT 588.400 227.600 589.200 228.400 ;
        RECT 590.000 224.200 590.800 235.800 ;
        RECT 591.600 224.200 592.400 237.800 ;
        RECT 593.200 224.200 594.000 237.800 ;
        RECT 604.500 234.400 605.100 251.600 ;
        RECT 596.400 233.600 597.200 234.400 ;
        RECT 604.400 233.600 605.200 234.400 ;
        RECT 591.600 219.600 592.400 220.400 ;
        RECT 591.700 214.400 592.300 219.600 ;
        RECT 578.800 213.600 579.600 214.400 ;
        RECT 591.600 213.600 592.400 214.400 ;
        RECT 574.000 211.600 574.800 212.400 ;
        RECT 575.600 211.600 576.400 212.400 ;
        RECT 577.200 211.600 578.000 212.400 ;
        RECT 574.100 210.400 574.700 211.600 ;
        RECT 574.000 209.600 574.800 210.400 ;
        RECT 572.400 203.600 573.200 204.400 ;
        RECT 559.600 189.600 560.400 190.400 ;
        RECT 566.000 189.600 566.800 190.400 ;
        RECT 554.800 185.600 555.600 186.400 ;
        RECT 548.500 181.700 550.700 182.300 ;
        RECT 550.100 178.400 550.700 181.700 ;
        RECT 554.900 180.300 555.500 185.600 ;
        RECT 553.300 179.700 555.500 180.300 ;
        RECT 550.000 177.600 550.800 178.400 ;
        RECT 545.200 175.600 546.000 176.400 ;
        RECT 551.600 175.600 552.400 176.400 ;
        RECT 505.200 173.600 506.000 174.400 ;
        RECT 506.800 173.600 507.600 174.400 ;
        RECT 516.400 173.600 517.200 174.400 ;
        RECT 521.200 173.600 522.000 174.400 ;
        RECT 529.200 173.600 530.000 174.400 ;
        RECT 537.200 173.600 538.000 174.400 ;
        RECT 543.600 173.600 544.400 174.400 ;
        RECT 505.300 170.300 505.900 173.600 ;
        RECT 506.900 172.400 507.500 173.600 ;
        RECT 506.800 171.600 507.600 172.400 ;
        RECT 514.800 172.300 515.600 172.400 ;
        RECT 513.300 171.700 515.600 172.300 ;
        RECT 505.300 169.700 507.500 170.300 ;
        RECT 502.000 165.600 502.800 166.400 ;
        RECT 506.900 160.400 507.500 169.700 ;
        RECT 511.600 169.600 512.400 170.400 ;
        RECT 513.300 160.400 513.900 171.700 ;
        RECT 514.800 171.600 515.600 171.700 ;
        RECT 516.500 170.300 517.100 173.600 ;
        RECT 537.300 172.400 537.900 173.600 ;
        RECT 518.000 171.600 518.800 172.400 ;
        RECT 519.600 171.600 520.400 172.400 ;
        RECT 524.400 171.600 525.200 172.400 ;
        RECT 527.600 171.600 528.400 172.400 ;
        RECT 529.200 171.600 530.000 172.400 ;
        RECT 534.000 171.600 534.800 172.400 ;
        RECT 537.200 171.600 538.000 172.400 ;
        RECT 538.800 171.600 539.600 172.400 ;
        RECT 540.400 171.600 541.200 172.400 ;
        RECT 514.900 169.700 517.100 170.300 ;
        RECT 506.800 159.600 507.600 160.400 ;
        RECT 513.200 159.600 514.000 160.400 ;
        RECT 505.200 153.600 506.000 154.400 ;
        RECT 505.300 150.400 505.900 153.600 ;
        RECT 500.400 149.600 501.200 150.400 ;
        RECT 505.200 149.600 506.000 150.400 ;
        RECT 500.500 146.400 501.100 149.600 ;
        RECT 506.900 148.400 507.500 159.600 ;
        RECT 510.000 151.600 510.800 152.400 ;
        RECT 513.300 150.400 513.900 159.600 ;
        RECT 508.400 149.600 509.200 150.400 ;
        RECT 513.200 149.600 514.000 150.400 ;
        RECT 508.500 148.400 509.100 149.600 ;
        RECT 514.900 148.400 515.500 169.700 ;
        RECT 518.100 158.400 518.700 171.600 ;
        RECT 519.700 170.400 520.300 171.600 ;
        RECT 524.500 170.400 525.100 171.600 ;
        RECT 519.600 169.600 520.400 170.400 ;
        RECT 524.400 169.600 525.200 170.400 ;
        RECT 519.600 165.600 520.400 166.400 ;
        RECT 518.000 157.600 518.800 158.400 ;
        RECT 519.700 154.400 520.300 165.600 ;
        RECT 524.500 156.400 525.100 169.600 ;
        RECT 529.300 168.400 529.900 171.600 ;
        RECT 534.100 170.400 534.700 171.600 ;
        RECT 534.000 169.600 534.800 170.400 ;
        RECT 529.200 167.600 530.000 168.400 ;
        RECT 529.300 164.400 529.900 167.600 ;
        RECT 529.200 163.600 530.000 164.400 ;
        RECT 532.400 163.600 533.200 164.400 ;
        RECT 516.400 153.600 517.200 154.400 ;
        RECT 519.600 153.600 520.400 154.400 ;
        RECT 516.500 152.400 517.100 153.600 ;
        RECT 516.400 151.600 517.200 152.400 ;
        RECT 502.000 147.600 502.800 148.400 ;
        RECT 503.600 147.600 504.400 148.400 ;
        RECT 506.800 147.600 507.600 148.400 ;
        RECT 508.400 147.600 509.200 148.400 ;
        RECT 514.800 147.600 515.600 148.400 ;
        RECT 500.400 145.600 501.200 146.400 ;
        RECT 502.100 140.400 502.700 147.600 ;
        RECT 502.000 139.600 502.800 140.400 ;
        RECT 506.900 138.400 507.500 147.600 ;
        RECT 502.000 137.600 502.800 138.400 ;
        RECT 506.800 137.600 507.600 138.400 ;
        RECT 502.100 132.400 502.700 137.600 ;
        RECT 514.900 136.400 515.500 147.600 ;
        RECT 521.200 144.200 522.000 155.800 ;
        RECT 524.400 155.600 525.200 156.400 ;
        RECT 527.600 149.600 528.400 150.400 ;
        RECT 524.400 145.600 525.200 146.400 ;
        RECT 529.200 145.600 530.000 146.400 ;
        RECT 518.000 137.600 518.800 138.400 ;
        RECT 513.200 135.600 514.000 136.400 ;
        RECT 514.800 135.600 515.600 136.400 ;
        RECT 508.400 133.600 509.200 134.400 ;
        RECT 511.600 133.600 512.400 134.400 ;
        RECT 497.200 131.700 499.500 132.300 ;
        RECT 497.200 131.600 498.000 131.700 ;
        RECT 502.000 131.600 502.800 132.400 ;
        RECT 503.600 131.600 504.400 132.400 ;
        RECT 503.700 122.400 504.300 131.600 ;
        RECT 506.800 125.600 507.600 126.400 ;
        RECT 503.600 121.600 504.400 122.400 ;
        RECT 505.200 119.600 506.000 120.400 ;
        RECT 505.300 118.400 505.900 119.600 ;
        RECT 495.600 117.600 496.400 118.400 ;
        RECT 505.200 117.600 506.000 118.400 ;
        RECT 503.600 115.600 504.400 116.400 ;
        RECT 503.700 114.400 504.300 115.600 ;
        RECT 503.600 113.600 504.400 114.400 ;
        RECT 506.900 110.400 507.500 125.600 ;
        RECT 492.400 110.300 493.200 110.400 ;
        RECT 490.900 109.700 493.200 110.300 ;
        RECT 492.400 109.600 493.200 109.700 ;
        RECT 503.600 109.600 504.400 110.400 ;
        RECT 506.800 109.600 507.600 110.400 ;
        RECT 487.600 107.600 488.400 108.400 ;
        RECT 490.800 107.600 491.600 108.400 ;
        RECT 492.400 107.600 493.200 108.400 ;
        RECT 494.000 107.600 494.800 108.400 ;
        RECT 500.400 107.600 501.200 108.400 ;
        RECT 486.000 101.600 486.800 102.400 ;
        RECT 490.900 94.400 491.500 107.600 ;
        RECT 490.800 93.600 491.600 94.400 ;
        RECT 492.500 92.400 493.100 107.600 ;
        RECT 498.800 103.600 499.600 104.400 ;
        RECT 495.600 99.600 496.400 100.400 ;
        RECT 479.600 91.600 480.400 92.400 ;
        RECT 484.400 91.600 485.200 92.400 ;
        RECT 490.800 91.600 491.600 92.400 ;
        RECT 492.400 91.600 493.200 92.400 ;
        RECT 495.700 90.400 496.300 99.600 ;
        RECT 497.200 97.600 498.000 98.400 ;
        RECT 497.300 92.400 497.900 97.600 ;
        RECT 498.900 94.300 499.500 103.600 ;
        RECT 503.700 94.400 504.300 109.600 ;
        RECT 508.500 108.400 509.100 133.600 ;
        RECT 513.300 132.400 513.900 135.600 ;
        RECT 510.000 131.600 510.800 132.400 ;
        RECT 513.200 131.600 514.000 132.400 ;
        RECT 514.800 131.600 515.600 132.400 ;
        RECT 510.100 122.400 510.700 131.600 ;
        RECT 510.000 121.600 510.800 122.400 ;
        RECT 510.000 111.600 510.800 112.400 ;
        RECT 513.200 111.600 514.000 112.400 ;
        RECT 508.400 107.600 509.200 108.400 ;
        RECT 511.600 107.600 512.400 108.400 ;
        RECT 513.300 108.300 513.900 111.600 ;
        RECT 514.900 110.400 515.500 131.600 ;
        RECT 516.400 129.600 517.200 130.400 ;
        RECT 514.800 109.600 515.600 110.400 ;
        RECT 513.300 107.700 515.500 108.300 ;
        RECT 506.800 105.600 507.600 106.400 ;
        RECT 508.400 101.600 509.200 102.400 ;
        RECT 506.800 97.600 507.600 98.400 ;
        RECT 498.900 93.700 501.100 94.300 ;
        RECT 497.200 91.600 498.000 92.400 ;
        RECT 498.800 91.600 499.600 92.400 ;
        RECT 495.600 89.600 496.400 90.400 ;
        RECT 478.000 83.600 478.800 84.400 ;
        RECT 479.600 83.600 480.400 84.400 ;
        RECT 487.600 83.600 488.400 84.400 ;
        RECT 492.400 83.600 493.200 84.400 ;
        RECT 471.600 73.600 472.400 74.400 ;
        RECT 470.000 71.600 470.800 72.400 ;
        RECT 474.800 69.600 475.600 70.400 ;
        RECT 473.200 67.600 474.000 68.400 ;
        RECT 473.300 62.400 473.900 67.600 ;
        RECT 478.000 64.200 478.800 75.800 ;
        RECT 479.700 70.400 480.300 83.600 ;
        RECT 479.600 69.600 480.400 70.400 ;
        RECT 473.200 61.600 474.000 62.400 ;
        RECT 479.700 60.400 480.300 69.600 ;
        RECT 481.200 66.200 482.000 71.800 ;
        RECT 484.400 71.600 485.200 72.400 ;
        RECT 484.500 70.400 485.100 71.600 ;
        RECT 484.400 69.600 485.200 70.400 ;
        RECT 482.800 67.600 483.600 68.400 ;
        RECT 487.700 66.300 488.300 83.600 ;
        RECT 492.500 80.400 493.100 83.600 ;
        RECT 492.400 79.600 493.200 80.400 ;
        RECT 489.200 73.600 490.000 74.400 ;
        RECT 489.300 72.400 489.900 73.600 ;
        RECT 489.200 71.600 490.000 72.400 ;
        RECT 489.300 68.400 489.900 71.600 ;
        RECT 492.400 69.600 493.200 70.400 ;
        RECT 489.200 67.600 490.000 68.400 ;
        RECT 494.000 67.600 494.800 68.400 ;
        RECT 487.700 65.700 489.900 66.300 ;
        RECT 487.600 63.600 488.400 64.400 ;
        RECT 484.400 61.600 485.200 62.400 ;
        RECT 479.600 59.600 480.400 60.400 ;
        RECT 471.600 55.600 472.400 56.400 ;
        RECT 476.400 55.600 477.200 56.400 ;
        RECT 479.600 55.600 480.400 56.400 ;
        RECT 446.000 51.600 446.800 52.400 ;
        RECT 447.600 51.600 448.400 52.400 ;
        RECT 449.200 52.300 450.000 52.400 ;
        RECT 449.200 51.700 451.500 52.300 ;
        RECT 449.200 51.600 450.000 51.700 ;
        RECT 447.700 50.400 448.300 51.600 ;
        RECT 442.800 49.600 443.600 50.400 ;
        RECT 444.400 49.600 445.200 50.400 ;
        RECT 447.600 49.600 448.400 50.400 ;
        RECT 444.400 47.600 445.200 48.400 ;
        RECT 444.500 38.400 445.100 47.600 ;
        RECT 444.400 37.600 445.200 38.400 ;
        RECT 442.800 33.600 443.600 34.400 ;
        RECT 447.600 31.600 448.400 32.400 ;
        RECT 444.400 29.600 445.200 30.400 ;
        RECT 439.600 27.700 441.900 28.300 ;
        RECT 439.600 27.600 440.400 27.700 ;
        RECT 446.000 27.600 446.800 28.400 ;
        RECT 422.000 7.600 422.800 8.400 ;
        RECT 425.200 7.600 426.000 8.400 ;
        RECT 434.800 7.600 435.600 8.400 ;
        RECT 438.000 6.200 438.800 17.800 ;
        RECT 446.100 16.400 446.700 27.600 ;
        RECT 447.700 20.400 448.300 31.600 ;
        RECT 450.900 30.400 451.500 51.700 ;
        RECT 455.600 51.600 456.400 52.400 ;
        RECT 463.600 52.300 464.400 52.400 ;
        RECT 465.200 52.300 466.000 52.400 ;
        RECT 463.600 51.700 466.000 52.300 ;
        RECT 463.600 51.600 464.400 51.700 ;
        RECT 465.200 51.600 466.000 51.700 ;
        RECT 466.800 51.600 467.600 52.400 ;
        RECT 473.200 51.600 474.000 52.400 ;
        RECT 474.800 51.600 475.600 52.400 ;
        RECT 455.700 44.400 456.300 51.600 ;
        RECT 474.900 50.400 475.500 51.600 ;
        RECT 463.600 49.600 464.400 50.400 ;
        RECT 474.800 50.300 475.600 50.400 ;
        RECT 473.300 49.700 475.600 50.300 ;
        RECT 463.700 48.400 464.300 49.600 ;
        RECT 463.600 47.600 464.400 48.400 ;
        RECT 455.600 43.600 456.400 44.400 ;
        RECT 450.800 29.600 451.600 30.400 ;
        RECT 449.200 27.600 450.000 28.400 ;
        RECT 452.400 27.600 453.200 28.400 ;
        RECT 447.600 19.600 448.400 20.400 ;
        RECT 446.000 15.600 446.800 16.400 ;
        RECT 446.000 13.600 446.800 14.400 ;
        RECT 446.100 12.600 446.700 13.600 ;
        RECT 446.000 11.800 446.800 12.600 ;
        RECT 447.600 6.200 448.400 17.800 ;
        RECT 449.300 10.400 449.900 27.600 ;
        RECT 452.500 24.400 453.100 27.600 ;
        RECT 457.200 25.600 458.000 26.400 ;
        RECT 458.800 26.200 459.600 31.800 ;
        RECT 452.400 23.600 453.200 24.400 ;
        RECT 449.200 9.600 450.000 10.400 ;
        RECT 450.800 10.200 451.600 15.800 ;
        RECT 457.300 14.400 457.900 25.600 ;
        RECT 462.000 24.200 462.800 35.800 ;
        RECT 465.200 29.600 466.000 30.400 ;
        RECT 470.000 29.600 470.800 30.400 ;
        RECT 470.100 28.400 470.700 29.600 ;
        RECT 470.000 27.600 470.800 28.400 ;
        RECT 471.600 24.200 472.400 35.800 ;
        RECT 463.600 21.600 464.400 22.400 ;
        RECT 452.400 13.600 453.200 14.400 ;
        RECT 455.600 13.600 456.400 14.400 ;
        RECT 457.200 13.600 458.000 14.400 ;
        RECT 455.700 12.400 456.300 13.600 ;
        RECT 463.700 12.400 464.300 21.600 ;
        RECT 465.200 19.600 466.000 20.400 ;
        RECT 465.300 12.400 465.900 19.600 ;
        RECT 466.800 15.600 467.600 16.400 ;
        RECT 466.900 14.400 467.500 15.600 ;
        RECT 466.800 13.600 467.600 14.400 ;
        RECT 473.300 12.400 473.900 49.700 ;
        RECT 474.800 49.600 475.600 49.700 ;
        RECT 474.800 43.600 475.600 44.400 ;
        RECT 474.900 12.400 475.500 43.600 ;
        RECT 476.500 38.400 477.100 55.600 ;
        RECT 479.700 52.400 480.300 55.600 ;
        RECT 479.600 51.600 480.400 52.400 ;
        RECT 482.800 50.200 483.600 55.800 ;
        RECT 484.500 54.400 485.100 61.600 ;
        RECT 484.400 53.600 485.200 54.400 ;
        RECT 486.000 46.200 486.800 57.800 ;
        RECT 487.700 52.600 488.300 63.600 ;
        RECT 487.600 51.800 488.400 52.600 ;
        RECT 478.000 43.600 478.800 44.400 ;
        RECT 476.400 37.600 477.200 38.400 ;
        RECT 476.500 32.400 477.100 37.600 ;
        RECT 476.400 31.600 477.200 32.400 ;
        RECT 478.100 30.400 478.700 43.600 ;
        RECT 484.400 31.600 485.200 32.400 ;
        RECT 489.300 30.400 489.900 65.700 ;
        RECT 494.100 54.400 494.700 67.600 ;
        RECT 494.000 53.600 494.800 54.400 ;
        RECT 495.600 46.200 496.400 57.800 ;
        RECT 497.300 52.400 497.900 91.600 ;
        RECT 498.900 76.400 499.500 91.600 ;
        RECT 500.500 82.400 501.100 93.700 ;
        RECT 503.600 93.600 504.400 94.400 ;
        RECT 503.700 92.400 504.300 93.600 ;
        RECT 506.900 92.400 507.500 97.600 ;
        RECT 503.600 91.600 504.400 92.400 ;
        RECT 506.800 91.600 507.600 92.400 ;
        RECT 502.000 83.600 502.800 84.400 ;
        RECT 500.400 81.600 501.200 82.400 ;
        RECT 498.800 75.600 499.600 76.400 ;
        RECT 498.900 72.300 499.500 75.600 ;
        RECT 500.400 72.300 501.200 72.400 ;
        RECT 498.900 71.700 501.200 72.300 ;
        RECT 500.400 71.600 501.200 71.700 ;
        RECT 502.100 70.400 502.700 83.600 ;
        RECT 506.900 78.400 507.500 91.600 ;
        RECT 506.800 77.600 507.600 78.400 ;
        RECT 505.200 71.600 506.000 72.400 ;
        RECT 508.500 70.400 509.100 101.600 ;
        RECT 510.000 95.600 510.800 96.400 ;
        RECT 511.700 94.400 512.300 107.600 ;
        RECT 514.900 104.400 515.500 107.700 ;
        RECT 513.200 103.600 514.000 104.400 ;
        RECT 514.800 103.600 515.600 104.400 ;
        RECT 511.600 93.600 512.400 94.400 ;
        RECT 513.300 88.400 513.900 103.600 ;
        RECT 516.500 98.400 517.100 129.600 ;
        RECT 522.800 126.200 523.600 137.800 ;
        RECT 522.800 123.600 523.600 124.400 ;
        RECT 522.900 114.400 523.500 123.600 ;
        RECT 522.800 113.600 523.600 114.400 ;
        RECT 521.200 111.600 522.000 112.400 ;
        RECT 521.300 110.400 521.900 111.600 ;
        RECT 522.900 110.400 523.500 113.600 ;
        RECT 518.000 109.600 518.800 110.400 ;
        RECT 521.200 109.600 522.000 110.400 ;
        RECT 522.800 109.600 523.600 110.400 ;
        RECT 521.300 106.400 521.900 109.600 ;
        RECT 521.200 105.600 522.000 106.400 ;
        RECT 521.200 101.600 522.000 102.400 ;
        RECT 516.400 97.600 517.200 98.400 ;
        RECT 518.000 91.600 518.800 92.400 ;
        RECT 519.600 91.600 520.400 92.400 ;
        RECT 513.200 87.600 514.000 88.400 ;
        RECT 516.400 87.600 517.200 88.400 ;
        RECT 511.600 79.600 512.400 80.400 ;
        RECT 502.000 69.600 502.800 70.400 ;
        RECT 505.200 69.600 506.000 70.400 ;
        RECT 508.400 69.600 509.200 70.400 ;
        RECT 500.400 67.600 501.200 68.400 ;
        RECT 503.600 67.600 504.400 68.400 ;
        RECT 506.800 67.600 507.600 68.400 ;
        RECT 508.400 67.600 509.200 68.400 ;
        RECT 500.500 58.400 501.100 67.600 ;
        RECT 503.700 58.400 504.300 67.600 ;
        RECT 506.900 66.300 507.500 67.600 ;
        RECT 506.900 65.700 509.100 66.300 ;
        RECT 500.400 57.600 501.200 58.400 ;
        RECT 503.600 57.600 504.400 58.400 ;
        RECT 502.000 55.600 502.800 56.400 ;
        RECT 497.200 51.600 498.000 52.400 ;
        RECT 502.100 40.400 502.700 55.600 ;
        RECT 505.200 51.600 506.000 52.400 ;
        RECT 506.800 51.600 507.600 52.400 ;
        RECT 502.000 39.600 502.800 40.400 ;
        RECT 506.900 38.300 507.500 51.600 ;
        RECT 508.500 40.400 509.100 65.700 ;
        RECT 511.700 52.400 512.300 79.600 ;
        RECT 514.800 75.600 515.600 76.400 ;
        RECT 513.200 71.600 514.000 72.400 ;
        RECT 513.300 66.400 513.900 71.600 ;
        RECT 513.200 65.600 514.000 66.400 ;
        RECT 513.200 63.600 514.000 64.400 ;
        RECT 516.500 58.400 517.100 87.600 ;
        RECT 516.400 57.600 517.200 58.400 ;
        RECT 516.400 53.600 517.200 54.400 ;
        RECT 511.600 51.600 512.400 52.400 ;
        RECT 514.800 51.600 515.600 52.400 ;
        RECT 511.700 50.400 512.300 51.600 ;
        RECT 511.600 49.600 512.400 50.400 ;
        RECT 510.000 43.600 510.800 44.400 ;
        RECT 508.400 39.600 509.200 40.400 ;
        RECT 508.400 38.300 509.200 38.400 ;
        RECT 506.900 37.700 509.200 38.300 ;
        RECT 508.400 37.600 509.200 37.700 ;
        RECT 478.000 29.600 478.800 30.400 ;
        RECT 481.200 29.600 482.000 30.400 ;
        RECT 489.200 29.600 490.000 30.400 ;
        RECT 478.000 27.600 478.800 28.400 ;
        RECT 489.200 27.600 490.000 28.400 ;
        RECT 478.100 26.400 478.700 27.600 ;
        RECT 478.000 25.600 478.800 26.400 ;
        RECT 482.800 25.600 483.600 26.400 ;
        RECT 478.000 15.600 478.800 16.400 ;
        RECT 478.100 14.400 478.700 15.600 ;
        RECT 482.900 14.400 483.500 25.600 ;
        RECT 489.300 24.400 489.900 27.600 ;
        RECT 490.800 26.200 491.600 31.800 ;
        RECT 492.400 29.600 493.200 30.400 ;
        RECT 489.200 23.600 490.000 24.400 ;
        RECT 489.300 14.400 489.900 23.600 ;
        RECT 478.000 13.600 478.800 14.400 ;
        RECT 482.800 13.600 483.600 14.400 ;
        RECT 484.400 13.600 485.200 14.400 ;
        RECT 487.600 13.600 488.400 14.400 ;
        RECT 489.200 13.600 490.000 14.400 ;
        RECT 484.500 12.400 485.100 13.600 ;
        RECT 455.600 11.600 456.400 12.400 ;
        RECT 463.600 11.600 464.400 12.400 ;
        RECT 465.200 11.600 466.000 12.400 ;
        RECT 473.200 11.600 474.000 12.400 ;
        RECT 474.800 11.600 475.600 12.400 ;
        RECT 479.600 11.600 480.400 12.400 ;
        RECT 481.200 11.600 482.000 12.400 ;
        RECT 484.400 11.600 485.200 12.400 ;
        RECT 479.700 10.400 480.300 11.600 ;
        RECT 452.400 9.600 453.200 10.400 ;
        RECT 479.600 9.600 480.400 10.400 ;
        RECT 487.700 8.400 488.300 13.600 ;
        RECT 492.500 12.400 493.100 29.600 ;
        RECT 494.000 24.200 494.800 35.800 ;
        RECT 497.200 29.600 498.000 30.400 ;
        RECT 502.000 29.600 502.800 30.400 ;
        RECT 502.100 28.400 502.700 29.600 ;
        RECT 502.000 27.600 502.800 28.400 ;
        RECT 494.000 13.600 494.800 14.400 ;
        RECT 492.400 11.600 493.200 12.400 ;
        RECT 489.200 9.600 490.000 10.400 ;
        RECT 495.600 10.200 496.400 15.800 ;
        RECT 487.600 7.600 488.400 8.400 ;
        RECT 498.800 6.200 499.600 17.800 ;
        RECT 502.100 14.400 502.700 27.600 ;
        RECT 503.600 24.200 504.400 35.800 ;
        RECT 508.500 34.400 509.100 37.600 ;
        RECT 508.400 33.600 509.200 34.400 ;
        RECT 510.100 30.400 510.700 43.600 ;
        RECT 510.000 29.600 510.800 30.400 ;
        RECT 513.200 29.600 514.000 30.400 ;
        RECT 510.000 27.600 510.800 28.400 ;
        RECT 510.100 26.400 510.700 27.600 ;
        RECT 510.000 25.600 510.800 26.400 ;
        RECT 502.000 13.600 502.800 14.400 ;
        RECT 500.400 11.800 501.200 12.600 ;
        RECT 500.500 8.400 501.100 11.800 ;
        RECT 500.400 7.600 501.200 8.400 ;
        RECT 508.400 6.200 509.200 17.800 ;
        RECT 514.900 12.400 515.500 51.600 ;
        RECT 516.400 33.600 517.200 34.400 ;
        RECT 516.500 32.400 517.100 33.600 ;
        RECT 516.400 31.600 517.200 32.400 ;
        RECT 518.100 12.400 518.700 91.600 ;
        RECT 519.700 90.400 520.300 91.600 ;
        RECT 519.600 89.600 520.400 90.400 ;
        RECT 519.600 64.200 520.400 75.800 ;
        RECT 521.300 52.400 521.900 101.600 ;
        RECT 522.900 92.400 523.500 109.600 ;
        RECT 524.500 108.400 525.100 145.600 ;
        RECT 529.300 134.400 529.900 145.600 ;
        RECT 530.800 144.200 531.600 155.800 ;
        RECT 532.500 150.400 533.100 163.600 ;
        RECT 538.900 160.400 539.500 171.600 ;
        RECT 538.800 159.600 539.600 160.400 ;
        RECT 540.500 152.400 541.100 171.600 ;
        RECT 542.000 169.600 542.800 170.400 ;
        RECT 542.100 168.400 542.700 169.600 ;
        RECT 542.000 167.600 542.800 168.400 ;
        RECT 542.100 158.400 542.700 167.600 ;
        RECT 542.000 157.600 542.800 158.400 ;
        RECT 532.400 149.600 533.200 150.400 ;
        RECT 532.400 147.600 533.200 148.400 ;
        RECT 534.000 146.200 534.800 151.800 ;
        RECT 540.400 151.600 541.200 152.400 ;
        RECT 537.200 149.600 538.000 150.400 ;
        RECT 540.400 149.600 541.200 150.400 ;
        RECT 535.600 147.600 536.400 148.400 ;
        RECT 535.700 146.400 536.300 147.600 ;
        RECT 535.600 145.600 536.400 146.400 ;
        RECT 535.700 142.400 536.300 145.600 ;
        RECT 537.200 143.600 538.000 144.400 ;
        RECT 535.600 141.600 536.400 142.400 ;
        RECT 529.200 133.600 530.000 134.400 ;
        RECT 529.200 131.600 530.000 132.400 ;
        RECT 529.300 130.400 529.900 131.600 ;
        RECT 529.200 129.600 530.000 130.400 ;
        RECT 532.400 126.200 533.200 137.800 ;
        RECT 535.600 130.200 536.400 135.800 ;
        RECT 537.300 134.400 537.900 143.600 ;
        RECT 543.700 134.400 544.300 173.600 ;
        RECT 545.300 172.400 545.900 175.600 ;
        RECT 551.600 173.600 552.400 174.400 ;
        RECT 545.200 171.600 546.000 172.400 ;
        RECT 545.200 169.600 546.000 170.400 ;
        RECT 548.400 169.600 549.200 170.400 ;
        RECT 545.300 156.400 545.900 169.600 ;
        RECT 545.200 155.600 546.000 156.400 ;
        RECT 545.200 153.600 546.000 154.400 ;
        RECT 545.300 148.400 545.900 153.600 ;
        RECT 545.200 147.600 546.000 148.400 ;
        RECT 546.800 144.200 547.600 155.800 ;
        RECT 548.500 138.400 549.100 169.600 ;
        RECT 551.600 159.600 552.400 160.400 ;
        RECT 550.000 149.600 550.800 150.400 ;
        RECT 548.400 137.600 549.200 138.400 ;
        RECT 545.200 135.600 546.000 136.400 ;
        RECT 551.700 134.400 552.300 159.600 ;
        RECT 553.300 148.400 553.900 179.700 ;
        RECT 554.800 177.600 555.600 178.400 ;
        RECT 558.000 173.600 558.800 174.400 ;
        RECT 558.100 172.400 558.700 173.600 ;
        RECT 566.100 172.400 566.700 189.600 ;
        RECT 570.800 184.200 571.600 197.800 ;
        RECT 572.400 184.200 573.200 197.800 ;
        RECT 574.000 184.200 574.800 195.800 ;
        RECT 575.700 192.400 576.300 211.600 ;
        RECT 577.200 209.600 578.000 210.400 ;
        RECT 577.300 198.400 577.900 209.600 ;
        RECT 577.200 197.600 578.000 198.400 ;
        RECT 575.600 191.600 576.400 192.400 ;
        RECT 575.600 187.600 576.400 188.400 ;
        RECT 577.200 184.200 578.000 195.800 ;
        RECT 578.800 185.600 579.600 186.400 ;
        RECT 572.400 181.600 573.200 182.400 ;
        RECT 567.600 175.600 568.400 176.400 ;
        RECT 558.000 171.600 558.800 172.400 ;
        RECT 559.600 171.600 560.400 172.400 ;
        RECT 564.400 171.600 565.200 172.400 ;
        RECT 566.000 171.600 566.800 172.400 ;
        RECT 556.400 169.600 557.200 170.400 ;
        RECT 553.200 147.600 554.000 148.400 ;
        RECT 556.400 144.200 557.200 155.800 ;
        RECT 558.100 136.400 558.700 171.600 ;
        RECT 559.700 168.400 560.300 171.600 ;
        RECT 564.500 170.400 565.100 171.600 ;
        RECT 562.800 169.600 563.600 170.400 ;
        RECT 564.400 169.600 565.200 170.400 ;
        RECT 567.700 168.400 568.300 175.600 ;
        RECT 559.600 167.600 560.400 168.400 ;
        RECT 562.800 167.600 563.600 168.400 ;
        RECT 567.600 167.600 568.400 168.400 ;
        RECT 559.600 146.200 560.400 151.800 ;
        RECT 562.900 148.400 563.500 167.600 ;
        RECT 567.700 154.400 568.300 167.600 ;
        RECT 567.600 153.600 568.400 154.400 ;
        RECT 562.800 147.600 563.600 148.400 ;
        RECT 569.200 147.600 570.000 148.400 ;
        RECT 561.200 146.300 562.000 146.400 ;
        RECT 561.200 145.700 563.500 146.300 ;
        RECT 561.200 145.600 562.000 145.700 ;
        RECT 559.600 139.600 560.400 140.400 ;
        RECT 559.700 138.400 560.300 139.600 ;
        RECT 559.600 137.600 560.400 138.400 ;
        RECT 562.900 136.400 563.500 145.700 ;
        RECT 569.300 144.400 569.900 147.600 ;
        RECT 569.200 143.600 570.000 144.400 ;
        RECT 556.400 135.600 557.200 136.400 ;
        RECT 558.000 135.600 558.800 136.400 ;
        RECT 561.200 135.600 562.000 136.400 ;
        RECT 562.800 135.600 563.600 136.400 ;
        RECT 537.200 133.600 538.000 134.400 ;
        RECT 538.800 133.600 539.600 134.400 ;
        RECT 543.600 133.600 544.400 134.400 ;
        RECT 551.600 133.600 552.400 134.400 ;
        RECT 538.900 132.400 539.500 133.600 ;
        RECT 551.700 132.400 552.300 133.600 ;
        RECT 538.800 131.600 539.600 132.400 ;
        RECT 540.400 131.600 541.200 132.400 ;
        RECT 546.800 131.600 547.600 132.400 ;
        RECT 551.600 131.600 552.400 132.400 ;
        RECT 553.200 131.600 554.000 132.400 ;
        RECT 546.900 128.400 547.500 131.600 ;
        RECT 553.300 130.400 553.900 131.600 ;
        RECT 561.300 130.400 561.900 135.600 ;
        RECT 562.900 134.400 563.500 135.600 ;
        RECT 562.800 133.600 563.600 134.400 ;
        RECT 564.400 131.600 565.200 132.400 ;
        RECT 567.600 131.600 568.400 132.400 ;
        RECT 569.200 131.600 570.000 132.400 ;
        RECT 570.800 131.600 571.600 132.400 ;
        RECT 553.200 129.600 554.000 130.400 ;
        RECT 556.400 129.600 557.200 130.400 ;
        RECT 561.200 129.600 562.000 130.400 ;
        RECT 567.600 129.600 568.400 130.400 ;
        RECT 546.800 127.600 547.600 128.400 ;
        RECT 550.000 123.600 550.800 124.400 ;
        RECT 534.000 113.600 534.800 114.400 ;
        RECT 537.200 113.600 538.000 114.400 ;
        RECT 530.800 111.600 531.600 112.400 ;
        RECT 534.100 110.400 534.700 113.600 ;
        RECT 537.300 112.400 537.900 113.600 ;
        RECT 537.200 111.600 538.000 112.400 ;
        RECT 526.000 109.600 526.800 110.400 ;
        RECT 529.200 109.600 530.000 110.400 ;
        RECT 534.000 109.600 534.800 110.400 ;
        RECT 529.300 108.400 529.900 109.600 ;
        RECT 524.400 107.600 525.200 108.400 ;
        RECT 529.200 107.600 530.000 108.400 ;
        RECT 524.500 96.400 525.100 107.600 ;
        RECT 534.100 96.400 534.700 109.600 ;
        RECT 535.600 107.600 536.400 108.400 ;
        RECT 538.800 107.600 539.600 108.400 ;
        RECT 524.400 95.600 525.200 96.400 ;
        RECT 527.600 95.600 528.400 96.400 ;
        RECT 534.000 95.600 534.800 96.400 ;
        RECT 537.200 95.600 538.000 96.400 ;
        RECT 527.700 94.400 528.300 95.600 ;
        RECT 527.600 93.600 528.400 94.400 ;
        RECT 532.400 93.600 533.200 94.400 ;
        RECT 522.800 91.600 523.600 92.400 ;
        RECT 524.400 91.600 525.200 92.400 ;
        RECT 524.500 88.400 525.100 91.600 ;
        RECT 524.400 87.600 525.200 88.400 ;
        RECT 522.800 81.600 523.600 82.400 ;
        RECT 522.900 52.400 523.500 81.600 ;
        RECT 526.000 71.600 526.800 72.400 ;
        RECT 526.100 70.400 526.700 71.600 ;
        RECT 526.000 69.600 526.800 70.400 ;
        RECT 526.000 67.600 526.800 68.400 ;
        RECT 521.200 51.600 522.000 52.400 ;
        RECT 522.800 51.600 523.600 52.400 ;
        RECT 519.600 31.600 520.400 32.400 ;
        RECT 519.700 30.400 520.300 31.600 ;
        RECT 521.300 30.400 521.900 51.600 ;
        RECT 524.400 49.600 525.200 50.400 ;
        RECT 526.100 44.400 526.700 67.600 ;
        RECT 527.700 60.400 528.300 93.600 ;
        RECT 532.500 92.400 533.100 93.600 ;
        RECT 537.300 92.400 537.900 95.600 ;
        RECT 538.900 94.400 539.500 107.600 ;
        RECT 542.000 104.200 542.800 115.800 ;
        RECT 550.100 114.400 550.700 123.600 ;
        RECT 550.000 113.600 550.800 114.400 ;
        RECT 548.400 109.600 549.200 110.400 ;
        RECT 551.600 104.200 552.400 115.800 ;
        RECT 553.200 107.600 554.000 108.400 ;
        RECT 553.300 106.400 553.900 107.600 ;
        RECT 553.200 105.600 554.000 106.400 ;
        RECT 554.800 106.200 555.600 111.800 ;
        RECT 556.500 110.400 557.100 129.600 ;
        RECT 569.300 124.400 569.900 131.600 ;
        RECT 570.900 130.400 571.500 131.600 ;
        RECT 570.800 129.600 571.600 130.400 ;
        RECT 569.200 123.600 570.000 124.400 ;
        RECT 567.600 115.600 568.400 116.400 ;
        RECT 567.700 112.400 568.300 115.600 ;
        RECT 567.600 111.600 568.400 112.400 ;
        RECT 569.200 111.600 570.000 112.400 ;
        RECT 569.300 110.400 569.900 111.600 ;
        RECT 556.400 109.600 557.200 110.400 ;
        RECT 564.400 109.600 565.200 110.400 ;
        RECT 569.200 109.600 570.000 110.400 ;
        RECT 570.800 109.600 571.600 110.400 ;
        RECT 556.500 102.400 557.100 109.600 ;
        RECT 562.800 107.600 563.600 108.400 ;
        RECT 556.400 101.600 557.200 102.400 ;
        RECT 542.000 99.600 542.800 100.400 ;
        RECT 542.100 98.400 542.700 99.600 ;
        RECT 562.900 98.400 563.500 107.600 ;
        RECT 566.000 103.600 566.800 104.400 ;
        RECT 566.100 98.400 566.700 103.600 ;
        RECT 542.000 97.600 542.800 98.400 ;
        RECT 548.400 97.600 549.200 98.400 ;
        RECT 538.800 93.600 539.600 94.400 ;
        RECT 540.400 93.600 541.200 94.400 ;
        RECT 532.400 91.600 533.200 92.400 ;
        RECT 537.200 91.600 538.000 92.400 ;
        RECT 534.000 89.600 534.800 90.400 ;
        RECT 545.200 89.600 546.000 90.400 ;
        RECT 545.300 88.400 545.900 89.600 ;
        RECT 543.600 87.600 544.400 88.400 ;
        RECT 545.200 87.600 546.000 88.400 ;
        RECT 543.700 76.400 544.300 87.600 ;
        RECT 529.200 64.200 530.000 75.800 ;
        RECT 543.600 75.600 544.400 76.400 ;
        RECT 546.800 75.600 547.600 76.400 ;
        RECT 535.600 73.600 536.400 74.400 ;
        RECT 543.600 73.600 544.400 74.400 ;
        RECT 543.700 72.400 544.300 73.600 ;
        RECT 532.400 66.200 533.200 71.800 ;
        RECT 543.600 71.600 544.400 72.400 ;
        RECT 535.600 69.600 536.400 70.400 ;
        RECT 534.000 67.600 534.800 68.400 ;
        RECT 540.400 67.600 541.200 68.400 ;
        RECT 543.600 67.600 544.400 68.400 ;
        RECT 530.800 61.600 531.600 62.400 ;
        RECT 527.600 59.600 528.400 60.400 ;
        RECT 527.600 55.600 528.400 56.400 ;
        RECT 527.700 52.400 528.300 55.600 ;
        RECT 530.900 54.400 531.500 61.600 ;
        RECT 530.800 53.600 531.600 54.400 ;
        RECT 532.400 53.600 533.200 54.400 ;
        RECT 532.500 52.400 533.100 53.600 ;
        RECT 527.600 51.600 528.400 52.400 ;
        RECT 529.200 51.600 530.000 52.400 ;
        RECT 532.400 51.600 533.200 52.400 ;
        RECT 526.000 43.600 526.800 44.400 ;
        RECT 524.400 39.600 525.200 40.400 ;
        RECT 519.600 29.600 520.400 30.400 ;
        RECT 521.200 29.600 522.000 30.400 ;
        RECT 521.200 27.600 522.000 28.400 ;
        RECT 522.800 27.600 523.600 28.400 ;
        RECT 521.300 24.400 521.900 27.600 ;
        RECT 524.500 26.400 525.100 39.600 ;
        RECT 526.100 28.400 526.700 43.600 ;
        RECT 532.500 32.400 533.100 51.600 ;
        RECT 534.100 48.400 534.700 67.600 ;
        RECT 542.000 59.600 542.800 60.400 ;
        RECT 538.800 57.600 539.600 58.400 ;
        RECT 535.600 55.600 536.400 56.400 ;
        RECT 535.700 50.400 536.300 55.600 ;
        RECT 535.600 49.600 536.400 50.400 ;
        RECT 534.000 47.600 534.800 48.400 ;
        RECT 537.200 47.600 538.000 48.400 ;
        RECT 535.600 45.600 536.400 46.400 ;
        RECT 535.700 36.400 536.300 45.600 ;
        RECT 537.300 38.400 537.900 47.600 ;
        RECT 538.900 38.400 539.500 57.600 ;
        RECT 542.100 54.400 542.700 59.600 ;
        RECT 543.700 58.400 544.300 67.600 ;
        RECT 545.200 65.600 546.000 66.400 ;
        RECT 543.600 57.600 544.400 58.400 ;
        RECT 543.700 56.400 544.300 57.600 ;
        RECT 543.600 55.600 544.400 56.400 ;
        RECT 542.000 53.600 542.800 54.400 ;
        RECT 540.400 51.600 541.200 52.400 ;
        RECT 540.500 50.400 541.100 51.600 ;
        RECT 540.400 49.600 541.200 50.400 ;
        RECT 540.400 47.600 541.200 48.400 ;
        RECT 537.200 37.600 538.000 38.400 ;
        RECT 538.800 37.600 539.600 38.400 ;
        RECT 535.600 35.600 536.400 36.400 ;
        RECT 532.400 32.300 533.200 32.400 ;
        RECT 532.400 31.700 534.700 32.300 ;
        RECT 532.400 31.600 533.200 31.700 ;
        RECT 526.000 27.600 526.800 28.400 ;
        RECT 524.400 25.600 525.200 26.400 ;
        RECT 521.200 23.600 522.000 24.400 ;
        RECT 524.500 14.400 525.100 25.600 ;
        RECT 521.200 13.600 522.000 14.400 ;
        RECT 524.400 13.600 525.200 14.400 ;
        RECT 529.200 13.600 530.000 14.400 ;
        RECT 530.800 13.600 531.600 14.400 ;
        RECT 521.300 12.400 521.900 13.600 ;
        RECT 529.300 12.400 529.900 13.600 ;
        RECT 514.800 11.600 515.600 12.400 ;
        RECT 518.000 11.600 518.800 12.400 ;
        RECT 521.200 11.600 522.000 12.400 ;
        RECT 522.800 11.600 523.600 12.400 ;
        RECT 526.000 11.600 526.800 12.400 ;
        RECT 529.200 11.600 530.000 12.400 ;
        RECT 526.100 10.400 526.700 11.600 ;
        RECT 530.900 10.400 531.500 13.600 ;
        RECT 534.100 12.400 534.700 31.700 ;
        RECT 535.700 28.400 536.300 35.600 ;
        RECT 538.900 32.400 539.500 37.600 ;
        RECT 543.600 33.600 544.400 34.400 ;
        RECT 546.900 32.400 547.500 75.600 ;
        RECT 548.500 70.400 549.100 97.600 ;
        RECT 550.000 86.200 550.800 97.800 ;
        RECT 556.400 91.600 557.200 92.400 ;
        RECT 559.600 86.200 560.400 97.800 ;
        RECT 562.800 97.600 563.600 98.400 ;
        RECT 566.000 97.600 566.800 98.400 ;
        RECT 569.200 97.600 570.000 98.400 ;
        RECT 561.200 95.600 562.000 96.400 ;
        RECT 561.300 94.400 561.900 95.600 ;
        RECT 561.200 93.600 562.000 94.400 ;
        RECT 562.800 90.200 563.600 95.800 ;
        RECT 569.300 94.400 569.900 97.600 ;
        RECT 564.400 93.600 565.200 94.400 ;
        RECT 569.200 93.600 570.000 94.400 ;
        RECT 570.900 92.400 571.500 109.600 ;
        RECT 572.500 104.400 573.100 181.600 ;
        RECT 578.900 180.400 579.500 185.600 ;
        RECT 580.400 184.200 581.200 195.800 ;
        RECT 582.000 184.200 582.800 197.800 ;
        RECT 583.600 184.200 584.400 197.800 ;
        RECT 585.200 184.200 586.000 197.800 ;
        RECT 578.800 179.600 579.600 180.400 ;
        RECT 582.000 179.600 582.800 180.400 ;
        RECT 574.000 171.600 574.800 172.400 ;
        RECT 575.600 164.200 576.400 177.800 ;
        RECT 577.200 164.200 578.000 177.800 ;
        RECT 578.800 164.200 579.600 177.800 ;
        RECT 580.400 166.200 581.200 177.800 ;
        RECT 582.100 176.400 582.700 179.600 ;
        RECT 582.000 175.600 582.800 176.400 ;
        RECT 582.100 160.400 582.700 175.600 ;
        RECT 583.600 166.200 584.400 177.800 ;
        RECT 585.200 173.600 586.000 174.400 ;
        RECT 586.800 166.200 587.600 177.800 ;
        RECT 588.400 164.200 589.200 177.800 ;
        RECT 590.000 164.200 590.800 177.800 ;
        RECT 591.700 176.400 592.300 213.600 ;
        RECT 594.800 193.600 595.600 194.400 ;
        RECT 594.900 190.400 595.500 193.600 ;
        RECT 594.800 189.600 595.800 190.400 ;
        RECT 591.600 175.600 592.400 176.400 ;
        RECT 594.800 171.600 595.600 172.400 ;
        RECT 582.000 159.600 582.800 160.400 ;
        RECT 585.200 159.600 586.000 160.400 ;
        RECT 575.600 155.600 576.400 156.400 ;
        RECT 575.700 132.400 576.300 155.600 ;
        RECT 578.800 144.200 579.600 157.800 ;
        RECT 580.400 144.200 581.200 157.800 ;
        RECT 582.000 144.200 582.800 157.800 ;
        RECT 583.600 144.200 584.400 155.800 ;
        RECT 585.300 146.400 585.900 159.600 ;
        RECT 585.200 145.600 586.000 146.400 ;
        RECT 585.300 142.400 585.900 145.600 ;
        RECT 586.800 144.200 587.600 155.800 ;
        RECT 588.400 147.600 589.200 148.400 ;
        RECT 590.000 144.200 590.800 155.800 ;
        RECT 591.600 144.200 592.400 157.800 ;
        RECT 593.200 144.200 594.000 157.800 ;
        RECT 594.900 150.400 595.500 171.600 ;
        RECT 594.800 149.600 595.600 150.400 ;
        RECT 578.800 141.600 579.600 142.400 ;
        RECT 585.200 141.600 586.000 142.400 ;
        RECT 586.800 141.600 587.600 142.400 ;
        RECT 591.600 141.600 592.400 142.400 ;
        RECT 578.900 134.400 579.500 141.600 ;
        RECT 585.200 137.600 586.000 138.400 ;
        RECT 578.800 133.600 579.600 134.400 ;
        RECT 575.600 131.600 576.400 132.400 ;
        RECT 583.600 131.600 584.400 132.400 ;
        RECT 585.200 131.600 586.000 132.400 ;
        RECT 583.700 130.400 584.300 131.600 ;
        RECT 583.600 129.600 584.400 130.400 ;
        RECT 585.200 127.600 586.000 128.400 ;
        RECT 585.300 118.400 585.900 127.600 ;
        RECT 578.800 109.600 579.600 110.400 ;
        RECT 572.400 103.600 573.200 104.400 ;
        RECT 578.900 92.400 579.500 109.600 ;
        RECT 580.400 104.200 581.200 117.800 ;
        RECT 582.000 104.200 582.800 117.800 ;
        RECT 583.600 104.200 584.400 117.800 ;
        RECT 585.200 117.600 586.000 118.400 ;
        RECT 585.200 104.200 586.000 115.800 ;
        RECT 586.900 106.400 587.500 141.600 ;
        RECT 588.400 133.600 589.200 134.400 ;
        RECT 590.000 130.200 590.800 135.800 ;
        RECT 591.700 134.400 592.300 141.600 ;
        RECT 591.600 133.600 592.400 134.400 ;
        RECT 593.200 126.200 594.000 137.800 ;
        RECT 594.800 131.600 595.600 132.600 ;
        RECT 596.500 120.400 597.100 233.600 ;
        RECT 604.400 231.600 605.200 232.400 ;
        RECT 604.400 229.600 605.200 230.400 ;
        RECT 602.800 227.600 603.600 228.400 ;
        RECT 604.400 225.600 605.200 226.400 ;
        RECT 604.500 218.400 605.100 225.600 ;
        RECT 604.400 217.600 605.200 218.400 ;
        RECT 598.000 191.600 598.800 192.400 ;
        RECT 601.200 189.600 602.000 190.400 ;
        RECT 602.800 189.600 603.600 190.400 ;
        RECT 601.300 186.300 601.900 189.600 ;
        RECT 602.800 187.600 603.600 188.400 ;
        RECT 601.300 185.700 603.500 186.300 ;
        RECT 598.000 183.600 598.800 184.400 ;
        RECT 601.200 183.600 602.000 184.400 ;
        RECT 598.100 160.400 598.700 183.600 ;
        RECT 599.600 173.600 600.400 174.400 ;
        RECT 599.600 169.600 600.400 170.400 ;
        RECT 599.600 167.600 600.400 168.400 ;
        RECT 598.000 159.600 598.800 160.400 ;
        RECT 598.000 149.600 598.800 150.400 ;
        RECT 596.400 119.600 597.200 120.400 ;
        RECT 586.800 105.600 587.600 106.400 ;
        RECT 588.400 104.200 589.200 115.800 ;
        RECT 590.000 107.600 590.800 108.400 ;
        RECT 591.600 104.200 592.400 115.800 ;
        RECT 593.200 104.200 594.000 117.800 ;
        RECT 594.800 104.200 595.600 117.800 ;
        RECT 598.100 110.400 598.700 149.600 ;
        RECT 599.700 110.400 600.300 167.600 ;
        RECT 598.000 109.600 598.800 110.400 ;
        RECT 599.600 109.600 600.400 110.400 ;
        RECT 601.300 108.300 601.900 183.600 ;
        RECT 602.900 172.400 603.500 185.700 ;
        RECT 602.800 171.600 603.600 172.400 ;
        RECT 602.900 168.400 603.500 171.600 ;
        RECT 602.800 167.600 603.600 168.400 ;
        RECT 606.100 150.400 606.700 281.600 ;
        RECT 607.600 231.600 608.400 232.400 ;
        RECT 607.700 184.400 608.300 231.600 ;
        RECT 607.600 183.600 608.400 184.400 ;
        RECT 606.000 149.600 606.800 150.400 ;
        RECT 602.800 143.600 603.600 144.400 ;
        RECT 602.900 140.400 603.500 143.600 ;
        RECT 602.800 139.600 603.600 140.400 ;
        RECT 609.200 139.600 610.000 140.400 ;
        RECT 602.800 126.200 603.600 137.800 ;
        RECT 607.600 137.600 608.400 138.400 ;
        RECT 607.700 130.400 608.300 137.600 ;
        RECT 607.600 129.600 608.400 130.400 ;
        RECT 604.400 111.600 605.200 112.400 ;
        RECT 606.000 109.600 606.800 110.400 ;
        RECT 607.600 109.600 608.400 110.400 ;
        RECT 599.700 107.700 601.900 108.300 ;
        RECT 570.800 91.600 571.600 92.400 ;
        RECT 578.800 91.600 579.600 92.400 ;
        RECT 567.600 89.600 568.400 90.400 ;
        RECT 574.000 89.600 574.800 90.400 ;
        RECT 561.200 85.600 562.000 86.400 ;
        RECT 558.000 73.600 558.800 74.400 ;
        RECT 561.300 72.400 561.900 85.600 ;
        RECT 562.800 81.600 563.600 82.400 ;
        RECT 561.200 71.600 562.000 72.400 ;
        RECT 548.400 69.600 549.200 70.400 ;
        RECT 554.800 69.600 555.600 70.400 ;
        RECT 561.200 69.600 562.000 70.400 ;
        RECT 548.400 67.600 549.200 68.400 ;
        RECT 553.200 63.600 554.000 64.400 ;
        RECT 548.400 46.200 549.200 57.800 ;
        RECT 550.000 51.600 550.800 52.400 ;
        RECT 551.600 51.600 552.400 52.400 ;
        RECT 550.100 44.400 550.700 51.600 ;
        RECT 551.700 48.400 552.300 51.600 ;
        RECT 551.600 47.600 552.400 48.400 ;
        RECT 550.000 43.600 550.800 44.400 ;
        RECT 553.300 40.400 553.900 63.600 ;
        RECT 554.900 54.400 555.500 69.600 ;
        RECT 556.400 67.600 557.200 68.400 ;
        RECT 556.500 62.400 557.100 67.600 ;
        RECT 559.600 63.600 560.400 64.400 ;
        RECT 556.400 61.600 557.200 62.400 ;
        RECT 554.800 53.600 555.600 54.400 ;
        RECT 558.000 46.200 558.800 57.800 ;
        RECT 559.700 54.400 560.300 63.600 ;
        RECT 559.600 53.600 560.400 54.400 ;
        RECT 561.200 50.200 562.000 55.800 ;
        RECT 553.200 39.600 554.000 40.400 ;
        RECT 551.600 35.600 552.400 36.400 ;
        RECT 551.700 32.400 552.300 35.600 ;
        RECT 553.200 33.600 554.000 34.400 ;
        RECT 553.300 32.400 553.900 33.600 ;
        RECT 562.900 32.400 563.500 81.600 ;
        RECT 564.400 71.600 565.200 72.400 ;
        RECT 564.500 70.400 565.100 71.600 ;
        RECT 564.400 69.600 565.200 70.400 ;
        RECT 567.700 58.400 568.300 89.600 ;
        RECT 569.200 87.600 570.000 88.400 ;
        RECT 569.300 70.400 569.900 87.600 ;
        RECT 570.800 83.600 571.600 84.400 ;
        RECT 583.600 84.200 584.400 97.800 ;
        RECT 585.200 84.200 586.000 97.800 ;
        RECT 586.800 86.200 587.600 97.800 ;
        RECT 588.400 97.600 589.200 98.400 ;
        RECT 588.500 94.400 589.100 97.600 ;
        RECT 588.400 93.600 589.200 94.400 ;
        RECT 588.400 91.600 589.200 92.400 ;
        RECT 570.900 76.400 571.500 83.600 ;
        RECT 570.800 75.600 571.600 76.400 ;
        RECT 572.400 73.600 573.200 74.400 ;
        RECT 575.600 73.600 576.400 74.400 ;
        RECT 572.500 72.400 573.100 73.600 ;
        RECT 572.400 71.600 573.200 72.400 ;
        RECT 569.200 69.600 570.000 70.400 ;
        RECT 570.800 69.600 571.600 70.400 ;
        RECT 575.600 69.600 576.400 70.400 ;
        RECT 570.900 68.400 571.500 69.600 ;
        RECT 570.800 67.600 571.600 68.400 ;
        RECT 577.200 67.600 578.000 68.400 ;
        RECT 577.300 60.400 577.900 67.600 ;
        RECT 578.800 66.200 579.600 71.800 ;
        RECT 580.400 67.600 581.200 68.400 ;
        RECT 580.500 64.400 581.100 67.600 ;
        RECT 580.400 63.600 581.200 64.400 ;
        RECT 582.000 64.200 582.800 75.800 ;
        RECT 583.600 73.600 584.400 74.400 ;
        RECT 583.700 70.200 584.300 73.600 ;
        RECT 583.600 69.400 584.400 70.200 ;
        RECT 577.200 59.600 578.000 60.400 ;
        RECT 588.500 60.300 589.100 91.600 ;
        RECT 590.000 86.200 590.800 97.800 ;
        RECT 591.600 95.600 592.400 96.400 ;
        RECT 591.700 78.400 592.300 95.600 ;
        RECT 593.200 86.200 594.000 97.800 ;
        RECT 594.800 84.200 595.600 97.800 ;
        RECT 596.400 84.200 597.200 97.800 ;
        RECT 598.000 84.200 598.800 97.800 ;
        RECT 599.700 78.400 600.300 107.700 ;
        RECT 604.400 107.600 605.200 108.400 ;
        RECT 601.200 91.600 602.000 92.400 ;
        RECT 591.600 77.600 592.400 78.400 ;
        RECT 594.800 77.600 595.600 78.400 ;
        RECT 599.600 77.600 600.400 78.400 ;
        RECT 591.600 64.200 592.400 75.800 ;
        RECT 586.900 59.700 589.100 60.300 ;
        RECT 567.600 57.600 568.400 58.400 ;
        RECT 578.800 57.600 579.600 58.400 ;
        RECT 575.600 53.600 576.400 54.400 ;
        RECT 575.700 46.400 576.300 53.600 ;
        RECT 586.900 52.400 587.500 59.700 ;
        RECT 586.800 51.600 587.600 52.400 ;
        RECT 586.800 49.600 587.600 50.400 ;
        RECT 575.600 45.600 576.400 46.400 ;
        RECT 564.400 43.600 565.200 44.400 ;
        RECT 538.800 31.600 539.600 32.400 ;
        RECT 546.800 31.600 547.600 32.400 ;
        RECT 551.600 31.600 552.400 32.400 ;
        RECT 553.200 31.600 554.000 32.400 ;
        RECT 556.400 31.600 557.200 32.400 ;
        RECT 559.600 31.600 560.400 32.400 ;
        RECT 562.800 31.600 563.600 32.400 ;
        RECT 556.500 30.400 557.100 31.600 ;
        RECT 542.000 29.600 542.800 30.400 ;
        RECT 548.400 29.600 549.200 30.400 ;
        RECT 556.400 29.600 557.200 30.400 ;
        RECT 535.600 27.600 536.400 28.400 ;
        RECT 538.800 27.600 539.600 28.400 ;
        RECT 538.900 26.400 539.500 27.600 ;
        RECT 538.800 25.600 539.600 26.400 ;
        RECT 538.800 23.600 539.600 24.400 ;
        RECT 538.900 18.400 539.500 23.600 ;
        RECT 538.800 17.600 539.600 18.400 ;
        RECT 542.100 12.400 542.700 29.600 ;
        RECT 559.700 28.400 560.300 31.600 ;
        RECT 562.900 30.400 563.500 31.600 ;
        RECT 562.800 29.600 563.600 30.400 ;
        RECT 543.600 27.600 544.400 28.400 ;
        RECT 545.200 27.600 546.000 28.400 ;
        RECT 551.600 27.600 552.400 28.400 ;
        RECT 558.000 27.600 558.800 28.400 ;
        RECT 559.600 27.600 560.400 28.400 ;
        RECT 561.200 27.600 562.000 28.400 ;
        RECT 543.700 18.400 544.300 27.600 ;
        RECT 545.300 24.400 545.900 27.600 ;
        RECT 558.100 26.400 558.700 27.600 ;
        RECT 558.000 25.600 558.800 26.400 ;
        RECT 562.800 25.600 563.600 26.400 ;
        RECT 545.200 23.600 546.000 24.400 ;
        RECT 553.200 23.600 554.000 24.400 ;
        RECT 543.600 17.600 544.400 18.400 ;
        RECT 543.700 14.400 544.300 17.600 ;
        RECT 543.600 13.600 544.400 14.400 ;
        RECT 534.000 11.600 534.800 12.400 ;
        RECT 542.000 11.600 542.800 12.400 ;
        RECT 513.200 9.600 514.000 10.400 ;
        RECT 518.000 9.600 518.800 10.400 ;
        RECT 526.000 9.600 526.800 10.400 ;
        RECT 530.800 9.600 531.600 10.400 ;
        RECT 513.300 8.400 513.900 9.600 ;
        RECT 513.200 7.600 514.000 8.400 ;
        RECT 548.400 6.200 549.200 17.800 ;
        RECT 553.300 16.400 553.900 23.600 ;
        RECT 562.900 18.400 563.500 25.600 ;
        RECT 564.500 18.400 565.100 43.600 ;
        RECT 574.000 37.600 574.800 38.400 ;
        RECT 570.800 35.600 571.600 36.400 ;
        RECT 570.800 33.600 571.600 34.400 ;
        RECT 570.900 18.400 571.500 33.600 ;
        RECT 574.100 18.400 574.700 37.600 ;
        RECT 580.400 24.200 581.200 37.800 ;
        RECT 582.000 24.200 582.800 37.800 ;
        RECT 583.600 24.200 584.400 37.800 ;
        RECT 585.200 24.200 586.000 35.800 ;
        RECT 586.900 26.400 587.500 49.600 ;
        RECT 588.400 44.200 589.200 57.800 ;
        RECT 590.000 44.200 590.800 57.800 ;
        RECT 591.600 44.200 592.400 57.800 ;
        RECT 593.200 46.200 594.000 57.800 ;
        RECT 594.900 56.400 595.500 77.600 ;
        RECT 596.400 73.600 597.200 74.400 ;
        RECT 596.500 72.400 597.100 73.600 ;
        RECT 601.300 72.400 601.900 91.600 ;
        RECT 606.100 82.400 606.700 109.600 ;
        RECT 609.300 108.400 609.900 139.600 ;
        RECT 609.200 107.600 610.000 108.400 ;
        RECT 607.600 97.600 608.400 98.400 ;
        RECT 606.000 81.600 606.800 82.400 ;
        RECT 602.800 75.600 603.600 76.400 ;
        RECT 602.900 72.400 603.500 75.600 ;
        RECT 596.400 71.600 597.200 72.400 ;
        RECT 601.200 71.600 602.000 72.400 ;
        RECT 602.800 71.600 603.600 72.400 ;
        RECT 601.300 68.400 601.900 71.600 ;
        RECT 606.100 70.400 606.700 81.600 ;
        RECT 606.000 69.600 606.800 70.400 ;
        RECT 598.000 67.600 598.800 68.400 ;
        RECT 601.200 67.600 602.000 68.400 ;
        RECT 606.000 67.600 606.800 68.400 ;
        RECT 607.600 67.600 608.400 68.400 ;
        RECT 602.800 63.600 603.600 64.400 ;
        RECT 602.900 60.400 603.500 63.600 ;
        RECT 598.000 59.600 598.800 60.400 ;
        RECT 602.800 59.600 603.600 60.400 ;
        RECT 594.800 55.600 595.600 56.400 ;
        RECT 594.900 50.400 595.500 55.600 ;
        RECT 594.800 49.600 595.600 50.400 ;
        RECT 596.400 46.200 597.200 57.800 ;
        RECT 598.100 54.400 598.700 59.600 ;
        RECT 598.000 53.600 598.800 54.400 ;
        RECT 598.000 51.600 598.800 52.400 ;
        RECT 586.800 25.600 587.600 26.400 ;
        RECT 588.400 24.200 589.200 35.800 ;
        RECT 590.000 27.600 590.800 28.400 ;
        RECT 590.000 25.600 590.800 26.400 ;
        RECT 590.100 18.400 590.700 25.600 ;
        RECT 591.600 24.200 592.400 35.800 ;
        RECT 593.200 24.200 594.000 37.800 ;
        RECT 594.800 24.200 595.600 37.800 ;
        RECT 598.100 30.400 598.700 51.600 ;
        RECT 599.600 46.200 600.400 57.800 ;
        RECT 601.200 44.200 602.000 57.800 ;
        RECT 602.800 44.200 603.600 57.800 ;
        RECT 604.400 41.600 605.200 42.400 ;
        RECT 604.500 38.400 605.100 41.600 ;
        RECT 604.400 37.600 605.200 38.400 ;
        RECT 606.100 30.400 606.700 67.600 ;
        RECT 598.000 29.600 598.800 30.400 ;
        RECT 601.200 29.600 602.000 30.400 ;
        RECT 606.000 29.600 606.800 30.400 ;
        RECT 553.200 15.600 554.000 16.400 ;
        RECT 554.800 11.600 555.600 12.400 ;
        RECT 558.000 6.200 558.800 17.800 ;
        RECT 559.600 17.600 560.400 18.400 ;
        RECT 562.800 17.600 563.600 18.400 ;
        RECT 564.400 17.600 565.200 18.400 ;
        RECT 570.800 17.600 571.600 18.400 ;
        RECT 574.000 17.600 574.800 18.400 ;
        RECT 559.700 14.400 560.300 17.600 ;
        RECT 559.600 13.600 560.400 14.400 ;
        RECT 561.200 10.200 562.000 15.800 ;
        RECT 566.000 13.600 566.800 14.400 ;
        RECT 567.600 11.600 568.400 12.400 ;
        RECT 570.800 9.600 571.600 10.400 ;
        RECT 583.600 4.200 584.400 17.800 ;
        RECT 585.200 4.200 586.000 17.800 ;
        RECT 586.800 4.200 587.600 17.800 ;
        RECT 588.400 6.200 589.200 17.800 ;
        RECT 590.000 17.600 590.800 18.400 ;
        RECT 590.100 16.400 590.700 17.600 ;
        RECT 590.000 15.600 590.800 16.400 ;
        RECT 591.600 6.200 592.400 17.800 ;
        RECT 593.200 15.600 594.000 16.400 ;
        RECT 593.300 14.400 593.900 15.600 ;
        RECT 593.200 13.600 594.000 14.400 ;
        RECT 594.800 6.200 595.600 17.800 ;
        RECT 596.400 4.200 597.200 17.800 ;
        RECT 598.000 4.200 598.800 17.800 ;
        RECT 601.300 12.400 601.900 29.600 ;
        RECT 607.700 18.400 608.300 67.600 ;
        RECT 607.600 17.600 608.400 18.400 ;
        RECT 601.200 11.600 602.000 12.400 ;
      LAYER via2 ;
        RECT 124.400 549.600 125.200 550.400 ;
        RECT 175.600 547.600 176.400 548.400 ;
        RECT 316.400 509.600 317.200 510.400 ;
        RECT 338.800 509.600 339.600 510.400 ;
        RECT 431.600 549.600 432.400 550.400 ;
        RECT 76.400 229.600 77.200 230.400 ;
        RECT 76.400 149.600 77.200 150.400 ;
        RECT 474.800 549.600 475.600 550.400 ;
        RECT 233.200 309.600 234.000 310.400 ;
        RECT 207.600 267.600 208.400 268.400 ;
        RECT 318.000 349.600 318.800 350.400 ;
        RECT 298.800 307.600 299.600 308.400 ;
        RECT 263.600 227.600 264.400 228.400 ;
        RECT 162.800 69.600 163.600 70.400 ;
        RECT 153.200 29.600 154.000 30.400 ;
        RECT 250.800 111.600 251.600 112.400 ;
        RECT 495.600 413.600 496.400 414.400 ;
        RECT 550.000 389.600 550.800 390.400 ;
        RECT 460.400 347.600 461.200 348.400 ;
        RECT 316.400 93.600 317.200 94.400 ;
        RECT 303.600 27.600 304.400 28.400 ;
        RECT 598.000 349.600 598.800 350.400 ;
        RECT 418.800 109.600 419.600 110.400 ;
        RECT 479.600 189.600 480.400 190.400 ;
        RECT 594.800 189.600 595.600 190.400 ;
      LAYER metal3 ;
        RECT 591.600 556.300 592.400 556.400 ;
        RECT 607.600 556.300 608.400 556.400 ;
        RECT 591.600 555.700 608.400 556.300 ;
        RECT 591.600 555.600 592.400 555.700 ;
        RECT 607.600 555.600 608.400 555.700 ;
        RECT 47.600 554.300 48.400 554.400 ;
        RECT 63.600 554.300 64.400 554.400 ;
        RECT 47.600 553.700 64.400 554.300 ;
        RECT 47.600 553.600 48.400 553.700 ;
        RECT 63.600 553.600 64.400 553.700 ;
        RECT 156.400 554.300 157.200 554.400 ;
        RECT 190.000 554.300 190.800 554.400 ;
        RECT 156.400 553.700 190.800 554.300 ;
        RECT 156.400 553.600 157.200 553.700 ;
        RECT 190.000 553.600 190.800 553.700 ;
        RECT 406.000 554.300 406.800 554.400 ;
        RECT 425.200 554.300 426.000 554.400 ;
        RECT 406.000 553.700 426.000 554.300 ;
        RECT 406.000 553.600 406.800 553.700 ;
        RECT 425.200 553.600 426.000 553.700 ;
        RECT 57.200 552.300 58.000 552.400 ;
        RECT 60.400 552.300 61.200 552.400 ;
        RECT 57.200 551.700 61.200 552.300 ;
        RECT 57.200 551.600 58.000 551.700 ;
        RECT 60.400 551.600 61.200 551.700 ;
        RECT 186.800 552.300 187.600 552.400 ;
        RECT 193.200 552.300 194.000 552.400 ;
        RECT 186.800 551.700 194.000 552.300 ;
        RECT 186.800 551.600 187.600 551.700 ;
        RECT 193.200 551.600 194.000 551.700 ;
        RECT 361.200 552.300 362.000 552.400 ;
        RECT 364.400 552.300 365.200 552.400 ;
        RECT 361.200 551.700 365.200 552.300 ;
        RECT 361.200 551.600 362.000 551.700 ;
        RECT 364.400 551.600 365.200 551.700 ;
        RECT 420.400 552.300 421.200 552.400 ;
        RECT 444.400 552.300 445.200 552.400 ;
        RECT 420.400 551.700 445.200 552.300 ;
        RECT 420.400 551.600 421.200 551.700 ;
        RECT 444.400 551.600 445.200 551.700 ;
        RECT 463.600 552.300 464.400 552.400 ;
        RECT 487.600 552.300 488.400 552.400 ;
        RECT 494.000 552.300 494.800 552.400 ;
        RECT 463.600 551.700 494.800 552.300 ;
        RECT 463.600 551.600 464.400 551.700 ;
        RECT 487.600 551.600 488.400 551.700 ;
        RECT 494.000 551.600 494.800 551.700 ;
        RECT 518.000 552.300 518.800 552.400 ;
        RECT 521.200 552.300 522.000 552.400 ;
        RECT 518.000 551.700 522.000 552.300 ;
        RECT 518.000 551.600 518.800 551.700 ;
        RECT 521.200 551.600 522.000 551.700 ;
        RECT 532.400 552.300 533.200 552.400 ;
        RECT 550.000 552.300 550.800 552.400 ;
        RECT 532.400 551.700 550.800 552.300 ;
        RECT 532.400 551.600 533.200 551.700 ;
        RECT 550.000 551.600 550.800 551.700 ;
        RECT 33.200 550.300 34.000 550.400 ;
        RECT 44.400 550.300 45.200 550.400 ;
        RECT 60.400 550.300 61.200 550.400 ;
        RECT 33.200 549.700 61.200 550.300 ;
        RECT 33.200 549.600 34.000 549.700 ;
        RECT 44.400 549.600 45.200 549.700 ;
        RECT 60.400 549.600 61.200 549.700 ;
        RECT 122.800 550.300 123.600 550.400 ;
        RECT 124.400 550.300 125.200 550.400 ;
        RECT 122.800 549.700 125.200 550.300 ;
        RECT 122.800 549.600 123.600 549.700 ;
        RECT 124.400 549.600 125.200 549.700 ;
        RECT 167.600 550.300 168.400 550.400 ;
        RECT 177.200 550.300 178.000 550.400 ;
        RECT 167.600 549.700 178.000 550.300 ;
        RECT 167.600 549.600 168.400 549.700 ;
        RECT 177.200 549.600 178.000 549.700 ;
        RECT 186.800 550.300 187.600 550.400 ;
        RECT 190.000 550.300 190.800 550.400 ;
        RECT 186.800 549.700 190.800 550.300 ;
        RECT 186.800 549.600 187.600 549.700 ;
        RECT 190.000 549.600 190.800 549.700 ;
        RECT 215.600 550.300 216.400 550.400 ;
        RECT 244.400 550.300 245.200 550.400 ;
        RECT 215.600 549.700 245.200 550.300 ;
        RECT 215.600 549.600 216.400 549.700 ;
        RECT 244.400 549.600 245.200 549.700 ;
        RECT 332.400 550.300 333.200 550.400 ;
        RECT 345.200 550.300 346.000 550.400 ;
        RECT 332.400 549.700 346.000 550.300 ;
        RECT 332.400 549.600 333.200 549.700 ;
        RECT 345.200 549.600 346.000 549.700 ;
        RECT 362.800 550.300 363.600 550.400 ;
        RECT 390.000 550.300 390.800 550.400 ;
        RECT 362.800 549.700 390.800 550.300 ;
        RECT 362.800 549.600 363.600 549.700 ;
        RECT 390.000 549.600 390.800 549.700 ;
        RECT 399.600 550.300 400.400 550.400 ;
        RECT 412.400 550.300 413.200 550.400 ;
        RECT 399.600 549.700 413.200 550.300 ;
        RECT 399.600 549.600 400.400 549.700 ;
        RECT 412.400 549.600 413.200 549.700 ;
        RECT 431.600 550.300 432.400 550.400 ;
        RECT 441.200 550.300 442.000 550.400 ;
        RECT 431.600 549.700 442.000 550.300 ;
        RECT 431.600 549.600 432.400 549.700 ;
        RECT 441.200 549.600 442.000 549.700 ;
        RECT 474.800 550.300 475.600 550.400 ;
        RECT 478.000 550.300 478.800 550.400 ;
        RECT 474.800 549.700 478.800 550.300 ;
        RECT 474.800 549.600 475.600 549.700 ;
        RECT 478.000 549.600 478.800 549.700 ;
        RECT 486.000 550.300 486.800 550.400 ;
        RECT 505.200 550.300 506.000 550.400 ;
        RECT 486.000 549.700 506.000 550.300 ;
        RECT 486.000 549.600 486.800 549.700 ;
        RECT 505.200 549.600 506.000 549.700 ;
        RECT 527.600 550.300 528.400 550.400 ;
        RECT 532.400 550.300 533.200 550.400 ;
        RECT 527.600 549.700 533.200 550.300 ;
        RECT 527.600 549.600 528.400 549.700 ;
        RECT 532.400 549.600 533.200 549.700 ;
        RECT 2.800 548.300 3.600 548.400 ;
        RECT 17.200 548.300 18.000 548.400 ;
        RECT 2.800 547.700 18.000 548.300 ;
        RECT 2.800 547.600 3.600 547.700 ;
        RECT 17.200 547.600 18.000 547.700 ;
        RECT 57.200 548.300 58.000 548.400 ;
        RECT 86.000 548.300 86.800 548.400 ;
        RECT 57.200 547.700 86.800 548.300 ;
        RECT 57.200 547.600 58.000 547.700 ;
        RECT 86.000 547.600 86.800 547.700 ;
        RECT 111.600 548.300 112.400 548.400 ;
        RECT 121.200 548.300 122.000 548.400 ;
        RECT 111.600 547.700 122.000 548.300 ;
        RECT 111.600 547.600 112.400 547.700 ;
        RECT 121.200 547.600 122.000 547.700 ;
        RECT 175.600 548.300 176.400 548.400 ;
        RECT 183.600 548.300 184.400 548.400 ;
        RECT 175.600 547.700 184.400 548.300 ;
        RECT 175.600 547.600 176.400 547.700 ;
        RECT 183.600 547.600 184.400 547.700 ;
        RECT 226.800 548.300 227.600 548.400 ;
        RECT 262.000 548.300 262.800 548.400 ;
        RECT 226.800 547.700 262.800 548.300 ;
        RECT 226.800 547.600 227.600 547.700 ;
        RECT 262.000 547.600 262.800 547.700 ;
        RECT 322.800 548.300 323.600 548.400 ;
        RECT 343.600 548.300 344.400 548.400 ;
        RECT 322.800 547.700 344.400 548.300 ;
        RECT 322.800 547.600 323.600 547.700 ;
        RECT 343.600 547.600 344.400 547.700 ;
        RECT 350.000 548.300 350.800 548.400 ;
        RECT 364.400 548.300 365.200 548.400 ;
        RECT 457.200 548.300 458.000 548.400 ;
        RECT 350.000 547.700 458.000 548.300 ;
        RECT 350.000 547.600 350.800 547.700 ;
        RECT 364.400 547.600 365.200 547.700 ;
        RECT 457.200 547.600 458.000 547.700 ;
        RECT 518.000 548.300 518.800 548.400 ;
        RECT 529.200 548.300 530.000 548.400 ;
        RECT 518.000 547.700 530.000 548.300 ;
        RECT 518.000 547.600 518.800 547.700 ;
        RECT 529.200 547.600 530.000 547.700 ;
        RECT 578.800 548.300 579.600 548.400 ;
        RECT 593.200 548.300 594.000 548.400 ;
        RECT 578.800 547.700 594.000 548.300 ;
        RECT 578.800 547.600 579.600 547.700 ;
        RECT 593.200 547.600 594.000 547.700 ;
        RECT 17.200 546.300 18.000 546.400 ;
        RECT 20.400 546.300 21.200 546.400 ;
        RECT 17.200 545.700 21.200 546.300 ;
        RECT 17.200 545.600 18.000 545.700 ;
        RECT 20.400 545.600 21.200 545.700 ;
        RECT 28.400 546.300 29.200 546.400 ;
        RECT 33.200 546.300 34.000 546.400 ;
        RECT 74.800 546.300 75.600 546.400 ;
        RECT 28.400 545.700 75.600 546.300 ;
        RECT 28.400 545.600 29.200 545.700 ;
        RECT 33.200 545.600 34.000 545.700 ;
        RECT 74.800 545.600 75.600 545.700 ;
        RECT 95.600 546.300 96.400 546.400 ;
        RECT 145.200 546.300 146.000 546.400 ;
        RECT 95.600 545.700 146.000 546.300 ;
        RECT 95.600 545.600 96.400 545.700 ;
        RECT 145.200 545.600 146.000 545.700 ;
        RECT 238.000 546.300 238.800 546.400 ;
        RECT 255.600 546.300 256.400 546.400 ;
        RECT 238.000 545.700 256.400 546.300 ;
        RECT 238.000 545.600 238.800 545.700 ;
        RECT 255.600 545.600 256.400 545.700 ;
        RECT 351.600 546.300 352.400 546.400 ;
        RECT 362.800 546.300 363.600 546.400 ;
        RECT 366.000 546.300 366.800 546.400 ;
        RECT 351.600 545.700 366.800 546.300 ;
        RECT 351.600 545.600 352.400 545.700 ;
        RECT 362.800 545.600 363.600 545.700 ;
        RECT 366.000 545.600 366.800 545.700 ;
        RECT 417.200 546.300 418.000 546.400 ;
        RECT 430.000 546.300 430.800 546.400 ;
        RECT 417.200 545.700 430.800 546.300 ;
        RECT 417.200 545.600 418.000 545.700 ;
        RECT 430.000 545.600 430.800 545.700 ;
        RECT 449.200 546.300 450.000 546.400 ;
        RECT 455.600 546.300 456.400 546.400 ;
        RECT 449.200 545.700 456.400 546.300 ;
        RECT 449.200 545.600 450.000 545.700 ;
        RECT 455.600 545.600 456.400 545.700 ;
        RECT 522.800 546.300 523.600 546.400 ;
        RECT 538.800 546.300 539.600 546.400 ;
        RECT 522.800 545.700 539.600 546.300 ;
        RECT 522.800 545.600 523.600 545.700 ;
        RECT 538.800 545.600 539.600 545.700 ;
        RECT 554.800 546.300 555.600 546.400 ;
        RECT 561.200 546.300 562.000 546.400 ;
        RECT 575.600 546.300 576.400 546.400 ;
        RECT 586.800 546.300 587.600 546.400 ;
        RECT 554.800 545.700 587.600 546.300 ;
        RECT 554.800 545.600 555.600 545.700 ;
        RECT 561.200 545.600 562.000 545.700 ;
        RECT 575.600 545.600 576.400 545.700 ;
        RECT 586.800 545.600 587.600 545.700 ;
        RECT 110.000 544.300 110.800 544.400 ;
        RECT 118.000 544.300 118.800 544.400 ;
        RECT 110.000 543.700 118.800 544.300 ;
        RECT 110.000 543.600 110.800 543.700 ;
        RECT 118.000 543.600 118.800 543.700 ;
        RECT 250.800 543.600 251.600 544.400 ;
        RECT 434.800 544.300 435.600 544.400 ;
        RECT 468.400 544.300 469.200 544.400 ;
        RECT 434.800 543.700 469.200 544.300 ;
        RECT 434.800 543.600 435.600 543.700 ;
        RECT 468.400 543.600 469.200 543.700 ;
        RECT 486.000 544.300 486.800 544.400 ;
        RECT 492.400 544.300 493.200 544.400 ;
        RECT 513.200 544.300 514.000 544.400 ;
        RECT 527.600 544.300 528.400 544.400 ;
        RECT 486.000 543.700 528.400 544.300 ;
        RECT 486.000 543.600 486.800 543.700 ;
        RECT 492.400 543.600 493.200 543.700 ;
        RECT 513.200 543.600 514.000 543.700 ;
        RECT 527.600 543.600 528.400 543.700 ;
        RECT 558.000 544.300 558.800 544.400 ;
        RECT 559.600 544.300 560.400 544.400 ;
        RECT 558.000 543.700 560.400 544.300 ;
        RECT 558.000 543.600 558.800 543.700 ;
        RECT 559.600 543.600 560.400 543.700 ;
        RECT 118.000 542.300 118.800 542.400 ;
        RECT 122.800 542.300 123.600 542.400 ;
        RECT 118.000 541.700 123.600 542.300 ;
        RECT 118.000 541.600 118.800 541.700 ;
        RECT 122.800 541.600 123.600 541.700 ;
        RECT 193.200 542.300 194.000 542.400 ;
        RECT 220.400 542.300 221.200 542.400 ;
        RECT 241.200 542.300 242.000 542.400 ;
        RECT 247.600 542.300 248.400 542.400 ;
        RECT 292.400 542.300 293.200 542.400 ;
        RECT 298.800 542.300 299.600 542.400 ;
        RECT 193.200 541.700 299.600 542.300 ;
        RECT 468.500 542.300 469.100 543.600 ;
        RECT 502.000 542.300 502.800 542.400 ;
        RECT 468.500 541.700 502.800 542.300 ;
        RECT 193.200 541.600 194.000 541.700 ;
        RECT 220.400 541.600 221.200 541.700 ;
        RECT 241.200 541.600 242.000 541.700 ;
        RECT 247.600 541.600 248.400 541.700 ;
        RECT 292.400 541.600 293.200 541.700 ;
        RECT 298.800 541.600 299.600 541.700 ;
        RECT 502.000 541.600 502.800 541.700 ;
        RECT 510.000 542.300 510.800 542.400 ;
        RECT 532.400 542.300 533.200 542.400 ;
        RECT 545.200 542.300 546.000 542.400 ;
        RECT 510.000 541.700 546.000 542.300 ;
        RECT 510.000 541.600 510.800 541.700 ;
        RECT 532.400 541.600 533.200 541.700 ;
        RECT 545.200 541.600 546.000 541.700 ;
        RECT 116.400 540.300 117.200 540.400 ;
        RECT 137.200 540.300 138.000 540.400 ;
        RECT 116.400 539.700 138.000 540.300 ;
        RECT 116.400 539.600 117.200 539.700 ;
        RECT 137.200 539.600 138.000 539.700 ;
        RECT 196.400 540.300 197.200 540.400 ;
        RECT 226.800 540.300 227.600 540.400 ;
        RECT 196.400 539.700 227.600 540.300 ;
        RECT 196.400 539.600 197.200 539.700 ;
        RECT 226.800 539.600 227.600 539.700 ;
        RECT 270.000 539.600 270.800 540.400 ;
        RECT 342.000 540.300 342.800 540.400 ;
        RECT 353.200 540.300 354.000 540.400 ;
        RECT 358.000 540.300 358.800 540.400 ;
        RECT 377.200 540.300 378.000 540.400 ;
        RECT 450.800 540.300 451.600 540.400 ;
        RECT 538.800 540.300 539.600 540.400 ;
        RECT 594.800 540.300 595.600 540.400 ;
        RECT 602.800 540.300 603.600 540.400 ;
        RECT 342.000 539.700 603.600 540.300 ;
        RECT 342.000 539.600 342.800 539.700 ;
        RECT 353.200 539.600 354.000 539.700 ;
        RECT 358.000 539.600 358.800 539.700 ;
        RECT 377.200 539.600 378.000 539.700 ;
        RECT 450.800 539.600 451.600 539.700 ;
        RECT 538.800 539.600 539.600 539.700 ;
        RECT 594.800 539.600 595.600 539.700 ;
        RECT 602.800 539.600 603.600 539.700 ;
        RECT 201.200 538.300 202.000 538.400 ;
        RECT 207.600 538.300 208.400 538.400 ;
        RECT 201.200 537.700 208.400 538.300 ;
        RECT 270.100 538.300 270.700 539.600 ;
        RECT 302.000 538.300 302.800 538.400 ;
        RECT 270.100 537.700 302.800 538.300 ;
        RECT 201.200 537.600 202.000 537.700 ;
        RECT 207.600 537.600 208.400 537.700 ;
        RECT 302.000 537.600 302.800 537.700 ;
        RECT 370.800 538.300 371.600 538.400 ;
        RECT 372.400 538.300 373.200 538.400 ;
        RECT 370.800 537.700 373.200 538.300 ;
        RECT 370.800 537.600 371.600 537.700 ;
        RECT 372.400 537.600 373.200 537.700 ;
        RECT 438.000 538.300 438.800 538.400 ;
        RECT 450.800 538.300 451.600 538.400 ;
        RECT 474.800 538.300 475.600 538.400 ;
        RECT 481.200 538.300 482.000 538.400 ;
        RECT 487.600 538.300 488.400 538.400 ;
        RECT 534.000 538.300 534.800 538.400 ;
        RECT 438.000 537.700 534.800 538.300 ;
        RECT 438.000 537.600 438.800 537.700 ;
        RECT 450.800 537.600 451.600 537.700 ;
        RECT 474.800 537.600 475.600 537.700 ;
        RECT 481.200 537.600 482.000 537.700 ;
        RECT 487.600 537.600 488.400 537.700 ;
        RECT 534.000 537.600 534.800 537.700 ;
        RECT 34.800 536.300 35.600 536.400 ;
        RECT 42.800 536.300 43.600 536.400 ;
        RECT 34.800 535.700 43.600 536.300 ;
        RECT 34.800 535.600 35.600 535.700 ;
        RECT 42.800 535.600 43.600 535.700 ;
        RECT 46.000 535.600 46.800 536.400 ;
        RECT 103.600 536.300 104.400 536.400 ;
        RECT 108.400 536.300 109.200 536.400 ;
        RECT 103.600 535.700 109.200 536.300 ;
        RECT 103.600 535.600 104.400 535.700 ;
        RECT 108.400 535.600 109.200 535.700 ;
        RECT 188.400 536.300 189.200 536.400 ;
        RECT 217.200 536.300 218.000 536.400 ;
        RECT 188.400 535.700 218.000 536.300 ;
        RECT 188.400 535.600 189.200 535.700 ;
        RECT 217.200 535.600 218.000 535.700 ;
        RECT 218.800 536.300 219.600 536.400 ;
        RECT 242.800 536.300 243.600 536.400 ;
        RECT 244.400 536.300 245.200 536.400 ;
        RECT 218.800 535.700 245.200 536.300 ;
        RECT 218.800 535.600 219.600 535.700 ;
        RECT 242.800 535.600 243.600 535.700 ;
        RECT 244.400 535.600 245.200 535.700 ;
        RECT 265.200 536.300 266.000 536.400 ;
        RECT 273.200 536.300 274.000 536.400 ;
        RECT 276.400 536.300 277.200 536.400 ;
        RECT 265.200 535.700 277.200 536.300 ;
        RECT 265.200 535.600 266.000 535.700 ;
        RECT 273.200 535.600 274.000 535.700 ;
        RECT 276.400 535.600 277.200 535.700 ;
        RECT 289.200 536.300 290.000 536.400 ;
        RECT 295.600 536.300 296.400 536.400 ;
        RECT 289.200 535.700 296.400 536.300 ;
        RECT 289.200 535.600 290.000 535.700 ;
        RECT 295.600 535.600 296.400 535.700 ;
        RECT 298.800 536.300 299.600 536.400 ;
        RECT 310.000 536.300 310.800 536.400 ;
        RECT 298.800 535.700 310.800 536.300 ;
        RECT 298.800 535.600 299.600 535.700 ;
        RECT 310.000 535.600 310.800 535.700 ;
        RECT 319.600 536.300 320.400 536.400 ;
        RECT 332.400 536.300 333.200 536.400 ;
        RECT 319.600 535.700 333.200 536.300 ;
        RECT 319.600 535.600 320.400 535.700 ;
        RECT 332.400 535.600 333.200 535.700 ;
        RECT 335.600 536.300 336.400 536.400 ;
        RECT 350.000 536.300 350.800 536.400 ;
        RECT 335.600 535.700 350.800 536.300 ;
        RECT 335.600 535.600 336.400 535.700 ;
        RECT 350.000 535.600 350.800 535.700 ;
        RECT 367.600 536.300 368.400 536.400 ;
        RECT 386.800 536.300 387.600 536.400 ;
        RECT 399.600 536.300 400.400 536.400 ;
        RECT 417.200 536.300 418.000 536.400 ;
        RECT 367.600 535.700 418.000 536.300 ;
        RECT 367.600 535.600 368.400 535.700 ;
        RECT 386.800 535.600 387.600 535.700 ;
        RECT 399.600 535.600 400.400 535.700 ;
        RECT 417.200 535.600 418.000 535.700 ;
        RECT 455.600 536.300 456.400 536.400 ;
        RECT 466.800 536.300 467.600 536.400 ;
        RECT 492.400 536.300 493.200 536.400 ;
        RECT 498.800 536.300 499.600 536.400 ;
        RECT 455.600 535.700 499.600 536.300 ;
        RECT 455.600 535.600 456.400 535.700 ;
        RECT 466.800 535.600 467.600 535.700 ;
        RECT 492.400 535.600 493.200 535.700 ;
        RECT 498.800 535.600 499.600 535.700 ;
        RECT 526.000 535.600 526.800 536.400 ;
        RECT 543.600 536.300 544.400 536.400 ;
        RECT 564.400 536.300 565.200 536.400 ;
        RECT 543.600 535.700 565.200 536.300 ;
        RECT 543.600 535.600 544.400 535.700 ;
        RECT 564.400 535.600 565.200 535.700 ;
        RECT 14.000 534.300 14.800 534.400 ;
        RECT 36.400 534.300 37.200 534.400 ;
        RECT 14.000 533.700 37.200 534.300 ;
        RECT 14.000 533.600 14.800 533.700 ;
        RECT 36.400 533.600 37.200 533.700 ;
        RECT 41.200 534.300 42.000 534.400 ;
        RECT 46.000 534.300 46.800 534.400 ;
        RECT 41.200 533.700 46.800 534.300 ;
        RECT 41.200 533.600 42.000 533.700 ;
        RECT 46.000 533.600 46.800 533.700 ;
        RECT 55.600 534.300 56.400 534.400 ;
        RECT 84.400 534.300 85.200 534.400 ;
        RECT 55.600 533.700 85.200 534.300 ;
        RECT 55.600 533.600 56.400 533.700 ;
        RECT 84.400 533.600 85.200 533.700 ;
        RECT 97.200 534.300 98.000 534.400 ;
        RECT 105.200 534.300 106.000 534.400 ;
        RECT 111.600 534.300 112.400 534.400 ;
        RECT 97.200 533.700 112.400 534.300 ;
        RECT 97.200 533.600 98.000 533.700 ;
        RECT 105.200 533.600 106.000 533.700 ;
        RECT 111.600 533.600 112.400 533.700 ;
        RECT 146.800 534.300 147.600 534.400 ;
        RECT 158.000 534.300 158.800 534.400 ;
        RECT 191.600 534.300 192.400 534.400 ;
        RECT 146.800 533.700 192.400 534.300 ;
        RECT 146.800 533.600 147.600 533.700 ;
        RECT 158.000 533.600 158.800 533.700 ;
        RECT 191.600 533.600 192.400 533.700 ;
        RECT 214.000 534.300 214.800 534.400 ;
        RECT 220.400 534.300 221.200 534.400 ;
        RECT 214.000 533.700 221.200 534.300 ;
        RECT 214.000 533.600 214.800 533.700 ;
        RECT 220.400 533.600 221.200 533.700 ;
        RECT 242.800 534.300 243.600 534.400 ;
        RECT 246.000 534.300 246.800 534.400 ;
        RECT 242.800 533.700 246.800 534.300 ;
        RECT 242.800 533.600 243.600 533.700 ;
        RECT 246.000 533.600 246.800 533.700 ;
        RECT 350.000 534.300 350.800 534.400 ;
        RECT 358.000 534.300 358.800 534.400 ;
        RECT 350.000 533.700 358.800 534.300 ;
        RECT 350.000 533.600 350.800 533.700 ;
        RECT 358.000 533.600 358.800 533.700 ;
        RECT 382.000 534.300 382.800 534.400 ;
        RECT 402.800 534.300 403.600 534.400 ;
        RECT 382.000 533.700 403.600 534.300 ;
        RECT 382.000 533.600 382.800 533.700 ;
        RECT 402.800 533.600 403.600 533.700 ;
        RECT 418.800 534.300 419.600 534.400 ;
        RECT 434.800 534.300 435.600 534.400 ;
        RECT 438.000 534.300 438.800 534.400 ;
        RECT 418.800 533.700 438.800 534.300 ;
        RECT 418.800 533.600 419.600 533.700 ;
        RECT 434.800 533.600 435.600 533.700 ;
        RECT 438.000 533.600 438.800 533.700 ;
        RECT 447.600 534.300 448.400 534.400 ;
        RECT 465.200 534.300 466.000 534.400 ;
        RECT 471.600 534.300 472.400 534.400 ;
        RECT 484.400 534.300 485.200 534.400 ;
        RECT 490.800 534.300 491.600 534.400 ;
        RECT 497.200 534.300 498.000 534.400 ;
        RECT 514.800 534.300 515.600 534.400 ;
        RECT 447.600 533.700 515.600 534.300 ;
        RECT 447.600 533.600 448.400 533.700 ;
        RECT 465.200 533.600 466.000 533.700 ;
        RECT 471.600 533.600 472.400 533.700 ;
        RECT 484.400 533.600 485.200 533.700 ;
        RECT 490.800 533.600 491.600 533.700 ;
        RECT 497.200 533.600 498.000 533.700 ;
        RECT 514.800 533.600 515.600 533.700 ;
        RECT 561.200 534.300 562.000 534.400 ;
        RECT 578.800 534.300 579.600 534.400 ;
        RECT 561.200 533.700 579.600 534.300 ;
        RECT 561.200 533.600 562.000 533.700 ;
        RECT 578.800 533.600 579.600 533.700 ;
        RECT 598.000 534.300 598.800 534.400 ;
        RECT 612.400 534.300 613.200 534.400 ;
        RECT 598.000 533.700 613.200 534.300 ;
        RECT 598.000 533.600 598.800 533.700 ;
        RECT 612.400 533.600 613.200 533.700 ;
        RECT 39.600 532.300 40.400 532.400 ;
        RECT 44.400 532.300 45.200 532.400 ;
        RECT 52.400 532.300 53.200 532.400 ;
        RECT 39.600 531.700 53.200 532.300 ;
        RECT 39.600 531.600 40.400 531.700 ;
        RECT 44.400 531.600 45.200 531.700 ;
        RECT 52.400 531.600 53.200 531.700 ;
        RECT 105.200 532.300 106.000 532.400 ;
        RECT 113.200 532.300 114.000 532.400 ;
        RECT 105.200 531.700 114.000 532.300 ;
        RECT 105.200 531.600 106.000 531.700 ;
        RECT 113.200 531.600 114.000 531.700 ;
        RECT 140.400 532.300 141.200 532.400 ;
        RECT 161.200 532.300 162.000 532.400 ;
        RECT 140.400 531.700 162.000 532.300 ;
        RECT 140.400 531.600 141.200 531.700 ;
        RECT 161.200 531.600 162.000 531.700 ;
        RECT 199.600 532.300 200.400 532.400 ;
        RECT 204.400 532.300 205.200 532.400 ;
        RECT 199.600 531.700 205.200 532.300 ;
        RECT 199.600 531.600 200.400 531.700 ;
        RECT 204.400 531.600 205.200 531.700 ;
        RECT 345.200 532.300 346.000 532.400 ;
        RECT 391.600 532.300 392.400 532.400 ;
        RECT 345.200 531.700 392.400 532.300 ;
        RECT 345.200 531.600 346.000 531.700 ;
        RECT 391.600 531.600 392.400 531.700 ;
        RECT 433.200 532.300 434.000 532.400 ;
        RECT 452.400 532.300 453.200 532.400 ;
        RECT 433.200 531.700 453.200 532.300 ;
        RECT 433.200 531.600 434.000 531.700 ;
        RECT 452.400 531.600 453.200 531.700 ;
        RECT 454.000 532.300 454.800 532.400 ;
        RECT 458.800 532.300 459.600 532.400 ;
        RECT 474.800 532.300 475.600 532.400 ;
        RECT 482.800 532.300 483.600 532.400 ;
        RECT 454.000 531.700 473.900 532.300 ;
        RECT 454.000 531.600 454.800 531.700 ;
        RECT 458.800 531.600 459.600 531.700 ;
        RECT 33.200 530.300 34.000 530.400 ;
        RECT 36.400 530.300 37.200 530.400 ;
        RECT 42.800 530.300 43.600 530.400 ;
        RECT 33.200 529.700 43.600 530.300 ;
        RECT 33.200 529.600 34.000 529.700 ;
        RECT 36.400 529.600 37.200 529.700 ;
        RECT 42.800 529.600 43.600 529.700 ;
        RECT 55.600 530.300 56.400 530.400 ;
        RECT 58.800 530.300 59.600 530.400 ;
        RECT 55.600 529.700 59.600 530.300 ;
        RECT 55.600 529.600 56.400 529.700 ;
        RECT 58.800 529.600 59.600 529.700 ;
        RECT 98.800 530.300 99.600 530.400 ;
        RECT 124.400 530.300 125.200 530.400 ;
        RECT 172.400 530.300 173.200 530.400 ;
        RECT 98.800 529.700 173.200 530.300 ;
        RECT 98.800 529.600 99.600 529.700 ;
        RECT 124.400 529.600 125.200 529.700 ;
        RECT 172.400 529.600 173.200 529.700 ;
        RECT 318.000 530.300 318.800 530.400 ;
        RECT 359.600 530.300 360.400 530.400 ;
        RECT 318.000 529.700 360.400 530.300 ;
        RECT 318.000 529.600 318.800 529.700 ;
        RECT 359.600 529.600 360.400 529.700 ;
        RECT 372.400 530.300 373.200 530.400 ;
        RECT 380.400 530.300 381.200 530.400 ;
        RECT 372.400 529.700 381.200 530.300 ;
        RECT 372.400 529.600 373.200 529.700 ;
        RECT 380.400 529.600 381.200 529.700 ;
        RECT 438.000 530.300 438.800 530.400 ;
        RECT 462.000 530.300 462.800 530.400 ;
        RECT 438.000 529.700 462.800 530.300 ;
        RECT 473.300 530.300 473.900 531.700 ;
        RECT 474.800 531.700 483.600 532.300 ;
        RECT 474.800 531.600 475.600 531.700 ;
        RECT 482.800 531.600 483.600 531.700 ;
        RECT 492.400 532.300 493.200 532.400 ;
        RECT 505.200 532.300 506.000 532.400 ;
        RECT 492.400 531.700 506.000 532.300 ;
        RECT 492.400 531.600 493.200 531.700 ;
        RECT 505.200 531.600 506.000 531.700 ;
        RECT 519.600 531.600 520.400 532.400 ;
        RECT 481.200 530.300 482.000 530.400 ;
        RECT 473.300 529.700 482.000 530.300 ;
        RECT 438.000 529.600 438.800 529.700 ;
        RECT 462.000 529.600 462.800 529.700 ;
        RECT 481.200 529.600 482.000 529.700 ;
        RECT 498.800 530.300 499.600 530.400 ;
        RECT 530.800 530.300 531.600 530.400 ;
        RECT 498.800 529.700 531.600 530.300 ;
        RECT 498.800 529.600 499.600 529.700 ;
        RECT 530.800 529.600 531.600 529.700 ;
        RECT 590.000 530.300 590.800 530.400 ;
        RECT 599.600 530.300 600.400 530.400 ;
        RECT 590.000 529.700 600.400 530.300 ;
        RECT 590.000 529.600 590.800 529.700 ;
        RECT 599.600 529.600 600.400 529.700 ;
        RECT 2.800 528.300 3.600 528.400 ;
        RECT 52.400 528.300 53.200 528.400 ;
        RECT 2.800 527.700 53.200 528.300 ;
        RECT 2.800 527.600 3.600 527.700 ;
        RECT 52.400 527.600 53.200 527.700 ;
        RECT 100.400 528.300 101.200 528.400 ;
        RECT 132.400 528.300 133.200 528.400 ;
        RECT 100.400 527.700 133.200 528.300 ;
        RECT 100.400 527.600 101.200 527.700 ;
        RECT 132.400 527.600 133.200 527.700 ;
        RECT 356.400 528.300 357.200 528.400 ;
        RECT 370.800 528.300 371.600 528.400 ;
        RECT 383.600 528.300 384.400 528.400 ;
        RECT 356.400 527.700 384.400 528.300 ;
        RECT 356.400 527.600 357.200 527.700 ;
        RECT 370.800 527.600 371.600 527.700 ;
        RECT 383.600 527.600 384.400 527.700 ;
        RECT 417.200 528.300 418.000 528.400 ;
        RECT 439.600 528.300 440.400 528.400 ;
        RECT 417.200 527.700 440.400 528.300 ;
        RECT 417.200 527.600 418.000 527.700 ;
        RECT 439.600 527.600 440.400 527.700 ;
        RECT 444.400 528.300 445.200 528.400 ;
        RECT 452.400 528.300 453.200 528.400 ;
        RECT 444.400 527.700 453.200 528.300 ;
        RECT 444.400 527.600 445.200 527.700 ;
        RECT 452.400 527.600 453.200 527.700 ;
        RECT 457.200 528.300 458.000 528.400 ;
        RECT 487.600 528.300 488.400 528.400 ;
        RECT 457.200 527.700 488.400 528.300 ;
        RECT 457.200 527.600 458.000 527.700 ;
        RECT 487.600 527.600 488.400 527.700 ;
        RECT 490.800 528.300 491.600 528.400 ;
        RECT 494.000 528.300 494.800 528.400 ;
        RECT 518.000 528.300 518.800 528.400 ;
        RECT 490.800 527.700 518.800 528.300 ;
        RECT 490.800 527.600 491.600 527.700 ;
        RECT 494.000 527.600 494.800 527.700 ;
        RECT 518.000 527.600 518.800 527.700 ;
        RECT 452.400 526.300 453.200 526.400 ;
        RECT 473.200 526.300 474.000 526.400 ;
        RECT 452.400 525.700 474.000 526.300 ;
        RECT 452.400 525.600 453.200 525.700 ;
        RECT 473.200 525.600 474.000 525.700 ;
        RECT 583.600 526.300 584.400 526.400 ;
        RECT 599.600 526.300 600.400 526.400 ;
        RECT 583.600 525.700 600.400 526.300 ;
        RECT 583.600 525.600 584.400 525.700 ;
        RECT 599.600 525.600 600.400 525.700 ;
        RECT 65.200 523.600 66.000 524.400 ;
        RECT 159.600 524.300 160.400 524.400 ;
        RECT 167.600 524.300 168.400 524.400 ;
        RECT 159.600 523.700 168.400 524.300 ;
        RECT 159.600 523.600 160.400 523.700 ;
        RECT 167.600 523.600 168.400 523.700 ;
        RECT 226.800 524.300 227.600 524.400 ;
        RECT 233.200 524.300 234.000 524.400 ;
        RECT 226.800 523.700 234.000 524.300 ;
        RECT 226.800 523.600 227.600 523.700 ;
        RECT 233.200 523.600 234.000 523.700 ;
        RECT 412.400 524.300 413.200 524.400 ;
        RECT 572.400 524.300 573.200 524.400 ;
        RECT 583.600 524.300 584.400 524.400 ;
        RECT 588.400 524.300 589.200 524.400 ;
        RECT 412.400 523.700 589.200 524.300 ;
        RECT 412.400 523.600 413.200 523.700 ;
        RECT 572.400 523.600 573.200 523.700 ;
        RECT 583.600 523.600 584.400 523.700 ;
        RECT 588.400 523.600 589.200 523.700 ;
        RECT 31.600 522.300 32.400 522.400 ;
        RECT 41.200 522.300 42.000 522.400 ;
        RECT 57.200 522.300 58.000 522.400 ;
        RECT 31.600 521.700 58.000 522.300 ;
        RECT 31.600 521.600 32.400 521.700 ;
        RECT 41.200 521.600 42.000 521.700 ;
        RECT 57.200 521.600 58.000 521.700 ;
        RECT 89.200 522.300 90.000 522.400 ;
        RECT 105.200 522.300 106.000 522.400 ;
        RECT 89.200 521.700 106.000 522.300 ;
        RECT 89.200 521.600 90.000 521.700 ;
        RECT 105.200 521.600 106.000 521.700 ;
        RECT 273.200 522.300 274.000 522.400 ;
        RECT 281.200 522.300 282.000 522.400 ;
        RECT 273.200 521.700 282.000 522.300 ;
        RECT 273.200 521.600 274.000 521.700 ;
        RECT 281.200 521.600 282.000 521.700 ;
        RECT 300.400 522.300 301.200 522.400 ;
        RECT 329.200 522.300 330.000 522.400 ;
        RECT 346.800 522.300 347.600 522.400 ;
        RECT 300.400 521.700 347.600 522.300 ;
        RECT 300.400 521.600 301.200 521.700 ;
        RECT 329.200 521.600 330.000 521.700 ;
        RECT 346.800 521.600 347.600 521.700 ;
        RECT 366.000 522.300 366.800 522.400 ;
        RECT 369.200 522.300 370.000 522.400 ;
        RECT 406.000 522.300 406.800 522.400 ;
        RECT 366.000 521.700 406.800 522.300 ;
        RECT 366.000 521.600 366.800 521.700 ;
        RECT 369.200 521.600 370.000 521.700 ;
        RECT 406.000 521.600 406.800 521.700 ;
        RECT 430.000 522.300 430.800 522.400 ;
        RECT 442.800 522.300 443.600 522.400 ;
        RECT 430.000 521.700 443.600 522.300 ;
        RECT 430.000 521.600 430.800 521.700 ;
        RECT 442.800 521.600 443.600 521.700 ;
        RECT 465.200 522.300 466.000 522.400 ;
        RECT 519.600 522.300 520.400 522.400 ;
        RECT 465.200 521.700 520.400 522.300 ;
        RECT 465.200 521.600 466.000 521.700 ;
        RECT 519.600 521.600 520.400 521.700 ;
        RECT 431.600 520.300 432.400 520.400 ;
        RECT 438.000 520.300 438.800 520.400 ;
        RECT 431.600 519.700 438.800 520.300 ;
        RECT 431.600 519.600 432.400 519.700 ;
        RECT 438.000 519.600 438.800 519.700 ;
        RECT 516.400 520.300 517.200 520.400 ;
        RECT 521.200 520.300 522.000 520.400 ;
        RECT 516.400 519.700 522.000 520.300 ;
        RECT 516.400 519.600 517.200 519.700 ;
        RECT 521.200 519.600 522.000 519.700 ;
        RECT 594.800 520.300 595.600 520.400 ;
        RECT 598.000 520.300 598.800 520.400 ;
        RECT 594.800 519.700 598.800 520.300 ;
        RECT 594.800 519.600 595.600 519.700 ;
        RECT 598.000 519.600 598.800 519.700 ;
        RECT 410.800 518.300 411.600 518.400 ;
        RECT 498.800 518.300 499.600 518.400 ;
        RECT 410.800 517.700 499.600 518.300 ;
        RECT 410.800 517.600 411.600 517.700 ;
        RECT 498.800 517.600 499.600 517.700 ;
        RECT 503.600 518.300 504.400 518.400 ;
        RECT 542.000 518.300 542.800 518.400 ;
        RECT 575.600 518.300 576.400 518.400 ;
        RECT 503.600 517.700 576.400 518.300 ;
        RECT 503.600 517.600 504.400 517.700 ;
        RECT 542.000 517.600 542.800 517.700 ;
        RECT 575.600 517.600 576.400 517.700 ;
        RECT 482.800 516.300 483.600 516.400 ;
        RECT 542.000 516.300 542.800 516.400 ;
        RECT 545.200 516.300 546.000 516.400 ;
        RECT 482.800 515.700 546.000 516.300 ;
        RECT 482.800 515.600 483.600 515.700 ;
        RECT 542.000 515.600 542.800 515.700 ;
        RECT 545.200 515.600 546.000 515.700 ;
        RECT 46.000 514.300 46.800 514.400 ;
        RECT 44.500 513.700 46.800 514.300 ;
        RECT 26.800 510.300 27.600 510.400 ;
        RECT 42.800 510.300 43.600 510.400 ;
        RECT 26.800 509.700 43.600 510.300 ;
        RECT 44.500 510.300 45.100 513.700 ;
        RECT 46.000 513.600 46.800 513.700 ;
        RECT 81.200 514.300 82.000 514.400 ;
        RECT 86.000 514.300 86.800 514.400 ;
        RECT 102.000 514.300 102.800 514.400 ;
        RECT 105.200 514.300 106.000 514.400 ;
        RECT 153.200 514.300 154.000 514.400 ;
        RECT 81.200 513.700 154.000 514.300 ;
        RECT 81.200 513.600 82.000 513.700 ;
        RECT 86.000 513.600 86.800 513.700 ;
        RECT 102.000 513.600 102.800 513.700 ;
        RECT 105.200 513.600 106.000 513.700 ;
        RECT 153.200 513.600 154.000 513.700 ;
        RECT 372.400 514.300 373.200 514.400 ;
        RECT 393.200 514.300 394.000 514.400 ;
        RECT 372.400 513.700 394.000 514.300 ;
        RECT 372.400 513.600 373.200 513.700 ;
        RECT 393.200 513.600 394.000 513.700 ;
        RECT 398.000 514.300 398.800 514.400 ;
        RECT 409.200 514.300 410.000 514.400 ;
        RECT 484.400 514.300 485.200 514.400 ;
        RECT 505.200 514.300 506.000 514.400 ;
        RECT 522.800 514.300 523.600 514.400 ;
        RECT 398.000 513.700 523.600 514.300 ;
        RECT 398.000 513.600 398.800 513.700 ;
        RECT 409.200 513.600 410.000 513.700 ;
        RECT 484.400 513.600 485.200 513.700 ;
        RECT 505.200 513.600 506.000 513.700 ;
        RECT 522.800 513.600 523.600 513.700 ;
        RECT 535.600 514.300 536.400 514.400 ;
        RECT 545.200 514.300 546.000 514.400 ;
        RECT 535.600 513.700 546.000 514.300 ;
        RECT 535.600 513.600 536.400 513.700 ;
        RECT 545.200 513.600 546.000 513.700 ;
        RECT 46.000 512.300 46.800 512.400 ;
        RECT 54.000 512.300 54.800 512.400 ;
        RECT 46.000 511.700 54.800 512.300 ;
        RECT 46.000 511.600 46.800 511.700 ;
        RECT 54.000 511.600 54.800 511.700 ;
        RECT 71.600 512.300 72.400 512.400 ;
        RECT 79.600 512.300 80.400 512.400 ;
        RECT 71.600 511.700 80.400 512.300 ;
        RECT 71.600 511.600 72.400 511.700 ;
        RECT 79.600 511.600 80.400 511.700 ;
        RECT 110.000 512.300 110.800 512.400 ;
        RECT 114.800 512.300 115.600 512.400 ;
        RECT 130.800 512.300 131.600 512.400 ;
        RECT 110.000 511.700 131.600 512.300 ;
        RECT 110.000 511.600 110.800 511.700 ;
        RECT 114.800 511.600 115.600 511.700 ;
        RECT 130.800 511.600 131.600 511.700 ;
        RECT 319.600 512.300 320.400 512.400 ;
        RECT 335.600 512.300 336.400 512.400 ;
        RECT 319.600 511.700 336.400 512.300 ;
        RECT 319.600 511.600 320.400 511.700 ;
        RECT 335.600 511.600 336.400 511.700 ;
        RECT 375.600 512.300 376.400 512.400 ;
        RECT 378.800 512.300 379.600 512.400 ;
        RECT 398.000 512.300 398.800 512.400 ;
        RECT 410.800 512.300 411.600 512.400 ;
        RECT 375.600 511.700 411.600 512.300 ;
        RECT 375.600 511.600 376.400 511.700 ;
        RECT 378.800 511.600 379.600 511.700 ;
        RECT 398.000 511.600 398.800 511.700 ;
        RECT 410.800 511.600 411.600 511.700 ;
        RECT 436.400 512.300 437.200 512.400 ;
        RECT 439.600 512.300 440.400 512.400 ;
        RECT 465.200 512.300 466.000 512.400 ;
        RECT 436.400 511.700 466.000 512.300 ;
        RECT 436.400 511.600 437.200 511.700 ;
        RECT 439.600 511.600 440.400 511.700 ;
        RECT 465.200 511.600 466.000 511.700 ;
        RECT 468.400 512.300 469.200 512.400 ;
        RECT 490.800 512.300 491.600 512.400 ;
        RECT 468.400 511.700 491.600 512.300 ;
        RECT 468.400 511.600 469.200 511.700 ;
        RECT 490.800 511.600 491.600 511.700 ;
        RECT 511.600 512.300 512.400 512.400 ;
        RECT 518.000 512.300 518.800 512.400 ;
        RECT 511.600 511.700 518.800 512.300 ;
        RECT 511.600 511.600 512.400 511.700 ;
        RECT 518.000 511.600 518.800 511.700 ;
        RECT 522.800 512.300 523.600 512.400 ;
        RECT 548.400 512.300 549.200 512.400 ;
        RECT 522.800 511.700 549.200 512.300 ;
        RECT 522.800 511.600 523.600 511.700 ;
        RECT 548.400 511.600 549.200 511.700 ;
        RECT 569.200 512.300 570.000 512.400 ;
        RECT 578.800 512.300 579.600 512.400 ;
        RECT 569.200 511.700 579.600 512.300 ;
        RECT 569.200 511.600 570.000 511.700 ;
        RECT 578.800 511.600 579.600 511.700 ;
        RECT 46.000 510.300 46.800 510.400 ;
        RECT 44.500 509.700 46.800 510.300 ;
        RECT 26.800 509.600 27.600 509.700 ;
        RECT 42.800 509.600 43.600 509.700 ;
        RECT 46.000 509.600 46.800 509.700 ;
        RECT 52.400 510.300 53.200 510.400 ;
        RECT 121.200 510.300 122.000 510.400 ;
        RECT 52.400 509.700 122.000 510.300 ;
        RECT 52.400 509.600 53.200 509.700 ;
        RECT 121.200 509.600 122.000 509.700 ;
        RECT 170.800 510.300 171.600 510.400 ;
        RECT 183.600 510.300 184.400 510.400 ;
        RECT 170.800 509.700 184.400 510.300 ;
        RECT 170.800 509.600 171.600 509.700 ;
        RECT 183.600 509.600 184.400 509.700 ;
        RECT 236.400 510.300 237.200 510.400 ;
        RECT 241.200 510.300 242.000 510.400 ;
        RECT 236.400 509.700 242.000 510.300 ;
        RECT 236.400 509.600 237.200 509.700 ;
        RECT 241.200 509.600 242.000 509.700 ;
        RECT 279.600 510.300 280.400 510.400 ;
        RECT 313.200 510.300 314.000 510.400 ;
        RECT 316.400 510.300 317.200 510.400 ;
        RECT 279.600 509.700 317.200 510.300 ;
        RECT 279.600 509.600 280.400 509.700 ;
        RECT 313.200 509.600 314.000 509.700 ;
        RECT 316.400 509.600 317.200 509.700 ;
        RECT 329.200 510.300 330.000 510.400 ;
        RECT 338.800 510.300 339.600 510.400 ;
        RECT 329.200 509.700 339.600 510.300 ;
        RECT 329.200 509.600 330.000 509.700 ;
        RECT 338.800 509.600 339.600 509.700 ;
        RECT 364.400 510.300 365.200 510.400 ;
        RECT 390.000 510.300 390.800 510.400 ;
        RECT 364.400 509.700 390.800 510.300 ;
        RECT 364.400 509.600 365.200 509.700 ;
        RECT 390.000 509.600 390.800 509.700 ;
        RECT 391.600 510.300 392.400 510.400 ;
        RECT 396.400 510.300 397.200 510.400 ;
        RECT 391.600 509.700 397.200 510.300 ;
        RECT 391.600 509.600 392.400 509.700 ;
        RECT 396.400 509.600 397.200 509.700 ;
        RECT 414.000 510.300 414.800 510.400 ;
        RECT 415.600 510.300 416.400 510.400 ;
        RECT 414.000 509.700 416.400 510.300 ;
        RECT 414.000 509.600 414.800 509.700 ;
        RECT 415.600 509.600 416.400 509.700 ;
        RECT 434.800 510.300 435.600 510.400 ;
        RECT 441.200 510.300 442.000 510.400 ;
        RECT 466.800 510.300 467.600 510.400 ;
        RECT 434.800 509.700 467.600 510.300 ;
        RECT 434.800 509.600 435.600 509.700 ;
        RECT 441.200 509.600 442.000 509.700 ;
        RECT 466.800 509.600 467.600 509.700 ;
        RECT 476.400 510.300 477.200 510.400 ;
        RECT 486.000 510.300 486.800 510.400 ;
        RECT 476.400 509.700 486.800 510.300 ;
        RECT 476.400 509.600 477.200 509.700 ;
        RECT 486.000 509.600 486.800 509.700 ;
        RECT 487.600 510.300 488.400 510.400 ;
        RECT 538.800 510.300 539.600 510.400 ;
        RECT 569.300 510.300 569.900 511.600 ;
        RECT 487.600 509.700 569.900 510.300 ;
        RECT 487.600 509.600 488.400 509.700 ;
        RECT 538.800 509.600 539.600 509.700 ;
        RECT 12.400 508.300 13.200 508.400 ;
        RECT 17.200 508.300 18.000 508.400 ;
        RECT 22.000 508.300 22.800 508.400 ;
        RECT 12.400 507.700 22.800 508.300 ;
        RECT 12.400 507.600 13.200 507.700 ;
        RECT 17.200 507.600 18.000 507.700 ;
        RECT 22.000 507.600 22.800 507.700 ;
        RECT 38.000 508.300 38.800 508.400 ;
        RECT 47.600 508.300 48.400 508.400 ;
        RECT 55.600 508.300 56.400 508.400 ;
        RECT 79.600 508.300 80.400 508.400 ;
        RECT 38.000 507.700 80.400 508.300 ;
        RECT 38.000 507.600 38.800 507.700 ;
        RECT 47.600 507.600 48.400 507.700 ;
        RECT 55.600 507.600 56.400 507.700 ;
        RECT 79.600 507.600 80.400 507.700 ;
        RECT 116.400 508.300 117.200 508.400 ;
        RECT 126.000 508.300 126.800 508.400 ;
        RECT 116.400 507.700 126.800 508.300 ;
        RECT 116.400 507.600 117.200 507.700 ;
        RECT 126.000 507.600 126.800 507.700 ;
        RECT 164.400 508.300 165.200 508.400 ;
        RECT 185.200 508.300 186.000 508.400 ;
        RECT 190.000 508.300 190.800 508.400 ;
        RECT 164.400 507.700 190.800 508.300 ;
        RECT 164.400 507.600 165.200 507.700 ;
        RECT 185.200 507.600 186.000 507.700 ;
        RECT 190.000 507.600 190.800 507.700 ;
        RECT 239.600 508.300 240.400 508.400 ;
        RECT 246.000 508.300 246.800 508.400 ;
        RECT 239.600 507.700 246.800 508.300 ;
        RECT 239.600 507.600 240.400 507.700 ;
        RECT 246.000 507.600 246.800 507.700 ;
        RECT 247.600 508.300 248.400 508.400 ;
        RECT 262.000 508.300 262.800 508.400 ;
        RECT 247.600 507.700 262.800 508.300 ;
        RECT 247.600 507.600 248.400 507.700 ;
        RECT 262.000 507.600 262.800 507.700 ;
        RECT 289.200 508.300 290.000 508.400 ;
        RECT 297.200 508.300 298.000 508.400 ;
        RECT 289.200 507.700 298.000 508.300 ;
        RECT 289.200 507.600 290.000 507.700 ;
        RECT 297.200 507.600 298.000 507.700 ;
        RECT 327.600 508.300 328.400 508.400 ;
        RECT 332.400 508.300 333.200 508.400 ;
        RECT 353.200 508.300 354.000 508.400 ;
        RECT 396.400 508.300 397.200 508.400 ;
        RECT 327.600 507.700 397.200 508.300 ;
        RECT 327.600 507.600 328.400 507.700 ;
        RECT 332.400 507.600 333.200 507.700 ;
        RECT 353.200 507.600 354.000 507.700 ;
        RECT 396.400 507.600 397.200 507.700 ;
        RECT 414.000 508.300 414.800 508.400 ;
        RECT 423.600 508.300 424.400 508.400 ;
        RECT 414.000 507.700 424.400 508.300 ;
        RECT 414.000 507.600 414.800 507.700 ;
        RECT 423.600 507.600 424.400 507.700 ;
        RECT 428.400 508.300 429.200 508.400 ;
        RECT 436.400 508.300 437.200 508.400 ;
        RECT 428.400 507.700 437.200 508.300 ;
        RECT 428.400 507.600 429.200 507.700 ;
        RECT 436.400 507.600 437.200 507.700 ;
        RECT 439.600 508.300 440.400 508.400 ;
        RECT 454.000 508.300 454.800 508.400 ;
        RECT 439.600 507.700 454.800 508.300 ;
        RECT 439.600 507.600 440.400 507.700 ;
        RECT 454.000 507.600 454.800 507.700 ;
        RECT 487.600 508.300 488.400 508.400 ;
        RECT 521.200 508.300 522.000 508.400 ;
        RECT 487.600 507.700 522.000 508.300 ;
        RECT 487.600 507.600 488.400 507.700 ;
        RECT 521.200 507.600 522.000 507.700 ;
        RECT 526.000 508.300 526.800 508.400 ;
        RECT 527.600 508.300 528.400 508.400 ;
        RECT 526.000 507.700 528.400 508.300 ;
        RECT 526.000 507.600 526.800 507.700 ;
        RECT 527.600 507.600 528.400 507.700 ;
        RECT 543.600 508.300 544.400 508.400 ;
        RECT 572.400 508.300 573.200 508.400 ;
        RECT 575.600 508.300 576.400 508.400 ;
        RECT 543.600 507.700 576.400 508.300 ;
        RECT 543.600 507.600 544.400 507.700 ;
        RECT 572.400 507.600 573.200 507.700 ;
        RECT 575.600 507.600 576.400 507.700 ;
        RECT 41.200 506.300 42.000 506.400 ;
        RECT 49.200 506.300 50.000 506.400 ;
        RECT 41.200 505.700 50.000 506.300 ;
        RECT 41.200 505.600 42.000 505.700 ;
        RECT 49.200 505.600 50.000 505.700 ;
        RECT 119.600 506.300 120.400 506.400 ;
        RECT 130.800 506.300 131.600 506.400 ;
        RECT 138.800 506.300 139.600 506.400 ;
        RECT 166.000 506.300 166.800 506.400 ;
        RECT 119.600 505.700 166.800 506.300 ;
        RECT 119.600 505.600 120.400 505.700 ;
        RECT 130.800 505.600 131.600 505.700 ;
        RECT 138.800 505.600 139.600 505.700 ;
        RECT 166.000 505.600 166.800 505.700 ;
        RECT 167.600 506.300 168.400 506.400 ;
        RECT 174.000 506.300 174.800 506.400 ;
        RECT 167.600 505.700 174.800 506.300 ;
        RECT 167.600 505.600 168.400 505.700 ;
        RECT 174.000 505.600 174.800 505.700 ;
        RECT 238.000 506.300 238.800 506.400 ;
        RECT 241.200 506.300 242.000 506.400 ;
        RECT 238.000 505.700 242.000 506.300 ;
        RECT 238.000 505.600 238.800 505.700 ;
        RECT 241.200 505.600 242.000 505.700 ;
        RECT 247.600 506.300 248.400 506.400 ;
        RECT 252.400 506.300 253.200 506.400 ;
        RECT 247.600 505.700 253.200 506.300 ;
        RECT 247.600 505.600 248.400 505.700 ;
        RECT 252.400 505.600 253.200 505.700 ;
        RECT 265.200 506.300 266.000 506.400 ;
        RECT 300.400 506.300 301.200 506.400 ;
        RECT 319.600 506.300 320.400 506.400 ;
        RECT 265.200 505.700 320.400 506.300 ;
        RECT 265.200 505.600 266.000 505.700 ;
        RECT 300.400 505.600 301.200 505.700 ;
        RECT 319.600 505.600 320.400 505.700 ;
        RECT 335.600 506.300 336.400 506.400 ;
        RECT 434.800 506.300 435.600 506.400 ;
        RECT 335.600 505.700 435.600 506.300 ;
        RECT 335.600 505.600 336.400 505.700 ;
        RECT 434.800 505.600 435.600 505.700 ;
        RECT 463.600 506.300 464.400 506.400 ;
        RECT 471.600 506.300 472.400 506.400 ;
        RECT 463.600 505.700 472.400 506.300 ;
        RECT 463.600 505.600 464.400 505.700 ;
        RECT 471.600 505.600 472.400 505.700 ;
        RECT 479.600 506.300 480.400 506.400 ;
        RECT 500.400 506.300 501.200 506.400 ;
        RECT 479.600 505.700 501.200 506.300 ;
        RECT 479.600 505.600 480.400 505.700 ;
        RECT 500.400 505.600 501.200 505.700 ;
        RECT 519.600 506.300 520.400 506.400 ;
        RECT 522.800 506.300 523.600 506.400 ;
        RECT 519.600 505.700 523.600 506.300 ;
        RECT 519.600 505.600 520.400 505.700 ;
        RECT 522.800 505.600 523.600 505.700 ;
        RECT 535.600 506.300 536.400 506.400 ;
        RECT 561.200 506.300 562.000 506.400 ;
        RECT 535.600 505.700 562.000 506.300 ;
        RECT 535.600 505.600 536.400 505.700 ;
        RECT 561.200 505.600 562.000 505.700 ;
        RECT 1.200 504.300 2.000 504.400 ;
        RECT 6.000 504.300 6.800 504.400 ;
        RECT 1.200 503.700 6.800 504.300 ;
        RECT 1.200 503.600 2.000 503.700 ;
        RECT 6.000 503.600 6.800 503.700 ;
        RECT 73.200 504.300 74.000 504.400 ;
        RECT 90.800 504.300 91.600 504.400 ;
        RECT 73.200 503.700 91.600 504.300 ;
        RECT 73.200 503.600 74.000 503.700 ;
        RECT 90.800 503.600 91.600 503.700 ;
        RECT 94.000 504.300 94.800 504.400 ;
        RECT 100.400 504.300 101.200 504.400 ;
        RECT 94.000 503.700 101.200 504.300 ;
        RECT 94.000 503.600 94.800 503.700 ;
        RECT 100.400 503.600 101.200 503.700 ;
        RECT 124.400 504.300 125.200 504.400 ;
        RECT 150.000 504.300 150.800 504.400 ;
        RECT 169.200 504.300 170.000 504.400 ;
        RECT 124.400 503.700 170.000 504.300 ;
        RECT 124.400 503.600 125.200 503.700 ;
        RECT 150.000 503.600 150.800 503.700 ;
        RECT 169.200 503.600 170.000 503.700 ;
        RECT 225.200 504.300 226.000 504.400 ;
        RECT 231.600 504.300 232.400 504.400 ;
        RECT 236.400 504.300 237.200 504.400 ;
        RECT 225.200 503.700 237.200 504.300 ;
        RECT 225.200 503.600 226.000 503.700 ;
        RECT 231.600 503.600 232.400 503.700 ;
        RECT 236.400 503.600 237.200 503.700 ;
        RECT 295.600 504.300 296.400 504.400 ;
        RECT 354.800 504.300 355.600 504.400 ;
        RECT 295.600 503.700 355.600 504.300 ;
        RECT 295.600 503.600 296.400 503.700 ;
        RECT 354.800 503.600 355.600 503.700 ;
        RECT 378.800 504.300 379.600 504.400 ;
        RECT 422.000 504.300 422.800 504.400 ;
        RECT 378.800 503.700 422.800 504.300 ;
        RECT 378.800 503.600 379.600 503.700 ;
        RECT 422.000 503.600 422.800 503.700 ;
        RECT 449.200 504.300 450.000 504.400 ;
        RECT 470.000 504.300 470.800 504.400 ;
        RECT 487.600 504.300 488.400 504.400 ;
        RECT 449.200 503.700 488.400 504.300 ;
        RECT 449.200 503.600 450.000 503.700 ;
        RECT 470.000 503.600 470.800 503.700 ;
        RECT 487.600 503.600 488.400 503.700 ;
        RECT 506.800 504.300 507.600 504.400 ;
        RECT 529.200 504.300 530.000 504.400 ;
        RECT 538.800 504.300 539.600 504.400 ;
        RECT 506.800 503.700 539.600 504.300 ;
        RECT 506.800 503.600 507.600 503.700 ;
        RECT 529.200 503.600 530.000 503.700 ;
        RECT 538.800 503.600 539.600 503.700 ;
        RECT 18.800 502.300 19.600 502.400 ;
        RECT 74.800 502.300 75.600 502.400 ;
        RECT 18.800 501.700 75.600 502.300 ;
        RECT 18.800 501.600 19.600 501.700 ;
        RECT 74.800 501.600 75.600 501.700 ;
        RECT 170.800 502.300 171.600 502.400 ;
        RECT 172.400 502.300 173.200 502.400 ;
        RECT 170.800 501.700 173.200 502.300 ;
        RECT 170.800 501.600 171.600 501.700 ;
        RECT 172.400 501.600 173.200 501.700 ;
        RECT 223.600 502.300 224.400 502.400 ;
        RECT 247.600 502.300 248.400 502.400 ;
        RECT 223.600 501.700 248.400 502.300 ;
        RECT 223.600 501.600 224.400 501.700 ;
        RECT 247.600 501.600 248.400 501.700 ;
        RECT 314.800 502.300 315.600 502.400 ;
        RECT 383.600 502.300 384.400 502.400 ;
        RECT 314.800 501.700 384.400 502.300 ;
        RECT 314.800 501.600 315.600 501.700 ;
        RECT 383.600 501.600 384.400 501.700 ;
        RECT 391.600 502.300 392.400 502.400 ;
        RECT 404.400 502.300 405.200 502.400 ;
        RECT 391.600 501.700 405.200 502.300 ;
        RECT 391.600 501.600 392.400 501.700 ;
        RECT 404.400 501.600 405.200 501.700 ;
        RECT 422.000 502.300 422.800 502.400 ;
        RECT 455.600 502.300 456.400 502.400 ;
        RECT 422.000 501.700 456.400 502.300 ;
        RECT 422.000 501.600 422.800 501.700 ;
        RECT 455.600 501.600 456.400 501.700 ;
        RECT 490.800 502.300 491.600 502.400 ;
        RECT 532.400 502.300 533.200 502.400 ;
        RECT 490.800 501.700 533.200 502.300 ;
        RECT 490.800 501.600 491.600 501.700 ;
        RECT 532.400 501.600 533.200 501.700 ;
        RECT 15.600 500.300 16.400 500.400 ;
        RECT 46.000 500.300 46.800 500.400 ;
        RECT 15.600 499.700 46.800 500.300 ;
        RECT 15.600 499.600 16.400 499.700 ;
        RECT 46.000 499.600 46.800 499.700 ;
        RECT 66.800 500.300 67.600 500.400 ;
        RECT 84.400 500.300 85.200 500.400 ;
        RECT 92.400 500.300 93.200 500.400 ;
        RECT 66.800 499.700 93.200 500.300 ;
        RECT 66.800 499.600 67.600 499.700 ;
        RECT 84.400 499.600 85.200 499.700 ;
        RECT 92.400 499.600 93.200 499.700 ;
        RECT 105.200 500.300 106.000 500.400 ;
        RECT 113.200 500.300 114.000 500.400 ;
        RECT 105.200 499.700 114.000 500.300 ;
        RECT 105.200 499.600 106.000 499.700 ;
        RECT 113.200 499.600 114.000 499.700 ;
        RECT 129.200 500.300 130.000 500.400 ;
        RECT 140.400 500.300 141.200 500.400 ;
        RECT 129.200 499.700 141.200 500.300 ;
        RECT 129.200 499.600 130.000 499.700 ;
        RECT 140.400 499.600 141.200 499.700 ;
        RECT 191.600 500.300 192.400 500.400 ;
        RECT 196.400 500.300 197.200 500.400 ;
        RECT 215.600 500.300 216.400 500.400 ;
        RECT 191.600 499.700 216.400 500.300 ;
        RECT 191.600 499.600 192.400 499.700 ;
        RECT 196.400 499.600 197.200 499.700 ;
        RECT 215.600 499.600 216.400 499.700 ;
        RECT 342.000 500.300 342.800 500.400 ;
        RECT 351.600 500.300 352.400 500.400 ;
        RECT 342.000 499.700 352.400 500.300 ;
        RECT 342.000 499.600 342.800 499.700 ;
        RECT 351.600 499.600 352.400 499.700 ;
        RECT 391.600 500.300 392.400 500.400 ;
        RECT 393.200 500.300 394.000 500.400 ;
        RECT 391.600 499.700 394.000 500.300 ;
        RECT 391.600 499.600 392.400 499.700 ;
        RECT 393.200 499.600 394.000 499.700 ;
        RECT 508.400 500.300 509.200 500.400 ;
        RECT 518.000 500.300 518.800 500.400 ;
        RECT 537.200 500.300 538.000 500.400 ;
        RECT 543.600 500.300 544.400 500.400 ;
        RECT 508.400 499.700 544.400 500.300 ;
        RECT 508.400 499.600 509.200 499.700 ;
        RECT 518.000 499.600 518.800 499.700 ;
        RECT 537.200 499.600 538.000 499.700 ;
        RECT 543.600 499.600 544.400 499.700 ;
        RECT 567.600 500.300 568.400 500.400 ;
        RECT 591.600 500.300 592.400 500.400 ;
        RECT 594.800 500.300 595.600 500.400 ;
        RECT 567.600 499.700 595.600 500.300 ;
        RECT 567.600 499.600 568.400 499.700 ;
        RECT 591.600 499.600 592.400 499.700 ;
        RECT 594.800 499.600 595.600 499.700 ;
        RECT 55.600 498.300 56.400 498.400 ;
        RECT 106.800 498.300 107.600 498.400 ;
        RECT 55.600 497.700 107.600 498.300 ;
        RECT 55.600 497.600 56.400 497.700 ;
        RECT 106.800 497.600 107.600 497.700 ;
        RECT 182.000 498.300 182.800 498.400 ;
        RECT 225.200 498.300 226.000 498.400 ;
        RECT 244.400 498.300 245.200 498.400 ;
        RECT 182.000 497.700 245.200 498.300 ;
        RECT 182.000 497.600 182.800 497.700 ;
        RECT 225.200 497.600 226.000 497.700 ;
        RECT 244.400 497.600 245.200 497.700 ;
        RECT 281.200 498.300 282.000 498.400 ;
        RECT 294.000 498.300 294.800 498.400 ;
        RECT 281.200 497.700 294.800 498.300 ;
        RECT 281.200 497.600 282.000 497.700 ;
        RECT 294.000 497.600 294.800 497.700 ;
        RECT 302.000 498.300 302.800 498.400 ;
        RECT 319.600 498.300 320.400 498.400 ;
        RECT 302.000 497.700 320.400 498.300 ;
        RECT 302.000 497.600 302.800 497.700 ;
        RECT 319.600 497.600 320.400 497.700 ;
        RECT 330.800 497.600 331.600 498.400 ;
        RECT 383.600 498.300 384.400 498.400 ;
        RECT 433.200 498.300 434.000 498.400 ;
        RECT 447.600 498.300 448.400 498.400 ;
        RECT 383.600 497.700 448.400 498.300 ;
        RECT 383.600 497.600 384.400 497.700 ;
        RECT 433.200 497.600 434.000 497.700 ;
        RECT 447.600 497.600 448.400 497.700 ;
        RECT 452.400 498.300 453.200 498.400 ;
        RECT 476.400 498.300 477.200 498.400 ;
        RECT 495.600 498.300 496.400 498.400 ;
        RECT 506.800 498.300 507.600 498.400 ;
        RECT 452.400 497.700 507.600 498.300 ;
        RECT 452.400 497.600 453.200 497.700 ;
        RECT 476.400 497.600 477.200 497.700 ;
        RECT 495.600 497.600 496.400 497.700 ;
        RECT 506.800 497.600 507.600 497.700 ;
        RECT 516.400 498.300 517.200 498.400 ;
        RECT 527.600 498.300 528.400 498.400 ;
        RECT 516.400 497.700 528.400 498.300 ;
        RECT 516.400 497.600 517.200 497.700 ;
        RECT 527.600 497.600 528.400 497.700 ;
        RECT 34.800 496.300 35.600 496.400 ;
        RECT 65.200 496.300 66.000 496.400 ;
        RECT 90.800 496.300 91.600 496.400 ;
        RECT 127.600 496.300 128.400 496.400 ;
        RECT 34.800 495.700 128.400 496.300 ;
        RECT 34.800 495.600 35.600 495.700 ;
        RECT 65.200 495.600 66.000 495.700 ;
        RECT 90.800 495.600 91.600 495.700 ;
        RECT 127.600 495.600 128.400 495.700 ;
        RECT 201.200 496.300 202.000 496.400 ;
        RECT 226.800 496.300 227.600 496.400 ;
        RECT 244.400 496.300 245.200 496.400 ;
        RECT 250.800 496.300 251.600 496.400 ;
        RECT 201.200 495.700 251.600 496.300 ;
        RECT 201.200 495.600 202.000 495.700 ;
        RECT 226.800 495.600 227.600 495.700 ;
        RECT 244.400 495.600 245.200 495.700 ;
        RECT 250.800 495.600 251.600 495.700 ;
        RECT 295.600 496.300 296.400 496.400 ;
        RECT 314.800 496.300 315.600 496.400 ;
        RECT 295.600 495.700 315.600 496.300 ;
        RECT 295.600 495.600 296.400 495.700 ;
        RECT 314.800 495.600 315.600 495.700 ;
        RECT 319.600 496.300 320.400 496.400 ;
        RECT 324.400 496.300 325.200 496.400 ;
        RECT 358.000 496.300 358.800 496.400 ;
        RECT 386.800 496.300 387.600 496.400 ;
        RECT 319.600 495.700 387.600 496.300 ;
        RECT 319.600 495.600 320.400 495.700 ;
        RECT 324.400 495.600 325.200 495.700 ;
        RECT 358.000 495.600 358.800 495.700 ;
        RECT 386.800 495.600 387.600 495.700 ;
        RECT 393.200 496.300 394.000 496.400 ;
        RECT 418.800 496.300 419.600 496.400 ;
        RECT 393.200 495.700 419.600 496.300 ;
        RECT 393.200 495.600 394.000 495.700 ;
        RECT 418.800 495.600 419.600 495.700 ;
        RECT 420.400 496.300 421.200 496.400 ;
        RECT 447.600 496.300 448.400 496.400 ;
        RECT 420.400 495.700 448.400 496.300 ;
        RECT 420.400 495.600 421.200 495.700 ;
        RECT 447.600 495.600 448.400 495.700 ;
        RECT 454.000 496.300 454.800 496.400 ;
        RECT 457.200 496.300 458.000 496.400 ;
        RECT 454.000 495.700 458.000 496.300 ;
        RECT 454.000 495.600 454.800 495.700 ;
        RECT 457.200 495.600 458.000 495.700 ;
        RECT 471.600 496.300 472.400 496.400 ;
        RECT 489.200 496.300 490.000 496.400 ;
        RECT 471.600 495.700 490.000 496.300 ;
        RECT 471.600 495.600 472.400 495.700 ;
        RECT 489.200 495.600 490.000 495.700 ;
        RECT 503.600 495.600 504.400 496.400 ;
        RECT 511.600 496.300 512.400 496.400 ;
        RECT 529.200 496.300 530.000 496.400 ;
        RECT 511.600 495.700 530.000 496.300 ;
        RECT 511.600 495.600 512.400 495.700 ;
        RECT 529.200 495.600 530.000 495.700 ;
        RECT 543.600 496.300 544.400 496.400 ;
        RECT 562.800 496.300 563.600 496.400 ;
        RECT 543.600 495.700 563.600 496.300 ;
        RECT 543.600 495.600 544.400 495.700 ;
        RECT 562.800 495.600 563.600 495.700 ;
        RECT 44.400 494.300 45.200 494.400 ;
        RECT 49.200 494.300 50.000 494.400 ;
        RECT 44.400 493.700 50.000 494.300 ;
        RECT 44.400 493.600 45.200 493.700 ;
        RECT 49.200 493.600 50.000 493.700 ;
        RECT 63.600 494.300 64.400 494.400 ;
        RECT 87.600 494.300 88.400 494.400 ;
        RECT 97.200 494.300 98.000 494.400 ;
        RECT 63.600 493.700 98.000 494.300 ;
        RECT 63.600 493.600 64.400 493.700 ;
        RECT 87.600 493.600 88.400 493.700 ;
        RECT 97.200 493.600 98.000 493.700 ;
        RECT 102.000 494.300 102.800 494.400 ;
        RECT 111.600 494.300 112.400 494.400 ;
        RECT 102.000 493.700 112.400 494.300 ;
        RECT 102.000 493.600 102.800 493.700 ;
        RECT 111.600 493.600 112.400 493.700 ;
        RECT 150.000 494.300 150.800 494.400 ;
        RECT 177.200 494.300 178.000 494.400 ;
        RECT 150.000 493.700 178.000 494.300 ;
        RECT 150.000 493.600 150.800 493.700 ;
        RECT 177.200 493.600 178.000 493.700 ;
        RECT 194.800 494.300 195.600 494.400 ;
        RECT 214.000 494.300 214.800 494.400 ;
        RECT 194.800 493.700 214.800 494.300 ;
        RECT 194.800 493.600 195.600 493.700 ;
        RECT 214.000 493.600 214.800 493.700 ;
        RECT 263.600 494.300 264.400 494.400 ;
        RECT 276.400 494.300 277.200 494.400 ;
        RECT 278.000 494.300 278.800 494.400 ;
        RECT 263.600 493.700 278.800 494.300 ;
        RECT 263.600 493.600 264.400 493.700 ;
        RECT 276.400 493.600 277.200 493.700 ;
        RECT 278.000 493.600 278.800 493.700 ;
        RECT 281.200 494.300 282.000 494.400 ;
        RECT 286.000 494.300 286.800 494.400 ;
        RECT 281.200 493.700 286.800 494.300 ;
        RECT 281.200 493.600 282.000 493.700 ;
        RECT 286.000 493.600 286.800 493.700 ;
        RECT 290.800 494.300 291.600 494.400 ;
        RECT 297.200 494.300 298.000 494.400 ;
        RECT 334.000 494.300 334.800 494.400 ;
        RECT 290.800 493.700 334.800 494.300 ;
        RECT 290.800 493.600 291.600 493.700 ;
        RECT 297.200 493.600 298.000 493.700 ;
        RECT 334.000 493.600 334.800 493.700 ;
        RECT 346.800 494.300 347.600 494.400 ;
        RECT 369.200 494.300 370.000 494.400 ;
        RECT 346.800 493.700 370.000 494.300 ;
        RECT 346.800 493.600 347.600 493.700 ;
        RECT 369.200 493.600 370.000 493.700 ;
        RECT 396.400 494.300 397.200 494.400 ;
        RECT 473.200 494.300 474.000 494.400 ;
        RECT 479.600 494.300 480.400 494.400 ;
        RECT 396.400 493.700 480.400 494.300 ;
        RECT 396.400 493.600 397.200 493.700 ;
        RECT 473.200 493.600 474.000 493.700 ;
        RECT 479.600 493.600 480.400 493.700 ;
        RECT 500.400 494.300 501.200 494.400 ;
        RECT 558.000 494.300 558.800 494.400 ;
        RECT 574.000 494.300 574.800 494.400 ;
        RECT 500.400 493.700 574.800 494.300 ;
        RECT 500.400 493.600 501.200 493.700 ;
        RECT 558.000 493.600 558.800 493.700 ;
        RECT 574.000 493.600 574.800 493.700 ;
        RECT 1.200 492.300 2.000 492.400 ;
        RECT 17.200 492.300 18.000 492.400 ;
        RECT 1.200 491.700 18.000 492.300 ;
        RECT 1.200 491.600 2.000 491.700 ;
        RECT 17.200 491.600 18.000 491.700 ;
        RECT 30.000 492.300 30.800 492.400 ;
        RECT 46.000 492.300 46.800 492.400 ;
        RECT 30.000 491.700 46.800 492.300 ;
        RECT 30.000 491.600 30.800 491.700 ;
        RECT 46.000 491.600 46.800 491.700 ;
        RECT 47.600 492.300 48.400 492.400 ;
        RECT 58.800 492.300 59.600 492.400 ;
        RECT 47.600 491.700 59.600 492.300 ;
        RECT 47.600 491.600 48.400 491.700 ;
        RECT 58.800 491.600 59.600 491.700 ;
        RECT 62.000 492.300 62.800 492.400 ;
        RECT 87.600 492.300 88.400 492.400 ;
        RECT 89.200 492.300 90.000 492.400 ;
        RECT 62.000 491.700 90.000 492.300 ;
        RECT 62.000 491.600 62.800 491.700 ;
        RECT 87.600 491.600 88.400 491.700 ;
        RECT 89.200 491.600 90.000 491.700 ;
        RECT 103.600 492.300 104.400 492.400 ;
        RECT 116.400 492.300 117.200 492.400 ;
        RECT 146.800 492.300 147.600 492.400 ;
        RECT 103.600 491.700 147.600 492.300 ;
        RECT 103.600 491.600 104.400 491.700 ;
        RECT 116.400 491.600 117.200 491.700 ;
        RECT 146.800 491.600 147.600 491.700 ;
        RECT 159.600 492.300 160.400 492.400 ;
        RECT 183.600 492.300 184.400 492.400 ;
        RECT 159.600 491.700 184.400 492.300 ;
        RECT 159.600 491.600 160.400 491.700 ;
        RECT 183.600 491.600 184.400 491.700 ;
        RECT 282.800 492.300 283.600 492.400 ;
        RECT 298.800 492.300 299.600 492.400 ;
        RECT 282.800 491.700 299.600 492.300 ;
        RECT 282.800 491.600 283.600 491.700 ;
        RECT 298.800 491.600 299.600 491.700 ;
        RECT 311.600 492.300 312.400 492.400 ;
        RECT 326.000 492.300 326.800 492.400 ;
        RECT 311.600 491.700 326.800 492.300 ;
        RECT 311.600 491.600 312.400 491.700 ;
        RECT 326.000 491.600 326.800 491.700 ;
        RECT 332.400 492.300 333.200 492.400 ;
        RECT 335.600 492.300 336.400 492.400 ;
        RECT 332.400 491.700 336.400 492.300 ;
        RECT 332.400 491.600 333.200 491.700 ;
        RECT 335.600 491.600 336.400 491.700 ;
        RECT 340.400 492.300 341.200 492.400 ;
        RECT 345.200 492.300 346.000 492.400 ;
        RECT 340.400 491.700 346.000 492.300 ;
        RECT 340.400 491.600 341.200 491.700 ;
        RECT 345.200 491.600 346.000 491.700 ;
        RECT 351.600 492.300 352.400 492.400 ;
        RECT 359.600 492.300 360.400 492.400 ;
        RECT 351.600 491.700 360.400 492.300 ;
        RECT 351.600 491.600 352.400 491.700 ;
        RECT 359.600 491.600 360.400 491.700 ;
        RECT 374.000 492.300 374.800 492.400 ;
        RECT 401.200 492.300 402.000 492.400 ;
        RECT 374.000 491.700 402.000 492.300 ;
        RECT 374.000 491.600 374.800 491.700 ;
        RECT 401.200 491.600 402.000 491.700 ;
        RECT 409.200 492.300 410.000 492.400 ;
        RECT 444.400 492.300 445.200 492.400 ;
        RECT 466.800 492.300 467.600 492.400 ;
        RECT 516.400 492.300 517.200 492.400 ;
        RECT 546.800 492.300 547.600 492.400 ;
        RECT 409.200 491.700 547.600 492.300 ;
        RECT 409.200 491.600 410.000 491.700 ;
        RECT 444.400 491.600 445.200 491.700 ;
        RECT 466.800 491.600 467.600 491.700 ;
        RECT 516.400 491.600 517.200 491.700 ;
        RECT 546.800 491.600 547.600 491.700 ;
        RECT 572.400 492.300 573.200 492.400 ;
        RECT 598.000 492.300 598.800 492.400 ;
        RECT 572.400 491.700 598.800 492.300 ;
        RECT 572.400 491.600 573.200 491.700 ;
        RECT 598.000 491.600 598.800 491.700 ;
        RECT 103.700 490.400 104.300 491.600 ;
        RECT 14.000 490.300 14.800 490.400 ;
        RECT 17.200 490.300 18.000 490.400 ;
        RECT 14.000 489.700 18.000 490.300 ;
        RECT 14.000 489.600 14.800 489.700 ;
        RECT 17.200 489.600 18.000 489.700 ;
        RECT 20.400 490.300 21.200 490.400 ;
        RECT 30.000 490.300 30.800 490.400 ;
        RECT 20.400 489.700 30.800 490.300 ;
        RECT 20.400 489.600 21.200 489.700 ;
        RECT 30.000 489.600 30.800 489.700 ;
        RECT 41.200 490.300 42.000 490.400 ;
        RECT 55.600 490.300 56.400 490.400 ;
        RECT 58.800 490.300 59.600 490.400 ;
        RECT 41.200 489.700 59.600 490.300 ;
        RECT 41.200 489.600 42.000 489.700 ;
        RECT 55.600 489.600 56.400 489.700 ;
        RECT 58.800 489.600 59.600 489.700 ;
        RECT 65.200 490.300 66.000 490.400 ;
        RECT 74.800 490.300 75.600 490.400 ;
        RECT 65.200 489.700 75.600 490.300 ;
        RECT 65.200 489.600 66.000 489.700 ;
        RECT 74.800 489.600 75.600 489.700 ;
        RECT 78.000 490.300 78.800 490.400 ;
        RECT 82.800 490.300 83.600 490.400 ;
        RECT 78.000 489.700 83.600 490.300 ;
        RECT 78.000 489.600 78.800 489.700 ;
        RECT 82.800 489.600 83.600 489.700 ;
        RECT 84.400 490.300 85.200 490.400 ;
        RECT 100.400 490.300 101.200 490.400 ;
        RECT 84.400 489.700 101.200 490.300 ;
        RECT 84.400 489.600 85.200 489.700 ;
        RECT 100.400 489.600 101.200 489.700 ;
        RECT 103.600 489.600 104.400 490.400 ;
        RECT 295.600 489.600 296.400 490.400 ;
        RECT 310.000 490.300 310.800 490.400 ;
        RECT 342.000 490.300 342.800 490.400 ;
        RECT 310.000 489.700 342.800 490.300 ;
        RECT 310.000 489.600 310.800 489.700 ;
        RECT 342.000 489.600 342.800 489.700 ;
        RECT 356.400 490.300 357.200 490.400 ;
        RECT 378.800 490.300 379.600 490.400 ;
        RECT 356.400 489.700 379.600 490.300 ;
        RECT 356.400 489.600 357.200 489.700 ;
        RECT 378.800 489.600 379.600 489.700 ;
        RECT 386.800 490.300 387.600 490.400 ;
        RECT 399.600 490.300 400.400 490.400 ;
        RECT 426.800 490.300 427.600 490.400 ;
        RECT 386.800 489.700 427.600 490.300 ;
        RECT 386.800 489.600 387.600 489.700 ;
        RECT 399.600 489.600 400.400 489.700 ;
        RECT 426.800 489.600 427.600 489.700 ;
        RECT 455.600 490.300 456.400 490.400 ;
        RECT 466.800 490.300 467.600 490.400 ;
        RECT 455.600 489.700 467.600 490.300 ;
        RECT 455.600 489.600 456.400 489.700 ;
        RECT 466.800 489.600 467.600 489.700 ;
        RECT 474.800 490.300 475.600 490.400 ;
        RECT 489.200 490.300 490.000 490.400 ;
        RECT 474.800 489.700 490.000 490.300 ;
        RECT 474.800 489.600 475.600 489.700 ;
        RECT 489.200 489.600 490.000 489.700 ;
        RECT 497.200 490.300 498.000 490.400 ;
        RECT 506.800 490.300 507.600 490.400 ;
        RECT 497.200 489.700 507.600 490.300 ;
        RECT 497.200 489.600 498.000 489.700 ;
        RECT 506.800 489.600 507.600 489.700 ;
        RECT 511.600 490.300 512.400 490.400 ;
        RECT 521.200 490.300 522.000 490.400 ;
        RECT 511.600 489.700 522.000 490.300 ;
        RECT 511.600 489.600 512.400 489.700 ;
        RECT 521.200 489.600 522.000 489.700 ;
        RECT 543.600 490.300 544.400 490.400 ;
        RECT 546.800 490.300 547.600 490.400 ;
        RECT 543.600 489.700 547.600 490.300 ;
        RECT 543.600 489.600 544.400 489.700 ;
        RECT 546.800 489.600 547.600 489.700 ;
        RECT 52.400 488.300 53.200 488.400 ;
        RECT 65.200 488.300 66.000 488.400 ;
        RECT 52.400 487.700 66.000 488.300 ;
        RECT 52.400 487.600 53.200 487.700 ;
        RECT 65.200 487.600 66.000 487.700 ;
        RECT 81.200 488.300 82.000 488.400 ;
        RECT 113.200 488.300 114.000 488.400 ;
        RECT 81.200 487.700 114.000 488.300 ;
        RECT 81.200 487.600 82.000 487.700 ;
        RECT 113.200 487.600 114.000 487.700 ;
        RECT 246.000 488.300 246.800 488.400 ;
        RECT 284.400 488.300 285.200 488.400 ;
        RECT 300.400 488.300 301.200 488.400 ;
        RECT 246.000 487.700 301.200 488.300 ;
        RECT 246.000 487.600 246.800 487.700 ;
        RECT 284.400 487.600 285.200 487.700 ;
        RECT 300.400 487.600 301.200 487.700 ;
        RECT 329.200 488.300 330.000 488.400 ;
        RECT 345.200 488.300 346.000 488.400 ;
        RECT 329.200 487.700 346.000 488.300 ;
        RECT 329.200 487.600 330.000 487.700 ;
        RECT 345.200 487.600 346.000 487.700 ;
        RECT 354.800 488.300 355.600 488.400 ;
        RECT 364.400 488.300 365.200 488.400 ;
        RECT 354.800 487.700 365.200 488.300 ;
        RECT 354.800 487.600 355.600 487.700 ;
        RECT 364.400 487.600 365.200 487.700 ;
        RECT 377.200 488.300 378.000 488.400 ;
        RECT 380.400 488.300 381.200 488.400 ;
        RECT 406.000 488.300 406.800 488.400 ;
        RECT 377.200 487.700 406.800 488.300 ;
        RECT 377.200 487.600 378.000 487.700 ;
        RECT 380.400 487.600 381.200 487.700 ;
        RECT 406.000 487.600 406.800 487.700 ;
        RECT 430.000 488.300 430.800 488.400 ;
        RECT 446.000 488.300 446.800 488.400 ;
        RECT 430.000 487.700 446.800 488.300 ;
        RECT 430.000 487.600 430.800 487.700 ;
        RECT 446.000 487.600 446.800 487.700 ;
        RECT 470.000 488.300 470.800 488.400 ;
        RECT 478.000 488.300 478.800 488.400 ;
        RECT 470.000 487.700 478.800 488.300 ;
        RECT 470.000 487.600 470.800 487.700 ;
        RECT 478.000 487.600 478.800 487.700 ;
        RECT 498.800 488.300 499.600 488.400 ;
        RECT 502.000 488.300 502.800 488.400 ;
        RECT 498.800 487.700 502.800 488.300 ;
        RECT 498.800 487.600 499.600 487.700 ;
        RECT 502.000 487.600 502.800 487.700 ;
        RECT 503.600 488.300 504.400 488.400 ;
        RECT 513.200 488.300 514.000 488.400 ;
        RECT 519.600 488.300 520.400 488.400 ;
        RECT 503.600 487.700 520.400 488.300 ;
        RECT 503.600 487.600 504.400 487.700 ;
        RECT 513.200 487.600 514.000 487.700 ;
        RECT 519.600 487.600 520.400 487.700 ;
        RECT 6.000 486.300 6.800 486.400 ;
        RECT 20.400 486.300 21.200 486.400 ;
        RECT 39.600 486.300 40.400 486.400 ;
        RECT 42.800 486.300 43.600 486.400 ;
        RECT 73.200 486.300 74.000 486.400 ;
        RECT 6.000 485.700 74.000 486.300 ;
        RECT 6.000 485.600 6.800 485.700 ;
        RECT 20.400 485.600 21.200 485.700 ;
        RECT 39.600 485.600 40.400 485.700 ;
        RECT 42.800 485.600 43.600 485.700 ;
        RECT 73.200 485.600 74.000 485.700 ;
        RECT 103.600 486.300 104.400 486.400 ;
        RECT 196.400 486.300 197.200 486.400 ;
        RECT 103.600 485.700 197.200 486.300 ;
        RECT 103.600 485.600 104.400 485.700 ;
        RECT 196.400 485.600 197.200 485.700 ;
        RECT 284.400 486.300 285.200 486.400 ;
        RECT 292.400 486.300 293.200 486.400 ;
        RECT 284.400 485.700 293.200 486.300 ;
        RECT 284.400 485.600 285.200 485.700 ;
        RECT 292.400 485.600 293.200 485.700 ;
        RECT 322.800 486.300 323.600 486.400 ;
        RECT 337.200 486.300 338.000 486.400 ;
        RECT 410.800 486.300 411.600 486.400 ;
        RECT 322.800 485.700 411.600 486.300 ;
        RECT 322.800 485.600 323.600 485.700 ;
        RECT 337.200 485.600 338.000 485.700 ;
        RECT 410.800 485.600 411.600 485.700 ;
        RECT 430.000 486.300 430.800 486.400 ;
        RECT 439.600 486.300 440.400 486.400 ;
        RECT 430.000 485.700 440.400 486.300 ;
        RECT 430.000 485.600 430.800 485.700 ;
        RECT 439.600 485.600 440.400 485.700 ;
        RECT 15.600 484.300 16.400 484.400 ;
        RECT 17.200 484.300 18.000 484.400 ;
        RECT 15.600 483.700 18.000 484.300 ;
        RECT 15.600 483.600 16.400 483.700 ;
        RECT 17.200 483.600 18.000 483.700 ;
        RECT 47.600 484.300 48.400 484.400 ;
        RECT 71.600 484.300 72.400 484.400 ;
        RECT 47.600 483.700 72.400 484.300 ;
        RECT 47.600 483.600 48.400 483.700 ;
        RECT 71.600 483.600 72.400 483.700 ;
        RECT 87.600 484.300 88.400 484.400 ;
        RECT 121.200 484.300 122.000 484.400 ;
        RECT 87.600 483.700 122.000 484.300 ;
        RECT 87.600 483.600 88.400 483.700 ;
        RECT 121.200 483.600 122.000 483.700 ;
        RECT 212.400 484.300 213.200 484.400 ;
        RECT 225.200 484.300 226.000 484.400 ;
        RECT 212.400 483.700 226.000 484.300 ;
        RECT 212.400 483.600 213.200 483.700 ;
        RECT 225.200 483.600 226.000 483.700 ;
        RECT 330.800 484.300 331.600 484.400 ;
        RECT 335.600 484.300 336.400 484.400 ;
        RECT 330.800 483.700 336.400 484.300 ;
        RECT 330.800 483.600 331.600 483.700 ;
        RECT 335.600 483.600 336.400 483.700 ;
        RECT 343.600 484.300 344.400 484.400 ;
        RECT 372.400 484.300 373.200 484.400 ;
        RECT 343.600 483.700 373.200 484.300 ;
        RECT 343.600 483.600 344.400 483.700 ;
        RECT 372.400 483.600 373.200 483.700 ;
        RECT 406.000 484.300 406.800 484.400 ;
        RECT 425.200 484.300 426.000 484.400 ;
        RECT 406.000 483.700 426.000 484.300 ;
        RECT 406.000 483.600 406.800 483.700 ;
        RECT 425.200 483.600 426.000 483.700 ;
        RECT 426.800 484.300 427.600 484.400 ;
        RECT 454.000 484.300 454.800 484.400 ;
        RECT 426.800 483.700 454.800 484.300 ;
        RECT 426.800 483.600 427.600 483.700 ;
        RECT 454.000 483.600 454.800 483.700 ;
        RECT 455.600 484.300 456.400 484.400 ;
        RECT 492.400 484.300 493.200 484.400 ;
        RECT 455.600 483.700 493.200 484.300 ;
        RECT 455.600 483.600 456.400 483.700 ;
        RECT 492.400 483.600 493.200 483.700 ;
        RECT 494.000 484.300 494.800 484.400 ;
        RECT 516.400 484.300 517.200 484.400 ;
        RECT 519.600 484.300 520.400 484.400 ;
        RECT 494.000 483.700 520.400 484.300 ;
        RECT 494.000 483.600 494.800 483.700 ;
        RECT 516.400 483.600 517.200 483.700 ;
        RECT 519.600 483.600 520.400 483.700 ;
        RECT 524.400 484.300 525.200 484.400 ;
        RECT 540.400 484.300 541.200 484.400 ;
        RECT 524.400 483.700 541.200 484.300 ;
        RECT 524.400 483.600 525.200 483.700 ;
        RECT 540.400 483.600 541.200 483.700 ;
        RECT 578.800 484.300 579.600 484.400 ;
        RECT 602.800 484.300 603.600 484.400 ;
        RECT 578.800 483.700 603.600 484.300 ;
        RECT 578.800 483.600 579.600 483.700 ;
        RECT 602.800 483.600 603.600 483.700 ;
        RECT 57.200 482.300 58.000 482.400 ;
        RECT 73.200 482.300 74.000 482.400 ;
        RECT 57.200 481.700 74.000 482.300 ;
        RECT 57.200 481.600 58.000 481.700 ;
        RECT 73.200 481.600 74.000 481.700 ;
        RECT 86.000 482.300 86.800 482.400 ;
        RECT 92.400 482.300 93.200 482.400 ;
        RECT 102.000 482.300 102.800 482.400 ;
        RECT 86.000 481.700 91.500 482.300 ;
        RECT 86.000 481.600 86.800 481.700 ;
        RECT 22.000 480.300 22.800 480.400 ;
        RECT 31.600 480.300 32.400 480.400 ;
        RECT 22.000 479.700 32.400 480.300 ;
        RECT 22.000 479.600 22.800 479.700 ;
        RECT 31.600 479.600 32.400 479.700 ;
        RECT 71.600 480.300 72.400 480.400 ;
        RECT 86.000 480.300 86.800 480.400 ;
        RECT 71.600 479.700 86.800 480.300 ;
        RECT 90.900 480.300 91.500 481.700 ;
        RECT 92.400 481.700 102.800 482.300 ;
        RECT 92.400 481.600 93.200 481.700 ;
        RECT 102.000 481.600 102.800 481.700 ;
        RECT 298.800 482.300 299.600 482.400 ;
        RECT 449.200 482.300 450.000 482.400 ;
        RECT 298.800 481.700 450.000 482.300 ;
        RECT 298.800 481.600 299.600 481.700 ;
        RECT 449.200 481.600 450.000 481.700 ;
        RECT 465.200 482.300 466.000 482.400 ;
        RECT 471.600 482.300 472.400 482.400 ;
        RECT 465.200 481.700 472.400 482.300 ;
        RECT 465.200 481.600 466.000 481.700 ;
        RECT 471.600 481.600 472.400 481.700 ;
        RECT 478.000 482.300 478.800 482.400 ;
        RECT 495.600 482.300 496.400 482.400 ;
        RECT 478.000 481.700 496.400 482.300 ;
        RECT 478.000 481.600 478.800 481.700 ;
        RECT 495.600 481.600 496.400 481.700 ;
        RECT 116.400 480.300 117.200 480.400 ;
        RECT 135.600 480.300 136.400 480.400 ;
        RECT 90.900 479.700 115.500 480.300 ;
        RECT 71.600 479.600 72.400 479.700 ;
        RECT 86.000 479.600 86.800 479.700 ;
        RECT 82.800 478.300 83.600 478.400 ;
        RECT 97.200 478.300 98.000 478.400 ;
        RECT 82.800 477.700 98.000 478.300 ;
        RECT 114.900 478.300 115.500 479.700 ;
        RECT 116.400 479.700 136.400 480.300 ;
        RECT 116.400 479.600 117.200 479.700 ;
        RECT 135.600 479.600 136.400 479.700 ;
        RECT 356.400 480.300 357.200 480.400 ;
        RECT 370.800 480.300 371.600 480.400 ;
        RECT 356.400 479.700 371.600 480.300 ;
        RECT 356.400 479.600 357.200 479.700 ;
        RECT 370.800 479.600 371.600 479.700 ;
        RECT 391.600 480.300 392.400 480.400 ;
        RECT 398.000 480.300 398.800 480.400 ;
        RECT 391.600 479.700 398.800 480.300 ;
        RECT 391.600 479.600 392.400 479.700 ;
        RECT 398.000 479.600 398.800 479.700 ;
        RECT 426.800 480.300 427.600 480.400 ;
        RECT 430.000 480.300 430.800 480.400 ;
        RECT 426.800 479.700 430.800 480.300 ;
        RECT 426.800 479.600 427.600 479.700 ;
        RECT 430.000 479.600 430.800 479.700 ;
        RECT 433.200 480.300 434.000 480.400 ;
        RECT 447.600 480.300 448.400 480.400 ;
        RECT 433.200 479.700 448.400 480.300 ;
        RECT 433.200 479.600 434.000 479.700 ;
        RECT 447.600 479.600 448.400 479.700 ;
        RECT 145.200 478.300 146.000 478.400 ;
        RECT 114.900 477.700 146.000 478.300 ;
        RECT 82.800 477.600 83.600 477.700 ;
        RECT 97.200 477.600 98.000 477.700 ;
        RECT 145.200 477.600 146.000 477.700 ;
        RECT 366.000 478.300 366.800 478.400 ;
        RECT 375.600 478.300 376.400 478.400 ;
        RECT 407.600 478.300 408.400 478.400 ;
        RECT 449.200 478.300 450.000 478.400 ;
        RECT 366.000 477.700 450.000 478.300 ;
        RECT 366.000 477.600 366.800 477.700 ;
        RECT 375.600 477.600 376.400 477.700 ;
        RECT 407.600 477.600 408.400 477.700 ;
        RECT 449.200 477.600 450.000 477.700 ;
        RECT 466.800 478.300 467.600 478.400 ;
        RECT 494.000 478.300 494.800 478.400 ;
        RECT 466.800 477.700 494.800 478.300 ;
        RECT 466.800 477.600 467.600 477.700 ;
        RECT 494.000 477.600 494.800 477.700 ;
        RECT 50.800 476.300 51.600 476.400 ;
        RECT 57.200 476.300 58.000 476.400 ;
        RECT 50.800 475.700 58.000 476.300 ;
        RECT 50.800 475.600 51.600 475.700 ;
        RECT 57.200 475.600 58.000 475.700 ;
        RECT 111.600 476.300 112.400 476.400 ;
        RECT 121.200 476.300 122.000 476.400 ;
        RECT 111.600 475.700 122.000 476.300 ;
        RECT 111.600 475.600 112.400 475.700 ;
        RECT 121.200 475.600 122.000 475.700 ;
        RECT 124.400 476.300 125.200 476.400 ;
        RECT 178.800 476.300 179.600 476.400 ;
        RECT 124.400 475.700 179.600 476.300 ;
        RECT 124.400 475.600 125.200 475.700 ;
        RECT 178.800 475.600 179.600 475.700 ;
        RECT 316.400 476.300 317.200 476.400 ;
        RECT 354.800 476.300 355.600 476.400 ;
        RECT 316.400 475.700 355.600 476.300 ;
        RECT 316.400 475.600 317.200 475.700 ;
        RECT 354.800 475.600 355.600 475.700 ;
        RECT 364.400 476.300 365.200 476.400 ;
        RECT 382.000 476.300 382.800 476.400 ;
        RECT 385.200 476.300 386.000 476.400 ;
        RECT 364.400 475.700 386.000 476.300 ;
        RECT 364.400 475.600 365.200 475.700 ;
        RECT 382.000 475.600 382.800 475.700 ;
        RECT 385.200 475.600 386.000 475.700 ;
        RECT 391.600 476.300 392.400 476.400 ;
        RECT 393.200 476.300 394.000 476.400 ;
        RECT 391.600 475.700 394.000 476.300 ;
        RECT 391.600 475.600 392.400 475.700 ;
        RECT 393.200 475.600 394.000 475.700 ;
        RECT 409.200 476.300 410.000 476.400 ;
        RECT 434.800 476.300 435.600 476.400 ;
        RECT 409.200 475.700 435.600 476.300 ;
        RECT 409.200 475.600 410.000 475.700 ;
        RECT 434.800 475.600 435.600 475.700 ;
        RECT 438.000 476.300 438.800 476.400 ;
        RECT 447.600 476.300 448.400 476.400 ;
        RECT 438.000 475.700 448.400 476.300 ;
        RECT 438.000 475.600 438.800 475.700 ;
        RECT 447.600 475.600 448.400 475.700 ;
        RECT 449.200 476.300 450.000 476.400 ;
        RECT 486.000 476.300 486.800 476.400 ;
        RECT 487.600 476.300 488.400 476.400 ;
        RECT 449.200 475.700 488.400 476.300 ;
        RECT 449.200 475.600 450.000 475.700 ;
        RECT 486.000 475.600 486.800 475.700 ;
        RECT 487.600 475.600 488.400 475.700 ;
        RECT 545.200 475.600 546.000 476.400 ;
        RECT 18.800 474.300 19.600 474.400 ;
        RECT 26.800 474.300 27.600 474.400 ;
        RECT 71.600 474.300 72.400 474.400 ;
        RECT 114.800 474.300 115.600 474.400 ;
        RECT 18.800 473.700 115.600 474.300 ;
        RECT 18.800 473.600 19.600 473.700 ;
        RECT 26.800 473.600 27.600 473.700 ;
        RECT 71.600 473.600 72.400 473.700 ;
        RECT 114.800 473.600 115.600 473.700 ;
        RECT 119.600 474.300 120.400 474.400 ;
        RECT 127.600 474.300 128.400 474.400 ;
        RECT 119.600 473.700 128.400 474.300 ;
        RECT 119.600 473.600 120.400 473.700 ;
        RECT 127.600 473.600 128.400 473.700 ;
        RECT 135.600 474.300 136.400 474.400 ;
        RECT 289.200 474.300 290.000 474.400 ;
        RECT 292.400 474.300 293.200 474.400 ;
        RECT 135.600 473.700 293.200 474.300 ;
        RECT 135.600 473.600 136.400 473.700 ;
        RECT 289.200 473.600 290.000 473.700 ;
        RECT 292.400 473.600 293.200 473.700 ;
        RECT 327.600 474.300 328.400 474.400 ;
        RECT 354.800 474.300 355.600 474.400 ;
        RECT 361.200 474.300 362.000 474.400 ;
        RECT 327.600 473.700 350.700 474.300 ;
        RECT 327.600 473.600 328.400 473.700 ;
        RECT 350.100 472.400 350.700 473.700 ;
        RECT 354.800 473.700 362.000 474.300 ;
        RECT 354.800 473.600 355.600 473.700 ;
        RECT 361.200 473.600 362.000 473.700 ;
        RECT 367.600 474.300 368.400 474.400 ;
        RECT 402.800 474.300 403.600 474.400 ;
        RECT 414.000 474.300 414.800 474.400 ;
        RECT 431.600 474.300 432.400 474.400 ;
        RECT 441.200 474.300 442.000 474.400 ;
        RECT 367.600 473.700 442.000 474.300 ;
        RECT 367.600 473.600 368.400 473.700 ;
        RECT 402.800 473.600 403.600 473.700 ;
        RECT 414.000 473.600 414.800 473.700 ;
        RECT 431.600 473.600 432.400 473.700 ;
        RECT 441.200 473.600 442.000 473.700 ;
        RECT 446.000 474.300 446.800 474.400 ;
        RECT 468.400 474.300 469.200 474.400 ;
        RECT 446.000 473.700 469.200 474.300 ;
        RECT 446.000 473.600 446.800 473.700 ;
        RECT 468.400 473.600 469.200 473.700 ;
        RECT 478.000 474.300 478.800 474.400 ;
        RECT 481.200 474.300 482.000 474.400 ;
        RECT 478.000 473.700 482.000 474.300 ;
        RECT 478.000 473.600 478.800 473.700 ;
        RECT 481.200 473.600 482.000 473.700 ;
        RECT 518.000 474.300 518.800 474.400 ;
        RECT 554.800 474.300 555.600 474.400 ;
        RECT 518.000 473.700 555.600 474.300 ;
        RECT 518.000 473.600 518.800 473.700 ;
        RECT 554.800 473.600 555.600 473.700 ;
        RECT 39.600 472.300 40.400 472.400 ;
        RECT 58.800 472.300 59.600 472.400 ;
        RECT 39.600 471.700 59.600 472.300 ;
        RECT 39.600 471.600 40.400 471.700 ;
        RECT 58.800 471.600 59.600 471.700 ;
        RECT 94.000 472.300 94.800 472.400 ;
        RECT 111.600 472.300 112.400 472.400 ;
        RECT 154.800 472.300 155.600 472.400 ;
        RECT 94.000 471.700 155.600 472.300 ;
        RECT 94.000 471.600 94.800 471.700 ;
        RECT 111.600 471.600 112.400 471.700 ;
        RECT 154.800 471.600 155.600 471.700 ;
        RECT 169.200 472.300 170.000 472.400 ;
        RECT 185.200 472.300 186.000 472.400 ;
        RECT 169.200 471.700 186.000 472.300 ;
        RECT 169.200 471.600 170.000 471.700 ;
        RECT 185.200 471.600 186.000 471.700 ;
        RECT 210.800 472.300 211.600 472.400 ;
        RECT 223.600 472.300 224.400 472.400 ;
        RECT 210.800 471.700 224.400 472.300 ;
        RECT 210.800 471.600 211.600 471.700 ;
        RECT 223.600 471.600 224.400 471.700 ;
        RECT 238.000 472.300 238.800 472.400 ;
        RECT 250.800 472.300 251.600 472.400 ;
        RECT 257.200 472.300 258.000 472.400 ;
        RECT 287.600 472.300 288.400 472.400 ;
        RECT 238.000 471.700 288.400 472.300 ;
        RECT 238.000 471.600 238.800 471.700 ;
        RECT 250.800 471.600 251.600 471.700 ;
        RECT 257.200 471.600 258.000 471.700 ;
        RECT 287.600 471.600 288.400 471.700 ;
        RECT 329.200 472.300 330.000 472.400 ;
        RECT 330.800 472.300 331.600 472.400 ;
        RECT 329.200 471.700 331.600 472.300 ;
        RECT 329.200 471.600 330.000 471.700 ;
        RECT 330.800 471.600 331.600 471.700 ;
        RECT 350.000 472.300 350.800 472.400 ;
        RECT 364.400 472.300 365.200 472.400 ;
        RECT 350.000 471.700 365.200 472.300 ;
        RECT 350.000 471.600 350.800 471.700 ;
        RECT 364.400 471.600 365.200 471.700 ;
        RECT 372.400 472.300 373.200 472.400 ;
        RECT 404.400 472.300 405.200 472.400 ;
        RECT 372.400 471.700 405.200 472.300 ;
        RECT 372.400 471.600 373.200 471.700 ;
        RECT 404.400 471.600 405.200 471.700 ;
        RECT 410.800 472.300 411.600 472.400 ;
        RECT 442.800 472.300 443.600 472.400 ;
        RECT 465.200 472.300 466.000 472.400 ;
        RECT 468.400 472.300 469.200 472.400 ;
        RECT 481.200 472.300 482.000 472.400 ;
        RECT 410.800 471.700 482.000 472.300 ;
        RECT 410.800 471.600 411.600 471.700 ;
        RECT 442.800 471.600 443.600 471.700 ;
        RECT 465.200 471.600 466.000 471.700 ;
        RECT 468.400 471.600 469.200 471.700 ;
        RECT 481.200 471.600 482.000 471.700 ;
        RECT 486.000 472.300 486.800 472.400 ;
        RECT 497.200 472.300 498.000 472.400 ;
        RECT 486.000 471.700 498.000 472.300 ;
        RECT 486.000 471.600 486.800 471.700 ;
        RECT 497.200 471.600 498.000 471.700 ;
        RECT 503.600 471.600 504.400 472.400 ;
        RECT 508.400 472.300 509.200 472.400 ;
        RECT 529.200 472.300 530.000 472.400 ;
        RECT 553.200 472.300 554.000 472.400 ;
        RECT 508.400 471.700 554.000 472.300 ;
        RECT 508.400 471.600 509.200 471.700 ;
        RECT 529.200 471.600 530.000 471.700 ;
        RECT 553.200 471.600 554.000 471.700 ;
        RECT 7.600 470.300 8.400 470.400 ;
        RECT 23.600 470.300 24.400 470.400 ;
        RECT 7.600 469.700 24.400 470.300 ;
        RECT 7.600 469.600 8.400 469.700 ;
        RECT 23.600 469.600 24.400 469.700 ;
        RECT 30.000 470.300 30.800 470.400 ;
        RECT 54.000 470.300 54.800 470.400 ;
        RECT 30.000 469.700 54.800 470.300 ;
        RECT 30.000 469.600 30.800 469.700 ;
        RECT 54.000 469.600 54.800 469.700 ;
        RECT 73.200 470.300 74.000 470.400 ;
        RECT 103.600 470.300 104.400 470.400 ;
        RECT 73.200 469.700 104.400 470.300 ;
        RECT 73.200 469.600 74.000 469.700 ;
        RECT 103.600 469.600 104.400 469.700 ;
        RECT 113.200 470.300 114.000 470.400 ;
        RECT 126.000 470.300 126.800 470.400 ;
        RECT 113.200 469.700 126.800 470.300 ;
        RECT 113.200 469.600 114.000 469.700 ;
        RECT 126.000 469.600 126.800 469.700 ;
        RECT 127.600 470.300 128.400 470.400 ;
        RECT 130.800 470.300 131.600 470.400 ;
        RECT 127.600 469.700 131.600 470.300 ;
        RECT 127.600 469.600 128.400 469.700 ;
        RECT 130.800 469.600 131.600 469.700 ;
        RECT 135.600 469.600 136.400 470.400 ;
        RECT 166.000 470.300 166.800 470.400 ;
        RECT 172.400 470.300 173.200 470.400 ;
        RECT 166.000 469.700 173.200 470.300 ;
        RECT 166.000 469.600 166.800 469.700 ;
        RECT 172.400 469.600 173.200 469.700 ;
        RECT 174.000 470.300 174.800 470.400 ;
        RECT 177.200 470.300 178.000 470.400 ;
        RECT 174.000 469.700 178.000 470.300 ;
        RECT 174.000 469.600 174.800 469.700 ;
        RECT 177.200 469.600 178.000 469.700 ;
        RECT 204.400 470.300 205.200 470.400 ;
        RECT 218.800 470.300 219.600 470.400 ;
        RECT 204.400 469.700 219.600 470.300 ;
        RECT 204.400 469.600 205.200 469.700 ;
        RECT 218.800 469.600 219.600 469.700 ;
        RECT 241.200 470.300 242.000 470.400 ;
        RECT 254.000 470.300 254.800 470.400 ;
        RECT 241.200 469.700 254.800 470.300 ;
        RECT 241.200 469.600 242.000 469.700 ;
        RECT 254.000 469.600 254.800 469.700 ;
        RECT 330.800 470.300 331.600 470.400 ;
        RECT 356.400 470.300 357.200 470.400 ;
        RECT 330.800 469.700 357.200 470.300 ;
        RECT 330.800 469.600 331.600 469.700 ;
        RECT 356.400 469.600 357.200 469.700 ;
        RECT 359.600 470.300 360.400 470.400 ;
        RECT 374.000 470.300 374.800 470.400 ;
        RECT 359.600 469.700 374.800 470.300 ;
        RECT 359.600 469.600 360.400 469.700 ;
        RECT 374.000 469.600 374.800 469.700 ;
        RECT 378.800 470.300 379.600 470.400 ;
        RECT 439.600 470.300 440.400 470.400 ;
        RECT 444.400 470.300 445.200 470.400 ;
        RECT 482.800 470.300 483.600 470.400 ;
        RECT 519.600 470.300 520.400 470.400 ;
        RECT 530.800 470.300 531.600 470.400 ;
        RECT 378.800 469.700 531.600 470.300 ;
        RECT 378.800 469.600 379.600 469.700 ;
        RECT 439.600 469.600 440.400 469.700 ;
        RECT 444.400 469.600 445.200 469.700 ;
        RECT 482.800 469.600 483.600 469.700 ;
        RECT 519.600 469.600 520.400 469.700 ;
        RECT 530.800 469.600 531.600 469.700 ;
        RECT 554.800 470.300 555.600 470.400 ;
        RECT 577.200 470.300 578.000 470.400 ;
        RECT 554.800 469.700 578.000 470.300 ;
        RECT 554.800 469.600 555.600 469.700 ;
        RECT 577.200 469.600 578.000 469.700 ;
        RECT 31.600 468.300 32.400 468.400 ;
        RECT 41.200 468.300 42.000 468.400 ;
        RECT 52.400 468.300 53.200 468.400 ;
        RECT 31.600 467.700 53.200 468.300 ;
        RECT 31.600 467.600 32.400 467.700 ;
        RECT 41.200 467.600 42.000 467.700 ;
        RECT 52.400 467.600 53.200 467.700 ;
        RECT 57.200 468.300 58.000 468.400 ;
        RECT 81.200 468.300 82.000 468.400 ;
        RECT 57.200 467.700 82.000 468.300 ;
        RECT 57.200 467.600 58.000 467.700 ;
        RECT 81.200 467.600 82.000 467.700 ;
        RECT 94.000 467.600 94.800 468.400 ;
        RECT 103.600 468.300 104.400 468.400 ;
        RECT 148.400 468.300 149.200 468.400 ;
        RECT 103.600 467.700 149.200 468.300 ;
        RECT 103.600 467.600 104.400 467.700 ;
        RECT 148.400 467.600 149.200 467.700 ;
        RECT 162.800 468.300 163.600 468.400 ;
        RECT 170.800 468.300 171.600 468.400 ;
        RECT 172.400 468.300 173.200 468.400 ;
        RECT 162.800 467.700 173.200 468.300 ;
        RECT 162.800 467.600 163.600 467.700 ;
        RECT 170.800 467.600 171.600 467.700 ;
        RECT 172.400 467.600 173.200 467.700 ;
        RECT 177.200 468.300 178.000 468.400 ;
        RECT 196.400 468.300 197.200 468.400 ;
        RECT 177.200 467.700 197.200 468.300 ;
        RECT 177.200 467.600 178.000 467.700 ;
        RECT 196.400 467.600 197.200 467.700 ;
        RECT 212.400 468.300 213.200 468.400 ;
        RECT 222.000 468.300 222.800 468.400 ;
        RECT 212.400 467.700 222.800 468.300 ;
        RECT 212.400 467.600 213.200 467.700 ;
        RECT 222.000 467.600 222.800 467.700 ;
        RECT 234.800 468.300 235.600 468.400 ;
        RECT 242.800 468.300 243.600 468.400 ;
        RECT 234.800 467.700 243.600 468.300 ;
        RECT 234.800 467.600 235.600 467.700 ;
        RECT 242.800 467.600 243.600 467.700 ;
        RECT 327.600 468.300 328.400 468.400 ;
        RECT 332.400 468.300 333.200 468.400 ;
        RECT 327.600 467.700 333.200 468.300 ;
        RECT 327.600 467.600 328.400 467.700 ;
        RECT 332.400 467.600 333.200 467.700 ;
        RECT 345.200 468.300 346.000 468.400 ;
        RECT 388.400 468.300 389.200 468.400 ;
        RECT 399.600 468.300 400.400 468.400 ;
        RECT 345.200 467.700 389.200 468.300 ;
        RECT 345.200 467.600 346.000 467.700 ;
        RECT 388.400 467.600 389.200 467.700 ;
        RECT 396.500 467.700 400.400 468.300 ;
        RECT 62.000 466.300 62.800 466.400 ;
        RECT 79.600 466.300 80.400 466.400 ;
        RECT 62.000 465.700 80.400 466.300 ;
        RECT 81.300 466.300 81.900 467.600 ;
        RECT 111.600 466.300 112.400 466.400 ;
        RECT 81.300 465.700 112.400 466.300 ;
        RECT 62.000 465.600 62.800 465.700 ;
        RECT 79.600 465.600 80.400 465.700 ;
        RECT 111.600 465.600 112.400 465.700 ;
        RECT 127.600 466.300 128.400 466.400 ;
        RECT 134.000 466.300 134.800 466.400 ;
        RECT 127.600 465.700 134.800 466.300 ;
        RECT 127.600 465.600 128.400 465.700 ;
        RECT 134.000 465.600 134.800 465.700 ;
        RECT 153.200 466.300 154.000 466.400 ;
        RECT 180.400 466.300 181.200 466.400 ;
        RECT 153.200 465.700 181.200 466.300 ;
        RECT 153.200 465.600 154.000 465.700 ;
        RECT 180.400 465.600 181.200 465.700 ;
        RECT 183.600 466.300 184.400 466.400 ;
        RECT 228.400 466.300 229.200 466.400 ;
        RECT 183.600 465.700 229.200 466.300 ;
        RECT 183.600 465.600 184.400 465.700 ;
        RECT 228.400 465.600 229.200 465.700 ;
        RECT 241.200 466.300 242.000 466.400 ;
        RECT 246.000 466.300 246.800 466.400 ;
        RECT 241.200 465.700 246.800 466.300 ;
        RECT 241.200 465.600 242.000 465.700 ;
        RECT 246.000 465.600 246.800 465.700 ;
        RECT 252.400 466.300 253.200 466.400 ;
        RECT 270.000 466.300 270.800 466.400 ;
        RECT 252.400 465.700 270.800 466.300 ;
        RECT 252.400 465.600 253.200 465.700 ;
        RECT 270.000 465.600 270.800 465.700 ;
        RECT 364.400 466.300 365.200 466.400 ;
        RECT 396.500 466.300 397.100 467.700 ;
        RECT 399.600 467.600 400.400 467.700 ;
        RECT 426.800 468.300 427.600 468.400 ;
        RECT 431.600 468.300 432.400 468.400 ;
        RECT 426.800 467.700 432.400 468.300 ;
        RECT 426.800 467.600 427.600 467.700 ;
        RECT 431.600 467.600 432.400 467.700 ;
        RECT 438.000 468.300 438.800 468.400 ;
        RECT 446.000 468.300 446.800 468.400 ;
        RECT 438.000 467.700 446.800 468.300 ;
        RECT 438.000 467.600 438.800 467.700 ;
        RECT 446.000 467.600 446.800 467.700 ;
        RECT 465.200 468.300 466.000 468.400 ;
        RECT 468.400 468.300 469.200 468.400 ;
        RECT 465.200 467.700 469.200 468.300 ;
        RECT 465.200 467.600 466.000 467.700 ;
        RECT 468.400 467.600 469.200 467.700 ;
        RECT 494.000 468.300 494.800 468.400 ;
        RECT 500.400 468.300 501.200 468.400 ;
        RECT 494.000 467.700 501.200 468.300 ;
        RECT 494.000 467.600 494.800 467.700 ;
        RECT 500.400 467.600 501.200 467.700 ;
        RECT 502.000 468.300 502.800 468.400 ;
        RECT 526.000 468.300 526.800 468.400 ;
        RECT 502.000 467.700 526.800 468.300 ;
        RECT 502.000 467.600 502.800 467.700 ;
        RECT 526.000 467.600 526.800 467.700 ;
        RECT 548.400 468.300 549.200 468.400 ;
        RECT 567.600 468.300 568.400 468.400 ;
        RECT 548.400 467.700 568.400 468.300 ;
        RECT 548.400 467.600 549.200 467.700 ;
        RECT 567.600 467.600 568.400 467.700 ;
        RECT 578.800 468.300 579.600 468.400 ;
        RECT 599.600 468.300 600.400 468.400 ;
        RECT 578.800 467.700 600.400 468.300 ;
        RECT 578.800 467.600 579.600 467.700 ;
        RECT 599.600 467.600 600.400 467.700 ;
        RECT 364.400 465.700 397.100 466.300 ;
        RECT 398.000 466.300 398.800 466.400 ;
        RECT 404.400 466.300 405.200 466.400 ;
        RECT 398.000 465.700 405.200 466.300 ;
        RECT 364.400 465.600 365.200 465.700 ;
        RECT 398.000 465.600 398.800 465.700 ;
        RECT 404.400 465.600 405.200 465.700 ;
        RECT 420.400 466.300 421.200 466.400 ;
        RECT 438.100 466.300 438.700 467.600 ;
        RECT 420.400 465.700 438.700 466.300 ;
        RECT 471.600 466.300 472.400 466.400 ;
        RECT 506.800 466.300 507.600 466.400 ;
        RECT 471.600 465.700 507.600 466.300 ;
        RECT 420.400 465.600 421.200 465.700 ;
        RECT 471.600 465.600 472.400 465.700 ;
        RECT 506.800 465.600 507.600 465.700 ;
        RECT 519.600 466.300 520.400 466.400 ;
        RECT 556.400 466.300 557.200 466.400 ;
        RECT 519.600 465.700 557.200 466.300 ;
        RECT 519.600 465.600 520.400 465.700 ;
        RECT 556.400 465.600 557.200 465.700 ;
        RECT 583.600 466.300 584.400 466.400 ;
        RECT 588.400 466.300 589.200 466.400 ;
        RECT 583.600 465.700 589.200 466.300 ;
        RECT 583.600 465.600 584.400 465.700 ;
        RECT 588.400 465.600 589.200 465.700 ;
        RECT 22.000 464.300 22.800 464.400 ;
        RECT 68.400 464.300 69.200 464.400 ;
        RECT 22.000 463.700 69.200 464.300 ;
        RECT 22.000 463.600 22.800 463.700 ;
        RECT 68.400 463.600 69.200 463.700 ;
        RECT 118.000 464.300 118.800 464.400 ;
        RECT 143.600 464.300 144.400 464.400 ;
        RECT 166.000 464.300 166.800 464.400 ;
        RECT 118.000 463.700 166.800 464.300 ;
        RECT 118.000 463.600 118.800 463.700 ;
        RECT 143.600 463.600 144.400 463.700 ;
        RECT 166.000 463.600 166.800 463.700 ;
        RECT 207.600 464.300 208.400 464.400 ;
        RECT 214.000 464.300 214.800 464.400 ;
        RECT 207.600 463.700 214.800 464.300 ;
        RECT 207.600 463.600 208.400 463.700 ;
        RECT 214.000 463.600 214.800 463.700 ;
        RECT 230.000 464.300 230.800 464.400 ;
        RECT 244.400 464.300 245.200 464.400 ;
        RECT 247.600 464.300 248.400 464.400 ;
        RECT 230.000 463.700 248.400 464.300 ;
        RECT 230.000 463.600 230.800 463.700 ;
        RECT 244.400 463.600 245.200 463.700 ;
        RECT 247.600 463.600 248.400 463.700 ;
        RECT 278.000 464.300 278.800 464.400 ;
        RECT 286.000 464.300 286.800 464.400 ;
        RECT 303.600 464.300 304.400 464.400 ;
        RECT 278.000 463.700 304.400 464.300 ;
        RECT 278.000 463.600 278.800 463.700 ;
        RECT 286.000 463.600 286.800 463.700 ;
        RECT 303.600 463.600 304.400 463.700 ;
        RECT 335.600 464.300 336.400 464.400 ;
        RECT 340.400 464.300 341.200 464.400 ;
        RECT 335.600 463.700 341.200 464.300 ;
        RECT 335.600 463.600 336.400 463.700 ;
        RECT 340.400 463.600 341.200 463.700 ;
        RECT 348.400 464.300 349.200 464.400 ;
        RECT 393.200 464.300 394.000 464.400 ;
        RECT 414.000 464.300 414.800 464.400 ;
        RECT 348.400 463.700 414.800 464.300 ;
        RECT 348.400 463.600 349.200 463.700 ;
        RECT 393.200 463.600 394.000 463.700 ;
        RECT 414.000 463.600 414.800 463.700 ;
        RECT 460.400 464.300 461.200 464.400 ;
        RECT 478.000 464.300 478.800 464.400 ;
        RECT 460.400 463.700 478.800 464.300 ;
        RECT 460.400 463.600 461.200 463.700 ;
        RECT 478.000 463.600 478.800 463.700 ;
        RECT 63.600 462.300 64.400 462.400 ;
        RECT 81.200 462.300 82.000 462.400 ;
        RECT 106.800 462.300 107.600 462.400 ;
        RECT 63.600 461.700 107.600 462.300 ;
        RECT 63.600 461.600 64.400 461.700 ;
        RECT 81.200 461.600 82.000 461.700 ;
        RECT 106.800 461.600 107.600 461.700 ;
        RECT 116.400 462.300 117.200 462.400 ;
        RECT 140.400 462.300 141.200 462.400 ;
        RECT 167.600 462.300 168.400 462.400 ;
        RECT 116.400 461.700 168.400 462.300 ;
        RECT 116.400 461.600 117.200 461.700 ;
        RECT 140.400 461.600 141.200 461.700 ;
        RECT 167.600 461.600 168.400 461.700 ;
        RECT 340.400 462.300 341.200 462.400 ;
        RECT 353.200 462.300 354.000 462.400 ;
        RECT 340.400 461.700 354.000 462.300 ;
        RECT 340.400 461.600 341.200 461.700 ;
        RECT 353.200 461.600 354.000 461.700 ;
        RECT 396.400 462.300 397.200 462.400 ;
        RECT 398.000 462.300 398.800 462.400 ;
        RECT 396.400 461.700 398.800 462.300 ;
        RECT 396.400 461.600 397.200 461.700 ;
        RECT 398.000 461.600 398.800 461.700 ;
        RECT 410.800 462.300 411.600 462.400 ;
        RECT 415.600 462.300 416.400 462.400 ;
        RECT 410.800 461.700 416.400 462.300 ;
        RECT 410.800 461.600 411.600 461.700 ;
        RECT 415.600 461.600 416.400 461.700 ;
        RECT 430.000 462.300 430.800 462.400 ;
        RECT 434.800 462.300 435.600 462.400 ;
        RECT 430.000 461.700 435.600 462.300 ;
        RECT 430.000 461.600 430.800 461.700 ;
        RECT 434.800 461.600 435.600 461.700 ;
        RECT 441.200 462.300 442.000 462.400 ;
        RECT 471.600 462.300 472.400 462.400 ;
        RECT 441.200 461.700 472.400 462.300 ;
        RECT 441.200 461.600 442.000 461.700 ;
        RECT 471.600 461.600 472.400 461.700 ;
        RECT 38.000 460.300 38.800 460.400 ;
        RECT 100.400 460.300 101.200 460.400 ;
        RECT 38.000 459.700 101.200 460.300 ;
        RECT 38.000 459.600 38.800 459.700 ;
        RECT 100.400 459.600 101.200 459.700 ;
        RECT 135.600 460.300 136.400 460.400 ;
        RECT 138.800 460.300 139.600 460.400 ;
        RECT 143.600 460.300 144.400 460.400 ;
        RECT 177.200 460.300 178.000 460.400 ;
        RECT 183.600 460.300 184.400 460.400 ;
        RECT 135.600 459.700 184.400 460.300 ;
        RECT 135.600 459.600 136.400 459.700 ;
        RECT 138.800 459.600 139.600 459.700 ;
        RECT 143.600 459.600 144.400 459.700 ;
        RECT 177.200 459.600 178.000 459.700 ;
        RECT 183.600 459.600 184.400 459.700 ;
        RECT 185.200 460.300 186.000 460.400 ;
        RECT 196.400 460.300 197.200 460.400 ;
        RECT 185.200 459.700 197.200 460.300 ;
        RECT 185.200 459.600 186.000 459.700 ;
        RECT 196.400 459.600 197.200 459.700 ;
        RECT 246.000 460.300 246.800 460.400 ;
        RECT 250.800 460.300 251.600 460.400 ;
        RECT 246.000 459.700 251.600 460.300 ;
        RECT 246.000 459.600 246.800 459.700 ;
        RECT 250.800 459.600 251.600 459.700 ;
        RECT 318.000 460.300 318.800 460.400 ;
        RECT 375.600 460.300 376.400 460.400 ;
        RECT 396.400 460.300 397.200 460.400 ;
        RECT 486.000 460.300 486.800 460.400 ;
        RECT 318.000 459.700 486.800 460.300 ;
        RECT 318.000 459.600 318.800 459.700 ;
        RECT 375.600 459.600 376.400 459.700 ;
        RECT 396.400 459.600 397.200 459.700 ;
        RECT 486.000 459.600 486.800 459.700 ;
        RECT 516.400 460.300 517.200 460.400 ;
        RECT 521.200 460.300 522.000 460.400 ;
        RECT 551.600 460.300 552.400 460.400 ;
        RECT 516.400 459.700 552.400 460.300 ;
        RECT 516.400 459.600 517.200 459.700 ;
        RECT 521.200 459.600 522.000 459.700 ;
        RECT 551.600 459.600 552.400 459.700 ;
        RECT 562.800 460.300 563.600 460.400 ;
        RECT 583.600 460.300 584.400 460.400 ;
        RECT 562.800 459.700 584.400 460.300 ;
        RECT 562.800 459.600 563.600 459.700 ;
        RECT 583.600 459.600 584.400 459.700 ;
        RECT 591.600 460.300 592.400 460.400 ;
        RECT 596.400 460.300 597.200 460.400 ;
        RECT 591.600 459.700 597.200 460.300 ;
        RECT 591.600 459.600 592.400 459.700 ;
        RECT 596.400 459.600 597.200 459.700 ;
        RECT 46.000 457.600 46.800 458.400 ;
        RECT 89.200 458.300 90.000 458.400 ;
        RECT 95.600 458.300 96.400 458.400 ;
        RECT 89.200 457.700 96.400 458.300 ;
        RECT 89.200 457.600 90.000 457.700 ;
        RECT 95.600 457.600 96.400 457.700 ;
        RECT 146.800 458.300 147.600 458.400 ;
        RECT 159.600 458.300 160.400 458.400 ;
        RECT 207.600 458.300 208.400 458.400 ;
        RECT 146.800 457.700 208.400 458.300 ;
        RECT 146.800 457.600 147.600 457.700 ;
        RECT 159.600 457.600 160.400 457.700 ;
        RECT 207.600 457.600 208.400 457.700 ;
        RECT 372.400 458.300 373.200 458.400 ;
        RECT 377.200 458.300 378.000 458.400 ;
        RECT 460.400 458.300 461.200 458.400 ;
        RECT 372.400 457.700 461.200 458.300 ;
        RECT 372.400 457.600 373.200 457.700 ;
        RECT 377.200 457.600 378.000 457.700 ;
        RECT 460.400 457.600 461.200 457.700 ;
        RECT 505.200 458.300 506.000 458.400 ;
        RECT 514.800 458.300 515.600 458.400 ;
        RECT 535.600 458.300 536.400 458.400 ;
        RECT 540.400 458.300 541.200 458.400 ;
        RECT 505.200 457.700 541.200 458.300 ;
        RECT 505.200 457.600 506.000 457.700 ;
        RECT 514.800 457.600 515.600 457.700 ;
        RECT 535.600 457.600 536.400 457.700 ;
        RECT 540.400 457.600 541.200 457.700 ;
        RECT 543.600 458.300 544.400 458.400 ;
        RECT 559.600 458.300 560.400 458.400 ;
        RECT 543.600 457.700 560.400 458.300 ;
        RECT 543.600 457.600 544.400 457.700 ;
        RECT 559.600 457.600 560.400 457.700 ;
        RECT 17.200 456.300 18.000 456.400 ;
        RECT 54.000 456.300 54.800 456.400 ;
        RECT 17.200 455.700 54.800 456.300 ;
        RECT 17.200 455.600 18.000 455.700 ;
        RECT 54.000 455.600 54.800 455.700 ;
        RECT 105.200 456.300 106.000 456.400 ;
        RECT 140.400 456.300 141.200 456.400 ;
        RECT 105.200 455.700 141.200 456.300 ;
        RECT 105.200 455.600 106.000 455.700 ;
        RECT 140.400 455.600 141.200 455.700 ;
        RECT 167.600 456.300 168.400 456.400 ;
        RECT 175.600 456.300 176.400 456.400 ;
        RECT 198.000 456.300 198.800 456.400 ;
        RECT 167.600 455.700 198.800 456.300 ;
        RECT 167.600 455.600 168.400 455.700 ;
        RECT 175.600 455.600 176.400 455.700 ;
        RECT 198.000 455.600 198.800 455.700 ;
        RECT 274.800 456.300 275.600 456.400 ;
        RECT 281.200 456.300 282.000 456.400 ;
        RECT 274.800 455.700 282.000 456.300 ;
        RECT 274.800 455.600 275.600 455.700 ;
        RECT 281.200 455.600 282.000 455.700 ;
        RECT 286.000 456.300 286.800 456.400 ;
        RECT 295.600 456.300 296.400 456.400 ;
        RECT 286.000 455.700 296.400 456.300 ;
        RECT 286.000 455.600 286.800 455.700 ;
        RECT 295.600 455.600 296.400 455.700 ;
        RECT 342.000 456.300 342.800 456.400 ;
        RECT 350.000 456.300 350.800 456.400 ;
        RECT 342.000 455.700 350.800 456.300 ;
        RECT 342.000 455.600 342.800 455.700 ;
        RECT 350.000 455.600 350.800 455.700 ;
        RECT 364.400 456.300 365.200 456.400 ;
        RECT 410.800 456.300 411.600 456.400 ;
        RECT 364.400 455.700 411.600 456.300 ;
        RECT 364.400 455.600 365.200 455.700 ;
        RECT 410.800 455.600 411.600 455.700 ;
        RECT 412.400 456.300 413.200 456.400 ;
        RECT 455.600 456.300 456.400 456.400 ;
        RECT 412.400 455.700 456.400 456.300 ;
        RECT 412.400 455.600 413.200 455.700 ;
        RECT 455.600 455.600 456.400 455.700 ;
        RECT 476.400 456.300 477.200 456.400 ;
        RECT 481.200 456.300 482.000 456.400 ;
        RECT 476.400 455.700 482.000 456.300 ;
        RECT 476.400 455.600 477.200 455.700 ;
        RECT 481.200 455.600 482.000 455.700 ;
        RECT 484.400 456.300 485.200 456.400 ;
        RECT 506.800 456.300 507.600 456.400 ;
        RECT 484.400 455.700 507.600 456.300 ;
        RECT 484.400 455.600 485.200 455.700 ;
        RECT 506.800 455.600 507.600 455.700 ;
        RECT 556.400 456.300 557.200 456.400 ;
        RECT 591.600 456.300 592.400 456.400 ;
        RECT 556.400 455.700 592.400 456.300 ;
        RECT 556.400 455.600 557.200 455.700 ;
        RECT 591.600 455.600 592.400 455.700 ;
        RECT 22.000 454.300 22.800 454.400 ;
        RECT 26.800 454.300 27.600 454.400 ;
        RECT 22.000 453.700 27.600 454.300 ;
        RECT 22.000 453.600 22.800 453.700 ;
        RECT 26.800 453.600 27.600 453.700 ;
        RECT 33.200 454.300 34.000 454.400 ;
        RECT 36.400 454.300 37.200 454.400 ;
        RECT 33.200 453.700 37.200 454.300 ;
        RECT 33.200 453.600 34.000 453.700 ;
        RECT 36.400 453.600 37.200 453.700 ;
        RECT 42.800 454.300 43.600 454.400 ;
        RECT 50.800 454.300 51.600 454.400 ;
        RECT 52.400 454.300 53.200 454.400 ;
        RECT 78.000 454.300 78.800 454.400 ;
        RECT 42.800 453.700 78.800 454.300 ;
        RECT 42.800 453.600 43.600 453.700 ;
        RECT 50.800 453.600 51.600 453.700 ;
        RECT 52.400 453.600 53.200 453.700 ;
        RECT 78.000 453.600 78.800 453.700 ;
        RECT 79.600 454.300 80.400 454.400 ;
        RECT 82.800 454.300 83.600 454.400 ;
        RECT 79.600 453.700 83.600 454.300 ;
        RECT 79.600 453.600 80.400 453.700 ;
        RECT 82.800 453.600 83.600 453.700 ;
        RECT 86.000 454.300 86.800 454.400 ;
        RECT 121.200 454.300 122.000 454.400 ;
        RECT 86.000 453.700 122.000 454.300 ;
        RECT 86.000 453.600 86.800 453.700 ;
        RECT 121.200 453.600 122.000 453.700 ;
        RECT 126.000 454.300 126.800 454.400 ;
        RECT 145.200 454.300 146.000 454.400 ;
        RECT 177.200 454.300 178.000 454.400 ;
        RECT 185.200 454.300 186.000 454.400 ;
        RECT 126.000 453.700 178.000 454.300 ;
        RECT 126.000 453.600 126.800 453.700 ;
        RECT 145.200 453.600 146.000 453.700 ;
        RECT 177.200 453.600 178.000 453.700 ;
        RECT 178.900 453.700 186.000 454.300 ;
        RECT 14.000 452.300 14.800 452.400 ;
        RECT 23.600 452.300 24.400 452.400 ;
        RECT 14.000 451.700 24.400 452.300 ;
        RECT 14.000 451.600 14.800 451.700 ;
        RECT 23.600 451.600 24.400 451.700 ;
        RECT 28.400 452.300 29.200 452.400 ;
        RECT 79.600 452.300 80.400 452.400 ;
        RECT 28.400 451.700 80.400 452.300 ;
        RECT 28.400 451.600 29.200 451.700 ;
        RECT 79.600 451.600 80.400 451.700 ;
        RECT 100.400 452.300 101.200 452.400 ;
        RECT 103.600 452.300 104.400 452.400 ;
        RECT 100.400 451.700 104.400 452.300 ;
        RECT 100.400 451.600 101.200 451.700 ;
        RECT 103.600 451.600 104.400 451.700 ;
        RECT 108.400 452.300 109.200 452.400 ;
        RECT 114.800 452.300 115.600 452.400 ;
        RECT 108.400 451.700 115.600 452.300 ;
        RECT 108.400 451.600 109.200 451.700 ;
        RECT 114.800 451.600 115.600 451.700 ;
        RECT 148.400 452.300 149.200 452.400 ;
        RECT 162.800 452.300 163.600 452.400 ;
        RECT 169.200 452.300 170.000 452.400 ;
        RECT 148.400 451.700 170.000 452.300 ;
        RECT 148.400 451.600 149.200 451.700 ;
        RECT 162.800 451.600 163.600 451.700 ;
        RECT 169.200 451.600 170.000 451.700 ;
        RECT 175.600 452.300 176.400 452.400 ;
        RECT 178.900 452.300 179.500 453.700 ;
        RECT 185.200 453.600 186.000 453.700 ;
        RECT 193.200 454.300 194.000 454.400 ;
        RECT 222.000 454.300 222.800 454.400 ;
        RECT 193.200 453.700 222.800 454.300 ;
        RECT 193.200 453.600 194.000 453.700 ;
        RECT 222.000 453.600 222.800 453.700 ;
        RECT 228.400 454.300 229.200 454.400 ;
        RECT 236.400 454.300 237.200 454.400 ;
        RECT 228.400 453.700 237.200 454.300 ;
        RECT 228.400 453.600 229.200 453.700 ;
        RECT 236.400 453.600 237.200 453.700 ;
        RECT 239.600 454.300 240.400 454.400 ;
        RECT 276.400 454.300 277.200 454.400 ;
        RECT 282.800 454.300 283.600 454.400 ;
        RECT 286.000 454.300 286.800 454.400 ;
        RECT 239.600 453.700 286.800 454.300 ;
        RECT 239.600 453.600 240.400 453.700 ;
        RECT 276.400 453.600 277.200 453.700 ;
        RECT 282.800 453.600 283.600 453.700 ;
        RECT 286.000 453.600 286.800 453.700 ;
        RECT 292.400 454.300 293.200 454.400 ;
        RECT 316.400 454.300 317.200 454.400 ;
        RECT 292.400 453.700 317.200 454.300 ;
        RECT 292.400 453.600 293.200 453.700 ;
        RECT 316.400 453.600 317.200 453.700 ;
        RECT 361.200 454.300 362.000 454.400 ;
        RECT 369.200 454.300 370.000 454.400 ;
        RECT 361.200 453.700 370.000 454.300 ;
        RECT 361.200 453.600 362.000 453.700 ;
        RECT 369.200 453.600 370.000 453.700 ;
        RECT 382.000 454.300 382.800 454.400 ;
        RECT 386.800 454.300 387.600 454.400 ;
        RECT 382.000 453.700 387.600 454.300 ;
        RECT 382.000 453.600 382.800 453.700 ;
        RECT 386.800 453.600 387.600 453.700 ;
        RECT 390.000 454.300 390.800 454.400 ;
        RECT 399.600 454.300 400.400 454.400 ;
        RECT 390.000 453.700 400.400 454.300 ;
        RECT 390.000 453.600 390.800 453.700 ;
        RECT 399.600 453.600 400.400 453.700 ;
        RECT 415.600 454.300 416.400 454.400 ;
        RECT 422.000 454.300 422.800 454.400 ;
        RECT 415.600 453.700 422.800 454.300 ;
        RECT 415.600 453.600 416.400 453.700 ;
        RECT 422.000 453.600 422.800 453.700 ;
        RECT 428.400 454.300 429.200 454.400 ;
        RECT 439.600 454.300 440.400 454.400 ;
        RECT 428.400 453.700 440.400 454.300 ;
        RECT 428.400 453.600 429.200 453.700 ;
        RECT 439.600 453.600 440.400 453.700 ;
        RECT 468.400 454.300 469.200 454.400 ;
        RECT 470.000 454.300 470.800 454.400 ;
        RECT 468.400 453.700 470.800 454.300 ;
        RECT 468.400 453.600 469.200 453.700 ;
        RECT 470.000 453.600 470.800 453.700 ;
        RECT 474.800 453.600 475.600 454.400 ;
        RECT 479.600 454.300 480.400 454.400 ;
        RECT 486.000 454.300 486.800 454.400 ;
        RECT 479.600 453.700 486.800 454.300 ;
        RECT 479.600 453.600 480.400 453.700 ;
        RECT 486.000 453.600 486.800 453.700 ;
        RECT 494.000 454.300 494.800 454.400 ;
        RECT 498.800 454.300 499.600 454.400 ;
        RECT 494.000 453.700 499.600 454.300 ;
        RECT 494.000 453.600 494.800 453.700 ;
        RECT 498.800 453.600 499.600 453.700 ;
        RECT 505.200 454.300 506.000 454.400 ;
        RECT 572.400 454.300 573.200 454.400 ;
        RECT 505.200 453.700 573.200 454.300 ;
        RECT 505.200 453.600 506.000 453.700 ;
        RECT 572.400 453.600 573.200 453.700 ;
        RECT 175.600 451.700 179.500 452.300 ;
        RECT 180.400 452.300 181.200 452.400 ;
        RECT 188.400 452.300 189.200 452.400 ;
        RECT 180.400 451.700 189.200 452.300 ;
        RECT 175.600 451.600 176.400 451.700 ;
        RECT 180.400 451.600 181.200 451.700 ;
        RECT 188.400 451.600 189.200 451.700 ;
        RECT 198.000 452.300 198.800 452.400 ;
        RECT 202.800 452.300 203.600 452.400 ;
        RECT 198.000 451.700 203.600 452.300 ;
        RECT 198.000 451.600 198.800 451.700 ;
        RECT 202.800 451.600 203.600 451.700 ;
        RECT 257.200 452.300 258.000 452.400 ;
        RECT 273.200 452.300 274.000 452.400 ;
        RECT 257.200 451.700 274.000 452.300 ;
        RECT 257.200 451.600 258.000 451.700 ;
        RECT 273.200 451.600 274.000 451.700 ;
        RECT 343.600 452.300 344.400 452.400 ;
        RECT 362.800 452.300 363.600 452.400 ;
        RECT 343.600 451.700 363.600 452.300 ;
        RECT 343.600 451.600 344.400 451.700 ;
        RECT 362.800 451.600 363.600 451.700 ;
        RECT 367.600 452.300 368.400 452.400 ;
        RECT 410.800 452.300 411.600 452.400 ;
        RECT 367.600 451.700 411.600 452.300 ;
        RECT 367.600 451.600 368.400 451.700 ;
        RECT 410.800 451.600 411.600 451.700 ;
        RECT 414.000 452.300 414.800 452.400 ;
        RECT 420.400 452.300 421.200 452.400 ;
        RECT 414.000 451.700 421.200 452.300 ;
        RECT 414.000 451.600 414.800 451.700 ;
        RECT 420.400 451.600 421.200 451.700 ;
        RECT 444.400 452.300 445.200 452.400 ;
        RECT 450.800 452.300 451.600 452.400 ;
        RECT 444.400 451.700 451.600 452.300 ;
        RECT 444.400 451.600 445.200 451.700 ;
        RECT 450.800 451.600 451.600 451.700 ;
        RECT 474.800 452.300 475.600 452.400 ;
        RECT 484.400 452.300 485.200 452.400 ;
        RECT 474.800 451.700 485.200 452.300 ;
        RECT 474.800 451.600 475.600 451.700 ;
        RECT 484.400 451.600 485.200 451.700 ;
        RECT 492.400 452.300 493.200 452.400 ;
        RECT 500.400 452.300 501.200 452.400 ;
        RECT 492.400 451.700 501.200 452.300 ;
        RECT 492.400 451.600 493.200 451.700 ;
        RECT 500.400 451.600 501.200 451.700 ;
        RECT 508.400 452.300 509.200 452.400 ;
        RECT 513.200 452.300 514.000 452.400 ;
        RECT 508.400 451.700 514.000 452.300 ;
        RECT 508.400 451.600 509.200 451.700 ;
        RECT 513.200 451.600 514.000 451.700 ;
        RECT 514.800 452.300 515.600 452.400 ;
        RECT 516.400 452.300 517.200 452.400 ;
        RECT 514.800 451.700 517.200 452.300 ;
        RECT 514.800 451.600 515.600 451.700 ;
        RECT 516.400 451.600 517.200 451.700 ;
        RECT 518.000 452.300 518.800 452.400 ;
        RECT 530.800 452.300 531.600 452.400 ;
        RECT 518.000 451.700 531.600 452.300 ;
        RECT 518.000 451.600 518.800 451.700 ;
        RECT 530.800 451.600 531.600 451.700 ;
        RECT 542.000 452.300 542.800 452.400 ;
        RECT 559.600 452.300 560.400 452.400 ;
        RECT 542.000 451.700 560.400 452.300 ;
        RECT 542.000 451.600 542.800 451.700 ;
        RECT 559.600 451.600 560.400 451.700 ;
        RECT 590.000 452.300 590.800 452.400 ;
        RECT 593.200 452.300 594.000 452.400 ;
        RECT 590.000 451.700 594.000 452.300 ;
        RECT 590.000 451.600 590.800 451.700 ;
        RECT 593.200 451.600 594.000 451.700 ;
        RECT 25.200 450.300 26.000 450.400 ;
        RECT 28.400 450.300 29.200 450.400 ;
        RECT 25.200 449.700 29.200 450.300 ;
        RECT 25.200 449.600 26.000 449.700 ;
        RECT 28.400 449.600 29.200 449.700 ;
        RECT 58.800 450.300 59.600 450.400 ;
        RECT 82.800 450.300 83.600 450.400 ;
        RECT 58.800 449.700 83.600 450.300 ;
        RECT 58.800 449.600 59.600 449.700 ;
        RECT 82.800 449.600 83.600 449.700 ;
        RECT 102.000 450.300 102.800 450.400 ;
        RECT 113.200 450.300 114.000 450.400 ;
        RECT 102.000 449.700 114.000 450.300 ;
        RECT 102.000 449.600 102.800 449.700 ;
        RECT 113.200 449.600 114.000 449.700 ;
        RECT 114.800 450.300 115.600 450.400 ;
        RECT 138.800 450.300 139.600 450.400 ;
        RECT 114.800 449.700 139.600 450.300 ;
        RECT 114.800 449.600 115.600 449.700 ;
        RECT 138.800 449.600 139.600 449.700 ;
        RECT 142.000 450.300 142.800 450.400 ;
        RECT 148.400 450.300 149.200 450.400 ;
        RECT 142.000 449.700 149.200 450.300 ;
        RECT 142.000 449.600 142.800 449.700 ;
        RECT 148.400 449.600 149.200 449.700 ;
        RECT 161.200 450.300 162.000 450.400 ;
        RECT 162.800 450.300 163.600 450.400 ;
        RECT 169.200 450.300 170.000 450.400 ;
        RECT 183.600 450.300 184.400 450.400 ;
        RECT 161.200 449.700 184.400 450.300 ;
        RECT 161.200 449.600 162.000 449.700 ;
        RECT 162.800 449.600 163.600 449.700 ;
        RECT 169.200 449.600 170.000 449.700 ;
        RECT 183.600 449.600 184.400 449.700 ;
        RECT 190.000 450.300 190.800 450.400 ;
        RECT 210.800 450.300 211.600 450.400 ;
        RECT 276.400 450.300 277.200 450.400 ;
        RECT 190.000 449.700 277.200 450.300 ;
        RECT 190.000 449.600 190.800 449.700 ;
        RECT 210.800 449.600 211.600 449.700 ;
        RECT 276.400 449.600 277.200 449.700 ;
        RECT 330.800 450.300 331.600 450.400 ;
        RECT 367.600 450.300 368.400 450.400 ;
        RECT 330.800 449.700 368.400 450.300 ;
        RECT 330.800 449.600 331.600 449.700 ;
        RECT 367.600 449.600 368.400 449.700 ;
        RECT 382.000 450.300 382.800 450.400 ;
        RECT 390.000 450.300 390.800 450.400 ;
        RECT 382.000 449.700 390.800 450.300 ;
        RECT 382.000 449.600 382.800 449.700 ;
        RECT 390.000 449.600 390.800 449.700 ;
        RECT 401.200 450.300 402.000 450.400 ;
        RECT 430.000 450.300 430.800 450.400 ;
        RECT 401.200 449.700 430.800 450.300 ;
        RECT 401.200 449.600 402.000 449.700 ;
        RECT 430.000 449.600 430.800 449.700 ;
        RECT 471.600 450.300 472.400 450.400 ;
        RECT 492.400 450.300 493.200 450.400 ;
        RECT 471.600 449.700 493.200 450.300 ;
        RECT 471.600 449.600 472.400 449.700 ;
        RECT 492.400 449.600 493.200 449.700 ;
        RECT 503.600 450.300 504.400 450.400 ;
        RECT 526.000 450.300 526.800 450.400 ;
        RECT 503.600 449.700 526.800 450.300 ;
        RECT 503.600 449.600 504.400 449.700 ;
        RECT 526.000 449.600 526.800 449.700 ;
        RECT 559.600 450.300 560.400 450.400 ;
        RECT 594.800 450.300 595.600 450.400 ;
        RECT 559.600 449.700 595.600 450.300 ;
        RECT 559.600 449.600 560.400 449.700 ;
        RECT 594.800 449.600 595.600 449.700 ;
        RECT 9.200 448.300 10.000 448.400 ;
        RECT 26.800 448.300 27.600 448.400 ;
        RECT 9.200 447.700 27.600 448.300 ;
        RECT 9.200 447.600 10.000 447.700 ;
        RECT 26.800 447.600 27.600 447.700 ;
        RECT 46.000 448.300 46.800 448.400 ;
        RECT 49.200 448.300 50.000 448.400 ;
        RECT 46.000 447.700 50.000 448.300 ;
        RECT 46.000 447.600 46.800 447.700 ;
        RECT 49.200 447.600 50.000 447.700 ;
        RECT 70.000 448.300 70.800 448.400 ;
        RECT 73.200 448.300 74.000 448.400 ;
        RECT 87.600 448.300 88.400 448.400 ;
        RECT 106.800 448.300 107.600 448.400 ;
        RECT 70.000 447.700 107.600 448.300 ;
        RECT 70.000 447.600 70.800 447.700 ;
        RECT 73.200 447.600 74.000 447.700 ;
        RECT 87.600 447.600 88.400 447.700 ;
        RECT 106.800 447.600 107.600 447.700 ;
        RECT 110.000 448.300 110.800 448.400 ;
        RECT 116.400 448.300 117.200 448.400 ;
        RECT 110.000 447.700 117.200 448.300 ;
        RECT 110.000 447.600 110.800 447.700 ;
        RECT 116.400 447.600 117.200 447.700 ;
        RECT 166.000 448.300 166.800 448.400 ;
        RECT 199.600 448.300 200.400 448.400 ;
        RECT 209.200 448.300 210.000 448.400 ;
        RECT 166.000 447.700 210.000 448.300 ;
        RECT 166.000 447.600 166.800 447.700 ;
        RECT 199.600 447.600 200.400 447.700 ;
        RECT 209.200 447.600 210.000 447.700 ;
        RECT 246.000 448.300 246.800 448.400 ;
        RECT 265.200 448.300 266.000 448.400 ;
        RECT 246.000 447.700 266.000 448.300 ;
        RECT 246.000 447.600 246.800 447.700 ;
        RECT 265.200 447.600 266.000 447.700 ;
        RECT 351.600 448.300 352.400 448.400 ;
        RECT 436.400 448.300 437.200 448.400 ;
        RECT 351.600 447.700 437.200 448.300 ;
        RECT 351.600 447.600 352.400 447.700 ;
        RECT 436.400 447.600 437.200 447.700 ;
        RECT 446.000 448.300 446.800 448.400 ;
        RECT 452.400 448.300 453.200 448.400 ;
        RECT 446.000 447.700 453.200 448.300 ;
        RECT 446.000 447.600 446.800 447.700 ;
        RECT 452.400 447.600 453.200 447.700 ;
        RECT 505.200 448.300 506.000 448.400 ;
        RECT 511.600 448.300 512.400 448.400 ;
        RECT 505.200 447.700 512.400 448.300 ;
        RECT 505.200 447.600 506.000 447.700 ;
        RECT 511.600 447.600 512.400 447.700 ;
        RECT 513.200 448.300 514.000 448.400 ;
        RECT 516.400 448.300 517.200 448.400 ;
        RECT 513.200 447.700 517.200 448.300 ;
        RECT 513.200 447.600 514.000 447.700 ;
        RECT 516.400 447.600 517.200 447.700 ;
        RECT 78.000 446.300 78.800 446.400 ;
        RECT 94.000 446.300 94.800 446.400 ;
        RECT 78.000 445.700 94.800 446.300 ;
        RECT 78.000 445.600 78.800 445.700 ;
        RECT 94.000 445.600 94.800 445.700 ;
        RECT 132.400 446.300 133.200 446.400 ;
        RECT 137.200 446.300 138.000 446.400 ;
        RECT 164.400 446.300 165.200 446.400 ;
        RECT 132.400 445.700 165.200 446.300 ;
        RECT 132.400 445.600 133.200 445.700 ;
        RECT 137.200 445.600 138.000 445.700 ;
        RECT 164.400 445.600 165.200 445.700 ;
        RECT 297.200 446.300 298.000 446.400 ;
        RECT 298.800 446.300 299.600 446.400 ;
        RECT 297.200 445.700 299.600 446.300 ;
        RECT 297.200 445.600 298.000 445.700 ;
        RECT 298.800 445.600 299.600 445.700 ;
        RECT 431.600 446.300 432.400 446.400 ;
        RECT 454.000 446.300 454.800 446.400 ;
        RECT 463.600 446.300 464.400 446.400 ;
        RECT 510.000 446.300 510.800 446.400 ;
        RECT 431.600 445.700 510.800 446.300 ;
        RECT 431.600 445.600 432.400 445.700 ;
        RECT 454.000 445.600 454.800 445.700 ;
        RECT 463.600 445.600 464.400 445.700 ;
        RECT 510.000 445.600 510.800 445.700 ;
        RECT 44.400 444.300 45.200 444.400 ;
        RECT 98.800 444.300 99.600 444.400 ;
        RECT 44.400 443.700 99.600 444.300 ;
        RECT 44.400 443.600 45.200 443.700 ;
        RECT 98.800 443.600 99.600 443.700 ;
        RECT 154.800 444.300 155.600 444.400 ;
        RECT 161.200 444.300 162.000 444.400 ;
        RECT 154.800 443.700 162.000 444.300 ;
        RECT 154.800 443.600 155.600 443.700 ;
        RECT 161.200 443.600 162.000 443.700 ;
        RECT 233.200 444.300 234.000 444.400 ;
        RECT 295.600 444.300 296.400 444.400 ;
        RECT 305.200 444.300 306.000 444.400 ;
        RECT 233.200 443.700 306.000 444.300 ;
        RECT 233.200 443.600 234.000 443.700 ;
        RECT 295.600 443.600 296.400 443.700 ;
        RECT 305.200 443.600 306.000 443.700 ;
        RECT 348.400 444.300 349.200 444.400 ;
        RECT 375.600 444.300 376.400 444.400 ;
        RECT 348.400 443.700 376.400 444.300 ;
        RECT 348.400 443.600 349.200 443.700 ;
        RECT 375.600 443.600 376.400 443.700 ;
        RECT 385.200 444.300 386.000 444.400 ;
        RECT 409.200 444.300 410.000 444.400 ;
        RECT 434.800 444.300 435.600 444.400 ;
        RECT 385.200 443.700 435.600 444.300 ;
        RECT 385.200 443.600 386.000 443.700 ;
        RECT 409.200 443.600 410.000 443.700 ;
        RECT 434.800 443.600 435.600 443.700 ;
        RECT 441.200 444.300 442.000 444.400 ;
        RECT 450.800 444.300 451.600 444.400 ;
        RECT 441.200 443.700 451.600 444.300 ;
        RECT 441.200 443.600 442.000 443.700 ;
        RECT 450.800 443.600 451.600 443.700 ;
        RECT 495.600 444.300 496.400 444.400 ;
        RECT 519.600 444.300 520.400 444.400 ;
        RECT 495.600 443.700 520.400 444.300 ;
        RECT 495.600 443.600 496.400 443.700 ;
        RECT 519.600 443.600 520.400 443.700 ;
        RECT 87.600 442.300 88.400 442.400 ;
        RECT 116.400 442.300 117.200 442.400 ;
        RECT 87.600 441.700 117.200 442.300 ;
        RECT 87.600 441.600 88.400 441.700 ;
        RECT 116.400 441.600 117.200 441.700 ;
        RECT 134.000 442.300 134.800 442.400 ;
        RECT 135.600 442.300 136.400 442.400 ;
        RECT 134.000 441.700 136.400 442.300 ;
        RECT 134.000 441.600 134.800 441.700 ;
        RECT 135.600 441.600 136.400 441.700 ;
        RECT 249.200 442.300 250.000 442.400 ;
        RECT 250.800 442.300 251.600 442.400 ;
        RECT 249.200 441.700 251.600 442.300 ;
        RECT 249.200 441.600 250.000 441.700 ;
        RECT 250.800 441.600 251.600 441.700 ;
        RECT 522.800 442.300 523.600 442.400 ;
        RECT 566.000 442.300 566.800 442.400 ;
        RECT 522.800 441.700 566.800 442.300 ;
        RECT 522.800 441.600 523.600 441.700 ;
        RECT 566.000 441.600 566.800 441.700 ;
        RECT 574.000 442.300 574.800 442.400 ;
        RECT 580.400 442.300 581.200 442.400 ;
        RECT 574.000 441.700 581.200 442.300 ;
        RECT 574.000 441.600 574.800 441.700 ;
        RECT 580.400 441.600 581.200 441.700 ;
        RECT 599.600 442.300 600.400 442.400 ;
        RECT 606.000 442.300 606.800 442.400 ;
        RECT 599.600 441.700 606.800 442.300 ;
        RECT 599.600 441.600 600.400 441.700 ;
        RECT 606.000 441.600 606.800 441.700 ;
        RECT 12.400 440.300 13.200 440.400 ;
        RECT 22.000 440.300 22.800 440.400 ;
        RECT 12.400 439.700 22.800 440.300 ;
        RECT 12.400 439.600 13.200 439.700 ;
        RECT 22.000 439.600 22.800 439.700 ;
        RECT 129.200 440.300 130.000 440.400 ;
        RECT 134.000 440.300 134.800 440.400 ;
        RECT 129.200 439.700 134.800 440.300 ;
        RECT 129.200 439.600 130.000 439.700 ;
        RECT 134.000 439.600 134.800 439.700 ;
        RECT 295.600 440.300 296.400 440.400 ;
        RECT 297.200 440.300 298.000 440.400 ;
        RECT 295.600 439.700 298.000 440.300 ;
        RECT 295.600 439.600 296.400 439.700 ;
        RECT 297.200 439.600 298.000 439.700 ;
        RECT 535.600 440.300 536.400 440.400 ;
        RECT 545.200 440.300 546.000 440.400 ;
        RECT 548.400 440.300 549.200 440.400 ;
        RECT 535.600 439.700 549.200 440.300 ;
        RECT 535.600 439.600 536.400 439.700 ;
        RECT 545.200 439.600 546.000 439.700 ;
        RECT 548.400 439.600 549.200 439.700 ;
        RECT 551.600 440.300 552.400 440.400 ;
        RECT 575.600 440.300 576.400 440.400 ;
        RECT 551.600 439.700 576.400 440.300 ;
        RECT 551.600 439.600 552.400 439.700 ;
        RECT 575.600 439.600 576.400 439.700 ;
        RECT 167.600 437.600 168.400 438.400 ;
        RECT 214.000 438.300 214.800 438.400 ;
        RECT 242.800 438.300 243.600 438.400 ;
        RECT 214.000 437.700 243.600 438.300 ;
        RECT 214.000 437.600 214.800 437.700 ;
        RECT 242.800 437.600 243.600 437.700 ;
        RECT 266.800 438.300 267.600 438.400 ;
        RECT 278.000 438.300 278.800 438.400 ;
        RECT 266.800 437.700 278.800 438.300 ;
        RECT 266.800 437.600 267.600 437.700 ;
        RECT 278.000 437.600 278.800 437.700 ;
        RECT 350.000 438.300 350.800 438.400 ;
        RECT 356.400 438.300 357.200 438.400 ;
        RECT 372.400 438.300 373.200 438.400 ;
        RECT 350.000 437.700 373.200 438.300 ;
        RECT 350.000 437.600 350.800 437.700 ;
        RECT 356.400 437.600 357.200 437.700 ;
        RECT 372.400 437.600 373.200 437.700 ;
        RECT 414.000 438.300 414.800 438.400 ;
        RECT 420.400 438.300 421.200 438.400 ;
        RECT 414.000 437.700 421.200 438.300 ;
        RECT 414.000 437.600 414.800 437.700 ;
        RECT 420.400 437.600 421.200 437.700 ;
        RECT 454.000 438.300 454.800 438.400 ;
        RECT 476.400 438.300 477.200 438.400 ;
        RECT 454.000 437.700 477.200 438.300 ;
        RECT 454.000 437.600 454.800 437.700 ;
        RECT 476.400 437.600 477.200 437.700 ;
        RECT 506.800 438.300 507.600 438.400 ;
        RECT 511.600 438.300 512.400 438.400 ;
        RECT 506.800 437.700 512.400 438.300 ;
        RECT 506.800 437.600 507.600 437.700 ;
        RECT 511.600 437.600 512.400 437.700 ;
        RECT 529.200 438.300 530.000 438.400 ;
        RECT 535.600 438.300 536.400 438.400 ;
        RECT 529.200 437.700 536.400 438.300 ;
        RECT 529.200 437.600 530.000 437.700 ;
        RECT 535.600 437.600 536.400 437.700 ;
        RECT 17.200 436.300 18.000 436.400 ;
        RECT 49.200 436.300 50.000 436.400 ;
        RECT 71.600 436.300 72.400 436.400 ;
        RECT 127.600 436.300 128.400 436.400 ;
        RECT 137.200 436.300 138.000 436.400 ;
        RECT 17.200 435.700 138.000 436.300 ;
        RECT 17.200 435.600 18.000 435.700 ;
        RECT 49.200 435.600 50.000 435.700 ;
        RECT 71.600 435.600 72.400 435.700 ;
        RECT 127.600 435.600 128.400 435.700 ;
        RECT 137.200 435.600 138.000 435.700 ;
        RECT 140.400 436.300 141.200 436.400 ;
        RECT 225.200 436.300 226.000 436.400 ;
        RECT 278.000 436.300 278.800 436.400 ;
        RECT 140.400 435.700 278.800 436.300 ;
        RECT 140.400 435.600 141.200 435.700 ;
        RECT 225.200 435.600 226.000 435.700 ;
        RECT 278.000 435.600 278.800 435.700 ;
        RECT 346.800 436.300 347.600 436.400 ;
        RECT 356.400 436.300 357.200 436.400 ;
        RECT 367.600 436.300 368.400 436.400 ;
        RECT 382.000 436.300 382.800 436.400 ;
        RECT 346.800 435.700 382.800 436.300 ;
        RECT 346.800 435.600 347.600 435.700 ;
        RECT 356.400 435.600 357.200 435.700 ;
        RECT 367.600 435.600 368.400 435.700 ;
        RECT 382.000 435.600 382.800 435.700 ;
        RECT 452.400 436.300 453.200 436.400 ;
        RECT 470.000 436.300 470.800 436.400 ;
        RECT 505.200 436.300 506.000 436.400 ;
        RECT 452.400 435.700 506.000 436.300 ;
        RECT 452.400 435.600 453.200 435.700 ;
        RECT 470.000 435.600 470.800 435.700 ;
        RECT 505.200 435.600 506.000 435.700 ;
        RECT 70.000 434.300 70.800 434.400 ;
        RECT 73.200 434.300 74.000 434.400 ;
        RECT 70.000 433.700 74.000 434.300 ;
        RECT 70.000 433.600 70.800 433.700 ;
        RECT 73.200 433.600 74.000 433.700 ;
        RECT 81.200 434.300 82.000 434.400 ;
        RECT 108.400 434.300 109.200 434.400 ;
        RECT 81.200 433.700 109.200 434.300 ;
        RECT 81.200 433.600 82.000 433.700 ;
        RECT 108.400 433.600 109.200 433.700 ;
        RECT 118.000 434.300 118.800 434.400 ;
        RECT 129.200 434.300 130.000 434.400 ;
        RECT 118.000 433.700 130.000 434.300 ;
        RECT 118.000 433.600 118.800 433.700 ;
        RECT 129.200 433.600 130.000 433.700 ;
        RECT 167.600 434.300 168.400 434.400 ;
        RECT 194.800 434.300 195.600 434.400 ;
        RECT 167.600 433.700 195.600 434.300 ;
        RECT 167.600 433.600 168.400 433.700 ;
        RECT 194.800 433.600 195.600 433.700 ;
        RECT 201.200 434.300 202.000 434.400 ;
        RECT 207.600 434.300 208.400 434.400 ;
        RECT 201.200 433.700 208.400 434.300 ;
        RECT 201.200 433.600 202.000 433.700 ;
        RECT 207.600 433.600 208.400 433.700 ;
        RECT 212.400 434.300 213.200 434.400 ;
        RECT 220.400 434.300 221.200 434.400 ;
        RECT 268.400 434.300 269.200 434.400 ;
        RECT 271.600 434.300 272.400 434.400 ;
        RECT 212.400 433.700 272.400 434.300 ;
        RECT 212.400 433.600 213.200 433.700 ;
        RECT 220.400 433.600 221.200 433.700 ;
        RECT 268.400 433.600 269.200 433.700 ;
        RECT 271.600 433.600 272.400 433.700 ;
        RECT 406.000 434.300 406.800 434.400 ;
        RECT 412.400 434.300 413.200 434.400 ;
        RECT 415.600 434.300 416.400 434.400 ;
        RECT 406.000 433.700 416.400 434.300 ;
        RECT 406.000 433.600 406.800 433.700 ;
        RECT 412.400 433.600 413.200 433.700 ;
        RECT 415.600 433.600 416.400 433.700 ;
        RECT 462.000 434.300 462.800 434.400 ;
        RECT 474.800 434.300 475.600 434.400 ;
        RECT 462.000 433.700 475.600 434.300 ;
        RECT 462.000 433.600 462.800 433.700 ;
        RECT 474.800 433.600 475.600 433.700 ;
        RECT 1.200 432.300 2.000 432.400 ;
        RECT 25.200 432.300 26.000 432.400 ;
        RECT 33.200 432.300 34.000 432.400 ;
        RECT 1.200 431.700 34.000 432.300 ;
        RECT 1.200 431.600 2.000 431.700 ;
        RECT 25.200 431.600 26.000 431.700 ;
        RECT 33.200 431.600 34.000 431.700 ;
        RECT 73.200 432.300 74.000 432.400 ;
        RECT 87.600 432.300 88.400 432.400 ;
        RECT 94.000 432.300 94.800 432.400 ;
        RECT 73.200 431.700 94.800 432.300 ;
        RECT 73.200 431.600 74.000 431.700 ;
        RECT 87.600 431.600 88.400 431.700 ;
        RECT 94.000 431.600 94.800 431.700 ;
        RECT 113.200 432.300 114.000 432.400 ;
        RECT 145.200 432.300 146.000 432.400 ;
        RECT 113.200 431.700 146.000 432.300 ;
        RECT 113.200 431.600 114.000 431.700 ;
        RECT 145.200 431.600 146.000 431.700 ;
        RECT 146.800 432.300 147.600 432.400 ;
        RECT 156.400 432.300 157.200 432.400 ;
        RECT 146.800 431.700 157.200 432.300 ;
        RECT 146.800 431.600 147.600 431.700 ;
        RECT 156.400 431.600 157.200 431.700 ;
        RECT 158.000 432.300 158.800 432.400 ;
        RECT 167.600 432.300 168.400 432.400 ;
        RECT 158.000 431.700 168.400 432.300 ;
        RECT 158.000 431.600 158.800 431.700 ;
        RECT 167.600 431.600 168.400 431.700 ;
        RECT 215.600 432.300 216.400 432.400 ;
        RECT 218.800 432.300 219.600 432.400 ;
        RECT 215.600 431.700 219.600 432.300 ;
        RECT 215.600 431.600 216.400 431.700 ;
        RECT 218.800 431.600 219.600 431.700 ;
        RECT 222.000 432.300 222.800 432.400 ;
        RECT 230.000 432.300 230.800 432.400 ;
        RECT 222.000 431.700 230.800 432.300 ;
        RECT 222.000 431.600 222.800 431.700 ;
        RECT 230.000 431.600 230.800 431.700 ;
        RECT 241.200 432.300 242.000 432.400 ;
        RECT 255.600 432.300 256.400 432.400 ;
        RECT 276.400 432.300 277.200 432.400 ;
        RECT 287.600 432.300 288.400 432.400 ;
        RECT 241.200 431.700 288.400 432.300 ;
        RECT 241.200 431.600 242.000 431.700 ;
        RECT 255.600 431.600 256.400 431.700 ;
        RECT 276.400 431.600 277.200 431.700 ;
        RECT 287.600 431.600 288.400 431.700 ;
        RECT 346.800 432.300 347.600 432.400 ;
        RECT 354.800 432.300 355.600 432.400 ;
        RECT 364.400 432.300 365.200 432.400 ;
        RECT 346.800 431.700 365.200 432.300 ;
        RECT 346.800 431.600 347.600 431.700 ;
        RECT 354.800 431.600 355.600 431.700 ;
        RECT 364.400 431.600 365.200 431.700 ;
        RECT 398.000 432.300 398.800 432.400 ;
        RECT 494.000 432.300 494.800 432.400 ;
        RECT 398.000 431.700 494.800 432.300 ;
        RECT 398.000 431.600 398.800 431.700 ;
        RECT 494.000 431.600 494.800 431.700 ;
        RECT 2.800 430.300 3.600 430.400 ;
        RECT 6.000 430.300 6.800 430.400 ;
        RECT 36.400 430.300 37.200 430.400 ;
        RECT 2.800 429.700 37.200 430.300 ;
        RECT 2.800 429.600 3.600 429.700 ;
        RECT 6.000 429.600 6.800 429.700 ;
        RECT 36.400 429.600 37.200 429.700 ;
        RECT 44.400 430.300 45.200 430.400 ;
        RECT 58.800 430.300 59.600 430.400 ;
        RECT 44.400 429.700 59.600 430.300 ;
        RECT 44.400 429.600 45.200 429.700 ;
        RECT 58.800 429.600 59.600 429.700 ;
        RECT 60.400 430.300 61.200 430.400 ;
        RECT 84.400 430.300 85.200 430.400 ;
        RECT 60.400 429.700 85.200 430.300 ;
        RECT 60.400 429.600 61.200 429.700 ;
        RECT 84.400 429.600 85.200 429.700 ;
        RECT 89.200 430.300 90.000 430.400 ;
        RECT 98.800 430.300 99.600 430.400 ;
        RECT 89.200 429.700 99.600 430.300 ;
        RECT 89.200 429.600 90.000 429.700 ;
        RECT 98.800 429.600 99.600 429.700 ;
        RECT 106.800 430.300 107.600 430.400 ;
        RECT 114.800 430.300 115.600 430.400 ;
        RECT 134.000 430.300 134.800 430.400 ;
        RECT 106.800 429.700 134.800 430.300 ;
        RECT 106.800 429.600 107.600 429.700 ;
        RECT 114.800 429.600 115.600 429.700 ;
        RECT 134.000 429.600 134.800 429.700 ;
        RECT 156.400 430.300 157.200 430.400 ;
        RECT 172.400 430.300 173.200 430.400 ;
        RECT 156.400 429.700 173.200 430.300 ;
        RECT 156.400 429.600 157.200 429.700 ;
        RECT 172.400 429.600 173.200 429.700 ;
        RECT 196.400 430.300 197.200 430.400 ;
        RECT 210.800 430.300 211.600 430.400 ;
        RECT 196.400 429.700 211.600 430.300 ;
        RECT 196.400 429.600 197.200 429.700 ;
        RECT 210.800 429.600 211.600 429.700 ;
        RECT 223.600 430.300 224.400 430.400 ;
        RECT 226.800 430.300 227.600 430.400 ;
        RECT 242.800 430.300 243.600 430.400 ;
        RECT 223.600 429.700 227.600 430.300 ;
        RECT 223.600 429.600 224.400 429.700 ;
        RECT 226.800 429.600 227.600 429.700 ;
        RECT 228.500 429.700 243.600 430.300 ;
        RECT 10.800 428.300 11.600 428.400 ;
        RECT 14.000 428.300 14.800 428.400 ;
        RECT 10.800 427.700 14.800 428.300 ;
        RECT 10.800 427.600 11.600 427.700 ;
        RECT 14.000 427.600 14.800 427.700 ;
        RECT 33.200 428.300 34.000 428.400 ;
        RECT 36.400 428.300 37.200 428.400 ;
        RECT 39.600 428.300 40.400 428.400 ;
        RECT 33.200 427.700 40.400 428.300 ;
        RECT 33.200 427.600 34.000 427.700 ;
        RECT 36.400 427.600 37.200 427.700 ;
        RECT 39.600 427.600 40.400 427.700 ;
        RECT 50.800 428.300 51.600 428.400 ;
        RECT 54.000 428.300 54.800 428.400 ;
        RECT 50.800 427.700 54.800 428.300 ;
        RECT 50.800 427.600 51.600 427.700 ;
        RECT 54.000 427.600 54.800 427.700 ;
        RECT 63.600 428.300 64.400 428.400 ;
        RECT 100.400 428.300 101.200 428.400 ;
        RECT 63.600 427.700 101.200 428.300 ;
        RECT 63.600 427.600 64.400 427.700 ;
        RECT 100.400 427.600 101.200 427.700 ;
        RECT 106.800 428.300 107.600 428.400 ;
        RECT 110.000 428.300 110.800 428.400 ;
        RECT 106.800 427.700 110.800 428.300 ;
        RECT 106.800 427.600 107.600 427.700 ;
        RECT 110.000 427.600 110.800 427.700 ;
        RECT 124.400 428.300 125.200 428.400 ;
        RECT 156.400 428.300 157.200 428.400 ;
        RECT 124.400 427.700 157.200 428.300 ;
        RECT 124.400 427.600 125.200 427.700 ;
        RECT 156.400 427.600 157.200 427.700 ;
        RECT 158.000 428.300 158.800 428.400 ;
        RECT 170.800 428.300 171.600 428.400 ;
        RECT 158.000 427.700 171.600 428.300 ;
        RECT 158.000 427.600 158.800 427.700 ;
        RECT 170.800 427.600 171.600 427.700 ;
        RECT 202.800 427.600 203.600 428.400 ;
        RECT 218.800 428.300 219.600 428.400 ;
        RECT 228.500 428.300 229.100 429.700 ;
        RECT 242.800 429.600 243.600 429.700 ;
        RECT 254.000 430.300 254.800 430.400 ;
        RECT 260.400 430.300 261.200 430.400 ;
        RECT 254.000 429.700 261.200 430.300 ;
        RECT 254.000 429.600 254.800 429.700 ;
        RECT 260.400 429.600 261.200 429.700 ;
        RECT 265.200 430.300 266.000 430.400 ;
        RECT 274.800 430.300 275.600 430.400 ;
        RECT 265.200 429.700 275.600 430.300 ;
        RECT 265.200 429.600 266.000 429.700 ;
        RECT 274.800 429.600 275.600 429.700 ;
        RECT 281.200 430.300 282.000 430.400 ;
        RECT 284.400 430.300 285.200 430.400 ;
        RECT 281.200 429.700 285.200 430.300 ;
        RECT 281.200 429.600 282.000 429.700 ;
        RECT 284.400 429.600 285.200 429.700 ;
        RECT 335.600 430.300 336.400 430.400 ;
        RECT 361.200 430.300 362.000 430.400 ;
        RECT 335.600 429.700 362.000 430.300 ;
        RECT 335.600 429.600 336.400 429.700 ;
        RECT 361.200 429.600 362.000 429.700 ;
        RECT 393.200 430.300 394.000 430.400 ;
        RECT 401.200 430.300 402.000 430.400 ;
        RECT 393.200 429.700 402.000 430.300 ;
        RECT 393.200 429.600 394.000 429.700 ;
        RECT 401.200 429.600 402.000 429.700 ;
        RECT 402.800 430.300 403.600 430.400 ;
        RECT 410.800 430.300 411.600 430.400 ;
        RECT 402.800 429.700 411.600 430.300 ;
        RECT 402.800 429.600 403.600 429.700 ;
        RECT 410.800 429.600 411.600 429.700 ;
        RECT 414.000 430.300 414.800 430.400 ;
        RECT 425.200 430.300 426.000 430.400 ;
        RECT 414.000 429.700 426.000 430.300 ;
        RECT 414.000 429.600 414.800 429.700 ;
        RECT 425.200 429.600 426.000 429.700 ;
        RECT 439.600 430.300 440.400 430.400 ;
        RECT 450.800 430.300 451.600 430.400 ;
        RECT 495.600 430.300 496.400 430.400 ;
        RECT 439.600 429.700 496.400 430.300 ;
        RECT 439.600 429.600 440.400 429.700 ;
        RECT 450.800 429.600 451.600 429.700 ;
        RECT 495.600 429.600 496.400 429.700 ;
        RECT 505.200 430.300 506.000 430.400 ;
        RECT 519.600 430.300 520.400 430.400 ;
        RECT 505.200 429.700 520.400 430.300 ;
        RECT 505.200 429.600 506.000 429.700 ;
        RECT 519.600 429.600 520.400 429.700 ;
        RECT 546.800 430.300 547.600 430.400 ;
        RECT 556.400 430.300 557.200 430.400 ;
        RECT 546.800 429.700 557.200 430.300 ;
        RECT 546.800 429.600 547.600 429.700 ;
        RECT 556.400 429.600 557.200 429.700 ;
        RECT 218.800 427.700 229.100 428.300 ;
        RECT 238.000 428.300 238.800 428.400 ;
        RECT 257.200 428.300 258.000 428.400 ;
        RECT 266.800 428.300 267.600 428.400 ;
        RECT 238.000 427.700 267.600 428.300 ;
        RECT 218.800 427.600 219.600 427.700 ;
        RECT 238.000 427.600 238.800 427.700 ;
        RECT 257.200 427.600 258.000 427.700 ;
        RECT 266.800 427.600 267.600 427.700 ;
        RECT 273.200 428.300 274.000 428.400 ;
        RECT 306.800 428.300 307.600 428.400 ;
        RECT 273.200 427.700 307.600 428.300 ;
        RECT 273.200 427.600 274.000 427.700 ;
        RECT 306.800 427.600 307.600 427.700 ;
        RECT 354.800 428.300 355.600 428.400 ;
        RECT 369.200 428.300 370.000 428.400 ;
        RECT 380.400 428.300 381.200 428.400 ;
        RECT 388.400 428.300 389.200 428.400 ;
        RECT 354.800 427.700 389.200 428.300 ;
        RECT 354.800 427.600 355.600 427.700 ;
        RECT 369.200 427.600 370.000 427.700 ;
        RECT 380.400 427.600 381.200 427.700 ;
        RECT 388.400 427.600 389.200 427.700 ;
        RECT 398.000 427.600 398.800 428.400 ;
        RECT 425.200 428.300 426.000 428.400 ;
        RECT 446.000 428.300 446.800 428.400 ;
        RECT 425.200 427.700 446.800 428.300 ;
        RECT 425.200 427.600 426.000 427.700 ;
        RECT 446.000 427.600 446.800 427.700 ;
        RECT 481.200 428.300 482.000 428.400 ;
        RECT 495.600 428.300 496.400 428.400 ;
        RECT 481.200 427.700 496.400 428.300 ;
        RECT 481.200 427.600 482.000 427.700 ;
        RECT 495.600 427.600 496.400 427.700 ;
        RECT 553.200 428.300 554.000 428.400 ;
        RECT 561.200 428.300 562.000 428.400 ;
        RECT 553.200 427.700 562.000 428.300 ;
        RECT 553.200 427.600 554.000 427.700 ;
        RECT 561.200 427.600 562.000 427.700 ;
        RECT 570.800 428.300 571.600 428.400 ;
        RECT 582.000 428.300 582.800 428.400 ;
        RECT 570.800 427.700 582.800 428.300 ;
        RECT 570.800 427.600 571.600 427.700 ;
        RECT 582.000 427.600 582.800 427.700 ;
        RECT 14.100 426.300 14.700 427.600 ;
        RECT 38.000 426.300 38.800 426.400 ;
        RECT 14.100 425.700 38.800 426.300 ;
        RECT 38.000 425.600 38.800 425.700 ;
        RECT 100.400 426.300 101.200 426.400 ;
        RECT 105.200 426.300 106.000 426.400 ;
        RECT 100.400 425.700 106.000 426.300 ;
        RECT 100.400 425.600 101.200 425.700 ;
        RECT 105.200 425.600 106.000 425.700 ;
        RECT 122.800 426.300 123.600 426.400 ;
        RECT 169.200 426.300 170.000 426.400 ;
        RECT 172.400 426.300 173.200 426.400 ;
        RECT 182.000 426.300 182.800 426.400 ;
        RECT 225.200 426.300 226.000 426.400 ;
        RECT 231.600 426.300 232.400 426.400 ;
        RECT 258.800 426.300 259.600 426.400 ;
        RECT 122.800 425.700 168.300 426.300 ;
        RECT 122.800 425.600 123.600 425.700 ;
        RECT 9.200 424.300 10.000 424.400 ;
        RECT 36.400 424.300 37.200 424.400 ;
        RECT 9.200 423.700 37.200 424.300 ;
        RECT 9.200 423.600 10.000 423.700 ;
        RECT 36.400 423.600 37.200 423.700 ;
        RECT 52.400 424.300 53.200 424.400 ;
        RECT 63.600 424.300 64.400 424.400 ;
        RECT 52.400 423.700 64.400 424.300 ;
        RECT 52.400 423.600 53.200 423.700 ;
        RECT 63.600 423.600 64.400 423.700 ;
        RECT 92.400 424.300 93.200 424.400 ;
        RECT 119.600 424.300 120.400 424.400 ;
        RECT 92.400 423.700 120.400 424.300 ;
        RECT 92.400 423.600 93.200 423.700 ;
        RECT 119.600 423.600 120.400 423.700 ;
        RECT 126.000 424.300 126.800 424.400 ;
        RECT 135.600 424.300 136.400 424.400 ;
        RECT 167.700 424.300 168.300 425.700 ;
        RECT 169.200 425.700 259.600 426.300 ;
        RECT 169.200 425.600 170.000 425.700 ;
        RECT 172.400 425.600 173.200 425.700 ;
        RECT 182.000 425.600 182.800 425.700 ;
        RECT 225.200 425.600 226.000 425.700 ;
        RECT 231.600 425.600 232.400 425.700 ;
        RECT 258.800 425.600 259.600 425.700 ;
        RECT 303.600 426.300 304.400 426.400 ;
        RECT 313.200 426.300 314.000 426.400 ;
        RECT 316.400 426.300 317.200 426.400 ;
        RECT 303.600 425.700 317.200 426.300 ;
        RECT 303.600 425.600 304.400 425.700 ;
        RECT 313.200 425.600 314.000 425.700 ;
        RECT 316.400 425.600 317.200 425.700 ;
        RECT 492.400 426.300 493.200 426.400 ;
        RECT 527.600 426.300 528.400 426.400 ;
        RECT 582.000 426.300 582.800 426.400 ;
        RECT 492.400 425.700 582.800 426.300 ;
        RECT 492.400 425.600 493.200 425.700 ;
        RECT 527.600 425.600 528.400 425.700 ;
        RECT 582.000 425.600 582.800 425.700 ;
        RECT 180.400 424.300 181.200 424.400 ;
        RECT 126.000 423.700 165.100 424.300 ;
        RECT 167.700 423.700 181.200 424.300 ;
        RECT 126.000 423.600 126.800 423.700 ;
        RECT 135.600 423.600 136.400 423.700 ;
        RECT 164.500 422.400 165.100 423.700 ;
        RECT 180.400 423.600 181.200 423.700 ;
        RECT 217.200 424.300 218.000 424.400 ;
        RECT 230.000 424.300 230.800 424.400 ;
        RECT 233.200 424.300 234.000 424.400 ;
        RECT 247.600 424.300 248.400 424.400 ;
        RECT 252.400 424.300 253.200 424.400 ;
        RECT 217.200 423.700 253.200 424.300 ;
        RECT 217.200 423.600 218.000 423.700 ;
        RECT 230.000 423.600 230.800 423.700 ;
        RECT 233.200 423.600 234.000 423.700 ;
        RECT 247.600 423.600 248.400 423.700 ;
        RECT 252.400 423.600 253.200 423.700 ;
        RECT 254.000 424.300 254.800 424.400 ;
        RECT 270.000 424.300 270.800 424.400 ;
        RECT 254.000 423.700 270.800 424.300 ;
        RECT 254.000 423.600 254.800 423.700 ;
        RECT 270.000 423.600 270.800 423.700 ;
        RECT 388.400 424.300 389.200 424.400 ;
        RECT 553.200 424.300 554.000 424.400 ;
        RECT 561.200 424.300 562.000 424.400 ;
        RECT 388.400 423.700 408.300 424.300 ;
        RECT 388.400 423.600 389.200 423.700 ;
        RECT 407.700 422.400 408.300 423.700 ;
        RECT 553.200 423.700 562.000 424.300 ;
        RECT 553.200 423.600 554.000 423.700 ;
        RECT 561.200 423.600 562.000 423.700 ;
        RECT 566.000 424.300 566.800 424.400 ;
        RECT 569.200 424.300 570.000 424.400 ;
        RECT 566.000 423.700 570.000 424.300 ;
        RECT 566.000 423.600 566.800 423.700 ;
        RECT 569.200 423.600 570.000 423.700 ;
        RECT 31.600 422.300 32.400 422.400 ;
        RECT 42.800 422.300 43.600 422.400 ;
        RECT 31.600 421.700 43.600 422.300 ;
        RECT 31.600 421.600 32.400 421.700 ;
        RECT 42.800 421.600 43.600 421.700 ;
        RECT 90.800 422.300 91.600 422.400 ;
        RECT 118.000 422.300 118.800 422.400 ;
        RECT 124.400 422.300 125.200 422.400 ;
        RECT 90.800 421.700 125.200 422.300 ;
        RECT 90.800 421.600 91.600 421.700 ;
        RECT 118.000 421.600 118.800 421.700 ;
        RECT 124.400 421.600 125.200 421.700 ;
        RECT 129.200 422.300 130.000 422.400 ;
        RECT 130.800 422.300 131.600 422.400 ;
        RECT 129.200 421.700 131.600 422.300 ;
        RECT 129.200 421.600 130.000 421.700 ;
        RECT 130.800 421.600 131.600 421.700 ;
        RECT 164.400 422.300 165.200 422.400 ;
        RECT 204.400 422.300 205.200 422.400 ;
        RECT 164.400 421.700 205.200 422.300 ;
        RECT 164.400 421.600 165.200 421.700 ;
        RECT 204.400 421.600 205.200 421.700 ;
        RECT 231.600 422.300 232.400 422.400 ;
        RECT 282.800 422.300 283.600 422.400 ;
        RECT 231.600 421.700 283.600 422.300 ;
        RECT 231.600 421.600 232.400 421.700 ;
        RECT 282.800 421.600 283.600 421.700 ;
        RECT 337.200 422.300 338.000 422.400 ;
        RECT 396.400 422.300 397.200 422.400 ;
        RECT 337.200 421.700 397.200 422.300 ;
        RECT 337.200 421.600 338.000 421.700 ;
        RECT 396.400 421.600 397.200 421.700 ;
        RECT 407.600 422.300 408.400 422.400 ;
        RECT 438.000 422.300 438.800 422.400 ;
        RECT 407.600 421.700 438.800 422.300 ;
        RECT 407.600 421.600 408.400 421.700 ;
        RECT 438.000 421.600 438.800 421.700 ;
        RECT 526.000 422.300 526.800 422.400 ;
        RECT 530.800 422.300 531.600 422.400 ;
        RECT 526.000 421.700 531.600 422.300 ;
        RECT 526.000 421.600 526.800 421.700 ;
        RECT 530.800 421.600 531.600 421.700 ;
        RECT 566.000 422.300 566.800 422.400 ;
        RECT 585.200 422.300 586.000 422.400 ;
        RECT 566.000 421.700 586.000 422.300 ;
        RECT 566.000 421.600 566.800 421.700 ;
        RECT 585.200 421.600 586.000 421.700 ;
        RECT 95.600 420.300 96.400 420.400 ;
        RECT 106.800 420.300 107.600 420.400 ;
        RECT 95.600 419.700 107.600 420.300 ;
        RECT 95.600 419.600 96.400 419.700 ;
        RECT 106.800 419.600 107.600 419.700 ;
        RECT 150.000 420.300 150.800 420.400 ;
        RECT 190.000 420.300 190.800 420.400 ;
        RECT 193.200 420.300 194.000 420.400 ;
        RECT 198.000 420.300 198.800 420.400 ;
        RECT 150.000 419.700 198.800 420.300 ;
        RECT 150.000 419.600 150.800 419.700 ;
        RECT 190.000 419.600 190.800 419.700 ;
        RECT 193.200 419.600 194.000 419.700 ;
        RECT 198.000 419.600 198.800 419.700 ;
        RECT 214.000 420.300 214.800 420.400 ;
        RECT 294.000 420.300 294.800 420.400 ;
        RECT 214.000 419.700 294.800 420.300 ;
        RECT 214.000 419.600 214.800 419.700 ;
        RECT 294.000 419.600 294.800 419.700 ;
        RECT 364.400 420.300 365.200 420.400 ;
        RECT 367.600 420.300 368.400 420.400 ;
        RECT 364.400 419.700 368.400 420.300 ;
        RECT 364.400 419.600 365.200 419.700 ;
        RECT 367.600 419.600 368.400 419.700 ;
        RECT 377.200 420.300 378.000 420.400 ;
        RECT 399.600 420.300 400.400 420.400 ;
        RECT 377.200 419.700 400.400 420.300 ;
        RECT 377.200 419.600 378.000 419.700 ;
        RECT 399.600 419.600 400.400 419.700 ;
        RECT 420.400 420.300 421.200 420.400 ;
        RECT 426.800 420.300 427.600 420.400 ;
        RECT 420.400 419.700 427.600 420.300 ;
        RECT 420.400 419.600 421.200 419.700 ;
        RECT 426.800 419.600 427.600 419.700 ;
        RECT 498.800 420.300 499.600 420.400 ;
        RECT 545.200 420.300 546.000 420.400 ;
        RECT 558.000 420.300 558.800 420.400 ;
        RECT 498.800 419.700 558.800 420.300 ;
        RECT 498.800 419.600 499.600 419.700 ;
        RECT 545.200 419.600 546.000 419.700 ;
        RECT 558.000 419.600 558.800 419.700 ;
        RECT 97.200 418.300 98.000 418.400 ;
        RECT 103.600 418.300 104.400 418.400 ;
        RECT 142.000 418.300 142.800 418.400 ;
        RECT 150.000 418.300 150.800 418.400 ;
        RECT 97.200 417.700 150.800 418.300 ;
        RECT 97.200 417.600 98.000 417.700 ;
        RECT 103.600 417.600 104.400 417.700 ;
        RECT 142.000 417.600 142.800 417.700 ;
        RECT 150.000 417.600 150.800 417.700 ;
        RECT 279.600 418.300 280.400 418.400 ;
        RECT 282.800 418.300 283.600 418.400 ;
        RECT 279.600 417.700 283.600 418.300 ;
        RECT 279.600 417.600 280.400 417.700 ;
        RECT 282.800 417.600 283.600 417.700 ;
        RECT 358.000 418.300 358.800 418.400 ;
        RECT 366.000 418.300 366.800 418.400 ;
        RECT 382.000 418.300 382.800 418.400 ;
        RECT 409.200 418.300 410.000 418.400 ;
        RECT 358.000 417.700 410.000 418.300 ;
        RECT 358.000 417.600 358.800 417.700 ;
        RECT 366.000 417.600 366.800 417.700 ;
        RECT 382.000 417.600 382.800 417.700 ;
        RECT 409.200 417.600 410.000 417.700 ;
        RECT 410.800 418.300 411.600 418.400 ;
        RECT 428.400 418.300 429.200 418.400 ;
        RECT 410.800 417.700 429.200 418.300 ;
        RECT 410.800 417.600 411.600 417.700 ;
        RECT 428.400 417.600 429.200 417.700 ;
        RECT 444.400 418.300 445.200 418.400 ;
        RECT 465.200 418.300 466.000 418.400 ;
        RECT 444.400 417.700 466.000 418.300 ;
        RECT 444.400 417.600 445.200 417.700 ;
        RECT 465.200 417.600 466.000 417.700 ;
        RECT 542.000 418.300 542.800 418.400 ;
        RECT 546.800 418.300 547.600 418.400 ;
        RECT 542.000 417.700 547.600 418.300 ;
        RECT 542.000 417.600 542.800 417.700 ;
        RECT 546.800 417.600 547.600 417.700 ;
        RECT 28.400 416.300 29.200 416.400 ;
        RECT 44.400 416.300 45.200 416.400 ;
        RECT 71.600 416.300 72.400 416.400 ;
        RECT 28.400 415.700 72.400 416.300 ;
        RECT 28.400 415.600 29.200 415.700 ;
        RECT 44.400 415.600 45.200 415.700 ;
        RECT 71.600 415.600 72.400 415.700 ;
        RECT 92.400 416.300 93.200 416.400 ;
        RECT 95.600 416.300 96.400 416.400 ;
        RECT 92.400 415.700 96.400 416.300 ;
        RECT 92.400 415.600 93.200 415.700 ;
        RECT 95.600 415.600 96.400 415.700 ;
        RECT 116.400 416.300 117.200 416.400 ;
        RECT 121.200 416.300 122.000 416.400 ;
        RECT 116.400 415.700 122.000 416.300 ;
        RECT 116.400 415.600 117.200 415.700 ;
        RECT 121.200 415.600 122.000 415.700 ;
        RECT 129.200 416.300 130.000 416.400 ;
        RECT 156.400 416.300 157.200 416.400 ;
        RECT 129.200 415.700 157.200 416.300 ;
        RECT 129.200 415.600 130.000 415.700 ;
        RECT 156.400 415.600 157.200 415.700 ;
        RECT 161.200 416.300 162.000 416.400 ;
        RECT 174.000 416.300 174.800 416.400 ;
        RECT 161.200 415.700 174.800 416.300 ;
        RECT 161.200 415.600 162.000 415.700 ;
        RECT 174.000 415.600 174.800 415.700 ;
        RECT 262.000 416.300 262.800 416.400 ;
        RECT 266.800 416.300 267.600 416.400 ;
        RECT 262.000 415.700 267.600 416.300 ;
        RECT 262.000 415.600 262.800 415.700 ;
        RECT 266.800 415.600 267.600 415.700 ;
        RECT 278.000 416.300 278.800 416.400 ;
        RECT 284.400 416.300 285.200 416.400 ;
        RECT 278.000 415.700 285.200 416.300 ;
        RECT 278.000 415.600 278.800 415.700 ;
        RECT 284.400 415.600 285.200 415.700 ;
        RECT 289.200 416.300 290.000 416.400 ;
        RECT 295.600 416.300 296.400 416.400 ;
        RECT 303.600 416.300 304.400 416.400 ;
        RECT 289.200 415.700 304.400 416.300 ;
        RECT 289.200 415.600 290.000 415.700 ;
        RECT 295.600 415.600 296.400 415.700 ;
        RECT 303.600 415.600 304.400 415.700 ;
        RECT 342.000 416.300 342.800 416.400 ;
        RECT 361.200 416.300 362.000 416.400 ;
        RECT 342.000 415.700 362.000 416.300 ;
        RECT 342.000 415.600 342.800 415.700 ;
        RECT 361.200 415.600 362.000 415.700 ;
        RECT 364.400 416.300 365.200 416.400 ;
        RECT 374.000 416.300 374.800 416.400 ;
        RECT 364.400 415.700 374.800 416.300 ;
        RECT 364.400 415.600 365.200 415.700 ;
        RECT 374.000 415.600 374.800 415.700 ;
        RECT 380.400 416.300 381.200 416.400 ;
        RECT 390.000 416.300 390.800 416.400 ;
        RECT 380.400 415.700 390.800 416.300 ;
        RECT 380.400 415.600 381.200 415.700 ;
        RECT 390.000 415.600 390.800 415.700 ;
        RECT 391.600 416.300 392.400 416.400 ;
        RECT 415.600 416.300 416.400 416.400 ;
        RECT 391.600 415.700 416.400 416.300 ;
        RECT 391.600 415.600 392.400 415.700 ;
        RECT 415.600 415.600 416.400 415.700 ;
        RECT 417.200 416.300 418.000 416.400 ;
        RECT 436.400 416.300 437.200 416.400 ;
        RECT 417.200 415.700 437.200 416.300 ;
        RECT 417.200 415.600 418.000 415.700 ;
        RECT 436.400 415.600 437.200 415.700 ;
        RECT 441.200 416.300 442.000 416.400 ;
        RECT 449.200 416.300 450.000 416.400 ;
        RECT 457.200 416.300 458.000 416.400 ;
        RECT 471.600 416.300 472.400 416.400 ;
        RECT 490.800 416.300 491.600 416.400 ;
        RECT 508.400 416.300 509.200 416.400 ;
        RECT 441.200 415.700 509.200 416.300 ;
        RECT 441.200 415.600 442.000 415.700 ;
        RECT 449.200 415.600 450.000 415.700 ;
        RECT 457.200 415.600 458.000 415.700 ;
        RECT 471.600 415.600 472.400 415.700 ;
        RECT 490.800 415.600 491.600 415.700 ;
        RECT 508.400 415.600 509.200 415.700 ;
        RECT 510.000 416.300 510.800 416.400 ;
        RECT 521.200 416.300 522.000 416.400 ;
        RECT 550.000 416.300 550.800 416.400 ;
        RECT 510.000 415.700 550.800 416.300 ;
        RECT 510.000 415.600 510.800 415.700 ;
        RECT 521.200 415.600 522.000 415.700 ;
        RECT 550.000 415.600 550.800 415.700 ;
        RECT 582.000 416.300 582.800 416.400 ;
        RECT 591.600 416.300 592.400 416.400 ;
        RECT 601.200 416.300 602.000 416.400 ;
        RECT 582.000 415.700 602.000 416.300 ;
        RECT 582.000 415.600 582.800 415.700 ;
        RECT 591.600 415.600 592.400 415.700 ;
        RECT 601.200 415.600 602.000 415.700 ;
        RECT 7.600 414.300 8.400 414.400 ;
        RECT 14.000 414.300 14.800 414.400 ;
        RECT 7.600 413.700 14.800 414.300 ;
        RECT 7.600 413.600 8.400 413.700 ;
        RECT 14.000 413.600 14.800 413.700 ;
        RECT 55.600 414.300 56.400 414.400 ;
        RECT 62.000 414.300 62.800 414.400 ;
        RECT 55.600 413.700 62.800 414.300 ;
        RECT 55.600 413.600 56.400 413.700 ;
        RECT 62.000 413.600 62.800 413.700 ;
        RECT 63.600 414.300 64.400 414.400 ;
        RECT 81.200 414.300 82.000 414.400 ;
        RECT 84.400 414.300 85.200 414.400 ;
        RECT 63.600 413.700 85.200 414.300 ;
        RECT 63.600 413.600 64.400 413.700 ;
        RECT 81.200 413.600 82.000 413.700 ;
        RECT 84.400 413.600 85.200 413.700 ;
        RECT 108.400 414.300 109.200 414.400 ;
        RECT 132.400 414.300 133.200 414.400 ;
        RECT 108.400 413.700 133.200 414.300 ;
        RECT 108.400 413.600 109.200 413.700 ;
        RECT 132.400 413.600 133.200 413.700 ;
        RECT 138.800 414.300 139.600 414.400 ;
        RECT 145.200 414.300 146.000 414.400 ;
        RECT 138.800 413.700 146.000 414.300 ;
        RECT 138.800 413.600 139.600 413.700 ;
        RECT 145.200 413.600 146.000 413.700 ;
        RECT 167.600 414.300 168.400 414.400 ;
        RECT 175.600 414.300 176.400 414.400 ;
        RECT 167.600 413.700 176.400 414.300 ;
        RECT 167.600 413.600 168.400 413.700 ;
        RECT 175.600 413.600 176.400 413.700 ;
        RECT 194.800 414.300 195.600 414.400 ;
        RECT 215.600 414.300 216.400 414.400 ;
        RECT 194.800 413.700 216.400 414.300 ;
        RECT 194.800 413.600 195.600 413.700 ;
        RECT 215.600 413.600 216.400 413.700 ;
        RECT 230.000 414.300 230.800 414.400 ;
        RECT 234.800 414.300 235.600 414.400 ;
        RECT 230.000 413.700 235.600 414.300 ;
        RECT 230.000 413.600 230.800 413.700 ;
        RECT 234.800 413.600 235.600 413.700 ;
        RECT 238.000 414.300 238.800 414.400 ;
        RECT 247.600 414.300 248.400 414.400 ;
        RECT 238.000 413.700 248.400 414.300 ;
        RECT 238.000 413.600 238.800 413.700 ;
        RECT 247.600 413.600 248.400 413.700 ;
        RECT 263.600 414.300 264.400 414.400 ;
        RECT 298.800 414.300 299.600 414.400 ;
        RECT 313.200 414.300 314.000 414.400 ;
        RECT 263.600 413.700 280.300 414.300 ;
        RECT 263.600 413.600 264.400 413.700 ;
        RECT 279.700 412.400 280.300 413.700 ;
        RECT 298.800 413.700 314.000 414.300 ;
        RECT 298.800 413.600 299.600 413.700 ;
        RECT 313.200 413.600 314.000 413.700 ;
        RECT 354.800 414.300 355.600 414.400 ;
        RECT 370.800 414.300 371.600 414.400 ;
        RECT 354.800 413.700 371.600 414.300 ;
        RECT 354.800 413.600 355.600 413.700 ;
        RECT 370.800 413.600 371.600 413.700 ;
        RECT 372.400 414.300 373.200 414.400 ;
        RECT 401.200 414.300 402.000 414.400 ;
        RECT 372.400 413.700 402.000 414.300 ;
        RECT 372.400 413.600 373.200 413.700 ;
        RECT 401.200 413.600 402.000 413.700 ;
        RECT 402.800 414.300 403.600 414.400 ;
        RECT 434.800 414.300 435.600 414.400 ;
        RECT 452.400 414.300 453.200 414.400 ;
        RECT 402.800 413.700 453.200 414.300 ;
        RECT 402.800 413.600 403.600 413.700 ;
        RECT 434.800 413.600 435.600 413.700 ;
        RECT 452.400 413.600 453.200 413.700 ;
        RECT 460.400 414.300 461.200 414.400 ;
        RECT 466.800 414.300 467.600 414.400 ;
        RECT 474.800 414.300 475.600 414.400 ;
        RECT 460.400 413.700 475.600 414.300 ;
        RECT 460.400 413.600 461.200 413.700 ;
        RECT 466.800 413.600 467.600 413.700 ;
        RECT 474.800 413.600 475.600 413.700 ;
        RECT 495.600 414.300 496.400 414.400 ;
        RECT 505.200 414.300 506.000 414.400 ;
        RECT 495.600 413.700 506.000 414.300 ;
        RECT 495.600 413.600 496.400 413.700 ;
        RECT 505.200 413.600 506.000 413.700 ;
        RECT 510.000 414.300 510.800 414.400 ;
        RECT 514.800 414.300 515.600 414.400 ;
        RECT 535.600 414.300 536.400 414.400 ;
        RECT 546.800 414.300 547.600 414.400 ;
        RECT 551.600 414.300 552.400 414.400 ;
        RECT 510.000 413.700 552.400 414.300 ;
        RECT 510.000 413.600 510.800 413.700 ;
        RECT 514.800 413.600 515.600 413.700 ;
        RECT 535.600 413.600 536.400 413.700 ;
        RECT 546.800 413.600 547.600 413.700 ;
        RECT 551.600 413.600 552.400 413.700 ;
        RECT 588.400 414.300 589.200 414.400 ;
        RECT 590.000 414.300 590.800 414.400 ;
        RECT 588.400 413.700 590.800 414.300 ;
        RECT 588.400 413.600 589.200 413.700 ;
        RECT 590.000 413.600 590.800 413.700 ;
        RECT 25.200 412.300 26.000 412.400 ;
        RECT 33.200 412.300 34.000 412.400 ;
        RECT 25.200 411.700 34.000 412.300 ;
        RECT 25.200 411.600 26.000 411.700 ;
        RECT 33.200 411.600 34.000 411.700 ;
        RECT 47.600 412.300 48.400 412.400 ;
        RECT 58.800 412.300 59.600 412.400 ;
        RECT 47.600 411.700 59.600 412.300 ;
        RECT 47.600 411.600 48.400 411.700 ;
        RECT 58.800 411.600 59.600 411.700 ;
        RECT 60.400 412.300 61.200 412.400 ;
        RECT 70.000 412.300 70.800 412.400 ;
        RECT 60.400 411.700 70.800 412.300 ;
        RECT 60.400 411.600 61.200 411.700 ;
        RECT 70.000 411.600 70.800 411.700 ;
        RECT 71.600 412.300 72.400 412.400 ;
        RECT 94.000 412.300 94.800 412.400 ;
        RECT 110.000 412.300 110.800 412.400 ;
        RECT 71.600 411.700 110.800 412.300 ;
        RECT 71.600 411.600 72.400 411.700 ;
        RECT 94.000 411.600 94.800 411.700 ;
        RECT 110.000 411.600 110.800 411.700 ;
        RECT 113.200 412.300 114.000 412.400 ;
        RECT 119.600 412.300 120.400 412.400 ;
        RECT 113.200 411.700 120.400 412.300 ;
        RECT 113.200 411.600 114.000 411.700 ;
        RECT 119.600 411.600 120.400 411.700 ;
        RECT 156.400 412.300 157.200 412.400 ;
        RECT 161.200 412.300 162.000 412.400 ;
        RECT 169.200 412.300 170.000 412.400 ;
        RECT 156.400 411.700 170.000 412.300 ;
        RECT 156.400 411.600 157.200 411.700 ;
        RECT 161.200 411.600 162.000 411.700 ;
        RECT 169.200 411.600 170.000 411.700 ;
        RECT 177.200 412.300 178.000 412.400 ;
        RECT 180.400 412.300 181.200 412.400 ;
        RECT 177.200 411.700 181.200 412.300 ;
        RECT 177.200 411.600 178.000 411.700 ;
        RECT 180.400 411.600 181.200 411.700 ;
        RECT 234.800 412.300 235.600 412.400 ;
        RECT 239.600 412.300 240.400 412.400 ;
        RECT 258.800 412.300 259.600 412.400 ;
        RECT 234.800 411.700 259.600 412.300 ;
        RECT 234.800 411.600 235.600 411.700 ;
        RECT 239.600 411.600 240.400 411.700 ;
        RECT 258.800 411.600 259.600 411.700 ;
        RECT 265.200 412.300 266.000 412.400 ;
        RECT 278.000 412.300 278.800 412.400 ;
        RECT 265.200 411.700 278.800 412.300 ;
        RECT 265.200 411.600 266.000 411.700 ;
        RECT 278.000 411.600 278.800 411.700 ;
        RECT 279.600 412.300 280.400 412.400 ;
        RECT 286.000 412.300 286.800 412.400 ;
        RECT 279.600 411.700 286.800 412.300 ;
        RECT 279.600 411.600 280.400 411.700 ;
        RECT 286.000 411.600 286.800 411.700 ;
        RECT 300.400 412.300 301.200 412.400 ;
        RECT 316.400 412.300 317.200 412.400 ;
        RECT 337.200 412.300 338.000 412.400 ;
        RECT 300.400 411.700 338.000 412.300 ;
        RECT 300.400 411.600 301.200 411.700 ;
        RECT 316.400 411.600 317.200 411.700 ;
        RECT 337.200 411.600 338.000 411.700 ;
        RECT 356.400 412.300 357.200 412.400 ;
        RECT 372.400 412.300 373.200 412.400 ;
        RECT 356.400 411.700 373.200 412.300 ;
        RECT 356.400 411.600 357.200 411.700 ;
        RECT 372.400 411.600 373.200 411.700 ;
        RECT 375.600 412.300 376.400 412.400 ;
        RECT 383.600 412.300 384.400 412.400 ;
        RECT 375.600 411.700 384.400 412.300 ;
        RECT 375.600 411.600 376.400 411.700 ;
        RECT 383.600 411.600 384.400 411.700 ;
        RECT 396.400 412.300 397.200 412.400 ;
        RECT 402.800 412.300 403.600 412.400 ;
        RECT 396.400 411.700 403.600 412.300 ;
        RECT 396.400 411.600 397.200 411.700 ;
        RECT 402.800 411.600 403.600 411.700 ;
        RECT 406.000 412.300 406.800 412.400 ;
        RECT 410.800 412.300 411.600 412.400 ;
        RECT 406.000 411.700 411.600 412.300 ;
        RECT 406.000 411.600 406.800 411.700 ;
        RECT 410.800 411.600 411.600 411.700 ;
        RECT 415.600 412.300 416.400 412.400 ;
        RECT 422.000 412.300 422.800 412.400 ;
        RECT 415.600 411.700 422.800 412.300 ;
        RECT 415.600 411.600 416.400 411.700 ;
        RECT 422.000 411.600 422.800 411.700 ;
        RECT 436.400 412.300 437.200 412.400 ;
        RECT 463.600 412.300 464.400 412.400 ;
        RECT 471.600 412.300 472.400 412.400 ;
        RECT 436.400 411.700 472.400 412.300 ;
        RECT 436.400 411.600 437.200 411.700 ;
        RECT 463.600 411.600 464.400 411.700 ;
        RECT 471.600 411.600 472.400 411.700 ;
        RECT 489.200 412.300 490.000 412.400 ;
        RECT 498.800 412.300 499.600 412.400 ;
        RECT 489.200 411.700 499.600 412.300 ;
        RECT 489.200 411.600 490.000 411.700 ;
        RECT 498.800 411.600 499.600 411.700 ;
        RECT 505.200 412.300 506.000 412.400 ;
        RECT 510.000 412.300 510.800 412.400 ;
        RECT 505.200 411.700 510.800 412.300 ;
        RECT 505.200 411.600 506.000 411.700 ;
        RECT 510.000 411.600 510.800 411.700 ;
        RECT 513.200 412.300 514.000 412.400 ;
        RECT 516.400 412.300 517.200 412.400 ;
        RECT 532.400 412.300 533.200 412.400 ;
        RECT 545.200 412.300 546.000 412.400 ;
        RECT 569.200 412.300 570.000 412.400 ;
        RECT 513.200 411.700 570.000 412.300 ;
        RECT 513.200 411.600 514.000 411.700 ;
        RECT 516.400 411.600 517.200 411.700 ;
        RECT 532.400 411.600 533.200 411.700 ;
        RECT 545.200 411.600 546.000 411.700 ;
        RECT 569.200 411.600 570.000 411.700 ;
        RECT 47.600 410.300 48.400 410.400 ;
        RECT 50.800 410.300 51.600 410.400 ;
        RECT 82.800 410.300 83.600 410.400 ;
        RECT 97.200 410.300 98.000 410.400 ;
        RECT 47.600 409.700 98.000 410.300 ;
        RECT 47.600 409.600 48.400 409.700 ;
        RECT 50.800 409.600 51.600 409.700 ;
        RECT 82.800 409.600 83.600 409.700 ;
        RECT 97.200 409.600 98.000 409.700 ;
        RECT 100.400 410.300 101.200 410.400 ;
        RECT 103.600 410.300 104.400 410.400 ;
        RECT 100.400 409.700 104.400 410.300 ;
        RECT 100.400 409.600 101.200 409.700 ;
        RECT 103.600 409.600 104.400 409.700 ;
        RECT 148.400 410.300 149.200 410.400 ;
        RECT 161.200 410.300 162.000 410.400 ;
        RECT 148.400 409.700 162.000 410.300 ;
        RECT 148.400 409.600 149.200 409.700 ;
        RECT 161.200 409.600 162.000 409.700 ;
        RECT 167.600 409.600 168.400 410.400 ;
        RECT 223.600 410.300 224.400 410.400 ;
        RECT 242.800 410.300 243.600 410.400 ;
        RECT 223.600 409.700 243.600 410.300 ;
        RECT 223.600 409.600 224.400 409.700 ;
        RECT 242.800 409.600 243.600 409.700 ;
        RECT 278.000 410.300 278.800 410.400 ;
        RECT 282.800 410.300 283.600 410.400 ;
        RECT 278.000 409.700 283.600 410.300 ;
        RECT 278.000 409.600 278.800 409.700 ;
        RECT 282.800 409.600 283.600 409.700 ;
        RECT 353.200 410.300 354.000 410.400 ;
        RECT 359.600 410.300 360.400 410.400 ;
        RECT 377.200 410.300 378.000 410.400 ;
        RECT 353.200 409.700 378.000 410.300 ;
        RECT 353.200 409.600 354.000 409.700 ;
        RECT 359.600 409.600 360.400 409.700 ;
        RECT 377.200 409.600 378.000 409.700 ;
        RECT 382.000 410.300 382.800 410.400 ;
        RECT 393.200 410.300 394.000 410.400 ;
        RECT 382.000 409.700 394.000 410.300 ;
        RECT 382.000 409.600 382.800 409.700 ;
        RECT 393.200 409.600 394.000 409.700 ;
        RECT 394.800 410.300 395.600 410.400 ;
        RECT 401.200 410.300 402.000 410.400 ;
        RECT 441.200 410.300 442.000 410.400 ;
        RECT 394.800 409.700 442.000 410.300 ;
        RECT 394.800 409.600 395.600 409.700 ;
        RECT 401.200 409.600 402.000 409.700 ;
        RECT 441.200 409.600 442.000 409.700 ;
        RECT 447.600 410.300 448.400 410.400 ;
        RECT 484.400 410.300 485.200 410.400 ;
        RECT 447.600 409.700 485.200 410.300 ;
        RECT 447.600 409.600 448.400 409.700 ;
        RECT 484.400 409.600 485.200 409.700 ;
        RECT 502.000 410.300 502.800 410.400 ;
        RECT 516.400 410.300 517.200 410.400 ;
        RECT 502.000 409.700 517.200 410.300 ;
        RECT 502.000 409.600 502.800 409.700 ;
        RECT 516.400 409.600 517.200 409.700 ;
        RECT 518.000 410.300 518.800 410.400 ;
        RECT 521.200 410.300 522.000 410.400 ;
        RECT 518.000 409.700 522.000 410.300 ;
        RECT 518.000 409.600 518.800 409.700 ;
        RECT 521.200 409.600 522.000 409.700 ;
        RECT 161.200 408.300 162.000 408.400 ;
        RECT 170.800 408.300 171.600 408.400 ;
        RECT 161.200 407.700 171.600 408.300 ;
        RECT 161.200 407.600 162.000 407.700 ;
        RECT 170.800 407.600 171.600 407.700 ;
        RECT 218.800 408.300 219.600 408.400 ;
        RECT 233.200 408.300 234.000 408.400 ;
        RECT 218.800 407.700 234.000 408.300 ;
        RECT 218.800 407.600 219.600 407.700 ;
        RECT 233.200 407.600 234.000 407.700 ;
        RECT 290.800 408.300 291.600 408.400 ;
        RECT 332.400 408.300 333.200 408.400 ;
        RECT 343.600 408.300 344.400 408.400 ;
        RECT 290.800 407.700 344.400 408.300 ;
        RECT 290.800 407.600 291.600 407.700 ;
        RECT 332.400 407.600 333.200 407.700 ;
        RECT 343.600 407.600 344.400 407.700 ;
        RECT 391.600 408.300 392.400 408.400 ;
        RECT 394.800 408.300 395.600 408.400 ;
        RECT 391.600 407.700 395.600 408.300 ;
        RECT 391.600 407.600 392.400 407.700 ;
        RECT 394.800 407.600 395.600 407.700 ;
        RECT 423.600 408.300 424.400 408.400 ;
        RECT 426.800 408.300 427.600 408.400 ;
        RECT 433.200 408.300 434.000 408.400 ;
        RECT 447.700 408.300 448.300 409.600 ;
        RECT 423.600 407.700 448.300 408.300 ;
        RECT 465.200 408.300 466.000 408.400 ;
        RECT 473.200 408.300 474.000 408.400 ;
        RECT 486.000 408.300 486.800 408.400 ;
        RECT 556.400 408.300 557.200 408.400 ;
        RECT 567.600 408.300 568.400 408.400 ;
        RECT 465.200 407.700 568.400 408.300 ;
        RECT 423.600 407.600 424.400 407.700 ;
        RECT 426.800 407.600 427.600 407.700 ;
        RECT 433.200 407.600 434.000 407.700 ;
        RECT 465.200 407.600 466.000 407.700 ;
        RECT 473.200 407.600 474.000 407.700 ;
        RECT 486.000 407.600 486.800 407.700 ;
        RECT 556.400 407.600 557.200 407.700 ;
        RECT 567.600 407.600 568.400 407.700 ;
        RECT 86.000 406.300 86.800 406.400 ;
        RECT 92.400 406.300 93.200 406.400 ;
        RECT 86.000 405.700 93.200 406.300 ;
        RECT 86.000 405.600 86.800 405.700 ;
        RECT 92.400 405.600 93.200 405.700 ;
        RECT 158.000 406.300 158.800 406.400 ;
        RECT 162.800 406.300 163.600 406.400 ;
        RECT 158.000 405.700 163.600 406.300 ;
        RECT 158.000 405.600 158.800 405.700 ;
        RECT 162.800 405.600 163.600 405.700 ;
        RECT 399.600 406.300 400.400 406.400 ;
        RECT 474.800 406.300 475.600 406.400 ;
        RECT 399.600 405.700 475.600 406.300 ;
        RECT 399.600 405.600 400.400 405.700 ;
        RECT 474.800 405.600 475.600 405.700 ;
        RECT 65.200 404.300 66.000 404.400 ;
        RECT 90.800 404.300 91.600 404.400 ;
        RECT 95.600 404.300 96.400 404.400 ;
        RECT 127.600 404.300 128.400 404.400 ;
        RECT 65.200 403.700 128.400 404.300 ;
        RECT 65.200 403.600 66.000 403.700 ;
        RECT 90.800 403.600 91.600 403.700 ;
        RECT 95.600 403.600 96.400 403.700 ;
        RECT 127.600 403.600 128.400 403.700 ;
        RECT 257.200 404.300 258.000 404.400 ;
        RECT 263.600 404.300 264.400 404.400 ;
        RECT 257.200 403.700 264.400 404.300 ;
        RECT 257.200 403.600 258.000 403.700 ;
        RECT 263.600 403.600 264.400 403.700 ;
        RECT 423.600 404.300 424.400 404.400 ;
        RECT 490.800 404.300 491.600 404.400 ;
        RECT 423.600 403.700 491.600 404.300 ;
        RECT 423.600 403.600 424.400 403.700 ;
        RECT 490.800 403.600 491.600 403.700 ;
        RECT 55.600 402.300 56.400 402.400 ;
        RECT 74.800 402.300 75.600 402.400 ;
        RECT 79.600 402.300 80.400 402.400 ;
        RECT 55.600 401.700 80.400 402.300 ;
        RECT 55.600 401.600 56.400 401.700 ;
        RECT 74.800 401.600 75.600 401.700 ;
        RECT 79.600 401.600 80.400 401.700 ;
        RECT 202.800 401.600 203.600 402.400 ;
        RECT 508.400 402.300 509.200 402.400 ;
        RECT 554.800 402.300 555.600 402.400 ;
        RECT 508.400 401.700 555.600 402.300 ;
        RECT 508.400 401.600 509.200 401.700 ;
        RECT 554.800 401.600 555.600 401.700 ;
        RECT 177.200 400.300 178.000 400.400 ;
        RECT 186.800 400.300 187.600 400.400 ;
        RECT 222.000 400.300 222.800 400.400 ;
        RECT 177.200 399.700 185.900 400.300 ;
        RECT 177.200 399.600 178.000 399.700 ;
        RECT 46.000 397.600 46.800 398.400 ;
        RECT 66.800 398.300 67.600 398.400 ;
        RECT 167.600 398.300 168.400 398.400 ;
        RECT 66.800 397.700 168.400 398.300 ;
        RECT 185.300 398.300 185.900 399.700 ;
        RECT 186.800 399.700 222.800 400.300 ;
        RECT 186.800 399.600 187.600 399.700 ;
        RECT 222.000 399.600 222.800 399.700 ;
        RECT 326.000 400.300 326.800 400.400 ;
        RECT 337.200 400.300 338.000 400.400 ;
        RECT 326.000 399.700 338.000 400.300 ;
        RECT 326.000 399.600 326.800 399.700 ;
        RECT 337.200 399.600 338.000 399.700 ;
        RECT 370.800 400.300 371.600 400.400 ;
        RECT 382.000 400.300 382.800 400.400 ;
        RECT 370.800 399.700 382.800 400.300 ;
        RECT 370.800 399.600 371.600 399.700 ;
        RECT 382.000 399.600 382.800 399.700 ;
        RECT 484.400 400.300 485.200 400.400 ;
        RECT 503.600 400.300 504.400 400.400 ;
        RECT 510.000 400.300 510.800 400.400 ;
        RECT 558.000 400.300 558.800 400.400 ;
        RECT 484.400 399.700 558.800 400.300 ;
        RECT 484.400 399.600 485.200 399.700 ;
        RECT 503.600 399.600 504.400 399.700 ;
        RECT 510.000 399.600 510.800 399.700 ;
        RECT 558.000 399.600 558.800 399.700 ;
        RECT 599.600 400.300 600.400 400.400 ;
        RECT 604.400 400.300 605.200 400.400 ;
        RECT 606.000 400.300 606.800 400.400 ;
        RECT 599.600 399.700 606.800 400.300 ;
        RECT 599.600 399.600 600.400 399.700 ;
        RECT 604.400 399.600 605.200 399.700 ;
        RECT 606.000 399.600 606.800 399.700 ;
        RECT 204.400 398.300 205.200 398.400 ;
        RECT 185.300 397.700 205.200 398.300 ;
        RECT 66.800 397.600 67.600 397.700 ;
        RECT 167.600 397.600 168.400 397.700 ;
        RECT 204.400 397.600 205.200 397.700 ;
        RECT 282.800 398.300 283.600 398.400 ;
        RECT 292.400 398.300 293.200 398.400 ;
        RECT 297.200 398.300 298.000 398.400 ;
        RECT 282.800 397.700 298.000 398.300 ;
        RECT 282.800 397.600 283.600 397.700 ;
        RECT 292.400 397.600 293.200 397.700 ;
        RECT 297.200 397.600 298.000 397.700 ;
        RECT 329.200 398.300 330.000 398.400 ;
        RECT 340.400 398.300 341.200 398.400 ;
        RECT 342.000 398.300 342.800 398.400 ;
        RECT 329.200 397.700 342.800 398.300 ;
        RECT 329.200 397.600 330.000 397.700 ;
        RECT 340.400 397.600 341.200 397.700 ;
        RECT 342.000 397.600 342.800 397.700 ;
        RECT 383.600 398.300 384.400 398.400 ;
        RECT 393.200 398.300 394.000 398.400 ;
        RECT 383.600 397.700 394.000 398.300 ;
        RECT 383.600 397.600 384.400 397.700 ;
        RECT 393.200 397.600 394.000 397.700 ;
        RECT 430.000 398.300 430.800 398.400 ;
        RECT 442.800 398.300 443.600 398.400 ;
        RECT 430.000 397.700 443.600 398.300 ;
        RECT 430.000 397.600 430.800 397.700 ;
        RECT 442.800 397.600 443.600 397.700 ;
        RECT 529.200 398.300 530.000 398.400 ;
        RECT 551.600 398.300 552.400 398.400 ;
        RECT 529.200 397.700 552.400 398.300 ;
        RECT 529.200 397.600 530.000 397.700 ;
        RECT 551.600 397.600 552.400 397.700 ;
        RECT 506.800 396.300 507.600 396.400 ;
        RECT 612.400 396.300 613.200 396.400 ;
        RECT 506.800 395.700 613.200 396.300 ;
        RECT 506.800 395.600 507.600 395.700 ;
        RECT 612.400 395.600 613.200 395.700 ;
        RECT 132.400 394.300 133.200 394.400 ;
        RECT 209.200 394.300 210.000 394.400 ;
        RECT 132.400 393.700 210.000 394.300 ;
        RECT 132.400 393.600 133.200 393.700 ;
        RECT 209.200 393.600 210.000 393.700 ;
        RECT 246.000 394.300 246.800 394.400 ;
        RECT 249.200 394.300 250.000 394.400 ;
        RECT 254.000 394.300 254.800 394.400 ;
        RECT 246.000 393.700 254.800 394.300 ;
        RECT 246.000 393.600 246.800 393.700 ;
        RECT 249.200 393.600 250.000 393.700 ;
        RECT 254.000 393.600 254.800 393.700 ;
        RECT 409.200 394.300 410.000 394.400 ;
        RECT 446.000 394.300 446.800 394.400 ;
        RECT 409.200 393.700 446.800 394.300 ;
        RECT 409.200 393.600 410.000 393.700 ;
        RECT 446.000 393.600 446.800 393.700 ;
        RECT 516.400 394.300 517.200 394.400 ;
        RECT 561.200 394.300 562.000 394.400 ;
        RECT 516.400 393.700 562.000 394.300 ;
        RECT 516.400 393.600 517.200 393.700 ;
        RECT 561.200 393.600 562.000 393.700 ;
        RECT 54.000 392.300 54.800 392.400 ;
        RECT 86.000 392.300 86.800 392.400 ;
        RECT 54.000 391.700 86.800 392.300 ;
        RECT 54.000 391.600 54.800 391.700 ;
        RECT 86.000 391.600 86.800 391.700 ;
        RECT 90.800 392.300 91.600 392.400 ;
        RECT 97.200 392.300 98.000 392.400 ;
        RECT 90.800 391.700 98.000 392.300 ;
        RECT 90.800 391.600 91.600 391.700 ;
        RECT 97.200 391.600 98.000 391.700 ;
        RECT 106.800 392.300 107.600 392.400 ;
        RECT 111.600 392.300 112.400 392.400 ;
        RECT 106.800 391.700 112.400 392.300 ;
        RECT 106.800 391.600 107.600 391.700 ;
        RECT 111.600 391.600 112.400 391.700 ;
        RECT 130.800 392.300 131.600 392.400 ;
        RECT 137.200 392.300 138.000 392.400 ;
        RECT 130.800 391.700 138.000 392.300 ;
        RECT 130.800 391.600 131.600 391.700 ;
        RECT 137.200 391.600 138.000 391.700 ;
        RECT 212.400 392.300 213.200 392.400 ;
        RECT 225.200 392.300 226.000 392.400 ;
        RECT 252.400 392.300 253.200 392.400 ;
        RECT 212.400 391.700 219.500 392.300 ;
        RECT 212.400 391.600 213.200 391.700 ;
        RECT 36.400 390.300 37.200 390.400 ;
        RECT 39.600 390.300 40.400 390.400 ;
        RECT 36.400 389.700 40.400 390.300 ;
        RECT 36.400 389.600 37.200 389.700 ;
        RECT 39.600 389.600 40.400 389.700 ;
        RECT 46.000 390.300 46.800 390.400 ;
        RECT 58.800 390.300 59.600 390.400 ;
        RECT 66.800 390.300 67.600 390.400 ;
        RECT 46.000 389.700 67.600 390.300 ;
        RECT 46.000 389.600 46.800 389.700 ;
        RECT 58.800 389.600 59.600 389.700 ;
        RECT 66.800 389.600 67.600 389.700 ;
        RECT 74.800 390.300 75.600 390.400 ;
        RECT 86.000 390.300 86.800 390.400 ;
        RECT 74.800 389.700 86.800 390.300 ;
        RECT 74.800 389.600 75.600 389.700 ;
        RECT 86.000 389.600 86.800 389.700 ;
        RECT 108.400 390.300 109.200 390.400 ;
        RECT 118.000 390.300 118.800 390.400 ;
        RECT 108.400 389.700 118.800 390.300 ;
        RECT 108.400 389.600 109.200 389.700 ;
        RECT 118.000 389.600 118.800 389.700 ;
        RECT 119.600 390.300 120.400 390.400 ;
        RECT 138.800 390.300 139.600 390.400 ;
        RECT 119.600 389.700 139.600 390.300 ;
        RECT 119.600 389.600 120.400 389.700 ;
        RECT 138.800 389.600 139.600 389.700 ;
        RECT 198.000 390.300 198.800 390.400 ;
        RECT 217.200 390.300 218.000 390.400 ;
        RECT 198.000 389.700 218.000 390.300 ;
        RECT 218.900 390.300 219.500 391.700 ;
        RECT 225.200 391.700 253.200 392.300 ;
        RECT 225.200 391.600 226.000 391.700 ;
        RECT 252.400 391.600 253.200 391.700 ;
        RECT 489.200 392.300 490.000 392.400 ;
        RECT 513.200 392.300 514.000 392.400 ;
        RECT 489.200 391.700 514.000 392.300 ;
        RECT 489.200 391.600 490.000 391.700 ;
        RECT 513.200 391.600 514.000 391.700 ;
        RECT 548.400 392.300 549.200 392.400 ;
        RECT 566.000 392.300 566.800 392.400 ;
        RECT 548.400 391.700 566.800 392.300 ;
        RECT 548.400 391.600 549.200 391.700 ;
        RECT 566.000 391.600 566.800 391.700 ;
        RECT 252.400 390.300 253.200 390.400 ;
        RECT 218.900 389.700 253.200 390.300 ;
        RECT 198.000 389.600 198.800 389.700 ;
        RECT 217.200 389.600 218.000 389.700 ;
        RECT 252.400 389.600 253.200 389.700 ;
        RECT 263.600 390.300 264.400 390.400 ;
        RECT 266.800 390.300 267.600 390.400 ;
        RECT 401.200 390.300 402.000 390.400 ;
        RECT 263.600 389.700 402.000 390.300 ;
        RECT 263.600 389.600 264.400 389.700 ;
        RECT 266.800 389.600 267.600 389.700 ;
        RECT 401.200 389.600 402.000 389.700 ;
        RECT 450.800 390.300 451.600 390.400 ;
        RECT 508.400 390.300 509.200 390.400 ;
        RECT 450.800 389.700 509.200 390.300 ;
        RECT 450.800 389.600 451.600 389.700 ;
        RECT 508.400 389.600 509.200 389.700 ;
        RECT 550.000 390.300 550.800 390.400 ;
        RECT 556.400 390.300 557.200 390.400 ;
        RECT 550.000 389.700 557.200 390.300 ;
        RECT 550.000 389.600 550.800 389.700 ;
        RECT 556.400 389.600 557.200 389.700 ;
        RECT 558.000 390.300 558.800 390.400 ;
        RECT 561.200 390.300 562.000 390.400 ;
        RECT 558.000 389.700 562.000 390.300 ;
        RECT 558.000 389.600 558.800 389.700 ;
        RECT 561.200 389.600 562.000 389.700 ;
        RECT 572.400 390.300 573.200 390.400 ;
        RECT 586.800 390.300 587.600 390.400 ;
        RECT 572.400 389.700 587.600 390.300 ;
        RECT 572.400 389.600 573.200 389.700 ;
        RECT 586.800 389.600 587.600 389.700 ;
        RECT 39.600 388.300 40.400 388.400 ;
        RECT 42.800 388.300 43.600 388.400 ;
        RECT 55.600 388.300 56.400 388.400 ;
        RECT 78.000 388.300 78.800 388.400 ;
        RECT 98.800 388.300 99.600 388.400 ;
        RECT 108.500 388.300 109.100 389.600 ;
        RECT 39.600 387.700 109.100 388.300 ;
        RECT 114.800 388.300 115.600 388.400 ;
        RECT 156.400 388.300 157.200 388.400 ;
        RECT 114.800 387.700 157.200 388.300 ;
        RECT 39.600 387.600 40.400 387.700 ;
        RECT 42.800 387.600 43.600 387.700 ;
        RECT 55.600 387.600 56.400 387.700 ;
        RECT 78.000 387.600 78.800 387.700 ;
        RECT 98.800 387.600 99.600 387.700 ;
        RECT 114.800 387.600 115.600 387.700 ;
        RECT 156.400 387.600 157.200 387.700 ;
        RECT 210.800 388.300 211.600 388.400 ;
        RECT 226.800 388.300 227.600 388.400 ;
        RECT 210.800 387.700 227.600 388.300 ;
        RECT 210.800 387.600 211.600 387.700 ;
        RECT 226.800 387.600 227.600 387.700 ;
        RECT 428.400 388.300 429.200 388.400 ;
        RECT 442.800 388.300 443.600 388.400 ;
        RECT 428.400 387.700 443.600 388.300 ;
        RECT 428.400 387.600 429.200 387.700 ;
        RECT 442.800 387.600 443.600 387.700 ;
        RECT 474.800 388.300 475.600 388.400 ;
        RECT 494.000 388.300 494.800 388.400 ;
        RECT 474.800 387.700 494.800 388.300 ;
        RECT 474.800 387.600 475.600 387.700 ;
        RECT 494.000 387.600 494.800 387.700 ;
        RECT 514.800 388.300 515.600 388.400 ;
        RECT 530.800 388.300 531.600 388.400 ;
        RECT 514.800 387.700 531.600 388.300 ;
        RECT 514.800 387.600 515.600 387.700 ;
        RECT 530.800 387.600 531.600 387.700 ;
        RECT 554.800 388.300 555.600 388.400 ;
        RECT 559.600 388.300 560.400 388.400 ;
        RECT 567.600 388.300 568.400 388.400 ;
        RECT 572.400 388.300 573.200 388.400 ;
        RECT 574.000 388.300 574.800 388.400 ;
        RECT 554.800 387.700 574.800 388.300 ;
        RECT 554.800 387.600 555.600 387.700 ;
        RECT 559.600 387.600 560.400 387.700 ;
        RECT 567.600 387.600 568.400 387.700 ;
        RECT 572.400 387.600 573.200 387.700 ;
        RECT 574.000 387.600 574.800 387.700 ;
        RECT 111.600 386.300 112.400 386.400 ;
        RECT 119.600 386.300 120.400 386.400 ;
        RECT 111.600 385.700 120.400 386.300 ;
        RECT 111.600 385.600 112.400 385.700 ;
        RECT 119.600 385.600 120.400 385.700 ;
        RECT 121.200 386.300 122.000 386.400 ;
        RECT 166.000 386.300 166.800 386.400 ;
        RECT 183.600 386.300 184.400 386.400 ;
        RECT 121.200 385.700 184.400 386.300 ;
        RECT 121.200 385.600 122.000 385.700 ;
        RECT 166.000 385.600 166.800 385.700 ;
        RECT 183.600 385.600 184.400 385.700 ;
        RECT 207.600 386.300 208.400 386.400 ;
        RECT 214.000 386.300 214.800 386.400 ;
        RECT 207.600 385.700 214.800 386.300 ;
        RECT 207.600 385.600 208.400 385.700 ;
        RECT 214.000 385.600 214.800 385.700 ;
        RECT 281.200 386.300 282.000 386.400 ;
        RECT 321.200 386.300 322.000 386.400 ;
        RECT 281.200 385.700 322.000 386.300 ;
        RECT 281.200 385.600 282.000 385.700 ;
        RECT 321.200 385.600 322.000 385.700 ;
        RECT 350.000 386.300 350.800 386.400 ;
        RECT 358.000 386.300 358.800 386.400 ;
        RECT 350.000 385.700 358.800 386.300 ;
        RECT 350.000 385.600 350.800 385.700 ;
        RECT 358.000 385.600 358.800 385.700 ;
        RECT 444.400 386.300 445.200 386.400 ;
        RECT 561.200 386.300 562.000 386.400 ;
        RECT 444.400 385.700 562.000 386.300 ;
        RECT 444.400 385.600 445.200 385.700 ;
        RECT 561.200 385.600 562.000 385.700 ;
        RECT 46.000 384.300 46.800 384.400 ;
        RECT 47.600 384.300 48.400 384.400 ;
        RECT 46.000 383.700 48.400 384.300 ;
        RECT 46.000 383.600 46.800 383.700 ;
        RECT 47.600 383.600 48.400 383.700 ;
        RECT 89.200 384.300 90.000 384.400 ;
        RECT 127.600 384.300 128.400 384.400 ;
        RECT 89.200 383.700 128.400 384.300 ;
        RECT 89.200 383.600 90.000 383.700 ;
        RECT 127.600 383.600 128.400 383.700 ;
        RECT 134.000 384.300 134.800 384.400 ;
        RECT 138.800 384.300 139.600 384.400 ;
        RECT 134.000 383.700 139.600 384.300 ;
        RECT 134.000 383.600 134.800 383.700 ;
        RECT 138.800 383.600 139.600 383.700 ;
        RECT 172.400 384.300 173.200 384.400 ;
        RECT 201.200 384.300 202.000 384.400 ;
        RECT 172.400 383.700 202.000 384.300 ;
        RECT 172.400 383.600 173.200 383.700 ;
        RECT 201.200 383.600 202.000 383.700 ;
        RECT 321.200 384.300 322.000 384.400 ;
        RECT 361.200 384.300 362.000 384.400 ;
        RECT 321.200 383.700 362.000 384.300 ;
        RECT 321.200 383.600 322.000 383.700 ;
        RECT 361.200 383.600 362.000 383.700 ;
        RECT 425.200 384.300 426.000 384.400 ;
        RECT 474.800 384.300 475.600 384.400 ;
        RECT 425.200 383.700 475.600 384.300 ;
        RECT 425.200 383.600 426.000 383.700 ;
        RECT 474.800 383.600 475.600 383.700 ;
        RECT 484.400 384.300 485.200 384.400 ;
        RECT 511.600 384.300 512.400 384.400 ;
        RECT 514.800 384.300 515.600 384.400 ;
        RECT 484.400 383.700 515.600 384.300 ;
        RECT 484.400 383.600 485.200 383.700 ;
        RECT 511.600 383.600 512.400 383.700 ;
        RECT 514.800 383.600 515.600 383.700 ;
        RECT 553.200 384.300 554.000 384.400 ;
        RECT 566.000 384.300 566.800 384.400 ;
        RECT 570.800 384.300 571.600 384.400 ;
        RECT 553.200 383.700 571.600 384.300 ;
        RECT 553.200 383.600 554.000 383.700 ;
        RECT 566.000 383.600 566.800 383.700 ;
        RECT 570.800 383.600 571.600 383.700 ;
        RECT 26.800 382.300 27.600 382.400 ;
        RECT 39.600 382.300 40.400 382.400 ;
        RECT 106.800 382.300 107.600 382.400 ;
        RECT 26.800 381.700 107.600 382.300 ;
        RECT 26.800 381.600 27.600 381.700 ;
        RECT 39.600 381.600 40.400 381.700 ;
        RECT 106.800 381.600 107.600 381.700 ;
        RECT 108.400 382.300 109.200 382.400 ;
        RECT 121.200 382.300 122.000 382.400 ;
        RECT 108.400 381.700 122.000 382.300 ;
        RECT 108.400 381.600 109.200 381.700 ;
        RECT 121.200 381.600 122.000 381.700 ;
        RECT 228.400 382.300 229.200 382.400 ;
        RECT 257.200 382.300 258.000 382.400 ;
        RECT 228.400 381.700 258.000 382.300 ;
        RECT 228.400 381.600 229.200 381.700 ;
        RECT 257.200 381.600 258.000 381.700 ;
        RECT 282.800 382.300 283.600 382.400 ;
        RECT 284.400 382.300 285.200 382.400 ;
        RECT 282.800 381.700 285.200 382.300 ;
        RECT 282.800 381.600 283.600 381.700 ;
        RECT 284.400 381.600 285.200 381.700 ;
        RECT 313.200 382.300 314.000 382.400 ;
        RECT 318.000 382.300 318.800 382.400 ;
        RECT 313.200 381.700 318.800 382.300 ;
        RECT 313.200 381.600 314.000 381.700 ;
        RECT 318.000 381.600 318.800 381.700 ;
        RECT 359.600 382.300 360.400 382.400 ;
        RECT 386.800 382.300 387.600 382.400 ;
        RECT 396.400 382.300 397.200 382.400 ;
        RECT 425.300 382.300 425.900 383.600 ;
        RECT 359.600 381.700 425.900 382.300 ;
        RECT 431.600 382.300 432.400 382.400 ;
        RECT 452.400 382.300 453.200 382.400 ;
        RECT 484.400 382.300 485.200 382.400 ;
        RECT 431.600 381.700 485.200 382.300 ;
        RECT 359.600 381.600 360.400 381.700 ;
        RECT 386.800 381.600 387.600 381.700 ;
        RECT 396.400 381.600 397.200 381.700 ;
        RECT 431.600 381.600 432.400 381.700 ;
        RECT 452.400 381.600 453.200 381.700 ;
        RECT 484.400 381.600 485.200 381.700 ;
        RECT 508.400 382.300 509.200 382.400 ;
        RECT 521.200 382.300 522.000 382.400 ;
        RECT 508.400 381.700 522.000 382.300 ;
        RECT 508.400 381.600 509.200 381.700 ;
        RECT 521.200 381.600 522.000 381.700 ;
        RECT 534.000 382.300 534.800 382.400 ;
        RECT 537.200 382.300 538.000 382.400 ;
        RECT 534.000 381.700 538.000 382.300 ;
        RECT 534.000 381.600 534.800 381.700 ;
        RECT 537.200 381.600 538.000 381.700 ;
        RECT 78.000 380.300 78.800 380.400 ;
        RECT 94.000 380.300 94.800 380.400 ;
        RECT 111.600 380.300 112.400 380.400 ;
        RECT 132.400 380.300 133.200 380.400 ;
        RECT 78.000 379.700 133.200 380.300 ;
        RECT 78.000 379.600 78.800 379.700 ;
        RECT 94.000 379.600 94.800 379.700 ;
        RECT 111.600 379.600 112.400 379.700 ;
        RECT 132.400 379.600 133.200 379.700 ;
        RECT 231.600 380.300 232.400 380.400 ;
        RECT 249.200 380.300 250.000 380.400 ;
        RECT 231.600 379.700 250.000 380.300 ;
        RECT 231.600 379.600 232.400 379.700 ;
        RECT 249.200 379.600 250.000 379.700 ;
        RECT 250.800 380.300 251.600 380.400 ;
        RECT 281.200 380.300 282.000 380.400 ;
        RECT 286.000 380.300 286.800 380.400 ;
        RECT 250.800 379.700 286.800 380.300 ;
        RECT 250.800 379.600 251.600 379.700 ;
        RECT 281.200 379.600 282.000 379.700 ;
        RECT 286.000 379.600 286.800 379.700 ;
        RECT 342.000 380.300 342.800 380.400 ;
        RECT 375.600 380.300 376.400 380.400 ;
        RECT 394.800 380.300 395.600 380.400 ;
        RECT 398.000 380.300 398.800 380.400 ;
        RECT 342.000 379.700 395.600 380.300 ;
        RECT 342.000 379.600 342.800 379.700 ;
        RECT 375.600 379.600 376.400 379.700 ;
        RECT 394.800 379.600 395.600 379.700 ;
        RECT 396.500 379.700 398.800 380.300 ;
        RECT 81.200 378.300 82.000 378.400 ;
        RECT 84.400 378.300 85.200 378.400 ;
        RECT 92.400 378.300 93.200 378.400 ;
        RECT 129.200 378.300 130.000 378.400 ;
        RECT 81.200 377.700 130.000 378.300 ;
        RECT 81.200 377.600 82.000 377.700 ;
        RECT 84.400 377.600 85.200 377.700 ;
        RECT 92.400 377.600 93.200 377.700 ;
        RECT 129.200 377.600 130.000 377.700 ;
        RECT 142.000 378.300 142.800 378.400 ;
        RECT 148.400 378.300 149.200 378.400 ;
        RECT 142.000 377.700 149.200 378.300 ;
        RECT 142.000 377.600 142.800 377.700 ;
        RECT 148.400 377.600 149.200 377.700 ;
        RECT 218.800 378.300 219.600 378.400 ;
        RECT 226.800 378.300 227.600 378.400 ;
        RECT 218.800 377.700 227.600 378.300 ;
        RECT 218.800 377.600 219.600 377.700 ;
        RECT 226.800 377.600 227.600 377.700 ;
        RECT 281.200 378.300 282.000 378.400 ;
        RECT 396.500 378.300 397.100 379.700 ;
        RECT 398.000 379.600 398.800 379.700 ;
        RECT 404.400 380.300 405.200 380.400 ;
        RECT 474.800 380.300 475.600 380.400 ;
        RECT 404.400 379.700 475.600 380.300 ;
        RECT 404.400 379.600 405.200 379.700 ;
        RECT 474.800 379.600 475.600 379.700 ;
        RECT 542.000 380.300 542.800 380.400 ;
        RECT 546.800 380.300 547.600 380.400 ;
        RECT 542.000 379.700 547.600 380.300 ;
        RECT 542.000 379.600 542.800 379.700 ;
        RECT 546.800 379.600 547.600 379.700 ;
        RECT 281.200 377.700 397.100 378.300 ;
        RECT 407.600 378.300 408.400 378.400 ;
        RECT 438.000 378.300 438.800 378.400 ;
        RECT 457.200 378.300 458.000 378.400 ;
        RECT 407.600 377.700 458.000 378.300 ;
        RECT 281.200 377.600 282.000 377.700 ;
        RECT 407.600 377.600 408.400 377.700 ;
        RECT 438.000 377.600 438.800 377.700 ;
        RECT 457.200 377.600 458.000 377.700 ;
        RECT 6.000 376.300 6.800 376.400 ;
        RECT 9.200 376.300 10.000 376.400 ;
        RECT 6.000 375.700 10.000 376.300 ;
        RECT 6.000 375.600 6.800 375.700 ;
        RECT 9.200 375.600 10.000 375.700 ;
        RECT 12.400 376.300 13.200 376.400 ;
        RECT 33.200 376.300 34.000 376.400 ;
        RECT 12.400 375.700 34.000 376.300 ;
        RECT 12.400 375.600 13.200 375.700 ;
        RECT 33.200 375.600 34.000 375.700 ;
        RECT 70.000 376.300 70.800 376.400 ;
        RECT 78.000 376.300 78.800 376.400 ;
        RECT 70.000 375.700 78.800 376.300 ;
        RECT 70.000 375.600 70.800 375.700 ;
        RECT 78.000 375.600 78.800 375.700 ;
        RECT 82.800 376.300 83.600 376.400 ;
        RECT 89.200 376.300 90.000 376.400 ;
        RECT 82.800 375.700 90.000 376.300 ;
        RECT 82.800 375.600 83.600 375.700 ;
        RECT 89.200 375.600 90.000 375.700 ;
        RECT 106.800 376.300 107.600 376.400 ;
        RECT 129.200 376.300 130.000 376.400 ;
        RECT 132.400 376.300 133.200 376.400 ;
        RECT 106.800 375.700 133.200 376.300 ;
        RECT 106.800 375.600 107.600 375.700 ;
        RECT 129.200 375.600 130.000 375.700 ;
        RECT 132.400 375.600 133.200 375.700 ;
        RECT 142.000 376.300 142.800 376.400 ;
        RECT 172.400 376.300 173.200 376.400 ;
        RECT 142.000 375.700 173.200 376.300 ;
        RECT 142.000 375.600 142.800 375.700 ;
        RECT 172.400 375.600 173.200 375.700 ;
        RECT 190.000 376.300 190.800 376.400 ;
        RECT 230.000 376.300 230.800 376.400 ;
        RECT 190.000 375.700 230.800 376.300 ;
        RECT 190.000 375.600 190.800 375.700 ;
        RECT 230.000 375.600 230.800 375.700 ;
        RECT 319.600 376.300 320.400 376.400 ;
        RECT 337.200 376.300 338.000 376.400 ;
        RECT 319.600 375.700 338.000 376.300 ;
        RECT 319.600 375.600 320.400 375.700 ;
        RECT 337.200 375.600 338.000 375.700 ;
        RECT 417.200 376.300 418.000 376.400 ;
        RECT 442.800 376.300 443.600 376.400 ;
        RECT 498.800 376.300 499.600 376.400 ;
        RECT 506.800 376.300 507.600 376.400 ;
        RECT 417.200 375.700 507.600 376.300 ;
        RECT 417.200 375.600 418.000 375.700 ;
        RECT 442.800 375.600 443.600 375.700 ;
        RECT 498.800 375.600 499.600 375.700 ;
        RECT 506.800 375.600 507.600 375.700 ;
        RECT 562.800 376.300 563.600 376.400 ;
        RECT 593.200 376.300 594.000 376.400 ;
        RECT 562.800 375.700 594.000 376.300 ;
        RECT 562.800 375.600 563.600 375.700 ;
        RECT 593.200 375.600 594.000 375.700 ;
        RECT 6.000 374.300 6.800 374.400 ;
        RECT 14.000 374.300 14.800 374.400 ;
        RECT 6.000 373.700 14.800 374.300 ;
        RECT 6.000 373.600 6.800 373.700 ;
        RECT 14.000 373.600 14.800 373.700 ;
        RECT 26.800 374.300 27.600 374.400 ;
        RECT 38.000 374.300 38.800 374.400 ;
        RECT 42.800 374.300 43.600 374.400 ;
        RECT 26.800 373.700 43.600 374.300 ;
        RECT 26.800 373.600 27.600 373.700 ;
        RECT 38.000 373.600 38.800 373.700 ;
        RECT 42.800 373.600 43.600 373.700 ;
        RECT 44.400 374.300 45.200 374.400 ;
        RECT 49.200 374.300 50.000 374.400 ;
        RECT 55.600 374.300 56.400 374.400 ;
        RECT 44.400 373.700 56.400 374.300 ;
        RECT 44.400 373.600 45.200 373.700 ;
        RECT 49.200 373.600 50.000 373.700 ;
        RECT 55.600 373.600 56.400 373.700 ;
        RECT 57.200 374.300 58.000 374.400 ;
        RECT 90.800 374.300 91.600 374.400 ;
        RECT 57.200 373.700 91.600 374.300 ;
        RECT 57.200 373.600 58.000 373.700 ;
        RECT 90.800 373.600 91.600 373.700 ;
        RECT 121.200 374.300 122.000 374.400 ;
        RECT 124.400 374.300 125.200 374.400 ;
        RECT 137.200 374.300 138.000 374.400 ;
        RECT 161.200 374.300 162.000 374.400 ;
        RECT 121.200 373.700 162.000 374.300 ;
        RECT 121.200 373.600 122.000 373.700 ;
        RECT 124.400 373.600 125.200 373.700 ;
        RECT 137.200 373.600 138.000 373.700 ;
        RECT 161.200 373.600 162.000 373.700 ;
        RECT 186.800 374.300 187.600 374.400 ;
        RECT 204.400 374.300 205.200 374.400 ;
        RECT 186.800 373.700 205.200 374.300 ;
        RECT 186.800 373.600 187.600 373.700 ;
        RECT 204.400 373.600 205.200 373.700 ;
        RECT 212.400 374.300 213.200 374.400 ;
        RECT 220.400 374.300 221.200 374.400 ;
        RECT 212.400 373.700 221.200 374.300 ;
        RECT 212.400 373.600 213.200 373.700 ;
        RECT 220.400 373.600 221.200 373.700 ;
        RECT 226.800 374.300 227.600 374.400 ;
        RECT 260.400 374.300 261.200 374.400 ;
        RECT 226.800 373.700 261.200 374.300 ;
        RECT 226.800 373.600 227.600 373.700 ;
        RECT 260.400 373.600 261.200 373.700 ;
        RECT 270.000 374.300 270.800 374.400 ;
        RECT 274.800 374.300 275.600 374.400 ;
        RECT 276.400 374.300 277.200 374.400 ;
        RECT 289.200 374.300 290.000 374.400 ;
        RECT 270.000 373.700 290.000 374.300 ;
        RECT 270.000 373.600 270.800 373.700 ;
        RECT 274.800 373.600 275.600 373.700 ;
        RECT 276.400 373.600 277.200 373.700 ;
        RECT 289.200 373.600 290.000 373.700 ;
        RECT 338.800 374.300 339.600 374.400 ;
        RECT 356.400 374.300 357.200 374.400 ;
        RECT 338.800 373.700 357.200 374.300 ;
        RECT 338.800 373.600 339.600 373.700 ;
        RECT 356.400 373.600 357.200 373.700 ;
        RECT 399.600 374.300 400.400 374.400 ;
        RECT 418.800 374.300 419.600 374.400 ;
        RECT 399.600 373.700 419.600 374.300 ;
        RECT 399.600 373.600 400.400 373.700 ;
        RECT 418.800 373.600 419.600 373.700 ;
        RECT 447.600 374.300 448.400 374.400 ;
        RECT 468.400 374.300 469.200 374.400 ;
        RECT 447.600 373.700 469.200 374.300 ;
        RECT 447.600 373.600 448.400 373.700 ;
        RECT 468.400 373.600 469.200 373.700 ;
        RECT 478.000 374.300 478.800 374.400 ;
        RECT 482.800 374.300 483.600 374.400 ;
        RECT 500.400 374.300 501.200 374.400 ;
        RECT 478.000 373.700 501.200 374.300 ;
        RECT 478.000 373.600 478.800 373.700 ;
        RECT 482.800 373.600 483.600 373.700 ;
        RECT 500.400 373.600 501.200 373.700 ;
        RECT 540.400 374.300 541.200 374.400 ;
        RECT 554.800 374.300 555.600 374.400 ;
        RECT 540.400 373.700 555.600 374.300 ;
        RECT 540.400 373.600 541.200 373.700 ;
        RECT 554.800 373.600 555.600 373.700 ;
        RECT 564.400 374.300 565.200 374.400 ;
        RECT 569.200 374.300 570.000 374.400 ;
        RECT 564.400 373.700 570.000 374.300 ;
        RECT 564.400 373.600 565.200 373.700 ;
        RECT 569.200 373.600 570.000 373.700 ;
        RECT 4.400 372.300 5.200 372.400 ;
        RECT 7.600 372.300 8.400 372.400 ;
        RECT 4.400 371.700 8.400 372.300 ;
        RECT 4.400 371.600 5.200 371.700 ;
        RECT 7.600 371.600 8.400 371.700 ;
        RECT 9.200 372.300 10.000 372.400 ;
        RECT 15.600 372.300 16.400 372.400 ;
        RECT 9.200 371.700 16.400 372.300 ;
        RECT 9.200 371.600 10.000 371.700 ;
        RECT 15.600 371.600 16.400 371.700 ;
        RECT 28.400 372.300 29.200 372.400 ;
        RECT 36.400 372.300 37.200 372.400 ;
        RECT 28.400 371.700 37.200 372.300 ;
        RECT 28.400 371.600 29.200 371.700 ;
        RECT 36.400 371.600 37.200 371.700 ;
        RECT 42.800 372.300 43.600 372.400 ;
        RECT 49.200 372.300 50.000 372.400 ;
        RECT 42.800 371.700 50.000 372.300 ;
        RECT 42.800 371.600 43.600 371.700 ;
        RECT 49.200 371.600 50.000 371.700 ;
        RECT 81.200 372.300 82.000 372.400 ;
        RECT 103.600 372.300 104.400 372.400 ;
        RECT 121.200 372.300 122.000 372.400 ;
        RECT 122.800 372.300 123.600 372.400 ;
        RECT 81.200 371.700 123.600 372.300 ;
        RECT 81.200 371.600 82.000 371.700 ;
        RECT 103.600 371.600 104.400 371.700 ;
        RECT 121.200 371.600 122.000 371.700 ;
        RECT 122.800 371.600 123.600 371.700 ;
        RECT 137.200 372.300 138.000 372.400 ;
        RECT 142.000 372.300 142.800 372.400 ;
        RECT 137.200 371.700 142.800 372.300 ;
        RECT 137.200 371.600 138.000 371.700 ;
        RECT 142.000 371.600 142.800 371.700 ;
        RECT 153.200 372.300 154.000 372.400 ;
        RECT 159.600 372.300 160.400 372.400 ;
        RECT 153.200 371.700 160.400 372.300 ;
        RECT 153.200 371.600 154.000 371.700 ;
        RECT 159.600 371.600 160.400 371.700 ;
        RECT 218.800 372.300 219.600 372.400 ;
        RECT 228.400 372.300 229.200 372.400 ;
        RECT 218.800 371.700 229.200 372.300 ;
        RECT 218.800 371.600 219.600 371.700 ;
        RECT 228.400 371.600 229.200 371.700 ;
        RECT 263.600 372.300 264.400 372.400 ;
        RECT 266.800 372.300 267.600 372.400 ;
        RECT 263.600 371.700 267.600 372.300 ;
        RECT 263.600 371.600 264.400 371.700 ;
        RECT 266.800 371.600 267.600 371.700 ;
        RECT 311.600 372.300 312.400 372.400 ;
        RECT 343.600 372.300 344.400 372.400 ;
        RECT 346.800 372.300 347.600 372.400 ;
        RECT 311.600 371.700 347.600 372.300 ;
        RECT 311.600 371.600 312.400 371.700 ;
        RECT 343.600 371.600 344.400 371.700 ;
        RECT 346.800 371.600 347.600 371.700 ;
        RECT 420.400 371.600 421.200 372.400 ;
        RECT 433.200 372.300 434.000 372.400 ;
        RECT 450.800 372.300 451.600 372.400 ;
        RECT 433.200 371.700 451.600 372.300 ;
        RECT 433.200 371.600 434.000 371.700 ;
        RECT 450.800 371.600 451.600 371.700 ;
        RECT 465.200 372.300 466.000 372.400 ;
        RECT 476.400 372.300 477.200 372.400 ;
        RECT 486.000 372.300 486.800 372.400 ;
        RECT 465.200 371.700 486.800 372.300 ;
        RECT 465.200 371.600 466.000 371.700 ;
        RECT 476.400 371.600 477.200 371.700 ;
        RECT 486.000 371.600 486.800 371.700 ;
        RECT 558.000 372.300 558.800 372.400 ;
        RECT 577.200 372.300 578.000 372.400 ;
        RECT 582.000 372.300 582.800 372.400 ;
        RECT 558.000 371.700 582.800 372.300 ;
        RECT 558.000 371.600 558.800 371.700 ;
        RECT 577.200 371.600 578.000 371.700 ;
        RECT 582.000 371.600 582.800 371.700 ;
        RECT 590.000 372.300 590.800 372.400 ;
        RECT 593.200 372.300 594.000 372.400 ;
        RECT 590.000 371.700 594.000 372.300 ;
        RECT 590.000 371.600 590.800 371.700 ;
        RECT 593.200 371.600 594.000 371.700 ;
        RECT 33.200 370.300 34.000 370.400 ;
        RECT 34.800 370.300 35.600 370.400 ;
        RECT 46.000 370.300 46.800 370.400 ;
        RECT 33.200 369.700 46.800 370.300 ;
        RECT 33.200 369.600 34.000 369.700 ;
        RECT 34.800 369.600 35.600 369.700 ;
        RECT 46.000 369.600 46.800 369.700 ;
        RECT 58.800 370.300 59.600 370.400 ;
        RECT 73.200 370.300 74.000 370.400 ;
        RECT 78.000 370.300 78.800 370.400 ;
        RECT 58.800 369.700 78.800 370.300 ;
        RECT 58.800 369.600 59.600 369.700 ;
        RECT 73.200 369.600 74.000 369.700 ;
        RECT 78.000 369.600 78.800 369.700 ;
        RECT 89.200 370.300 90.000 370.400 ;
        RECT 102.000 370.300 102.800 370.400 ;
        RECT 89.200 369.700 102.800 370.300 ;
        RECT 122.900 370.300 123.500 371.600 ;
        RECT 138.800 370.300 139.600 370.400 ;
        RECT 122.900 369.700 139.600 370.300 ;
        RECT 89.200 369.600 90.000 369.700 ;
        RECT 102.000 369.600 102.800 369.700 ;
        RECT 138.800 369.600 139.600 369.700 ;
        RECT 206.000 370.300 206.800 370.400 ;
        RECT 212.400 370.300 213.200 370.400 ;
        RECT 238.000 370.300 238.800 370.400 ;
        RECT 206.000 369.700 238.800 370.300 ;
        RECT 206.000 369.600 206.800 369.700 ;
        RECT 212.400 369.600 213.200 369.700 ;
        RECT 238.000 369.600 238.800 369.700 ;
        RECT 270.000 370.300 270.800 370.400 ;
        RECT 308.400 370.300 309.200 370.400 ;
        RECT 321.200 370.300 322.000 370.400 ;
        RECT 330.800 370.300 331.600 370.400 ;
        RECT 270.000 369.700 331.600 370.300 ;
        RECT 270.000 369.600 270.800 369.700 ;
        RECT 308.400 369.600 309.200 369.700 ;
        RECT 321.200 369.600 322.000 369.700 ;
        RECT 330.800 369.600 331.600 369.700 ;
        RECT 378.800 370.300 379.600 370.400 ;
        RECT 380.400 370.300 381.200 370.400 ;
        RECT 423.600 370.300 424.400 370.400 ;
        RECT 378.800 369.700 424.400 370.300 ;
        RECT 378.800 369.600 379.600 369.700 ;
        RECT 380.400 369.600 381.200 369.700 ;
        RECT 423.600 369.600 424.400 369.700 ;
        RECT 438.000 370.300 438.800 370.400 ;
        RECT 449.200 370.300 450.000 370.400 ;
        RECT 438.000 369.700 450.000 370.300 ;
        RECT 438.000 369.600 438.800 369.700 ;
        RECT 449.200 369.600 450.000 369.700 ;
        RECT 31.600 368.300 32.400 368.400 ;
        RECT 34.800 368.300 35.600 368.400 ;
        RECT 31.600 367.700 35.600 368.300 ;
        RECT 31.600 367.600 32.400 367.700 ;
        RECT 34.800 367.600 35.600 367.700 ;
        RECT 78.000 368.300 78.800 368.400 ;
        RECT 100.400 368.300 101.200 368.400 ;
        RECT 78.000 367.700 101.200 368.300 ;
        RECT 78.000 367.600 78.800 367.700 ;
        RECT 100.400 367.600 101.200 367.700 ;
        RECT 132.400 368.300 133.200 368.400 ;
        RECT 145.200 368.300 146.000 368.400 ;
        RECT 132.400 367.700 146.000 368.300 ;
        RECT 132.400 367.600 133.200 367.700 ;
        RECT 145.200 367.600 146.000 367.700 ;
        RECT 66.800 366.300 67.600 366.400 ;
        RECT 90.800 366.300 91.600 366.400 ;
        RECT 130.800 366.300 131.600 366.400 ;
        RECT 143.600 366.300 144.400 366.400 ;
        RECT 66.800 365.700 144.400 366.300 ;
        RECT 66.800 365.600 67.600 365.700 ;
        RECT 90.800 365.600 91.600 365.700 ;
        RECT 130.800 365.600 131.600 365.700 ;
        RECT 143.600 365.600 144.400 365.700 ;
        RECT 244.400 366.300 245.200 366.400 ;
        RECT 310.000 366.300 310.800 366.400 ;
        RECT 244.400 365.700 310.800 366.300 ;
        RECT 244.400 365.600 245.200 365.700 ;
        RECT 310.000 365.600 310.800 365.700 ;
        RECT 505.200 366.300 506.000 366.400 ;
        RECT 511.600 366.300 512.400 366.400 ;
        RECT 551.600 366.300 552.400 366.400 ;
        RECT 554.800 366.300 555.600 366.400 ;
        RECT 505.200 365.700 555.600 366.300 ;
        RECT 505.200 365.600 506.000 365.700 ;
        RECT 511.600 365.600 512.400 365.700 ;
        RECT 551.600 365.600 552.400 365.700 ;
        RECT 554.800 365.600 555.600 365.700 ;
        RECT 63.600 364.300 64.400 364.400 ;
        RECT 76.400 364.300 77.200 364.400 ;
        RECT 90.800 364.300 91.600 364.400 ;
        RECT 63.600 363.700 91.600 364.300 ;
        RECT 63.600 363.600 64.400 363.700 ;
        RECT 76.400 363.600 77.200 363.700 ;
        RECT 90.800 363.600 91.600 363.700 ;
        RECT 126.000 364.300 126.800 364.400 ;
        RECT 142.000 364.300 142.800 364.400 ;
        RECT 151.600 364.300 152.400 364.400 ;
        RECT 126.000 363.700 152.400 364.300 ;
        RECT 126.000 363.600 126.800 363.700 ;
        RECT 142.000 363.600 142.800 363.700 ;
        RECT 151.600 363.600 152.400 363.700 ;
        RECT 20.400 362.300 21.200 362.400 ;
        RECT 42.800 362.300 43.600 362.400 ;
        RECT 20.400 361.700 43.600 362.300 ;
        RECT 20.400 361.600 21.200 361.700 ;
        RECT 42.800 361.600 43.600 361.700 ;
        RECT 198.000 362.300 198.800 362.400 ;
        RECT 202.800 362.300 203.600 362.400 ;
        RECT 198.000 361.700 203.600 362.300 ;
        RECT 198.000 361.600 198.800 361.700 ;
        RECT 202.800 361.600 203.600 361.700 ;
        RECT 218.800 362.300 219.600 362.400 ;
        RECT 222.000 362.300 222.800 362.400 ;
        RECT 218.800 361.700 222.800 362.300 ;
        RECT 218.800 361.600 219.600 361.700 ;
        RECT 222.000 361.600 222.800 361.700 ;
        RECT 538.800 362.300 539.600 362.400 ;
        RECT 574.000 362.300 574.800 362.400 ;
        RECT 538.800 361.700 574.800 362.300 ;
        RECT 538.800 361.600 539.600 361.700 ;
        RECT 574.000 361.600 574.800 361.700 ;
        RECT 6.000 360.300 6.800 360.400 ;
        RECT 9.200 360.300 10.000 360.400 ;
        RECT 6.000 359.700 10.000 360.300 ;
        RECT 6.000 359.600 6.800 359.700 ;
        RECT 9.200 359.600 10.000 359.700 ;
        RECT 191.600 360.300 192.400 360.400 ;
        RECT 210.800 360.300 211.600 360.400 ;
        RECT 191.600 359.700 211.600 360.300 ;
        RECT 191.600 359.600 192.400 359.700 ;
        RECT 210.800 359.600 211.600 359.700 ;
        RECT 234.800 360.300 235.600 360.400 ;
        RECT 241.200 360.300 242.000 360.400 ;
        RECT 234.800 359.700 242.000 360.300 ;
        RECT 234.800 359.600 235.600 359.700 ;
        RECT 241.200 359.600 242.000 359.700 ;
        RECT 367.600 360.300 368.400 360.400 ;
        RECT 438.000 360.300 438.800 360.400 ;
        RECT 367.600 359.700 438.800 360.300 ;
        RECT 367.600 359.600 368.400 359.700 ;
        RECT 438.000 359.600 438.800 359.700 ;
        RECT 479.600 360.300 480.400 360.400 ;
        RECT 482.800 360.300 483.600 360.400 ;
        RECT 479.600 359.700 483.600 360.300 ;
        RECT 479.600 359.600 480.400 359.700 ;
        RECT 482.800 359.600 483.600 359.700 ;
        RECT 532.400 360.300 533.200 360.400 ;
        RECT 554.800 360.300 555.600 360.400 ;
        RECT 532.400 359.700 555.600 360.300 ;
        RECT 532.400 359.600 533.200 359.700 ;
        RECT 554.800 359.600 555.600 359.700 ;
        RECT 9.200 358.300 10.000 358.400 ;
        RECT 28.400 358.300 29.200 358.400 ;
        RECT 9.200 357.700 29.200 358.300 ;
        RECT 9.200 357.600 10.000 357.700 ;
        RECT 28.400 357.600 29.200 357.700 ;
        RECT 119.600 358.300 120.400 358.400 ;
        RECT 129.200 358.300 130.000 358.400 ;
        RECT 119.600 357.700 130.000 358.300 ;
        RECT 119.600 357.600 120.400 357.700 ;
        RECT 129.200 357.600 130.000 357.700 ;
        RECT 153.200 358.300 154.000 358.400 ;
        RECT 156.400 358.300 157.200 358.400 ;
        RECT 153.200 357.700 157.200 358.300 ;
        RECT 153.200 357.600 154.000 357.700 ;
        RECT 156.400 357.600 157.200 357.700 ;
        RECT 210.800 358.300 211.600 358.400 ;
        RECT 220.400 358.300 221.200 358.400 ;
        RECT 210.800 357.700 221.200 358.300 ;
        RECT 210.800 357.600 211.600 357.700 ;
        RECT 220.400 357.600 221.200 357.700 ;
        RECT 266.800 358.300 267.600 358.400 ;
        RECT 281.200 358.300 282.000 358.400 ;
        RECT 266.800 357.700 282.000 358.300 ;
        RECT 266.800 357.600 267.600 357.700 ;
        RECT 281.200 357.600 282.000 357.700 ;
        RECT 542.000 357.600 542.800 358.400 ;
        RECT 538.800 356.300 539.600 356.400 ;
        RECT 551.600 356.300 552.400 356.400 ;
        RECT 538.800 355.700 552.400 356.300 ;
        RECT 538.800 355.600 539.600 355.700 ;
        RECT 551.600 355.600 552.400 355.700 ;
        RECT 55.600 354.300 56.400 354.400 ;
        RECT 94.000 354.300 94.800 354.400 ;
        RECT 55.600 353.700 94.800 354.300 ;
        RECT 55.600 353.600 56.400 353.700 ;
        RECT 94.000 353.600 94.800 353.700 ;
        RECT 97.200 354.300 98.000 354.400 ;
        RECT 134.000 354.300 134.800 354.400 ;
        RECT 146.800 354.300 147.600 354.400 ;
        RECT 97.200 353.700 147.600 354.300 ;
        RECT 97.200 353.600 98.000 353.700 ;
        RECT 134.000 353.600 134.800 353.700 ;
        RECT 146.800 353.600 147.600 353.700 ;
        RECT 161.200 354.300 162.000 354.400 ;
        RECT 393.200 354.300 394.000 354.400 ;
        RECT 161.200 353.700 394.000 354.300 ;
        RECT 161.200 353.600 162.000 353.700 ;
        RECT 393.200 353.600 394.000 353.700 ;
        RECT 490.800 354.300 491.600 354.400 ;
        RECT 532.400 354.300 533.200 354.400 ;
        RECT 490.800 353.700 533.200 354.300 ;
        RECT 490.800 353.600 491.600 353.700 ;
        RECT 532.400 353.600 533.200 353.700 ;
        RECT 534.000 354.300 534.800 354.400 ;
        RECT 559.600 354.300 560.400 354.400 ;
        RECT 534.000 353.700 560.400 354.300 ;
        RECT 534.000 353.600 534.800 353.700 ;
        RECT 559.600 353.600 560.400 353.700 ;
        RECT 42.800 352.300 43.600 352.400 ;
        RECT 81.200 352.300 82.000 352.400 ;
        RECT 42.800 351.700 82.000 352.300 ;
        RECT 42.800 351.600 43.600 351.700 ;
        RECT 81.200 351.600 82.000 351.700 ;
        RECT 90.800 352.300 91.600 352.400 ;
        RECT 105.200 352.300 106.000 352.400 ;
        RECT 90.800 351.700 106.000 352.300 ;
        RECT 90.800 351.600 91.600 351.700 ;
        RECT 105.200 351.600 106.000 351.700 ;
        RECT 113.200 352.300 114.000 352.400 ;
        RECT 116.400 352.300 117.200 352.400 ;
        RECT 119.600 352.300 120.400 352.400 ;
        RECT 113.200 351.700 120.400 352.300 ;
        RECT 113.200 351.600 114.000 351.700 ;
        RECT 116.400 351.600 117.200 351.700 ;
        RECT 119.600 351.600 120.400 351.700 ;
        RECT 122.800 352.300 123.600 352.400 ;
        RECT 126.000 352.300 126.800 352.400 ;
        RECT 122.800 351.700 126.800 352.300 ;
        RECT 122.800 351.600 123.600 351.700 ;
        RECT 126.000 351.600 126.800 351.700 ;
        RECT 258.800 352.300 259.600 352.400 ;
        RECT 289.200 352.300 290.000 352.400 ;
        RECT 258.800 351.700 290.000 352.300 ;
        RECT 258.800 351.600 259.600 351.700 ;
        RECT 289.200 351.600 290.000 351.700 ;
        RECT 394.800 352.300 395.600 352.400 ;
        RECT 401.200 352.300 402.000 352.400 ;
        RECT 394.800 351.700 402.000 352.300 ;
        RECT 394.800 351.600 395.600 351.700 ;
        RECT 401.200 351.600 402.000 351.700 ;
        RECT 407.600 352.300 408.400 352.400 ;
        RECT 412.400 352.300 413.200 352.400 ;
        RECT 434.800 352.300 435.600 352.400 ;
        RECT 446.000 352.300 446.800 352.400 ;
        RECT 407.600 351.700 446.800 352.300 ;
        RECT 407.600 351.600 408.400 351.700 ;
        RECT 412.400 351.600 413.200 351.700 ;
        RECT 434.800 351.600 435.600 351.700 ;
        RECT 446.000 351.600 446.800 351.700 ;
        RECT 521.200 352.300 522.000 352.400 ;
        RECT 540.400 352.300 541.200 352.400 ;
        RECT 521.200 351.700 541.200 352.300 ;
        RECT 521.200 351.600 522.000 351.700 ;
        RECT 540.400 351.600 541.200 351.700 ;
        RECT 558.000 352.300 558.800 352.400 ;
        RECT 561.200 352.300 562.000 352.400 ;
        RECT 558.000 351.700 562.000 352.300 ;
        RECT 558.000 351.600 558.800 351.700 ;
        RECT 561.200 351.600 562.000 351.700 ;
        RECT 103.600 350.300 104.400 350.400 ;
        RECT 127.600 350.300 128.400 350.400 ;
        RECT 132.400 350.300 133.200 350.400 ;
        RECT 103.600 349.700 133.200 350.300 ;
        RECT 103.600 349.600 104.400 349.700 ;
        RECT 127.600 349.600 128.400 349.700 ;
        RECT 132.400 349.600 133.200 349.700 ;
        RECT 158.000 350.300 158.800 350.400 ;
        RECT 170.800 350.300 171.600 350.400 ;
        RECT 158.000 349.700 171.600 350.300 ;
        RECT 158.000 349.600 158.800 349.700 ;
        RECT 170.800 349.600 171.600 349.700 ;
        RECT 202.800 350.300 203.600 350.400 ;
        RECT 212.400 350.300 213.200 350.400 ;
        RECT 202.800 349.700 213.200 350.300 ;
        RECT 202.800 349.600 203.600 349.700 ;
        RECT 212.400 349.600 213.200 349.700 ;
        RECT 228.400 349.600 229.200 350.400 ;
        RECT 233.200 350.300 234.000 350.400 ;
        RECT 238.000 350.300 238.800 350.400 ;
        RECT 233.200 349.700 238.800 350.300 ;
        RECT 233.200 349.600 234.000 349.700 ;
        RECT 238.000 349.600 238.800 349.700 ;
        RECT 286.000 350.300 286.800 350.400 ;
        RECT 302.000 350.300 302.800 350.400 ;
        RECT 286.000 349.700 302.800 350.300 ;
        RECT 286.000 349.600 286.800 349.700 ;
        RECT 302.000 349.600 302.800 349.700 ;
        RECT 318.000 350.300 318.800 350.400 ;
        RECT 346.800 350.300 347.600 350.400 ;
        RECT 388.400 350.300 389.200 350.400 ;
        RECT 318.000 349.700 337.900 350.300 ;
        RECT 318.000 349.600 318.800 349.700 ;
        RECT 337.300 348.400 337.900 349.700 ;
        RECT 346.800 349.700 389.200 350.300 ;
        RECT 346.800 349.600 347.600 349.700 ;
        RECT 388.400 349.600 389.200 349.700 ;
        RECT 390.000 350.300 390.800 350.400 ;
        RECT 399.600 350.300 400.400 350.400 ;
        RECT 390.000 349.700 400.400 350.300 ;
        RECT 390.000 349.600 390.800 349.700 ;
        RECT 399.600 349.600 400.400 349.700 ;
        RECT 404.400 350.300 405.200 350.400 ;
        RECT 409.200 350.300 410.000 350.400 ;
        RECT 404.400 349.700 410.000 350.300 ;
        RECT 404.400 349.600 405.200 349.700 ;
        RECT 409.200 349.600 410.000 349.700 ;
        RECT 489.200 350.300 490.000 350.400 ;
        RECT 495.600 350.300 496.400 350.400 ;
        RECT 489.200 349.700 496.400 350.300 ;
        RECT 489.200 349.600 490.000 349.700 ;
        RECT 495.600 349.600 496.400 349.700 ;
        RECT 518.000 350.300 518.800 350.400 ;
        RECT 567.600 350.300 568.400 350.400 ;
        RECT 518.000 349.700 568.400 350.300 ;
        RECT 518.000 349.600 518.800 349.700 ;
        RECT 567.600 349.600 568.400 349.700 ;
        RECT 598.000 350.300 598.800 350.400 ;
        RECT 604.400 350.300 605.200 350.400 ;
        RECT 598.000 349.700 605.200 350.300 ;
        RECT 598.000 349.600 598.800 349.700 ;
        RECT 604.400 349.600 605.200 349.700 ;
        RECT 15.600 348.300 16.400 348.400 ;
        RECT 23.600 348.300 24.400 348.400 ;
        RECT 15.600 347.700 24.400 348.300 ;
        RECT 15.600 347.600 16.400 347.700 ;
        RECT 23.600 347.600 24.400 347.700 ;
        RECT 34.800 348.300 35.600 348.400 ;
        RECT 50.800 348.300 51.600 348.400 ;
        RECT 34.800 347.700 51.600 348.300 ;
        RECT 34.800 347.600 35.600 347.700 ;
        RECT 50.800 347.600 51.600 347.700 ;
        RECT 55.600 348.300 56.400 348.400 ;
        RECT 86.000 348.300 86.800 348.400 ;
        RECT 92.400 348.300 93.200 348.400 ;
        RECT 98.800 348.300 99.600 348.400 ;
        RECT 55.600 347.700 99.600 348.300 ;
        RECT 55.600 347.600 56.400 347.700 ;
        RECT 86.000 347.600 86.800 347.700 ;
        RECT 92.400 347.600 93.200 347.700 ;
        RECT 98.800 347.600 99.600 347.700 ;
        RECT 113.200 348.300 114.000 348.400 ;
        RECT 130.800 348.300 131.600 348.400 ;
        RECT 113.200 347.700 131.600 348.300 ;
        RECT 113.200 347.600 114.000 347.700 ;
        RECT 130.800 347.600 131.600 347.700 ;
        RECT 247.600 348.300 248.400 348.400 ;
        RECT 273.200 348.300 274.000 348.400 ;
        RECT 247.600 347.700 274.000 348.300 ;
        RECT 247.600 347.600 248.400 347.700 ;
        RECT 273.200 347.600 274.000 347.700 ;
        RECT 298.800 348.300 299.600 348.400 ;
        RECT 329.200 348.300 330.000 348.400 ;
        RECT 298.800 347.700 330.000 348.300 ;
        RECT 298.800 347.600 299.600 347.700 ;
        RECT 329.200 347.600 330.000 347.700 ;
        RECT 337.200 347.600 338.000 348.400 ;
        RECT 374.000 348.300 374.800 348.400 ;
        RECT 404.400 348.300 405.200 348.400 ;
        RECT 409.200 348.300 410.000 348.400 ;
        RECT 374.000 347.700 410.000 348.300 ;
        RECT 374.000 347.600 374.800 347.700 ;
        RECT 404.400 347.600 405.200 347.700 ;
        RECT 409.200 347.600 410.000 347.700 ;
        RECT 460.400 348.300 461.200 348.400 ;
        RECT 506.800 348.300 507.600 348.400 ;
        RECT 460.400 347.700 507.600 348.300 ;
        RECT 460.400 347.600 461.200 347.700 ;
        RECT 506.800 347.600 507.600 347.700 ;
        RECT 543.600 348.300 544.400 348.400 ;
        RECT 559.600 348.300 560.400 348.400 ;
        RECT 566.000 348.300 566.800 348.400 ;
        RECT 543.600 347.700 566.800 348.300 ;
        RECT 543.600 347.600 544.400 347.700 ;
        RECT 559.600 347.600 560.400 347.700 ;
        RECT 566.000 347.600 566.800 347.700 ;
        RECT 590.000 348.300 590.800 348.400 ;
        RECT 601.200 348.300 602.000 348.400 ;
        RECT 606.000 348.300 606.800 348.400 ;
        RECT 590.000 347.700 606.800 348.300 ;
        RECT 590.000 347.600 590.800 347.700 ;
        RECT 601.200 347.600 602.000 347.700 ;
        RECT 606.000 347.600 606.800 347.700 ;
        RECT 17.200 346.300 18.000 346.400 ;
        RECT 26.800 346.300 27.600 346.400 ;
        RECT 17.200 345.700 27.600 346.300 ;
        RECT 17.200 345.600 18.000 345.700 ;
        RECT 26.800 345.600 27.600 345.700 ;
        RECT 52.400 346.300 53.200 346.400 ;
        RECT 236.400 346.300 237.200 346.400 ;
        RECT 327.600 346.300 328.400 346.400 ;
        RECT 345.200 346.300 346.000 346.400 ;
        RECT 52.400 345.700 346.000 346.300 ;
        RECT 52.400 345.600 53.200 345.700 ;
        RECT 236.400 345.600 237.200 345.700 ;
        RECT 327.600 345.600 328.400 345.700 ;
        RECT 345.200 345.600 346.000 345.700 ;
        RECT 351.600 346.300 352.400 346.400 ;
        RECT 378.800 346.300 379.600 346.400 ;
        RECT 351.600 345.700 379.600 346.300 ;
        RECT 351.600 345.600 352.400 345.700 ;
        RECT 378.800 345.600 379.600 345.700 ;
        RECT 401.200 346.300 402.000 346.400 ;
        RECT 407.600 346.300 408.400 346.400 ;
        RECT 415.600 346.300 416.400 346.400 ;
        RECT 401.200 345.700 416.400 346.300 ;
        RECT 401.200 345.600 402.000 345.700 ;
        RECT 407.600 345.600 408.400 345.700 ;
        RECT 415.600 345.600 416.400 345.700 ;
        RECT 476.400 346.300 477.200 346.400 ;
        RECT 510.000 346.300 510.800 346.400 ;
        RECT 522.800 346.300 523.600 346.400 ;
        RECT 476.400 345.700 523.600 346.300 ;
        RECT 476.400 345.600 477.200 345.700 ;
        RECT 510.000 345.600 510.800 345.700 ;
        RECT 522.800 345.600 523.600 345.700 ;
        RECT 529.200 345.600 530.000 346.400 ;
        RECT 129.200 344.300 130.000 344.400 ;
        RECT 135.600 344.300 136.400 344.400 ;
        RECT 129.200 343.700 136.400 344.300 ;
        RECT 129.200 343.600 130.000 343.700 ;
        RECT 135.600 343.600 136.400 343.700 ;
        RECT 174.000 344.300 174.800 344.400 ;
        RECT 196.400 344.300 197.200 344.400 ;
        RECT 174.000 343.700 197.200 344.300 ;
        RECT 174.000 343.600 174.800 343.700 ;
        RECT 196.400 343.600 197.200 343.700 ;
        RECT 321.200 344.300 322.000 344.400 ;
        RECT 326.000 344.300 326.800 344.400 ;
        RECT 321.200 343.700 326.800 344.300 ;
        RECT 321.200 343.600 322.000 343.700 ;
        RECT 326.000 343.600 326.800 343.700 ;
        RECT 370.800 344.300 371.600 344.400 ;
        RECT 449.200 344.300 450.000 344.400 ;
        RECT 370.800 343.700 450.000 344.300 ;
        RECT 370.800 343.600 371.600 343.700 ;
        RECT 449.200 343.600 450.000 343.700 ;
        RECT 9.200 342.300 10.000 342.400 ;
        RECT 14.000 342.300 14.800 342.400 ;
        RECT 9.200 341.700 14.800 342.300 ;
        RECT 9.200 341.600 10.000 341.700 ;
        RECT 14.000 341.600 14.800 341.700 ;
        RECT 60.400 342.300 61.200 342.400 ;
        RECT 81.200 342.300 82.000 342.400 ;
        RECT 94.000 342.300 94.800 342.400 ;
        RECT 60.400 341.700 94.800 342.300 ;
        RECT 60.400 341.600 61.200 341.700 ;
        RECT 81.200 341.600 82.000 341.700 ;
        RECT 94.000 341.600 94.800 341.700 ;
        RECT 119.600 342.300 120.400 342.400 ;
        RECT 124.400 342.300 125.200 342.400 ;
        RECT 119.600 341.700 125.200 342.300 ;
        RECT 119.600 341.600 120.400 341.700 ;
        RECT 124.400 341.600 125.200 341.700 ;
        RECT 169.200 342.300 170.000 342.400 ;
        RECT 174.000 342.300 174.800 342.400 ;
        RECT 169.200 341.700 174.800 342.300 ;
        RECT 169.200 341.600 170.000 341.700 ;
        RECT 174.000 341.600 174.800 341.700 ;
        RECT 194.800 342.300 195.600 342.400 ;
        RECT 210.800 342.300 211.600 342.400 ;
        RECT 194.800 341.700 211.600 342.300 ;
        RECT 194.800 341.600 195.600 341.700 ;
        RECT 210.800 341.600 211.600 341.700 ;
        RECT 226.800 342.300 227.600 342.400 ;
        RECT 231.600 342.300 232.400 342.400 ;
        RECT 238.000 342.300 238.800 342.400 ;
        RECT 226.800 341.700 238.800 342.300 ;
        RECT 226.800 341.600 227.600 341.700 ;
        RECT 231.600 341.600 232.400 341.700 ;
        RECT 238.000 341.600 238.800 341.700 ;
        RECT 324.400 342.300 325.200 342.400 ;
        RECT 335.600 342.300 336.400 342.400 ;
        RECT 324.400 341.700 336.400 342.300 ;
        RECT 324.400 341.600 325.200 341.700 ;
        RECT 335.600 341.600 336.400 341.700 ;
        RECT 410.800 341.600 411.600 342.400 ;
        RECT 414.000 342.300 414.800 342.400 ;
        RECT 431.600 342.300 432.400 342.400 ;
        RECT 414.000 341.700 432.400 342.300 ;
        RECT 414.000 341.600 414.800 341.700 ;
        RECT 431.600 341.600 432.400 341.700 ;
        RECT 526.000 342.300 526.800 342.400 ;
        RECT 585.200 342.300 586.000 342.400 ;
        RECT 526.000 341.700 586.000 342.300 ;
        RECT 526.000 341.600 526.800 341.700 ;
        RECT 585.200 341.600 586.000 341.700 ;
        RECT 7.600 340.300 8.400 340.400 ;
        RECT 12.400 340.300 13.200 340.400 ;
        RECT 7.600 339.700 13.200 340.300 ;
        RECT 7.600 339.600 8.400 339.700 ;
        RECT 12.400 339.600 13.200 339.700 ;
        RECT 90.800 340.300 91.600 340.400 ;
        RECT 145.200 340.300 146.000 340.400 ;
        RECT 90.800 339.700 146.000 340.300 ;
        RECT 90.800 339.600 91.600 339.700 ;
        RECT 145.200 339.600 146.000 339.700 ;
        RECT 172.400 340.300 173.200 340.400 ;
        RECT 196.400 340.300 197.200 340.400 ;
        RECT 172.400 339.700 197.200 340.300 ;
        RECT 172.400 339.600 173.200 339.700 ;
        RECT 196.400 339.600 197.200 339.700 ;
        RECT 250.800 340.300 251.600 340.400 ;
        RECT 257.200 340.300 258.000 340.400 ;
        RECT 250.800 339.700 258.000 340.300 ;
        RECT 250.800 339.600 251.600 339.700 ;
        RECT 257.200 339.600 258.000 339.700 ;
        RECT 270.000 340.300 270.800 340.400 ;
        RECT 271.600 340.300 272.400 340.400 ;
        RECT 270.000 339.700 272.400 340.300 ;
        RECT 270.000 339.600 270.800 339.700 ;
        RECT 271.600 339.600 272.400 339.700 ;
        RECT 292.400 340.300 293.200 340.400 ;
        RECT 294.000 340.300 294.800 340.400 ;
        RECT 292.400 339.700 294.800 340.300 ;
        RECT 292.400 339.600 293.200 339.700 ;
        RECT 294.000 339.600 294.800 339.700 ;
        RECT 343.600 340.300 344.400 340.400 ;
        RECT 382.000 340.300 382.800 340.400 ;
        RECT 343.600 339.700 382.800 340.300 ;
        RECT 343.600 339.600 344.400 339.700 ;
        RECT 382.000 339.600 382.800 339.700 ;
        RECT 402.800 340.300 403.600 340.400 ;
        RECT 452.400 340.300 453.200 340.400 ;
        RECT 462.000 340.300 462.800 340.400 ;
        RECT 402.800 339.700 462.800 340.300 ;
        RECT 402.800 339.600 403.600 339.700 ;
        RECT 452.400 339.600 453.200 339.700 ;
        RECT 462.000 339.600 462.800 339.700 ;
        RECT 526.000 340.300 526.800 340.400 ;
        RECT 530.800 340.300 531.600 340.400 ;
        RECT 526.000 339.700 531.600 340.300 ;
        RECT 526.000 339.600 526.800 339.700 ;
        RECT 530.800 339.600 531.600 339.700 ;
        RECT 292.400 338.300 293.200 338.400 ;
        RECT 332.400 338.300 333.200 338.400 ;
        RECT 292.400 337.700 333.200 338.300 ;
        RECT 292.400 337.600 293.200 337.700 ;
        RECT 332.400 337.600 333.200 337.700 ;
        RECT 353.200 338.300 354.000 338.400 ;
        RECT 414.000 338.300 414.800 338.400 ;
        RECT 353.200 337.700 414.800 338.300 ;
        RECT 353.200 337.600 354.000 337.700 ;
        RECT 414.000 337.600 414.800 337.700 ;
        RECT 431.600 338.300 432.400 338.400 ;
        RECT 434.800 338.300 435.600 338.400 ;
        RECT 431.600 337.700 435.600 338.300 ;
        RECT 431.600 337.600 432.400 337.700 ;
        RECT 434.800 337.600 435.600 337.700 ;
        RECT 564.400 338.300 565.200 338.400 ;
        RECT 572.400 338.300 573.200 338.400 ;
        RECT 564.400 337.700 573.200 338.300 ;
        RECT 564.400 337.600 565.200 337.700 ;
        RECT 572.400 337.600 573.200 337.700 ;
        RECT 594.800 338.300 595.600 338.400 ;
        RECT 602.800 338.300 603.600 338.400 ;
        RECT 594.800 337.700 603.600 338.300 ;
        RECT 594.800 337.600 595.600 337.700 ;
        RECT 602.800 337.600 603.600 337.700 ;
        RECT 50.800 336.300 51.600 336.400 ;
        RECT 55.600 336.300 56.400 336.400 ;
        RECT 50.800 335.700 56.400 336.300 ;
        RECT 50.800 335.600 51.600 335.700 ;
        RECT 55.600 335.600 56.400 335.700 ;
        RECT 68.400 336.300 69.200 336.400 ;
        RECT 76.400 336.300 77.200 336.400 ;
        RECT 108.400 336.300 109.200 336.400 ;
        RECT 68.400 335.700 109.200 336.300 ;
        RECT 68.400 335.600 69.200 335.700 ;
        RECT 76.400 335.600 77.200 335.700 ;
        RECT 108.400 335.600 109.200 335.700 ;
        RECT 134.000 336.300 134.800 336.400 ;
        RECT 153.200 336.300 154.000 336.400 ;
        RECT 170.800 336.300 171.600 336.400 ;
        RECT 134.000 335.700 171.600 336.300 ;
        RECT 134.000 335.600 134.800 335.700 ;
        RECT 153.200 335.600 154.000 335.700 ;
        RECT 170.800 335.600 171.600 335.700 ;
        RECT 273.200 336.300 274.000 336.400 ;
        RECT 278.000 336.300 278.800 336.400 ;
        RECT 282.800 336.300 283.600 336.400 ;
        RECT 273.200 335.700 283.600 336.300 ;
        RECT 273.200 335.600 274.000 335.700 ;
        RECT 278.000 335.600 278.800 335.700 ;
        RECT 282.800 335.600 283.600 335.700 ;
        RECT 380.400 336.300 381.200 336.400 ;
        RECT 455.600 336.300 456.400 336.400 ;
        RECT 380.400 335.700 456.400 336.300 ;
        RECT 380.400 335.600 381.200 335.700 ;
        RECT 455.600 335.600 456.400 335.700 ;
        RECT 466.800 336.300 467.600 336.400 ;
        RECT 490.800 336.300 491.600 336.400 ;
        RECT 466.800 335.700 491.600 336.300 ;
        RECT 466.800 335.600 467.600 335.700 ;
        RECT 490.800 335.600 491.600 335.700 ;
        RECT 522.800 336.300 523.600 336.400 ;
        RECT 537.200 336.300 538.000 336.400 ;
        RECT 556.400 336.300 557.200 336.400 ;
        RECT 522.800 335.700 557.200 336.300 ;
        RECT 522.800 335.600 523.600 335.700 ;
        RECT 537.200 335.600 538.000 335.700 ;
        RECT 556.400 335.600 557.200 335.700 ;
        RECT 588.400 336.300 589.200 336.400 ;
        RECT 598.000 336.300 598.800 336.400 ;
        RECT 588.400 335.700 598.800 336.300 ;
        RECT 588.400 335.600 589.200 335.700 ;
        RECT 598.000 335.600 598.800 335.700 ;
        RECT 602.800 336.300 603.600 336.400 ;
        RECT 607.600 336.300 608.400 336.400 ;
        RECT 602.800 335.700 608.400 336.300 ;
        RECT 602.800 335.600 603.600 335.700 ;
        RECT 607.600 335.600 608.400 335.700 ;
        RECT 79.600 334.300 80.400 334.400 ;
        RECT 97.200 334.300 98.000 334.400 ;
        RECT 79.600 333.700 98.000 334.300 ;
        RECT 79.600 333.600 80.400 333.700 ;
        RECT 97.200 333.600 98.000 333.700 ;
        RECT 254.000 334.300 254.800 334.400 ;
        RECT 268.400 334.300 269.200 334.400 ;
        RECT 254.000 333.700 269.200 334.300 ;
        RECT 254.000 333.600 254.800 333.700 ;
        RECT 268.400 333.600 269.200 333.700 ;
        RECT 326.000 334.300 326.800 334.400 ;
        RECT 356.400 334.300 357.200 334.400 ;
        RECT 326.000 333.700 357.200 334.300 ;
        RECT 326.000 333.600 326.800 333.700 ;
        RECT 356.400 333.600 357.200 333.700 ;
        RECT 375.600 334.300 376.400 334.400 ;
        RECT 391.600 334.300 392.400 334.400 ;
        RECT 375.600 333.700 392.400 334.300 ;
        RECT 375.600 333.600 376.400 333.700 ;
        RECT 391.600 333.600 392.400 333.700 ;
        RECT 401.200 334.300 402.000 334.400 ;
        RECT 439.600 334.300 440.400 334.400 ;
        RECT 401.200 333.700 440.400 334.300 ;
        RECT 401.200 333.600 402.000 333.700 ;
        RECT 439.600 333.600 440.400 333.700 ;
        RECT 450.800 334.300 451.600 334.400 ;
        RECT 465.200 334.300 466.000 334.400 ;
        RECT 450.800 333.700 466.000 334.300 ;
        RECT 450.800 333.600 451.600 333.700 ;
        RECT 465.200 333.600 466.000 333.700 ;
        RECT 468.400 334.300 469.200 334.400 ;
        RECT 489.200 334.300 490.000 334.400 ;
        RECT 468.400 333.700 490.000 334.300 ;
        RECT 468.400 333.600 469.200 333.700 ;
        RECT 489.200 333.600 490.000 333.700 ;
        RECT 537.200 334.300 538.000 334.400 ;
        RECT 538.800 334.300 539.600 334.400 ;
        RECT 537.200 333.700 539.600 334.300 ;
        RECT 537.200 333.600 538.000 333.700 ;
        RECT 538.800 333.600 539.600 333.700 ;
        RECT 570.800 334.300 571.600 334.400 ;
        RECT 590.000 334.300 590.800 334.400 ;
        RECT 570.800 333.700 590.800 334.300 ;
        RECT 570.800 333.600 571.600 333.700 ;
        RECT 590.000 333.600 590.800 333.700 ;
        RECT 54.000 332.300 54.800 332.400 ;
        RECT 95.600 332.300 96.400 332.400 ;
        RECT 105.200 332.300 106.000 332.400 ;
        RECT 54.000 331.700 106.000 332.300 ;
        RECT 54.000 331.600 54.800 331.700 ;
        RECT 95.600 331.600 96.400 331.700 ;
        RECT 105.200 331.600 106.000 331.700 ;
        RECT 127.600 332.300 128.400 332.400 ;
        RECT 130.800 332.300 131.600 332.400 ;
        RECT 127.600 331.700 131.600 332.300 ;
        RECT 127.600 331.600 128.400 331.700 ;
        RECT 130.800 331.600 131.600 331.700 ;
        RECT 183.600 332.300 184.400 332.400 ;
        RECT 191.600 332.300 192.400 332.400 ;
        RECT 183.600 331.700 192.400 332.300 ;
        RECT 183.600 331.600 184.400 331.700 ;
        RECT 191.600 331.600 192.400 331.700 ;
        RECT 220.400 332.300 221.200 332.400 ;
        RECT 287.600 332.300 288.400 332.400 ;
        RECT 220.400 331.700 288.400 332.300 ;
        RECT 220.400 331.600 221.200 331.700 ;
        RECT 287.600 331.600 288.400 331.700 ;
        RECT 290.800 332.300 291.600 332.400 ;
        RECT 297.200 332.300 298.000 332.400 ;
        RECT 305.200 332.300 306.000 332.400 ;
        RECT 316.400 332.300 317.200 332.400 ;
        RECT 290.800 331.700 317.200 332.300 ;
        RECT 290.800 331.600 291.600 331.700 ;
        RECT 297.200 331.600 298.000 331.700 ;
        RECT 305.200 331.600 306.000 331.700 ;
        RECT 316.400 331.600 317.200 331.700 ;
        RECT 326.000 332.300 326.800 332.400 ;
        RECT 329.200 332.300 330.000 332.400 ;
        RECT 326.000 331.700 330.000 332.300 ;
        RECT 326.000 331.600 326.800 331.700 ;
        RECT 329.200 331.600 330.000 331.700 ;
        RECT 332.400 332.300 333.200 332.400 ;
        RECT 364.400 332.300 365.200 332.400 ;
        RECT 374.000 332.300 374.800 332.400 ;
        RECT 332.400 331.700 374.800 332.300 ;
        RECT 332.400 331.600 333.200 331.700 ;
        RECT 364.400 331.600 365.200 331.700 ;
        RECT 374.000 331.600 374.800 331.700 ;
        RECT 398.000 332.300 398.800 332.400 ;
        RECT 406.000 332.300 406.800 332.400 ;
        RECT 398.000 331.700 406.800 332.300 ;
        RECT 398.000 331.600 398.800 331.700 ;
        RECT 406.000 331.600 406.800 331.700 ;
        RECT 417.200 332.300 418.000 332.400 ;
        RECT 439.700 332.300 440.300 333.600 ;
        RECT 478.000 332.300 478.800 332.400 ;
        RECT 484.400 332.300 485.200 332.400 ;
        RECT 417.200 331.700 438.700 332.300 ;
        RECT 439.700 331.700 485.200 332.300 ;
        RECT 417.200 331.600 418.000 331.700 ;
        RECT 188.400 330.300 189.200 330.400 ;
        RECT 228.400 330.300 229.200 330.400 ;
        RECT 188.400 329.700 229.200 330.300 ;
        RECT 188.400 329.600 189.200 329.700 ;
        RECT 228.400 329.600 229.200 329.700 ;
        RECT 231.600 330.300 232.400 330.400 ;
        RECT 281.200 330.300 282.000 330.400 ;
        RECT 231.600 329.700 282.000 330.300 ;
        RECT 231.600 329.600 232.400 329.700 ;
        RECT 281.200 329.600 282.000 329.700 ;
        RECT 284.400 330.300 285.200 330.400 ;
        RECT 290.800 330.300 291.600 330.400 ;
        RECT 284.400 329.700 291.600 330.300 ;
        RECT 284.400 329.600 285.200 329.700 ;
        RECT 290.800 329.600 291.600 329.700 ;
        RECT 298.800 330.300 299.600 330.400 ;
        RECT 329.200 330.300 330.000 330.400 ;
        RECT 337.200 330.300 338.000 330.400 ;
        RECT 298.800 329.700 338.000 330.300 ;
        RECT 298.800 329.600 299.600 329.700 ;
        RECT 329.200 329.600 330.000 329.700 ;
        RECT 337.200 329.600 338.000 329.700 ;
        RECT 372.400 330.300 373.200 330.400 ;
        RECT 385.200 330.300 386.000 330.400 ;
        RECT 372.400 329.700 386.000 330.300 ;
        RECT 372.400 329.600 373.200 329.700 ;
        RECT 385.200 329.600 386.000 329.700 ;
        RECT 391.600 330.300 392.400 330.400 ;
        RECT 436.400 330.300 437.200 330.400 ;
        RECT 391.600 329.700 437.200 330.300 ;
        RECT 438.100 330.300 438.700 331.700 ;
        RECT 478.000 331.600 478.800 331.700 ;
        RECT 484.400 331.600 485.200 331.700 ;
        RECT 494.000 332.300 494.800 332.400 ;
        RECT 495.600 332.300 496.400 332.400 ;
        RECT 494.000 331.700 496.400 332.300 ;
        RECT 494.000 331.600 494.800 331.700 ;
        RECT 495.600 331.600 496.400 331.700 ;
        RECT 500.400 332.300 501.200 332.400 ;
        RECT 510.000 332.300 510.800 332.400 ;
        RECT 500.400 331.700 510.800 332.300 ;
        RECT 500.400 331.600 501.200 331.700 ;
        RECT 510.000 331.600 510.800 331.700 ;
        RECT 526.000 332.300 526.800 332.400 ;
        RECT 529.200 332.300 530.000 332.400 ;
        RECT 526.000 331.700 530.000 332.300 ;
        RECT 526.000 331.600 526.800 331.700 ;
        RECT 529.200 331.600 530.000 331.700 ;
        RECT 535.600 332.300 536.400 332.400 ;
        RECT 543.600 332.300 544.400 332.400 ;
        RECT 554.800 332.300 555.600 332.400 ;
        RECT 535.600 331.700 555.600 332.300 ;
        RECT 535.600 331.600 536.400 331.700 ;
        RECT 543.600 331.600 544.400 331.700 ;
        RECT 554.800 331.600 555.600 331.700 ;
        RECT 578.800 332.300 579.600 332.400 ;
        RECT 585.200 332.300 586.000 332.400 ;
        RECT 593.200 332.300 594.000 332.400 ;
        RECT 599.600 332.300 600.400 332.400 ;
        RECT 578.800 331.700 600.400 332.300 ;
        RECT 578.800 331.600 579.600 331.700 ;
        RECT 585.200 331.600 586.000 331.700 ;
        RECT 593.200 331.600 594.000 331.700 ;
        RECT 599.600 331.600 600.400 331.700 ;
        RECT 441.200 330.300 442.000 330.400 ;
        RECT 438.100 329.700 442.000 330.300 ;
        RECT 391.600 329.600 392.400 329.700 ;
        RECT 436.400 329.600 437.200 329.700 ;
        RECT 441.200 329.600 442.000 329.700 ;
        RECT 447.600 330.300 448.400 330.400 ;
        RECT 449.200 330.300 450.000 330.400 ;
        RECT 447.600 329.700 450.000 330.300 ;
        RECT 447.600 329.600 448.400 329.700 ;
        RECT 449.200 329.600 450.000 329.700 ;
        RECT 450.800 330.300 451.600 330.400 ;
        RECT 468.400 330.300 469.200 330.400 ;
        RECT 450.800 329.700 469.200 330.300 ;
        RECT 450.800 329.600 451.600 329.700 ;
        RECT 468.400 329.600 469.200 329.700 ;
        RECT 470.000 330.300 470.800 330.400 ;
        RECT 482.800 330.300 483.600 330.400 ;
        RECT 505.200 330.300 506.000 330.400 ;
        RECT 470.000 329.700 506.000 330.300 ;
        RECT 470.000 329.600 470.800 329.700 ;
        RECT 482.800 329.600 483.600 329.700 ;
        RECT 505.200 329.600 506.000 329.700 ;
        RECT 295.600 328.300 296.400 328.400 ;
        RECT 300.400 328.300 301.200 328.400 ;
        RECT 295.600 327.700 301.200 328.300 ;
        RECT 295.600 327.600 296.400 327.700 ;
        RECT 300.400 327.600 301.200 327.700 ;
        RECT 327.600 328.300 328.400 328.400 ;
        RECT 337.200 328.300 338.000 328.400 ;
        RECT 327.600 327.700 338.000 328.300 ;
        RECT 327.600 327.600 328.400 327.700 ;
        RECT 337.200 327.600 338.000 327.700 ;
        RECT 374.000 328.300 374.800 328.400 ;
        RECT 378.800 328.300 379.600 328.400 ;
        RECT 374.000 327.700 379.600 328.300 ;
        RECT 374.000 327.600 374.800 327.700 ;
        RECT 378.800 327.600 379.600 327.700 ;
        RECT 399.600 328.300 400.400 328.400 ;
        RECT 434.800 328.300 435.600 328.400 ;
        RECT 454.000 328.300 454.800 328.400 ;
        RECT 399.600 327.700 454.800 328.300 ;
        RECT 399.600 327.600 400.400 327.700 ;
        RECT 434.800 327.600 435.600 327.700 ;
        RECT 454.000 327.600 454.800 327.700 ;
        RECT 466.800 328.300 467.600 328.400 ;
        RECT 494.000 328.300 494.800 328.400 ;
        RECT 466.800 327.700 494.800 328.300 ;
        RECT 466.800 327.600 467.600 327.700 ;
        RECT 494.000 327.600 494.800 327.700 ;
        RECT 218.800 326.300 219.600 326.400 ;
        RECT 254.000 326.300 254.800 326.400 ;
        RECT 218.800 325.700 254.800 326.300 ;
        RECT 218.800 325.600 219.600 325.700 ;
        RECT 254.000 325.600 254.800 325.700 ;
        RECT 321.200 326.300 322.000 326.400 ;
        RECT 340.400 326.300 341.200 326.400 ;
        RECT 321.200 325.700 341.200 326.300 ;
        RECT 321.200 325.600 322.000 325.700 ;
        RECT 340.400 325.600 341.200 325.700 ;
        RECT 375.600 326.300 376.400 326.400 ;
        RECT 378.800 326.300 379.600 326.400 ;
        RECT 375.600 325.700 379.600 326.300 ;
        RECT 375.600 325.600 376.400 325.700 ;
        RECT 378.800 325.600 379.600 325.700 ;
        RECT 460.400 326.300 461.200 326.400 ;
        RECT 471.600 326.300 472.400 326.400 ;
        RECT 487.600 326.300 488.400 326.400 ;
        RECT 460.400 325.700 488.400 326.300 ;
        RECT 460.400 325.600 461.200 325.700 ;
        RECT 471.600 325.600 472.400 325.700 ;
        RECT 487.600 325.600 488.400 325.700 ;
        RECT 12.400 324.300 13.200 324.400 ;
        RECT 17.200 324.300 18.000 324.400 ;
        RECT 31.600 324.300 32.400 324.400 ;
        RECT 12.400 323.700 32.400 324.300 ;
        RECT 12.400 323.600 13.200 323.700 ;
        RECT 17.200 323.600 18.000 323.700 ;
        RECT 31.600 323.600 32.400 323.700 ;
        RECT 207.600 324.300 208.400 324.400 ;
        RECT 258.800 324.300 259.600 324.400 ;
        RECT 207.600 323.700 259.600 324.300 ;
        RECT 207.600 323.600 208.400 323.700 ;
        RECT 258.800 323.600 259.600 323.700 ;
        RECT 337.200 324.300 338.000 324.400 ;
        RECT 377.200 324.300 378.000 324.400 ;
        RECT 337.200 323.700 378.000 324.300 ;
        RECT 337.200 323.600 338.000 323.700 ;
        RECT 377.200 323.600 378.000 323.700 ;
        RECT 442.800 324.300 443.600 324.400 ;
        RECT 449.200 324.300 450.000 324.400 ;
        RECT 546.800 324.300 547.600 324.400 ;
        RECT 442.800 323.700 547.600 324.300 ;
        RECT 442.800 323.600 443.600 323.700 ;
        RECT 449.200 323.600 450.000 323.700 ;
        RECT 546.800 323.600 547.600 323.700 ;
        RECT 52.400 322.300 53.200 322.400 ;
        RECT 60.400 322.300 61.200 322.400 ;
        RECT 52.400 321.700 61.200 322.300 ;
        RECT 52.400 321.600 53.200 321.700 ;
        RECT 60.400 321.600 61.200 321.700 ;
        RECT 103.600 322.300 104.400 322.400 ;
        RECT 110.000 322.300 110.800 322.400 ;
        RECT 103.600 321.700 110.800 322.300 ;
        RECT 103.600 321.600 104.400 321.700 ;
        RECT 110.000 321.600 110.800 321.700 ;
        RECT 210.800 322.300 211.600 322.400 ;
        RECT 217.200 322.300 218.000 322.400 ;
        RECT 210.800 321.700 218.000 322.300 ;
        RECT 210.800 321.600 211.600 321.700 ;
        RECT 217.200 321.600 218.000 321.700 ;
        RECT 314.800 322.300 315.600 322.400 ;
        RECT 324.400 322.300 325.200 322.400 ;
        RECT 314.800 321.700 325.200 322.300 ;
        RECT 314.800 321.600 315.600 321.700 ;
        RECT 324.400 321.600 325.200 321.700 ;
        RECT 340.400 322.300 341.200 322.400 ;
        RECT 383.600 322.300 384.400 322.400 ;
        RECT 340.400 321.700 384.400 322.300 ;
        RECT 340.400 321.600 341.200 321.700 ;
        RECT 383.600 321.600 384.400 321.700 ;
        RECT 490.800 322.300 491.600 322.400 ;
        RECT 510.000 322.300 510.800 322.400 ;
        RECT 518.000 322.300 518.800 322.400 ;
        RECT 490.800 321.700 518.800 322.300 ;
        RECT 490.800 321.600 491.600 321.700 ;
        RECT 510.000 321.600 510.800 321.700 ;
        RECT 518.000 321.600 518.800 321.700 ;
        RECT 519.600 322.300 520.400 322.400 ;
        RECT 524.400 322.300 525.200 322.400 ;
        RECT 519.600 321.700 525.200 322.300 ;
        RECT 519.600 321.600 520.400 321.700 ;
        RECT 524.400 321.600 525.200 321.700 ;
        RECT 535.600 322.300 536.400 322.400 ;
        RECT 558.000 322.300 558.800 322.400 ;
        RECT 535.600 321.700 558.800 322.300 ;
        RECT 535.600 321.600 536.400 321.700 ;
        RECT 558.000 321.600 558.800 321.700 ;
        RECT 1.200 320.300 2.000 320.400 ;
        RECT 14.000 320.300 14.800 320.400 ;
        RECT 38.000 320.300 38.800 320.400 ;
        RECT 138.800 320.300 139.600 320.400 ;
        RECT 142.000 320.300 142.800 320.400 ;
        RECT 1.200 319.700 142.800 320.300 ;
        RECT 324.500 320.300 325.100 321.600 ;
        RECT 398.000 320.300 398.800 320.400 ;
        RECT 324.500 319.700 398.800 320.300 ;
        RECT 1.200 319.600 2.000 319.700 ;
        RECT 14.000 319.600 14.800 319.700 ;
        RECT 38.000 319.600 38.800 319.700 ;
        RECT 138.800 319.600 139.600 319.700 ;
        RECT 142.000 319.600 142.800 319.700 ;
        RECT 398.000 319.600 398.800 319.700 ;
        RECT 423.600 320.300 424.400 320.400 ;
        RECT 433.200 320.300 434.000 320.400 ;
        RECT 423.600 319.700 434.000 320.300 ;
        RECT 423.600 319.600 424.400 319.700 ;
        RECT 433.200 319.600 434.000 319.700 ;
        RECT 444.400 320.300 445.200 320.400 ;
        RECT 450.800 320.300 451.600 320.400 ;
        RECT 444.400 319.700 451.600 320.300 ;
        RECT 444.400 319.600 445.200 319.700 ;
        RECT 450.800 319.600 451.600 319.700 ;
        RECT 465.200 320.300 466.000 320.400 ;
        RECT 506.800 320.300 507.600 320.400 ;
        RECT 521.200 320.300 522.000 320.400 ;
        RECT 465.200 319.700 522.000 320.300 ;
        RECT 465.200 319.600 466.000 319.700 ;
        RECT 506.800 319.600 507.600 319.700 ;
        RECT 521.200 319.600 522.000 319.700 ;
        RECT 44.400 318.300 45.200 318.400 ;
        RECT 47.600 318.300 48.400 318.400 ;
        RECT 44.400 317.700 48.400 318.300 ;
        RECT 44.400 317.600 45.200 317.700 ;
        RECT 47.600 317.600 48.400 317.700 ;
        RECT 102.000 318.300 102.800 318.400 ;
        RECT 110.000 318.300 110.800 318.400 ;
        RECT 102.000 317.700 110.800 318.300 ;
        RECT 102.000 317.600 102.800 317.700 ;
        RECT 110.000 317.600 110.800 317.700 ;
        RECT 129.200 318.300 130.000 318.400 ;
        RECT 161.200 318.300 162.000 318.400 ;
        RECT 129.200 317.700 162.000 318.300 ;
        RECT 129.200 317.600 130.000 317.700 ;
        RECT 161.200 317.600 162.000 317.700 ;
        RECT 206.000 318.300 206.800 318.400 ;
        RECT 346.800 318.300 347.600 318.400 ;
        RECT 206.000 317.700 347.600 318.300 ;
        RECT 206.000 317.600 206.800 317.700 ;
        RECT 346.800 317.600 347.600 317.700 ;
        RECT 359.600 318.300 360.400 318.400 ;
        RECT 375.600 318.300 376.400 318.400 ;
        RECT 359.600 317.700 376.400 318.300 ;
        RECT 359.600 317.600 360.400 317.700 ;
        RECT 375.600 317.600 376.400 317.700 ;
        RECT 399.600 318.300 400.400 318.400 ;
        RECT 404.400 318.300 405.200 318.400 ;
        RECT 399.600 317.700 405.200 318.300 ;
        RECT 399.600 317.600 400.400 317.700 ;
        RECT 404.400 317.600 405.200 317.700 ;
        RECT 436.400 318.300 437.200 318.400 ;
        RECT 460.400 318.300 461.200 318.400 ;
        RECT 481.200 318.300 482.000 318.400 ;
        RECT 490.800 318.300 491.600 318.400 ;
        RECT 502.000 318.300 502.800 318.400 ;
        RECT 513.200 318.300 514.000 318.400 ;
        RECT 522.800 318.300 523.600 318.400 ;
        RECT 436.400 317.700 461.200 318.300 ;
        RECT 436.400 317.600 437.200 317.700 ;
        RECT 460.400 317.600 461.200 317.700 ;
        RECT 462.100 317.700 489.900 318.300 ;
        RECT 238.000 316.300 238.800 316.400 ;
        RECT 388.400 316.300 389.200 316.400 ;
        RECT 238.000 315.700 389.200 316.300 ;
        RECT 238.000 315.600 238.800 315.700 ;
        RECT 388.400 315.600 389.200 315.700 ;
        RECT 402.800 316.300 403.600 316.400 ;
        RECT 418.800 316.300 419.600 316.400 ;
        RECT 402.800 315.700 419.600 316.300 ;
        RECT 402.800 315.600 403.600 315.700 ;
        RECT 418.800 315.600 419.600 315.700 ;
        RECT 454.000 316.300 454.800 316.400 ;
        RECT 457.200 316.300 458.000 316.400 ;
        RECT 454.000 315.700 458.000 316.300 ;
        RECT 454.000 315.600 454.800 315.700 ;
        RECT 457.200 315.600 458.000 315.700 ;
        RECT 458.800 316.300 459.600 316.400 ;
        RECT 462.100 316.300 462.700 317.700 ;
        RECT 481.200 317.600 482.000 317.700 ;
        RECT 458.800 315.700 462.700 316.300 ;
        RECT 465.200 316.300 466.000 316.400 ;
        RECT 487.600 316.300 488.400 316.400 ;
        RECT 465.200 315.700 488.400 316.300 ;
        RECT 489.300 316.300 489.900 317.700 ;
        RECT 490.800 317.700 523.600 318.300 ;
        RECT 490.800 317.600 491.600 317.700 ;
        RECT 502.000 317.600 502.800 317.700 ;
        RECT 513.200 317.600 514.000 317.700 ;
        RECT 522.800 317.600 523.600 317.700 ;
        RECT 500.400 316.300 501.200 316.400 ;
        RECT 489.300 315.700 501.200 316.300 ;
        RECT 458.800 315.600 459.600 315.700 ;
        RECT 465.200 315.600 466.000 315.700 ;
        RECT 487.600 315.600 488.400 315.700 ;
        RECT 500.400 315.600 501.200 315.700 ;
        RECT 265.200 314.300 266.000 314.400 ;
        RECT 270.000 314.300 270.800 314.400 ;
        RECT 265.200 313.700 270.800 314.300 ;
        RECT 265.200 313.600 266.000 313.700 ;
        RECT 270.000 313.600 270.800 313.700 ;
        RECT 289.200 314.300 290.000 314.400 ;
        RECT 311.600 314.300 312.400 314.400 ;
        RECT 289.200 313.700 312.400 314.300 ;
        RECT 289.200 313.600 290.000 313.700 ;
        RECT 311.600 313.600 312.400 313.700 ;
        RECT 334.000 314.300 334.800 314.400 ;
        RECT 358.000 314.300 358.800 314.400 ;
        RECT 372.400 314.300 373.200 314.400 ;
        RECT 334.000 313.700 373.200 314.300 ;
        RECT 334.000 313.600 334.800 313.700 ;
        RECT 358.000 313.600 358.800 313.700 ;
        RECT 372.400 313.600 373.200 313.700 ;
        RECT 375.600 314.300 376.400 314.400 ;
        RECT 465.200 314.300 466.000 314.400 ;
        RECT 375.600 313.700 466.000 314.300 ;
        RECT 375.600 313.600 376.400 313.700 ;
        RECT 465.200 313.600 466.000 313.700 ;
        RECT 478.000 314.300 478.800 314.400 ;
        RECT 481.200 314.300 482.000 314.400 ;
        RECT 478.000 313.700 482.000 314.300 ;
        RECT 478.000 313.600 478.800 313.700 ;
        RECT 481.200 313.600 482.000 313.700 ;
        RECT 484.400 314.300 485.200 314.400 ;
        RECT 502.000 314.300 502.800 314.400 ;
        RECT 484.400 313.700 502.800 314.300 ;
        RECT 484.400 313.600 485.200 313.700 ;
        RECT 502.000 313.600 502.800 313.700 ;
        RECT 503.600 314.300 504.400 314.400 ;
        RECT 508.400 314.300 509.200 314.400 ;
        RECT 503.600 313.700 509.200 314.300 ;
        RECT 503.600 313.600 504.400 313.700 ;
        RECT 508.400 313.600 509.200 313.700 ;
        RECT 527.600 314.300 528.400 314.400 ;
        RECT 532.400 314.300 533.200 314.400 ;
        RECT 527.600 313.700 533.200 314.300 ;
        RECT 527.600 313.600 528.400 313.700 ;
        RECT 532.400 313.600 533.200 313.700 ;
        RECT 583.600 314.300 584.400 314.400 ;
        RECT 586.800 314.300 587.600 314.400 ;
        RECT 583.600 313.700 587.600 314.300 ;
        RECT 583.600 313.600 584.400 313.700 ;
        RECT 586.800 313.600 587.600 313.700 ;
        RECT 79.600 312.300 80.400 312.400 ;
        RECT 118.000 312.300 118.800 312.400 ;
        RECT 79.600 311.700 118.800 312.300 ;
        RECT 79.600 311.600 80.400 311.700 ;
        RECT 118.000 311.600 118.800 311.700 ;
        RECT 137.200 312.300 138.000 312.400 ;
        RECT 169.200 312.300 170.000 312.400 ;
        RECT 137.200 311.700 170.000 312.300 ;
        RECT 137.200 311.600 138.000 311.700 ;
        RECT 169.200 311.600 170.000 311.700 ;
        RECT 191.600 312.300 192.400 312.400 ;
        RECT 204.400 312.300 205.200 312.400 ;
        RECT 191.600 311.700 205.200 312.300 ;
        RECT 191.600 311.600 192.400 311.700 ;
        RECT 204.400 311.600 205.200 311.700 ;
        RECT 239.600 312.300 240.400 312.400 ;
        RECT 257.200 312.300 258.000 312.400 ;
        RECT 271.600 312.300 272.400 312.400 ;
        RECT 239.600 311.700 258.000 312.300 ;
        RECT 239.600 311.600 240.400 311.700 ;
        RECT 257.200 311.600 258.000 311.700 ;
        RECT 258.900 311.700 272.400 312.300 ;
        RECT 57.200 310.300 58.000 310.400 ;
        RECT 87.600 310.300 88.400 310.400 ;
        RECT 57.200 309.700 88.400 310.300 ;
        RECT 57.200 309.600 58.000 309.700 ;
        RECT 87.600 309.600 88.400 309.700 ;
        RECT 103.600 310.300 104.400 310.400 ;
        RECT 129.200 310.300 130.000 310.400 ;
        RECT 103.600 309.700 130.000 310.300 ;
        RECT 103.600 309.600 104.400 309.700 ;
        RECT 129.200 309.600 130.000 309.700 ;
        RECT 146.800 310.300 147.600 310.400 ;
        RECT 156.400 310.300 157.200 310.400 ;
        RECT 146.800 309.700 157.200 310.300 ;
        RECT 146.800 309.600 147.600 309.700 ;
        RECT 156.400 309.600 157.200 309.700 ;
        RECT 196.400 309.600 197.200 310.400 ;
        RECT 233.200 310.300 234.000 310.400 ;
        RECT 238.000 310.300 238.800 310.400 ;
        RECT 233.200 309.700 238.800 310.300 ;
        RECT 233.200 309.600 234.000 309.700 ;
        RECT 238.000 309.600 238.800 309.700 ;
        RECT 247.600 310.300 248.400 310.400 ;
        RECT 258.900 310.300 259.500 311.700 ;
        RECT 271.600 311.600 272.400 311.700 ;
        RECT 273.200 312.300 274.000 312.400 ;
        RECT 274.800 312.300 275.600 312.400 ;
        RECT 273.200 311.700 275.600 312.300 ;
        RECT 273.200 311.600 274.000 311.700 ;
        RECT 274.800 311.600 275.600 311.700 ;
        RECT 284.400 312.300 285.200 312.400 ;
        RECT 292.400 312.300 293.200 312.400 ;
        RECT 284.400 311.700 293.200 312.300 ;
        RECT 284.400 311.600 285.200 311.700 ;
        RECT 292.400 311.600 293.200 311.700 ;
        RECT 348.400 312.300 349.200 312.400 ;
        RECT 370.800 312.300 371.600 312.400 ;
        RECT 348.400 311.700 371.600 312.300 ;
        RECT 348.400 311.600 349.200 311.700 ;
        RECT 370.800 311.600 371.600 311.700 ;
        RECT 385.200 312.300 386.000 312.400 ;
        RECT 396.400 312.300 397.200 312.400 ;
        RECT 385.200 311.700 397.200 312.300 ;
        RECT 385.200 311.600 386.000 311.700 ;
        RECT 396.400 311.600 397.200 311.700 ;
        RECT 401.200 312.300 402.000 312.400 ;
        RECT 407.600 312.300 408.400 312.400 ;
        RECT 401.200 311.700 408.400 312.300 ;
        RECT 401.200 311.600 402.000 311.700 ;
        RECT 407.600 311.600 408.400 311.700 ;
        RECT 410.800 312.300 411.600 312.400 ;
        RECT 412.400 312.300 413.200 312.400 ;
        RECT 410.800 311.700 413.200 312.300 ;
        RECT 410.800 311.600 411.600 311.700 ;
        RECT 412.400 311.600 413.200 311.700 ;
        RECT 474.800 312.300 475.600 312.400 ;
        RECT 479.600 312.300 480.400 312.400 ;
        RECT 474.800 311.700 480.400 312.300 ;
        RECT 474.800 311.600 475.600 311.700 ;
        RECT 479.600 311.600 480.400 311.700 ;
        RECT 486.000 312.300 486.800 312.400 ;
        RECT 506.800 312.300 507.600 312.400 ;
        RECT 486.000 311.700 507.600 312.300 ;
        RECT 486.000 311.600 486.800 311.700 ;
        RECT 506.800 311.600 507.600 311.700 ;
        RECT 511.600 312.300 512.400 312.400 ;
        RECT 521.200 312.300 522.000 312.400 ;
        RECT 522.800 312.300 523.600 312.400 ;
        RECT 511.600 311.700 523.600 312.300 ;
        RECT 511.600 311.600 512.400 311.700 ;
        RECT 521.200 311.600 522.000 311.700 ;
        RECT 522.800 311.600 523.600 311.700 ;
        RECT 529.200 312.300 530.000 312.400 ;
        RECT 538.800 312.300 539.600 312.400 ;
        RECT 529.200 311.700 539.600 312.300 ;
        RECT 529.200 311.600 530.000 311.700 ;
        RECT 538.800 311.600 539.600 311.700 ;
        RECT 575.600 312.300 576.400 312.400 ;
        RECT 585.200 312.300 586.000 312.400 ;
        RECT 575.600 311.700 586.000 312.300 ;
        RECT 575.600 311.600 576.400 311.700 ;
        RECT 585.200 311.600 586.000 311.700 ;
        RECT 247.600 309.700 259.500 310.300 ;
        RECT 262.000 310.300 262.800 310.400 ;
        RECT 284.400 310.300 285.200 310.400 ;
        RECT 297.200 310.300 298.000 310.400 ;
        RECT 262.000 309.700 298.000 310.300 ;
        RECT 247.600 309.600 248.400 309.700 ;
        RECT 262.000 309.600 262.800 309.700 ;
        RECT 284.400 309.600 285.200 309.700 ;
        RECT 297.200 309.600 298.000 309.700 ;
        RECT 370.800 310.300 371.600 310.400 ;
        RECT 375.600 310.300 376.400 310.400 ;
        RECT 370.800 309.700 376.400 310.300 ;
        RECT 370.800 309.600 371.600 309.700 ;
        RECT 375.600 309.600 376.400 309.700 ;
        RECT 378.800 310.300 379.600 310.400 ;
        RECT 383.600 310.300 384.400 310.400 ;
        RECT 378.800 309.700 384.400 310.300 ;
        RECT 378.800 309.600 379.600 309.700 ;
        RECT 383.600 309.600 384.400 309.700 ;
        RECT 391.600 310.300 392.400 310.400 ;
        RECT 404.400 310.300 405.200 310.400 ;
        RECT 391.600 309.700 405.200 310.300 ;
        RECT 391.600 309.600 392.400 309.700 ;
        RECT 404.400 309.600 405.200 309.700 ;
        RECT 407.600 310.300 408.400 310.400 ;
        RECT 417.200 310.300 418.000 310.400 ;
        RECT 407.600 309.700 418.000 310.300 ;
        RECT 407.600 309.600 408.400 309.700 ;
        RECT 417.200 309.600 418.000 309.700 ;
        RECT 423.600 310.300 424.400 310.400 ;
        RECT 438.000 310.300 438.800 310.400 ;
        RECT 423.600 309.700 438.800 310.300 ;
        RECT 423.600 309.600 424.400 309.700 ;
        RECT 438.000 309.600 438.800 309.700 ;
        RECT 466.800 310.300 467.600 310.400 ;
        RECT 468.400 310.300 469.200 310.400 ;
        RECT 466.800 309.700 469.200 310.300 ;
        RECT 466.800 309.600 467.600 309.700 ;
        RECT 468.400 309.600 469.200 309.700 ;
        RECT 471.600 310.300 472.400 310.400 ;
        RECT 476.400 310.300 477.200 310.400 ;
        RECT 471.600 309.700 477.200 310.300 ;
        RECT 471.600 309.600 472.400 309.700 ;
        RECT 476.400 309.600 477.200 309.700 ;
        RECT 495.600 310.300 496.400 310.400 ;
        RECT 498.800 310.300 499.600 310.400 ;
        RECT 495.600 309.700 499.600 310.300 ;
        RECT 495.600 309.600 496.400 309.700 ;
        RECT 498.800 309.600 499.600 309.700 ;
        RECT 500.400 309.600 501.200 310.400 ;
        RECT 505.200 310.300 506.000 310.400 ;
        RECT 511.600 310.300 512.400 310.400 ;
        RECT 505.200 309.700 512.400 310.300 ;
        RECT 505.200 309.600 506.000 309.700 ;
        RECT 511.600 309.600 512.400 309.700 ;
        RECT 526.000 310.300 526.800 310.400 ;
        RECT 534.000 310.300 534.800 310.400 ;
        RECT 526.000 309.700 534.800 310.300 ;
        RECT 526.000 309.600 526.800 309.700 ;
        RECT 534.000 309.600 534.800 309.700 ;
        RECT 28.400 308.300 29.200 308.400 ;
        RECT 49.200 308.300 50.000 308.400 ;
        RECT 28.400 307.700 50.000 308.300 ;
        RECT 28.400 307.600 29.200 307.700 ;
        RECT 49.200 307.600 50.000 307.700 ;
        RECT 71.600 308.300 72.400 308.400 ;
        RECT 86.000 308.300 86.800 308.400 ;
        RECT 71.600 307.700 86.800 308.300 ;
        RECT 71.600 307.600 72.400 307.700 ;
        RECT 86.000 307.600 86.800 307.700 ;
        RECT 97.200 308.300 98.000 308.400 ;
        RECT 262.100 308.300 262.700 309.600 ;
        RECT 97.200 307.700 262.700 308.300 ;
        RECT 268.400 308.300 269.200 308.400 ;
        RECT 270.000 308.300 270.800 308.400 ;
        RECT 268.400 307.700 270.800 308.300 ;
        RECT 97.200 307.600 98.000 307.700 ;
        RECT 268.400 307.600 269.200 307.700 ;
        RECT 270.000 307.600 270.800 307.700 ;
        RECT 279.600 308.300 280.400 308.400 ;
        RECT 282.800 308.300 283.600 308.400 ;
        RECT 279.600 307.700 283.600 308.300 ;
        RECT 279.600 307.600 280.400 307.700 ;
        RECT 282.800 307.600 283.600 307.700 ;
        RECT 287.600 308.300 288.400 308.400 ;
        RECT 298.800 308.300 299.600 308.400 ;
        RECT 332.400 308.300 333.200 308.400 ;
        RECT 287.600 307.700 333.200 308.300 ;
        RECT 287.600 307.600 288.400 307.700 ;
        RECT 298.800 307.600 299.600 307.700 ;
        RECT 332.400 307.600 333.200 307.700 ;
        RECT 346.800 308.300 347.600 308.400 ;
        RECT 369.200 308.300 370.000 308.400 ;
        RECT 346.800 307.700 370.000 308.300 ;
        RECT 346.800 307.600 347.600 307.700 ;
        RECT 369.200 307.600 370.000 307.700 ;
        RECT 377.200 308.300 378.000 308.400 ;
        RECT 378.800 308.300 379.600 308.400 ;
        RECT 377.200 307.700 379.600 308.300 ;
        RECT 377.200 307.600 378.000 307.700 ;
        RECT 378.800 307.600 379.600 307.700 ;
        RECT 380.400 308.300 381.200 308.400 ;
        RECT 390.000 308.300 390.800 308.400 ;
        RECT 380.400 307.700 390.800 308.300 ;
        RECT 380.400 307.600 381.200 307.700 ;
        RECT 390.000 307.600 390.800 307.700 ;
        RECT 391.600 308.300 392.400 308.400 ;
        RECT 393.200 308.300 394.000 308.400 ;
        RECT 391.600 307.700 394.000 308.300 ;
        RECT 391.600 307.600 392.400 307.700 ;
        RECT 393.200 307.600 394.000 307.700 ;
        RECT 398.000 308.300 398.800 308.400 ;
        RECT 404.400 308.300 405.200 308.400 ;
        RECT 409.200 308.300 410.000 308.400 ;
        RECT 398.000 307.700 410.000 308.300 ;
        RECT 398.000 307.600 398.800 307.700 ;
        RECT 404.400 307.600 405.200 307.700 ;
        RECT 409.200 307.600 410.000 307.700 ;
        RECT 410.800 308.300 411.600 308.400 ;
        RECT 449.200 308.300 450.000 308.400 ;
        RECT 490.800 308.300 491.600 308.400 ;
        RECT 410.800 307.700 491.600 308.300 ;
        RECT 410.800 307.600 411.600 307.700 ;
        RECT 449.200 307.600 450.000 307.700 ;
        RECT 490.800 307.600 491.600 307.700 ;
        RECT 500.400 308.300 501.200 308.400 ;
        RECT 503.600 308.300 504.400 308.400 ;
        RECT 500.400 307.700 504.400 308.300 ;
        RECT 500.400 307.600 501.200 307.700 ;
        RECT 503.600 307.600 504.400 307.700 ;
        RECT 516.400 308.300 517.200 308.400 ;
        RECT 529.200 308.300 530.000 308.400 ;
        RECT 516.400 307.700 530.000 308.300 ;
        RECT 516.400 307.600 517.200 307.700 ;
        RECT 529.200 307.600 530.000 307.700 ;
        RECT 562.800 308.300 563.600 308.400 ;
        RECT 585.200 308.300 586.000 308.400 ;
        RECT 562.800 307.700 586.000 308.300 ;
        RECT 562.800 307.600 563.600 307.700 ;
        RECT 585.200 307.600 586.000 307.700 ;
        RECT 590.000 308.300 590.800 308.400 ;
        RECT 599.600 308.300 600.400 308.400 ;
        RECT 590.000 307.700 600.400 308.300 ;
        RECT 590.000 307.600 590.800 307.700 ;
        RECT 599.600 307.600 600.400 307.700 ;
        RECT 31.600 306.300 32.400 306.400 ;
        RECT 68.400 306.300 69.200 306.400 ;
        RECT 31.600 305.700 69.200 306.300 ;
        RECT 31.600 305.600 32.400 305.700 ;
        RECT 68.400 305.600 69.200 305.700 ;
        RECT 92.400 306.300 93.200 306.400 ;
        RECT 207.600 306.300 208.400 306.400 ;
        RECT 92.400 305.700 208.400 306.300 ;
        RECT 92.400 305.600 93.200 305.700 ;
        RECT 207.600 305.600 208.400 305.700 ;
        RECT 214.000 306.300 214.800 306.400 ;
        RECT 246.000 306.300 246.800 306.400 ;
        RECT 214.000 305.700 246.800 306.300 ;
        RECT 214.000 305.600 214.800 305.700 ;
        RECT 246.000 305.600 246.800 305.700 ;
        RECT 290.800 306.300 291.600 306.400 ;
        RECT 306.800 306.300 307.600 306.400 ;
        RECT 324.400 306.300 325.200 306.400 ;
        RECT 290.800 305.700 325.200 306.300 ;
        RECT 290.800 305.600 291.600 305.700 ;
        RECT 306.800 305.600 307.600 305.700 ;
        RECT 324.400 305.600 325.200 305.700 ;
        RECT 353.200 306.300 354.000 306.400 ;
        RECT 356.400 306.300 357.200 306.400 ;
        RECT 394.800 306.300 395.600 306.400 ;
        RECT 353.200 305.700 395.600 306.300 ;
        RECT 353.200 305.600 354.000 305.700 ;
        RECT 356.400 305.600 357.200 305.700 ;
        RECT 394.800 305.600 395.600 305.700 ;
        RECT 396.400 306.300 397.200 306.400 ;
        RECT 402.800 306.300 403.600 306.400 ;
        RECT 396.400 305.700 403.600 306.300 ;
        RECT 396.400 305.600 397.200 305.700 ;
        RECT 402.800 305.600 403.600 305.700 ;
        RECT 414.000 306.300 414.800 306.400 ;
        RECT 417.200 306.300 418.000 306.400 ;
        RECT 441.200 306.300 442.000 306.400 ;
        RECT 414.000 305.700 442.000 306.300 ;
        RECT 414.000 305.600 414.800 305.700 ;
        RECT 417.200 305.600 418.000 305.700 ;
        RECT 441.200 305.600 442.000 305.700 ;
        RECT 479.600 306.300 480.400 306.400 ;
        RECT 492.400 306.300 493.200 306.400 ;
        RECT 479.600 305.700 493.200 306.300 ;
        RECT 479.600 305.600 480.400 305.700 ;
        RECT 492.400 305.600 493.200 305.700 ;
        RECT 494.000 306.300 494.800 306.400 ;
        RECT 511.600 306.300 512.400 306.400 ;
        RECT 494.000 305.700 512.400 306.300 ;
        RECT 494.000 305.600 494.800 305.700 ;
        RECT 511.600 305.600 512.400 305.700 ;
        RECT 538.800 306.300 539.600 306.400 ;
        RECT 542.000 306.300 542.800 306.400 ;
        RECT 538.800 305.700 542.800 306.300 ;
        RECT 538.800 305.600 539.600 305.700 ;
        RECT 542.000 305.600 542.800 305.700 ;
        RECT 574.000 306.300 574.800 306.400 ;
        RECT 578.800 306.300 579.600 306.400 ;
        RECT 574.000 305.700 579.600 306.300 ;
        RECT 574.000 305.600 574.800 305.700 ;
        RECT 578.800 305.600 579.600 305.700 ;
        RECT 582.000 306.300 582.800 306.400 ;
        RECT 593.200 306.300 594.000 306.400 ;
        RECT 604.400 306.300 605.200 306.400 ;
        RECT 582.000 305.700 605.200 306.300 ;
        RECT 582.000 305.600 582.800 305.700 ;
        RECT 593.200 305.600 594.000 305.700 ;
        RECT 604.400 305.600 605.200 305.700 ;
        RECT 169.200 304.300 170.000 304.400 ;
        RECT 180.400 304.300 181.200 304.400 ;
        RECT 169.200 303.700 181.200 304.300 ;
        RECT 169.200 303.600 170.000 303.700 ;
        RECT 180.400 303.600 181.200 303.700 ;
        RECT 186.800 304.300 187.600 304.400 ;
        RECT 217.200 304.300 218.000 304.400 ;
        RECT 234.800 304.300 235.600 304.400 ;
        RECT 186.800 303.700 235.600 304.300 ;
        RECT 186.800 303.600 187.600 303.700 ;
        RECT 217.200 303.600 218.000 303.700 ;
        RECT 234.800 303.600 235.600 303.700 ;
        RECT 263.600 304.300 264.400 304.400 ;
        RECT 289.200 304.300 290.000 304.400 ;
        RECT 263.600 303.700 290.000 304.300 ;
        RECT 263.600 303.600 264.400 303.700 ;
        RECT 289.200 303.600 290.000 303.700 ;
        RECT 314.800 303.600 315.600 304.400 ;
        RECT 318.000 304.300 318.800 304.400 ;
        RECT 338.800 304.300 339.600 304.400 ;
        RECT 318.000 303.700 339.600 304.300 ;
        RECT 318.000 303.600 318.800 303.700 ;
        RECT 338.800 303.600 339.600 303.700 ;
        RECT 404.400 304.300 405.200 304.400 ;
        RECT 449.200 304.300 450.000 304.400 ;
        RECT 404.400 303.700 450.000 304.300 ;
        RECT 404.400 303.600 405.200 303.700 ;
        RECT 449.200 303.600 450.000 303.700 ;
        RECT 450.800 304.300 451.600 304.400 ;
        RECT 481.200 304.300 482.000 304.400 ;
        RECT 450.800 303.700 482.000 304.300 ;
        RECT 450.800 303.600 451.600 303.700 ;
        RECT 481.200 303.600 482.000 303.700 ;
        RECT 526.000 304.300 526.800 304.400 ;
        RECT 534.000 304.300 534.800 304.400 ;
        RECT 526.000 303.700 534.800 304.300 ;
        RECT 526.000 303.600 526.800 303.700 ;
        RECT 534.000 303.600 534.800 303.700 ;
        RECT 554.800 304.300 555.600 304.400 ;
        RECT 566.000 304.300 566.800 304.400 ;
        RECT 580.400 304.300 581.200 304.400 ;
        RECT 593.200 304.300 594.000 304.400 ;
        RECT 554.800 303.700 594.000 304.300 ;
        RECT 554.800 303.600 555.600 303.700 ;
        RECT 566.000 303.600 566.800 303.700 ;
        RECT 580.400 303.600 581.200 303.700 ;
        RECT 593.200 303.600 594.000 303.700 ;
        RECT 122.800 302.300 123.600 302.400 ;
        RECT 143.600 302.300 144.400 302.400 ;
        RECT 122.800 301.700 144.400 302.300 ;
        RECT 122.800 301.600 123.600 301.700 ;
        RECT 143.600 301.600 144.400 301.700 ;
        RECT 158.000 302.300 158.800 302.400 ;
        RECT 263.600 302.300 264.400 302.400 ;
        RECT 158.000 301.700 264.400 302.300 ;
        RECT 158.000 301.600 158.800 301.700 ;
        RECT 263.600 301.600 264.400 301.700 ;
        RECT 278.000 302.300 278.800 302.400 ;
        RECT 295.600 302.300 296.400 302.400 ;
        RECT 278.000 301.700 296.400 302.300 ;
        RECT 278.000 301.600 278.800 301.700 ;
        RECT 295.600 301.600 296.400 301.700 ;
        RECT 390.000 302.300 390.800 302.400 ;
        RECT 401.200 302.300 402.000 302.400 ;
        RECT 390.000 301.700 402.000 302.300 ;
        RECT 390.000 301.600 390.800 301.700 ;
        RECT 401.200 301.600 402.000 301.700 ;
        RECT 412.400 302.300 413.200 302.400 ;
        RECT 418.800 302.300 419.600 302.400 ;
        RECT 412.400 301.700 419.600 302.300 ;
        RECT 412.400 301.600 413.200 301.700 ;
        RECT 418.800 301.600 419.600 301.700 ;
        RECT 420.400 302.300 421.200 302.400 ;
        RECT 442.800 302.300 443.600 302.400 ;
        RECT 420.400 301.700 443.600 302.300 ;
        RECT 420.400 301.600 421.200 301.700 ;
        RECT 442.800 301.600 443.600 301.700 ;
        RECT 476.400 302.300 477.200 302.400 ;
        RECT 486.000 302.300 486.800 302.400 ;
        RECT 476.400 301.700 486.800 302.300 ;
        RECT 476.400 301.600 477.200 301.700 ;
        RECT 486.000 301.600 486.800 301.700 ;
        RECT 497.200 302.300 498.000 302.400 ;
        RECT 500.400 302.300 501.200 302.400 ;
        RECT 497.200 301.700 501.200 302.300 ;
        RECT 497.200 301.600 498.000 301.700 ;
        RECT 500.400 301.600 501.200 301.700 ;
        RECT 521.200 302.300 522.000 302.400 ;
        RECT 526.000 302.300 526.800 302.400 ;
        RECT 542.000 302.300 542.800 302.400 ;
        RECT 521.200 301.700 542.800 302.300 ;
        RECT 521.200 301.600 522.000 301.700 ;
        RECT 526.000 301.600 526.800 301.700 ;
        RECT 542.000 301.600 542.800 301.700 ;
        RECT 572.400 302.300 573.200 302.400 ;
        RECT 590.000 302.300 590.800 302.400 ;
        RECT 572.400 301.700 590.800 302.300 ;
        RECT 572.400 301.600 573.200 301.700 ;
        RECT 590.000 301.600 590.800 301.700 ;
        RECT 415.600 300.300 416.400 300.400 ;
        RECT 434.800 300.300 435.600 300.400 ;
        RECT 415.600 299.700 435.600 300.300 ;
        RECT 415.600 299.600 416.400 299.700 ;
        RECT 434.800 299.600 435.600 299.700 ;
        RECT 450.800 300.300 451.600 300.400 ;
        RECT 470.000 300.300 470.800 300.400 ;
        RECT 450.800 299.700 470.800 300.300 ;
        RECT 450.800 299.600 451.600 299.700 ;
        RECT 470.000 299.600 470.800 299.700 ;
        RECT 471.600 300.300 472.400 300.400 ;
        RECT 489.200 300.300 490.000 300.400 ;
        RECT 502.000 300.300 502.800 300.400 ;
        RECT 471.600 299.700 488.300 300.300 ;
        RECT 471.600 299.600 472.400 299.700 ;
        RECT 294.000 298.300 294.800 298.400 ;
        RECT 298.800 298.300 299.600 298.400 ;
        RECT 294.000 297.700 299.600 298.300 ;
        RECT 294.000 297.600 294.800 297.700 ;
        RECT 298.800 297.600 299.600 297.700 ;
        RECT 311.600 298.300 312.400 298.400 ;
        RECT 316.400 298.300 317.200 298.400 ;
        RECT 311.600 297.700 317.200 298.300 ;
        RECT 311.600 297.600 312.400 297.700 ;
        RECT 316.400 297.600 317.200 297.700 ;
        RECT 332.400 298.300 333.200 298.400 ;
        RECT 359.600 298.300 360.400 298.400 ;
        RECT 332.400 297.700 360.400 298.300 ;
        RECT 332.400 297.600 333.200 297.700 ;
        RECT 359.600 297.600 360.400 297.700 ;
        RECT 377.200 298.300 378.000 298.400 ;
        RECT 388.400 298.300 389.200 298.400 ;
        RECT 401.200 298.300 402.000 298.400 ;
        RECT 377.200 297.700 402.000 298.300 ;
        RECT 487.700 298.300 488.300 299.700 ;
        RECT 489.200 299.700 502.800 300.300 ;
        RECT 489.200 299.600 490.000 299.700 ;
        RECT 502.000 299.600 502.800 299.700 ;
        RECT 590.000 300.300 590.800 300.400 ;
        RECT 594.800 300.300 595.600 300.400 ;
        RECT 590.000 299.700 595.600 300.300 ;
        RECT 590.000 299.600 590.800 299.700 ;
        RECT 594.800 299.600 595.600 299.700 ;
        RECT 489.200 298.300 490.000 298.400 ;
        RECT 494.000 298.300 494.800 298.400 ;
        RECT 487.700 297.700 494.800 298.300 ;
        RECT 377.200 297.600 378.000 297.700 ;
        RECT 388.400 297.600 389.200 297.700 ;
        RECT 401.200 297.600 402.000 297.700 ;
        RECT 489.200 297.600 490.000 297.700 ;
        RECT 494.000 297.600 494.800 297.700 ;
        RECT 506.800 298.300 507.600 298.400 ;
        RECT 521.200 298.300 522.000 298.400 ;
        RECT 506.800 297.700 522.000 298.300 ;
        RECT 506.800 297.600 507.600 297.700 ;
        RECT 521.200 297.600 522.000 297.700 ;
        RECT 28.400 296.300 29.200 296.400 ;
        RECT 57.200 296.300 58.000 296.400 ;
        RECT 28.400 295.700 58.000 296.300 ;
        RECT 28.400 295.600 29.200 295.700 ;
        RECT 57.200 295.600 58.000 295.700 ;
        RECT 58.800 296.300 59.600 296.400 ;
        RECT 86.000 296.300 86.800 296.400 ;
        RECT 108.400 296.300 109.200 296.400 ;
        RECT 58.800 295.700 109.200 296.300 ;
        RECT 58.800 295.600 59.600 295.700 ;
        RECT 86.000 295.600 86.800 295.700 ;
        RECT 108.400 295.600 109.200 295.700 ;
        RECT 126.000 296.300 126.800 296.400 ;
        RECT 138.800 296.300 139.600 296.400 ;
        RECT 177.200 296.300 178.000 296.400 ;
        RECT 126.000 295.700 178.000 296.300 ;
        RECT 126.000 295.600 126.800 295.700 ;
        RECT 138.800 295.600 139.600 295.700 ;
        RECT 177.200 295.600 178.000 295.700 ;
        RECT 247.600 296.300 248.400 296.400 ;
        RECT 282.800 296.300 283.600 296.400 ;
        RECT 314.800 296.300 315.600 296.400 ;
        RECT 247.600 295.700 315.600 296.300 ;
        RECT 247.600 295.600 248.400 295.700 ;
        RECT 282.800 295.600 283.600 295.700 ;
        RECT 314.800 295.600 315.600 295.700 ;
        RECT 338.800 296.300 339.600 296.400 ;
        RECT 348.400 296.300 349.200 296.400 ;
        RECT 399.600 296.300 400.400 296.400 ;
        RECT 338.800 295.700 400.400 296.300 ;
        RECT 338.800 295.600 339.600 295.700 ;
        RECT 348.400 295.600 349.200 295.700 ;
        RECT 399.600 295.600 400.400 295.700 ;
        RECT 415.600 296.300 416.400 296.400 ;
        RECT 417.200 296.300 418.000 296.400 ;
        RECT 415.600 295.700 418.000 296.300 ;
        RECT 415.600 295.600 416.400 295.700 ;
        RECT 417.200 295.600 418.000 295.700 ;
        RECT 457.200 296.300 458.000 296.400 ;
        RECT 466.800 296.300 467.600 296.400 ;
        RECT 500.400 296.300 501.200 296.400 ;
        RECT 457.200 295.700 467.600 296.300 ;
        RECT 457.200 295.600 458.000 295.700 ;
        RECT 466.800 295.600 467.600 295.700 ;
        RECT 494.100 295.700 501.200 296.300 ;
        RECT 14.000 294.300 14.800 294.400 ;
        RECT 17.200 294.300 18.000 294.400 ;
        RECT 31.600 294.300 32.400 294.400 ;
        RECT 78.000 294.300 78.800 294.400 ;
        RECT 14.000 293.700 78.800 294.300 ;
        RECT 14.000 293.600 14.800 293.700 ;
        RECT 17.200 293.600 18.000 293.700 ;
        RECT 31.600 293.600 32.400 293.700 ;
        RECT 78.000 293.600 78.800 293.700 ;
        RECT 100.400 294.300 101.200 294.400 ;
        RECT 105.200 294.300 106.000 294.400 ;
        RECT 142.000 294.300 142.800 294.400 ;
        RECT 154.800 294.300 155.600 294.400 ;
        RECT 100.400 293.700 121.900 294.300 ;
        RECT 100.400 293.600 101.200 293.700 ;
        RECT 105.200 293.600 106.000 293.700 ;
        RECT 121.300 292.400 121.900 293.700 ;
        RECT 142.000 293.700 155.600 294.300 ;
        RECT 142.000 293.600 142.800 293.700 ;
        RECT 154.800 293.600 155.600 293.700 ;
        RECT 183.600 294.300 184.400 294.400 ;
        RECT 204.400 294.300 205.200 294.400 ;
        RECT 183.600 293.700 205.200 294.300 ;
        RECT 183.600 293.600 184.400 293.700 ;
        RECT 204.400 293.600 205.200 293.700 ;
        RECT 206.000 294.300 206.800 294.400 ;
        RECT 209.200 294.300 210.000 294.400 ;
        RECT 206.000 293.700 210.000 294.300 ;
        RECT 206.000 293.600 206.800 293.700 ;
        RECT 209.200 293.600 210.000 293.700 ;
        RECT 231.600 294.300 232.400 294.400 ;
        RECT 257.200 294.300 258.000 294.400 ;
        RECT 231.600 293.700 258.000 294.300 ;
        RECT 231.600 293.600 232.400 293.700 ;
        RECT 257.200 293.600 258.000 293.700 ;
        RECT 294.000 294.300 294.800 294.400 ;
        RECT 327.600 294.300 328.400 294.400 ;
        RECT 294.000 293.700 328.400 294.300 ;
        RECT 294.000 293.600 294.800 293.700 ;
        RECT 327.600 293.600 328.400 293.700 ;
        RECT 329.200 294.300 330.000 294.400 ;
        RECT 351.600 294.300 352.400 294.400 ;
        RECT 329.200 293.700 352.400 294.300 ;
        RECT 329.200 293.600 330.000 293.700 ;
        RECT 351.600 293.600 352.400 293.700 ;
        RECT 354.800 294.300 355.600 294.400 ;
        RECT 367.600 294.300 368.400 294.400 ;
        RECT 354.800 293.700 368.400 294.300 ;
        RECT 354.800 293.600 355.600 293.700 ;
        RECT 367.600 293.600 368.400 293.700 ;
        RECT 374.000 294.300 374.800 294.400 ;
        RECT 380.400 294.300 381.200 294.400 ;
        RECT 374.000 293.700 381.200 294.300 ;
        RECT 374.000 293.600 374.800 293.700 ;
        RECT 380.400 293.600 381.200 293.700 ;
        RECT 386.800 294.300 387.600 294.400 ;
        RECT 391.600 294.300 392.400 294.400 ;
        RECT 386.800 293.700 392.400 294.300 ;
        RECT 386.800 293.600 387.600 293.700 ;
        RECT 391.600 293.600 392.400 293.700 ;
        RECT 438.000 294.300 438.800 294.400 ;
        RECT 447.600 294.300 448.400 294.400 ;
        RECT 450.800 294.300 451.600 294.400 ;
        RECT 438.000 293.700 451.600 294.300 ;
        RECT 438.000 293.600 438.800 293.700 ;
        RECT 447.600 293.600 448.400 293.700 ;
        RECT 450.800 293.600 451.600 293.700 ;
        RECT 463.600 294.300 464.400 294.400 ;
        RECT 473.200 294.300 474.000 294.400 ;
        RECT 463.600 293.700 474.000 294.300 ;
        RECT 463.600 293.600 464.400 293.700 ;
        RECT 473.200 293.600 474.000 293.700 ;
        RECT 474.800 294.300 475.600 294.400 ;
        RECT 479.600 294.300 480.400 294.400 ;
        RECT 474.800 293.700 480.400 294.300 ;
        RECT 474.800 293.600 475.600 293.700 ;
        RECT 479.600 293.600 480.400 293.700 ;
        RECT 482.800 294.300 483.600 294.400 ;
        RECT 484.400 294.300 485.200 294.400 ;
        RECT 482.800 293.700 485.200 294.300 ;
        RECT 482.800 293.600 483.600 293.700 ;
        RECT 484.400 293.600 485.200 293.700 ;
        RECT 489.200 294.300 490.000 294.400 ;
        RECT 494.100 294.300 494.700 295.700 ;
        RECT 500.400 295.600 501.200 295.700 ;
        RECT 506.800 296.300 507.600 296.400 ;
        RECT 519.600 296.300 520.400 296.400 ;
        RECT 506.800 295.700 520.400 296.300 ;
        RECT 506.800 295.600 507.600 295.700 ;
        RECT 519.600 295.600 520.400 295.700 ;
        RECT 537.200 296.300 538.000 296.400 ;
        RECT 558.000 296.300 558.800 296.400 ;
        RECT 537.200 295.700 558.800 296.300 ;
        RECT 537.200 295.600 538.000 295.700 ;
        RECT 558.000 295.600 558.800 295.700 ;
        RECT 489.200 293.700 494.700 294.300 ;
        RECT 495.600 294.300 496.400 294.400 ;
        RECT 506.800 294.300 507.600 294.400 ;
        RECT 510.000 294.300 510.800 294.400 ;
        RECT 495.600 293.700 510.800 294.300 ;
        RECT 489.200 293.600 490.000 293.700 ;
        RECT 495.600 293.600 496.400 293.700 ;
        RECT 506.800 293.600 507.600 293.700 ;
        RECT 510.000 293.600 510.800 293.700 ;
        RECT 513.200 294.300 514.000 294.400 ;
        RECT 518.000 294.300 518.800 294.400 ;
        RECT 513.200 293.700 518.800 294.300 ;
        RECT 513.200 293.600 514.000 293.700 ;
        RECT 518.000 293.600 518.800 293.700 ;
        RECT 535.600 294.300 536.400 294.400 ;
        RECT 542.000 294.300 542.800 294.400 ;
        RECT 554.800 294.300 555.600 294.400 ;
        RECT 535.600 293.700 555.600 294.300 ;
        RECT 535.600 293.600 536.400 293.700 ;
        RECT 542.000 293.600 542.800 293.700 ;
        RECT 554.800 293.600 555.600 293.700 ;
        RECT 580.400 294.300 581.200 294.400 ;
        RECT 593.200 294.300 594.000 294.400 ;
        RECT 580.400 293.700 594.000 294.300 ;
        RECT 580.400 293.600 581.200 293.700 ;
        RECT 593.200 293.600 594.000 293.700 ;
        RECT 74.800 292.300 75.600 292.400 ;
        RECT 102.000 292.300 102.800 292.400 ;
        RECT 74.800 291.700 102.800 292.300 ;
        RECT 74.800 291.600 75.600 291.700 ;
        RECT 102.000 291.600 102.800 291.700 ;
        RECT 110.000 292.300 110.800 292.400 ;
        RECT 118.000 292.300 118.800 292.400 ;
        RECT 110.000 291.700 118.800 292.300 ;
        RECT 110.000 291.600 110.800 291.700 ;
        RECT 118.000 291.600 118.800 291.700 ;
        RECT 121.200 292.300 122.000 292.400 ;
        RECT 156.400 292.300 157.200 292.400 ;
        RECT 164.400 292.300 165.200 292.400 ;
        RECT 121.200 291.700 165.200 292.300 ;
        RECT 121.200 291.600 122.000 291.700 ;
        RECT 156.400 291.600 157.200 291.700 ;
        RECT 164.400 291.600 165.200 291.700 ;
        RECT 199.600 292.300 200.400 292.400 ;
        RECT 222.000 292.300 222.800 292.400 ;
        RECT 199.600 291.700 222.800 292.300 ;
        RECT 199.600 291.600 200.400 291.700 ;
        RECT 222.000 291.600 222.800 291.700 ;
        RECT 255.600 292.300 256.400 292.400 ;
        RECT 270.000 292.300 270.800 292.400 ;
        RECT 255.600 291.700 270.800 292.300 ;
        RECT 255.600 291.600 256.400 291.700 ;
        RECT 270.000 291.600 270.800 291.700 ;
        RECT 279.600 292.300 280.400 292.400 ;
        RECT 305.200 292.300 306.000 292.400 ;
        RECT 279.600 291.700 306.000 292.300 ;
        RECT 279.600 291.600 280.400 291.700 ;
        RECT 305.200 291.600 306.000 291.700 ;
        RECT 322.800 292.300 323.600 292.400 ;
        RECT 330.800 292.300 331.600 292.400 ;
        RECT 322.800 291.700 331.600 292.300 ;
        RECT 322.800 291.600 323.600 291.700 ;
        RECT 330.800 291.600 331.600 291.700 ;
        RECT 345.200 292.300 346.000 292.400 ;
        RECT 361.200 292.300 362.000 292.400 ;
        RECT 345.200 291.700 362.000 292.300 ;
        RECT 345.200 291.600 346.000 291.700 ;
        RECT 361.200 291.600 362.000 291.700 ;
        RECT 370.800 292.300 371.600 292.400 ;
        RECT 402.800 292.300 403.600 292.400 ;
        RECT 370.800 291.700 403.600 292.300 ;
        RECT 370.800 291.600 371.600 291.700 ;
        RECT 402.800 291.600 403.600 291.700 ;
        RECT 439.600 292.300 440.400 292.400 ;
        RECT 447.600 292.300 448.400 292.400 ;
        RECT 439.600 291.700 448.400 292.300 ;
        RECT 439.600 291.600 440.400 291.700 ;
        RECT 447.600 291.600 448.400 291.700 ;
        RECT 462.000 292.300 462.800 292.400 ;
        RECT 468.400 292.300 469.200 292.400 ;
        RECT 462.000 291.700 469.200 292.300 ;
        RECT 462.000 291.600 462.800 291.700 ;
        RECT 468.400 291.600 469.200 291.700 ;
        RECT 478.000 292.300 478.800 292.400 ;
        RECT 492.400 292.300 493.200 292.400 ;
        RECT 478.000 291.700 493.200 292.300 ;
        RECT 478.000 291.600 478.800 291.700 ;
        RECT 492.400 291.600 493.200 291.700 ;
        RECT 494.000 292.300 494.800 292.400 ;
        RECT 498.800 292.300 499.600 292.400 ;
        RECT 494.000 291.700 499.600 292.300 ;
        RECT 494.000 291.600 494.800 291.700 ;
        RECT 498.800 291.600 499.600 291.700 ;
        RECT 521.200 292.300 522.000 292.400 ;
        RECT 526.000 292.300 526.800 292.400 ;
        RECT 521.200 291.700 526.800 292.300 ;
        RECT 521.200 291.600 522.000 291.700 ;
        RECT 526.000 291.600 526.800 291.700 ;
        RECT 554.800 292.300 555.600 292.400 ;
        RECT 558.000 292.300 558.800 292.400 ;
        RECT 554.800 291.700 558.800 292.300 ;
        RECT 554.800 291.600 555.600 291.700 ;
        RECT 558.000 291.600 558.800 291.700 ;
        RECT 54.000 290.300 54.800 290.400 ;
        RECT 58.800 290.300 59.600 290.400 ;
        RECT 54.000 289.700 59.600 290.300 ;
        RECT 54.000 289.600 54.800 289.700 ;
        RECT 58.800 289.600 59.600 289.700 ;
        RECT 95.600 290.300 96.400 290.400 ;
        RECT 111.600 290.300 112.400 290.400 ;
        RECT 169.200 290.300 170.000 290.400 ;
        RECT 196.400 290.300 197.200 290.400 ;
        RECT 95.600 289.700 197.200 290.300 ;
        RECT 95.600 289.600 96.400 289.700 ;
        RECT 111.600 289.600 112.400 289.700 ;
        RECT 169.200 289.600 170.000 289.700 ;
        RECT 196.400 289.600 197.200 289.700 ;
        RECT 214.000 290.300 214.800 290.400 ;
        RECT 242.800 290.300 243.600 290.400 ;
        RECT 292.400 290.300 293.200 290.400 ;
        RECT 305.200 290.300 306.000 290.400 ;
        RECT 214.000 289.700 306.000 290.300 ;
        RECT 214.000 289.600 214.800 289.700 ;
        RECT 242.800 289.600 243.600 289.700 ;
        RECT 292.400 289.600 293.200 289.700 ;
        RECT 305.200 289.600 306.000 289.700 ;
        RECT 314.800 290.300 315.600 290.400 ;
        RECT 322.800 290.300 323.600 290.400 ;
        RECT 314.800 289.700 323.600 290.300 ;
        RECT 314.800 289.600 315.600 289.700 ;
        RECT 322.800 289.600 323.600 289.700 ;
        RECT 326.000 290.300 326.800 290.400 ;
        RECT 334.000 290.300 334.800 290.400 ;
        RECT 326.000 289.700 334.800 290.300 ;
        RECT 326.000 289.600 326.800 289.700 ;
        RECT 334.000 289.600 334.800 289.700 ;
        RECT 351.600 290.300 352.400 290.400 ;
        RECT 359.600 290.300 360.400 290.400 ;
        RECT 351.600 289.700 360.400 290.300 ;
        RECT 351.600 289.600 352.400 289.700 ;
        RECT 359.600 289.600 360.400 289.700 ;
        RECT 394.800 290.300 395.600 290.400 ;
        RECT 495.600 290.300 496.400 290.400 ;
        RECT 518.000 290.300 518.800 290.400 ;
        RECT 394.800 289.700 469.100 290.300 ;
        RECT 394.800 289.600 395.600 289.700 ;
        RECT 151.600 288.300 152.400 288.400 ;
        RECT 175.600 288.300 176.400 288.400 ;
        RECT 151.600 287.700 176.400 288.300 ;
        RECT 151.600 287.600 152.400 287.700 ;
        RECT 175.600 287.600 176.400 287.700 ;
        RECT 290.800 288.300 291.600 288.400 ;
        RECT 354.800 288.300 355.600 288.400 ;
        RECT 290.800 287.700 355.600 288.300 ;
        RECT 290.800 287.600 291.600 287.700 ;
        RECT 354.800 287.600 355.600 287.700 ;
        RECT 366.000 288.300 366.800 288.400 ;
        RECT 380.400 288.300 381.200 288.400 ;
        RECT 366.000 287.700 381.200 288.300 ;
        RECT 366.000 287.600 366.800 287.700 ;
        RECT 380.400 287.600 381.200 287.700 ;
        RECT 382.000 288.300 382.800 288.400 ;
        RECT 430.000 288.300 430.800 288.400 ;
        RECT 382.000 287.700 430.800 288.300 ;
        RECT 382.000 287.600 382.800 287.700 ;
        RECT 430.000 287.600 430.800 287.700 ;
        RECT 434.800 288.300 435.600 288.400 ;
        RECT 452.400 288.300 453.200 288.400 ;
        RECT 434.800 287.700 453.200 288.300 ;
        RECT 434.800 287.600 435.600 287.700 ;
        RECT 452.400 287.600 453.200 287.700 ;
        RECT 463.600 288.300 464.400 288.400 ;
        RECT 466.800 288.300 467.600 288.400 ;
        RECT 463.600 287.700 467.600 288.300 ;
        RECT 468.500 288.300 469.100 289.700 ;
        RECT 495.600 289.700 518.800 290.300 ;
        RECT 495.600 289.600 496.400 289.700 ;
        RECT 518.000 289.600 518.800 289.700 ;
        RECT 530.800 290.300 531.600 290.400 ;
        RECT 538.800 290.300 539.600 290.400 ;
        RECT 530.800 289.700 539.600 290.300 ;
        RECT 530.800 289.600 531.600 289.700 ;
        RECT 538.800 289.600 539.600 289.700 ;
        RECT 530.900 288.300 531.500 289.600 ;
        RECT 468.500 287.700 531.500 288.300 ;
        RECT 463.600 287.600 464.400 287.700 ;
        RECT 466.800 287.600 467.600 287.700 ;
        RECT 106.800 286.300 107.600 286.400 ;
        RECT 113.200 286.300 114.000 286.400 ;
        RECT 266.800 286.300 267.600 286.400 ;
        RECT 106.800 285.700 267.600 286.300 ;
        RECT 106.800 285.600 107.600 285.700 ;
        RECT 113.200 285.600 114.000 285.700 ;
        RECT 266.800 285.600 267.600 285.700 ;
        RECT 313.200 286.300 314.000 286.400 ;
        RECT 329.200 286.300 330.000 286.400 ;
        RECT 313.200 285.700 330.000 286.300 ;
        RECT 313.200 285.600 314.000 285.700 ;
        RECT 329.200 285.600 330.000 285.700 ;
        RECT 334.000 286.300 334.800 286.400 ;
        RECT 342.000 286.300 342.800 286.400 ;
        RECT 346.800 286.300 347.600 286.400 ;
        RECT 334.000 285.700 347.600 286.300 ;
        RECT 334.000 285.600 334.800 285.700 ;
        RECT 342.000 285.600 342.800 285.700 ;
        RECT 346.800 285.600 347.600 285.700 ;
        RECT 362.800 286.300 363.600 286.400 ;
        RECT 385.200 286.300 386.000 286.400 ;
        RECT 362.800 285.700 386.000 286.300 ;
        RECT 362.800 285.600 363.600 285.700 ;
        RECT 385.200 285.600 386.000 285.700 ;
        RECT 390.000 286.300 390.800 286.400 ;
        RECT 396.400 286.300 397.200 286.400 ;
        RECT 390.000 285.700 397.200 286.300 ;
        RECT 390.000 285.600 390.800 285.700 ;
        RECT 396.400 285.600 397.200 285.700 ;
        RECT 404.400 286.300 405.200 286.400 ;
        RECT 406.000 286.300 406.800 286.400 ;
        RECT 404.400 285.700 406.800 286.300 ;
        RECT 404.400 285.600 405.200 285.700 ;
        RECT 406.000 285.600 406.800 285.700 ;
        RECT 439.600 286.300 440.400 286.400 ;
        RECT 471.600 286.300 472.400 286.400 ;
        RECT 439.600 285.700 472.400 286.300 ;
        RECT 439.600 285.600 440.400 285.700 ;
        RECT 471.600 285.600 472.400 285.700 ;
        RECT 500.400 286.300 501.200 286.400 ;
        RECT 521.200 286.300 522.000 286.400 ;
        RECT 500.400 285.700 522.000 286.300 ;
        RECT 500.400 285.600 501.200 285.700 ;
        RECT 521.200 285.600 522.000 285.700 ;
        RECT 39.600 284.300 40.400 284.400 ;
        RECT 47.600 284.300 48.400 284.400 ;
        RECT 39.600 283.700 48.400 284.300 ;
        RECT 39.600 283.600 40.400 283.700 ;
        RECT 47.600 283.600 48.400 283.700 ;
        RECT 89.200 284.300 90.000 284.400 ;
        RECT 94.000 284.300 94.800 284.400 ;
        RECT 89.200 283.700 94.800 284.300 ;
        RECT 89.200 283.600 90.000 283.700 ;
        RECT 94.000 283.600 94.800 283.700 ;
        RECT 143.600 284.300 144.400 284.400 ;
        RECT 206.000 284.300 206.800 284.400 ;
        RECT 143.600 283.700 206.800 284.300 ;
        RECT 143.600 283.600 144.400 283.700 ;
        RECT 206.000 283.600 206.800 283.700 ;
        RECT 207.600 284.300 208.400 284.400 ;
        RECT 236.400 284.300 237.200 284.400 ;
        RECT 244.400 284.300 245.200 284.400 ;
        RECT 207.600 283.700 245.200 284.300 ;
        RECT 207.600 283.600 208.400 283.700 ;
        RECT 236.400 283.600 237.200 283.700 ;
        RECT 244.400 283.600 245.200 283.700 ;
        RECT 250.800 283.600 251.600 284.400 ;
        RECT 292.400 284.300 293.200 284.400 ;
        RECT 314.800 284.300 315.600 284.400 ;
        RECT 292.400 283.700 315.600 284.300 ;
        RECT 292.400 283.600 293.200 283.700 ;
        RECT 314.800 283.600 315.600 283.700 ;
        RECT 319.600 284.300 320.400 284.400 ;
        RECT 327.600 284.300 328.400 284.400 ;
        RECT 319.600 283.700 328.400 284.300 ;
        RECT 319.600 283.600 320.400 283.700 ;
        RECT 327.600 283.600 328.400 283.700 ;
        RECT 369.200 284.300 370.000 284.400 ;
        RECT 383.600 284.300 384.400 284.400 ;
        RECT 369.200 283.700 384.400 284.300 ;
        RECT 369.200 283.600 370.000 283.700 ;
        RECT 383.600 283.600 384.400 283.700 ;
        RECT 399.600 284.300 400.400 284.400 ;
        RECT 463.600 284.300 464.400 284.400 ;
        RECT 399.600 283.700 464.400 284.300 ;
        RECT 399.600 283.600 400.400 283.700 ;
        RECT 463.600 283.600 464.400 283.700 ;
        RECT 465.200 284.300 466.000 284.400 ;
        RECT 481.200 284.300 482.000 284.400 ;
        RECT 465.200 283.700 482.000 284.300 ;
        RECT 465.200 283.600 466.000 283.700 ;
        RECT 481.200 283.600 482.000 283.700 ;
        RECT 186.800 282.300 187.600 282.400 ;
        RECT 191.600 282.300 192.400 282.400 ;
        RECT 186.800 281.700 192.400 282.300 ;
        RECT 186.800 281.600 187.600 281.700 ;
        RECT 191.600 281.600 192.400 281.700 ;
        RECT 228.400 282.300 229.200 282.400 ;
        RECT 249.200 282.300 250.000 282.400 ;
        RECT 228.400 281.700 250.000 282.300 ;
        RECT 228.400 281.600 229.200 281.700 ;
        RECT 249.200 281.600 250.000 281.700 ;
        RECT 266.800 282.300 267.600 282.400 ;
        RECT 276.400 282.300 277.200 282.400 ;
        RECT 266.800 281.700 277.200 282.300 ;
        RECT 266.800 281.600 267.600 281.700 ;
        RECT 276.400 281.600 277.200 281.700 ;
        RECT 321.200 282.300 322.000 282.400 ;
        RECT 324.400 282.300 325.200 282.400 ;
        RECT 321.200 281.700 325.200 282.300 ;
        RECT 321.200 281.600 322.000 281.700 ;
        RECT 324.400 281.600 325.200 281.700 ;
        RECT 335.600 282.300 336.400 282.400 ;
        RECT 364.400 282.300 365.200 282.400 ;
        RECT 378.800 282.300 379.600 282.400 ;
        RECT 385.200 282.300 386.000 282.400 ;
        RECT 335.600 281.700 386.000 282.300 ;
        RECT 335.600 281.600 336.400 281.700 ;
        RECT 364.400 281.600 365.200 281.700 ;
        RECT 378.800 281.600 379.600 281.700 ;
        RECT 385.200 281.600 386.000 281.700 ;
        RECT 478.000 282.300 478.800 282.400 ;
        RECT 479.600 282.300 480.400 282.400 ;
        RECT 478.000 281.700 480.400 282.300 ;
        RECT 478.000 281.600 478.800 281.700 ;
        RECT 479.600 281.600 480.400 281.700 ;
        RECT 487.600 282.300 488.400 282.400 ;
        RECT 497.200 282.300 498.000 282.400 ;
        RECT 487.600 281.700 498.000 282.300 ;
        RECT 487.600 281.600 488.400 281.700 ;
        RECT 497.200 281.600 498.000 281.700 ;
        RECT 506.800 282.300 507.600 282.400 ;
        RECT 513.200 282.300 514.000 282.400 ;
        RECT 530.800 282.300 531.600 282.400 ;
        RECT 506.800 281.700 531.600 282.300 ;
        RECT 506.800 281.600 507.600 281.700 ;
        RECT 513.200 281.600 514.000 281.700 ;
        RECT 530.800 281.600 531.600 281.700 ;
        RECT 602.800 282.300 603.600 282.400 ;
        RECT 606.000 282.300 606.800 282.400 ;
        RECT 609.200 282.300 610.000 282.400 ;
        RECT 602.800 281.700 610.000 282.300 ;
        RECT 602.800 281.600 603.600 281.700 ;
        RECT 606.000 281.600 606.800 281.700 ;
        RECT 609.200 281.600 610.000 281.700 ;
        RECT 81.200 280.300 82.000 280.400 ;
        RECT 97.200 280.300 98.000 280.400 ;
        RECT 81.200 279.700 98.000 280.300 ;
        RECT 81.200 279.600 82.000 279.700 ;
        RECT 97.200 279.600 98.000 279.700 ;
        RECT 194.800 280.300 195.600 280.400 ;
        RECT 199.600 280.300 200.400 280.400 ;
        RECT 273.200 280.300 274.000 280.400 ;
        RECT 279.600 280.300 280.400 280.400 ;
        RECT 289.200 280.300 290.000 280.400 ;
        RECT 326.000 280.300 326.800 280.400 ;
        RECT 194.800 279.700 326.800 280.300 ;
        RECT 194.800 279.600 195.600 279.700 ;
        RECT 199.600 279.600 200.400 279.700 ;
        RECT 273.200 279.600 274.000 279.700 ;
        RECT 279.600 279.600 280.400 279.700 ;
        RECT 289.200 279.600 290.000 279.700 ;
        RECT 326.000 279.600 326.800 279.700 ;
        RECT 334.000 280.300 334.800 280.400 ;
        RECT 340.400 280.300 341.200 280.400 ;
        RECT 433.200 280.300 434.000 280.400 ;
        RECT 474.800 280.300 475.600 280.400 ;
        RECT 334.000 279.700 341.200 280.300 ;
        RECT 334.000 279.600 334.800 279.700 ;
        RECT 340.400 279.600 341.200 279.700 ;
        RECT 342.100 279.700 434.000 280.300 ;
        RECT 250.800 278.300 251.600 278.400 ;
        RECT 342.100 278.300 342.700 279.700 ;
        RECT 433.200 279.600 434.000 279.700 ;
        RECT 463.700 279.700 475.600 280.300 ;
        RECT 250.800 277.700 342.700 278.300 ;
        RECT 361.200 278.300 362.000 278.400 ;
        RECT 390.000 278.300 390.800 278.400 ;
        RECT 361.200 277.700 390.800 278.300 ;
        RECT 250.800 277.600 251.600 277.700 ;
        RECT 361.200 277.600 362.000 277.700 ;
        RECT 390.000 277.600 390.800 277.700 ;
        RECT 401.200 278.300 402.000 278.400 ;
        RECT 420.400 278.300 421.200 278.400 ;
        RECT 401.200 277.700 421.200 278.300 ;
        RECT 401.200 277.600 402.000 277.700 ;
        RECT 420.400 277.600 421.200 277.700 ;
        RECT 442.800 278.300 443.600 278.400 ;
        RECT 463.700 278.300 464.300 279.700 ;
        RECT 474.800 279.600 475.600 279.700 ;
        RECT 490.800 280.300 491.600 280.400 ;
        RECT 505.200 280.300 506.000 280.400 ;
        RECT 522.800 280.300 523.600 280.400 ;
        RECT 490.800 279.700 523.600 280.300 ;
        RECT 490.800 279.600 491.600 279.700 ;
        RECT 505.200 279.600 506.000 279.700 ;
        RECT 522.800 279.600 523.600 279.700 ;
        RECT 529.200 280.300 530.000 280.400 ;
        RECT 537.200 280.300 538.000 280.400 ;
        RECT 529.200 279.700 538.000 280.300 ;
        RECT 529.200 279.600 530.000 279.700 ;
        RECT 537.200 279.600 538.000 279.700 ;
        RECT 442.800 277.700 464.300 278.300 ;
        RECT 465.200 278.300 466.000 278.400 ;
        RECT 468.400 278.300 469.200 278.400 ;
        RECT 500.400 278.300 501.200 278.400 ;
        RECT 465.200 277.700 501.200 278.300 ;
        RECT 442.800 277.600 443.600 277.700 ;
        RECT 465.200 277.600 466.000 277.700 ;
        RECT 468.400 277.600 469.200 277.700 ;
        RECT 500.400 277.600 501.200 277.700 ;
        RECT 519.600 278.300 520.400 278.400 ;
        RECT 532.400 278.300 533.200 278.400 ;
        RECT 519.600 277.700 533.200 278.300 ;
        RECT 519.600 277.600 520.400 277.700 ;
        RECT 532.400 277.600 533.200 277.700 ;
        RECT 122.800 276.300 123.600 276.400 ;
        RECT 130.800 276.300 131.600 276.400 ;
        RECT 122.800 275.700 131.600 276.300 ;
        RECT 122.800 275.600 123.600 275.700 ;
        RECT 130.800 275.600 131.600 275.700 ;
        RECT 174.000 276.300 174.800 276.400 ;
        RECT 196.400 276.300 197.200 276.400 ;
        RECT 338.800 276.300 339.600 276.400 ;
        RECT 174.000 275.700 339.600 276.300 ;
        RECT 174.000 275.600 174.800 275.700 ;
        RECT 196.400 275.600 197.200 275.700 ;
        RECT 338.800 275.600 339.600 275.700 ;
        RECT 359.600 275.600 360.400 276.400 ;
        RECT 372.400 276.300 373.200 276.400 ;
        RECT 382.000 276.300 382.800 276.400 ;
        RECT 372.400 275.700 382.800 276.300 ;
        RECT 372.400 275.600 373.200 275.700 ;
        RECT 382.000 275.600 382.800 275.700 ;
        RECT 399.600 276.300 400.400 276.400 ;
        RECT 433.200 276.300 434.000 276.400 ;
        RECT 399.600 275.700 434.000 276.300 ;
        RECT 399.600 275.600 400.400 275.700 ;
        RECT 433.200 275.600 434.000 275.700 ;
        RECT 466.800 276.300 467.600 276.400 ;
        RECT 474.800 276.300 475.600 276.400 ;
        RECT 466.800 275.700 475.600 276.300 ;
        RECT 466.800 275.600 467.600 275.700 ;
        RECT 474.800 275.600 475.600 275.700 ;
        RECT 487.600 276.300 488.400 276.400 ;
        RECT 519.600 276.300 520.400 276.400 ;
        RECT 487.600 275.700 520.400 276.300 ;
        RECT 487.600 275.600 488.400 275.700 ;
        RECT 519.600 275.600 520.400 275.700 ;
        RECT 527.600 276.300 528.400 276.400 ;
        RECT 529.200 276.300 530.000 276.400 ;
        RECT 527.600 275.700 530.000 276.300 ;
        RECT 527.600 275.600 528.400 275.700 ;
        RECT 529.200 275.600 530.000 275.700 ;
        RECT 534.000 276.300 534.800 276.400 ;
        RECT 556.400 276.300 557.200 276.400 ;
        RECT 567.600 276.300 568.400 276.400 ;
        RECT 534.000 275.700 568.400 276.300 ;
        RECT 534.000 275.600 534.800 275.700 ;
        RECT 556.400 275.600 557.200 275.700 ;
        RECT 567.600 275.600 568.400 275.700 ;
        RECT 572.400 276.300 573.200 276.400 ;
        RECT 575.600 276.300 576.400 276.400 ;
        RECT 578.800 276.300 579.600 276.400 ;
        RECT 572.400 275.700 579.600 276.300 ;
        RECT 572.400 275.600 573.200 275.700 ;
        RECT 575.600 275.600 576.400 275.700 ;
        RECT 578.800 275.600 579.600 275.700 ;
        RECT 84.400 274.300 85.200 274.400 ;
        RECT 92.400 274.300 93.200 274.400 ;
        RECT 84.400 273.700 93.200 274.300 ;
        RECT 84.400 273.600 85.200 273.700 ;
        RECT 92.400 273.600 93.200 273.700 ;
        RECT 110.000 274.300 110.800 274.400 ;
        RECT 122.800 274.300 123.600 274.400 ;
        RECT 212.400 274.300 213.200 274.400 ;
        RECT 110.000 273.700 213.200 274.300 ;
        RECT 110.000 273.600 110.800 273.700 ;
        RECT 122.800 273.600 123.600 273.700 ;
        RECT 212.400 273.600 213.200 273.700 ;
        RECT 217.200 274.300 218.000 274.400 ;
        RECT 295.600 274.300 296.400 274.400 ;
        RECT 298.800 274.300 299.600 274.400 ;
        RECT 217.200 273.700 280.300 274.300 ;
        RECT 217.200 273.600 218.000 273.700 ;
        RECT 65.200 272.300 66.000 272.400 ;
        RECT 68.400 272.300 69.200 272.400 ;
        RECT 92.400 272.300 93.200 272.400 ;
        RECT 65.200 271.700 93.200 272.300 ;
        RECT 65.200 271.600 66.000 271.700 ;
        RECT 68.400 271.600 69.200 271.700 ;
        RECT 92.400 271.600 93.200 271.700 ;
        RECT 164.400 272.300 165.200 272.400 ;
        RECT 169.200 272.300 170.000 272.400 ;
        RECT 164.400 271.700 170.000 272.300 ;
        RECT 164.400 271.600 165.200 271.700 ;
        RECT 169.200 271.600 170.000 271.700 ;
        RECT 222.000 272.300 222.800 272.400 ;
        RECT 278.000 272.300 278.800 272.400 ;
        RECT 222.000 271.700 278.800 272.300 ;
        RECT 279.700 272.300 280.300 273.700 ;
        RECT 295.600 273.700 299.600 274.300 ;
        RECT 295.600 273.600 296.400 273.700 ;
        RECT 298.800 273.600 299.600 273.700 ;
        RECT 302.000 274.300 302.800 274.400 ;
        RECT 343.600 274.300 344.400 274.400 ;
        RECT 302.000 273.700 344.400 274.300 ;
        RECT 302.000 273.600 302.800 273.700 ;
        RECT 343.600 273.600 344.400 273.700 ;
        RECT 345.200 274.300 346.000 274.400 ;
        RECT 356.400 274.300 357.200 274.400 ;
        RECT 382.000 274.300 382.800 274.400 ;
        RECT 391.600 274.300 392.400 274.400 ;
        RECT 345.200 273.700 392.400 274.300 ;
        RECT 345.200 273.600 346.000 273.700 ;
        RECT 356.400 273.600 357.200 273.700 ;
        RECT 382.000 273.600 382.800 273.700 ;
        RECT 391.600 273.600 392.400 273.700 ;
        RECT 407.600 274.300 408.400 274.400 ;
        RECT 410.800 274.300 411.600 274.400 ;
        RECT 407.600 273.700 411.600 274.300 ;
        RECT 407.600 273.600 408.400 273.700 ;
        RECT 410.800 273.600 411.600 273.700 ;
        RECT 414.000 274.300 414.800 274.400 ;
        RECT 417.200 274.300 418.000 274.400 ;
        RECT 414.000 273.700 418.000 274.300 ;
        RECT 414.000 273.600 414.800 273.700 ;
        RECT 417.200 273.600 418.000 273.700 ;
        RECT 434.800 274.300 435.600 274.400 ;
        RECT 439.600 274.300 440.400 274.400 ;
        RECT 434.800 273.700 440.400 274.300 ;
        RECT 434.800 273.600 435.600 273.700 ;
        RECT 439.600 273.600 440.400 273.700 ;
        RECT 450.800 274.300 451.600 274.400 ;
        RECT 482.800 274.300 483.600 274.400 ;
        RECT 450.800 273.700 483.600 274.300 ;
        RECT 450.800 273.600 451.600 273.700 ;
        RECT 482.800 273.600 483.600 273.700 ;
        RECT 489.200 274.300 490.000 274.400 ;
        RECT 510.000 274.300 510.800 274.400 ;
        RECT 489.200 273.700 510.800 274.300 ;
        RECT 489.200 273.600 490.000 273.700 ;
        RECT 510.000 273.600 510.800 273.700 ;
        RECT 516.400 274.300 517.200 274.400 ;
        RECT 534.000 274.300 534.800 274.400 ;
        RECT 516.400 273.700 534.800 274.300 ;
        RECT 516.400 273.600 517.200 273.700 ;
        RECT 534.000 273.600 534.800 273.700 ;
        RECT 558.000 274.300 558.800 274.400 ;
        RECT 564.400 274.300 565.200 274.400 ;
        RECT 575.600 274.300 576.400 274.400 ;
        RECT 558.000 273.700 576.400 274.300 ;
        RECT 558.000 273.600 558.800 273.700 ;
        RECT 564.400 273.600 565.200 273.700 ;
        RECT 575.600 273.600 576.400 273.700 ;
        RECT 348.400 272.300 349.200 272.400 ;
        RECT 279.700 271.700 349.200 272.300 ;
        RECT 222.000 271.600 222.800 271.700 ;
        RECT 278.000 271.600 278.800 271.700 ;
        RECT 348.400 271.600 349.200 271.700 ;
        RECT 351.600 272.300 352.400 272.400 ;
        RECT 356.400 272.300 357.200 272.400 ;
        RECT 351.600 271.700 357.200 272.300 ;
        RECT 351.600 271.600 352.400 271.700 ;
        RECT 356.400 271.600 357.200 271.700 ;
        RECT 364.400 272.300 365.200 272.400 ;
        RECT 366.000 272.300 366.800 272.400 ;
        RECT 364.400 271.700 366.800 272.300 ;
        RECT 364.400 271.600 365.200 271.700 ;
        RECT 366.000 271.600 366.800 271.700 ;
        RECT 369.200 272.300 370.000 272.400 ;
        RECT 375.600 272.300 376.400 272.400 ;
        RECT 369.200 271.700 376.400 272.300 ;
        RECT 369.200 271.600 370.000 271.700 ;
        RECT 375.600 271.600 376.400 271.700 ;
        RECT 377.200 272.300 378.000 272.400 ;
        RECT 444.400 272.300 445.200 272.400 ;
        RECT 377.200 271.700 445.200 272.300 ;
        RECT 377.200 271.600 378.000 271.700 ;
        RECT 444.400 271.600 445.200 271.700 ;
        RECT 454.000 272.300 454.800 272.400 ;
        RECT 478.000 272.300 478.800 272.400 ;
        RECT 454.000 271.700 478.800 272.300 ;
        RECT 454.000 271.600 454.800 271.700 ;
        RECT 478.000 271.600 478.800 271.700 ;
        RECT 482.800 272.300 483.600 272.400 ;
        RECT 502.000 272.300 502.800 272.400 ;
        RECT 540.400 272.300 541.200 272.400 ;
        RECT 545.200 272.300 546.000 272.400 ;
        RECT 550.000 272.300 550.800 272.400 ;
        RECT 482.800 271.700 550.800 272.300 ;
        RECT 482.800 271.600 483.600 271.700 ;
        RECT 502.000 271.600 502.800 271.700 ;
        RECT 540.400 271.600 541.200 271.700 ;
        RECT 545.200 271.600 546.000 271.700 ;
        RECT 550.000 271.600 550.800 271.700 ;
        RECT 25.200 270.300 26.000 270.400 ;
        RECT 28.400 270.300 29.200 270.400 ;
        RECT 46.000 270.300 46.800 270.400 ;
        RECT 25.200 269.700 46.800 270.300 ;
        RECT 25.200 269.600 26.000 269.700 ;
        RECT 28.400 269.600 29.200 269.700 ;
        RECT 46.000 269.600 46.800 269.700 ;
        RECT 54.000 270.300 54.800 270.400 ;
        RECT 74.800 270.300 75.600 270.400 ;
        RECT 78.000 270.300 78.800 270.400 ;
        RECT 54.000 269.700 78.800 270.300 ;
        RECT 54.000 269.600 54.800 269.700 ;
        RECT 74.800 269.600 75.600 269.700 ;
        RECT 78.000 269.600 78.800 269.700 ;
        RECT 103.600 270.300 104.400 270.400 ;
        RECT 114.800 270.300 115.600 270.400 ;
        RECT 103.600 269.700 115.600 270.300 ;
        RECT 103.600 269.600 104.400 269.700 ;
        RECT 114.800 269.600 115.600 269.700 ;
        RECT 162.800 270.300 163.600 270.400 ;
        RECT 175.600 270.300 176.400 270.400 ;
        RECT 178.800 270.300 179.600 270.400 ;
        RECT 162.800 269.700 179.600 270.300 ;
        RECT 162.800 269.600 163.600 269.700 ;
        RECT 175.600 269.600 176.400 269.700 ;
        RECT 178.800 269.600 179.600 269.700 ;
        RECT 212.400 270.300 213.200 270.400 ;
        RECT 268.400 270.300 269.200 270.400 ;
        RECT 212.400 269.700 269.200 270.300 ;
        RECT 212.400 269.600 213.200 269.700 ;
        RECT 268.400 269.600 269.200 269.700 ;
        RECT 276.400 270.300 277.200 270.400 ;
        RECT 350.000 270.300 350.800 270.400 ;
        RECT 276.400 269.700 350.800 270.300 ;
        RECT 276.400 269.600 277.200 269.700 ;
        RECT 350.000 269.600 350.800 269.700 ;
        RECT 354.800 270.300 355.600 270.400 ;
        RECT 359.600 270.300 360.400 270.400 ;
        RECT 354.800 269.700 360.400 270.300 ;
        RECT 354.800 269.600 355.600 269.700 ;
        RECT 359.600 269.600 360.400 269.700 ;
        RECT 367.600 270.300 368.400 270.400 ;
        RECT 372.400 270.300 373.200 270.400 ;
        RECT 367.600 269.700 373.200 270.300 ;
        RECT 367.600 269.600 368.400 269.700 ;
        RECT 372.400 269.600 373.200 269.700 ;
        RECT 375.600 270.300 376.400 270.400 ;
        RECT 382.000 270.300 382.800 270.400 ;
        RECT 375.600 269.700 382.800 270.300 ;
        RECT 375.600 269.600 376.400 269.700 ;
        RECT 382.000 269.600 382.800 269.700 ;
        RECT 383.600 270.300 384.400 270.400 ;
        RECT 394.800 270.300 395.600 270.400 ;
        RECT 409.200 270.300 410.000 270.400 ;
        RECT 412.400 270.300 413.200 270.400 ;
        RECT 383.600 269.700 413.200 270.300 ;
        RECT 383.600 269.600 384.400 269.700 ;
        RECT 394.800 269.600 395.600 269.700 ;
        RECT 409.200 269.600 410.000 269.700 ;
        RECT 412.400 269.600 413.200 269.700 ;
        RECT 426.800 270.300 427.600 270.400 ;
        RECT 431.600 270.300 432.400 270.400 ;
        RECT 426.800 269.700 432.400 270.300 ;
        RECT 426.800 269.600 427.600 269.700 ;
        RECT 431.600 269.600 432.400 269.700 ;
        RECT 442.800 270.300 443.600 270.400 ;
        RECT 446.000 270.300 446.800 270.400 ;
        RECT 442.800 269.700 446.800 270.300 ;
        RECT 442.800 269.600 443.600 269.700 ;
        RECT 446.000 269.600 446.800 269.700 ;
        RECT 474.800 270.300 475.600 270.400 ;
        RECT 478.000 270.300 478.800 270.400 ;
        RECT 486.000 270.300 486.800 270.400 ;
        RECT 474.800 269.700 486.800 270.300 ;
        RECT 474.800 269.600 475.600 269.700 ;
        RECT 478.000 269.600 478.800 269.700 ;
        RECT 486.000 269.600 486.800 269.700 ;
        RECT 495.600 270.300 496.400 270.400 ;
        RECT 503.600 270.300 504.400 270.400 ;
        RECT 495.600 269.700 504.400 270.300 ;
        RECT 495.600 269.600 496.400 269.700 ;
        RECT 503.600 269.600 504.400 269.700 ;
        RECT 508.400 270.300 509.200 270.400 ;
        RECT 516.400 270.300 517.200 270.400 ;
        RECT 508.400 269.700 517.200 270.300 ;
        RECT 508.400 269.600 509.200 269.700 ;
        RECT 516.400 269.600 517.200 269.700 ;
        RECT 519.600 270.300 520.400 270.400 ;
        RECT 527.600 270.300 528.400 270.400 ;
        RECT 519.600 269.700 528.400 270.300 ;
        RECT 519.600 269.600 520.400 269.700 ;
        RECT 527.600 269.600 528.400 269.700 ;
        RECT 534.000 270.300 534.800 270.400 ;
        RECT 538.800 270.300 539.600 270.400 ;
        RECT 534.000 269.700 539.600 270.300 ;
        RECT 534.000 269.600 534.800 269.700 ;
        RECT 538.800 269.600 539.600 269.700 ;
        RECT 569.200 270.300 570.000 270.400 ;
        RECT 578.800 270.300 579.600 270.400 ;
        RECT 586.800 270.300 587.600 270.400 ;
        RECT 569.200 269.700 587.600 270.300 ;
        RECT 569.200 269.600 570.000 269.700 ;
        RECT 578.800 269.600 579.600 269.700 ;
        RECT 586.800 269.600 587.600 269.700 ;
        RECT 14.000 268.300 14.800 268.400 ;
        RECT 74.800 268.300 75.600 268.400 ;
        RECT 79.600 268.300 80.400 268.400 ;
        RECT 82.800 268.300 83.600 268.400 ;
        RECT 87.600 268.300 88.400 268.400 ;
        RECT 100.400 268.300 101.200 268.400 ;
        RECT 14.000 267.700 75.600 268.300 ;
        RECT 78.100 267.700 101.200 268.300 ;
        RECT 14.000 267.600 14.800 267.700 ;
        RECT 74.800 267.600 75.600 267.700 ;
        RECT 79.600 267.600 80.400 267.700 ;
        RECT 82.800 267.600 83.600 267.700 ;
        RECT 87.600 267.600 88.400 267.700 ;
        RECT 100.400 267.600 101.200 267.700 ;
        RECT 113.200 268.300 114.000 268.400 ;
        RECT 124.400 268.300 125.200 268.400 ;
        RECT 113.200 267.700 125.200 268.300 ;
        RECT 113.200 267.600 114.000 267.700 ;
        RECT 124.400 267.600 125.200 267.700 ;
        RECT 138.800 267.600 139.600 268.400 ;
        RECT 188.400 268.300 189.200 268.400 ;
        RECT 207.600 268.300 208.400 268.400 ;
        RECT 212.400 268.300 213.200 268.400 ;
        RECT 188.400 267.700 190.700 268.300 ;
        RECT 188.400 267.600 189.200 267.700 ;
        RECT 17.200 266.300 18.000 266.400 ;
        RECT 54.000 266.300 54.800 266.400 ;
        RECT 17.200 265.700 54.800 266.300 ;
        RECT 17.200 265.600 18.000 265.700 ;
        RECT 54.000 265.600 54.800 265.700 ;
        RECT 57.200 266.300 58.000 266.400 ;
        RECT 81.200 266.300 82.000 266.400 ;
        RECT 57.200 265.700 82.000 266.300 ;
        RECT 57.200 265.600 58.000 265.700 ;
        RECT 81.200 265.600 82.000 265.700 ;
        RECT 90.800 266.300 91.600 266.400 ;
        RECT 118.000 266.300 118.800 266.400 ;
        RECT 90.800 265.700 118.800 266.300 ;
        RECT 90.800 265.600 91.600 265.700 ;
        RECT 118.000 265.600 118.800 265.700 ;
        RECT 167.600 266.300 168.400 266.400 ;
        RECT 188.400 266.300 189.200 266.400 ;
        RECT 167.600 265.700 189.200 266.300 ;
        RECT 190.100 266.300 190.700 267.700 ;
        RECT 207.600 267.700 213.200 268.300 ;
        RECT 207.600 267.600 208.400 267.700 ;
        RECT 212.400 267.600 213.200 267.700 ;
        RECT 244.400 268.300 245.200 268.400 ;
        RECT 270.000 268.300 270.800 268.400 ;
        RECT 244.400 267.700 270.800 268.300 ;
        RECT 244.400 267.600 245.200 267.700 ;
        RECT 270.000 267.600 270.800 267.700 ;
        RECT 286.000 267.600 286.800 268.400 ;
        RECT 298.800 268.300 299.600 268.400 ;
        RECT 300.400 268.300 301.200 268.400 ;
        RECT 298.800 267.700 301.200 268.300 ;
        RECT 298.800 267.600 299.600 267.700 ;
        RECT 300.400 267.600 301.200 267.700 ;
        RECT 308.400 268.300 309.200 268.400 ;
        RECT 322.800 268.300 323.600 268.400 ;
        RECT 308.400 267.700 323.600 268.300 ;
        RECT 308.400 267.600 309.200 267.700 ;
        RECT 322.800 267.600 323.600 267.700 ;
        RECT 327.600 268.300 328.400 268.400 ;
        RECT 340.400 268.300 341.200 268.400 ;
        RECT 327.600 267.700 341.200 268.300 ;
        RECT 327.600 267.600 328.400 267.700 ;
        RECT 340.400 267.600 341.200 267.700 ;
        RECT 343.600 268.300 344.400 268.400 ;
        RECT 394.800 268.300 395.600 268.400 ;
        RECT 343.600 267.700 395.600 268.300 ;
        RECT 343.600 267.600 344.400 267.700 ;
        RECT 394.800 267.600 395.600 267.700 ;
        RECT 396.400 268.300 397.200 268.400 ;
        RECT 404.400 268.300 405.200 268.400 ;
        RECT 396.400 267.700 405.200 268.300 ;
        RECT 396.400 267.600 397.200 267.700 ;
        RECT 404.400 267.600 405.200 267.700 ;
        RECT 415.600 268.300 416.400 268.400 ;
        RECT 433.200 268.300 434.000 268.400 ;
        RECT 441.200 268.300 442.000 268.400 ;
        RECT 476.400 268.300 477.200 268.400 ;
        RECT 415.600 267.700 432.300 268.300 ;
        RECT 415.600 267.600 416.400 267.700 ;
        RECT 220.400 266.300 221.200 266.400 ;
        RECT 190.100 265.700 221.200 266.300 ;
        RECT 167.600 265.600 168.400 265.700 ;
        RECT 188.400 265.600 189.200 265.700 ;
        RECT 220.400 265.600 221.200 265.700 ;
        RECT 263.600 266.300 264.400 266.400 ;
        RECT 278.000 266.300 278.800 266.400 ;
        RECT 263.600 265.700 278.800 266.300 ;
        RECT 263.600 265.600 264.400 265.700 ;
        RECT 278.000 265.600 278.800 265.700 ;
        RECT 284.400 266.300 285.200 266.400 ;
        RECT 300.400 266.300 301.200 266.400 ;
        RECT 284.400 265.700 301.200 266.300 ;
        RECT 284.400 265.600 285.200 265.700 ;
        RECT 300.400 265.600 301.200 265.700 ;
        RECT 314.800 266.300 315.600 266.400 ;
        RECT 324.400 266.300 325.200 266.400 ;
        RECT 326.000 266.300 326.800 266.400 ;
        RECT 314.800 265.700 326.800 266.300 ;
        RECT 314.800 265.600 315.600 265.700 ;
        RECT 324.400 265.600 325.200 265.700 ;
        RECT 326.000 265.600 326.800 265.700 ;
        RECT 386.800 266.300 387.600 266.400 ;
        RECT 401.200 266.300 402.000 266.400 ;
        RECT 407.600 266.300 408.400 266.400 ;
        RECT 420.400 266.300 421.200 266.400 ;
        RECT 386.800 265.700 421.200 266.300 ;
        RECT 431.700 266.300 432.300 267.700 ;
        RECT 433.200 267.700 442.000 268.300 ;
        RECT 433.200 267.600 434.000 267.700 ;
        RECT 441.200 267.600 442.000 267.700 ;
        RECT 474.900 267.700 477.200 268.300 ;
        RECT 474.900 266.300 475.500 267.700 ;
        RECT 476.400 267.600 477.200 267.700 ;
        RECT 486.000 268.300 486.800 268.400 ;
        RECT 497.200 268.300 498.000 268.400 ;
        RECT 510.000 268.300 510.800 268.400 ;
        RECT 542.000 268.300 542.800 268.400 ;
        RECT 548.400 268.300 549.200 268.400 ;
        RECT 486.000 267.700 549.200 268.300 ;
        RECT 486.000 267.600 486.800 267.700 ;
        RECT 497.200 267.600 498.000 267.700 ;
        RECT 510.000 267.600 510.800 267.700 ;
        RECT 542.000 267.600 542.800 267.700 ;
        RECT 548.400 267.600 549.200 267.700 ;
        RECT 554.800 268.300 555.600 268.400 ;
        RECT 564.400 268.300 565.200 268.400 ;
        RECT 554.800 267.700 565.200 268.300 ;
        RECT 554.800 267.600 555.600 267.700 ;
        RECT 564.400 267.600 565.200 267.700 ;
        RECT 577.200 268.300 578.000 268.400 ;
        RECT 598.000 268.300 598.800 268.400 ;
        RECT 577.200 267.700 598.800 268.300 ;
        RECT 577.200 267.600 578.000 267.700 ;
        RECT 598.000 267.600 598.800 267.700 ;
        RECT 602.800 268.300 603.600 268.400 ;
        RECT 604.400 268.300 605.200 268.400 ;
        RECT 602.800 267.700 605.200 268.300 ;
        RECT 602.800 267.600 603.600 267.700 ;
        RECT 604.400 267.600 605.200 267.700 ;
        RECT 431.700 265.700 475.500 266.300 ;
        RECT 476.400 266.300 477.200 266.400 ;
        RECT 479.600 266.300 480.400 266.400 ;
        RECT 484.400 266.300 485.200 266.400 ;
        RECT 495.600 266.300 496.400 266.400 ;
        RECT 476.400 265.700 496.400 266.300 ;
        RECT 386.800 265.600 387.600 265.700 ;
        RECT 401.200 265.600 402.000 265.700 ;
        RECT 407.600 265.600 408.400 265.700 ;
        RECT 420.400 265.600 421.200 265.700 ;
        RECT 476.400 265.600 477.200 265.700 ;
        RECT 479.600 265.600 480.400 265.700 ;
        RECT 484.400 265.600 485.200 265.700 ;
        RECT 495.600 265.600 496.400 265.700 ;
        RECT 500.400 266.300 501.200 266.400 ;
        RECT 514.800 266.300 515.600 266.400 ;
        RECT 500.400 265.700 515.600 266.300 ;
        RECT 500.400 265.600 501.200 265.700 ;
        RECT 514.800 265.600 515.600 265.700 ;
        RECT 516.400 266.300 517.200 266.400 ;
        RECT 524.400 266.300 525.200 266.400 ;
        RECT 516.400 265.700 525.200 266.300 ;
        RECT 516.400 265.600 517.200 265.700 ;
        RECT 524.400 265.600 525.200 265.700 ;
        RECT 526.000 266.300 526.800 266.400 ;
        RECT 543.600 266.300 544.400 266.400 ;
        RECT 548.400 266.300 549.200 266.400 ;
        RECT 526.000 265.700 549.200 266.300 ;
        RECT 526.000 265.600 526.800 265.700 ;
        RECT 543.600 265.600 544.400 265.700 ;
        RECT 548.400 265.600 549.200 265.700 ;
        RECT 586.800 266.300 587.600 266.400 ;
        RECT 594.800 266.300 595.600 266.400 ;
        RECT 586.800 265.700 595.600 266.300 ;
        RECT 586.800 265.600 587.600 265.700 ;
        RECT 594.800 265.600 595.600 265.700 ;
        RECT 33.200 264.300 34.000 264.400 ;
        RECT 36.400 264.300 37.200 264.400 ;
        RECT 71.600 264.300 72.400 264.400 ;
        RECT 33.200 263.700 72.400 264.300 ;
        RECT 33.200 263.600 34.000 263.700 ;
        RECT 36.400 263.600 37.200 263.700 ;
        RECT 71.600 263.600 72.400 263.700 ;
        RECT 150.000 264.300 150.800 264.400 ;
        RECT 191.600 264.300 192.400 264.400 ;
        RECT 210.800 264.300 211.600 264.400 ;
        RECT 150.000 263.700 211.600 264.300 ;
        RECT 150.000 263.600 150.800 263.700 ;
        RECT 191.600 263.600 192.400 263.700 ;
        RECT 210.800 263.600 211.600 263.700 ;
        RECT 266.800 264.300 267.600 264.400 ;
        RECT 281.200 264.300 282.000 264.400 ;
        RECT 295.600 264.300 296.400 264.400 ;
        RECT 359.600 264.300 360.400 264.400 ;
        RECT 266.800 263.700 360.400 264.300 ;
        RECT 266.800 263.600 267.600 263.700 ;
        RECT 281.200 263.600 282.000 263.700 ;
        RECT 295.600 263.600 296.400 263.700 ;
        RECT 359.600 263.600 360.400 263.700 ;
        RECT 372.400 264.300 373.200 264.400 ;
        RECT 377.200 264.300 378.000 264.400 ;
        RECT 372.400 263.700 378.000 264.300 ;
        RECT 372.400 263.600 373.200 263.700 ;
        RECT 377.200 263.600 378.000 263.700 ;
        RECT 378.800 264.300 379.600 264.400 ;
        RECT 406.000 264.300 406.800 264.400 ;
        RECT 417.200 264.300 418.000 264.400 ;
        RECT 425.200 264.300 426.000 264.400 ;
        RECT 431.600 264.300 432.400 264.400 ;
        RECT 468.400 264.300 469.200 264.400 ;
        RECT 378.800 263.700 469.200 264.300 ;
        RECT 378.800 263.600 379.600 263.700 ;
        RECT 406.000 263.600 406.800 263.700 ;
        RECT 417.200 263.600 418.000 263.700 ;
        RECT 425.200 263.600 426.000 263.700 ;
        RECT 431.600 263.600 432.400 263.700 ;
        RECT 468.400 263.600 469.200 263.700 ;
        RECT 474.800 264.300 475.600 264.400 ;
        RECT 487.600 264.300 488.400 264.400 ;
        RECT 474.800 263.700 488.400 264.300 ;
        RECT 474.800 263.600 475.600 263.700 ;
        RECT 487.600 263.600 488.400 263.700 ;
        RECT 494.000 264.300 494.800 264.400 ;
        RECT 502.000 264.300 502.800 264.400 ;
        RECT 494.000 263.700 502.800 264.300 ;
        RECT 494.000 263.600 494.800 263.700 ;
        RECT 502.000 263.600 502.800 263.700 ;
        RECT 503.600 264.300 504.400 264.400 ;
        RECT 505.200 264.300 506.000 264.400 ;
        RECT 503.600 263.700 506.000 264.300 ;
        RECT 503.600 263.600 504.400 263.700 ;
        RECT 505.200 263.600 506.000 263.700 ;
        RECT 506.800 264.300 507.600 264.400 ;
        RECT 508.400 264.300 509.200 264.400 ;
        RECT 506.800 263.700 509.200 264.300 ;
        RECT 506.800 263.600 507.600 263.700 ;
        RECT 508.400 263.600 509.200 263.700 ;
        RECT 521.200 264.300 522.000 264.400 ;
        RECT 558.000 264.300 558.800 264.400 ;
        RECT 521.200 263.700 558.800 264.300 ;
        RECT 521.200 263.600 522.000 263.700 ;
        RECT 558.000 263.600 558.800 263.700 ;
        RECT 169.200 262.300 170.000 262.400 ;
        RECT 186.800 262.300 187.600 262.400 ;
        RECT 169.200 261.700 187.600 262.300 ;
        RECT 169.200 261.600 170.000 261.700 ;
        RECT 186.800 261.600 187.600 261.700 ;
        RECT 188.400 262.300 189.200 262.400 ;
        RECT 214.000 262.300 214.800 262.400 ;
        RECT 217.200 262.300 218.000 262.400 ;
        RECT 188.400 261.700 218.000 262.300 ;
        RECT 188.400 261.600 189.200 261.700 ;
        RECT 214.000 261.600 214.800 261.700 ;
        RECT 217.200 261.600 218.000 261.700 ;
        RECT 353.200 262.300 354.000 262.400 ;
        RECT 366.000 262.300 366.800 262.400 ;
        RECT 353.200 261.700 366.800 262.300 ;
        RECT 353.200 261.600 354.000 261.700 ;
        RECT 366.000 261.600 366.800 261.700 ;
        RECT 367.600 262.300 368.400 262.400 ;
        RECT 386.800 262.300 387.600 262.400 ;
        RECT 417.200 262.300 418.000 262.400 ;
        RECT 367.600 261.700 387.600 262.300 ;
        RECT 367.600 261.600 368.400 261.700 ;
        RECT 386.800 261.600 387.600 261.700 ;
        RECT 388.500 261.700 418.000 262.300 ;
        RECT 114.800 260.300 115.600 260.400 ;
        RECT 119.600 260.300 120.400 260.400 ;
        RECT 114.800 259.700 120.400 260.300 ;
        RECT 114.800 259.600 115.600 259.700 ;
        RECT 119.600 259.600 120.400 259.700 ;
        RECT 166.000 260.300 166.800 260.400 ;
        RECT 185.200 260.300 186.000 260.400 ;
        RECT 166.000 259.700 186.000 260.300 ;
        RECT 166.000 259.600 166.800 259.700 ;
        RECT 185.200 259.600 186.000 259.700 ;
        RECT 193.200 260.300 194.000 260.400 ;
        RECT 199.600 260.300 200.400 260.400 ;
        RECT 193.200 259.700 200.400 260.300 ;
        RECT 193.200 259.600 194.000 259.700 ;
        RECT 199.600 259.600 200.400 259.700 ;
        RECT 350.000 260.300 350.800 260.400 ;
        RECT 362.800 260.300 363.600 260.400 ;
        RECT 350.000 259.700 363.600 260.300 ;
        RECT 350.000 259.600 350.800 259.700 ;
        RECT 362.800 259.600 363.600 259.700 ;
        RECT 367.600 260.300 368.400 260.400 ;
        RECT 388.500 260.300 389.100 261.700 ;
        RECT 417.200 261.600 418.000 261.700 ;
        RECT 426.800 262.300 427.600 262.400 ;
        RECT 430.000 262.300 430.800 262.400 ;
        RECT 426.800 261.700 430.800 262.300 ;
        RECT 426.800 261.600 427.600 261.700 ;
        RECT 430.000 261.600 430.800 261.700 ;
        RECT 433.200 262.300 434.000 262.400 ;
        RECT 463.600 262.300 464.400 262.400 ;
        RECT 433.200 261.700 464.400 262.300 ;
        RECT 433.200 261.600 434.000 261.700 ;
        RECT 463.600 261.600 464.400 261.700 ;
        RECT 471.600 262.300 472.400 262.400 ;
        RECT 478.000 262.300 478.800 262.400 ;
        RECT 471.600 261.700 478.800 262.300 ;
        RECT 471.600 261.600 472.400 261.700 ;
        RECT 478.000 261.600 478.800 261.700 ;
        RECT 484.400 262.300 485.200 262.400 ;
        RECT 495.600 262.300 496.400 262.400 ;
        RECT 484.400 261.700 496.400 262.300 ;
        RECT 484.400 261.600 485.200 261.700 ;
        RECT 495.600 261.600 496.400 261.700 ;
        RECT 502.000 262.300 502.800 262.400 ;
        RECT 519.600 262.300 520.400 262.400 ;
        RECT 502.000 261.700 520.400 262.300 ;
        RECT 502.000 261.600 502.800 261.700 ;
        RECT 519.600 261.600 520.400 261.700 ;
        RECT 535.600 262.300 536.400 262.400 ;
        RECT 542.000 262.300 542.800 262.400 ;
        RECT 535.600 261.700 542.800 262.300 ;
        RECT 535.600 261.600 536.400 261.700 ;
        RECT 542.000 261.600 542.800 261.700 ;
        RECT 367.600 259.700 389.100 260.300 ;
        RECT 402.800 260.300 403.600 260.400 ;
        RECT 414.000 260.300 414.800 260.400 ;
        RECT 402.800 259.700 414.800 260.300 ;
        RECT 367.600 259.600 368.400 259.700 ;
        RECT 402.800 259.600 403.600 259.700 ;
        RECT 414.000 259.600 414.800 259.700 ;
        RECT 415.600 260.300 416.400 260.400 ;
        RECT 420.400 260.300 421.200 260.400 ;
        RECT 428.400 260.300 429.200 260.400 ;
        RECT 441.200 260.300 442.000 260.400 ;
        RECT 415.600 259.700 442.000 260.300 ;
        RECT 415.600 259.600 416.400 259.700 ;
        RECT 420.400 259.600 421.200 259.700 ;
        RECT 428.400 259.600 429.200 259.700 ;
        RECT 441.200 259.600 442.000 259.700 ;
        RECT 454.000 260.300 454.800 260.400 ;
        RECT 465.200 260.300 466.000 260.400 ;
        RECT 478.000 260.300 478.800 260.400 ;
        RECT 500.400 260.300 501.200 260.400 ;
        RECT 454.000 259.700 501.200 260.300 ;
        RECT 454.000 259.600 454.800 259.700 ;
        RECT 465.200 259.600 466.000 259.700 ;
        RECT 478.000 259.600 478.800 259.700 ;
        RECT 500.400 259.600 501.200 259.700 ;
        RECT 503.600 260.300 504.400 260.400 ;
        RECT 514.800 260.300 515.600 260.400 ;
        RECT 503.600 259.700 515.600 260.300 ;
        RECT 503.600 259.600 504.400 259.700 ;
        RECT 514.800 259.600 515.600 259.700 ;
        RECT 522.800 260.300 523.600 260.400 ;
        RECT 530.800 260.300 531.600 260.400 ;
        RECT 522.800 259.700 531.600 260.300 ;
        RECT 522.800 259.600 523.600 259.700 ;
        RECT 530.800 259.600 531.600 259.700 ;
        RECT 546.800 260.300 547.600 260.400 ;
        RECT 577.200 260.300 578.000 260.400 ;
        RECT 546.800 259.700 578.000 260.300 ;
        RECT 546.800 259.600 547.600 259.700 ;
        RECT 577.200 259.600 578.000 259.700 ;
        RECT 242.800 258.300 243.600 258.400 ;
        RECT 266.800 258.300 267.600 258.400 ;
        RECT 242.800 257.700 267.600 258.300 ;
        RECT 242.800 257.600 243.600 257.700 ;
        RECT 266.800 257.600 267.600 257.700 ;
        RECT 270.000 258.300 270.800 258.400 ;
        RECT 286.000 258.300 286.800 258.400 ;
        RECT 270.000 257.700 286.800 258.300 ;
        RECT 270.000 257.600 270.800 257.700 ;
        RECT 286.000 257.600 286.800 257.700 ;
        RECT 290.800 258.300 291.600 258.400 ;
        RECT 318.000 258.300 318.800 258.400 ;
        RECT 390.000 258.300 390.800 258.400 ;
        RECT 290.800 257.700 317.100 258.300 ;
        RECT 290.800 257.600 291.600 257.700 ;
        RECT 38.000 256.300 38.800 256.400 ;
        RECT 74.800 256.300 75.600 256.400 ;
        RECT 38.000 255.700 75.600 256.300 ;
        RECT 38.000 255.600 38.800 255.700 ;
        RECT 74.800 255.600 75.600 255.700 ;
        RECT 100.400 256.300 101.200 256.400 ;
        RECT 111.600 256.300 112.400 256.400 ;
        RECT 126.000 256.300 126.800 256.400 ;
        RECT 161.200 256.300 162.000 256.400 ;
        RECT 100.400 255.700 162.000 256.300 ;
        RECT 100.400 255.600 101.200 255.700 ;
        RECT 111.600 255.600 112.400 255.700 ;
        RECT 126.000 255.600 126.800 255.700 ;
        RECT 161.200 255.600 162.000 255.700 ;
        RECT 247.600 256.300 248.400 256.400 ;
        RECT 260.400 256.300 261.200 256.400 ;
        RECT 266.800 256.300 267.600 256.400 ;
        RECT 247.600 255.700 267.600 256.300 ;
        RECT 247.600 255.600 248.400 255.700 ;
        RECT 260.400 255.600 261.200 255.700 ;
        RECT 266.800 255.600 267.600 255.700 ;
        RECT 284.400 256.300 285.200 256.400 ;
        RECT 287.600 256.300 288.400 256.400 ;
        RECT 313.200 256.300 314.000 256.400 ;
        RECT 284.400 255.700 314.000 256.300 ;
        RECT 316.500 256.300 317.100 257.700 ;
        RECT 318.000 257.700 390.800 258.300 ;
        RECT 318.000 257.600 318.800 257.700 ;
        RECT 390.000 257.600 390.800 257.700 ;
        RECT 391.600 258.300 392.400 258.400 ;
        RECT 466.800 258.300 467.600 258.400 ;
        RECT 391.600 257.700 467.600 258.300 ;
        RECT 391.600 257.600 392.400 257.700 ;
        RECT 466.800 257.600 467.600 257.700 ;
        RECT 471.600 258.300 472.400 258.400 ;
        RECT 492.400 258.300 493.200 258.400 ;
        RECT 471.600 257.700 493.200 258.300 ;
        RECT 471.600 257.600 472.400 257.700 ;
        RECT 492.400 257.600 493.200 257.700 ;
        RECT 502.000 258.300 502.800 258.400 ;
        RECT 506.800 258.300 507.600 258.400 ;
        RECT 502.000 257.700 507.600 258.300 ;
        RECT 502.000 257.600 502.800 257.700 ;
        RECT 506.800 257.600 507.600 257.700 ;
        RECT 511.600 258.300 512.400 258.400 ;
        RECT 518.000 258.300 518.800 258.400 ;
        RECT 529.200 258.300 530.000 258.400 ;
        RECT 546.800 258.300 547.600 258.400 ;
        RECT 511.600 257.700 547.600 258.300 ;
        RECT 511.600 257.600 512.400 257.700 ;
        RECT 518.000 257.600 518.800 257.700 ;
        RECT 529.200 257.600 530.000 257.700 ;
        RECT 546.800 257.600 547.600 257.700 ;
        RECT 561.200 258.300 562.000 258.400 ;
        RECT 570.800 258.300 571.600 258.400 ;
        RECT 561.200 257.700 571.600 258.300 ;
        RECT 561.200 257.600 562.000 257.700 ;
        RECT 570.800 257.600 571.600 257.700 ;
        RECT 327.600 256.300 328.400 256.400 ;
        RECT 337.200 256.300 338.000 256.400 ;
        RECT 316.500 255.700 338.000 256.300 ;
        RECT 284.400 255.600 285.200 255.700 ;
        RECT 287.600 255.600 288.400 255.700 ;
        RECT 313.200 255.600 314.000 255.700 ;
        RECT 327.600 255.600 328.400 255.700 ;
        RECT 337.200 255.600 338.000 255.700 ;
        RECT 338.800 256.300 339.600 256.400 ;
        RECT 350.000 256.300 350.800 256.400 ;
        RECT 375.600 256.300 376.400 256.400 ;
        RECT 338.800 255.700 376.400 256.300 ;
        RECT 338.800 255.600 339.600 255.700 ;
        RECT 350.000 255.600 350.800 255.700 ;
        RECT 375.600 255.600 376.400 255.700 ;
        RECT 398.000 256.300 398.800 256.400 ;
        RECT 406.000 256.300 406.800 256.400 ;
        RECT 398.000 255.700 406.800 256.300 ;
        RECT 398.000 255.600 398.800 255.700 ;
        RECT 406.000 255.600 406.800 255.700 ;
        RECT 418.800 256.300 419.600 256.400 ;
        RECT 423.600 256.300 424.400 256.400 ;
        RECT 418.800 255.700 424.400 256.300 ;
        RECT 418.800 255.600 419.600 255.700 ;
        RECT 423.600 255.600 424.400 255.700 ;
        RECT 430.000 256.300 430.800 256.400 ;
        RECT 436.400 256.300 437.200 256.400 ;
        RECT 430.000 255.700 437.200 256.300 ;
        RECT 430.000 255.600 430.800 255.700 ;
        RECT 436.400 255.600 437.200 255.700 ;
        RECT 441.200 256.300 442.000 256.400 ;
        RECT 450.800 256.300 451.600 256.400 ;
        RECT 441.200 255.700 451.600 256.300 ;
        RECT 441.200 255.600 442.000 255.700 ;
        RECT 450.800 255.600 451.600 255.700 ;
        RECT 479.600 256.300 480.400 256.400 ;
        RECT 482.800 256.300 483.600 256.400 ;
        RECT 489.200 256.300 490.000 256.400 ;
        RECT 479.600 255.700 483.600 256.300 ;
        RECT 479.600 255.600 480.400 255.700 ;
        RECT 482.800 255.600 483.600 255.700 ;
        RECT 484.500 255.700 490.000 256.300 ;
        RECT 164.400 254.300 165.200 254.400 ;
        RECT 182.000 254.300 182.800 254.400 ;
        RECT 164.400 253.700 182.800 254.300 ;
        RECT 164.400 253.600 165.200 253.700 ;
        RECT 182.000 253.600 182.800 253.700 ;
        RECT 207.600 254.300 208.400 254.400 ;
        RECT 233.200 254.300 234.000 254.400 ;
        RECT 207.600 253.700 234.000 254.300 ;
        RECT 207.600 253.600 208.400 253.700 ;
        RECT 233.200 253.600 234.000 253.700 ;
        RECT 236.400 254.300 237.200 254.400 ;
        RECT 239.600 254.300 240.400 254.400 ;
        RECT 236.400 253.700 240.400 254.300 ;
        RECT 236.400 253.600 237.200 253.700 ;
        RECT 239.600 253.600 240.400 253.700 ;
        RECT 273.200 254.300 274.000 254.400 ;
        RECT 290.800 254.300 291.600 254.400 ;
        RECT 273.200 253.700 291.600 254.300 ;
        RECT 273.200 253.600 274.000 253.700 ;
        RECT 290.800 253.600 291.600 253.700 ;
        RECT 295.600 254.300 296.400 254.400 ;
        RECT 303.600 254.300 304.400 254.400 ;
        RECT 295.600 253.700 304.400 254.300 ;
        RECT 295.600 253.600 296.400 253.700 ;
        RECT 303.600 253.600 304.400 253.700 ;
        RECT 308.400 254.300 309.200 254.400 ;
        RECT 314.800 254.300 315.600 254.400 ;
        RECT 308.400 253.700 315.600 254.300 ;
        RECT 308.400 253.600 309.200 253.700 ;
        RECT 314.800 253.600 315.600 253.700 ;
        RECT 342.000 254.300 342.800 254.400 ;
        RECT 346.800 254.300 347.600 254.400 ;
        RECT 366.000 254.300 366.800 254.400 ;
        RECT 342.000 253.700 366.800 254.300 ;
        RECT 342.000 253.600 342.800 253.700 ;
        RECT 346.800 253.600 347.600 253.700 ;
        RECT 366.000 253.600 366.800 253.700 ;
        RECT 414.000 254.300 414.800 254.400 ;
        RECT 426.800 254.300 427.600 254.400 ;
        RECT 414.000 253.700 427.600 254.300 ;
        RECT 414.000 253.600 414.800 253.700 ;
        RECT 426.800 253.600 427.600 253.700 ;
        RECT 439.600 254.300 440.400 254.400 ;
        RECT 447.600 254.300 448.400 254.400 ;
        RECT 439.600 253.700 448.400 254.300 ;
        RECT 439.600 253.600 440.400 253.700 ;
        RECT 447.600 253.600 448.400 253.700 ;
        RECT 452.400 254.300 453.200 254.400 ;
        RECT 455.600 254.300 456.400 254.400 ;
        RECT 452.400 253.700 456.400 254.300 ;
        RECT 452.400 253.600 453.200 253.700 ;
        RECT 455.600 253.600 456.400 253.700 ;
        RECT 457.200 254.300 458.000 254.400 ;
        RECT 470.000 254.300 470.800 254.400 ;
        RECT 484.500 254.300 485.100 255.700 ;
        RECT 489.200 255.600 490.000 255.700 ;
        RECT 505.200 256.300 506.000 256.400 ;
        RECT 510.000 256.300 510.800 256.400 ;
        RECT 529.200 256.300 530.000 256.400 ;
        RECT 534.000 256.300 534.800 256.400 ;
        RECT 505.200 255.700 534.800 256.300 ;
        RECT 505.200 255.600 506.000 255.700 ;
        RECT 510.000 255.600 510.800 255.700 ;
        RECT 529.200 255.600 530.000 255.700 ;
        RECT 534.000 255.600 534.800 255.700 ;
        RECT 535.600 256.300 536.400 256.400 ;
        RECT 542.000 256.300 542.800 256.400 ;
        RECT 545.200 256.300 546.000 256.400 ;
        RECT 535.600 255.700 546.000 256.300 ;
        RECT 535.600 255.600 536.400 255.700 ;
        RECT 542.000 255.600 542.800 255.700 ;
        RECT 545.200 255.600 546.000 255.700 ;
        RECT 457.200 253.700 485.100 254.300 ;
        RECT 487.600 254.300 488.400 254.400 ;
        RECT 489.200 254.300 490.000 254.400 ;
        RECT 497.200 254.300 498.000 254.400 ;
        RECT 526.000 254.300 526.800 254.400 ;
        RECT 487.600 253.700 526.800 254.300 ;
        RECT 457.200 253.600 458.000 253.700 ;
        RECT 470.000 253.600 470.800 253.700 ;
        RECT 487.600 253.600 488.400 253.700 ;
        RECT 489.200 253.600 490.000 253.700 ;
        RECT 497.200 253.600 498.000 253.700 ;
        RECT 526.000 253.600 526.800 253.700 ;
        RECT 532.400 254.300 533.200 254.400 ;
        RECT 537.200 254.300 538.000 254.400 ;
        RECT 532.400 253.700 538.000 254.300 ;
        RECT 532.400 253.600 533.200 253.700 ;
        RECT 537.200 253.600 538.000 253.700 ;
        RECT 564.400 254.300 565.200 254.400 ;
        RECT 590.000 254.300 590.800 254.400 ;
        RECT 564.400 253.700 590.800 254.300 ;
        RECT 564.400 253.600 565.200 253.700 ;
        RECT 590.000 253.600 590.800 253.700 ;
        RECT 25.200 252.300 26.000 252.400 ;
        RECT 41.200 252.300 42.000 252.400 ;
        RECT 25.200 251.700 42.000 252.300 ;
        RECT 25.200 251.600 26.000 251.700 ;
        RECT 41.200 251.600 42.000 251.700 ;
        RECT 63.600 252.300 64.400 252.400 ;
        RECT 68.400 252.300 69.200 252.400 ;
        RECT 63.600 251.700 69.200 252.300 ;
        RECT 63.600 251.600 64.400 251.700 ;
        RECT 68.400 251.600 69.200 251.700 ;
        RECT 124.400 252.300 125.200 252.400 ;
        RECT 130.800 252.300 131.600 252.400 ;
        RECT 124.400 251.700 131.600 252.300 ;
        RECT 124.400 251.600 125.200 251.700 ;
        RECT 130.800 251.600 131.600 251.700 ;
        RECT 137.200 252.300 138.000 252.400 ;
        RECT 153.200 252.300 154.000 252.400 ;
        RECT 225.200 252.300 226.000 252.400 ;
        RECT 247.600 252.300 248.400 252.400 ;
        RECT 137.200 251.700 248.400 252.300 ;
        RECT 137.200 251.600 138.000 251.700 ;
        RECT 153.200 251.600 154.000 251.700 ;
        RECT 225.200 251.600 226.000 251.700 ;
        RECT 247.600 251.600 248.400 251.700 ;
        RECT 297.200 252.300 298.000 252.400 ;
        RECT 308.500 252.300 309.100 253.600 ;
        RECT 297.200 251.700 309.100 252.300 ;
        RECT 319.600 252.300 320.400 252.400 ;
        RECT 321.200 252.300 322.000 252.400 ;
        RECT 346.800 252.300 347.600 252.400 ;
        RECT 319.600 251.700 347.600 252.300 ;
        RECT 297.200 251.600 298.000 251.700 ;
        RECT 319.600 251.600 320.400 251.700 ;
        RECT 321.200 251.600 322.000 251.700 ;
        RECT 346.800 251.600 347.600 251.700 ;
        RECT 399.600 252.300 400.400 252.400 ;
        RECT 404.400 252.300 405.200 252.400 ;
        RECT 399.600 251.700 405.200 252.300 ;
        RECT 399.600 251.600 400.400 251.700 ;
        RECT 404.400 251.600 405.200 251.700 ;
        RECT 407.600 252.300 408.400 252.400 ;
        RECT 420.400 252.300 421.200 252.400 ;
        RECT 407.600 251.700 421.200 252.300 ;
        RECT 407.600 251.600 408.400 251.700 ;
        RECT 420.400 251.600 421.200 251.700 ;
        RECT 423.600 252.300 424.400 252.400 ;
        RECT 452.400 252.300 453.200 252.400 ;
        RECT 423.600 251.700 453.200 252.300 ;
        RECT 423.600 251.600 424.400 251.700 ;
        RECT 452.400 251.600 453.200 251.700 ;
        RECT 458.800 252.300 459.600 252.400 ;
        RECT 471.600 252.300 472.400 252.400 ;
        RECT 458.800 251.700 472.400 252.300 ;
        RECT 458.800 251.600 459.600 251.700 ;
        RECT 471.600 251.600 472.400 251.700 ;
        RECT 484.400 252.300 485.200 252.400 ;
        RECT 508.400 252.300 509.200 252.400 ;
        RECT 484.400 251.700 509.200 252.300 ;
        RECT 484.400 251.600 485.200 251.700 ;
        RECT 508.400 251.600 509.200 251.700 ;
        RECT 510.000 252.300 510.800 252.400 ;
        RECT 511.600 252.300 512.400 252.400 ;
        RECT 518.000 252.300 518.800 252.400 ;
        RECT 510.000 251.700 518.800 252.300 ;
        RECT 510.000 251.600 510.800 251.700 ;
        RECT 511.600 251.600 512.400 251.700 ;
        RECT 518.000 251.600 518.800 251.700 ;
        RECT 519.600 252.300 520.400 252.400 ;
        RECT 527.600 252.300 528.400 252.400 ;
        RECT 538.800 252.300 539.600 252.400 ;
        RECT 519.600 251.700 539.600 252.300 ;
        RECT 519.600 251.600 520.400 251.700 ;
        RECT 527.600 251.600 528.400 251.700 ;
        RECT 538.800 251.600 539.600 251.700 ;
        RECT 286.000 249.600 286.800 250.400 ;
        RECT 314.800 250.300 315.600 250.400 ;
        RECT 318.000 250.300 318.800 250.400 ;
        RECT 314.800 249.700 318.800 250.300 ;
        RECT 314.800 249.600 315.600 249.700 ;
        RECT 318.000 249.600 318.800 249.700 ;
        RECT 324.400 250.300 325.200 250.400 ;
        RECT 343.600 250.300 344.400 250.400 ;
        RECT 324.400 249.700 344.400 250.300 ;
        RECT 324.400 249.600 325.200 249.700 ;
        RECT 343.600 249.600 344.400 249.700 ;
        RECT 414.000 250.300 414.800 250.400 ;
        RECT 417.200 250.300 418.000 250.400 ;
        RECT 414.000 249.700 418.000 250.300 ;
        RECT 414.000 249.600 414.800 249.700 ;
        RECT 417.200 249.600 418.000 249.700 ;
        RECT 420.400 250.300 421.200 250.400 ;
        RECT 423.600 250.300 424.400 250.400 ;
        RECT 428.400 250.300 429.200 250.400 ;
        RECT 420.400 249.700 429.200 250.300 ;
        RECT 420.400 249.600 421.200 249.700 ;
        RECT 423.600 249.600 424.400 249.700 ;
        RECT 428.400 249.600 429.200 249.700 ;
        RECT 433.200 250.300 434.000 250.400 ;
        RECT 439.600 250.300 440.400 250.400 ;
        RECT 452.400 250.300 453.200 250.400 ;
        RECT 433.200 249.700 453.200 250.300 ;
        RECT 433.200 249.600 434.000 249.700 ;
        RECT 439.600 249.600 440.400 249.700 ;
        RECT 452.400 249.600 453.200 249.700 ;
        RECT 455.600 250.300 456.400 250.400 ;
        RECT 465.200 250.300 466.000 250.400 ;
        RECT 455.600 249.700 466.000 250.300 ;
        RECT 455.600 249.600 456.400 249.700 ;
        RECT 465.200 249.600 466.000 249.700 ;
        RECT 482.800 250.300 483.600 250.400 ;
        RECT 484.400 250.300 485.200 250.400 ;
        RECT 482.800 249.700 485.200 250.300 ;
        RECT 482.800 249.600 483.600 249.700 ;
        RECT 484.400 249.600 485.200 249.700 ;
        RECT 495.600 250.300 496.400 250.400 ;
        RECT 502.000 250.300 502.800 250.400 ;
        RECT 495.600 249.700 502.800 250.300 ;
        RECT 495.600 249.600 496.400 249.700 ;
        RECT 502.000 249.600 502.800 249.700 ;
        RECT 516.400 250.300 517.200 250.400 ;
        RECT 538.800 250.300 539.600 250.400 ;
        RECT 516.400 249.700 539.600 250.300 ;
        RECT 516.400 249.600 517.200 249.700 ;
        RECT 538.800 249.600 539.600 249.700 ;
        RECT 244.400 248.300 245.200 248.400 ;
        RECT 258.800 248.300 259.600 248.400 ;
        RECT 244.400 247.700 259.600 248.300 ;
        RECT 244.400 247.600 245.200 247.700 ;
        RECT 258.800 247.600 259.600 247.700 ;
        RECT 316.400 248.300 317.200 248.400 ;
        RECT 319.600 248.300 320.400 248.400 ;
        RECT 316.400 247.700 320.400 248.300 ;
        RECT 316.400 247.600 317.200 247.700 ;
        RECT 319.600 247.600 320.400 247.700 ;
        RECT 324.400 248.300 325.200 248.400 ;
        RECT 329.200 248.300 330.000 248.400 ;
        RECT 324.400 247.700 330.000 248.300 ;
        RECT 324.400 247.600 325.200 247.700 ;
        RECT 329.200 247.600 330.000 247.700 ;
        RECT 337.200 248.300 338.000 248.400 ;
        RECT 345.200 248.300 346.000 248.400 ;
        RECT 337.200 247.700 346.000 248.300 ;
        RECT 337.200 247.600 338.000 247.700 ;
        RECT 345.200 247.600 346.000 247.700 ;
        RECT 346.800 248.300 347.600 248.400 ;
        RECT 465.200 248.300 466.000 248.400 ;
        RECT 346.800 247.700 466.000 248.300 ;
        RECT 346.800 247.600 347.600 247.700 ;
        RECT 465.200 247.600 466.000 247.700 ;
        RECT 466.800 248.300 467.600 248.400 ;
        RECT 561.200 248.300 562.000 248.400 ;
        RECT 466.800 247.700 562.000 248.300 ;
        RECT 466.800 247.600 467.600 247.700 ;
        RECT 561.200 247.600 562.000 247.700 ;
        RECT 300.400 246.300 301.200 246.400 ;
        RECT 314.800 246.300 315.600 246.400 ;
        RECT 300.400 245.700 315.600 246.300 ;
        RECT 300.400 245.600 301.200 245.700 ;
        RECT 314.800 245.600 315.600 245.700 ;
        RECT 316.400 246.300 317.200 246.400 ;
        RECT 346.800 246.300 347.600 246.400 ;
        RECT 316.400 245.700 347.600 246.300 ;
        RECT 316.400 245.600 317.200 245.700 ;
        RECT 346.800 245.600 347.600 245.700 ;
        RECT 401.200 246.300 402.000 246.400 ;
        RECT 409.200 246.300 410.000 246.400 ;
        RECT 447.600 246.300 448.400 246.400 ;
        RECT 401.200 245.700 448.400 246.300 ;
        RECT 401.200 245.600 402.000 245.700 ;
        RECT 409.200 245.600 410.000 245.700 ;
        RECT 447.600 245.600 448.400 245.700 ;
        RECT 452.400 246.300 453.200 246.400 ;
        RECT 484.400 246.300 485.200 246.400 ;
        RECT 452.400 245.700 485.200 246.300 ;
        RECT 452.400 245.600 453.200 245.700 ;
        RECT 484.400 245.600 485.200 245.700 ;
        RECT 500.400 246.300 501.200 246.400 ;
        RECT 505.200 246.300 506.000 246.400 ;
        RECT 500.400 245.700 506.000 246.300 ;
        RECT 500.400 245.600 501.200 245.700 ;
        RECT 505.200 245.600 506.000 245.700 ;
        RECT 510.000 246.300 510.800 246.400 ;
        RECT 545.200 246.300 546.000 246.400 ;
        RECT 510.000 245.700 546.000 246.300 ;
        RECT 510.000 245.600 510.800 245.700 ;
        RECT 545.200 245.600 546.000 245.700 ;
        RECT 50.800 244.300 51.600 244.400 ;
        RECT 95.600 244.300 96.400 244.400 ;
        RECT 50.800 243.700 96.400 244.300 ;
        RECT 50.800 243.600 51.600 243.700 ;
        RECT 95.600 243.600 96.400 243.700 ;
        RECT 135.600 244.300 136.400 244.400 ;
        RECT 145.200 244.300 146.000 244.400 ;
        RECT 178.800 244.300 179.600 244.400 ;
        RECT 135.600 243.700 179.600 244.300 ;
        RECT 135.600 243.600 136.400 243.700 ;
        RECT 145.200 243.600 146.000 243.700 ;
        RECT 178.800 243.600 179.600 243.700 ;
        RECT 241.200 244.300 242.000 244.400 ;
        RECT 250.800 244.300 251.600 244.400 ;
        RECT 292.400 244.300 293.200 244.400 ;
        RECT 241.200 243.700 293.200 244.300 ;
        RECT 241.200 243.600 242.000 243.700 ;
        RECT 250.800 243.600 251.600 243.700 ;
        RECT 292.400 243.600 293.200 243.700 ;
        RECT 310.000 244.300 310.800 244.400 ;
        RECT 321.200 244.300 322.000 244.400 ;
        RECT 310.000 243.700 322.000 244.300 ;
        RECT 310.000 243.600 310.800 243.700 ;
        RECT 321.200 243.600 322.000 243.700 ;
        RECT 324.400 244.300 325.200 244.400 ;
        RECT 326.000 244.300 326.800 244.400 ;
        RECT 324.400 243.700 326.800 244.300 ;
        RECT 324.400 243.600 325.200 243.700 ;
        RECT 326.000 243.600 326.800 243.700 ;
        RECT 345.200 244.300 346.000 244.400 ;
        RECT 406.000 244.300 406.800 244.400 ;
        RECT 345.200 243.700 406.800 244.300 ;
        RECT 345.200 243.600 346.000 243.700 ;
        RECT 406.000 243.600 406.800 243.700 ;
        RECT 410.800 244.300 411.600 244.400 ;
        RECT 422.000 244.300 422.800 244.400 ;
        RECT 410.800 243.700 422.800 244.300 ;
        RECT 410.800 243.600 411.600 243.700 ;
        RECT 422.000 243.600 422.800 243.700 ;
        RECT 423.600 244.300 424.400 244.400 ;
        RECT 465.200 244.300 466.000 244.400 ;
        RECT 423.600 243.700 466.000 244.300 ;
        RECT 423.600 243.600 424.400 243.700 ;
        RECT 465.200 243.600 466.000 243.700 ;
        RECT 490.800 244.300 491.600 244.400 ;
        RECT 503.600 244.300 504.400 244.400 ;
        RECT 535.600 244.300 536.400 244.400 ;
        RECT 490.800 243.700 536.400 244.300 ;
        RECT 490.800 243.600 491.600 243.700 ;
        RECT 503.600 243.600 504.400 243.700 ;
        RECT 535.600 243.600 536.400 243.700 ;
        RECT 538.800 244.300 539.600 244.400 ;
        RECT 551.600 244.300 552.400 244.400 ;
        RECT 538.800 243.700 552.400 244.300 ;
        RECT 538.800 243.600 539.600 243.700 ;
        RECT 551.600 243.600 552.400 243.700 ;
        RECT 36.400 242.300 37.200 242.400 ;
        RECT 71.600 242.300 72.400 242.400 ;
        RECT 78.000 242.300 78.800 242.400 ;
        RECT 36.400 241.700 78.800 242.300 ;
        RECT 36.400 241.600 37.200 241.700 ;
        RECT 71.600 241.600 72.400 241.700 ;
        RECT 78.000 241.600 78.800 241.700 ;
        RECT 162.800 242.300 163.600 242.400 ;
        RECT 182.000 242.300 182.800 242.400 ;
        RECT 186.800 242.300 187.600 242.400 ;
        RECT 162.800 241.700 187.600 242.300 ;
        RECT 162.800 241.600 163.600 241.700 ;
        RECT 182.000 241.600 182.800 241.700 ;
        RECT 186.800 241.600 187.600 241.700 ;
        RECT 220.400 242.300 221.200 242.400 ;
        RECT 353.200 242.300 354.000 242.400 ;
        RECT 410.800 242.300 411.600 242.400 ;
        RECT 220.400 241.700 411.600 242.300 ;
        RECT 220.400 241.600 221.200 241.700 ;
        RECT 353.200 241.600 354.000 241.700 ;
        RECT 410.800 241.600 411.600 241.700 ;
        RECT 417.200 242.300 418.000 242.400 ;
        RECT 418.800 242.300 419.600 242.400 ;
        RECT 417.200 241.700 419.600 242.300 ;
        RECT 417.200 241.600 418.000 241.700 ;
        RECT 418.800 241.600 419.600 241.700 ;
        RECT 463.600 242.300 464.400 242.400 ;
        RECT 468.400 242.300 469.200 242.400 ;
        RECT 463.600 241.700 469.200 242.300 ;
        RECT 463.600 241.600 464.400 241.700 ;
        RECT 468.400 241.600 469.200 241.700 ;
        RECT 471.600 242.300 472.400 242.400 ;
        RECT 481.200 242.300 482.000 242.400 ;
        RECT 471.600 241.700 482.000 242.300 ;
        RECT 471.600 241.600 472.400 241.700 ;
        RECT 481.200 241.600 482.000 241.700 ;
        RECT 482.800 242.300 483.600 242.400 ;
        RECT 500.400 242.300 501.200 242.400 ;
        RECT 482.800 241.700 501.200 242.300 ;
        RECT 482.800 241.600 483.600 241.700 ;
        RECT 500.400 241.600 501.200 241.700 ;
        RECT 503.600 242.300 504.400 242.400 ;
        RECT 537.200 242.300 538.000 242.400 ;
        RECT 503.600 241.700 538.000 242.300 ;
        RECT 503.600 241.600 504.400 241.700 ;
        RECT 537.200 241.600 538.000 241.700 ;
        RECT 22.000 240.300 22.800 240.400 ;
        RECT 52.400 240.300 53.200 240.400 ;
        RECT 22.000 239.700 53.200 240.300 ;
        RECT 22.000 239.600 22.800 239.700 ;
        RECT 52.400 239.600 53.200 239.700 ;
        RECT 278.000 240.300 278.800 240.400 ;
        RECT 383.600 240.300 384.400 240.400 ;
        RECT 388.400 240.300 389.200 240.400 ;
        RECT 423.600 240.300 424.400 240.400 ;
        RECT 278.000 239.700 361.900 240.300 ;
        RECT 278.000 239.600 278.800 239.700 ;
        RECT 182.000 238.300 182.800 238.400 ;
        RECT 193.200 238.300 194.000 238.400 ;
        RECT 182.000 237.700 194.000 238.300 ;
        RECT 182.000 237.600 182.800 237.700 ;
        RECT 193.200 237.600 194.000 237.700 ;
        RECT 226.800 238.300 227.600 238.400 ;
        RECT 346.800 238.300 347.600 238.400 ;
        RECT 226.800 237.700 347.600 238.300 ;
        RECT 226.800 237.600 227.600 237.700 ;
        RECT 346.800 237.600 347.600 237.700 ;
        RECT 351.600 238.300 352.400 238.400 ;
        RECT 359.600 238.300 360.400 238.400 ;
        RECT 351.600 237.700 360.400 238.300 ;
        RECT 361.300 238.300 361.900 239.700 ;
        RECT 383.600 239.700 424.400 240.300 ;
        RECT 383.600 239.600 384.400 239.700 ;
        RECT 388.400 239.600 389.200 239.700 ;
        RECT 423.600 239.600 424.400 239.700 ;
        RECT 436.400 240.300 437.200 240.400 ;
        RECT 454.000 240.300 454.800 240.400 ;
        RECT 436.400 239.700 454.800 240.300 ;
        RECT 436.400 239.600 437.200 239.700 ;
        RECT 454.000 239.600 454.800 239.700 ;
        RECT 474.800 240.300 475.600 240.400 ;
        RECT 490.800 240.300 491.600 240.400 ;
        RECT 474.800 239.700 491.600 240.300 ;
        RECT 474.800 239.600 475.600 239.700 ;
        RECT 490.800 239.600 491.600 239.700 ;
        RECT 514.800 240.300 515.600 240.400 ;
        RECT 522.800 240.300 523.600 240.400 ;
        RECT 514.800 239.700 541.100 240.300 ;
        RECT 514.800 239.600 515.600 239.700 ;
        RECT 522.800 239.600 523.600 239.700 ;
        RECT 540.500 238.400 541.100 239.700 ;
        RECT 463.600 238.300 464.400 238.400 ;
        RECT 361.300 237.700 464.400 238.300 ;
        RECT 351.600 237.600 352.400 237.700 ;
        RECT 359.600 237.600 360.400 237.700 ;
        RECT 463.600 237.600 464.400 237.700 ;
        RECT 495.600 238.300 496.400 238.400 ;
        RECT 506.800 238.300 507.600 238.400 ;
        RECT 495.600 237.700 507.600 238.300 ;
        RECT 495.600 237.600 496.400 237.700 ;
        RECT 506.800 237.600 507.600 237.700 ;
        RECT 540.400 238.300 541.200 238.400 ;
        RECT 554.800 238.300 555.600 238.400 ;
        RECT 540.400 237.700 555.600 238.300 ;
        RECT 540.400 237.600 541.200 237.700 ;
        RECT 554.800 237.600 555.600 237.700 ;
        RECT 566.000 238.300 566.800 238.400 ;
        RECT 574.000 238.300 574.800 238.400 ;
        RECT 566.000 237.700 574.800 238.300 ;
        RECT 566.000 237.600 566.800 237.700 ;
        RECT 574.000 237.600 574.800 237.700 ;
        RECT 586.800 238.300 587.600 238.400 ;
        RECT 588.400 238.300 589.200 238.400 ;
        RECT 586.800 237.700 589.200 238.300 ;
        RECT 586.800 237.600 587.600 237.700 ;
        RECT 588.400 237.600 589.200 237.700 ;
        RECT 18.800 236.300 19.600 236.400 ;
        RECT 30.000 236.300 30.800 236.400 ;
        RECT 33.200 236.300 34.000 236.400 ;
        RECT 18.800 235.700 34.000 236.300 ;
        RECT 18.800 235.600 19.600 235.700 ;
        RECT 30.000 235.600 30.800 235.700 ;
        RECT 33.200 235.600 34.000 235.700 ;
        RECT 302.000 236.300 302.800 236.400 ;
        RECT 353.200 236.300 354.000 236.400 ;
        RECT 302.000 235.700 354.000 236.300 ;
        RECT 302.000 235.600 302.800 235.700 ;
        RECT 353.200 235.600 354.000 235.700 ;
        RECT 404.400 236.300 405.200 236.400 ;
        RECT 407.600 236.300 408.400 236.400 ;
        RECT 404.400 235.700 408.400 236.300 ;
        RECT 404.400 235.600 405.200 235.700 ;
        RECT 407.600 235.600 408.400 235.700 ;
        RECT 409.200 236.300 410.000 236.400 ;
        RECT 505.200 236.300 506.000 236.400 ;
        RECT 409.200 235.700 506.000 236.300 ;
        RECT 409.200 235.600 410.000 235.700 ;
        RECT 505.200 235.600 506.000 235.700 ;
        RECT 506.800 236.300 507.600 236.400 ;
        RECT 511.600 236.300 512.400 236.400 ;
        RECT 506.800 235.700 512.400 236.300 ;
        RECT 506.800 235.600 507.600 235.700 ;
        RECT 511.600 235.600 512.400 235.700 ;
        RECT 526.000 236.300 526.800 236.400 ;
        RECT 530.800 236.300 531.600 236.400 ;
        RECT 526.000 235.700 531.600 236.300 ;
        RECT 526.000 235.600 526.800 235.700 ;
        RECT 530.800 235.600 531.600 235.700 ;
        RECT 532.400 236.300 533.200 236.400 ;
        RECT 566.000 236.300 566.800 236.400 ;
        RECT 532.400 235.700 566.800 236.300 ;
        RECT 532.400 235.600 533.200 235.700 ;
        RECT 566.000 235.600 566.800 235.700 ;
        RECT 12.400 234.300 13.200 234.400 ;
        RECT 15.600 234.300 16.400 234.400 ;
        RECT 12.400 233.700 16.400 234.300 ;
        RECT 12.400 233.600 13.200 233.700 ;
        RECT 15.600 233.600 16.400 233.700 ;
        RECT 82.800 234.300 83.600 234.400 ;
        RECT 124.400 234.300 125.200 234.400 ;
        RECT 82.800 233.700 125.200 234.300 ;
        RECT 82.800 233.600 83.600 233.700 ;
        RECT 124.400 233.600 125.200 233.700 ;
        RECT 321.200 234.300 322.000 234.400 ;
        RECT 335.600 234.300 336.400 234.400 ;
        RECT 342.000 234.300 342.800 234.400 ;
        RECT 348.400 234.300 349.200 234.400 ;
        RECT 351.600 234.300 352.400 234.400 ;
        RECT 321.200 233.700 352.400 234.300 ;
        RECT 321.200 233.600 322.000 233.700 ;
        RECT 335.600 233.600 336.400 233.700 ;
        RECT 342.000 233.600 342.800 233.700 ;
        RECT 348.400 233.600 349.200 233.700 ;
        RECT 351.600 233.600 352.400 233.700 ;
        RECT 399.600 234.300 400.400 234.400 ;
        RECT 404.400 234.300 405.200 234.400 ;
        RECT 476.400 234.300 477.200 234.400 ;
        RECT 399.600 233.700 477.200 234.300 ;
        RECT 399.600 233.600 400.400 233.700 ;
        RECT 404.400 233.600 405.200 233.700 ;
        RECT 476.400 233.600 477.200 233.700 ;
        RECT 487.600 234.300 488.400 234.400 ;
        RECT 492.400 234.300 493.200 234.400 ;
        RECT 487.600 233.700 493.200 234.300 ;
        RECT 487.600 233.600 488.400 233.700 ;
        RECT 492.400 233.600 493.200 233.700 ;
        RECT 508.400 234.300 509.200 234.400 ;
        RECT 519.600 234.300 520.400 234.400 ;
        RECT 530.800 234.300 531.600 234.400 ;
        RECT 543.600 234.300 544.400 234.400 ;
        RECT 508.400 233.700 544.400 234.300 ;
        RECT 508.400 233.600 509.200 233.700 ;
        RECT 519.600 233.600 520.400 233.700 ;
        RECT 530.800 233.600 531.600 233.700 ;
        RECT 543.600 233.600 544.400 233.700 ;
        RECT 596.400 234.300 597.200 234.400 ;
        RECT 604.400 234.300 605.200 234.400 ;
        RECT 596.400 233.700 605.200 234.300 ;
        RECT 596.400 233.600 597.200 233.700 ;
        RECT 604.400 233.600 605.200 233.700 ;
        RECT 9.200 232.300 10.000 232.400 ;
        RECT 22.000 232.300 22.800 232.400 ;
        RECT 9.200 231.700 22.800 232.300 ;
        RECT 9.200 231.600 10.000 231.700 ;
        RECT 22.000 231.600 22.800 231.700 ;
        RECT 25.200 232.300 26.000 232.400 ;
        RECT 33.200 232.300 34.000 232.400 ;
        RECT 25.200 231.700 34.000 232.300 ;
        RECT 25.200 231.600 26.000 231.700 ;
        RECT 33.200 231.600 34.000 231.700 ;
        RECT 271.600 232.300 272.400 232.400 ;
        RECT 273.200 232.300 274.000 232.400 ;
        RECT 271.600 231.700 274.000 232.300 ;
        RECT 271.600 231.600 272.400 231.700 ;
        RECT 273.200 231.600 274.000 231.700 ;
        RECT 298.800 232.300 299.600 232.400 ;
        RECT 302.000 232.300 302.800 232.400 ;
        RECT 298.800 231.700 302.800 232.300 ;
        RECT 298.800 231.600 299.600 231.700 ;
        RECT 302.000 231.600 302.800 231.700 ;
        RECT 303.600 232.300 304.400 232.400 ;
        RECT 313.200 232.300 314.000 232.400 ;
        RECT 303.600 231.700 314.000 232.300 ;
        RECT 303.600 231.600 304.400 231.700 ;
        RECT 313.200 231.600 314.000 231.700 ;
        RECT 314.800 232.300 315.600 232.400 ;
        RECT 340.400 232.300 341.200 232.400 ;
        RECT 314.800 231.700 341.200 232.300 ;
        RECT 314.800 231.600 315.600 231.700 ;
        RECT 340.400 231.600 341.200 231.700 ;
        RECT 346.800 232.300 347.600 232.400 ;
        RECT 351.600 232.300 352.400 232.400 ;
        RECT 346.800 231.700 352.400 232.300 ;
        RECT 346.800 231.600 347.600 231.700 ;
        RECT 351.600 231.600 352.400 231.700 ;
        RECT 354.800 232.300 355.600 232.400 ;
        RECT 407.600 232.300 408.400 232.400 ;
        RECT 354.800 231.700 408.400 232.300 ;
        RECT 354.800 231.600 355.600 231.700 ;
        RECT 407.600 231.600 408.400 231.700 ;
        RECT 428.400 232.300 429.200 232.400 ;
        RECT 450.800 232.300 451.600 232.400 ;
        RECT 470.000 232.300 470.800 232.400 ;
        RECT 471.600 232.300 472.400 232.400 ;
        RECT 428.400 231.700 472.400 232.300 ;
        RECT 428.400 231.600 429.200 231.700 ;
        RECT 450.800 231.600 451.600 231.700 ;
        RECT 470.000 231.600 470.800 231.700 ;
        RECT 471.600 231.600 472.400 231.700 ;
        RECT 474.800 232.300 475.600 232.400 ;
        RECT 478.000 232.300 478.800 232.400 ;
        RECT 474.800 231.700 478.800 232.300 ;
        RECT 474.800 231.600 475.600 231.700 ;
        RECT 478.000 231.600 478.800 231.700 ;
        RECT 481.200 232.300 482.000 232.400 ;
        RECT 484.400 232.300 485.200 232.400 ;
        RECT 487.600 232.300 488.400 232.400 ;
        RECT 481.200 231.700 488.400 232.300 ;
        RECT 481.200 231.600 482.000 231.700 ;
        RECT 484.400 231.600 485.200 231.700 ;
        RECT 487.600 231.600 488.400 231.700 ;
        RECT 495.600 232.300 496.400 232.400 ;
        RECT 524.400 232.300 525.200 232.400 ;
        RECT 495.600 231.700 525.200 232.300 ;
        RECT 495.600 231.600 496.400 231.700 ;
        RECT 524.400 231.600 525.200 231.700 ;
        RECT 530.800 232.300 531.600 232.400 ;
        RECT 532.400 232.300 533.200 232.400 ;
        RECT 530.800 231.700 533.200 232.300 ;
        RECT 530.800 231.600 531.600 231.700 ;
        RECT 532.400 231.600 533.200 231.700 ;
        RECT 545.200 232.300 546.000 232.400 ;
        RECT 548.400 232.300 549.200 232.400 ;
        RECT 545.200 231.700 549.200 232.300 ;
        RECT 545.200 231.600 546.000 231.700 ;
        RECT 548.400 231.600 549.200 231.700 ;
        RECT 550.000 232.300 550.800 232.400 ;
        RECT 562.800 232.300 563.600 232.400 ;
        RECT 550.000 231.700 563.600 232.300 ;
        RECT 550.000 231.600 550.800 231.700 ;
        RECT 562.800 231.600 563.600 231.700 ;
        RECT 586.800 232.300 587.600 232.400 ;
        RECT 604.400 232.300 605.200 232.400 ;
        RECT 586.800 231.700 605.200 232.300 ;
        RECT 586.800 231.600 587.600 231.700 ;
        RECT 604.400 231.600 605.200 231.700 ;
        RECT 15.600 230.300 16.400 230.400 ;
        RECT 18.800 230.300 19.600 230.400 ;
        RECT 15.600 229.700 19.600 230.300 ;
        RECT 15.600 229.600 16.400 229.700 ;
        RECT 18.800 229.600 19.600 229.700 ;
        RECT 23.600 230.300 24.400 230.400 ;
        RECT 26.800 230.300 27.600 230.400 ;
        RECT 76.400 230.300 77.200 230.400 ;
        RECT 82.800 230.300 83.600 230.400 ;
        RECT 130.800 230.300 131.600 230.400 ;
        RECT 134.000 230.300 134.800 230.400 ;
        RECT 265.200 230.300 266.000 230.400 ;
        RECT 23.600 229.700 134.800 230.300 ;
        RECT 23.600 229.600 24.400 229.700 ;
        RECT 26.800 229.600 27.600 229.700 ;
        RECT 76.400 229.600 77.200 229.700 ;
        RECT 82.800 229.600 83.600 229.700 ;
        RECT 130.800 229.600 131.600 229.700 ;
        RECT 134.000 229.600 134.800 229.700 ;
        RECT 244.500 229.700 266.000 230.300 ;
        RECT 244.500 228.400 245.100 229.700 ;
        RECT 265.200 229.600 266.000 229.700 ;
        RECT 266.800 230.300 267.600 230.400 ;
        RECT 287.600 230.300 288.400 230.400 ;
        RECT 266.800 229.700 288.400 230.300 ;
        RECT 266.800 229.600 267.600 229.700 ;
        RECT 287.600 229.600 288.400 229.700 ;
        RECT 297.200 230.300 298.000 230.400 ;
        RECT 311.600 230.300 312.400 230.400 ;
        RECT 297.200 229.700 312.400 230.300 ;
        RECT 297.200 229.600 298.000 229.700 ;
        RECT 311.600 229.600 312.400 229.700 ;
        RECT 319.600 230.300 320.400 230.400 ;
        RECT 321.200 230.300 322.000 230.400 ;
        RECT 319.600 229.700 322.000 230.300 ;
        RECT 319.600 229.600 320.400 229.700 ;
        RECT 321.200 229.600 322.000 229.700 ;
        RECT 340.400 229.600 341.200 230.400 ;
        RECT 358.000 230.300 358.800 230.400 ;
        RECT 359.600 230.300 360.400 230.400 ;
        RECT 358.000 229.700 360.400 230.300 ;
        RECT 358.000 229.600 358.800 229.700 ;
        RECT 359.600 229.600 360.400 229.700 ;
        RECT 364.400 230.300 365.200 230.400 ;
        RECT 401.200 230.300 402.000 230.400 ;
        RECT 364.400 229.700 402.000 230.300 ;
        RECT 364.400 229.600 365.200 229.700 ;
        RECT 401.200 229.600 402.000 229.700 ;
        RECT 452.400 230.300 453.200 230.400 ;
        RECT 478.000 230.300 478.800 230.400 ;
        RECT 452.400 229.700 478.800 230.300 ;
        RECT 452.400 229.600 453.200 229.700 ;
        RECT 478.000 229.600 478.800 229.700 ;
        RECT 494.000 230.300 494.800 230.400 ;
        RECT 497.200 230.300 498.000 230.400 ;
        RECT 494.000 229.700 498.000 230.300 ;
        RECT 494.000 229.600 494.800 229.700 ;
        RECT 497.200 229.600 498.000 229.700 ;
        RECT 500.400 230.300 501.200 230.400 ;
        RECT 506.800 230.300 507.600 230.400 ;
        RECT 530.800 230.300 531.600 230.400 ;
        RECT 500.400 229.700 531.600 230.300 ;
        RECT 500.400 229.600 501.200 229.700 ;
        RECT 506.800 229.600 507.600 229.700 ;
        RECT 530.800 229.600 531.600 229.700 ;
        RECT 538.800 230.300 539.600 230.400 ;
        RECT 542.000 230.300 542.800 230.400 ;
        RECT 538.800 229.700 542.800 230.300 ;
        RECT 538.800 229.600 539.600 229.700 ;
        RECT 542.000 229.600 542.800 229.700 ;
        RECT 558.000 230.300 558.800 230.400 ;
        RECT 562.800 230.300 563.600 230.400 ;
        RECT 558.000 229.700 563.600 230.300 ;
        RECT 558.000 229.600 558.800 229.700 ;
        RECT 562.800 229.600 563.600 229.700 ;
        RECT 602.800 230.300 603.600 230.400 ;
        RECT 604.400 230.300 605.200 230.400 ;
        RECT 602.800 229.700 605.200 230.300 ;
        RECT 602.800 229.600 603.600 229.700 ;
        RECT 604.400 229.600 605.200 229.700 ;
        RECT 2.800 228.300 3.600 228.400 ;
        RECT 7.600 228.300 8.400 228.400 ;
        RECT 2.800 227.700 8.400 228.300 ;
        RECT 2.800 227.600 3.600 227.700 ;
        RECT 7.600 227.600 8.400 227.700 ;
        RECT 18.800 228.300 19.600 228.400 ;
        RECT 33.200 228.300 34.000 228.400 ;
        RECT 18.800 227.700 34.000 228.300 ;
        RECT 18.800 227.600 19.600 227.700 ;
        RECT 33.200 227.600 34.000 227.700 ;
        RECT 42.800 228.300 43.600 228.400 ;
        RECT 57.200 228.300 58.000 228.400 ;
        RECT 42.800 227.700 58.000 228.300 ;
        RECT 42.800 227.600 43.600 227.700 ;
        RECT 57.200 227.600 58.000 227.700 ;
        RECT 84.400 228.300 85.200 228.400 ;
        RECT 102.000 228.300 102.800 228.400 ;
        RECT 84.400 227.700 102.800 228.300 ;
        RECT 84.400 227.600 85.200 227.700 ;
        RECT 102.000 227.600 102.800 227.700 ;
        RECT 185.200 228.300 186.000 228.400 ;
        RECT 185.200 227.700 227.500 228.300 ;
        RECT 185.200 227.600 186.000 227.700 ;
        RECT 6.000 226.300 6.800 226.400 ;
        RECT 20.400 226.300 21.200 226.400 ;
        RECT 6.000 225.700 21.200 226.300 ;
        RECT 6.000 225.600 6.800 225.700 ;
        RECT 20.400 225.600 21.200 225.700 ;
        RECT 22.000 226.300 22.800 226.400 ;
        RECT 41.200 226.300 42.000 226.400 ;
        RECT 22.000 225.700 42.000 226.300 ;
        RECT 22.000 225.600 22.800 225.700 ;
        RECT 41.200 225.600 42.000 225.700 ;
        RECT 68.400 226.300 69.200 226.400 ;
        RECT 225.200 226.300 226.000 226.400 ;
        RECT 68.400 225.700 226.000 226.300 ;
        RECT 226.900 226.300 227.500 227.700 ;
        RECT 244.400 227.600 245.200 228.400 ;
        RECT 263.600 228.300 264.400 228.400 ;
        RECT 274.800 228.300 275.600 228.400 ;
        RECT 263.600 227.700 275.600 228.300 ;
        RECT 263.600 227.600 264.400 227.700 ;
        RECT 274.800 227.600 275.600 227.700 ;
        RECT 294.000 228.300 294.800 228.400 ;
        RECT 303.600 228.300 304.400 228.400 ;
        RECT 294.000 227.700 304.400 228.300 ;
        RECT 294.000 227.600 294.800 227.700 ;
        RECT 303.600 227.600 304.400 227.700 ;
        RECT 305.200 228.300 306.000 228.400 ;
        RECT 348.400 228.300 349.200 228.400 ;
        RECT 305.200 227.700 349.200 228.300 ;
        RECT 305.200 227.600 306.000 227.700 ;
        RECT 348.400 227.600 349.200 227.700 ;
        RECT 356.400 228.300 357.200 228.400 ;
        RECT 370.800 228.300 371.600 228.400 ;
        RECT 356.400 227.700 371.600 228.300 ;
        RECT 356.400 227.600 357.200 227.700 ;
        RECT 370.800 227.600 371.600 227.700 ;
        RECT 372.400 228.300 373.200 228.400 ;
        RECT 380.400 228.300 381.200 228.400 ;
        RECT 372.400 227.700 381.200 228.300 ;
        RECT 372.400 227.600 373.200 227.700 ;
        RECT 380.400 227.600 381.200 227.700 ;
        RECT 382.000 228.300 382.800 228.400 ;
        RECT 415.600 228.300 416.400 228.400 ;
        RECT 428.400 228.300 429.200 228.400 ;
        RECT 430.000 228.300 430.800 228.400 ;
        RECT 382.000 227.700 430.800 228.300 ;
        RECT 382.000 227.600 382.800 227.700 ;
        RECT 415.600 227.600 416.400 227.700 ;
        RECT 428.400 227.600 429.200 227.700 ;
        RECT 430.000 227.600 430.800 227.700 ;
        RECT 447.600 228.300 448.400 228.400 ;
        RECT 455.600 228.300 456.400 228.400 ;
        RECT 447.600 227.700 456.400 228.300 ;
        RECT 447.600 227.600 448.400 227.700 ;
        RECT 455.600 227.600 456.400 227.700 ;
        RECT 468.400 228.300 469.200 228.400 ;
        RECT 471.600 228.300 472.400 228.400 ;
        RECT 468.400 227.700 472.400 228.300 ;
        RECT 468.400 227.600 469.200 227.700 ;
        RECT 471.600 227.600 472.400 227.700 ;
        RECT 482.800 228.300 483.600 228.400 ;
        RECT 508.400 228.300 509.200 228.400 ;
        RECT 482.800 227.700 509.200 228.300 ;
        RECT 482.800 227.600 483.600 227.700 ;
        RECT 508.400 227.600 509.200 227.700 ;
        RECT 513.200 228.300 514.000 228.400 ;
        RECT 519.600 228.300 520.400 228.400 ;
        RECT 513.200 227.700 520.400 228.300 ;
        RECT 513.200 227.600 514.000 227.700 ;
        RECT 519.600 227.600 520.400 227.700 ;
        RECT 534.000 228.300 534.800 228.400 ;
        RECT 559.600 228.300 560.400 228.400 ;
        RECT 534.000 227.700 560.400 228.300 ;
        RECT 534.000 227.600 534.800 227.700 ;
        RECT 559.600 227.600 560.400 227.700 ;
        RECT 572.400 228.300 573.200 228.400 ;
        RECT 602.800 228.300 603.600 228.400 ;
        RECT 572.400 227.700 603.600 228.300 ;
        RECT 572.400 227.600 573.200 227.700 ;
        RECT 602.800 227.600 603.600 227.700 ;
        RECT 282.800 226.300 283.600 226.400 ;
        RECT 334.000 226.300 334.800 226.400 ;
        RECT 354.800 226.300 355.600 226.400 ;
        RECT 226.900 225.700 355.600 226.300 ;
        RECT 68.400 225.600 69.200 225.700 ;
        RECT 225.200 225.600 226.000 225.700 ;
        RECT 282.800 225.600 283.600 225.700 ;
        RECT 334.000 225.600 334.800 225.700 ;
        RECT 354.800 225.600 355.600 225.700 ;
        RECT 366.000 226.300 366.800 226.400 ;
        RECT 410.800 226.300 411.600 226.400 ;
        RECT 366.000 225.700 411.600 226.300 ;
        RECT 366.000 225.600 366.800 225.700 ;
        RECT 410.800 225.600 411.600 225.700 ;
        RECT 444.400 226.300 445.200 226.400 ;
        RECT 466.800 226.300 467.600 226.400 ;
        RECT 444.400 225.700 467.600 226.300 ;
        RECT 444.400 225.600 445.200 225.700 ;
        RECT 466.800 225.600 467.600 225.700 ;
        RECT 519.600 226.300 520.400 226.400 ;
        RECT 526.000 226.300 526.800 226.400 ;
        RECT 551.600 226.300 552.400 226.400 ;
        RECT 519.600 225.700 552.400 226.300 ;
        RECT 519.600 225.600 520.400 225.700 ;
        RECT 526.000 225.600 526.800 225.700 ;
        RECT 551.600 225.600 552.400 225.700 ;
        RECT 585.200 226.300 586.000 226.400 ;
        RECT 604.400 226.300 605.200 226.400 ;
        RECT 585.200 225.700 605.200 226.300 ;
        RECT 585.200 225.600 586.000 225.700 ;
        RECT 604.400 225.600 605.200 225.700 ;
        RECT 87.600 224.300 88.400 224.400 ;
        RECT 132.400 224.300 133.200 224.400 ;
        RECT 87.600 223.700 133.200 224.300 ;
        RECT 87.600 223.600 88.400 223.700 ;
        RECT 132.400 223.600 133.200 223.700 ;
        RECT 217.200 224.300 218.000 224.400 ;
        RECT 220.400 224.300 221.200 224.400 ;
        RECT 217.200 223.700 221.200 224.300 ;
        RECT 217.200 223.600 218.000 223.700 ;
        RECT 220.400 223.600 221.200 223.700 ;
        RECT 244.400 224.300 245.200 224.400 ;
        RECT 350.000 224.300 350.800 224.400 ;
        RECT 434.800 224.300 435.600 224.400 ;
        RECT 446.000 224.300 446.800 224.400 ;
        RECT 458.800 224.300 459.600 224.400 ;
        RECT 244.400 223.700 459.600 224.300 ;
        RECT 244.400 223.600 245.200 223.700 ;
        RECT 350.000 223.600 350.800 223.700 ;
        RECT 434.800 223.600 435.600 223.700 ;
        RECT 446.000 223.600 446.800 223.700 ;
        RECT 458.800 223.600 459.600 223.700 ;
        RECT 465.200 224.300 466.000 224.400 ;
        RECT 468.400 224.300 469.200 224.400 ;
        RECT 465.200 223.700 469.200 224.300 ;
        RECT 465.200 223.600 466.000 223.700 ;
        RECT 468.400 223.600 469.200 223.700 ;
        RECT 530.800 224.300 531.600 224.400 ;
        RECT 548.400 224.300 549.200 224.400 ;
        RECT 530.800 223.700 549.200 224.300 ;
        RECT 530.800 223.600 531.600 223.700 ;
        RECT 548.400 223.600 549.200 223.700 ;
        RECT 55.600 222.300 56.400 222.400 ;
        RECT 84.400 222.300 85.200 222.400 ;
        RECT 55.600 221.700 85.200 222.300 ;
        RECT 55.600 221.600 56.400 221.700 ;
        RECT 84.400 221.600 85.200 221.700 ;
        RECT 201.200 222.300 202.000 222.400 ;
        RECT 209.200 222.300 210.000 222.400 ;
        RECT 201.200 221.700 210.000 222.300 ;
        RECT 201.200 221.600 202.000 221.700 ;
        RECT 209.200 221.600 210.000 221.700 ;
        RECT 249.200 222.300 250.000 222.400 ;
        RECT 295.600 222.300 296.400 222.400 ;
        RECT 249.200 221.700 296.400 222.300 ;
        RECT 249.200 221.600 250.000 221.700 ;
        RECT 295.600 221.600 296.400 221.700 ;
        RECT 311.600 221.600 312.400 222.400 ;
        RECT 337.200 222.300 338.000 222.400 ;
        RECT 382.000 222.300 382.800 222.400 ;
        RECT 337.200 221.700 382.800 222.300 ;
        RECT 337.200 221.600 338.000 221.700 ;
        RECT 382.000 221.600 382.800 221.700 ;
        RECT 401.200 222.300 402.000 222.400 ;
        RECT 500.400 222.300 501.200 222.400 ;
        RECT 518.000 222.300 518.800 222.400 ;
        RECT 522.800 222.300 523.600 222.400 ;
        RECT 529.200 222.300 530.000 222.400 ;
        RECT 401.200 221.700 530.000 222.300 ;
        RECT 401.200 221.600 402.000 221.700 ;
        RECT 500.400 221.600 501.200 221.700 ;
        RECT 518.000 221.600 518.800 221.700 ;
        RECT 522.800 221.600 523.600 221.700 ;
        RECT 529.200 221.600 530.000 221.700 ;
        RECT 546.800 222.300 547.600 222.400 ;
        RECT 569.200 222.300 570.000 222.400 ;
        RECT 546.800 221.700 570.000 222.300 ;
        RECT 546.800 221.600 547.600 221.700 ;
        RECT 569.200 221.600 570.000 221.700 ;
        RECT 60.400 220.300 61.200 220.400 ;
        RECT 66.800 220.300 67.600 220.400 ;
        RECT 60.400 219.700 67.600 220.300 ;
        RECT 60.400 219.600 61.200 219.700 ;
        RECT 66.800 219.600 67.600 219.700 ;
        RECT 346.800 220.300 347.600 220.400 ;
        RECT 351.600 220.300 352.400 220.400 ;
        RECT 346.800 219.700 352.400 220.300 ;
        RECT 346.800 219.600 347.600 219.700 ;
        RECT 351.600 219.600 352.400 219.700 ;
        RECT 367.600 220.300 368.400 220.400 ;
        RECT 383.600 220.300 384.400 220.400 ;
        RECT 367.600 219.700 384.400 220.300 ;
        RECT 367.600 219.600 368.400 219.700 ;
        RECT 383.600 219.600 384.400 219.700 ;
        RECT 441.200 220.300 442.000 220.400 ;
        RECT 460.400 220.300 461.200 220.400 ;
        RECT 441.200 219.700 461.200 220.300 ;
        RECT 441.200 219.600 442.000 219.700 ;
        RECT 460.400 219.600 461.200 219.700 ;
        RECT 463.600 220.300 464.400 220.400 ;
        RECT 474.800 220.300 475.600 220.400 ;
        RECT 463.600 219.700 475.600 220.300 ;
        RECT 463.600 219.600 464.400 219.700 ;
        RECT 474.800 219.600 475.600 219.700 ;
        RECT 497.200 220.300 498.000 220.400 ;
        RECT 505.200 220.300 506.000 220.400 ;
        RECT 538.800 220.300 539.600 220.400 ;
        RECT 553.200 220.300 554.000 220.400 ;
        RECT 497.200 219.700 554.000 220.300 ;
        RECT 497.200 219.600 498.000 219.700 ;
        RECT 505.200 219.600 506.000 219.700 ;
        RECT 538.800 219.600 539.600 219.700 ;
        RECT 553.200 219.600 554.000 219.700 ;
        RECT 556.400 220.300 557.200 220.400 ;
        RECT 591.600 220.300 592.400 220.400 ;
        RECT 556.400 219.700 592.400 220.300 ;
        RECT 556.400 219.600 557.200 219.700 ;
        RECT 591.600 219.600 592.400 219.700 ;
        RECT 92.400 218.300 93.200 218.400 ;
        RECT 95.600 218.300 96.400 218.400 ;
        RECT 106.800 218.300 107.600 218.400 ;
        RECT 150.000 218.300 150.800 218.400 ;
        RECT 166.000 218.300 166.800 218.400 ;
        RECT 92.400 217.700 166.800 218.300 ;
        RECT 92.400 217.600 93.200 217.700 ;
        RECT 95.600 217.600 96.400 217.700 ;
        RECT 106.800 217.600 107.600 217.700 ;
        RECT 150.000 217.600 150.800 217.700 ;
        RECT 166.000 217.600 166.800 217.700 ;
        RECT 172.400 218.300 173.200 218.400 ;
        RECT 198.000 218.300 198.800 218.400 ;
        RECT 172.400 217.700 198.800 218.300 ;
        RECT 172.400 217.600 173.200 217.700 ;
        RECT 198.000 217.600 198.800 217.700 ;
        RECT 228.400 218.300 229.200 218.400 ;
        RECT 247.600 218.300 248.400 218.400 ;
        RECT 228.400 217.700 248.400 218.300 ;
        RECT 228.400 217.600 229.200 217.700 ;
        RECT 247.600 217.600 248.400 217.700 ;
        RECT 300.400 218.300 301.200 218.400 ;
        RECT 482.800 218.300 483.600 218.400 ;
        RECT 300.400 217.700 483.600 218.300 ;
        RECT 300.400 217.600 301.200 217.700 ;
        RECT 482.800 217.600 483.600 217.700 ;
        RECT 532.400 218.300 533.200 218.400 ;
        RECT 558.000 218.300 558.800 218.400 ;
        RECT 532.400 217.700 558.800 218.300 ;
        RECT 532.400 217.600 533.200 217.700 ;
        RECT 558.000 217.600 558.800 217.700 ;
        RECT 15.600 216.300 16.400 216.400 ;
        RECT 31.600 216.300 32.400 216.400 ;
        RECT 15.600 215.700 32.400 216.300 ;
        RECT 15.600 215.600 16.400 215.700 ;
        RECT 31.600 215.600 32.400 215.700 ;
        RECT 74.800 216.300 75.600 216.400 ;
        RECT 100.400 216.300 101.200 216.400 ;
        RECT 74.800 215.700 101.200 216.300 ;
        RECT 74.800 215.600 75.600 215.700 ;
        RECT 100.400 215.600 101.200 215.700 ;
        RECT 118.000 216.300 118.800 216.400 ;
        RECT 122.800 216.300 123.600 216.400 ;
        RECT 118.000 215.700 123.600 216.300 ;
        RECT 166.100 216.300 166.700 217.600 ;
        RECT 194.800 216.300 195.600 216.400 ;
        RECT 204.400 216.300 205.200 216.400 ;
        RECT 166.100 215.700 205.200 216.300 ;
        RECT 118.000 215.600 118.800 215.700 ;
        RECT 122.800 215.600 123.600 215.700 ;
        RECT 194.800 215.600 195.600 215.700 ;
        RECT 204.400 215.600 205.200 215.700 ;
        RECT 260.400 216.300 261.200 216.400 ;
        RECT 266.800 216.300 267.600 216.400 ;
        RECT 260.400 215.700 267.600 216.300 ;
        RECT 260.400 215.600 261.200 215.700 ;
        RECT 266.800 215.600 267.600 215.700 ;
        RECT 274.800 216.300 275.600 216.400 ;
        RECT 318.000 216.300 318.800 216.400 ;
        RECT 274.800 215.700 318.800 216.300 ;
        RECT 274.800 215.600 275.600 215.700 ;
        RECT 318.000 215.600 318.800 215.700 ;
        RECT 340.400 216.300 341.200 216.400 ;
        RECT 356.400 216.300 357.200 216.400 ;
        RECT 340.400 215.700 357.200 216.300 ;
        RECT 340.400 215.600 341.200 215.700 ;
        RECT 356.400 215.600 357.200 215.700 ;
        RECT 370.800 216.300 371.600 216.400 ;
        RECT 386.800 216.300 387.600 216.400 ;
        RECT 370.800 215.700 387.600 216.300 ;
        RECT 370.800 215.600 371.600 215.700 ;
        RECT 386.800 215.600 387.600 215.700 ;
        RECT 455.600 216.300 456.400 216.400 ;
        RECT 481.200 216.300 482.000 216.400 ;
        RECT 455.600 215.700 482.000 216.300 ;
        RECT 455.600 215.600 456.400 215.700 ;
        RECT 481.200 215.600 482.000 215.700 ;
        RECT 511.600 216.300 512.400 216.400 ;
        RECT 567.600 216.300 568.400 216.400 ;
        RECT 511.600 215.700 568.400 216.300 ;
        RECT 511.600 215.600 512.400 215.700 ;
        RECT 567.600 215.600 568.400 215.700 ;
        RECT 23.600 214.300 24.400 214.400 ;
        RECT 33.200 214.300 34.000 214.400 ;
        RECT 39.600 214.300 40.400 214.400 ;
        RECT 46.000 214.300 46.800 214.400 ;
        RECT 23.600 213.700 46.800 214.300 ;
        RECT 23.600 213.600 24.400 213.700 ;
        RECT 33.200 213.600 34.000 213.700 ;
        RECT 39.600 213.600 40.400 213.700 ;
        RECT 46.000 213.600 46.800 213.700 ;
        RECT 92.400 214.300 93.200 214.400 ;
        RECT 102.000 214.300 102.800 214.400 ;
        RECT 92.400 213.700 102.800 214.300 ;
        RECT 92.400 213.600 93.200 213.700 ;
        RECT 102.000 213.600 102.800 213.700 ;
        RECT 110.000 214.300 110.800 214.400 ;
        RECT 124.400 214.300 125.200 214.400 ;
        RECT 143.600 214.300 144.400 214.400 ;
        RECT 110.000 213.700 144.400 214.300 ;
        RECT 110.000 213.600 110.800 213.700 ;
        RECT 124.400 213.600 125.200 213.700 ;
        RECT 143.600 213.600 144.400 213.700 ;
        RECT 164.400 214.300 165.200 214.400 ;
        RECT 175.600 214.300 176.400 214.400 ;
        RECT 164.400 213.700 176.400 214.300 ;
        RECT 164.400 213.600 165.200 213.700 ;
        RECT 175.600 213.600 176.400 213.700 ;
        RECT 222.000 214.300 222.800 214.400 ;
        RECT 225.200 214.300 226.000 214.400 ;
        RECT 222.000 213.700 226.000 214.300 ;
        RECT 222.000 213.600 222.800 213.700 ;
        RECT 225.200 213.600 226.000 213.700 ;
        RECT 263.600 214.300 264.400 214.400 ;
        RECT 279.600 214.300 280.400 214.400 ;
        RECT 263.600 213.700 280.400 214.300 ;
        RECT 263.600 213.600 264.400 213.700 ;
        RECT 279.600 213.600 280.400 213.700 ;
        RECT 297.200 214.300 298.000 214.400 ;
        RECT 302.000 214.300 302.800 214.400 ;
        RECT 337.200 214.300 338.000 214.400 ;
        RECT 297.200 213.700 338.000 214.300 ;
        RECT 297.200 213.600 298.000 213.700 ;
        RECT 302.000 213.600 302.800 213.700 ;
        RECT 337.200 213.600 338.000 213.700 ;
        RECT 350.000 214.300 350.800 214.400 ;
        RECT 385.200 214.300 386.000 214.400 ;
        RECT 350.000 213.700 386.000 214.300 ;
        RECT 350.000 213.600 350.800 213.700 ;
        RECT 385.200 213.600 386.000 213.700 ;
        RECT 410.800 214.300 411.600 214.400 ;
        RECT 420.400 214.300 421.200 214.400 ;
        RECT 410.800 213.700 421.200 214.300 ;
        RECT 410.800 213.600 411.600 213.700 ;
        RECT 420.400 213.600 421.200 213.700 ;
        RECT 425.200 214.300 426.000 214.400 ;
        RECT 446.000 214.300 446.800 214.400 ;
        RECT 425.200 213.700 446.800 214.300 ;
        RECT 425.200 213.600 426.000 213.700 ;
        RECT 446.000 213.600 446.800 213.700 ;
        RECT 516.400 214.300 517.200 214.400 ;
        RECT 535.600 214.300 536.400 214.400 ;
        RECT 546.800 214.300 547.600 214.400 ;
        RECT 516.400 213.700 547.600 214.300 ;
        RECT 516.400 213.600 517.200 213.700 ;
        RECT 535.600 213.600 536.400 213.700 ;
        RECT 546.800 213.600 547.600 213.700 ;
        RECT 554.800 214.300 555.600 214.400 ;
        RECT 578.800 214.300 579.600 214.400 ;
        RECT 554.800 213.700 579.600 214.300 ;
        RECT 554.800 213.600 555.600 213.700 ;
        RECT 578.800 213.600 579.600 213.700 ;
        RECT 4.400 212.300 5.200 212.400 ;
        RECT 6.000 212.300 6.800 212.400 ;
        RECT 9.200 212.300 10.000 212.400 ;
        RECT 4.400 211.700 10.000 212.300 ;
        RECT 4.400 211.600 5.200 211.700 ;
        RECT 6.000 211.600 6.800 211.700 ;
        RECT 9.200 211.600 10.000 211.700 ;
        RECT 14.000 212.300 14.800 212.400 ;
        RECT 18.800 212.300 19.600 212.400 ;
        RECT 14.000 211.700 19.600 212.300 ;
        RECT 14.000 211.600 14.800 211.700 ;
        RECT 18.800 211.600 19.600 211.700 ;
        RECT 82.800 212.300 83.600 212.400 ;
        RECT 108.400 212.300 109.200 212.400 ;
        RECT 82.800 211.700 109.200 212.300 ;
        RECT 82.800 211.600 83.600 211.700 ;
        RECT 108.400 211.600 109.200 211.700 ;
        RECT 113.200 212.300 114.000 212.400 ;
        RECT 116.400 212.300 117.200 212.400 ;
        RECT 113.200 211.700 117.200 212.300 ;
        RECT 113.200 211.600 114.000 211.700 ;
        RECT 116.400 211.600 117.200 211.700 ;
        RECT 204.400 212.300 205.200 212.400 ;
        RECT 212.400 212.300 213.200 212.400 ;
        RECT 215.600 212.300 216.400 212.400 ;
        RECT 204.400 211.700 216.400 212.300 ;
        RECT 204.400 211.600 205.200 211.700 ;
        RECT 212.400 211.600 213.200 211.700 ;
        RECT 215.600 211.600 216.400 211.700 ;
        RECT 484.400 212.300 485.200 212.400 ;
        RECT 519.600 212.300 520.400 212.400 ;
        RECT 484.400 211.700 520.400 212.300 ;
        RECT 484.400 211.600 485.200 211.700 ;
        RECT 519.600 211.600 520.400 211.700 ;
        RECT 567.600 212.300 568.400 212.400 ;
        RECT 577.200 212.300 578.000 212.400 ;
        RECT 567.600 211.700 578.000 212.300 ;
        RECT 567.600 211.600 568.400 211.700 ;
        RECT 577.200 211.600 578.000 211.700 ;
        RECT 9.200 210.300 10.000 210.400 ;
        RECT 18.800 210.300 19.600 210.400 ;
        RECT 9.200 209.700 19.600 210.300 ;
        RECT 9.200 209.600 10.000 209.700 ;
        RECT 18.800 209.600 19.600 209.700 ;
        RECT 22.000 210.300 22.800 210.400 ;
        RECT 26.800 210.300 27.600 210.400 ;
        RECT 33.200 210.300 34.000 210.400 ;
        RECT 22.000 209.700 34.000 210.300 ;
        RECT 108.500 210.300 109.100 211.600 ;
        RECT 121.200 210.300 122.000 210.400 ;
        RECT 108.500 209.700 122.000 210.300 ;
        RECT 22.000 209.600 22.800 209.700 ;
        RECT 26.800 209.600 27.600 209.700 ;
        RECT 33.200 209.600 34.000 209.700 ;
        RECT 121.200 209.600 122.000 209.700 ;
        RECT 134.000 210.300 134.800 210.400 ;
        RECT 148.400 210.300 149.200 210.400 ;
        RECT 134.000 209.700 149.200 210.300 ;
        RECT 134.000 209.600 134.800 209.700 ;
        RECT 148.400 209.600 149.200 209.700 ;
        RECT 382.000 210.300 382.800 210.400 ;
        RECT 388.400 210.300 389.200 210.400 ;
        RECT 382.000 209.700 389.200 210.300 ;
        RECT 382.000 209.600 382.800 209.700 ;
        RECT 388.400 209.600 389.200 209.700 ;
        RECT 410.800 210.300 411.600 210.400 ;
        RECT 412.400 210.300 413.200 210.400 ;
        RECT 426.800 210.300 427.600 210.400 ;
        RECT 410.800 209.700 427.600 210.300 ;
        RECT 410.800 209.600 411.600 209.700 ;
        RECT 412.400 209.600 413.200 209.700 ;
        RECT 426.800 209.600 427.600 209.700 ;
        RECT 489.200 210.300 490.000 210.400 ;
        RECT 503.600 210.300 504.400 210.400 ;
        RECT 489.200 209.700 504.400 210.300 ;
        RECT 489.200 209.600 490.000 209.700 ;
        RECT 503.600 209.600 504.400 209.700 ;
        RECT 564.400 210.300 565.200 210.400 ;
        RECT 574.000 210.300 574.800 210.400 ;
        RECT 564.400 209.700 574.800 210.300 ;
        RECT 564.400 209.600 565.200 209.700 ;
        RECT 574.000 209.600 574.800 209.700 ;
        RECT 25.200 208.300 26.000 208.400 ;
        RECT 34.800 208.300 35.600 208.400 ;
        RECT 25.200 207.700 35.600 208.300 ;
        RECT 25.200 207.600 26.000 207.700 ;
        RECT 34.800 207.600 35.600 207.700 ;
        RECT 76.400 208.300 77.200 208.400 ;
        RECT 79.600 208.300 80.400 208.400 ;
        RECT 105.200 208.300 106.000 208.400 ;
        RECT 76.400 207.700 106.000 208.300 ;
        RECT 76.400 207.600 77.200 207.700 ;
        RECT 79.600 207.600 80.400 207.700 ;
        RECT 105.200 207.600 106.000 207.700 ;
        RECT 130.800 208.300 131.600 208.400 ;
        RECT 137.200 208.300 138.000 208.400 ;
        RECT 130.800 207.700 138.000 208.300 ;
        RECT 130.800 207.600 131.600 207.700 ;
        RECT 137.200 207.600 138.000 207.700 ;
        RECT 145.200 208.300 146.000 208.400 ;
        RECT 166.000 208.300 166.800 208.400 ;
        RECT 145.200 207.700 166.800 208.300 ;
        RECT 145.200 207.600 146.000 207.700 ;
        RECT 166.000 207.600 166.800 207.700 ;
        RECT 282.800 206.300 283.600 206.400 ;
        RECT 287.600 206.300 288.400 206.400 ;
        RECT 516.400 206.300 517.200 206.400 ;
        RECT 282.800 205.700 517.200 206.300 ;
        RECT 282.800 205.600 283.600 205.700 ;
        RECT 287.600 205.600 288.400 205.700 ;
        RECT 516.400 205.600 517.200 205.700 ;
        RECT 236.400 204.300 237.200 204.400 ;
        RECT 244.400 204.300 245.200 204.400 ;
        RECT 236.400 203.700 245.200 204.300 ;
        RECT 236.400 203.600 237.200 203.700 ;
        RECT 244.400 203.600 245.200 203.700 ;
        RECT 321.200 204.300 322.000 204.400 ;
        RECT 324.400 204.300 325.200 204.400 ;
        RECT 321.200 203.700 325.200 204.300 ;
        RECT 321.200 203.600 322.000 203.700 ;
        RECT 324.400 203.600 325.200 203.700 ;
        RECT 345.200 204.300 346.000 204.400 ;
        RECT 346.800 204.300 347.600 204.400 ;
        RECT 345.200 203.700 347.600 204.300 ;
        RECT 345.200 203.600 346.000 203.700 ;
        RECT 346.800 203.600 347.600 203.700 ;
        RECT 567.600 204.300 568.400 204.400 ;
        RECT 572.400 204.300 573.200 204.400 ;
        RECT 567.600 203.700 573.200 204.300 ;
        RECT 567.600 203.600 568.400 203.700 ;
        RECT 572.400 203.600 573.200 203.700 ;
        RECT 78.000 202.300 78.800 202.400 ;
        RECT 84.400 202.300 85.200 202.400 ;
        RECT 78.000 201.700 85.200 202.300 ;
        RECT 78.000 201.600 78.800 201.700 ;
        RECT 84.400 201.600 85.200 201.700 ;
        RECT 310.000 202.300 310.800 202.400 ;
        RECT 311.600 202.300 312.400 202.400 ;
        RECT 310.000 201.700 312.400 202.300 ;
        RECT 310.000 201.600 310.800 201.700 ;
        RECT 311.600 201.600 312.400 201.700 ;
        RECT 374.000 202.300 374.800 202.400 ;
        RECT 378.800 202.300 379.600 202.400 ;
        RECT 374.000 201.700 379.600 202.300 ;
        RECT 374.000 201.600 374.800 201.700 ;
        RECT 378.800 201.600 379.600 201.700 ;
        RECT 433.200 200.300 434.000 200.400 ;
        RECT 442.800 200.300 443.600 200.400 ;
        RECT 450.800 200.300 451.600 200.400 ;
        RECT 433.200 199.700 451.600 200.300 ;
        RECT 433.200 199.600 434.000 199.700 ;
        RECT 442.800 199.600 443.600 199.700 ;
        RECT 450.800 199.600 451.600 199.700 ;
        RECT 84.400 198.300 85.200 198.400 ;
        RECT 86.000 198.300 86.800 198.400 ;
        RECT 84.400 197.700 86.800 198.300 ;
        RECT 84.400 197.600 85.200 197.700 ;
        RECT 86.000 197.600 86.800 197.700 ;
        RECT 98.800 198.300 99.600 198.400 ;
        RECT 106.800 198.300 107.600 198.400 ;
        RECT 111.600 198.300 112.400 198.400 ;
        RECT 135.600 198.300 136.400 198.400 ;
        RECT 142.000 198.300 142.800 198.400 ;
        RECT 161.200 198.300 162.000 198.400 ;
        RECT 164.400 198.300 165.200 198.400 ;
        RECT 98.800 197.700 165.200 198.300 ;
        RECT 98.800 197.600 99.600 197.700 ;
        RECT 106.800 197.600 107.600 197.700 ;
        RECT 111.600 197.600 112.400 197.700 ;
        RECT 135.600 197.600 136.400 197.700 ;
        RECT 142.000 197.600 142.800 197.700 ;
        RECT 161.200 197.600 162.000 197.700 ;
        RECT 164.400 197.600 165.200 197.700 ;
        RECT 410.800 198.300 411.600 198.400 ;
        RECT 417.200 198.300 418.000 198.400 ;
        RECT 410.800 197.700 418.000 198.300 ;
        RECT 410.800 197.600 411.600 197.700 ;
        RECT 417.200 197.600 418.000 197.700 ;
        RECT 577.200 198.300 578.000 198.400 ;
        RECT 590.000 198.300 590.800 198.400 ;
        RECT 577.200 197.700 590.800 198.300 ;
        RECT 577.200 197.600 578.000 197.700 ;
        RECT 590.000 197.600 590.800 197.700 ;
        RECT 57.200 196.300 58.000 196.400 ;
        RECT 70.000 196.300 70.800 196.400 ;
        RECT 57.200 195.700 70.800 196.300 ;
        RECT 57.200 195.600 58.000 195.700 ;
        RECT 70.000 195.600 70.800 195.700 ;
        RECT 271.600 196.300 272.400 196.400 ;
        RECT 290.800 196.300 291.600 196.400 ;
        RECT 318.000 196.300 318.800 196.400 ;
        RECT 340.400 196.300 341.200 196.400 ;
        RECT 367.600 196.300 368.400 196.400 ;
        RECT 382.000 196.300 382.800 196.400 ;
        RECT 271.600 195.700 382.800 196.300 ;
        RECT 271.600 195.600 272.400 195.700 ;
        RECT 290.800 195.600 291.600 195.700 ;
        RECT 318.000 195.600 318.800 195.700 ;
        RECT 340.400 195.600 341.200 195.700 ;
        RECT 367.600 195.600 368.400 195.700 ;
        RECT 382.000 195.600 382.800 195.700 ;
        RECT 479.600 196.300 480.400 196.400 ;
        RECT 506.800 196.300 507.600 196.400 ;
        RECT 479.600 195.700 507.600 196.300 ;
        RECT 479.600 195.600 480.400 195.700 ;
        RECT 506.800 195.600 507.600 195.700 ;
        RECT 38.000 194.300 38.800 194.400 ;
        RECT 71.600 194.300 72.400 194.400 ;
        RECT 73.200 194.300 74.000 194.400 ;
        RECT 114.800 194.300 115.600 194.400 ;
        RECT 38.000 193.700 115.600 194.300 ;
        RECT 38.000 193.600 38.800 193.700 ;
        RECT 71.600 193.600 72.400 193.700 ;
        RECT 73.200 193.600 74.000 193.700 ;
        RECT 114.800 193.600 115.600 193.700 ;
        RECT 244.400 194.300 245.200 194.400 ;
        RECT 286.000 194.300 286.800 194.400 ;
        RECT 287.600 194.300 288.400 194.400 ;
        RECT 244.400 193.700 288.400 194.300 ;
        RECT 244.400 193.600 245.200 193.700 ;
        RECT 286.000 193.600 286.800 193.700 ;
        RECT 287.600 193.600 288.400 193.700 ;
        RECT 343.600 193.600 344.400 194.400 ;
        RECT 353.200 194.300 354.000 194.400 ;
        RECT 358.000 194.300 358.800 194.400 ;
        RECT 366.000 194.300 366.800 194.400 ;
        RECT 353.200 193.700 366.800 194.300 ;
        RECT 353.200 193.600 354.000 193.700 ;
        RECT 358.000 193.600 358.800 193.700 ;
        RECT 366.000 193.600 366.800 193.700 ;
        RECT 412.400 194.300 413.200 194.400 ;
        RECT 481.200 194.300 482.000 194.400 ;
        RECT 412.400 193.700 482.000 194.300 ;
        RECT 412.400 193.600 413.200 193.700 ;
        RECT 481.200 193.600 482.000 193.700 ;
        RECT 503.600 194.300 504.400 194.400 ;
        RECT 518.000 194.300 518.800 194.400 ;
        RECT 503.600 193.700 518.800 194.300 ;
        RECT 503.600 193.600 504.400 193.700 ;
        RECT 518.000 193.600 518.800 193.700 ;
        RECT 526.000 194.300 526.800 194.400 ;
        RECT 594.800 194.300 595.600 194.400 ;
        RECT 526.000 193.700 595.600 194.300 ;
        RECT 526.000 193.600 526.800 193.700 ;
        RECT 594.800 193.600 595.600 193.700 ;
        RECT 25.200 192.300 26.000 192.400 ;
        RECT 47.600 192.300 48.400 192.400 ;
        RECT 25.200 191.700 48.400 192.300 ;
        RECT 25.200 191.600 26.000 191.700 ;
        RECT 47.600 191.600 48.400 191.700 ;
        RECT 58.800 192.300 59.600 192.400 ;
        RECT 66.800 192.300 67.600 192.400 ;
        RECT 58.800 191.700 67.600 192.300 ;
        RECT 58.800 191.600 59.600 191.700 ;
        RECT 66.800 191.600 67.600 191.700 ;
        RECT 70.000 192.300 70.800 192.400 ;
        RECT 78.000 192.300 78.800 192.400 ;
        RECT 70.000 191.700 78.800 192.300 ;
        RECT 70.000 191.600 70.800 191.700 ;
        RECT 78.000 191.600 78.800 191.700 ;
        RECT 94.000 192.300 94.800 192.400 ;
        RECT 108.400 192.300 109.200 192.400 ;
        RECT 94.000 191.700 109.200 192.300 ;
        RECT 94.000 191.600 94.800 191.700 ;
        RECT 108.400 191.600 109.200 191.700 ;
        RECT 111.600 192.300 112.400 192.400 ;
        RECT 121.200 192.300 122.000 192.400 ;
        RECT 111.600 191.700 122.000 192.300 ;
        RECT 111.600 191.600 112.400 191.700 ;
        RECT 121.200 191.600 122.000 191.700 ;
        RECT 199.600 192.300 200.400 192.400 ;
        RECT 247.600 192.300 248.400 192.400 ;
        RECT 199.600 191.700 248.400 192.300 ;
        RECT 199.600 191.600 200.400 191.700 ;
        RECT 247.600 191.600 248.400 191.700 ;
        RECT 476.400 192.300 477.200 192.400 ;
        RECT 495.600 192.300 496.400 192.400 ;
        RECT 476.400 191.700 496.400 192.300 ;
        RECT 476.400 191.600 477.200 191.700 ;
        RECT 495.600 191.600 496.400 191.700 ;
        RECT 498.800 192.300 499.600 192.400 ;
        RECT 502.000 192.300 502.800 192.400 ;
        RECT 498.800 191.700 502.800 192.300 ;
        RECT 498.800 191.600 499.600 191.700 ;
        RECT 502.000 191.600 502.800 191.700 ;
        RECT 510.000 192.300 510.800 192.400 ;
        RECT 537.200 192.300 538.000 192.400 ;
        RECT 510.000 191.700 538.000 192.300 ;
        RECT 510.000 191.600 510.800 191.700 ;
        RECT 537.200 191.600 538.000 191.700 ;
        RECT 575.600 192.300 576.400 192.400 ;
        RECT 598.000 192.300 598.800 192.400 ;
        RECT 575.600 191.700 598.800 192.300 ;
        RECT 575.600 191.600 576.400 191.700 ;
        RECT 598.000 191.600 598.800 191.700 ;
        RECT 14.000 189.600 14.800 190.400 ;
        RECT 47.600 190.300 48.400 190.400 ;
        RECT 58.800 190.300 59.600 190.400 ;
        RECT 47.600 189.700 59.600 190.300 ;
        RECT 47.600 189.600 48.400 189.700 ;
        RECT 58.800 189.600 59.600 189.700 ;
        RECT 62.000 190.300 62.800 190.400 ;
        RECT 71.600 190.300 72.400 190.400 ;
        RECT 62.000 189.700 72.400 190.300 ;
        RECT 62.000 189.600 62.800 189.700 ;
        RECT 71.600 189.600 72.400 189.700 ;
        RECT 102.000 190.300 102.800 190.400 ;
        RECT 108.400 190.300 109.200 190.400 ;
        RECT 102.000 189.700 109.200 190.300 ;
        RECT 102.000 189.600 102.800 189.700 ;
        RECT 108.400 189.600 109.200 189.700 ;
        RECT 127.600 190.300 128.400 190.400 ;
        RECT 135.600 190.300 136.400 190.400 ;
        RECT 145.200 190.300 146.000 190.400 ;
        RECT 127.600 189.700 146.000 190.300 ;
        RECT 127.600 189.600 128.400 189.700 ;
        RECT 135.600 189.600 136.400 189.700 ;
        RECT 145.200 189.600 146.000 189.700 ;
        RECT 151.600 190.300 152.400 190.400 ;
        RECT 159.600 190.300 160.400 190.400 ;
        RECT 170.800 190.300 171.600 190.400 ;
        RECT 151.600 189.700 171.600 190.300 ;
        RECT 151.600 189.600 152.400 189.700 ;
        RECT 159.600 189.600 160.400 189.700 ;
        RECT 170.800 189.600 171.600 189.700 ;
        RECT 206.000 190.300 206.800 190.400 ;
        RECT 207.600 190.300 208.400 190.400 ;
        RECT 206.000 189.700 208.400 190.300 ;
        RECT 206.000 189.600 206.800 189.700 ;
        RECT 207.600 189.600 208.400 189.700 ;
        RECT 209.200 190.300 210.000 190.400 ;
        RECT 234.800 190.300 235.600 190.400 ;
        RECT 209.200 189.700 235.600 190.300 ;
        RECT 209.200 189.600 210.000 189.700 ;
        RECT 234.800 189.600 235.600 189.700 ;
        RECT 249.200 190.300 250.000 190.400 ;
        RECT 258.800 190.300 259.600 190.400 ;
        RECT 249.200 189.700 259.600 190.300 ;
        RECT 249.200 189.600 250.000 189.700 ;
        RECT 258.800 189.600 259.600 189.700 ;
        RECT 286.000 190.300 286.800 190.400 ;
        RECT 295.600 190.300 296.400 190.400 ;
        RECT 286.000 189.700 296.400 190.300 ;
        RECT 286.000 189.600 286.800 189.700 ;
        RECT 295.600 189.600 296.400 189.700 ;
        RECT 311.600 190.300 312.400 190.400 ;
        RECT 313.200 190.300 314.000 190.400 ;
        RECT 318.000 190.300 318.800 190.400 ;
        RECT 346.800 190.300 347.600 190.400 ;
        RECT 361.200 190.300 362.000 190.400 ;
        RECT 366.000 190.300 366.800 190.400 ;
        RECT 402.800 190.300 403.600 190.400 ;
        RECT 311.600 189.700 403.600 190.300 ;
        RECT 311.600 189.600 312.400 189.700 ;
        RECT 313.200 189.600 314.000 189.700 ;
        RECT 318.000 189.600 318.800 189.700 ;
        RECT 346.800 189.600 347.600 189.700 ;
        RECT 361.200 189.600 362.000 189.700 ;
        RECT 366.000 189.600 366.800 189.700 ;
        RECT 402.800 189.600 403.600 189.700 ;
        RECT 466.800 190.300 467.600 190.400 ;
        RECT 468.400 190.300 469.200 190.400 ;
        RECT 466.800 189.700 469.200 190.300 ;
        RECT 466.800 189.600 467.600 189.700 ;
        RECT 468.400 189.600 469.200 189.700 ;
        RECT 476.400 190.300 477.200 190.400 ;
        RECT 479.600 190.300 480.400 190.400 ;
        RECT 476.400 189.700 480.400 190.300 ;
        RECT 476.400 189.600 477.200 189.700 ;
        RECT 479.600 189.600 480.400 189.700 ;
        RECT 494.000 190.300 494.800 190.400 ;
        RECT 513.200 190.300 514.000 190.400 ;
        RECT 529.200 190.300 530.000 190.400 ;
        RECT 494.000 189.700 530.000 190.300 ;
        RECT 494.000 189.600 494.800 189.700 ;
        RECT 513.200 189.600 514.000 189.700 ;
        RECT 529.200 189.600 530.000 189.700 ;
        RECT 559.600 190.300 560.400 190.400 ;
        RECT 566.000 190.300 566.800 190.400 ;
        RECT 559.600 189.700 566.800 190.300 ;
        RECT 559.600 189.600 560.400 189.700 ;
        RECT 566.000 189.600 566.800 189.700 ;
        RECT 594.800 190.300 595.600 190.400 ;
        RECT 602.800 190.300 603.600 190.400 ;
        RECT 594.800 189.700 603.600 190.300 ;
        RECT 594.800 189.600 595.600 189.700 ;
        RECT 602.800 189.600 603.600 189.700 ;
        RECT 6.000 188.300 6.800 188.400 ;
        RECT 14.000 188.300 14.800 188.400 ;
        RECT 6.000 187.700 14.800 188.300 ;
        RECT 6.000 187.600 6.800 187.700 ;
        RECT 14.000 187.600 14.800 187.700 ;
        RECT 33.200 188.300 34.000 188.400 ;
        RECT 38.000 188.300 38.800 188.400 ;
        RECT 33.200 187.700 38.800 188.300 ;
        RECT 33.200 187.600 34.000 187.700 ;
        RECT 38.000 187.600 38.800 187.700 ;
        RECT 68.400 188.300 69.200 188.400 ;
        RECT 89.200 188.300 90.000 188.400 ;
        RECT 68.400 187.700 90.000 188.300 ;
        RECT 68.400 187.600 69.200 187.700 ;
        RECT 89.200 187.600 90.000 187.700 ;
        RECT 92.400 188.300 93.200 188.400 ;
        RECT 124.400 188.300 125.200 188.400 ;
        RECT 127.600 188.300 128.400 188.400 ;
        RECT 132.400 188.300 133.200 188.400 ;
        RECT 92.400 187.700 133.200 188.300 ;
        RECT 92.400 187.600 93.200 187.700 ;
        RECT 124.400 187.600 125.200 187.700 ;
        RECT 127.600 187.600 128.400 187.700 ;
        RECT 132.400 187.600 133.200 187.700 ;
        RECT 172.400 188.300 173.200 188.400 ;
        RECT 193.200 188.300 194.000 188.400 ;
        RECT 172.400 187.700 194.000 188.300 ;
        RECT 172.400 187.600 173.200 187.700 ;
        RECT 193.200 187.600 194.000 187.700 ;
        RECT 210.800 188.300 211.600 188.400 ;
        RECT 215.600 188.300 216.400 188.400 ;
        RECT 210.800 187.700 216.400 188.300 ;
        RECT 210.800 187.600 211.600 187.700 ;
        RECT 215.600 187.600 216.400 187.700 ;
        RECT 223.600 188.300 224.400 188.400 ;
        RECT 231.600 188.300 232.400 188.400 ;
        RECT 238.000 188.300 238.800 188.400 ;
        RECT 223.600 187.700 238.800 188.300 ;
        RECT 223.600 187.600 224.400 187.700 ;
        RECT 231.600 187.600 232.400 187.700 ;
        RECT 238.000 187.600 238.800 187.700 ;
        RECT 247.600 188.300 248.400 188.400 ;
        RECT 268.400 188.300 269.200 188.400 ;
        RECT 247.600 187.700 269.200 188.300 ;
        RECT 247.600 187.600 248.400 187.700 ;
        RECT 268.400 187.600 269.200 187.700 ;
        RECT 295.600 188.300 296.400 188.400 ;
        RECT 300.400 188.300 301.200 188.400 ;
        RECT 295.600 187.700 301.200 188.300 ;
        RECT 295.600 187.600 296.400 187.700 ;
        RECT 300.400 187.600 301.200 187.700 ;
        RECT 362.800 188.300 363.600 188.400 ;
        RECT 385.200 188.300 386.000 188.400 ;
        RECT 362.800 187.700 386.000 188.300 ;
        RECT 362.800 187.600 363.600 187.700 ;
        RECT 385.200 187.600 386.000 187.700 ;
        RECT 396.400 188.300 397.200 188.400 ;
        RECT 404.400 188.300 405.200 188.400 ;
        RECT 434.800 188.300 435.600 188.400 ;
        RECT 438.000 188.300 438.800 188.400 ;
        RECT 396.400 187.700 438.800 188.300 ;
        RECT 396.400 187.600 397.200 187.700 ;
        RECT 404.400 187.600 405.200 187.700 ;
        RECT 434.800 187.600 435.600 187.700 ;
        RECT 438.000 187.600 438.800 187.700 ;
        RECT 450.800 188.300 451.600 188.400 ;
        RECT 481.200 188.300 482.000 188.400 ;
        RECT 450.800 187.700 482.000 188.300 ;
        RECT 450.800 187.600 451.600 187.700 ;
        RECT 481.200 187.600 482.000 187.700 ;
        RECT 519.600 188.300 520.400 188.400 ;
        RECT 575.600 188.300 576.400 188.400 ;
        RECT 519.600 187.700 576.400 188.300 ;
        RECT 519.600 187.600 520.400 187.700 ;
        RECT 575.600 187.600 576.400 187.700 ;
        RECT 602.800 188.300 603.600 188.400 ;
        RECT 609.200 188.300 610.000 188.400 ;
        RECT 602.800 187.700 610.000 188.300 ;
        RECT 602.800 187.600 603.600 187.700 ;
        RECT 609.200 187.600 610.000 187.700 ;
        RECT 6.000 186.300 6.800 186.400 ;
        RECT 17.200 186.300 18.000 186.400 ;
        RECT 41.200 186.300 42.000 186.400 ;
        RECT 6.000 185.700 42.000 186.300 ;
        RECT 6.000 185.600 6.800 185.700 ;
        RECT 17.200 185.600 18.000 185.700 ;
        RECT 41.200 185.600 42.000 185.700 ;
        RECT 49.200 186.300 50.000 186.400 ;
        RECT 79.600 186.300 80.400 186.400 ;
        RECT 134.000 186.300 134.800 186.400 ;
        RECT 150.000 186.300 150.800 186.400 ;
        RECT 49.200 185.700 150.800 186.300 ;
        RECT 49.200 185.600 50.000 185.700 ;
        RECT 79.600 185.600 80.400 185.700 ;
        RECT 134.000 185.600 134.800 185.700 ;
        RECT 150.000 185.600 150.800 185.700 ;
        RECT 177.200 186.300 178.000 186.400 ;
        RECT 190.000 186.300 190.800 186.400 ;
        RECT 177.200 185.700 190.800 186.300 ;
        RECT 177.200 185.600 178.000 185.700 ;
        RECT 190.000 185.600 190.800 185.700 ;
        RECT 206.000 186.300 206.800 186.400 ;
        RECT 212.400 186.300 213.200 186.400 ;
        RECT 223.700 186.300 224.300 187.600 ;
        RECT 206.000 185.700 224.300 186.300 ;
        RECT 292.400 186.300 293.200 186.400 ;
        RECT 308.400 186.300 309.200 186.400 ;
        RECT 292.400 185.700 309.200 186.300 ;
        RECT 206.000 185.600 206.800 185.700 ;
        RECT 212.400 185.600 213.200 185.700 ;
        RECT 292.400 185.600 293.200 185.700 ;
        RECT 308.400 185.600 309.200 185.700 ;
        RECT 382.000 186.300 382.800 186.400 ;
        RECT 415.600 186.300 416.400 186.400 ;
        RECT 382.000 185.700 416.400 186.300 ;
        RECT 382.000 185.600 382.800 185.700 ;
        RECT 415.600 185.600 416.400 185.700 ;
        RECT 438.000 186.300 438.800 186.400 ;
        RECT 503.600 186.300 504.400 186.400 ;
        RECT 522.800 186.300 523.600 186.400 ;
        RECT 438.000 185.700 523.600 186.300 ;
        RECT 438.000 185.600 438.800 185.700 ;
        RECT 503.600 185.600 504.400 185.700 ;
        RECT 522.800 185.600 523.600 185.700 ;
        RECT 545.200 186.300 546.000 186.400 ;
        RECT 554.800 186.300 555.600 186.400 ;
        RECT 545.200 185.700 555.600 186.300 ;
        RECT 545.200 185.600 546.000 185.700 ;
        RECT 554.800 185.600 555.600 185.700 ;
        RECT 574.000 186.300 574.800 186.400 ;
        RECT 578.800 186.300 579.600 186.400 ;
        RECT 574.000 185.700 579.600 186.300 ;
        RECT 574.000 185.600 574.800 185.700 ;
        RECT 578.800 185.600 579.600 185.700 ;
        RECT 36.400 184.300 37.200 184.400 ;
        RECT 38.000 184.300 38.800 184.400 ;
        RECT 36.400 183.700 38.800 184.300 ;
        RECT 36.400 183.600 37.200 183.700 ;
        RECT 38.000 183.600 38.800 183.700 ;
        RECT 113.200 184.300 114.000 184.400 ;
        RECT 121.200 184.300 122.000 184.400 ;
        RECT 113.200 183.700 122.000 184.300 ;
        RECT 113.200 183.600 114.000 183.700 ;
        RECT 121.200 183.600 122.000 183.700 ;
        RECT 204.400 184.300 205.200 184.400 ;
        RECT 214.000 184.300 214.800 184.400 ;
        RECT 233.200 184.300 234.000 184.400 ;
        RECT 239.600 184.300 240.400 184.400 ;
        RECT 294.000 184.300 294.800 184.400 ;
        RECT 204.400 183.700 294.800 184.300 ;
        RECT 204.400 183.600 205.200 183.700 ;
        RECT 214.000 183.600 214.800 183.700 ;
        RECT 233.200 183.600 234.000 183.700 ;
        RECT 239.600 183.600 240.400 183.700 ;
        RECT 294.000 183.600 294.800 183.700 ;
        RECT 340.400 184.300 341.200 184.400 ;
        RECT 343.600 184.300 344.400 184.400 ;
        RECT 340.400 183.700 344.400 184.300 ;
        RECT 340.400 183.600 341.200 183.700 ;
        RECT 343.600 183.600 344.400 183.700 ;
        RECT 404.400 184.300 405.200 184.400 ;
        RECT 407.600 184.300 408.400 184.400 ;
        RECT 404.400 183.700 408.400 184.300 ;
        RECT 404.400 183.600 405.200 183.700 ;
        RECT 407.600 183.600 408.400 183.700 ;
        RECT 431.600 184.300 432.400 184.400 ;
        RECT 500.400 184.300 501.200 184.400 ;
        RECT 431.600 183.700 501.200 184.300 ;
        RECT 431.600 183.600 432.400 183.700 ;
        RECT 500.400 183.600 501.200 183.700 ;
        RECT 516.400 184.300 517.200 184.400 ;
        RECT 522.800 184.300 523.600 184.400 ;
        RECT 516.400 183.700 523.600 184.300 ;
        RECT 516.400 183.600 517.200 183.700 ;
        RECT 522.800 183.600 523.600 183.700 ;
        RECT 601.200 184.300 602.000 184.400 ;
        RECT 607.600 184.300 608.400 184.400 ;
        RECT 601.200 183.700 608.400 184.300 ;
        RECT 601.200 183.600 602.000 183.700 ;
        RECT 607.600 183.600 608.400 183.700 ;
        RECT 31.600 182.300 32.400 182.400 ;
        RECT 38.000 182.300 38.800 182.400 ;
        RECT 65.200 182.300 66.000 182.400 ;
        RECT 31.600 181.700 66.000 182.300 ;
        RECT 31.600 181.600 32.400 181.700 ;
        RECT 38.000 181.600 38.800 181.700 ;
        RECT 65.200 181.600 66.000 181.700 ;
        RECT 66.800 182.300 67.600 182.400 ;
        RECT 82.800 182.300 83.600 182.400 ;
        RECT 66.800 181.700 83.600 182.300 ;
        RECT 66.800 181.600 67.600 181.700 ;
        RECT 82.800 181.600 83.600 181.700 ;
        RECT 190.000 182.300 190.800 182.400 ;
        RECT 225.200 182.300 226.000 182.400 ;
        RECT 254.000 182.300 254.800 182.400 ;
        RECT 190.000 181.700 254.800 182.300 ;
        RECT 190.000 181.600 190.800 181.700 ;
        RECT 225.200 181.600 226.000 181.700 ;
        RECT 254.000 181.600 254.800 181.700 ;
        RECT 316.400 182.300 317.200 182.400 ;
        RECT 343.600 182.300 344.400 182.400 ;
        RECT 346.800 182.300 347.600 182.400 ;
        RECT 316.400 181.700 347.600 182.300 ;
        RECT 316.400 181.600 317.200 181.700 ;
        RECT 343.600 181.600 344.400 181.700 ;
        RECT 346.800 181.600 347.600 181.700 ;
        RECT 380.400 182.300 381.200 182.400 ;
        RECT 412.400 182.300 413.200 182.400 ;
        RECT 380.400 181.700 413.200 182.300 ;
        RECT 380.400 181.600 381.200 181.700 ;
        RECT 412.400 181.600 413.200 181.700 ;
        RECT 447.600 182.300 448.400 182.400 ;
        RECT 450.800 182.300 451.600 182.400 ;
        RECT 447.600 181.700 451.600 182.300 ;
        RECT 447.600 181.600 448.400 181.700 ;
        RECT 450.800 181.600 451.600 181.700 ;
        RECT 514.800 182.300 515.600 182.400 ;
        RECT 519.600 182.300 520.400 182.400 ;
        RECT 514.800 181.700 520.400 182.300 ;
        RECT 514.800 181.600 515.600 181.700 ;
        RECT 519.600 181.600 520.400 181.700 ;
        RECT 572.400 182.300 573.200 182.400 ;
        RECT 580.400 182.300 581.200 182.400 ;
        RECT 572.400 181.700 581.200 182.300 ;
        RECT 572.400 181.600 573.200 181.700 ;
        RECT 580.400 181.600 581.200 181.700 ;
        RECT 78.000 180.300 78.800 180.400 ;
        RECT 110.000 180.300 110.800 180.400 ;
        RECT 78.000 179.700 110.800 180.300 ;
        RECT 78.000 179.600 78.800 179.700 ;
        RECT 110.000 179.600 110.800 179.700 ;
        RECT 122.800 180.300 123.600 180.400 ;
        RECT 138.800 180.300 139.600 180.400 ;
        RECT 122.800 179.700 139.600 180.300 ;
        RECT 122.800 179.600 123.600 179.700 ;
        RECT 138.800 179.600 139.600 179.700 ;
        RECT 207.600 180.300 208.400 180.400 ;
        RECT 218.800 180.300 219.600 180.400 ;
        RECT 286.000 180.300 286.800 180.400 ;
        RECT 207.600 179.700 286.800 180.300 ;
        RECT 207.600 179.600 208.400 179.700 ;
        RECT 218.800 179.600 219.600 179.700 ;
        RECT 286.000 179.600 286.800 179.700 ;
        RECT 321.200 180.300 322.000 180.400 ;
        RECT 337.200 180.300 338.000 180.400 ;
        RECT 321.200 179.700 338.000 180.300 ;
        RECT 321.200 179.600 322.000 179.700 ;
        RECT 337.200 179.600 338.000 179.700 ;
        RECT 353.200 180.300 354.000 180.400 ;
        RECT 398.000 180.300 398.800 180.400 ;
        RECT 353.200 179.700 398.800 180.300 ;
        RECT 353.200 179.600 354.000 179.700 ;
        RECT 398.000 179.600 398.800 179.700 ;
        RECT 497.200 180.300 498.000 180.400 ;
        RECT 510.000 180.300 510.800 180.400 ;
        RECT 497.200 179.700 510.800 180.300 ;
        RECT 497.200 179.600 498.000 179.700 ;
        RECT 510.000 179.600 510.800 179.700 ;
        RECT 578.800 180.300 579.600 180.400 ;
        RECT 582.000 180.300 582.800 180.400 ;
        RECT 578.800 179.700 582.800 180.300 ;
        RECT 578.800 179.600 579.600 179.700 ;
        RECT 582.000 179.600 582.800 179.700 ;
        RECT 30.000 178.300 30.800 178.400 ;
        RECT 39.600 178.300 40.400 178.400 ;
        RECT 30.000 177.700 40.400 178.300 ;
        RECT 30.000 177.600 30.800 177.700 ;
        RECT 39.600 177.600 40.400 177.700 ;
        RECT 52.400 178.300 53.200 178.400 ;
        RECT 73.200 178.300 74.000 178.400 ;
        RECT 87.600 178.300 88.400 178.400 ;
        RECT 94.000 178.300 94.800 178.400 ;
        RECT 52.400 177.700 94.800 178.300 ;
        RECT 52.400 177.600 53.200 177.700 ;
        RECT 73.200 177.600 74.000 177.700 ;
        RECT 87.600 177.600 88.400 177.700 ;
        RECT 94.000 177.600 94.800 177.700 ;
        RECT 103.600 178.300 104.400 178.400 ;
        RECT 114.800 178.300 115.600 178.400 ;
        RECT 122.800 178.300 123.600 178.400 ;
        RECT 103.600 177.700 123.600 178.300 ;
        RECT 103.600 177.600 104.400 177.700 ;
        RECT 114.800 177.600 115.600 177.700 ;
        RECT 122.800 177.600 123.600 177.700 ;
        RECT 193.200 178.300 194.000 178.400 ;
        RECT 222.000 178.300 222.800 178.400 ;
        RECT 193.200 177.700 222.800 178.300 ;
        RECT 193.200 177.600 194.000 177.700 ;
        RECT 222.000 177.600 222.800 177.700 ;
        RECT 225.200 178.300 226.000 178.400 ;
        RECT 228.400 178.300 229.200 178.400 ;
        RECT 225.200 177.700 229.200 178.300 ;
        RECT 225.200 177.600 226.000 177.700 ;
        RECT 228.400 177.600 229.200 177.700 ;
        RECT 274.800 178.300 275.600 178.400 ;
        RECT 289.200 178.300 290.000 178.400 ;
        RECT 274.800 177.700 290.000 178.300 ;
        RECT 274.800 177.600 275.600 177.700 ;
        RECT 289.200 177.600 290.000 177.700 ;
        RECT 346.800 178.300 347.600 178.400 ;
        RECT 356.400 178.300 357.200 178.400 ;
        RECT 346.800 177.700 357.200 178.300 ;
        RECT 346.800 177.600 347.600 177.700 ;
        RECT 356.400 177.600 357.200 177.700 ;
        RECT 370.800 178.300 371.600 178.400 ;
        RECT 391.600 178.300 392.400 178.400 ;
        RECT 370.800 177.700 392.400 178.300 ;
        RECT 370.800 177.600 371.600 177.700 ;
        RECT 391.600 177.600 392.400 177.700 ;
        RECT 423.600 178.300 424.400 178.400 ;
        RECT 474.800 178.300 475.600 178.400 ;
        RECT 498.800 178.300 499.600 178.400 ;
        RECT 423.600 177.700 499.600 178.300 ;
        RECT 423.600 177.600 424.400 177.700 ;
        RECT 474.800 177.600 475.600 177.700 ;
        RECT 498.800 177.600 499.600 177.700 ;
        RECT 502.000 178.300 502.800 178.400 ;
        RECT 554.800 178.300 555.600 178.400 ;
        RECT 502.000 177.700 555.600 178.300 ;
        RECT 502.000 177.600 502.800 177.700 ;
        RECT 554.800 177.600 555.600 177.700 ;
        RECT 25.200 176.300 26.000 176.400 ;
        RECT 30.000 176.300 30.800 176.400 ;
        RECT 25.200 175.700 30.800 176.300 ;
        RECT 25.200 175.600 26.000 175.700 ;
        RECT 30.000 175.600 30.800 175.700 ;
        RECT 63.600 176.300 64.400 176.400 ;
        RECT 81.200 176.300 82.000 176.400 ;
        RECT 63.600 175.700 82.000 176.300 ;
        RECT 63.600 175.600 64.400 175.700 ;
        RECT 81.200 175.600 82.000 175.700 ;
        RECT 82.800 176.300 83.600 176.400 ;
        RECT 90.800 176.300 91.600 176.400 ;
        RECT 82.800 175.700 91.600 176.300 ;
        RECT 82.800 175.600 83.600 175.700 ;
        RECT 90.800 175.600 91.600 175.700 ;
        RECT 126.000 176.300 126.800 176.400 ;
        RECT 146.800 176.300 147.600 176.400 ;
        RECT 178.800 176.300 179.600 176.400 ;
        RECT 126.000 175.700 179.600 176.300 ;
        RECT 126.000 175.600 126.800 175.700 ;
        RECT 146.800 175.600 147.600 175.700 ;
        RECT 178.800 175.600 179.600 175.700 ;
        RECT 194.800 176.300 195.600 176.400 ;
        RECT 209.200 176.300 210.000 176.400 ;
        RECT 194.800 175.700 210.000 176.300 ;
        RECT 194.800 175.600 195.600 175.700 ;
        RECT 209.200 175.600 210.000 175.700 ;
        RECT 212.400 176.300 213.200 176.400 ;
        RECT 241.200 176.300 242.000 176.400 ;
        RECT 212.400 175.700 242.000 176.300 ;
        RECT 212.400 175.600 213.200 175.700 ;
        RECT 241.200 175.600 242.000 175.700 ;
        RECT 298.800 176.300 299.600 176.400 ;
        RECT 314.800 176.300 315.600 176.400 ;
        RECT 298.800 175.700 315.600 176.300 ;
        RECT 298.800 175.600 299.600 175.700 ;
        RECT 314.800 175.600 315.600 175.700 ;
        RECT 318.000 175.600 318.800 176.400 ;
        RECT 350.000 176.300 350.800 176.400 ;
        RECT 319.700 175.700 350.800 176.300 ;
        RECT 76.400 174.300 77.200 174.400 ;
        RECT 82.800 174.300 83.600 174.400 ;
        RECT 76.400 173.700 83.600 174.300 ;
        RECT 76.400 173.600 77.200 173.700 ;
        RECT 82.800 173.600 83.600 173.700 ;
        RECT 84.400 174.300 85.200 174.400 ;
        RECT 105.200 174.300 106.000 174.400 ;
        RECT 129.200 174.300 130.000 174.400 ;
        RECT 84.400 173.700 130.000 174.300 ;
        RECT 84.400 173.600 85.200 173.700 ;
        RECT 105.200 173.600 106.000 173.700 ;
        RECT 129.200 173.600 130.000 173.700 ;
        RECT 193.200 174.300 194.000 174.400 ;
        RECT 246.000 174.300 246.800 174.400 ;
        RECT 193.200 173.700 246.800 174.300 ;
        RECT 193.200 173.600 194.000 173.700 ;
        RECT 246.000 173.600 246.800 173.700 ;
        RECT 255.600 174.300 256.400 174.400 ;
        RECT 276.400 174.300 277.200 174.400 ;
        RECT 255.600 173.700 277.200 174.300 ;
        RECT 255.600 173.600 256.400 173.700 ;
        RECT 276.400 173.600 277.200 173.700 ;
        RECT 281.200 174.300 282.000 174.400 ;
        RECT 290.800 174.300 291.600 174.400 ;
        RECT 281.200 173.700 291.600 174.300 ;
        RECT 281.200 173.600 282.000 173.700 ;
        RECT 290.800 173.600 291.600 173.700 ;
        RECT 314.800 174.300 315.600 174.400 ;
        RECT 319.700 174.300 320.300 175.700 ;
        RECT 350.000 175.600 350.800 175.700 ;
        RECT 398.000 176.300 398.800 176.400 ;
        RECT 410.800 176.300 411.600 176.400 ;
        RECT 398.000 175.700 411.600 176.300 ;
        RECT 398.000 175.600 398.800 175.700 ;
        RECT 410.800 175.600 411.600 175.700 ;
        RECT 414.000 176.300 414.800 176.400 ;
        RECT 417.200 176.300 418.000 176.400 ;
        RECT 414.000 175.700 418.000 176.300 ;
        RECT 414.000 175.600 414.800 175.700 ;
        RECT 417.200 175.600 418.000 175.700 ;
        RECT 470.000 176.300 470.800 176.400 ;
        RECT 545.200 176.300 546.000 176.400 ;
        RECT 470.000 175.700 546.000 176.300 ;
        RECT 470.000 175.600 470.800 175.700 ;
        RECT 545.200 175.600 546.000 175.700 ;
        RECT 551.600 176.300 552.400 176.400 ;
        RECT 567.600 176.300 568.400 176.400 ;
        RECT 551.600 175.700 568.400 176.300 ;
        RECT 551.600 175.600 552.400 175.700 ;
        RECT 567.600 175.600 568.400 175.700 ;
        RECT 580.400 176.300 581.200 176.400 ;
        RECT 591.600 176.300 592.400 176.400 ;
        RECT 580.400 175.700 592.400 176.300 ;
        RECT 580.400 175.600 581.200 175.700 ;
        RECT 591.600 175.600 592.400 175.700 ;
        RECT 314.800 173.700 320.300 174.300 ;
        RECT 343.600 174.300 344.400 174.400 ;
        RECT 348.400 174.300 349.200 174.400 ;
        RECT 343.600 173.700 349.200 174.300 ;
        RECT 314.800 173.600 315.600 173.700 ;
        RECT 343.600 173.600 344.400 173.700 ;
        RECT 348.400 173.600 349.200 173.700 ;
        RECT 356.400 174.300 357.200 174.400 ;
        RECT 364.400 174.300 365.200 174.400 ;
        RECT 356.400 173.700 365.200 174.300 ;
        RECT 356.400 173.600 357.200 173.700 ;
        RECT 364.400 173.600 365.200 173.700 ;
        RECT 369.200 174.300 370.000 174.400 ;
        RECT 377.200 174.300 378.000 174.400 ;
        RECT 369.200 173.700 378.000 174.300 ;
        RECT 369.200 173.600 370.000 173.700 ;
        RECT 377.200 173.600 378.000 173.700 ;
        RECT 401.200 174.300 402.000 174.400 ;
        RECT 433.200 174.300 434.000 174.400 ;
        RECT 401.200 173.700 434.000 174.300 ;
        RECT 401.200 173.600 402.000 173.700 ;
        RECT 433.200 173.600 434.000 173.700 ;
        RECT 446.000 174.300 446.800 174.400 ;
        RECT 470.000 174.300 470.800 174.400 ;
        RECT 446.000 173.700 470.800 174.300 ;
        RECT 446.000 173.600 446.800 173.700 ;
        RECT 470.000 173.600 470.800 173.700 ;
        RECT 482.800 174.300 483.600 174.400 ;
        RECT 492.400 174.300 493.200 174.400 ;
        RECT 482.800 173.700 493.200 174.300 ;
        RECT 482.800 173.600 483.600 173.700 ;
        RECT 492.400 173.600 493.200 173.700 ;
        RECT 506.800 174.300 507.600 174.400 ;
        RECT 521.200 174.300 522.000 174.400 ;
        RECT 506.800 173.700 522.000 174.300 ;
        RECT 506.800 173.600 507.600 173.700 ;
        RECT 521.200 173.600 522.000 173.700 ;
        RECT 529.200 174.300 530.000 174.400 ;
        RECT 543.600 174.300 544.400 174.400 ;
        RECT 551.600 174.300 552.400 174.400 ;
        RECT 529.200 173.700 552.400 174.300 ;
        RECT 529.200 173.600 530.000 173.700 ;
        RECT 543.600 173.600 544.400 173.700 ;
        RECT 551.600 173.600 552.400 173.700 ;
        RECT 585.200 174.300 586.000 174.400 ;
        RECT 599.600 174.300 600.400 174.400 ;
        RECT 585.200 173.700 600.400 174.300 ;
        RECT 585.200 173.600 586.000 173.700 ;
        RECT 599.600 173.600 600.400 173.700 ;
        RECT 9.200 172.300 10.000 172.400 ;
        RECT 20.400 172.300 21.200 172.400 ;
        RECT 9.200 171.700 21.200 172.300 ;
        RECT 9.200 171.600 10.000 171.700 ;
        RECT 20.400 171.600 21.200 171.700 ;
        RECT 23.600 172.300 24.400 172.400 ;
        RECT 31.600 172.300 32.400 172.400 ;
        RECT 23.600 171.700 32.400 172.300 ;
        RECT 23.600 171.600 24.400 171.700 ;
        RECT 31.600 171.600 32.400 171.700 ;
        RECT 79.600 172.300 80.400 172.400 ;
        RECT 81.200 172.300 82.000 172.400 ;
        RECT 113.200 172.300 114.000 172.400 ;
        RECT 79.600 171.700 114.000 172.300 ;
        RECT 79.600 171.600 80.400 171.700 ;
        RECT 81.200 171.600 82.000 171.700 ;
        RECT 113.200 171.600 114.000 171.700 ;
        RECT 121.200 172.300 122.000 172.400 ;
        RECT 129.200 172.300 130.000 172.400 ;
        RECT 140.400 172.300 141.200 172.400 ;
        RECT 156.400 172.300 157.200 172.400 ;
        RECT 121.200 171.700 157.200 172.300 ;
        RECT 121.200 171.600 122.000 171.700 ;
        RECT 129.200 171.600 130.000 171.700 ;
        RECT 140.400 171.600 141.200 171.700 ;
        RECT 156.400 171.600 157.200 171.700 ;
        RECT 180.400 172.300 181.200 172.400 ;
        RECT 182.000 172.300 182.800 172.400 ;
        RECT 185.200 172.300 186.000 172.400 ;
        RECT 180.400 171.700 186.000 172.300 ;
        RECT 180.400 171.600 181.200 171.700 ;
        RECT 182.000 171.600 182.800 171.700 ;
        RECT 185.200 171.600 186.000 171.700 ;
        RECT 201.200 172.300 202.000 172.400 ;
        RECT 228.400 172.300 229.200 172.400 ;
        RECT 201.200 171.700 229.200 172.300 ;
        RECT 201.200 171.600 202.000 171.700 ;
        RECT 228.400 171.600 229.200 171.700 ;
        RECT 326.000 172.300 326.800 172.400 ;
        RECT 332.400 172.300 333.200 172.400 ;
        RECT 326.000 171.700 333.200 172.300 ;
        RECT 326.000 171.600 326.800 171.700 ;
        RECT 332.400 171.600 333.200 171.700 ;
        RECT 345.200 172.300 346.000 172.400 ;
        RECT 364.400 172.300 365.200 172.400 ;
        RECT 345.200 171.700 365.200 172.300 ;
        RECT 345.200 171.600 346.000 171.700 ;
        RECT 364.400 171.600 365.200 171.700 ;
        RECT 369.200 172.300 370.000 172.400 ;
        RECT 431.600 172.300 432.400 172.400 ;
        RECT 369.200 171.700 432.400 172.300 ;
        RECT 369.200 171.600 370.000 171.700 ;
        RECT 431.600 171.600 432.400 171.700 ;
        RECT 433.200 172.300 434.000 172.400 ;
        RECT 449.200 172.300 450.000 172.400 ;
        RECT 433.200 171.700 450.000 172.300 ;
        RECT 433.200 171.600 434.000 171.700 ;
        RECT 449.200 171.600 450.000 171.700 ;
        RECT 471.600 172.300 472.400 172.400 ;
        RECT 478.000 172.300 478.800 172.400 ;
        RECT 471.600 171.700 478.800 172.300 ;
        RECT 471.600 171.600 472.400 171.700 ;
        RECT 478.000 171.600 478.800 171.700 ;
        RECT 503.600 172.300 504.400 172.400 ;
        RECT 527.600 172.300 528.400 172.400 ;
        RECT 503.600 171.700 528.400 172.300 ;
        RECT 503.600 171.600 504.400 171.700 ;
        RECT 527.600 171.600 528.400 171.700 ;
        RECT 537.200 172.300 538.000 172.400 ;
        RECT 558.000 172.300 558.800 172.400 ;
        RECT 537.200 171.700 558.800 172.300 ;
        RECT 537.200 171.600 538.000 171.700 ;
        RECT 558.000 171.600 558.800 171.700 ;
        RECT 566.000 172.300 566.800 172.400 ;
        RECT 574.000 172.300 574.800 172.400 ;
        RECT 566.000 171.700 574.800 172.300 ;
        RECT 566.000 171.600 566.800 171.700 ;
        RECT 574.000 171.600 574.800 171.700 ;
        RECT 20.400 170.300 21.200 170.400 ;
        RECT 23.600 170.300 24.400 170.400 ;
        RECT 20.400 169.700 24.400 170.300 ;
        RECT 20.400 169.600 21.200 169.700 ;
        RECT 23.600 169.600 24.400 169.700 ;
        RECT 65.200 170.300 66.000 170.400 ;
        RECT 82.800 170.300 83.600 170.400 ;
        RECT 65.200 169.700 83.600 170.300 ;
        RECT 65.200 169.600 66.000 169.700 ;
        RECT 82.800 169.600 83.600 169.700 ;
        RECT 137.200 170.300 138.000 170.400 ;
        RECT 196.400 170.300 197.200 170.400 ;
        RECT 199.600 170.300 200.400 170.400 ;
        RECT 137.200 169.700 200.400 170.300 ;
        RECT 137.200 169.600 138.000 169.700 ;
        RECT 196.400 169.600 197.200 169.700 ;
        RECT 199.600 169.600 200.400 169.700 ;
        RECT 201.200 170.300 202.000 170.400 ;
        RECT 209.200 170.300 210.000 170.400 ;
        RECT 215.600 170.300 216.400 170.400 ;
        RECT 201.200 169.700 216.400 170.300 ;
        RECT 201.200 169.600 202.000 169.700 ;
        RECT 209.200 169.600 210.000 169.700 ;
        RECT 215.600 169.600 216.400 169.700 ;
        RECT 334.000 170.300 334.800 170.400 ;
        RECT 340.400 170.300 341.200 170.400 ;
        RECT 342.000 170.300 342.800 170.400 ;
        RECT 334.000 169.700 342.800 170.300 ;
        RECT 334.000 169.600 334.800 169.700 ;
        RECT 340.400 169.600 341.200 169.700 ;
        RECT 342.000 169.600 342.800 169.700 ;
        RECT 354.800 170.300 355.600 170.400 ;
        RECT 362.800 170.300 363.600 170.400 ;
        RECT 374.000 170.300 374.800 170.400 ;
        RECT 354.800 169.700 374.800 170.300 ;
        RECT 354.800 169.600 355.600 169.700 ;
        RECT 362.800 169.600 363.600 169.700 ;
        RECT 374.000 169.600 374.800 169.700 ;
        RECT 380.400 170.300 381.200 170.400 ;
        RECT 382.000 170.300 382.800 170.400 ;
        RECT 380.400 169.700 382.800 170.300 ;
        RECT 380.400 169.600 381.200 169.700 ;
        RECT 382.000 169.600 382.800 169.700 ;
        RECT 385.200 170.300 386.000 170.400 ;
        RECT 409.200 170.300 410.000 170.400 ;
        RECT 417.200 170.300 418.000 170.400 ;
        RECT 385.200 169.700 418.000 170.300 ;
        RECT 385.200 169.600 386.000 169.700 ;
        RECT 409.200 169.600 410.000 169.700 ;
        RECT 417.200 169.600 418.000 169.700 ;
        RECT 444.400 170.300 445.200 170.400 ;
        RECT 452.400 170.300 453.200 170.400 ;
        RECT 444.400 169.700 453.200 170.300 ;
        RECT 444.400 169.600 445.200 169.700 ;
        RECT 452.400 169.600 453.200 169.700 ;
        RECT 465.200 170.300 466.000 170.400 ;
        RECT 474.800 170.300 475.600 170.400 ;
        RECT 465.200 169.700 475.600 170.300 ;
        RECT 465.200 169.600 466.000 169.700 ;
        RECT 474.800 169.600 475.600 169.700 ;
        RECT 476.400 170.300 477.200 170.400 ;
        RECT 489.200 170.300 490.000 170.400 ;
        RECT 476.400 169.700 490.000 170.300 ;
        RECT 476.400 169.600 477.200 169.700 ;
        RECT 489.200 169.600 490.000 169.700 ;
        RECT 511.600 170.300 512.400 170.400 ;
        RECT 519.600 170.300 520.400 170.400 ;
        RECT 511.600 169.700 520.400 170.300 ;
        RECT 511.600 169.600 512.400 169.700 ;
        RECT 519.600 169.600 520.400 169.700 ;
        RECT 524.400 170.300 525.200 170.400 ;
        RECT 534.000 170.300 534.800 170.400 ;
        RECT 545.200 170.300 546.000 170.400 ;
        RECT 524.400 169.700 546.000 170.300 ;
        RECT 524.400 169.600 525.200 169.700 ;
        RECT 534.000 169.600 534.800 169.700 ;
        RECT 545.200 169.600 546.000 169.700 ;
        RECT 556.400 170.300 557.200 170.400 ;
        RECT 562.800 170.300 563.600 170.400 ;
        RECT 556.400 169.700 563.600 170.300 ;
        RECT 556.400 169.600 557.200 169.700 ;
        RECT 562.800 169.600 563.600 169.700 ;
        RECT 564.400 170.300 565.200 170.400 ;
        RECT 599.600 170.300 600.400 170.400 ;
        RECT 564.400 169.700 600.400 170.300 ;
        RECT 564.400 169.600 565.200 169.700 ;
        RECT 599.600 169.600 600.400 169.700 ;
        RECT 18.800 168.300 19.600 168.400 ;
        RECT 20.400 168.300 21.200 168.400 ;
        RECT 28.400 168.300 29.200 168.400 ;
        RECT 18.800 167.700 29.200 168.300 ;
        RECT 18.800 167.600 19.600 167.700 ;
        RECT 20.400 167.600 21.200 167.700 ;
        RECT 28.400 167.600 29.200 167.700 ;
        RECT 41.200 168.300 42.000 168.400 ;
        RECT 135.600 168.300 136.400 168.400 ;
        RECT 158.000 168.300 158.800 168.400 ;
        RECT 41.200 167.700 158.800 168.300 ;
        RECT 41.200 167.600 42.000 167.700 ;
        RECT 135.600 167.600 136.400 167.700 ;
        RECT 158.000 167.600 158.800 167.700 ;
        RECT 167.600 168.300 168.400 168.400 ;
        RECT 177.200 168.300 178.000 168.400 ;
        RECT 225.200 168.300 226.000 168.400 ;
        RECT 167.600 167.700 226.000 168.300 ;
        RECT 167.600 167.600 168.400 167.700 ;
        RECT 177.200 167.600 178.000 167.700 ;
        RECT 225.200 167.600 226.000 167.700 ;
        RECT 351.600 168.300 352.400 168.400 ;
        RECT 361.200 168.300 362.000 168.400 ;
        RECT 351.600 167.700 362.000 168.300 ;
        RECT 351.600 167.600 352.400 167.700 ;
        RECT 361.200 167.600 362.000 167.700 ;
        RECT 415.600 168.300 416.400 168.400 ;
        RECT 420.400 168.300 421.200 168.400 ;
        RECT 446.000 168.300 446.800 168.400 ;
        RECT 415.600 167.700 446.800 168.300 ;
        RECT 415.600 167.600 416.400 167.700 ;
        RECT 420.400 167.600 421.200 167.700 ;
        RECT 446.000 167.600 446.800 167.700 ;
        RECT 452.400 168.300 453.200 168.400 ;
        RECT 457.200 168.300 458.000 168.400 ;
        RECT 452.400 167.700 458.000 168.300 ;
        RECT 452.400 167.600 453.200 167.700 ;
        RECT 457.200 167.600 458.000 167.700 ;
        RECT 484.400 167.600 485.200 168.400 ;
        RECT 486.000 168.300 486.800 168.400 ;
        RECT 492.400 168.300 493.200 168.400 ;
        RECT 511.700 168.300 512.300 169.600 ;
        RECT 486.000 167.700 512.300 168.300 ;
        RECT 529.200 168.300 530.000 168.400 ;
        RECT 542.000 168.300 542.800 168.400 ;
        RECT 529.200 167.700 542.800 168.300 ;
        RECT 486.000 167.600 486.800 167.700 ;
        RECT 492.400 167.600 493.200 167.700 ;
        RECT 529.200 167.600 530.000 167.700 ;
        RECT 542.000 167.600 542.800 167.700 ;
        RECT 559.600 168.300 560.400 168.400 ;
        RECT 562.800 168.300 563.600 168.400 ;
        RECT 564.400 168.300 565.200 168.400 ;
        RECT 559.600 167.700 565.200 168.300 ;
        RECT 559.600 167.600 560.400 167.700 ;
        RECT 562.800 167.600 563.600 167.700 ;
        RECT 564.400 167.600 565.200 167.700 ;
        RECT 567.600 168.300 568.400 168.400 ;
        RECT 599.600 168.300 600.400 168.400 ;
        RECT 602.800 168.300 603.600 168.400 ;
        RECT 567.600 167.700 603.600 168.300 ;
        RECT 567.600 167.600 568.400 167.700 ;
        RECT 599.600 167.600 600.400 167.700 ;
        RECT 602.800 167.600 603.600 167.700 ;
        RECT 78.000 166.300 78.800 166.400 ;
        RECT 98.800 166.300 99.600 166.400 ;
        RECT 78.000 165.700 99.600 166.300 ;
        RECT 78.000 165.600 78.800 165.700 ;
        RECT 98.800 165.600 99.600 165.700 ;
        RECT 106.800 166.300 107.600 166.400 ;
        RECT 142.000 166.300 142.800 166.400 ;
        RECT 151.600 166.300 152.400 166.400 ;
        RECT 106.800 165.700 152.400 166.300 ;
        RECT 106.800 165.600 107.600 165.700 ;
        RECT 142.000 165.600 142.800 165.700 ;
        RECT 151.600 165.600 152.400 165.700 ;
        RECT 318.000 166.300 318.800 166.400 ;
        RECT 340.400 166.300 341.200 166.400 ;
        RECT 380.400 166.300 381.200 166.400 ;
        RECT 318.000 165.700 381.200 166.300 ;
        RECT 318.000 165.600 318.800 165.700 ;
        RECT 340.400 165.600 341.200 165.700 ;
        RECT 380.400 165.600 381.200 165.700 ;
        RECT 454.000 166.300 454.800 166.400 ;
        RECT 468.400 166.300 469.200 166.400 ;
        RECT 482.800 166.300 483.600 166.400 ;
        RECT 454.000 165.700 483.600 166.300 ;
        RECT 454.000 165.600 454.800 165.700 ;
        RECT 468.400 165.600 469.200 165.700 ;
        RECT 482.800 165.600 483.600 165.700 ;
        RECT 502.000 166.300 502.800 166.400 ;
        RECT 519.600 166.300 520.400 166.400 ;
        RECT 502.000 165.700 520.400 166.300 ;
        RECT 502.000 165.600 502.800 165.700 ;
        RECT 519.600 165.600 520.400 165.700 ;
        RECT 142.000 164.300 142.800 164.400 ;
        RECT 206.000 164.300 206.800 164.400 ;
        RECT 142.000 163.700 206.800 164.300 ;
        RECT 142.000 163.600 142.800 163.700 ;
        RECT 206.000 163.600 206.800 163.700 ;
        RECT 407.600 164.300 408.400 164.400 ;
        RECT 529.200 164.300 530.000 164.400 ;
        RECT 407.600 163.700 530.000 164.300 ;
        RECT 407.600 163.600 408.400 163.700 ;
        RECT 529.200 163.600 530.000 163.700 ;
        RECT 161.200 162.300 162.000 162.400 ;
        RECT 191.600 162.300 192.400 162.400 ;
        RECT 161.200 161.700 192.400 162.300 ;
        RECT 161.200 161.600 162.000 161.700 ;
        RECT 191.600 161.600 192.400 161.700 ;
        RECT 406.000 162.300 406.800 162.400 ;
        RECT 410.800 162.300 411.600 162.400 ;
        RECT 406.000 161.700 411.600 162.300 ;
        RECT 406.000 161.600 406.800 161.700 ;
        RECT 410.800 161.600 411.600 161.700 ;
        RECT 26.800 160.300 27.600 160.400 ;
        RECT 42.800 160.300 43.600 160.400 ;
        RECT 57.200 160.300 58.000 160.400 ;
        RECT 140.400 160.300 141.200 160.400 ;
        RECT 26.800 159.700 141.200 160.300 ;
        RECT 26.800 159.600 27.600 159.700 ;
        RECT 42.800 159.600 43.600 159.700 ;
        RECT 57.200 159.600 58.000 159.700 ;
        RECT 140.400 159.600 141.200 159.700 ;
        RECT 170.800 159.600 171.600 160.400 ;
        RECT 241.200 160.300 242.000 160.400 ;
        RECT 258.800 160.300 259.600 160.400 ;
        RECT 281.200 160.300 282.000 160.400 ;
        RECT 284.400 160.300 285.200 160.400 ;
        RECT 241.200 159.700 285.200 160.300 ;
        RECT 241.200 159.600 242.000 159.700 ;
        RECT 258.800 159.600 259.600 159.700 ;
        RECT 281.200 159.600 282.000 159.700 ;
        RECT 284.400 159.600 285.200 159.700 ;
        RECT 297.200 160.300 298.000 160.400 ;
        RECT 319.600 160.300 320.400 160.400 ;
        RECT 297.200 159.700 320.400 160.300 ;
        RECT 297.200 159.600 298.000 159.700 ;
        RECT 319.600 159.600 320.400 159.700 ;
        RECT 470.000 160.300 470.800 160.400 ;
        RECT 506.800 160.300 507.600 160.400 ;
        RECT 470.000 159.700 507.600 160.300 ;
        RECT 470.000 159.600 470.800 159.700 ;
        RECT 506.800 159.600 507.600 159.700 ;
        RECT 513.200 160.300 514.000 160.400 ;
        RECT 538.800 160.300 539.600 160.400 ;
        RECT 551.600 160.300 552.400 160.400 ;
        RECT 513.200 159.700 552.400 160.300 ;
        RECT 513.200 159.600 514.000 159.700 ;
        RECT 538.800 159.600 539.600 159.700 ;
        RECT 551.600 159.600 552.400 159.700 ;
        RECT 582.000 160.300 582.800 160.400 ;
        RECT 585.200 160.300 586.000 160.400 ;
        RECT 582.000 159.700 586.000 160.300 ;
        RECT 582.000 159.600 582.800 159.700 ;
        RECT 585.200 159.600 586.000 159.700 ;
        RECT 596.400 160.300 597.200 160.400 ;
        RECT 598.000 160.300 598.800 160.400 ;
        RECT 596.400 159.700 598.800 160.300 ;
        RECT 596.400 159.600 597.200 159.700 ;
        RECT 598.000 159.600 598.800 159.700 ;
        RECT 28.400 158.300 29.200 158.400 ;
        RECT 103.600 158.300 104.400 158.400 ;
        RECT 28.400 157.700 104.400 158.300 ;
        RECT 28.400 157.600 29.200 157.700 ;
        RECT 103.600 157.600 104.400 157.700 ;
        RECT 151.600 158.300 152.400 158.400 ;
        RECT 170.900 158.300 171.500 159.600 ;
        RECT 151.600 157.700 171.500 158.300 ;
        RECT 404.400 158.300 405.200 158.400 ;
        RECT 409.200 158.300 410.000 158.400 ;
        RECT 404.400 157.700 410.000 158.300 ;
        RECT 151.600 157.600 152.400 157.700 ;
        RECT 404.400 157.600 405.200 157.700 ;
        RECT 409.200 157.600 410.000 157.700 ;
        RECT 412.400 158.300 413.200 158.400 ;
        RECT 479.600 158.300 480.400 158.400 ;
        RECT 412.400 157.700 480.400 158.300 ;
        RECT 412.400 157.600 413.200 157.700 ;
        RECT 479.600 157.600 480.400 157.700 ;
        RECT 484.400 158.300 485.200 158.400 ;
        RECT 518.000 158.300 518.800 158.400 ;
        RECT 484.400 157.700 518.800 158.300 ;
        RECT 484.400 157.600 485.200 157.700 ;
        RECT 518.000 157.600 518.800 157.700 ;
        RECT 68.400 156.300 69.200 156.400 ;
        RECT 73.200 156.300 74.000 156.400 ;
        RECT 68.400 155.700 74.000 156.300 ;
        RECT 68.400 155.600 69.200 155.700 ;
        RECT 73.200 155.600 74.000 155.700 ;
        RECT 94.000 156.300 94.800 156.400 ;
        RECT 106.800 156.300 107.600 156.400 ;
        RECT 94.000 155.700 107.600 156.300 ;
        RECT 94.000 155.600 94.800 155.700 ;
        RECT 106.800 155.600 107.600 155.700 ;
        RECT 111.600 156.300 112.400 156.400 ;
        RECT 114.800 156.300 115.600 156.400 ;
        RECT 111.600 155.700 115.600 156.300 ;
        RECT 111.600 155.600 112.400 155.700 ;
        RECT 114.800 155.600 115.600 155.700 ;
        RECT 116.400 156.300 117.200 156.400 ;
        RECT 122.800 156.300 123.600 156.400 ;
        RECT 116.400 155.700 123.600 156.300 ;
        RECT 116.400 155.600 117.200 155.700 ;
        RECT 122.800 155.600 123.600 155.700 ;
        RECT 134.000 156.300 134.800 156.400 ;
        RECT 135.600 156.300 136.400 156.400 ;
        RECT 134.000 155.700 136.400 156.300 ;
        RECT 134.000 155.600 134.800 155.700 ;
        RECT 135.600 155.600 136.400 155.700 ;
        RECT 140.400 156.300 141.200 156.400 ;
        RECT 161.200 156.300 162.000 156.400 ;
        RECT 140.400 155.700 162.000 156.300 ;
        RECT 140.400 155.600 141.200 155.700 ;
        RECT 161.200 155.600 162.000 155.700 ;
        RECT 223.600 156.300 224.400 156.400 ;
        RECT 257.200 156.300 258.000 156.400 ;
        RECT 292.400 156.300 293.200 156.400 ;
        RECT 223.600 155.700 293.200 156.300 ;
        RECT 223.600 155.600 224.400 155.700 ;
        RECT 257.200 155.600 258.000 155.700 ;
        RECT 292.400 155.600 293.200 155.700 ;
        RECT 356.400 156.300 357.200 156.400 ;
        RECT 370.800 156.300 371.600 156.400 ;
        RECT 356.400 155.700 371.600 156.300 ;
        RECT 356.400 155.600 357.200 155.700 ;
        RECT 370.800 155.600 371.600 155.700 ;
        RECT 390.000 156.300 390.800 156.400 ;
        RECT 402.800 156.300 403.600 156.400 ;
        RECT 390.000 155.700 403.600 156.300 ;
        RECT 390.000 155.600 390.800 155.700 ;
        RECT 402.800 155.600 403.600 155.700 ;
        RECT 428.400 156.300 429.200 156.400 ;
        RECT 460.400 156.300 461.200 156.400 ;
        RECT 428.400 155.700 461.200 156.300 ;
        RECT 428.400 155.600 429.200 155.700 ;
        RECT 460.400 155.600 461.200 155.700 ;
        RECT 466.800 156.300 467.600 156.400 ;
        RECT 470.000 156.300 470.800 156.400 ;
        RECT 466.800 155.700 470.800 156.300 ;
        RECT 466.800 155.600 467.600 155.700 ;
        RECT 470.000 155.600 470.800 155.700 ;
        RECT 484.400 156.300 485.200 156.400 ;
        RECT 524.400 156.300 525.200 156.400 ;
        RECT 484.400 155.700 525.200 156.300 ;
        RECT 484.400 155.600 485.200 155.700 ;
        RECT 524.400 155.600 525.200 155.700 ;
        RECT 545.200 156.300 546.000 156.400 ;
        RECT 575.600 156.300 576.400 156.400 ;
        RECT 545.200 155.700 576.400 156.300 ;
        RECT 545.200 155.600 546.000 155.700 ;
        RECT 575.600 155.600 576.400 155.700 ;
        RECT 26.800 154.300 27.600 154.400 ;
        RECT 38.000 154.300 38.800 154.400 ;
        RECT 26.800 153.700 38.800 154.300 ;
        RECT 26.800 153.600 27.600 153.700 ;
        RECT 38.000 153.600 38.800 153.700 ;
        RECT 55.600 154.300 56.400 154.400 ;
        RECT 63.600 154.300 64.400 154.400 ;
        RECT 89.200 154.300 90.000 154.400 ;
        RECT 55.600 153.700 90.000 154.300 ;
        RECT 55.600 153.600 56.400 153.700 ;
        RECT 63.600 153.600 64.400 153.700 ;
        RECT 89.200 153.600 90.000 153.700 ;
        RECT 111.600 154.300 112.400 154.400 ;
        RECT 129.200 154.300 130.000 154.400 ;
        RECT 111.600 153.700 130.000 154.300 ;
        RECT 111.600 153.600 112.400 153.700 ;
        RECT 129.200 153.600 130.000 153.700 ;
        RECT 271.600 154.300 272.400 154.400 ;
        RECT 278.000 154.300 278.800 154.400 ;
        RECT 271.600 153.700 278.800 154.300 ;
        RECT 271.600 153.600 272.400 153.700 ;
        RECT 278.000 153.600 278.800 153.700 ;
        RECT 351.600 154.300 352.400 154.400 ;
        RECT 358.000 154.300 358.800 154.400 ;
        RECT 366.000 154.300 366.800 154.400 ;
        RECT 351.600 153.700 366.800 154.300 ;
        RECT 351.600 153.600 352.400 153.700 ;
        RECT 358.000 153.600 358.800 153.700 ;
        RECT 366.000 153.600 366.800 153.700 ;
        RECT 398.000 154.300 398.800 154.400 ;
        RECT 404.400 154.300 405.200 154.400 ;
        RECT 398.000 153.700 405.200 154.300 ;
        RECT 398.000 153.600 398.800 153.700 ;
        RECT 404.400 153.600 405.200 153.700 ;
        RECT 450.800 154.300 451.600 154.400 ;
        RECT 455.600 154.300 456.400 154.400 ;
        RECT 450.800 153.700 456.400 154.300 ;
        RECT 450.800 153.600 451.600 153.700 ;
        RECT 455.600 153.600 456.400 153.700 ;
        RECT 487.600 154.300 488.400 154.400 ;
        RECT 505.200 154.300 506.000 154.400 ;
        RECT 487.600 153.700 506.000 154.300 ;
        RECT 487.600 153.600 488.400 153.700 ;
        RECT 505.200 153.600 506.000 153.700 ;
        RECT 36.400 151.600 37.200 152.400 ;
        RECT 46.000 152.300 46.800 152.400 ;
        RECT 50.800 152.300 51.600 152.400 ;
        RECT 78.000 152.300 78.800 152.400 ;
        RECT 46.000 151.700 78.800 152.300 ;
        RECT 46.000 151.600 46.800 151.700 ;
        RECT 50.800 151.600 51.600 151.700 ;
        RECT 78.000 151.600 78.800 151.700 ;
        RECT 95.600 152.300 96.400 152.400 ;
        RECT 102.000 152.300 102.800 152.400 ;
        RECT 95.600 151.700 102.800 152.300 ;
        RECT 95.600 151.600 96.400 151.700 ;
        RECT 102.000 151.600 102.800 151.700 ;
        RECT 108.400 152.300 109.200 152.400 ;
        RECT 116.400 152.300 117.200 152.400 ;
        RECT 108.400 151.700 117.200 152.300 ;
        RECT 108.400 151.600 109.200 151.700 ;
        RECT 116.400 151.600 117.200 151.700 ;
        RECT 130.800 152.300 131.600 152.400 ;
        RECT 214.000 152.300 214.800 152.400 ;
        RECT 260.400 152.300 261.200 152.400 ;
        RECT 130.800 151.700 261.200 152.300 ;
        RECT 130.800 151.600 131.600 151.700 ;
        RECT 214.000 151.600 214.800 151.700 ;
        RECT 260.400 151.600 261.200 151.700 ;
        RECT 370.800 152.300 371.600 152.400 ;
        RECT 377.200 152.300 378.000 152.400 ;
        RECT 385.200 152.300 386.000 152.400 ;
        RECT 370.800 151.700 378.000 152.300 ;
        RECT 370.800 151.600 371.600 151.700 ;
        RECT 377.200 151.600 378.000 151.700 ;
        RECT 378.900 151.700 386.000 152.300 ;
        RECT 7.600 150.300 8.400 150.400 ;
        RECT 33.200 150.300 34.000 150.400 ;
        RECT 7.600 149.700 34.000 150.300 ;
        RECT 7.600 149.600 8.400 149.700 ;
        RECT 33.200 149.600 34.000 149.700 ;
        RECT 39.600 150.300 40.400 150.400 ;
        RECT 63.600 150.300 64.400 150.400 ;
        RECT 39.600 149.700 64.400 150.300 ;
        RECT 39.600 149.600 40.400 149.700 ;
        RECT 63.600 149.600 64.400 149.700 ;
        RECT 66.800 150.300 67.600 150.400 ;
        RECT 76.400 150.300 77.200 150.400 ;
        RECT 66.800 149.700 77.200 150.300 ;
        RECT 66.800 149.600 67.600 149.700 ;
        RECT 76.400 149.600 77.200 149.700 ;
        RECT 92.400 150.300 93.200 150.400 ;
        RECT 105.200 150.300 106.000 150.400 ;
        RECT 92.400 149.700 106.000 150.300 ;
        RECT 92.400 149.600 93.200 149.700 ;
        RECT 105.200 149.600 106.000 149.700 ;
        RECT 118.000 150.300 118.800 150.400 ;
        RECT 127.600 150.300 128.400 150.400 ;
        RECT 118.000 149.700 128.400 150.300 ;
        RECT 118.000 149.600 118.800 149.700 ;
        RECT 127.600 149.600 128.400 149.700 ;
        RECT 201.200 150.300 202.000 150.400 ;
        RECT 204.400 150.300 205.200 150.400 ;
        RECT 214.000 150.300 214.800 150.400 ;
        RECT 220.400 150.300 221.200 150.400 ;
        RECT 252.400 150.300 253.200 150.400 ;
        RECT 201.200 149.700 253.200 150.300 ;
        RECT 201.200 149.600 202.000 149.700 ;
        RECT 204.400 149.600 205.200 149.700 ;
        RECT 214.000 149.600 214.800 149.700 ;
        RECT 220.400 149.600 221.200 149.700 ;
        RECT 252.400 149.600 253.200 149.700 ;
        RECT 310.000 150.300 310.800 150.400 ;
        RECT 311.600 150.300 312.400 150.400 ;
        RECT 310.000 149.700 312.400 150.300 ;
        RECT 310.000 149.600 310.800 149.700 ;
        RECT 311.600 149.600 312.400 149.700 ;
        RECT 343.600 150.300 344.400 150.400 ;
        RECT 359.600 150.300 360.400 150.400 ;
        RECT 343.600 149.700 360.400 150.300 ;
        RECT 343.600 149.600 344.400 149.700 ;
        RECT 359.600 149.600 360.400 149.700 ;
        RECT 375.600 150.300 376.400 150.400 ;
        RECT 378.900 150.300 379.500 151.700 ;
        RECT 385.200 151.600 386.000 151.700 ;
        RECT 388.400 152.300 389.200 152.400 ;
        RECT 396.400 152.300 397.200 152.400 ;
        RECT 388.400 151.700 397.200 152.300 ;
        RECT 388.400 151.600 389.200 151.700 ;
        RECT 396.400 151.600 397.200 151.700 ;
        RECT 401.200 152.300 402.000 152.400 ;
        RECT 414.000 152.300 414.800 152.400 ;
        RECT 428.400 152.300 429.200 152.400 ;
        RECT 401.200 151.700 429.200 152.300 ;
        RECT 401.200 151.600 402.000 151.700 ;
        RECT 414.000 151.600 414.800 151.700 ;
        RECT 428.400 151.600 429.200 151.700 ;
        RECT 431.600 152.300 432.400 152.400 ;
        RECT 447.600 152.300 448.400 152.400 ;
        RECT 431.600 151.700 448.400 152.300 ;
        RECT 431.600 151.600 432.400 151.700 ;
        RECT 447.600 151.600 448.400 151.700 ;
        RECT 449.200 152.300 450.000 152.400 ;
        RECT 450.800 152.300 451.600 152.400 ;
        RECT 449.200 151.700 451.600 152.300 ;
        RECT 449.200 151.600 450.000 151.700 ;
        RECT 450.800 151.600 451.600 151.700 ;
        RECT 489.200 152.300 490.000 152.400 ;
        RECT 510.000 152.300 510.800 152.400 ;
        RECT 516.400 152.300 517.200 152.400 ;
        RECT 489.200 151.700 517.200 152.300 ;
        RECT 489.200 151.600 490.000 151.700 ;
        RECT 510.000 151.600 510.800 151.700 ;
        RECT 516.400 151.600 517.200 151.700 ;
        RECT 375.600 149.700 379.500 150.300 ;
        RECT 385.200 150.300 386.000 150.400 ;
        RECT 393.200 150.300 394.000 150.400 ;
        RECT 385.200 149.700 394.000 150.300 ;
        RECT 375.600 149.600 376.400 149.700 ;
        RECT 385.200 149.600 386.000 149.700 ;
        RECT 393.200 149.600 394.000 149.700 ;
        RECT 399.600 150.300 400.400 150.400 ;
        RECT 406.000 150.300 406.800 150.400 ;
        RECT 399.600 149.700 406.800 150.300 ;
        RECT 399.600 149.600 400.400 149.700 ;
        RECT 406.000 149.600 406.800 149.700 ;
        RECT 430.000 150.300 430.800 150.400 ;
        RECT 441.200 150.300 442.000 150.400 ;
        RECT 430.000 149.700 442.000 150.300 ;
        RECT 430.000 149.600 430.800 149.700 ;
        RECT 441.200 149.600 442.000 149.700 ;
        RECT 447.600 150.300 448.400 150.400 ;
        RECT 466.800 150.300 467.600 150.400 ;
        RECT 447.600 149.700 467.600 150.300 ;
        RECT 447.600 149.600 448.400 149.700 ;
        RECT 466.800 149.600 467.600 149.700 ;
        RECT 481.200 150.300 482.000 150.400 ;
        RECT 490.800 150.300 491.600 150.400 ;
        RECT 481.200 149.700 491.600 150.300 ;
        RECT 481.200 149.600 482.000 149.700 ;
        RECT 490.800 149.600 491.600 149.700 ;
        RECT 508.400 150.300 509.200 150.400 ;
        RECT 527.600 150.300 528.400 150.400 ;
        RECT 508.400 149.700 528.400 150.300 ;
        RECT 508.400 149.600 509.200 149.700 ;
        RECT 527.600 149.600 528.400 149.700 ;
        RECT 532.400 150.300 533.200 150.400 ;
        RECT 537.200 150.300 538.000 150.400 ;
        RECT 532.400 149.700 538.000 150.300 ;
        RECT 532.400 149.600 533.200 149.700 ;
        RECT 537.200 149.600 538.000 149.700 ;
        RECT 540.400 150.300 541.200 150.400 ;
        RECT 550.000 150.300 550.800 150.400 ;
        RECT 540.400 149.700 550.800 150.300 ;
        RECT 540.400 149.600 541.200 149.700 ;
        RECT 550.000 149.600 550.800 149.700 ;
        RECT 18.800 148.300 19.600 148.400 ;
        RECT 31.600 148.300 32.400 148.400 ;
        RECT 46.000 148.300 46.800 148.400 ;
        RECT 18.800 147.700 46.800 148.300 ;
        RECT 18.800 147.600 19.600 147.700 ;
        RECT 31.600 147.600 32.400 147.700 ;
        RECT 46.000 147.600 46.800 147.700 ;
        RECT 54.000 148.300 54.800 148.400 ;
        RECT 68.400 148.300 69.200 148.400 ;
        RECT 54.000 147.700 69.200 148.300 ;
        RECT 54.000 147.600 54.800 147.700 ;
        RECT 68.400 147.600 69.200 147.700 ;
        RECT 111.600 148.300 112.400 148.400 ;
        RECT 124.400 148.300 125.200 148.400 ;
        RECT 111.600 147.700 125.200 148.300 ;
        RECT 111.600 147.600 112.400 147.700 ;
        RECT 124.400 147.600 125.200 147.700 ;
        RECT 127.600 148.300 128.400 148.400 ;
        RECT 137.200 148.300 138.000 148.400 ;
        RECT 127.600 147.700 138.000 148.300 ;
        RECT 127.600 147.600 128.400 147.700 ;
        RECT 137.200 147.600 138.000 147.700 ;
        RECT 174.000 148.300 174.800 148.400 ;
        RECT 198.000 148.300 198.800 148.400 ;
        RECT 174.000 147.700 198.800 148.300 ;
        RECT 174.000 147.600 174.800 147.700 ;
        RECT 198.000 147.600 198.800 147.700 ;
        RECT 217.200 148.300 218.000 148.400 ;
        RECT 222.000 148.300 222.800 148.400 ;
        RECT 217.200 147.700 222.800 148.300 ;
        RECT 217.200 147.600 218.000 147.700 ;
        RECT 222.000 147.600 222.800 147.700 ;
        RECT 278.000 148.300 278.800 148.400 ;
        RECT 298.800 148.300 299.600 148.400 ;
        RECT 278.000 147.700 299.600 148.300 ;
        RECT 278.000 147.600 278.800 147.700 ;
        RECT 298.800 147.600 299.600 147.700 ;
        RECT 332.400 148.300 333.200 148.400 ;
        RECT 354.800 148.300 355.600 148.400 ;
        RECT 332.400 147.700 355.600 148.300 ;
        RECT 332.400 147.600 333.200 147.700 ;
        RECT 354.800 147.600 355.600 147.700 ;
        RECT 382.000 148.300 382.800 148.400 ;
        RECT 390.000 148.300 390.800 148.400 ;
        RECT 382.000 147.700 390.800 148.300 ;
        RECT 382.000 147.600 382.800 147.700 ;
        RECT 390.000 147.600 390.800 147.700 ;
        RECT 394.800 148.300 395.600 148.400 ;
        RECT 412.400 148.300 413.200 148.400 ;
        RECT 394.800 147.700 413.200 148.300 ;
        RECT 394.800 147.600 395.600 147.700 ;
        RECT 412.400 147.600 413.200 147.700 ;
        RECT 417.200 148.300 418.000 148.400 ;
        RECT 471.600 148.300 472.400 148.400 ;
        RECT 417.200 147.700 472.400 148.300 ;
        RECT 417.200 147.600 418.000 147.700 ;
        RECT 471.600 147.600 472.400 147.700 ;
        RECT 481.200 148.300 482.000 148.400 ;
        RECT 489.200 148.300 490.000 148.400 ;
        RECT 481.200 147.700 490.000 148.300 ;
        RECT 481.200 147.600 482.000 147.700 ;
        RECT 489.200 147.600 490.000 147.700 ;
        RECT 503.600 148.300 504.400 148.400 ;
        RECT 506.800 148.300 507.600 148.400 ;
        RECT 503.600 147.700 507.600 148.300 ;
        RECT 503.600 147.600 504.400 147.700 ;
        RECT 506.800 147.600 507.600 147.700 ;
        RECT 532.400 148.300 533.200 148.400 ;
        RECT 545.200 148.300 546.000 148.400 ;
        RECT 532.400 147.700 546.000 148.300 ;
        RECT 532.400 147.600 533.200 147.700 ;
        RECT 545.200 147.600 546.000 147.700 ;
        RECT 562.800 148.300 563.600 148.400 ;
        RECT 569.200 148.300 570.000 148.400 ;
        RECT 562.800 147.700 570.000 148.300 ;
        RECT 562.800 147.600 563.600 147.700 ;
        RECT 569.200 147.600 570.000 147.700 ;
        RECT 586.800 148.300 587.600 148.400 ;
        RECT 588.400 148.300 589.200 148.400 ;
        RECT 586.800 147.700 589.200 148.300 ;
        RECT 586.800 147.600 587.600 147.700 ;
        RECT 588.400 147.600 589.200 147.700 ;
        RECT 36.400 146.300 37.200 146.400 ;
        RECT 39.600 146.300 40.400 146.400 ;
        RECT 36.400 145.700 40.400 146.300 ;
        RECT 36.400 145.600 37.200 145.700 ;
        RECT 39.600 145.600 40.400 145.700 ;
        RECT 98.800 146.300 99.600 146.400 ;
        RECT 119.600 146.300 120.400 146.400 ;
        RECT 98.800 145.700 120.400 146.300 ;
        RECT 98.800 145.600 99.600 145.700 ;
        RECT 119.600 145.600 120.400 145.700 ;
        RECT 122.800 146.300 123.600 146.400 ;
        RECT 126.000 146.300 126.800 146.400 ;
        RECT 122.800 145.700 126.800 146.300 ;
        RECT 122.800 145.600 123.600 145.700 ;
        RECT 126.000 145.600 126.800 145.700 ;
        RECT 134.000 146.300 134.800 146.400 ;
        RECT 140.400 146.300 141.200 146.400 ;
        RECT 148.400 146.300 149.200 146.400 ;
        RECT 134.000 145.700 149.200 146.300 ;
        RECT 134.000 145.600 134.800 145.700 ;
        RECT 140.400 145.600 141.200 145.700 ;
        RECT 148.400 145.600 149.200 145.700 ;
        RECT 204.400 146.300 205.200 146.400 ;
        RECT 218.800 146.300 219.600 146.400 ;
        RECT 249.200 146.300 250.000 146.400 ;
        RECT 204.400 145.700 250.000 146.300 ;
        RECT 204.400 145.600 205.200 145.700 ;
        RECT 218.800 145.600 219.600 145.700 ;
        RECT 249.200 145.600 250.000 145.700 ;
        RECT 289.200 146.300 290.000 146.400 ;
        RECT 322.800 146.300 323.600 146.400 ;
        RECT 289.200 145.700 323.600 146.300 ;
        RECT 289.200 145.600 290.000 145.700 ;
        RECT 322.800 145.600 323.600 145.700 ;
        RECT 335.600 146.300 336.400 146.400 ;
        RECT 348.400 146.300 349.200 146.400 ;
        RECT 335.600 145.700 349.200 146.300 ;
        RECT 335.600 145.600 336.400 145.700 ;
        RECT 348.400 145.600 349.200 145.700 ;
        RECT 354.800 146.300 355.600 146.400 ;
        RECT 369.200 146.300 370.000 146.400 ;
        RECT 438.000 146.300 438.800 146.400 ;
        RECT 354.800 145.700 438.800 146.300 ;
        RECT 354.800 145.600 355.600 145.700 ;
        RECT 369.200 145.600 370.000 145.700 ;
        RECT 438.000 145.600 438.800 145.700 ;
        RECT 471.600 146.300 472.400 146.400 ;
        RECT 482.800 146.300 483.600 146.400 ;
        RECT 471.600 145.700 483.600 146.300 ;
        RECT 471.600 145.600 472.400 145.700 ;
        RECT 482.800 145.600 483.600 145.700 ;
        RECT 486.000 146.300 486.800 146.400 ;
        RECT 500.400 146.300 501.200 146.400 ;
        RECT 486.000 145.700 501.200 146.300 ;
        RECT 486.000 145.600 486.800 145.700 ;
        RECT 500.400 145.600 501.200 145.700 ;
        RECT 524.400 146.300 525.200 146.400 ;
        RECT 535.600 146.300 536.400 146.400 ;
        RECT 524.400 145.700 536.400 146.300 ;
        RECT 524.400 145.600 525.200 145.700 ;
        RECT 535.600 145.600 536.400 145.700 ;
        RECT 25.200 144.300 26.000 144.400 ;
        RECT 38.000 144.300 38.800 144.400 ;
        RECT 68.400 144.300 69.200 144.400 ;
        RECT 25.200 143.700 69.200 144.300 ;
        RECT 25.200 143.600 26.000 143.700 ;
        RECT 38.000 143.600 38.800 143.700 ;
        RECT 68.400 143.600 69.200 143.700 ;
        RECT 102.000 144.300 102.800 144.400 ;
        RECT 135.600 144.300 136.400 144.400 ;
        RECT 102.000 143.700 136.400 144.300 ;
        RECT 102.000 143.600 102.800 143.700 ;
        RECT 135.600 143.600 136.400 143.700 ;
        RECT 215.600 144.300 216.400 144.400 ;
        RECT 238.000 144.300 238.800 144.400 ;
        RECT 215.600 143.700 238.800 144.300 ;
        RECT 215.600 143.600 216.400 143.700 ;
        RECT 238.000 143.600 238.800 143.700 ;
        RECT 308.400 144.300 309.200 144.400 ;
        RECT 364.400 144.300 365.200 144.400 ;
        RECT 308.400 143.700 365.200 144.300 ;
        RECT 308.400 143.600 309.200 143.700 ;
        RECT 364.400 143.600 365.200 143.700 ;
        RECT 374.000 144.300 374.800 144.400 ;
        RECT 431.600 144.300 432.400 144.400 ;
        RECT 374.000 143.700 432.400 144.300 ;
        RECT 374.000 143.600 374.800 143.700 ;
        RECT 431.600 143.600 432.400 143.700 ;
        RECT 463.600 144.300 464.400 144.400 ;
        RECT 478.000 144.300 478.800 144.400 ;
        RECT 463.600 143.700 478.800 144.300 ;
        RECT 463.600 143.600 464.400 143.700 ;
        RECT 478.000 143.600 478.800 143.700 ;
        RECT 522.800 144.300 523.600 144.400 ;
        RECT 537.200 144.300 538.000 144.400 ;
        RECT 522.800 143.700 538.000 144.300 ;
        RECT 522.800 143.600 523.600 143.700 ;
        RECT 537.200 143.600 538.000 143.700 ;
        RECT 569.200 144.300 570.000 144.400 ;
        RECT 570.800 144.300 571.600 144.400 ;
        RECT 569.200 143.700 571.600 144.300 ;
        RECT 569.200 143.600 570.000 143.700 ;
        RECT 570.800 143.600 571.600 143.700 ;
        RECT 38.000 142.300 38.800 142.400 ;
        RECT 41.200 142.300 42.000 142.400 ;
        RECT 38.000 141.700 42.000 142.300 ;
        RECT 38.000 141.600 38.800 141.700 ;
        RECT 41.200 141.600 42.000 141.700 ;
        RECT 71.600 142.300 72.400 142.400 ;
        RECT 82.800 142.300 83.600 142.400 ;
        RECT 71.600 141.700 83.600 142.300 ;
        RECT 71.600 141.600 72.400 141.700 ;
        RECT 82.800 141.600 83.600 141.700 ;
        RECT 177.200 142.300 178.000 142.400 ;
        RECT 180.400 142.300 181.200 142.400 ;
        RECT 177.200 141.700 181.200 142.300 ;
        RECT 177.200 141.600 178.000 141.700 ;
        RECT 180.400 141.600 181.200 141.700 ;
        RECT 380.400 142.300 381.200 142.400 ;
        RECT 497.200 142.300 498.000 142.400 ;
        RECT 380.400 141.700 498.000 142.300 ;
        RECT 380.400 141.600 381.200 141.700 ;
        RECT 497.200 141.600 498.000 141.700 ;
        RECT 535.600 142.300 536.400 142.400 ;
        RECT 578.800 142.300 579.600 142.400 ;
        RECT 535.600 141.700 579.600 142.300 ;
        RECT 535.600 141.600 536.400 141.700 ;
        RECT 578.800 141.600 579.600 141.700 ;
        RECT 585.200 142.300 586.000 142.400 ;
        RECT 586.800 142.300 587.600 142.400 ;
        RECT 591.600 142.300 592.400 142.400 ;
        RECT 585.200 141.700 592.400 142.300 ;
        RECT 585.200 141.600 586.000 141.700 ;
        RECT 586.800 141.600 587.600 141.700 ;
        RECT 591.600 141.600 592.400 141.700 ;
        RECT 46.000 140.300 46.800 140.400 ;
        RECT 129.200 140.300 130.000 140.400 ;
        RECT 46.000 139.700 130.000 140.300 ;
        RECT 46.000 139.600 46.800 139.700 ;
        RECT 129.200 139.600 130.000 139.700 ;
        RECT 138.800 140.300 139.600 140.400 ;
        RECT 143.600 140.300 144.400 140.400 ;
        RECT 138.800 139.700 144.400 140.300 ;
        RECT 138.800 139.600 139.600 139.700 ;
        RECT 143.600 139.600 144.400 139.700 ;
        RECT 185.200 140.300 186.000 140.400 ;
        RECT 193.200 140.300 194.000 140.400 ;
        RECT 185.200 139.700 194.000 140.300 ;
        RECT 185.200 139.600 186.000 139.700 ;
        RECT 193.200 139.600 194.000 139.700 ;
        RECT 281.200 140.300 282.000 140.400 ;
        RECT 281.200 139.700 293.100 140.300 ;
        RECT 281.200 139.600 282.000 139.700 ;
        RECT 78.000 138.300 78.800 138.400 ;
        RECT 86.000 138.300 86.800 138.400 ;
        RECT 78.000 137.700 86.800 138.300 ;
        RECT 78.000 137.600 78.800 137.700 ;
        RECT 86.000 137.600 86.800 137.700 ;
        RECT 95.600 138.300 96.400 138.400 ;
        RECT 156.400 138.300 157.200 138.400 ;
        RECT 95.600 137.700 157.200 138.300 ;
        RECT 292.500 138.300 293.100 139.700 ;
        RECT 369.200 139.600 370.000 140.400 ;
        RECT 393.200 140.300 394.000 140.400 ;
        RECT 412.400 140.300 413.200 140.400 ;
        RECT 393.200 139.700 413.200 140.300 ;
        RECT 393.200 139.600 394.000 139.700 ;
        RECT 412.400 139.600 413.200 139.700 ;
        RECT 439.600 140.300 440.400 140.400 ;
        RECT 502.000 140.300 502.800 140.400 ;
        RECT 559.600 140.300 560.400 140.400 ;
        RECT 439.600 139.700 481.900 140.300 ;
        RECT 439.600 139.600 440.400 139.700 ;
        RECT 481.300 138.400 481.900 139.700 ;
        RECT 502.000 139.700 560.400 140.300 ;
        RECT 502.000 139.600 502.800 139.700 ;
        RECT 559.600 139.600 560.400 139.700 ;
        RECT 602.800 140.300 603.600 140.400 ;
        RECT 609.200 140.300 610.000 140.400 ;
        RECT 602.800 139.700 610.000 140.300 ;
        RECT 602.800 139.600 603.600 139.700 ;
        RECT 609.200 139.600 610.000 139.700 ;
        RECT 337.200 138.300 338.000 138.400 ;
        RECT 292.500 137.700 338.000 138.300 ;
        RECT 95.600 137.600 96.400 137.700 ;
        RECT 156.400 137.600 157.200 137.700 ;
        RECT 337.200 137.600 338.000 137.700 ;
        RECT 362.800 138.300 363.600 138.400 ;
        RECT 369.200 138.300 370.000 138.400 ;
        RECT 362.800 137.700 370.000 138.300 ;
        RECT 362.800 137.600 363.600 137.700 ;
        RECT 369.200 137.600 370.000 137.700 ;
        RECT 410.800 138.300 411.600 138.400 ;
        RECT 431.600 138.300 432.400 138.400 ;
        RECT 463.600 138.300 464.400 138.400 ;
        RECT 410.800 137.700 464.400 138.300 ;
        RECT 410.800 137.600 411.600 137.700 ;
        RECT 431.600 137.600 432.400 137.700 ;
        RECT 463.600 137.600 464.400 137.700 ;
        RECT 473.200 138.300 474.000 138.400 ;
        RECT 479.600 138.300 480.400 138.400 ;
        RECT 473.200 137.700 480.400 138.300 ;
        RECT 473.200 137.600 474.000 137.700 ;
        RECT 479.600 137.600 480.400 137.700 ;
        RECT 481.200 138.300 482.000 138.400 ;
        RECT 502.000 138.300 502.800 138.400 ;
        RECT 518.000 138.300 518.800 138.400 ;
        RECT 481.200 137.700 518.800 138.300 ;
        RECT 481.200 137.600 482.000 137.700 ;
        RECT 502.000 137.600 502.800 137.700 ;
        RECT 518.000 137.600 518.800 137.700 ;
        RECT 548.400 138.300 549.200 138.400 ;
        RECT 585.200 138.300 586.000 138.400 ;
        RECT 548.400 137.700 586.000 138.300 ;
        RECT 548.400 137.600 549.200 137.700 ;
        RECT 585.200 137.600 586.000 137.700 ;
        RECT 6.000 136.300 6.800 136.400 ;
        RECT 18.800 136.300 19.600 136.400 ;
        RECT 6.000 135.700 19.600 136.300 ;
        RECT 6.000 135.600 6.800 135.700 ;
        RECT 18.800 135.600 19.600 135.700 ;
        RECT 22.000 136.300 22.800 136.400 ;
        RECT 41.200 136.300 42.000 136.400 ;
        RECT 22.000 135.700 42.000 136.300 ;
        RECT 22.000 135.600 22.800 135.700 ;
        RECT 41.200 135.600 42.000 135.700 ;
        RECT 68.400 136.300 69.200 136.400 ;
        RECT 81.200 136.300 82.000 136.400 ;
        RECT 89.200 136.300 90.000 136.400 ;
        RECT 68.400 135.700 90.000 136.300 ;
        RECT 68.400 135.600 69.200 135.700 ;
        RECT 81.200 135.600 82.000 135.700 ;
        RECT 89.200 135.600 90.000 135.700 ;
        RECT 138.800 136.300 139.600 136.400 ;
        RECT 158.000 136.300 158.800 136.400 ;
        RECT 138.800 135.700 158.800 136.300 ;
        RECT 138.800 135.600 139.600 135.700 ;
        RECT 158.000 135.600 158.800 135.700 ;
        RECT 190.000 136.300 190.800 136.400 ;
        RECT 207.600 136.300 208.400 136.400 ;
        RECT 254.000 136.300 254.800 136.400 ;
        RECT 190.000 135.700 254.800 136.300 ;
        RECT 190.000 135.600 190.800 135.700 ;
        RECT 207.600 135.600 208.400 135.700 ;
        RECT 254.000 135.600 254.800 135.700 ;
        RECT 359.600 136.300 360.400 136.400 ;
        RECT 382.000 136.300 382.800 136.400 ;
        RECT 359.600 135.700 382.800 136.300 ;
        RECT 359.600 135.600 360.400 135.700 ;
        RECT 382.000 135.600 382.800 135.700 ;
        RECT 394.800 136.300 395.600 136.400 ;
        RECT 414.000 136.300 414.800 136.400 ;
        RECT 394.800 135.700 414.800 136.300 ;
        RECT 394.800 135.600 395.600 135.700 ;
        RECT 414.000 135.600 414.800 135.700 ;
        RECT 441.200 136.300 442.000 136.400 ;
        RECT 473.200 136.300 474.000 136.400 ;
        RECT 503.600 136.300 504.400 136.400 ;
        RECT 441.200 135.700 504.400 136.300 ;
        RECT 441.200 135.600 442.000 135.700 ;
        RECT 473.200 135.600 474.000 135.700 ;
        RECT 503.600 135.600 504.400 135.700 ;
        RECT 506.800 136.300 507.600 136.400 ;
        RECT 513.200 136.300 514.000 136.400 ;
        RECT 506.800 135.700 514.000 136.300 ;
        RECT 506.800 135.600 507.600 135.700 ;
        RECT 513.200 135.600 514.000 135.700 ;
        RECT 514.800 136.300 515.600 136.400 ;
        RECT 545.200 136.300 546.000 136.400 ;
        RECT 556.400 136.300 557.200 136.400 ;
        RECT 558.000 136.300 558.800 136.400 ;
        RECT 562.800 136.300 563.600 136.400 ;
        RECT 514.800 135.700 563.600 136.300 ;
        RECT 514.800 135.600 515.600 135.700 ;
        RECT 545.200 135.600 546.000 135.700 ;
        RECT 556.400 135.600 557.200 135.700 ;
        RECT 558.000 135.600 558.800 135.700 ;
        RECT 562.800 135.600 563.600 135.700 ;
        RECT 36.400 134.300 37.200 134.400 ;
        RECT 46.000 134.300 46.800 134.400 ;
        RECT 57.200 134.300 58.000 134.400 ;
        RECT 36.400 133.700 58.000 134.300 ;
        RECT 36.400 133.600 37.200 133.700 ;
        RECT 46.000 133.600 46.800 133.700 ;
        RECT 57.200 133.600 58.000 133.700 ;
        RECT 76.400 134.300 77.200 134.400 ;
        RECT 103.600 134.300 104.400 134.400 ;
        RECT 76.400 133.700 104.400 134.300 ;
        RECT 76.400 133.600 77.200 133.700 ;
        RECT 103.600 133.600 104.400 133.700 ;
        RECT 127.600 134.300 128.400 134.400 ;
        RECT 134.000 134.300 134.800 134.400 ;
        RECT 127.600 133.700 134.800 134.300 ;
        RECT 127.600 133.600 128.400 133.700 ;
        RECT 134.000 133.600 134.800 133.700 ;
        RECT 142.000 134.300 142.800 134.400 ;
        RECT 150.000 134.300 150.800 134.400 ;
        RECT 142.000 133.700 150.800 134.300 ;
        RECT 142.000 133.600 142.800 133.700 ;
        RECT 150.000 133.600 150.800 133.700 ;
        RECT 183.600 133.600 184.400 134.400 ;
        RECT 196.400 134.300 197.200 134.400 ;
        RECT 201.200 134.300 202.000 134.400 ;
        RECT 196.400 133.700 202.000 134.300 ;
        RECT 196.400 133.600 197.200 133.700 ;
        RECT 201.200 133.600 202.000 133.700 ;
        RECT 202.800 134.300 203.600 134.400 ;
        RECT 218.800 134.300 219.600 134.400 ;
        RECT 202.800 133.700 219.600 134.300 ;
        RECT 202.800 133.600 203.600 133.700 ;
        RECT 218.800 133.600 219.600 133.700 ;
        RECT 230.000 134.300 230.800 134.400 ;
        RECT 244.400 134.300 245.200 134.400 ;
        RECT 230.000 133.700 245.200 134.300 ;
        RECT 230.000 133.600 230.800 133.700 ;
        RECT 244.400 133.600 245.200 133.700 ;
        RECT 249.200 134.300 250.000 134.400 ;
        RECT 260.400 134.300 261.200 134.400 ;
        RECT 249.200 133.700 261.200 134.300 ;
        RECT 249.200 133.600 250.000 133.700 ;
        RECT 260.400 133.600 261.200 133.700 ;
        RECT 262.000 134.300 262.800 134.400 ;
        RECT 287.600 134.300 288.400 134.400 ;
        RECT 262.000 133.700 288.400 134.300 ;
        RECT 262.000 133.600 262.800 133.700 ;
        RECT 287.600 133.600 288.400 133.700 ;
        RECT 297.200 134.300 298.000 134.400 ;
        RECT 334.000 134.300 334.800 134.400 ;
        RECT 297.200 133.700 334.800 134.300 ;
        RECT 297.200 133.600 298.000 133.700 ;
        RECT 334.000 133.600 334.800 133.700 ;
        RECT 362.800 134.300 363.600 134.400 ;
        RECT 364.400 134.300 365.200 134.400 ;
        RECT 367.600 134.300 368.400 134.400 ;
        RECT 362.800 133.700 368.400 134.300 ;
        RECT 362.800 133.600 363.600 133.700 ;
        RECT 364.400 133.600 365.200 133.700 ;
        RECT 367.600 133.600 368.400 133.700 ;
        RECT 377.200 134.300 378.000 134.400 ;
        RECT 391.600 134.300 392.400 134.400 ;
        RECT 377.200 133.700 392.400 134.300 ;
        RECT 377.200 133.600 378.000 133.700 ;
        RECT 391.600 133.600 392.400 133.700 ;
        RECT 409.200 134.300 410.000 134.400 ;
        RECT 433.200 134.300 434.000 134.400 ;
        RECT 438.000 134.300 438.800 134.400 ;
        RECT 452.400 134.300 453.200 134.400 ;
        RECT 476.400 134.300 477.200 134.400 ;
        RECT 409.200 133.700 477.200 134.300 ;
        RECT 409.200 133.600 410.000 133.700 ;
        RECT 433.200 133.600 434.000 133.700 ;
        RECT 438.000 133.600 438.800 133.700 ;
        RECT 452.400 133.600 453.200 133.700 ;
        RECT 476.400 133.600 477.200 133.700 ;
        RECT 478.000 134.300 478.800 134.400 ;
        RECT 482.800 134.300 483.600 134.400 ;
        RECT 478.000 133.700 483.600 134.300 ;
        RECT 478.000 133.600 478.800 133.700 ;
        RECT 482.800 133.600 483.600 133.700 ;
        RECT 484.400 134.300 485.200 134.400 ;
        RECT 489.200 134.300 490.000 134.400 ;
        RECT 484.400 133.700 490.000 134.300 ;
        RECT 484.400 133.600 485.200 133.700 ;
        RECT 489.200 133.600 490.000 133.700 ;
        RECT 508.400 134.300 509.200 134.400 ;
        RECT 511.600 134.300 512.400 134.400 ;
        RECT 538.800 134.300 539.600 134.400 ;
        RECT 543.600 134.300 544.400 134.400 ;
        RECT 588.400 134.300 589.200 134.400 ;
        RECT 602.800 134.300 603.600 134.400 ;
        RECT 508.400 133.700 603.600 134.300 ;
        RECT 508.400 133.600 509.200 133.700 ;
        RECT 511.600 133.600 512.400 133.700 ;
        RECT 538.800 133.600 539.600 133.700 ;
        RECT 543.600 133.600 544.400 133.700 ;
        RECT 588.400 133.600 589.200 133.700 ;
        RECT 602.800 133.600 603.600 133.700 ;
        RECT 33.200 132.300 34.000 132.400 ;
        RECT 44.400 132.300 45.200 132.400 ;
        RECT 33.200 131.700 45.200 132.300 ;
        RECT 33.200 131.600 34.000 131.700 ;
        RECT 44.400 131.600 45.200 131.700 ;
        RECT 47.600 132.300 48.400 132.400 ;
        RECT 55.600 132.300 56.400 132.400 ;
        RECT 47.600 131.700 56.400 132.300 ;
        RECT 47.600 131.600 48.400 131.700 ;
        RECT 55.600 131.600 56.400 131.700 ;
        RECT 65.200 132.300 66.000 132.400 ;
        RECT 74.800 132.300 75.600 132.400 ;
        RECT 65.200 131.700 75.600 132.300 ;
        RECT 65.200 131.600 66.000 131.700 ;
        RECT 74.800 131.600 75.600 131.700 ;
        RECT 94.000 131.600 94.800 132.400 ;
        RECT 97.200 132.300 98.000 132.400 ;
        RECT 100.400 132.300 101.200 132.400 ;
        RECT 97.200 131.700 101.200 132.300 ;
        RECT 97.200 131.600 98.000 131.700 ;
        RECT 100.400 131.600 101.200 131.700 ;
        RECT 110.000 132.300 110.800 132.400 ;
        RECT 124.400 132.300 125.200 132.400 ;
        RECT 135.600 132.300 136.400 132.400 ;
        RECT 142.000 132.300 142.800 132.400 ;
        RECT 145.200 132.300 146.000 132.400 ;
        RECT 110.000 131.700 146.000 132.300 ;
        RECT 110.000 131.600 110.800 131.700 ;
        RECT 124.400 131.600 125.200 131.700 ;
        RECT 135.600 131.600 136.400 131.700 ;
        RECT 142.000 131.600 142.800 131.700 ;
        RECT 145.200 131.600 146.000 131.700 ;
        RECT 156.400 132.300 157.200 132.400 ;
        RECT 183.700 132.300 184.300 133.600 ;
        RECT 156.400 131.700 184.300 132.300 ;
        RECT 193.200 132.300 194.000 132.400 ;
        RECT 202.800 132.300 203.600 132.400 ;
        RECT 193.200 131.700 203.600 132.300 ;
        RECT 156.400 131.600 157.200 131.700 ;
        RECT 193.200 131.600 194.000 131.700 ;
        RECT 202.800 131.600 203.600 131.700 ;
        RECT 206.000 132.300 206.800 132.400 ;
        RECT 209.200 132.300 210.000 132.400 ;
        RECT 206.000 131.700 210.000 132.300 ;
        RECT 206.000 131.600 206.800 131.700 ;
        RECT 209.200 131.600 210.000 131.700 ;
        RECT 252.400 132.300 253.200 132.400 ;
        RECT 262.000 132.300 262.800 132.400 ;
        RECT 252.400 131.700 262.800 132.300 ;
        RECT 252.400 131.600 253.200 131.700 ;
        RECT 262.000 131.600 262.800 131.700 ;
        RECT 284.400 132.300 285.200 132.400 ;
        RECT 306.800 132.300 307.600 132.400 ;
        RECT 284.400 131.700 307.600 132.300 ;
        RECT 284.400 131.600 285.200 131.700 ;
        RECT 306.800 131.600 307.600 131.700 ;
        RECT 334.000 132.300 334.800 132.400 ;
        RECT 353.200 132.300 354.000 132.400 ;
        RECT 366.000 132.300 366.800 132.400 ;
        RECT 334.000 131.700 366.800 132.300 ;
        RECT 334.000 131.600 334.800 131.700 ;
        RECT 353.200 131.600 354.000 131.700 ;
        RECT 366.000 131.600 366.800 131.700 ;
        RECT 406.000 132.300 406.800 132.400 ;
        RECT 444.400 132.300 445.200 132.400 ;
        RECT 449.200 132.300 450.000 132.400 ;
        RECT 406.000 131.700 450.000 132.300 ;
        RECT 406.000 131.600 406.800 131.700 ;
        RECT 444.400 131.600 445.200 131.700 ;
        RECT 449.200 131.600 450.000 131.700 ;
        RECT 450.800 132.300 451.600 132.400 ;
        RECT 494.000 132.300 494.800 132.400 ;
        RECT 450.800 131.700 494.800 132.300 ;
        RECT 450.800 131.600 451.600 131.700 ;
        RECT 494.000 131.600 494.800 131.700 ;
        RECT 510.000 132.300 510.800 132.400 ;
        RECT 540.400 132.300 541.200 132.400 ;
        RECT 510.000 131.700 541.200 132.300 ;
        RECT 510.000 131.600 510.800 131.700 ;
        RECT 540.400 131.600 541.200 131.700 ;
        RECT 551.600 132.300 552.400 132.400 ;
        RECT 564.400 132.300 565.200 132.400 ;
        RECT 551.600 131.700 565.200 132.300 ;
        RECT 551.600 131.600 552.400 131.700 ;
        RECT 564.400 131.600 565.200 131.700 ;
        RECT 567.600 132.300 568.400 132.400 ;
        RECT 583.600 132.300 584.400 132.400 ;
        RECT 567.600 131.700 584.400 132.300 ;
        RECT 567.600 131.600 568.400 131.700 ;
        RECT 583.600 131.600 584.400 131.700 ;
        RECT 585.200 132.300 586.000 132.400 ;
        RECT 594.800 132.300 595.600 132.400 ;
        RECT 585.200 131.700 595.600 132.300 ;
        RECT 585.200 131.600 586.000 131.700 ;
        RECT 594.800 131.600 595.600 131.700 ;
        RECT 2.800 130.300 3.600 130.400 ;
        RECT 14.000 130.300 14.800 130.400 ;
        RECT 39.600 130.300 40.400 130.400 ;
        RECT 2.800 129.700 40.400 130.300 ;
        RECT 2.800 129.600 3.600 129.700 ;
        RECT 14.000 129.600 14.800 129.700 ;
        RECT 39.600 129.600 40.400 129.700 ;
        RECT 57.200 130.300 58.000 130.400 ;
        RECT 106.800 130.300 107.600 130.400 ;
        RECT 57.200 129.700 107.600 130.300 ;
        RECT 57.200 129.600 58.000 129.700 ;
        RECT 106.800 129.600 107.600 129.700 ;
        RECT 113.200 130.300 114.000 130.400 ;
        RECT 124.400 130.300 125.200 130.400 ;
        RECT 132.400 130.300 133.200 130.400 ;
        RECT 113.200 129.700 133.200 130.300 ;
        RECT 113.200 129.600 114.000 129.700 ;
        RECT 124.400 129.600 125.200 129.700 ;
        RECT 132.400 129.600 133.200 129.700 ;
        RECT 134.000 130.300 134.800 130.400 ;
        RECT 146.800 130.300 147.600 130.400 ;
        RECT 134.000 129.700 147.600 130.300 ;
        RECT 134.000 129.600 134.800 129.700 ;
        RECT 146.800 129.600 147.600 129.700 ;
        RECT 158.000 130.300 158.800 130.400 ;
        RECT 209.200 130.300 210.000 130.400 ;
        RECT 158.000 129.700 210.000 130.300 ;
        RECT 158.000 129.600 158.800 129.700 ;
        RECT 209.200 129.600 210.000 129.700 ;
        RECT 257.200 130.300 258.000 130.400 ;
        RECT 276.400 130.300 277.200 130.400 ;
        RECT 257.200 129.700 277.200 130.300 ;
        RECT 257.200 129.600 258.000 129.700 ;
        RECT 276.400 129.600 277.200 129.700 ;
        RECT 404.400 130.300 405.200 130.400 ;
        RECT 433.200 130.300 434.000 130.400 ;
        RECT 452.400 130.300 453.200 130.400 ;
        RECT 404.400 129.700 453.200 130.300 ;
        RECT 404.400 129.600 405.200 129.700 ;
        RECT 433.200 129.600 434.000 129.700 ;
        RECT 452.400 129.600 453.200 129.700 ;
        RECT 484.400 130.300 485.200 130.400 ;
        RECT 487.600 130.300 488.400 130.400 ;
        RECT 484.400 129.700 488.400 130.300 ;
        RECT 484.400 129.600 485.200 129.700 ;
        RECT 487.600 129.600 488.400 129.700 ;
        RECT 492.400 130.300 493.200 130.400 ;
        RECT 529.200 130.300 530.000 130.400 ;
        RECT 492.400 129.700 530.000 130.300 ;
        RECT 492.400 129.600 493.200 129.700 ;
        RECT 529.200 129.600 530.000 129.700 ;
        RECT 553.200 130.300 554.000 130.400 ;
        RECT 556.400 130.300 557.200 130.400 ;
        RECT 553.200 129.700 557.200 130.300 ;
        RECT 553.200 129.600 554.000 129.700 ;
        RECT 556.400 129.600 557.200 129.700 ;
        RECT 561.200 130.300 562.000 130.400 ;
        RECT 567.600 130.300 568.400 130.400 ;
        RECT 570.800 130.300 571.600 130.400 ;
        RECT 607.600 130.300 608.400 130.400 ;
        RECT 561.200 129.700 608.400 130.300 ;
        RECT 561.200 129.600 562.000 129.700 ;
        RECT 567.600 129.600 568.400 129.700 ;
        RECT 570.800 129.600 571.600 129.700 ;
        RECT 607.600 129.600 608.400 129.700 ;
        RECT 42.800 128.300 43.600 128.400 ;
        RECT 66.800 128.300 67.600 128.400 ;
        RECT 42.800 127.700 67.600 128.300 ;
        RECT 42.800 127.600 43.600 127.700 ;
        RECT 66.800 127.600 67.600 127.700 ;
        RECT 130.800 128.300 131.600 128.400 ;
        RECT 138.800 128.300 139.600 128.400 ;
        RECT 130.800 127.700 139.600 128.300 ;
        RECT 130.800 127.600 131.600 127.700 ;
        RECT 138.800 127.600 139.600 127.700 ;
        RECT 154.800 128.300 155.600 128.400 ;
        RECT 161.200 128.300 162.000 128.400 ;
        RECT 238.000 128.300 238.800 128.400 ;
        RECT 154.800 127.700 238.800 128.300 ;
        RECT 154.800 127.600 155.600 127.700 ;
        RECT 161.200 127.600 162.000 127.700 ;
        RECT 238.000 127.600 238.800 127.700 ;
        RECT 372.400 128.300 373.200 128.400 ;
        RECT 374.000 128.300 374.800 128.400 ;
        RECT 410.800 128.300 411.600 128.400 ;
        RECT 372.400 127.700 411.600 128.300 ;
        RECT 372.400 127.600 373.200 127.700 ;
        RECT 374.000 127.600 374.800 127.700 ;
        RECT 410.800 127.600 411.600 127.700 ;
        RECT 433.200 128.300 434.000 128.400 ;
        RECT 450.800 128.300 451.600 128.400 ;
        RECT 474.800 128.300 475.600 128.400 ;
        RECT 433.200 127.700 451.600 128.300 ;
        RECT 433.200 127.600 434.000 127.700 ;
        RECT 450.800 127.600 451.600 127.700 ;
        RECT 466.900 127.700 475.600 128.300 ;
        RECT 487.700 128.300 488.300 129.600 ;
        RECT 519.600 128.300 520.400 128.400 ;
        RECT 546.800 128.300 547.600 128.400 ;
        RECT 487.700 127.700 547.600 128.300 ;
        RECT 54.000 126.300 54.800 126.400 ;
        RECT 121.200 126.300 122.000 126.400 ;
        RECT 54.000 125.700 122.000 126.300 ;
        RECT 54.000 125.600 54.800 125.700 ;
        RECT 121.200 125.600 122.000 125.700 ;
        RECT 135.600 126.300 136.400 126.400 ;
        RECT 154.900 126.300 155.500 127.600 ;
        RECT 135.600 125.700 155.500 126.300 ;
        RECT 426.800 126.300 427.600 126.400 ;
        RECT 447.600 126.300 448.400 126.400 ;
        RECT 466.900 126.300 467.500 127.700 ;
        RECT 474.800 127.600 475.600 127.700 ;
        RECT 519.600 127.600 520.400 127.700 ;
        RECT 546.800 127.600 547.600 127.700 ;
        RECT 426.800 125.700 467.500 126.300 ;
        RECT 468.400 126.300 469.200 126.400 ;
        RECT 506.800 126.300 507.600 126.400 ;
        RECT 468.400 125.700 507.600 126.300 ;
        RECT 135.600 125.600 136.400 125.700 ;
        RECT 426.800 125.600 427.600 125.700 ;
        RECT 447.600 125.600 448.400 125.700 ;
        RECT 468.400 125.600 469.200 125.700 ;
        RECT 506.800 125.600 507.600 125.700 ;
        RECT 41.200 124.300 42.000 124.400 ;
        RECT 42.800 124.300 43.600 124.400 ;
        RECT 41.200 123.700 43.600 124.300 ;
        RECT 41.200 123.600 42.000 123.700 ;
        RECT 42.800 123.600 43.600 123.700 ;
        RECT 46.000 124.300 46.800 124.400 ;
        RECT 62.000 124.300 62.800 124.400 ;
        RECT 46.000 123.700 62.800 124.300 ;
        RECT 46.000 123.600 46.800 123.700 ;
        RECT 62.000 123.600 62.800 123.700 ;
        RECT 68.400 124.300 69.200 124.400 ;
        RECT 119.600 124.300 120.400 124.400 ;
        RECT 126.000 124.300 126.800 124.400 ;
        RECT 68.400 123.700 126.800 124.300 ;
        RECT 68.400 123.600 69.200 123.700 ;
        RECT 119.600 123.600 120.400 123.700 ;
        RECT 126.000 123.600 126.800 123.700 ;
        RECT 146.800 124.300 147.600 124.400 ;
        RECT 150.000 124.300 150.800 124.400 ;
        RECT 146.800 123.700 150.800 124.300 ;
        RECT 146.800 123.600 147.600 123.700 ;
        RECT 150.000 123.600 150.800 123.700 ;
        RECT 153.200 124.300 154.000 124.400 ;
        RECT 158.000 124.300 158.800 124.400 ;
        RECT 153.200 123.700 158.800 124.300 ;
        RECT 153.200 123.600 154.000 123.700 ;
        RECT 158.000 123.600 158.800 123.700 ;
        RECT 345.200 124.300 346.000 124.400 ;
        RECT 394.800 124.300 395.600 124.400 ;
        RECT 510.000 124.300 510.800 124.400 ;
        RECT 345.200 123.700 510.800 124.300 ;
        RECT 345.200 123.600 346.000 123.700 ;
        RECT 394.800 123.600 395.600 123.700 ;
        RECT 510.000 123.600 510.800 123.700 ;
        RECT 522.800 124.300 523.600 124.400 ;
        RECT 569.200 124.300 570.000 124.400 ;
        RECT 522.800 123.700 570.000 124.300 ;
        RECT 522.800 123.600 523.600 123.700 ;
        RECT 569.200 123.600 570.000 123.700 ;
        RECT 62.100 122.300 62.700 123.600 ;
        RECT 84.400 122.300 85.200 122.400 ;
        RECT 87.600 122.300 88.400 122.400 ;
        RECT 62.100 121.700 88.400 122.300 ;
        RECT 84.400 121.600 85.200 121.700 ;
        RECT 87.600 121.600 88.400 121.700 ;
        RECT 98.800 122.300 99.600 122.400 ;
        RECT 100.400 122.300 101.200 122.400 ;
        RECT 98.800 121.700 101.200 122.300 ;
        RECT 98.800 121.600 99.600 121.700 ;
        RECT 100.400 121.600 101.200 121.700 ;
        RECT 103.600 122.300 104.400 122.400 ;
        RECT 142.000 122.300 142.800 122.400 ;
        RECT 103.600 121.700 142.800 122.300 ;
        RECT 103.600 121.600 104.400 121.700 ;
        RECT 142.000 121.600 142.800 121.700 ;
        RECT 228.400 122.300 229.200 122.400 ;
        RECT 265.200 122.300 266.000 122.400 ;
        RECT 228.400 121.700 266.000 122.300 ;
        RECT 228.400 121.600 229.200 121.700 ;
        RECT 265.200 121.600 266.000 121.700 ;
        RECT 377.200 122.300 378.000 122.400 ;
        RECT 401.200 122.300 402.000 122.400 ;
        RECT 377.200 121.700 402.000 122.300 ;
        RECT 377.200 121.600 378.000 121.700 ;
        RECT 401.200 121.600 402.000 121.700 ;
        RECT 406.000 122.300 406.800 122.400 ;
        RECT 428.400 122.300 429.200 122.400 ;
        RECT 436.400 122.300 437.200 122.400 ;
        RECT 406.000 121.700 437.200 122.300 ;
        RECT 406.000 121.600 406.800 121.700 ;
        RECT 428.400 121.600 429.200 121.700 ;
        RECT 436.400 121.600 437.200 121.700 ;
        RECT 481.200 122.300 482.000 122.400 ;
        RECT 503.600 122.300 504.400 122.400 ;
        RECT 481.200 121.700 504.400 122.300 ;
        RECT 481.200 121.600 482.000 121.700 ;
        RECT 503.600 121.600 504.400 121.700 ;
        RECT 506.800 122.300 507.600 122.400 ;
        RECT 510.000 122.300 510.800 122.400 ;
        RECT 506.800 121.700 510.800 122.300 ;
        RECT 506.800 121.600 507.600 121.700 ;
        RECT 510.000 121.600 510.800 121.700 ;
        RECT 170.800 120.300 171.600 120.400 ;
        RECT 180.400 120.300 181.200 120.400 ;
        RECT 170.800 119.700 181.200 120.300 ;
        RECT 170.800 119.600 171.600 119.700 ;
        RECT 180.400 119.600 181.200 119.700 ;
        RECT 223.600 120.300 224.400 120.400 ;
        RECT 247.600 120.300 248.400 120.400 ;
        RECT 223.600 119.700 248.400 120.300 ;
        RECT 223.600 119.600 224.400 119.700 ;
        RECT 247.600 119.600 248.400 119.700 ;
        RECT 257.200 120.300 258.000 120.400 ;
        RECT 266.800 120.300 267.600 120.400 ;
        RECT 257.200 119.700 267.600 120.300 ;
        RECT 257.200 119.600 258.000 119.700 ;
        RECT 266.800 119.600 267.600 119.700 ;
        RECT 330.800 120.300 331.600 120.400 ;
        RECT 337.200 120.300 338.000 120.400 ;
        RECT 330.800 119.700 338.000 120.300 ;
        RECT 330.800 119.600 331.600 119.700 ;
        RECT 337.200 119.600 338.000 119.700 ;
        RECT 425.200 120.300 426.000 120.400 ;
        RECT 446.000 120.300 446.800 120.400 ;
        RECT 425.200 119.700 446.800 120.300 ;
        RECT 425.200 119.600 426.000 119.700 ;
        RECT 446.000 119.600 446.800 119.700 ;
        RECT 487.600 120.300 488.400 120.400 ;
        RECT 505.200 120.300 506.000 120.400 ;
        RECT 487.600 119.700 506.000 120.300 ;
        RECT 487.600 119.600 488.400 119.700 ;
        RECT 505.200 119.600 506.000 119.700 ;
        RECT 583.600 120.300 584.400 120.400 ;
        RECT 596.400 120.300 597.200 120.400 ;
        RECT 583.600 119.700 597.200 120.300 ;
        RECT 583.600 119.600 584.400 119.700 ;
        RECT 596.400 119.600 597.200 119.700 ;
        RECT 193.200 118.300 194.000 118.400 ;
        RECT 226.800 118.300 227.600 118.400 ;
        RECT 193.200 117.700 227.600 118.300 ;
        RECT 193.200 117.600 194.000 117.700 ;
        RECT 226.800 117.600 227.600 117.700 ;
        RECT 249.200 118.300 250.000 118.400 ;
        RECT 262.000 118.300 262.800 118.400 ;
        RECT 282.800 118.300 283.600 118.400 ;
        RECT 249.200 117.700 283.600 118.300 ;
        RECT 249.200 117.600 250.000 117.700 ;
        RECT 262.000 117.600 262.800 117.700 ;
        RECT 282.800 117.600 283.600 117.700 ;
        RECT 422.000 118.300 422.800 118.400 ;
        RECT 442.800 118.300 443.600 118.400 ;
        RECT 422.000 117.700 443.600 118.300 ;
        RECT 422.000 117.600 422.800 117.700 ;
        RECT 442.800 117.600 443.600 117.700 ;
        RECT 449.200 118.300 450.000 118.400 ;
        RECT 489.200 118.300 490.000 118.400 ;
        RECT 495.600 118.300 496.400 118.400 ;
        RECT 542.000 118.300 542.800 118.400 ;
        RECT 449.200 117.700 542.800 118.300 ;
        RECT 449.200 117.600 450.000 117.700 ;
        RECT 489.200 117.600 490.000 117.700 ;
        RECT 495.600 117.600 496.400 117.700 ;
        RECT 542.000 117.600 542.800 117.700 ;
        RECT 585.200 118.300 586.000 118.400 ;
        RECT 590.000 118.300 590.800 118.400 ;
        RECT 602.800 118.300 603.600 118.400 ;
        RECT 585.200 117.700 603.600 118.300 ;
        RECT 585.200 117.600 586.000 117.700 ;
        RECT 590.000 117.600 590.800 117.700 ;
        RECT 602.800 117.600 603.600 117.700 ;
        RECT 23.600 116.300 24.400 116.400 ;
        RECT 50.800 116.300 51.600 116.400 ;
        RECT 23.600 115.700 51.600 116.300 ;
        RECT 23.600 115.600 24.400 115.700 ;
        RECT 50.800 115.600 51.600 115.700 ;
        RECT 87.600 116.300 88.400 116.400 ;
        RECT 113.200 116.300 114.000 116.400 ;
        RECT 87.600 115.700 114.000 116.300 ;
        RECT 87.600 115.600 88.400 115.700 ;
        RECT 113.200 115.600 114.000 115.700 ;
        RECT 118.000 116.300 118.800 116.400 ;
        RECT 193.200 116.300 194.000 116.400 ;
        RECT 198.000 116.300 198.800 116.400 ;
        RECT 118.000 115.700 198.800 116.300 ;
        RECT 118.000 115.600 118.800 115.700 ;
        RECT 193.200 115.600 194.000 115.700 ;
        RECT 198.000 115.600 198.800 115.700 ;
        RECT 238.000 116.300 238.800 116.400 ;
        RECT 250.800 116.300 251.600 116.400 ;
        RECT 238.000 115.700 251.600 116.300 ;
        RECT 238.000 115.600 238.800 115.700 ;
        RECT 250.800 115.600 251.600 115.700 ;
        RECT 366.000 116.300 366.800 116.400 ;
        RECT 369.200 116.300 370.000 116.400 ;
        RECT 366.000 115.700 370.000 116.300 ;
        RECT 366.000 115.600 366.800 115.700 ;
        RECT 369.200 115.600 370.000 115.700 ;
        RECT 428.400 116.300 429.200 116.400 ;
        RECT 431.600 116.300 432.400 116.400 ;
        RECT 428.400 115.700 432.400 116.300 ;
        RECT 428.400 115.600 429.200 115.700 ;
        RECT 431.600 115.600 432.400 115.700 ;
        RECT 444.400 116.300 445.200 116.400 ;
        RECT 450.800 116.300 451.600 116.400 ;
        RECT 444.400 115.700 451.600 116.300 ;
        RECT 444.400 115.600 445.200 115.700 ;
        RECT 450.800 115.600 451.600 115.700 ;
        RECT 503.600 116.300 504.400 116.400 ;
        RECT 567.600 116.300 568.400 116.400 ;
        RECT 503.600 115.700 568.400 116.300 ;
        RECT 503.600 115.600 504.400 115.700 ;
        RECT 567.600 115.600 568.400 115.700 ;
        RECT 18.800 114.300 19.600 114.400 ;
        RECT 26.800 114.300 27.600 114.400 ;
        RECT 54.000 114.300 54.800 114.400 ;
        RECT 18.800 113.700 54.800 114.300 ;
        RECT 18.800 113.600 19.600 113.700 ;
        RECT 26.800 113.600 27.600 113.700 ;
        RECT 54.000 113.600 54.800 113.700 ;
        RECT 86.000 114.300 86.800 114.400 ;
        RECT 95.600 114.300 96.400 114.400 ;
        RECT 86.000 113.700 96.400 114.300 ;
        RECT 86.000 113.600 86.800 113.700 ;
        RECT 95.600 113.600 96.400 113.700 ;
        RECT 106.800 114.300 107.600 114.400 ;
        RECT 119.600 114.300 120.400 114.400 ;
        RECT 135.600 114.300 136.400 114.400 ;
        RECT 106.800 113.700 136.400 114.300 ;
        RECT 106.800 113.600 107.600 113.700 ;
        RECT 119.600 113.600 120.400 113.700 ;
        RECT 135.600 113.600 136.400 113.700 ;
        RECT 220.400 114.300 221.200 114.400 ;
        RECT 223.600 114.300 224.400 114.400 ;
        RECT 220.400 113.700 224.400 114.300 ;
        RECT 220.400 113.600 221.200 113.700 ;
        RECT 223.600 113.600 224.400 113.700 ;
        RECT 226.800 114.300 227.600 114.400 ;
        RECT 260.400 114.300 261.200 114.400 ;
        RECT 226.800 113.700 261.200 114.300 ;
        RECT 226.800 113.600 227.600 113.700 ;
        RECT 260.400 113.600 261.200 113.700 ;
        RECT 276.400 114.300 277.200 114.400 ;
        RECT 286.000 114.300 286.800 114.400 ;
        RECT 290.800 114.300 291.600 114.400 ;
        RECT 276.400 113.700 291.600 114.300 ;
        RECT 276.400 113.600 277.200 113.700 ;
        RECT 286.000 113.600 286.800 113.700 ;
        RECT 290.800 113.600 291.600 113.700 ;
        RECT 369.200 113.600 370.000 114.400 ;
        RECT 430.000 114.300 430.800 114.400 ;
        RECT 441.200 114.300 442.000 114.400 ;
        RECT 430.000 113.700 442.000 114.300 ;
        RECT 430.000 113.600 430.800 113.700 ;
        RECT 441.200 113.600 442.000 113.700 ;
        RECT 446.000 114.300 446.800 114.400 ;
        RECT 471.600 114.300 472.400 114.400 ;
        RECT 446.000 113.700 472.400 114.300 ;
        RECT 446.000 113.600 446.800 113.700 ;
        RECT 471.600 113.600 472.400 113.700 ;
        RECT 503.600 114.300 504.400 114.400 ;
        RECT 522.800 114.300 523.600 114.400 ;
        RECT 503.600 113.700 523.600 114.300 ;
        RECT 503.600 113.600 504.400 113.700 ;
        RECT 522.800 113.600 523.600 113.700 ;
        RECT 534.000 114.300 534.800 114.400 ;
        RECT 550.000 114.300 550.800 114.400 ;
        RECT 534.000 113.700 550.800 114.300 ;
        RECT 534.000 113.600 534.800 113.700 ;
        RECT 550.000 113.600 550.800 113.700 ;
        RECT 30.000 112.300 30.800 112.400 ;
        RECT 50.800 112.300 51.600 112.400 ;
        RECT 58.800 112.300 59.600 112.400 ;
        RECT 73.200 112.300 74.000 112.400 ;
        RECT 30.000 111.700 74.000 112.300 ;
        RECT 30.000 111.600 30.800 111.700 ;
        RECT 50.800 111.600 51.600 111.700 ;
        RECT 58.800 111.600 59.600 111.700 ;
        RECT 73.200 111.600 74.000 111.700 ;
        RECT 82.800 112.300 83.600 112.400 ;
        RECT 94.000 112.300 94.800 112.400 ;
        RECT 121.200 112.300 122.000 112.400 ;
        RECT 122.800 112.300 123.600 112.400 ;
        RECT 82.800 111.700 123.600 112.300 ;
        RECT 82.800 111.600 83.600 111.700 ;
        RECT 94.000 111.600 94.800 111.700 ;
        RECT 121.200 111.600 122.000 111.700 ;
        RECT 122.800 111.600 123.600 111.700 ;
        RECT 132.400 112.300 133.200 112.400 ;
        RECT 142.000 112.300 142.800 112.400 ;
        RECT 150.000 112.300 150.800 112.400 ;
        RECT 164.400 112.300 165.200 112.400 ;
        RECT 132.400 111.700 165.200 112.300 ;
        RECT 132.400 111.600 133.200 111.700 ;
        RECT 142.000 111.600 142.800 111.700 ;
        RECT 150.000 111.600 150.800 111.700 ;
        RECT 164.400 111.600 165.200 111.700 ;
        RECT 214.000 112.300 214.800 112.400 ;
        RECT 218.800 112.300 219.600 112.400 ;
        RECT 214.000 111.700 219.600 112.300 ;
        RECT 214.000 111.600 214.800 111.700 ;
        RECT 218.800 111.600 219.600 111.700 ;
        RECT 250.800 112.300 251.600 112.400 ;
        RECT 257.200 112.300 258.000 112.400 ;
        RECT 250.800 111.700 258.000 112.300 ;
        RECT 250.800 111.600 251.600 111.700 ;
        RECT 257.200 111.600 258.000 111.700 ;
        RECT 422.000 112.300 422.800 112.400 ;
        RECT 439.600 112.300 440.400 112.400 ;
        RECT 422.000 111.700 440.400 112.300 ;
        RECT 422.000 111.600 422.800 111.700 ;
        RECT 439.600 111.600 440.400 111.700 ;
        RECT 444.400 112.300 445.200 112.400 ;
        RECT 446.000 112.300 446.800 112.400 ;
        RECT 510.000 112.300 510.800 112.400 ;
        RECT 444.400 111.700 446.800 112.300 ;
        RECT 444.400 111.600 445.200 111.700 ;
        RECT 446.000 111.600 446.800 111.700 ;
        RECT 447.700 111.700 510.800 112.300 ;
        RECT 9.200 110.300 10.000 110.400 ;
        RECT 22.000 110.300 22.800 110.400 ;
        RECT 9.200 109.700 22.800 110.300 ;
        RECT 9.200 109.600 10.000 109.700 ;
        RECT 22.000 109.600 22.800 109.700 ;
        RECT 54.000 110.300 54.800 110.400 ;
        RECT 68.400 110.300 69.200 110.400 ;
        RECT 54.000 109.700 69.200 110.300 ;
        RECT 54.000 109.600 54.800 109.700 ;
        RECT 68.400 109.600 69.200 109.700 ;
        RECT 98.800 110.300 99.600 110.400 ;
        RECT 110.000 110.300 110.800 110.400 ;
        RECT 98.800 109.700 110.800 110.300 ;
        RECT 98.800 109.600 99.600 109.700 ;
        RECT 110.000 109.600 110.800 109.700 ;
        RECT 142.000 110.300 142.800 110.400 ;
        RECT 153.200 110.300 154.000 110.400 ;
        RECT 142.000 109.700 154.000 110.300 ;
        RECT 142.000 109.600 142.800 109.700 ;
        RECT 153.200 109.600 154.000 109.700 ;
        RECT 175.600 110.300 176.400 110.400 ;
        RECT 185.200 110.300 186.000 110.400 ;
        RECT 198.000 110.300 198.800 110.400 ;
        RECT 175.600 109.700 198.800 110.300 ;
        RECT 175.600 109.600 176.400 109.700 ;
        RECT 185.200 109.600 186.000 109.700 ;
        RECT 198.000 109.600 198.800 109.700 ;
        RECT 202.800 110.300 203.600 110.400 ;
        RECT 218.800 110.300 219.600 110.400 ;
        RECT 222.000 110.300 222.800 110.400 ;
        RECT 225.200 110.300 226.000 110.400 ;
        RECT 202.800 109.700 226.000 110.300 ;
        RECT 202.800 109.600 203.600 109.700 ;
        RECT 218.800 109.600 219.600 109.700 ;
        RECT 222.000 109.600 222.800 109.700 ;
        RECT 225.200 109.600 226.000 109.700 ;
        RECT 233.200 110.300 234.000 110.400 ;
        RECT 236.400 110.300 237.200 110.400 ;
        RECT 244.400 110.300 245.200 110.400 ;
        RECT 233.200 109.700 245.200 110.300 ;
        RECT 233.200 109.600 234.000 109.700 ;
        RECT 236.400 109.600 237.200 109.700 ;
        RECT 244.400 109.600 245.200 109.700 ;
        RECT 260.400 110.300 261.200 110.400 ;
        RECT 284.400 110.300 285.200 110.400 ;
        RECT 260.400 109.700 285.200 110.300 ;
        RECT 260.400 109.600 261.200 109.700 ;
        RECT 284.400 109.600 285.200 109.700 ;
        RECT 343.600 110.300 344.400 110.400 ;
        RECT 350.000 110.300 350.800 110.400 ;
        RECT 343.600 109.700 350.800 110.300 ;
        RECT 343.600 109.600 344.400 109.700 ;
        RECT 350.000 109.600 350.800 109.700 ;
        RECT 386.800 110.300 387.600 110.400 ;
        RECT 415.600 110.300 416.400 110.400 ;
        RECT 386.800 109.700 416.400 110.300 ;
        RECT 386.800 109.600 387.600 109.700 ;
        RECT 415.600 109.600 416.400 109.700 ;
        RECT 418.800 110.300 419.600 110.400 ;
        RECT 428.400 110.300 429.200 110.400 ;
        RECT 418.800 109.700 429.200 110.300 ;
        RECT 418.800 109.600 419.600 109.700 ;
        RECT 428.400 109.600 429.200 109.700 ;
        RECT 441.200 110.300 442.000 110.400 ;
        RECT 447.700 110.300 448.300 111.700 ;
        RECT 510.000 111.600 510.800 111.700 ;
        RECT 521.200 112.300 522.000 112.400 ;
        RECT 530.800 112.300 531.600 112.400 ;
        RECT 537.200 112.300 538.000 112.400 ;
        RECT 521.200 111.700 538.000 112.300 ;
        RECT 521.200 111.600 522.000 111.700 ;
        RECT 530.800 111.600 531.600 111.700 ;
        RECT 537.200 111.600 538.000 111.700 ;
        RECT 569.200 112.300 570.000 112.400 ;
        RECT 604.400 112.300 605.200 112.400 ;
        RECT 569.200 111.700 605.200 112.300 ;
        RECT 569.200 111.600 570.000 111.700 ;
        RECT 604.400 111.600 605.200 111.700 ;
        RECT 441.200 109.700 448.300 110.300 ;
        RECT 455.600 110.300 456.400 110.400 ;
        RECT 468.400 110.300 469.200 110.400 ;
        RECT 455.600 109.700 469.200 110.300 ;
        RECT 441.200 109.600 442.000 109.700 ;
        RECT 455.600 109.600 456.400 109.700 ;
        RECT 468.400 109.600 469.200 109.700 ;
        RECT 476.400 110.300 477.200 110.400 ;
        RECT 481.200 110.300 482.000 110.400 ;
        RECT 476.400 109.700 482.000 110.300 ;
        RECT 476.400 109.600 477.200 109.700 ;
        RECT 481.200 109.600 482.000 109.700 ;
        RECT 482.800 110.300 483.600 110.400 ;
        RECT 489.200 110.300 490.000 110.400 ;
        RECT 482.800 109.700 490.000 110.300 ;
        RECT 482.800 109.600 483.600 109.700 ;
        RECT 489.200 109.600 490.000 109.700 ;
        RECT 503.600 110.300 504.400 110.400 ;
        RECT 514.800 110.300 515.600 110.400 ;
        RECT 503.600 109.700 515.600 110.300 ;
        RECT 503.600 109.600 504.400 109.700 ;
        RECT 514.800 109.600 515.600 109.700 ;
        RECT 518.000 110.300 518.800 110.400 ;
        RECT 526.000 110.300 526.800 110.400 ;
        RECT 518.000 109.700 526.800 110.300 ;
        RECT 518.000 109.600 518.800 109.700 ;
        RECT 526.000 109.600 526.800 109.700 ;
        RECT 529.200 110.300 530.000 110.400 ;
        RECT 548.400 110.300 549.200 110.400 ;
        RECT 529.200 109.700 549.200 110.300 ;
        RECT 529.200 109.600 530.000 109.700 ;
        RECT 548.400 109.600 549.200 109.700 ;
        RECT 564.400 110.300 565.200 110.400 ;
        RECT 570.800 110.300 571.600 110.400 ;
        RECT 564.400 109.700 571.600 110.300 ;
        RECT 564.400 109.600 565.200 109.700 ;
        RECT 570.800 109.600 571.600 109.700 ;
        RECT 599.600 110.300 600.400 110.400 ;
        RECT 606.000 110.300 606.800 110.400 ;
        RECT 607.600 110.300 608.400 110.400 ;
        RECT 599.600 109.700 608.400 110.300 ;
        RECT 599.600 109.600 600.400 109.700 ;
        RECT 606.000 109.600 606.800 109.700 ;
        RECT 607.600 109.600 608.400 109.700 ;
        RECT 20.400 108.300 21.200 108.400 ;
        RECT 26.800 108.300 27.600 108.400 ;
        RECT 20.400 107.700 27.600 108.300 ;
        RECT 20.400 107.600 21.200 107.700 ;
        RECT 26.800 107.600 27.600 107.700 ;
        RECT 34.800 108.300 35.600 108.400 ;
        RECT 47.600 108.300 48.400 108.400 ;
        RECT 49.200 108.300 50.000 108.400 ;
        RECT 34.800 107.700 50.000 108.300 ;
        RECT 34.800 107.600 35.600 107.700 ;
        RECT 47.600 107.600 48.400 107.700 ;
        RECT 49.200 107.600 50.000 107.700 ;
        RECT 97.200 108.300 98.000 108.400 ;
        RECT 102.000 108.300 102.800 108.400 ;
        RECT 97.200 107.700 102.800 108.300 ;
        RECT 97.200 107.600 98.000 107.700 ;
        RECT 102.000 107.600 102.800 107.700 ;
        RECT 113.200 108.300 114.000 108.400 ;
        RECT 121.200 108.300 122.000 108.400 ;
        RECT 113.200 107.700 122.000 108.300 ;
        RECT 113.200 107.600 114.000 107.700 ;
        RECT 121.200 107.600 122.000 107.700 ;
        RECT 127.600 108.300 128.400 108.400 ;
        RECT 138.800 108.300 139.600 108.400 ;
        RECT 146.800 108.300 147.600 108.400 ;
        RECT 127.600 107.700 147.600 108.300 ;
        RECT 127.600 107.600 128.400 107.700 ;
        RECT 138.800 107.600 139.600 107.700 ;
        RECT 146.800 107.600 147.600 107.700 ;
        RECT 180.400 108.300 181.200 108.400 ;
        RECT 186.800 108.300 187.600 108.400 ;
        RECT 180.400 107.700 187.600 108.300 ;
        RECT 180.400 107.600 181.200 107.700 ;
        RECT 186.800 107.600 187.600 107.700 ;
        RECT 191.600 108.300 192.400 108.400 ;
        RECT 209.200 108.300 210.000 108.400 ;
        RECT 217.200 108.300 218.000 108.400 ;
        RECT 218.800 108.300 219.600 108.400 ;
        RECT 226.800 108.300 227.600 108.400 ;
        RECT 279.600 108.300 280.400 108.400 ;
        RECT 191.600 107.700 227.600 108.300 ;
        RECT 191.600 107.600 192.400 107.700 ;
        RECT 209.200 107.600 210.000 107.700 ;
        RECT 217.200 107.600 218.000 107.700 ;
        RECT 218.800 107.600 219.600 107.700 ;
        RECT 226.800 107.600 227.600 107.700 ;
        RECT 234.900 107.700 280.400 108.300 ;
        RECT 234.900 106.400 235.500 107.700 ;
        RECT 279.600 107.600 280.400 107.700 ;
        RECT 281.200 108.300 282.000 108.400 ;
        RECT 292.400 108.300 293.200 108.400 ;
        RECT 281.200 107.700 293.200 108.300 ;
        RECT 281.200 107.600 282.000 107.700 ;
        RECT 292.400 107.600 293.200 107.700 ;
        RECT 295.600 108.300 296.400 108.400 ;
        RECT 302.000 108.300 302.800 108.400 ;
        RECT 295.600 107.700 302.800 108.300 ;
        RECT 295.600 107.600 296.400 107.700 ;
        RECT 302.000 107.600 302.800 107.700 ;
        RECT 318.000 108.300 318.800 108.400 ;
        RECT 334.000 108.300 334.800 108.400 ;
        RECT 318.000 107.700 334.800 108.300 ;
        RECT 318.000 107.600 318.800 107.700 ;
        RECT 334.000 107.600 334.800 107.700 ;
        RECT 353.200 108.300 354.000 108.400 ;
        RECT 364.400 108.300 365.200 108.400 ;
        RECT 353.200 107.700 365.200 108.300 ;
        RECT 353.200 107.600 354.000 107.700 ;
        RECT 364.400 107.600 365.200 107.700 ;
        RECT 369.200 108.300 370.000 108.400 ;
        RECT 383.600 108.300 384.400 108.400 ;
        RECT 369.200 107.700 384.400 108.300 ;
        RECT 369.200 107.600 370.000 107.700 ;
        RECT 383.600 107.600 384.400 107.700 ;
        RECT 407.600 108.300 408.400 108.400 ;
        RECT 410.800 108.300 411.600 108.400 ;
        RECT 407.600 107.700 411.600 108.300 ;
        RECT 407.600 107.600 408.400 107.700 ;
        RECT 410.800 107.600 411.600 107.700 ;
        RECT 442.800 108.300 443.600 108.400 ;
        RECT 462.000 108.300 462.800 108.400 ;
        RECT 442.800 107.700 462.800 108.300 ;
        RECT 442.800 107.600 443.600 107.700 ;
        RECT 462.000 107.600 462.800 107.700 ;
        RECT 471.600 108.300 472.400 108.400 ;
        RECT 478.000 108.300 478.800 108.400 ;
        RECT 471.600 107.700 478.800 108.300 ;
        RECT 471.600 107.600 472.400 107.700 ;
        RECT 478.000 107.600 478.800 107.700 ;
        RECT 490.800 108.300 491.600 108.400 ;
        RECT 494.000 108.300 494.800 108.400 ;
        RECT 500.400 108.300 501.200 108.400 ;
        RECT 508.400 108.300 509.200 108.400 ;
        RECT 511.600 108.300 512.400 108.400 ;
        RECT 490.800 107.700 512.400 108.300 ;
        RECT 490.800 107.600 491.600 107.700 ;
        RECT 494.000 107.600 494.800 107.700 ;
        RECT 500.400 107.600 501.200 107.700 ;
        RECT 508.400 107.600 509.200 107.700 ;
        RECT 511.600 107.600 512.400 107.700 ;
        RECT 535.600 108.300 536.400 108.400 ;
        RECT 538.800 108.300 539.600 108.400 ;
        RECT 562.800 108.300 563.600 108.400 ;
        RECT 567.600 108.300 568.400 108.400 ;
        RECT 535.600 107.700 568.400 108.300 ;
        RECT 535.600 107.600 536.400 107.700 ;
        RECT 538.800 107.600 539.600 107.700 ;
        RECT 562.800 107.600 563.600 107.700 ;
        RECT 567.600 107.600 568.400 107.700 ;
        RECT 590.000 108.300 590.800 108.400 ;
        RECT 604.400 108.300 605.200 108.400 ;
        RECT 590.000 107.700 605.200 108.300 ;
        RECT 590.000 107.600 590.800 107.700 ;
        RECT 604.400 107.600 605.200 107.700 ;
        RECT 25.200 106.300 26.000 106.400 ;
        RECT 26.800 106.300 27.600 106.400 ;
        RECT 60.400 106.300 61.200 106.400 ;
        RECT 25.200 105.700 61.200 106.300 ;
        RECT 25.200 105.600 26.000 105.700 ;
        RECT 26.800 105.600 27.600 105.700 ;
        RECT 60.400 105.600 61.200 105.700 ;
        RECT 106.800 106.300 107.600 106.400 ;
        RECT 108.400 106.300 109.200 106.400 ;
        RECT 106.800 105.700 109.200 106.300 ;
        RECT 106.800 105.600 107.600 105.700 ;
        RECT 108.400 105.600 109.200 105.700 ;
        RECT 124.400 106.300 125.200 106.400 ;
        RECT 156.400 106.300 157.200 106.400 ;
        RECT 183.600 106.300 184.400 106.400 ;
        RECT 210.800 106.300 211.600 106.400 ;
        RECT 234.800 106.300 235.600 106.400 ;
        RECT 124.400 105.700 235.600 106.300 ;
        RECT 124.400 105.600 125.200 105.700 ;
        RECT 156.400 105.600 157.200 105.700 ;
        RECT 183.600 105.600 184.400 105.700 ;
        RECT 210.800 105.600 211.600 105.700 ;
        RECT 234.800 105.600 235.600 105.700 ;
        RECT 236.400 106.300 237.200 106.400 ;
        RECT 241.200 106.300 242.000 106.400 ;
        RECT 257.200 106.300 258.000 106.400 ;
        RECT 236.400 105.700 258.000 106.300 ;
        RECT 236.400 105.600 237.200 105.700 ;
        RECT 241.200 105.600 242.000 105.700 ;
        RECT 257.200 105.600 258.000 105.700 ;
        RECT 289.200 106.300 290.000 106.400 ;
        RECT 308.400 106.300 309.200 106.400 ;
        RECT 353.300 106.300 353.900 107.600 ;
        RECT 289.200 105.700 353.900 106.300 ;
        RECT 382.000 106.300 382.800 106.400 ;
        RECT 444.400 106.300 445.200 106.400 ;
        RECT 382.000 105.700 445.200 106.300 ;
        RECT 289.200 105.600 290.000 105.700 ;
        RECT 308.400 105.600 309.200 105.700 ;
        RECT 382.000 105.600 382.800 105.700 ;
        RECT 444.400 105.600 445.200 105.700 ;
        RECT 447.600 106.300 448.400 106.400 ;
        RECT 449.200 106.300 450.000 106.400 ;
        RECT 468.400 106.300 469.200 106.400 ;
        RECT 447.600 105.700 469.200 106.300 ;
        RECT 447.600 105.600 448.400 105.700 ;
        RECT 449.200 105.600 450.000 105.700 ;
        RECT 468.400 105.600 469.200 105.700 ;
        RECT 506.800 106.300 507.600 106.400 ;
        RECT 521.200 106.300 522.000 106.400 ;
        RECT 506.800 105.700 522.000 106.300 ;
        RECT 506.800 105.600 507.600 105.700 ;
        RECT 521.200 105.600 522.000 105.700 ;
        RECT 553.200 106.300 554.000 106.400 ;
        RECT 586.800 106.300 587.600 106.400 ;
        RECT 553.200 105.700 587.600 106.300 ;
        RECT 553.200 105.600 554.000 105.700 ;
        RECT 586.800 105.600 587.600 105.700 ;
        RECT 20.400 104.300 21.200 104.400 ;
        RECT 39.600 104.300 40.400 104.400 ;
        RECT 20.400 103.700 40.400 104.300 ;
        RECT 20.400 103.600 21.200 103.700 ;
        RECT 39.600 103.600 40.400 103.700 ;
        RECT 44.400 104.300 45.200 104.400 ;
        RECT 46.000 104.300 46.800 104.400 ;
        RECT 44.400 103.700 46.800 104.300 ;
        RECT 44.400 103.600 45.200 103.700 ;
        RECT 46.000 103.600 46.800 103.700 ;
        RECT 145.200 104.300 146.000 104.400 ;
        RECT 158.000 104.300 158.800 104.400 ;
        RECT 174.000 104.300 174.800 104.400 ;
        RECT 204.400 104.300 205.200 104.400 ;
        RECT 145.200 103.700 205.200 104.300 ;
        RECT 145.200 103.600 146.000 103.700 ;
        RECT 158.000 103.600 158.800 103.700 ;
        RECT 174.000 103.600 174.800 103.700 ;
        RECT 204.400 103.600 205.200 103.700 ;
        RECT 215.600 104.300 216.400 104.400 ;
        RECT 223.600 104.300 224.400 104.400 ;
        RECT 215.600 103.700 224.400 104.300 ;
        RECT 215.600 103.600 216.400 103.700 ;
        RECT 223.600 103.600 224.400 103.700 ;
        RECT 242.800 104.300 243.600 104.400 ;
        RECT 247.600 104.300 248.400 104.400 ;
        RECT 242.800 103.700 248.400 104.300 ;
        RECT 242.800 103.600 243.600 103.700 ;
        RECT 247.600 103.600 248.400 103.700 ;
        RECT 404.400 104.300 405.200 104.400 ;
        RECT 449.200 104.300 450.000 104.400 ;
        RECT 404.400 103.700 450.000 104.300 ;
        RECT 404.400 103.600 405.200 103.700 ;
        RECT 449.200 103.600 450.000 103.700 ;
        RECT 452.400 104.300 453.200 104.400 ;
        RECT 514.800 104.300 515.600 104.400 ;
        RECT 566.000 104.300 566.800 104.400 ;
        RECT 452.400 103.700 510.700 104.300 ;
        RECT 452.400 103.600 453.200 103.700 ;
        RECT 39.600 102.300 40.400 102.400 ;
        RECT 89.200 102.300 90.000 102.400 ;
        RECT 271.600 102.300 272.400 102.400 ;
        RECT 39.600 101.700 90.000 102.300 ;
        RECT 39.600 101.600 40.400 101.700 ;
        RECT 89.200 101.600 90.000 101.700 ;
        RECT 255.700 101.700 272.400 102.300 ;
        RECT 255.700 100.400 256.300 101.700 ;
        RECT 271.600 101.600 272.400 101.700 ;
        RECT 362.800 102.300 363.600 102.400 ;
        RECT 401.200 102.300 402.000 102.400 ;
        RECT 402.800 102.300 403.600 102.400 ;
        RECT 362.800 101.700 403.600 102.300 ;
        RECT 362.800 101.600 363.600 101.700 ;
        RECT 401.200 101.600 402.000 101.700 ;
        RECT 402.800 101.600 403.600 101.700 ;
        RECT 410.800 102.300 411.600 102.400 ;
        RECT 434.800 102.300 435.600 102.400 ;
        RECT 463.600 102.300 464.400 102.400 ;
        RECT 486.000 102.300 486.800 102.400 ;
        RECT 508.400 102.300 509.200 102.400 ;
        RECT 410.800 101.700 509.200 102.300 ;
        RECT 510.100 102.300 510.700 103.700 ;
        RECT 514.800 103.700 566.800 104.300 ;
        RECT 514.800 103.600 515.600 103.700 ;
        RECT 566.000 103.600 566.800 103.700 ;
        RECT 570.800 104.300 571.600 104.400 ;
        RECT 572.400 104.300 573.200 104.400 ;
        RECT 570.800 103.700 573.200 104.300 ;
        RECT 570.800 103.600 571.600 103.700 ;
        RECT 572.400 103.600 573.200 103.700 ;
        RECT 521.200 102.300 522.000 102.400 ;
        RECT 556.400 102.300 557.200 102.400 ;
        RECT 510.100 101.700 557.200 102.300 ;
        RECT 410.800 101.600 411.600 101.700 ;
        RECT 434.800 101.600 435.600 101.700 ;
        RECT 463.600 101.600 464.400 101.700 ;
        RECT 486.000 101.600 486.800 101.700 ;
        RECT 508.400 101.600 509.200 101.700 ;
        RECT 521.200 101.600 522.000 101.700 ;
        RECT 556.400 101.600 557.200 101.700 ;
        RECT 137.200 100.300 138.000 100.400 ;
        RECT 255.600 100.300 256.400 100.400 ;
        RECT 137.200 99.700 256.400 100.300 ;
        RECT 137.200 99.600 138.000 99.700 ;
        RECT 255.600 99.600 256.400 99.700 ;
        RECT 260.400 100.300 261.200 100.400 ;
        RECT 266.800 100.300 267.600 100.400 ;
        RECT 260.400 99.700 267.600 100.300 ;
        RECT 260.400 99.600 261.200 99.700 ;
        RECT 266.800 99.600 267.600 99.700 ;
        RECT 348.400 100.300 349.200 100.400 ;
        RECT 382.000 100.300 382.800 100.400 ;
        RECT 386.800 100.300 387.600 100.400 ;
        RECT 348.400 99.700 387.600 100.300 ;
        RECT 348.400 99.600 349.200 99.700 ;
        RECT 382.000 99.600 382.800 99.700 ;
        RECT 386.800 99.600 387.600 99.700 ;
        RECT 418.800 100.300 419.600 100.400 ;
        RECT 441.200 100.300 442.000 100.400 ;
        RECT 418.800 99.700 442.000 100.300 ;
        RECT 418.800 99.600 419.600 99.700 ;
        RECT 441.200 99.600 442.000 99.700 ;
        RECT 450.800 100.300 451.600 100.400 ;
        RECT 482.800 100.300 483.600 100.400 ;
        RECT 450.800 99.700 483.600 100.300 ;
        RECT 450.800 99.600 451.600 99.700 ;
        RECT 482.800 99.600 483.600 99.700 ;
        RECT 495.600 100.300 496.400 100.400 ;
        RECT 542.000 100.300 542.800 100.400 ;
        RECT 495.600 99.700 542.800 100.300 ;
        RECT 495.600 99.600 496.400 99.700 ;
        RECT 542.000 99.600 542.800 99.700 ;
        RECT 31.600 98.300 32.400 98.400 ;
        RECT 42.800 98.300 43.600 98.400 ;
        RECT 31.600 97.700 43.600 98.300 ;
        RECT 31.600 97.600 32.400 97.700 ;
        RECT 42.800 97.600 43.600 97.700 ;
        RECT 60.400 98.300 61.200 98.400 ;
        RECT 73.200 98.300 74.000 98.400 ;
        RECT 79.600 98.300 80.400 98.400 ;
        RECT 60.400 97.700 80.400 98.300 ;
        RECT 60.400 97.600 61.200 97.700 ;
        RECT 73.200 97.600 74.000 97.700 ;
        RECT 79.600 97.600 80.400 97.700 ;
        RECT 226.800 98.300 227.600 98.400 ;
        RECT 239.600 98.300 240.400 98.400 ;
        RECT 226.800 97.700 240.400 98.300 ;
        RECT 226.800 97.600 227.600 97.700 ;
        RECT 239.600 97.600 240.400 97.700 ;
        RECT 332.400 98.300 333.200 98.400 ;
        RECT 334.000 98.300 334.800 98.400 ;
        RECT 332.400 97.700 334.800 98.300 ;
        RECT 332.400 97.600 333.200 97.700 ;
        RECT 334.000 97.600 334.800 97.700 ;
        RECT 428.400 98.300 429.200 98.400 ;
        RECT 484.400 98.300 485.200 98.400 ;
        RECT 497.200 98.300 498.000 98.400 ;
        RECT 428.400 97.700 498.000 98.300 ;
        RECT 428.400 97.600 429.200 97.700 ;
        RECT 484.400 97.600 485.200 97.700 ;
        RECT 497.200 97.600 498.000 97.700 ;
        RECT 506.800 98.300 507.600 98.400 ;
        RECT 548.400 98.300 549.200 98.400 ;
        RECT 506.800 97.700 549.200 98.300 ;
        RECT 506.800 97.600 507.600 97.700 ;
        RECT 548.400 97.600 549.200 97.700 ;
        RECT 562.800 98.300 563.600 98.400 ;
        RECT 569.200 98.300 570.000 98.400 ;
        RECT 586.800 98.300 587.600 98.400 ;
        RECT 562.800 97.700 587.600 98.300 ;
        RECT 562.800 97.600 563.600 97.700 ;
        RECT 569.200 97.600 570.000 97.700 ;
        RECT 586.800 97.600 587.600 97.700 ;
        RECT 588.400 98.300 589.200 98.400 ;
        RECT 596.400 98.300 597.200 98.400 ;
        RECT 588.400 97.700 597.200 98.300 ;
        RECT 588.400 97.600 589.200 97.700 ;
        RECT 596.400 97.600 597.200 97.700 ;
        RECT 602.800 98.300 603.600 98.400 ;
        RECT 607.600 98.300 608.400 98.400 ;
        RECT 602.800 97.700 608.400 98.300 ;
        RECT 602.800 97.600 603.600 97.700 ;
        RECT 607.600 97.600 608.400 97.700 ;
        RECT 23.600 96.300 24.400 96.400 ;
        RECT 36.400 96.300 37.200 96.400 ;
        RECT 23.600 95.700 37.200 96.300 ;
        RECT 23.600 95.600 24.400 95.700 ;
        RECT 36.400 95.600 37.200 95.700 ;
        RECT 58.800 96.300 59.600 96.400 ;
        RECT 68.400 96.300 69.200 96.400 ;
        RECT 58.800 95.700 69.200 96.300 ;
        RECT 58.800 95.600 59.600 95.700 ;
        RECT 68.400 95.600 69.200 95.700 ;
        RECT 71.600 96.300 72.400 96.400 ;
        RECT 79.600 96.300 80.400 96.400 ;
        RECT 71.600 95.700 80.400 96.300 ;
        RECT 71.600 95.600 72.400 95.700 ;
        RECT 79.600 95.600 80.400 95.700 ;
        RECT 92.400 96.300 93.200 96.400 ;
        RECT 105.200 96.300 106.000 96.400 ;
        RECT 113.200 96.300 114.000 96.400 ;
        RECT 132.400 96.300 133.200 96.400 ;
        RECT 92.400 95.700 133.200 96.300 ;
        RECT 92.400 95.600 93.200 95.700 ;
        RECT 105.200 95.600 106.000 95.700 ;
        RECT 113.200 95.600 114.000 95.700 ;
        RECT 132.400 95.600 133.200 95.700 ;
        RECT 226.800 96.300 227.600 96.400 ;
        RECT 231.600 96.300 232.400 96.400 ;
        RECT 244.400 96.300 245.200 96.400 ;
        RECT 250.800 96.300 251.600 96.400 ;
        RECT 226.800 95.700 251.600 96.300 ;
        RECT 226.800 95.600 227.600 95.700 ;
        RECT 231.600 95.600 232.400 95.700 ;
        RECT 244.400 95.600 245.200 95.700 ;
        RECT 250.800 95.600 251.600 95.700 ;
        RECT 300.400 96.300 301.200 96.400 ;
        RECT 330.800 96.300 331.600 96.400 ;
        RECT 300.400 95.700 331.600 96.300 ;
        RECT 300.400 95.600 301.200 95.700 ;
        RECT 330.800 95.600 331.600 95.700 ;
        RECT 420.400 96.300 421.200 96.400 ;
        RECT 447.600 96.300 448.400 96.400 ;
        RECT 420.400 95.700 448.400 96.300 ;
        RECT 420.400 95.600 421.200 95.700 ;
        RECT 447.600 95.600 448.400 95.700 ;
        RECT 452.400 96.300 453.200 96.400 ;
        RECT 463.600 96.300 464.400 96.400 ;
        RECT 452.400 95.700 464.400 96.300 ;
        RECT 452.400 95.600 453.200 95.700 ;
        RECT 463.600 95.600 464.400 95.700 ;
        RECT 466.800 96.300 467.600 96.400 ;
        RECT 510.000 96.300 510.800 96.400 ;
        RECT 524.400 96.300 525.200 96.400 ;
        RECT 527.600 96.300 528.400 96.400 ;
        RECT 466.800 95.700 475.500 96.300 ;
        RECT 466.800 95.600 467.600 95.700 ;
        RECT 22.000 94.300 22.800 94.400 ;
        RECT 25.200 94.300 26.000 94.400 ;
        RECT 33.200 94.300 34.000 94.400 ;
        RECT 22.000 93.700 34.000 94.300 ;
        RECT 22.000 93.600 22.800 93.700 ;
        RECT 25.200 93.600 26.000 93.700 ;
        RECT 33.200 93.600 34.000 93.700 ;
        RECT 34.800 94.300 35.600 94.400 ;
        RECT 63.600 94.300 64.400 94.400 ;
        RECT 34.800 93.700 64.400 94.300 ;
        RECT 34.800 93.600 35.600 93.700 ;
        RECT 63.600 93.600 64.400 93.700 ;
        RECT 81.200 94.300 82.000 94.400 ;
        RECT 82.800 94.300 83.600 94.400 ;
        RECT 81.200 93.700 83.600 94.300 ;
        RECT 81.200 93.600 82.000 93.700 ;
        RECT 82.800 93.600 83.600 93.700 ;
        RECT 97.200 93.600 98.000 94.400 ;
        RECT 119.600 94.300 120.400 94.400 ;
        RECT 127.600 94.300 128.400 94.400 ;
        RECT 119.600 93.700 128.400 94.300 ;
        RECT 119.600 93.600 120.400 93.700 ;
        RECT 127.600 93.600 128.400 93.700 ;
        RECT 178.800 94.300 179.600 94.400 ;
        RECT 190.000 94.300 190.800 94.400 ;
        RECT 178.800 93.700 190.800 94.300 ;
        RECT 178.800 93.600 179.600 93.700 ;
        RECT 190.000 93.600 190.800 93.700 ;
        RECT 222.000 94.300 222.800 94.400 ;
        RECT 241.200 94.300 242.000 94.400 ;
        RECT 295.600 94.300 296.400 94.400 ;
        RECT 316.400 94.300 317.200 94.400 ;
        RECT 222.000 93.700 317.200 94.300 ;
        RECT 222.000 93.600 222.800 93.700 ;
        RECT 241.200 93.600 242.000 93.700 ;
        RECT 295.600 93.600 296.400 93.700 ;
        RECT 316.400 93.600 317.200 93.700 ;
        RECT 351.600 94.300 352.400 94.400 ;
        RECT 359.600 94.300 360.400 94.400 ;
        RECT 351.600 93.700 360.400 94.300 ;
        RECT 351.600 93.600 352.400 93.700 ;
        RECT 359.600 93.600 360.400 93.700 ;
        RECT 407.600 94.300 408.400 94.400 ;
        RECT 414.000 94.300 414.800 94.400 ;
        RECT 407.600 93.700 414.800 94.300 ;
        RECT 407.600 93.600 408.400 93.700 ;
        RECT 414.000 93.600 414.800 93.700 ;
        RECT 433.200 94.300 434.000 94.400 ;
        RECT 438.000 94.300 438.800 94.400 ;
        RECT 447.600 94.300 448.400 94.400 ;
        RECT 433.200 93.700 448.400 94.300 ;
        RECT 433.200 93.600 434.000 93.700 ;
        RECT 438.000 93.600 438.800 93.700 ;
        RECT 447.600 93.600 448.400 93.700 ;
        RECT 455.600 94.300 456.400 94.400 ;
        RECT 473.200 94.300 474.000 94.400 ;
        RECT 455.600 93.700 474.000 94.300 ;
        RECT 474.900 94.300 475.500 95.700 ;
        RECT 510.000 95.700 528.400 96.300 ;
        RECT 510.000 95.600 510.800 95.700 ;
        RECT 524.400 95.600 525.200 95.700 ;
        RECT 527.600 95.600 528.400 95.700 ;
        RECT 534.000 96.300 534.800 96.400 ;
        RECT 537.200 96.300 538.000 96.400 ;
        RECT 534.000 95.700 538.000 96.300 ;
        RECT 534.000 95.600 534.800 95.700 ;
        RECT 537.200 95.600 538.000 95.700 ;
        RECT 561.200 96.300 562.000 96.400 ;
        RECT 591.600 96.300 592.400 96.400 ;
        RECT 561.200 95.700 592.400 96.300 ;
        RECT 561.200 95.600 562.000 95.700 ;
        RECT 591.600 95.600 592.400 95.700 ;
        RECT 503.600 94.300 504.400 94.400 ;
        RECT 474.900 93.700 504.400 94.300 ;
        RECT 455.600 93.600 456.400 93.700 ;
        RECT 473.200 93.600 474.000 93.700 ;
        RECT 503.600 93.600 504.400 93.700 ;
        RECT 511.600 94.300 512.400 94.400 ;
        RECT 540.400 94.300 541.200 94.400 ;
        RECT 564.400 94.300 565.200 94.400 ;
        RECT 511.600 93.700 565.200 94.300 ;
        RECT 511.600 93.600 512.400 93.700 ;
        RECT 540.400 93.600 541.200 93.700 ;
        RECT 564.400 93.600 565.200 93.700 ;
        RECT 28.400 92.300 29.200 92.400 ;
        RECT 36.400 92.300 37.200 92.400 ;
        RECT 28.400 91.700 37.200 92.300 ;
        RECT 28.400 91.600 29.200 91.700 ;
        RECT 36.400 91.600 37.200 91.700 ;
        RECT 41.200 92.300 42.000 92.400 ;
        RECT 74.800 92.300 75.600 92.400 ;
        RECT 41.200 91.700 75.600 92.300 ;
        RECT 41.200 91.600 42.000 91.700 ;
        RECT 74.800 91.600 75.600 91.700 ;
        RECT 84.400 92.300 85.200 92.400 ;
        RECT 87.600 92.300 88.400 92.400 ;
        RECT 84.400 91.700 88.400 92.300 ;
        RECT 84.400 91.600 85.200 91.700 ;
        RECT 87.600 91.600 88.400 91.700 ;
        RECT 100.400 92.300 101.200 92.400 ;
        RECT 118.000 92.300 118.800 92.400 ;
        RECT 129.200 92.300 130.000 92.400 ;
        RECT 137.200 92.300 138.000 92.400 ;
        RECT 100.400 91.700 138.000 92.300 ;
        RECT 100.400 91.600 101.200 91.700 ;
        RECT 118.000 91.600 118.800 91.700 ;
        RECT 129.200 91.600 130.000 91.700 ;
        RECT 137.200 91.600 138.000 91.700 ;
        RECT 212.400 92.300 213.200 92.400 ;
        RECT 215.600 92.300 216.400 92.400 ;
        RECT 212.400 91.700 216.400 92.300 ;
        RECT 212.400 91.600 213.200 91.700 ;
        RECT 215.600 91.600 216.400 91.700 ;
        RECT 217.200 92.300 218.000 92.400 ;
        RECT 226.800 92.300 227.600 92.400 ;
        RECT 217.200 91.700 227.600 92.300 ;
        RECT 217.200 91.600 218.000 91.700 ;
        RECT 226.800 91.600 227.600 91.700 ;
        RECT 239.600 92.300 240.400 92.400 ;
        RECT 270.000 92.300 270.800 92.400 ;
        RECT 239.600 91.700 270.800 92.300 ;
        RECT 239.600 91.600 240.400 91.700 ;
        RECT 270.000 91.600 270.800 91.700 ;
        RECT 279.600 92.300 280.400 92.400 ;
        RECT 287.600 92.300 288.400 92.400 ;
        RECT 279.600 91.700 288.400 92.300 ;
        RECT 279.600 91.600 280.400 91.700 ;
        RECT 287.600 91.600 288.400 91.700 ;
        RECT 358.000 92.300 358.800 92.400 ;
        RECT 366.000 92.300 366.800 92.400 ;
        RECT 369.200 92.300 370.000 92.400 ;
        RECT 358.000 91.700 370.000 92.300 ;
        RECT 358.000 91.600 358.800 91.700 ;
        RECT 366.000 91.600 366.800 91.700 ;
        RECT 369.200 91.600 370.000 91.700 ;
        RECT 425.200 92.300 426.000 92.400 ;
        RECT 430.000 92.300 430.800 92.400 ;
        RECT 433.200 92.300 434.000 92.400 ;
        RECT 425.200 91.700 434.000 92.300 ;
        RECT 425.200 91.600 426.000 91.700 ;
        RECT 430.000 91.600 430.800 91.700 ;
        RECT 433.200 91.600 434.000 91.700 ;
        RECT 436.400 91.600 437.200 92.400 ;
        RECT 441.200 92.300 442.000 92.400 ;
        RECT 442.800 92.300 443.600 92.400 ;
        RECT 441.200 91.700 443.600 92.300 ;
        RECT 441.200 91.600 442.000 91.700 ;
        RECT 442.800 91.600 443.600 91.700 ;
        RECT 449.200 92.300 450.000 92.400 ;
        RECT 455.600 92.300 456.400 92.400 ;
        RECT 449.200 91.700 456.400 92.300 ;
        RECT 449.200 91.600 450.000 91.700 ;
        RECT 455.600 91.600 456.400 91.700 ;
        RECT 465.200 92.300 466.000 92.400 ;
        RECT 474.800 92.300 475.600 92.400 ;
        RECT 465.200 91.700 475.600 92.300 ;
        RECT 465.200 91.600 466.000 91.700 ;
        RECT 474.800 91.600 475.600 91.700 ;
        RECT 479.600 92.300 480.400 92.400 ;
        RECT 490.800 92.300 491.600 92.400 ;
        RECT 479.600 91.700 491.600 92.300 ;
        RECT 479.600 91.600 480.400 91.700 ;
        RECT 490.800 91.600 491.600 91.700 ;
        RECT 492.400 92.300 493.200 92.400 ;
        RECT 498.800 92.300 499.600 92.400 ;
        RECT 492.400 91.700 499.600 92.300 ;
        RECT 492.400 91.600 493.200 91.700 ;
        RECT 498.800 91.600 499.600 91.700 ;
        RECT 518.000 92.300 518.800 92.400 ;
        RECT 522.800 92.300 523.600 92.400 ;
        RECT 518.000 91.700 523.600 92.300 ;
        RECT 518.000 91.600 518.800 91.700 ;
        RECT 522.800 91.600 523.600 91.700 ;
        RECT 532.400 92.300 533.200 92.400 ;
        RECT 556.400 92.300 557.200 92.400 ;
        RECT 532.400 91.700 557.200 92.300 ;
        RECT 532.400 91.600 533.200 91.700 ;
        RECT 556.400 91.600 557.200 91.700 ;
        RECT 570.800 92.300 571.600 92.400 ;
        RECT 601.200 92.300 602.000 92.400 ;
        RECT 570.800 91.700 602.000 92.300 ;
        RECT 570.800 91.600 571.600 91.700 ;
        RECT 601.200 91.600 602.000 91.700 ;
        RECT 14.000 90.300 14.800 90.400 ;
        RECT 28.400 90.300 29.200 90.400 ;
        RECT 14.000 89.700 29.200 90.300 ;
        RECT 14.000 89.600 14.800 89.700 ;
        RECT 28.400 89.600 29.200 89.700 ;
        RECT 39.600 90.300 40.400 90.400 ;
        RECT 42.800 90.300 43.600 90.400 ;
        RECT 39.600 89.700 43.600 90.300 ;
        RECT 39.600 89.600 40.400 89.700 ;
        RECT 42.800 89.600 43.600 89.700 ;
        RECT 66.800 90.300 67.600 90.400 ;
        RECT 76.400 90.300 77.200 90.400 ;
        RECT 66.800 89.700 77.200 90.300 ;
        RECT 66.800 89.600 67.600 89.700 ;
        RECT 76.400 89.600 77.200 89.700 ;
        RECT 94.000 90.300 94.800 90.400 ;
        RECT 106.800 90.300 107.600 90.400 ;
        RECT 110.000 90.300 110.800 90.400 ;
        RECT 94.000 89.700 110.800 90.300 ;
        RECT 94.000 89.600 94.800 89.700 ;
        RECT 106.800 89.600 107.600 89.700 ;
        RECT 110.000 89.600 110.800 89.700 ;
        RECT 111.600 90.300 112.400 90.400 ;
        RECT 121.200 90.300 122.000 90.400 ;
        RECT 130.800 90.300 131.600 90.400 ;
        RECT 142.000 90.300 142.800 90.400 ;
        RECT 111.600 89.700 142.800 90.300 ;
        RECT 111.600 89.600 112.400 89.700 ;
        RECT 121.200 89.600 122.000 89.700 ;
        RECT 130.800 89.600 131.600 89.700 ;
        RECT 142.000 89.600 142.800 89.700 ;
        RECT 204.400 90.300 205.200 90.400 ;
        RECT 212.400 90.300 213.200 90.400 ;
        RECT 204.400 89.700 213.200 90.300 ;
        RECT 204.400 89.600 205.200 89.700 ;
        RECT 212.400 89.600 213.200 89.700 ;
        RECT 215.600 90.300 216.400 90.400 ;
        RECT 234.800 90.300 235.600 90.400 ;
        RECT 215.600 89.700 235.600 90.300 ;
        RECT 215.600 89.600 216.400 89.700 ;
        RECT 234.800 89.600 235.600 89.700 ;
        RECT 425.200 90.300 426.000 90.400 ;
        RECT 444.400 90.300 445.200 90.400 ;
        RECT 425.200 89.700 445.200 90.300 ;
        RECT 425.200 89.600 426.000 89.700 ;
        RECT 444.400 89.600 445.200 89.700 ;
        RECT 449.200 90.300 450.000 90.400 ;
        RECT 457.200 90.300 458.000 90.400 ;
        RECT 449.200 89.700 458.000 90.300 ;
        RECT 449.200 89.600 450.000 89.700 ;
        RECT 457.200 89.600 458.000 89.700 ;
        RECT 476.400 90.300 477.200 90.400 ;
        RECT 519.600 90.300 520.400 90.400 ;
        RECT 534.000 90.300 534.800 90.400 ;
        RECT 545.200 90.300 546.000 90.400 ;
        RECT 476.400 89.700 546.000 90.300 ;
        RECT 476.400 89.600 477.200 89.700 ;
        RECT 519.600 89.600 520.400 89.700 ;
        RECT 534.000 89.600 534.800 89.700 ;
        RECT 545.200 89.600 546.000 89.700 ;
        RECT 567.600 90.300 568.400 90.400 ;
        RECT 574.000 90.300 574.800 90.400 ;
        RECT 567.600 89.700 574.800 90.300 ;
        RECT 567.600 89.600 568.400 89.700 ;
        RECT 574.000 89.600 574.800 89.700 ;
        RECT 1.200 88.300 2.000 88.400 ;
        RECT 39.700 88.300 40.300 89.600 ;
        RECT 1.200 87.700 40.300 88.300 ;
        RECT 65.200 88.300 66.000 88.400 ;
        RECT 68.400 88.300 69.200 88.400 ;
        RECT 65.200 87.700 69.200 88.300 ;
        RECT 76.500 88.300 77.100 89.600 ;
        RECT 103.600 88.300 104.400 88.400 ;
        RECT 76.500 87.700 104.400 88.300 ;
        RECT 1.200 87.600 2.000 87.700 ;
        RECT 65.200 87.600 66.000 87.700 ;
        RECT 68.400 87.600 69.200 87.700 ;
        RECT 103.600 87.600 104.400 87.700 ;
        RECT 108.400 88.300 109.200 88.400 ;
        RECT 114.800 88.300 115.600 88.400 ;
        RECT 108.400 87.700 115.600 88.300 ;
        RECT 108.400 87.600 109.200 87.700 ;
        RECT 114.800 87.600 115.600 87.700 ;
        RECT 124.400 88.300 125.200 88.400 ;
        RECT 132.400 88.300 133.200 88.400 ;
        RECT 124.400 87.700 133.200 88.300 ;
        RECT 124.400 87.600 125.200 87.700 ;
        RECT 132.400 87.600 133.200 87.700 ;
        RECT 135.600 87.600 136.400 88.400 ;
        RECT 140.400 88.300 141.200 88.400 ;
        RECT 146.800 88.300 147.600 88.400 ;
        RECT 140.400 87.700 147.600 88.300 ;
        RECT 140.400 87.600 141.200 87.700 ;
        RECT 146.800 87.600 147.600 87.700 ;
        RECT 415.600 88.300 416.400 88.400 ;
        RECT 428.400 88.300 429.200 88.400 ;
        RECT 415.600 87.700 429.200 88.300 ;
        RECT 415.600 87.600 416.400 87.700 ;
        RECT 428.400 87.600 429.200 87.700 ;
        RECT 513.200 88.300 514.000 88.400 ;
        RECT 524.400 88.300 525.200 88.400 ;
        RECT 569.200 88.300 570.000 88.400 ;
        RECT 513.200 87.700 570.000 88.300 ;
        RECT 513.200 87.600 514.000 87.700 ;
        RECT 524.400 87.600 525.200 87.700 ;
        RECT 569.200 87.600 570.000 87.700 ;
        RECT 73.200 86.300 74.000 86.400 ;
        RECT 84.400 86.300 85.200 86.400 ;
        RECT 73.200 85.700 85.200 86.300 ;
        RECT 73.200 85.600 74.000 85.700 ;
        RECT 84.400 85.600 85.200 85.700 ;
        RECT 106.800 85.600 107.600 86.400 ;
        RECT 132.500 86.300 133.100 87.600 ;
        RECT 143.600 86.300 144.400 86.400 ;
        RECT 175.600 86.300 176.400 86.400 ;
        RECT 132.500 85.700 176.400 86.300 ;
        RECT 143.600 85.600 144.400 85.700 ;
        RECT 175.600 85.600 176.400 85.700 ;
        RECT 458.800 86.300 459.600 86.400 ;
        RECT 561.200 86.300 562.000 86.400 ;
        RECT 458.800 85.700 562.000 86.300 ;
        RECT 458.800 85.600 459.600 85.700 ;
        RECT 561.200 85.600 562.000 85.700 ;
        RECT 62.000 84.300 62.800 84.400 ;
        RECT 90.800 84.300 91.600 84.400 ;
        RECT 62.000 83.700 91.600 84.300 ;
        RECT 62.000 83.600 62.800 83.700 ;
        RECT 90.800 83.600 91.600 83.700 ;
        RECT 398.000 84.300 398.800 84.400 ;
        RECT 406.000 84.300 406.800 84.400 ;
        RECT 425.200 84.300 426.000 84.400 ;
        RECT 398.000 83.700 426.000 84.300 ;
        RECT 398.000 83.600 398.800 83.700 ;
        RECT 406.000 83.600 406.800 83.700 ;
        RECT 425.200 83.600 426.000 83.700 ;
        RECT 430.000 84.300 430.800 84.400 ;
        RECT 478.000 84.300 478.800 84.400 ;
        RECT 430.000 83.700 478.800 84.300 ;
        RECT 430.000 83.600 430.800 83.700 ;
        RECT 478.000 83.600 478.800 83.700 ;
        RECT 38.000 82.300 38.800 82.400 ;
        RECT 52.400 82.300 53.200 82.400 ;
        RECT 38.000 81.700 53.200 82.300 ;
        RECT 38.000 81.600 38.800 81.700 ;
        RECT 52.400 81.600 53.200 81.700 ;
        RECT 78.000 82.300 78.800 82.400 ;
        RECT 98.800 82.300 99.600 82.400 ;
        RECT 78.000 81.700 99.600 82.300 ;
        RECT 78.000 81.600 78.800 81.700 ;
        RECT 98.800 81.600 99.600 81.700 ;
        RECT 122.800 82.300 123.600 82.400 ;
        RECT 138.800 82.300 139.600 82.400 ;
        RECT 122.800 81.700 139.600 82.300 ;
        RECT 122.800 81.600 123.600 81.700 ;
        RECT 138.800 81.600 139.600 81.700 ;
        RECT 170.800 82.300 171.600 82.400 ;
        RECT 186.800 82.300 187.600 82.400 ;
        RECT 170.800 81.700 187.600 82.300 ;
        RECT 170.800 81.600 171.600 81.700 ;
        RECT 186.800 81.600 187.600 81.700 ;
        RECT 378.800 82.300 379.600 82.400 ;
        RECT 398.000 82.300 398.800 82.400 ;
        RECT 378.800 81.700 398.800 82.300 ;
        RECT 378.800 81.600 379.600 81.700 ;
        RECT 398.000 81.600 398.800 81.700 ;
        RECT 465.200 82.300 466.000 82.400 ;
        RECT 500.400 82.300 501.200 82.400 ;
        RECT 522.800 82.300 523.600 82.400 ;
        RECT 465.200 81.700 523.600 82.300 ;
        RECT 465.200 81.600 466.000 81.700 ;
        RECT 500.400 81.600 501.200 81.700 ;
        RECT 522.800 81.600 523.600 81.700 ;
        RECT 562.800 82.300 563.600 82.400 ;
        RECT 606.000 82.300 606.800 82.400 ;
        RECT 562.800 81.700 606.800 82.300 ;
        RECT 562.800 81.600 563.600 81.700 ;
        RECT 606.000 81.600 606.800 81.700 ;
        RECT 161.200 80.300 162.000 80.400 ;
        RECT 190.000 80.300 190.800 80.400 ;
        RECT 161.200 79.700 190.800 80.300 ;
        RECT 161.200 79.600 162.000 79.700 ;
        RECT 190.000 79.600 190.800 79.700 ;
        RECT 207.600 80.300 208.400 80.400 ;
        RECT 246.000 80.300 246.800 80.400 ;
        RECT 284.400 80.300 285.200 80.400 ;
        RECT 207.600 79.700 285.200 80.300 ;
        RECT 207.600 79.600 208.400 79.700 ;
        RECT 246.000 79.600 246.800 79.700 ;
        RECT 284.400 79.600 285.200 79.700 ;
        RECT 326.000 80.300 326.800 80.400 ;
        RECT 337.200 80.300 338.000 80.400 ;
        RECT 359.600 80.300 360.400 80.400 ;
        RECT 367.600 80.300 368.400 80.400 ;
        RECT 326.000 79.700 368.400 80.300 ;
        RECT 326.000 79.600 326.800 79.700 ;
        RECT 337.200 79.600 338.000 79.700 ;
        RECT 359.600 79.600 360.400 79.700 ;
        RECT 367.600 79.600 368.400 79.700 ;
        RECT 423.600 80.300 424.400 80.400 ;
        RECT 446.000 80.300 446.800 80.400 ;
        RECT 423.600 79.700 446.800 80.300 ;
        RECT 423.600 79.600 424.400 79.700 ;
        RECT 446.000 79.600 446.800 79.700 ;
        RECT 492.400 80.300 493.200 80.400 ;
        RECT 511.600 80.300 512.400 80.400 ;
        RECT 492.400 79.700 512.400 80.300 ;
        RECT 492.400 79.600 493.200 79.700 ;
        RECT 511.600 79.600 512.400 79.700 ;
        RECT 158.000 78.300 158.800 78.400 ;
        RECT 182.000 78.300 182.800 78.400 ;
        RECT 158.000 77.700 182.800 78.300 ;
        RECT 158.000 77.600 158.800 77.700 ;
        RECT 182.000 77.600 182.800 77.700 ;
        RECT 361.200 78.300 362.000 78.400 ;
        RECT 364.400 78.300 365.200 78.400 ;
        RECT 436.400 78.300 437.200 78.400 ;
        RECT 438.000 78.300 438.800 78.400 ;
        RECT 506.800 78.300 507.600 78.400 ;
        RECT 361.200 77.700 429.100 78.300 ;
        RECT 361.200 77.600 362.000 77.700 ;
        RECT 364.400 77.600 365.200 77.700 ;
        RECT 30.000 76.300 30.800 76.400 ;
        RECT 41.200 76.300 42.000 76.400 ;
        RECT 30.000 75.700 42.000 76.300 ;
        RECT 30.000 75.600 30.800 75.700 ;
        RECT 41.200 75.600 42.000 75.700 ;
        RECT 130.800 76.300 131.600 76.400 ;
        RECT 150.000 76.300 150.800 76.400 ;
        RECT 130.800 75.700 150.800 76.300 ;
        RECT 130.800 75.600 131.600 75.700 ;
        RECT 150.000 75.600 150.800 75.700 ;
        RECT 318.000 76.300 318.800 76.400 ;
        RECT 426.800 76.300 427.600 76.400 ;
        RECT 318.000 75.700 427.600 76.300 ;
        RECT 428.500 76.300 429.100 77.700 ;
        RECT 436.400 77.700 507.600 78.300 ;
        RECT 436.400 77.600 437.200 77.700 ;
        RECT 438.000 77.600 438.800 77.700 ;
        RECT 506.800 77.600 507.600 77.700 ;
        RECT 591.600 78.300 592.400 78.400 ;
        RECT 594.800 78.300 595.600 78.400 ;
        RECT 591.600 77.700 595.600 78.300 ;
        RECT 591.600 77.600 592.400 77.700 ;
        RECT 594.800 77.600 595.600 77.700 ;
        RECT 455.600 76.300 456.400 76.400 ;
        RECT 428.500 75.700 456.400 76.300 ;
        RECT 318.000 75.600 318.800 75.700 ;
        RECT 426.800 75.600 427.600 75.700 ;
        RECT 455.600 75.600 456.400 75.700 ;
        RECT 457.200 76.300 458.000 76.400 ;
        RECT 498.800 76.300 499.600 76.400 ;
        RECT 514.800 76.300 515.600 76.400 ;
        RECT 457.200 75.700 491.500 76.300 ;
        RECT 457.200 75.600 458.000 75.700 ;
        RECT 7.600 74.300 8.400 74.400 ;
        RECT 10.800 74.300 11.600 74.400 ;
        RECT 7.600 73.700 11.600 74.300 ;
        RECT 7.600 73.600 8.400 73.700 ;
        RECT 10.800 73.600 11.600 73.700 ;
        RECT 28.400 74.300 29.200 74.400 ;
        RECT 38.000 74.300 38.800 74.400 ;
        RECT 62.000 74.300 62.800 74.400 ;
        RECT 28.400 73.700 62.800 74.300 ;
        RECT 28.400 73.600 29.200 73.700 ;
        RECT 38.000 73.600 38.800 73.700 ;
        RECT 62.000 73.600 62.800 73.700 ;
        RECT 63.600 74.300 64.400 74.400 ;
        RECT 78.000 74.300 78.800 74.400 ;
        RECT 63.600 73.700 78.800 74.300 ;
        RECT 63.600 73.600 64.400 73.700 ;
        RECT 78.000 73.600 78.800 73.700 ;
        RECT 79.600 74.300 80.400 74.400 ;
        RECT 119.600 74.300 120.400 74.400 ;
        RECT 79.600 73.700 120.400 74.300 ;
        RECT 79.600 73.600 80.400 73.700 ;
        RECT 119.600 73.600 120.400 73.700 ;
        RECT 145.200 74.300 146.000 74.400 ;
        RECT 148.400 74.300 149.200 74.400 ;
        RECT 145.200 73.700 149.200 74.300 ;
        RECT 145.200 73.600 146.000 73.700 ;
        RECT 148.400 73.600 149.200 73.700 ;
        RECT 156.400 74.300 157.200 74.400 ;
        RECT 188.400 74.300 189.200 74.400 ;
        RECT 156.400 73.700 189.200 74.300 ;
        RECT 156.400 73.600 157.200 73.700 ;
        RECT 188.400 73.600 189.200 73.700 ;
        RECT 193.200 74.300 194.000 74.400 ;
        RECT 199.600 74.300 200.400 74.400 ;
        RECT 193.200 73.700 200.400 74.300 ;
        RECT 193.200 73.600 194.000 73.700 ;
        RECT 199.600 73.600 200.400 73.700 ;
        RECT 252.400 74.300 253.200 74.400 ;
        RECT 258.800 74.300 259.600 74.400 ;
        RECT 252.400 73.700 259.600 74.300 ;
        RECT 252.400 73.600 253.200 73.700 ;
        RECT 258.800 73.600 259.600 73.700 ;
        RECT 303.600 74.300 304.400 74.400 ;
        RECT 354.800 74.300 355.600 74.400 ;
        RECT 303.600 73.700 355.600 74.300 ;
        RECT 303.600 73.600 304.400 73.700 ;
        RECT 354.800 73.600 355.600 73.700 ;
        RECT 386.800 74.300 387.600 74.400 ;
        RECT 390.000 74.300 390.800 74.400 ;
        RECT 386.800 73.700 390.800 74.300 ;
        RECT 386.800 73.600 387.600 73.700 ;
        RECT 390.000 73.600 390.800 73.700 ;
        RECT 394.800 74.300 395.600 74.400 ;
        RECT 410.800 74.300 411.600 74.400 ;
        RECT 444.400 74.300 445.200 74.400 ;
        RECT 394.800 73.700 411.600 74.300 ;
        RECT 394.800 73.600 395.600 73.700 ;
        RECT 410.800 73.600 411.600 73.700 ;
        RECT 412.500 73.700 445.200 74.300 ;
        RECT 10.800 72.300 11.600 72.400 ;
        RECT 17.200 72.300 18.000 72.400 ;
        RECT 10.800 71.700 18.000 72.300 ;
        RECT 10.800 71.600 11.600 71.700 ;
        RECT 17.200 71.600 18.000 71.700 ;
        RECT 26.800 72.300 27.600 72.400 ;
        RECT 31.600 72.300 32.400 72.400 ;
        RECT 26.800 71.700 32.400 72.300 ;
        RECT 26.800 71.600 27.600 71.700 ;
        RECT 31.600 71.600 32.400 71.700 ;
        RECT 36.400 72.300 37.200 72.400 ;
        RECT 49.200 72.300 50.000 72.400 ;
        RECT 36.400 71.700 50.000 72.300 ;
        RECT 36.400 71.600 37.200 71.700 ;
        RECT 49.200 71.600 50.000 71.700 ;
        RECT 70.000 72.300 70.800 72.400 ;
        RECT 71.600 72.300 72.400 72.400 ;
        RECT 70.000 71.700 72.400 72.300 ;
        RECT 70.000 71.600 70.800 71.700 ;
        RECT 71.600 71.600 72.400 71.700 ;
        RECT 82.800 72.300 83.600 72.400 ;
        RECT 121.200 72.300 122.000 72.400 ;
        RECT 82.800 71.700 122.000 72.300 ;
        RECT 82.800 71.600 83.600 71.700 ;
        RECT 121.200 71.600 122.000 71.700 ;
        RECT 145.200 72.300 146.000 72.400 ;
        RECT 196.400 72.300 197.200 72.400 ;
        RECT 145.200 71.700 197.200 72.300 ;
        RECT 145.200 71.600 146.000 71.700 ;
        RECT 196.400 71.600 197.200 71.700 ;
        RECT 202.800 72.300 203.600 72.400 ;
        RECT 238.000 72.300 238.800 72.400 ;
        RECT 202.800 71.700 238.800 72.300 ;
        RECT 202.800 71.600 203.600 71.700 ;
        RECT 238.000 71.600 238.800 71.700 ;
        RECT 370.800 72.300 371.600 72.400 ;
        RECT 374.000 72.300 374.800 72.400 ;
        RECT 382.000 72.300 382.800 72.400 ;
        RECT 394.800 72.300 395.600 72.400 ;
        RECT 401.200 72.300 402.000 72.400 ;
        RECT 412.500 72.300 413.100 73.700 ;
        RECT 444.400 73.600 445.200 73.700 ;
        RECT 446.000 74.300 446.800 74.400 ;
        RECT 463.600 74.300 464.400 74.400 ;
        RECT 446.000 73.700 464.400 74.300 ;
        RECT 446.000 73.600 446.800 73.700 ;
        RECT 463.600 73.600 464.400 73.700 ;
        RECT 471.600 74.300 472.400 74.400 ;
        RECT 489.200 74.300 490.000 74.400 ;
        RECT 471.600 73.700 490.000 74.300 ;
        RECT 490.900 74.300 491.500 75.700 ;
        RECT 498.800 75.700 515.600 76.300 ;
        RECT 498.800 75.600 499.600 75.700 ;
        RECT 514.800 75.600 515.600 75.700 ;
        RECT 543.600 76.300 544.400 76.400 ;
        RECT 546.800 76.300 547.600 76.400 ;
        RECT 543.600 75.700 547.600 76.300 ;
        RECT 543.600 75.600 544.400 75.700 ;
        RECT 546.800 75.600 547.600 75.700 ;
        RECT 570.800 76.300 571.600 76.400 ;
        RECT 602.800 76.300 603.600 76.400 ;
        RECT 570.800 75.700 603.600 76.300 ;
        RECT 570.800 75.600 571.600 75.700 ;
        RECT 602.800 75.600 603.600 75.700 ;
        RECT 535.600 74.300 536.400 74.400 ;
        RECT 490.900 73.700 536.400 74.300 ;
        RECT 471.600 73.600 472.400 73.700 ;
        RECT 489.200 73.600 490.000 73.700 ;
        RECT 535.600 73.600 536.400 73.700 ;
        RECT 542.000 74.300 542.800 74.400 ;
        RECT 543.600 74.300 544.400 74.400 ;
        RECT 542.000 73.700 544.400 74.300 ;
        RECT 542.000 73.600 542.800 73.700 ;
        RECT 543.600 73.600 544.400 73.700 ;
        RECT 558.000 74.300 558.800 74.400 ;
        RECT 572.400 74.300 573.200 74.400 ;
        RECT 558.000 73.700 573.200 74.300 ;
        RECT 558.000 73.600 558.800 73.700 ;
        RECT 572.400 73.600 573.200 73.700 ;
        RECT 575.600 74.300 576.400 74.400 ;
        RECT 583.600 74.300 584.400 74.400 ;
        RECT 575.600 73.700 584.400 74.300 ;
        RECT 575.600 73.600 576.400 73.700 ;
        RECT 583.600 73.600 584.400 73.700 ;
        RECT 370.800 71.700 413.100 72.300 ;
        RECT 414.000 72.300 414.800 72.400 ;
        RECT 417.200 72.300 418.000 72.400 ;
        RECT 414.000 71.700 418.000 72.300 ;
        RECT 370.800 71.600 371.600 71.700 ;
        RECT 374.000 71.600 374.800 71.700 ;
        RECT 382.000 71.600 382.800 71.700 ;
        RECT 394.800 71.600 395.600 71.700 ;
        RECT 401.200 71.600 402.000 71.700 ;
        RECT 414.000 71.600 414.800 71.700 ;
        RECT 417.200 71.600 418.000 71.700 ;
        RECT 420.400 72.300 421.200 72.400 ;
        RECT 425.200 72.300 426.000 72.400 ;
        RECT 420.400 71.700 426.000 72.300 ;
        RECT 420.400 71.600 421.200 71.700 ;
        RECT 425.200 71.600 426.000 71.700 ;
        RECT 444.400 72.300 445.200 72.400 ;
        RECT 446.000 72.300 446.800 72.400 ;
        RECT 452.400 72.300 453.200 72.400 ;
        RECT 444.400 71.700 453.200 72.300 ;
        RECT 444.400 71.600 445.200 71.700 ;
        RECT 446.000 71.600 446.800 71.700 ;
        RECT 452.400 71.600 453.200 71.700 ;
        RECT 470.000 72.300 470.800 72.400 ;
        RECT 484.400 72.300 485.200 72.400 ;
        RECT 470.000 71.700 485.200 72.300 ;
        RECT 470.000 71.600 470.800 71.700 ;
        RECT 484.400 71.600 485.200 71.700 ;
        RECT 505.200 72.300 506.000 72.400 ;
        RECT 526.000 72.300 526.800 72.400 ;
        RECT 505.200 71.700 526.800 72.300 ;
        RECT 505.200 71.600 506.000 71.700 ;
        RECT 526.000 71.600 526.800 71.700 ;
        RECT 561.200 72.300 562.000 72.400 ;
        RECT 564.400 72.300 565.200 72.400 ;
        RECT 596.400 72.300 597.200 72.400 ;
        RECT 561.200 71.700 597.200 72.300 ;
        RECT 561.200 71.600 562.000 71.700 ;
        RECT 564.400 71.600 565.200 71.700 ;
        RECT 596.400 71.600 597.200 71.700 ;
        RECT 4.400 70.300 5.200 70.400 ;
        RECT 6.000 70.300 6.800 70.400 ;
        RECT 4.400 69.700 6.800 70.300 ;
        RECT 4.400 69.600 5.200 69.700 ;
        RECT 6.000 69.600 6.800 69.700 ;
        RECT 25.200 70.300 26.000 70.400 ;
        RECT 33.200 70.300 34.000 70.400 ;
        RECT 25.200 69.700 34.000 70.300 ;
        RECT 25.200 69.600 26.000 69.700 ;
        RECT 33.200 69.600 34.000 69.700 ;
        RECT 41.200 70.300 42.000 70.400 ;
        RECT 46.000 70.300 46.800 70.400 ;
        RECT 52.400 70.300 53.200 70.400 ;
        RECT 65.200 70.300 66.000 70.400 ;
        RECT 71.600 70.300 72.400 70.400 ;
        RECT 90.800 70.300 91.600 70.400 ;
        RECT 41.200 69.700 91.600 70.300 ;
        RECT 41.200 69.600 42.000 69.700 ;
        RECT 46.000 69.600 46.800 69.700 ;
        RECT 52.400 69.600 53.200 69.700 ;
        RECT 65.200 69.600 66.000 69.700 ;
        RECT 71.600 69.600 72.400 69.700 ;
        RECT 90.800 69.600 91.600 69.700 ;
        RECT 98.800 70.300 99.600 70.400 ;
        RECT 134.000 70.300 134.800 70.400 ;
        RECT 98.800 69.700 134.800 70.300 ;
        RECT 98.800 69.600 99.600 69.700 ;
        RECT 134.000 69.600 134.800 69.700 ;
        RECT 146.800 70.300 147.600 70.400 ;
        RECT 162.800 70.300 163.600 70.400 ;
        RECT 146.800 69.700 163.600 70.300 ;
        RECT 146.800 69.600 147.600 69.700 ;
        RECT 162.800 69.600 163.600 69.700 ;
        RECT 182.000 70.300 182.800 70.400 ;
        RECT 191.600 70.300 192.400 70.400 ;
        RECT 182.000 69.700 192.400 70.300 ;
        RECT 182.000 69.600 182.800 69.700 ;
        RECT 191.600 69.600 192.400 69.700 ;
        RECT 201.200 70.300 202.000 70.400 ;
        RECT 207.600 70.300 208.400 70.400 ;
        RECT 201.200 69.700 208.400 70.300 ;
        RECT 201.200 69.600 202.000 69.700 ;
        RECT 207.600 69.600 208.400 69.700 ;
        RECT 338.800 70.300 339.600 70.400 ;
        RECT 358.000 70.300 358.800 70.400 ;
        RECT 366.000 70.300 366.800 70.400 ;
        RECT 375.600 70.300 376.400 70.400 ;
        RECT 338.800 69.700 376.400 70.300 ;
        RECT 338.800 69.600 339.600 69.700 ;
        RECT 358.000 69.600 358.800 69.700 ;
        RECT 366.000 69.600 366.800 69.700 ;
        RECT 375.600 69.600 376.400 69.700 ;
        RECT 410.800 69.600 411.600 70.400 ;
        RECT 423.600 70.300 424.400 70.400 ;
        RECT 426.800 70.300 427.600 70.400 ;
        RECT 423.600 69.700 427.600 70.300 ;
        RECT 423.600 69.600 424.400 69.700 ;
        RECT 426.800 69.600 427.600 69.700 ;
        RECT 439.600 70.300 440.400 70.400 ;
        RECT 474.800 70.300 475.600 70.400 ;
        RECT 439.600 69.700 475.600 70.300 ;
        RECT 439.600 69.600 440.400 69.700 ;
        RECT 474.800 69.600 475.600 69.700 ;
        RECT 479.600 70.300 480.400 70.400 ;
        RECT 492.400 70.300 493.200 70.400 ;
        RECT 479.600 69.700 493.200 70.300 ;
        RECT 479.600 69.600 480.400 69.700 ;
        RECT 492.400 69.600 493.200 69.700 ;
        RECT 502.000 70.300 502.800 70.400 ;
        RECT 505.200 70.300 506.000 70.400 ;
        RECT 502.000 69.700 506.000 70.300 ;
        RECT 502.000 69.600 502.800 69.700 ;
        RECT 505.200 69.600 506.000 69.700 ;
        RECT 508.400 70.300 509.200 70.400 ;
        RECT 535.600 70.300 536.400 70.400 ;
        RECT 508.400 69.700 536.400 70.300 ;
        RECT 508.400 69.600 509.200 69.700 ;
        RECT 535.600 69.600 536.400 69.700 ;
        RECT 554.800 70.300 555.600 70.400 ;
        RECT 561.200 70.300 562.000 70.400 ;
        RECT 554.800 69.700 562.000 70.300 ;
        RECT 554.800 69.600 555.600 69.700 ;
        RECT 561.200 69.600 562.000 69.700 ;
        RECT 570.800 70.300 571.600 70.400 ;
        RECT 575.600 70.300 576.400 70.400 ;
        RECT 570.800 69.700 576.400 70.300 ;
        RECT 570.800 69.600 571.600 69.700 ;
        RECT 575.600 69.600 576.400 69.700 ;
        RECT 22.000 68.300 22.800 68.400 ;
        RECT 46.000 68.300 46.800 68.400 ;
        RECT 22.000 67.700 46.800 68.300 ;
        RECT 22.000 67.600 22.800 67.700 ;
        RECT 46.000 67.600 46.800 67.700 ;
        RECT 71.600 67.600 72.400 68.400 ;
        RECT 74.800 68.300 75.600 68.400 ;
        RECT 92.400 68.300 93.200 68.400 ;
        RECT 74.800 67.700 93.200 68.300 ;
        RECT 74.800 67.600 75.600 67.700 ;
        RECT 92.400 67.600 93.200 67.700 ;
        RECT 100.400 68.300 101.200 68.400 ;
        RECT 118.000 68.300 118.800 68.400 ;
        RECT 100.400 67.700 118.800 68.300 ;
        RECT 100.400 67.600 101.200 67.700 ;
        RECT 118.000 67.600 118.800 67.700 ;
        RECT 140.400 68.300 141.200 68.400 ;
        RECT 164.400 68.300 165.200 68.400 ;
        RECT 177.200 68.300 178.000 68.400 ;
        RECT 140.400 67.700 178.000 68.300 ;
        RECT 140.400 67.600 141.200 67.700 ;
        RECT 164.400 67.600 165.200 67.700 ;
        RECT 177.200 67.600 178.000 67.700 ;
        RECT 186.800 68.300 187.600 68.400 ;
        RECT 193.200 68.300 194.000 68.400 ;
        RECT 186.800 67.700 194.000 68.300 ;
        RECT 186.800 67.600 187.600 67.700 ;
        RECT 193.200 67.600 194.000 67.700 ;
        RECT 201.200 68.300 202.000 68.400 ;
        RECT 217.200 68.300 218.000 68.400 ;
        RECT 201.200 67.700 218.000 68.300 ;
        RECT 201.200 67.600 202.000 67.700 ;
        RECT 217.200 67.600 218.000 67.700 ;
        RECT 257.200 68.300 258.000 68.400 ;
        RECT 278.000 68.300 278.800 68.400 ;
        RECT 257.200 67.700 278.800 68.300 ;
        RECT 257.200 67.600 258.000 67.700 ;
        RECT 278.000 67.600 278.800 67.700 ;
        RECT 289.200 68.300 290.000 68.400 ;
        RECT 292.400 68.300 293.200 68.400 ;
        RECT 289.200 67.700 293.200 68.300 ;
        RECT 289.200 67.600 290.000 67.700 ;
        RECT 292.400 67.600 293.200 67.700 ;
        RECT 343.600 68.300 344.400 68.400 ;
        RECT 353.200 68.300 354.000 68.400 ;
        RECT 343.600 67.700 354.000 68.300 ;
        RECT 343.600 67.600 344.400 67.700 ;
        RECT 353.200 67.600 354.000 67.700 ;
        RECT 356.400 68.300 357.200 68.400 ;
        RECT 361.200 68.300 362.000 68.400 ;
        RECT 356.400 67.700 362.000 68.300 ;
        RECT 356.400 67.600 357.200 67.700 ;
        RECT 361.200 67.600 362.000 67.700 ;
        RECT 407.600 68.300 408.400 68.400 ;
        RECT 415.600 68.300 416.400 68.400 ;
        RECT 422.000 68.300 422.800 68.400 ;
        RECT 407.600 67.700 422.800 68.300 ;
        RECT 407.600 67.600 408.400 67.700 ;
        RECT 415.600 67.600 416.400 67.700 ;
        RECT 422.000 67.600 422.800 67.700 ;
        RECT 425.200 68.300 426.000 68.400 ;
        RECT 428.400 68.300 429.200 68.400 ;
        RECT 425.200 67.700 429.200 68.300 ;
        RECT 425.200 67.600 426.000 67.700 ;
        RECT 428.400 67.600 429.200 67.700 ;
        RECT 447.600 68.300 448.400 68.400 ;
        RECT 482.800 68.300 483.600 68.400 ;
        RECT 447.600 67.700 483.600 68.300 ;
        RECT 447.600 67.600 448.400 67.700 ;
        RECT 482.800 67.600 483.600 67.700 ;
        RECT 489.200 68.300 490.000 68.400 ;
        RECT 500.400 68.300 501.200 68.400 ;
        RECT 489.200 67.700 501.200 68.300 ;
        RECT 489.200 67.600 490.000 67.700 ;
        RECT 500.400 67.600 501.200 67.700 ;
        RECT 503.600 68.300 504.400 68.400 ;
        RECT 508.400 68.300 509.200 68.400 ;
        RECT 503.600 67.700 509.200 68.300 ;
        RECT 503.600 67.600 504.400 67.700 ;
        RECT 508.400 67.600 509.200 67.700 ;
        RECT 516.400 68.300 517.200 68.400 ;
        RECT 540.400 68.300 541.200 68.400 ;
        RECT 516.400 67.700 541.200 68.300 ;
        RECT 516.400 67.600 517.200 67.700 ;
        RECT 540.400 67.600 541.200 67.700 ;
        RECT 543.600 68.300 544.400 68.400 ;
        RECT 548.400 68.300 549.200 68.400 ;
        RECT 543.600 67.700 549.200 68.300 ;
        RECT 543.600 67.600 544.400 67.700 ;
        RECT 548.400 67.600 549.200 67.700 ;
        RECT 586.800 68.300 587.600 68.400 ;
        RECT 598.000 68.300 598.800 68.400 ;
        RECT 586.800 67.700 598.800 68.300 ;
        RECT 586.800 67.600 587.600 67.700 ;
        RECT 598.000 67.600 598.800 67.700 ;
        RECT 601.200 68.300 602.000 68.400 ;
        RECT 606.000 68.300 606.800 68.400 ;
        RECT 601.200 67.700 606.800 68.300 ;
        RECT 601.200 67.600 602.000 67.700 ;
        RECT 606.000 67.600 606.800 67.700 ;
        RECT 17.200 66.300 18.000 66.400 ;
        RECT 33.200 66.300 34.000 66.400 ;
        RECT 17.200 65.700 34.000 66.300 ;
        RECT 17.200 65.600 18.000 65.700 ;
        RECT 33.200 65.600 34.000 65.700 ;
        RECT 36.400 66.300 37.200 66.400 ;
        RECT 42.800 66.300 43.600 66.400 ;
        RECT 63.600 66.300 64.400 66.400 ;
        RECT 70.000 66.300 70.800 66.400 ;
        RECT 36.400 65.700 70.800 66.300 ;
        RECT 36.400 65.600 37.200 65.700 ;
        RECT 42.800 65.600 43.600 65.700 ;
        RECT 63.600 65.600 64.400 65.700 ;
        RECT 70.000 65.600 70.800 65.700 ;
        RECT 79.600 66.300 80.400 66.400 ;
        RECT 86.000 66.300 86.800 66.400 ;
        RECT 79.600 65.700 86.800 66.300 ;
        RECT 79.600 65.600 80.400 65.700 ;
        RECT 86.000 65.600 86.800 65.700 ;
        RECT 92.400 66.300 93.200 66.400 ;
        RECT 102.000 66.300 102.800 66.400 ;
        RECT 108.400 66.300 109.200 66.400 ;
        RECT 92.400 65.700 109.200 66.300 ;
        RECT 92.400 65.600 93.200 65.700 ;
        RECT 102.000 65.600 102.800 65.700 ;
        RECT 108.400 65.600 109.200 65.700 ;
        RECT 196.400 66.300 197.200 66.400 ;
        RECT 220.400 66.300 221.200 66.400 ;
        RECT 196.400 65.700 221.200 66.300 ;
        RECT 196.400 65.600 197.200 65.700 ;
        RECT 220.400 65.600 221.200 65.700 ;
        RECT 266.800 66.300 267.600 66.400 ;
        RECT 274.800 66.300 275.600 66.400 ;
        RECT 319.600 66.300 320.400 66.400 ;
        RECT 266.800 65.700 320.400 66.300 ;
        RECT 266.800 65.600 267.600 65.700 ;
        RECT 274.800 65.600 275.600 65.700 ;
        RECT 319.600 65.600 320.400 65.700 ;
        RECT 322.800 66.300 323.600 66.400 ;
        RECT 362.800 66.300 363.600 66.400 ;
        RECT 322.800 65.700 363.600 66.300 ;
        RECT 322.800 65.600 323.600 65.700 ;
        RECT 362.800 65.600 363.600 65.700 ;
        RECT 367.600 66.300 368.400 66.400 ;
        RECT 372.400 66.300 373.200 66.400 ;
        RECT 367.600 65.700 373.200 66.300 ;
        RECT 367.600 65.600 368.400 65.700 ;
        RECT 372.400 65.600 373.200 65.700 ;
        RECT 412.400 66.300 413.200 66.400 ;
        RECT 423.600 66.300 424.400 66.400 ;
        RECT 454.000 66.300 454.800 66.400 ;
        RECT 466.800 66.300 467.600 66.400 ;
        RECT 412.400 65.700 467.600 66.300 ;
        RECT 412.400 65.600 413.200 65.700 ;
        RECT 423.600 65.600 424.400 65.700 ;
        RECT 454.000 65.600 454.800 65.700 ;
        RECT 466.800 65.600 467.600 65.700 ;
        RECT 513.200 66.300 514.000 66.400 ;
        RECT 545.200 66.300 546.000 66.400 ;
        RECT 513.200 65.700 546.000 66.300 ;
        RECT 513.200 65.600 514.000 65.700 ;
        RECT 545.200 65.600 546.000 65.700 ;
        RECT 2.800 64.300 3.600 64.400 ;
        RECT 14.000 64.300 14.800 64.400 ;
        RECT 34.800 64.300 35.600 64.400 ;
        RECT 2.800 63.700 35.600 64.300 ;
        RECT 2.800 63.600 3.600 63.700 ;
        RECT 14.000 63.600 14.800 63.700 ;
        RECT 34.800 63.600 35.600 63.700 ;
        RECT 44.400 64.300 45.200 64.400 ;
        RECT 46.000 64.300 46.800 64.400 ;
        RECT 44.400 63.700 46.800 64.300 ;
        RECT 44.400 63.600 45.200 63.700 ;
        RECT 46.000 63.600 46.800 63.700 ;
        RECT 68.400 64.300 69.200 64.400 ;
        RECT 98.800 64.300 99.600 64.400 ;
        RECT 68.400 63.700 99.600 64.300 ;
        RECT 68.400 63.600 69.200 63.700 ;
        RECT 98.800 63.600 99.600 63.700 ;
        RECT 284.400 64.300 285.200 64.400 ;
        RECT 310.000 64.300 310.800 64.400 ;
        RECT 284.400 63.700 310.800 64.300 ;
        RECT 284.400 63.600 285.200 63.700 ;
        RECT 310.000 63.600 310.800 63.700 ;
        RECT 338.800 64.300 339.600 64.400 ;
        RECT 370.800 64.300 371.600 64.400 ;
        RECT 393.200 64.300 394.000 64.400 ;
        RECT 409.200 64.300 410.000 64.400 ;
        RECT 417.200 64.300 418.000 64.400 ;
        RECT 338.800 63.700 418.000 64.300 ;
        RECT 338.800 63.600 339.600 63.700 ;
        RECT 370.800 63.600 371.600 63.700 ;
        RECT 393.200 63.600 394.000 63.700 ;
        RECT 409.200 63.600 410.000 63.700 ;
        RECT 417.200 63.600 418.000 63.700 ;
        RECT 441.200 64.300 442.000 64.400 ;
        RECT 513.200 64.300 514.000 64.400 ;
        RECT 441.200 63.700 514.000 64.300 ;
        RECT 441.200 63.600 442.000 63.700 ;
        RECT 513.200 63.600 514.000 63.700 ;
        RECT 559.600 64.300 560.400 64.400 ;
        RECT 580.400 64.300 581.200 64.400 ;
        RECT 559.600 63.700 581.200 64.300 ;
        RECT 559.600 63.600 560.400 63.700 ;
        RECT 580.400 63.600 581.200 63.700 ;
        RECT 9.200 62.300 10.000 62.400 ;
        RECT 14.000 62.300 14.800 62.400 ;
        RECT 9.200 61.700 14.800 62.300 ;
        RECT 9.200 61.600 10.000 61.700 ;
        RECT 14.000 61.600 14.800 61.700 ;
        RECT 15.600 62.300 16.400 62.400 ;
        RECT 36.400 62.300 37.200 62.400 ;
        RECT 15.600 61.700 37.200 62.300 ;
        RECT 15.600 61.600 16.400 61.700 ;
        RECT 36.400 61.600 37.200 61.700 ;
        RECT 74.800 62.300 75.600 62.400 ;
        RECT 89.200 62.300 90.000 62.400 ;
        RECT 74.800 61.700 90.000 62.300 ;
        RECT 74.800 61.600 75.600 61.700 ;
        RECT 89.200 61.600 90.000 61.700 ;
        RECT 174.000 62.300 174.800 62.400 ;
        RECT 252.400 62.300 253.200 62.400 ;
        RECT 174.000 61.700 253.200 62.300 ;
        RECT 174.000 61.600 174.800 61.700 ;
        RECT 252.400 61.600 253.200 61.700 ;
        RECT 370.800 62.300 371.600 62.400 ;
        RECT 377.200 62.300 378.000 62.400 ;
        RECT 370.800 61.700 378.000 62.300 ;
        RECT 370.800 61.600 371.600 61.700 ;
        RECT 377.200 61.600 378.000 61.700 ;
        RECT 399.600 62.300 400.400 62.400 ;
        RECT 401.200 62.300 402.000 62.400 ;
        RECT 399.600 61.700 402.000 62.300 ;
        RECT 399.600 61.600 400.400 61.700 ;
        RECT 401.200 61.600 402.000 61.700 ;
        RECT 418.800 62.300 419.600 62.400 ;
        RECT 473.200 62.300 474.000 62.400 ;
        RECT 484.400 62.300 485.200 62.400 ;
        RECT 418.800 61.700 485.200 62.300 ;
        RECT 418.800 61.600 419.600 61.700 ;
        RECT 473.200 61.600 474.000 61.700 ;
        RECT 484.400 61.600 485.200 61.700 ;
        RECT 530.800 62.300 531.600 62.400 ;
        RECT 556.400 62.300 557.200 62.400 ;
        RECT 530.800 61.700 557.200 62.300 ;
        RECT 530.800 61.600 531.600 61.700 ;
        RECT 556.400 61.600 557.200 61.700 ;
        RECT 12.400 60.300 13.200 60.400 ;
        RECT 17.200 60.300 18.000 60.400 ;
        RECT 12.400 59.700 18.000 60.300 ;
        RECT 12.400 59.600 13.200 59.700 ;
        RECT 17.200 59.600 18.000 59.700 ;
        RECT 23.600 60.300 24.400 60.400 ;
        RECT 63.600 60.300 64.400 60.400 ;
        RECT 84.400 60.300 85.200 60.400 ;
        RECT 23.600 59.700 85.200 60.300 ;
        RECT 23.600 59.600 24.400 59.700 ;
        RECT 63.600 59.600 64.400 59.700 ;
        RECT 84.400 59.600 85.200 59.700 ;
        RECT 162.800 60.300 163.600 60.400 ;
        RECT 178.800 60.300 179.600 60.400 ;
        RECT 162.800 59.700 179.600 60.300 ;
        RECT 162.800 59.600 163.600 59.700 ;
        RECT 178.800 59.600 179.600 59.700 ;
        RECT 353.200 60.300 354.000 60.400 ;
        RECT 390.000 60.300 390.800 60.400 ;
        RECT 353.200 59.700 390.800 60.300 ;
        RECT 353.200 59.600 354.000 59.700 ;
        RECT 390.000 59.600 390.800 59.700 ;
        RECT 404.400 60.300 405.200 60.400 ;
        RECT 420.400 60.300 421.200 60.400 ;
        RECT 404.400 59.700 421.200 60.300 ;
        RECT 404.400 59.600 405.200 59.700 ;
        RECT 420.400 59.600 421.200 59.700 ;
        RECT 422.000 60.300 422.800 60.400 ;
        RECT 434.800 60.300 435.600 60.400 ;
        RECT 422.000 59.700 435.600 60.300 ;
        RECT 422.000 59.600 422.800 59.700 ;
        RECT 434.800 59.600 435.600 59.700 ;
        RECT 449.200 60.300 450.000 60.400 ;
        RECT 479.600 60.300 480.400 60.400 ;
        RECT 449.200 59.700 480.400 60.300 ;
        RECT 449.200 59.600 450.000 59.700 ;
        RECT 479.600 59.600 480.400 59.700 ;
        RECT 527.600 60.300 528.400 60.400 ;
        RECT 542.000 60.300 542.800 60.400 ;
        RECT 577.200 60.300 578.000 60.400 ;
        RECT 527.600 59.700 578.000 60.300 ;
        RECT 527.600 59.600 528.400 59.700 ;
        RECT 542.000 59.600 542.800 59.700 ;
        RECT 577.200 59.600 578.000 59.700 ;
        RECT 598.000 60.300 598.800 60.400 ;
        RECT 602.800 60.300 603.600 60.400 ;
        RECT 598.000 59.700 603.600 60.300 ;
        RECT 598.000 59.600 598.800 59.700 ;
        RECT 602.800 59.600 603.600 59.700 ;
        RECT 92.400 58.300 93.200 58.400 ;
        RECT 105.200 58.300 106.000 58.400 ;
        RECT 92.400 57.700 106.000 58.300 ;
        RECT 92.400 57.600 93.200 57.700 ;
        RECT 105.200 57.600 106.000 57.700 ;
        RECT 206.000 58.300 206.800 58.400 ;
        RECT 212.400 58.300 213.200 58.400 ;
        RECT 206.000 57.700 213.200 58.300 ;
        RECT 206.000 57.600 206.800 57.700 ;
        RECT 212.400 57.600 213.200 57.700 ;
        RECT 222.000 58.300 222.800 58.400 ;
        RECT 246.000 58.300 246.800 58.400 ;
        RECT 222.000 57.700 246.800 58.300 ;
        RECT 222.000 57.600 222.800 57.700 ;
        RECT 246.000 57.600 246.800 57.700 ;
        RECT 311.600 58.300 312.400 58.400 ;
        RECT 319.600 58.300 320.400 58.400 ;
        RECT 311.600 57.700 320.400 58.300 ;
        RECT 311.600 57.600 312.400 57.700 ;
        RECT 319.600 57.600 320.400 57.700 ;
        RECT 326.000 58.300 326.800 58.400 ;
        RECT 342.000 58.300 342.800 58.400 ;
        RECT 354.800 58.300 355.600 58.400 ;
        RECT 362.800 58.300 363.600 58.400 ;
        RECT 326.000 57.700 363.600 58.300 ;
        RECT 326.000 57.600 326.800 57.700 ;
        RECT 342.000 57.600 342.800 57.700 ;
        RECT 354.800 57.600 355.600 57.700 ;
        RECT 362.800 57.600 363.600 57.700 ;
        RECT 367.600 58.300 368.400 58.400 ;
        RECT 388.400 58.300 389.200 58.400 ;
        RECT 367.600 57.700 389.200 58.300 ;
        RECT 367.600 57.600 368.400 57.700 ;
        RECT 388.400 57.600 389.200 57.700 ;
        RECT 434.800 58.300 435.600 58.400 ;
        RECT 439.600 58.300 440.400 58.400 ;
        RECT 434.800 57.700 440.400 58.300 ;
        RECT 434.800 57.600 435.600 57.700 ;
        RECT 439.600 57.600 440.400 57.700 ;
        RECT 516.400 58.300 517.200 58.400 ;
        RECT 538.800 58.300 539.600 58.400 ;
        RECT 516.400 57.700 539.600 58.300 ;
        RECT 516.400 57.600 517.200 57.700 ;
        RECT 538.800 57.600 539.600 57.700 ;
        RECT 567.600 58.300 568.400 58.400 ;
        RECT 578.800 58.300 579.600 58.400 ;
        RECT 567.600 57.700 579.600 58.300 ;
        RECT 567.600 57.600 568.400 57.700 ;
        RECT 578.800 57.600 579.600 57.700 ;
        RECT 17.200 56.300 18.000 56.400 ;
        RECT 49.200 56.300 50.000 56.400 ;
        RECT 17.200 55.700 50.000 56.300 ;
        RECT 17.200 55.600 18.000 55.700 ;
        RECT 49.200 55.600 50.000 55.700 ;
        RECT 55.600 56.300 56.400 56.400 ;
        RECT 60.400 56.300 61.200 56.400 ;
        RECT 111.600 56.300 112.400 56.400 ;
        RECT 55.600 55.700 112.400 56.300 ;
        RECT 55.600 55.600 56.400 55.700 ;
        RECT 60.400 55.600 61.200 55.700 ;
        RECT 111.600 55.600 112.400 55.700 ;
        RECT 119.600 56.300 120.400 56.400 ;
        RECT 140.400 56.300 141.200 56.400 ;
        RECT 145.200 56.300 146.000 56.400 ;
        RECT 119.600 55.700 146.000 56.300 ;
        RECT 119.600 55.600 120.400 55.700 ;
        RECT 140.400 55.600 141.200 55.700 ;
        RECT 145.200 55.600 146.000 55.700 ;
        RECT 146.800 56.300 147.600 56.400 ;
        RECT 154.800 56.300 155.600 56.400 ;
        RECT 146.800 55.700 155.600 56.300 ;
        RECT 146.800 55.600 147.600 55.700 ;
        RECT 154.800 55.600 155.600 55.700 ;
        RECT 193.200 56.300 194.000 56.400 ;
        RECT 220.400 56.300 221.200 56.400 ;
        RECT 193.200 55.700 221.200 56.300 ;
        RECT 193.200 55.600 194.000 55.700 ;
        RECT 220.400 55.600 221.200 55.700 ;
        RECT 231.600 56.300 232.400 56.400 ;
        RECT 236.400 56.300 237.200 56.400 ;
        RECT 231.600 55.700 237.200 56.300 ;
        RECT 231.600 55.600 232.400 55.700 ;
        RECT 236.400 55.600 237.200 55.700 ;
        RECT 241.200 56.300 242.000 56.400 ;
        RECT 274.800 56.300 275.600 56.400 ;
        RECT 241.200 55.700 275.600 56.300 ;
        RECT 241.200 55.600 242.000 55.700 ;
        RECT 274.800 55.600 275.600 55.700 ;
        RECT 361.200 56.300 362.000 56.400 ;
        RECT 369.200 56.300 370.000 56.400 ;
        RECT 361.200 55.700 370.000 56.300 ;
        RECT 361.200 55.600 362.000 55.700 ;
        RECT 369.200 55.600 370.000 55.700 ;
        RECT 382.000 56.300 382.800 56.400 ;
        RECT 385.200 56.300 386.000 56.400 ;
        RECT 382.000 55.700 386.000 56.300 ;
        RECT 382.000 55.600 382.800 55.700 ;
        RECT 385.200 55.600 386.000 55.700 ;
        RECT 388.400 56.300 389.200 56.400 ;
        RECT 409.200 56.300 410.000 56.400 ;
        RECT 388.400 55.700 410.000 56.300 ;
        RECT 388.400 55.600 389.200 55.700 ;
        RECT 409.200 55.600 410.000 55.700 ;
        RECT 426.800 56.300 427.600 56.400 ;
        RECT 436.400 56.300 437.200 56.400 ;
        RECT 444.400 56.300 445.200 56.400 ;
        RECT 426.800 55.700 445.200 56.300 ;
        RECT 426.800 55.600 427.600 55.700 ;
        RECT 436.400 55.600 437.200 55.700 ;
        RECT 444.400 55.600 445.200 55.700 ;
        RECT 446.000 56.300 446.800 56.400 ;
        RECT 452.400 56.300 453.200 56.400 ;
        RECT 446.000 55.700 453.200 56.300 ;
        RECT 446.000 55.600 446.800 55.700 ;
        RECT 452.400 55.600 453.200 55.700 ;
        RECT 455.600 56.300 456.400 56.400 ;
        RECT 465.200 56.300 466.000 56.400 ;
        RECT 455.600 55.700 466.000 56.300 ;
        RECT 455.600 55.600 456.400 55.700 ;
        RECT 465.200 55.600 466.000 55.700 ;
        RECT 471.600 56.300 472.400 56.400 ;
        RECT 476.400 56.300 477.200 56.400 ;
        RECT 479.600 56.300 480.400 56.400 ;
        RECT 471.600 55.700 480.400 56.300 ;
        RECT 471.600 55.600 472.400 55.700 ;
        RECT 476.400 55.600 477.200 55.700 ;
        RECT 479.600 55.600 480.400 55.700 ;
        RECT 527.600 56.300 528.400 56.400 ;
        RECT 535.600 56.300 536.400 56.400 ;
        RECT 543.600 56.300 544.400 56.400 ;
        RECT 527.600 55.700 544.400 56.300 ;
        RECT 527.600 55.600 528.400 55.700 ;
        RECT 535.600 55.600 536.400 55.700 ;
        RECT 543.600 55.600 544.400 55.700 ;
        RECT 46.000 54.300 46.800 54.400 ;
        RECT 74.800 54.300 75.600 54.400 ;
        RECT 46.000 53.700 75.600 54.300 ;
        RECT 46.000 53.600 46.800 53.700 ;
        RECT 74.800 53.600 75.600 53.700 ;
        RECT 76.400 54.300 77.200 54.400 ;
        RECT 82.800 54.300 83.600 54.400 ;
        RECT 76.400 53.700 83.600 54.300 ;
        RECT 76.400 53.600 77.200 53.700 ;
        RECT 82.800 53.600 83.600 53.700 ;
        RECT 86.000 54.300 86.800 54.400 ;
        RECT 95.600 54.300 96.400 54.400 ;
        RECT 86.000 53.700 96.400 54.300 ;
        RECT 86.000 53.600 86.800 53.700 ;
        RECT 95.600 53.600 96.400 53.700 ;
        RECT 111.600 54.300 112.400 54.400 ;
        RECT 159.600 54.300 160.400 54.400 ;
        RECT 166.000 54.300 166.800 54.400 ;
        RECT 111.600 53.700 166.800 54.300 ;
        RECT 111.600 53.600 112.400 53.700 ;
        RECT 159.600 53.600 160.400 53.700 ;
        RECT 166.000 53.600 166.800 53.700 ;
        RECT 169.200 54.300 170.000 54.400 ;
        RECT 178.800 54.300 179.600 54.400 ;
        RECT 196.400 54.300 197.200 54.400 ;
        RECT 169.200 53.700 197.200 54.300 ;
        RECT 169.200 53.600 170.000 53.700 ;
        RECT 178.800 53.600 179.600 53.700 ;
        RECT 196.400 53.600 197.200 53.700 ;
        RECT 215.600 53.600 216.400 54.400 ;
        RECT 218.800 54.300 219.600 54.400 ;
        RECT 223.600 54.300 224.400 54.400 ;
        RECT 228.400 54.300 229.200 54.400 ;
        RECT 238.000 54.300 238.800 54.400 ;
        RECT 218.800 53.700 238.800 54.300 ;
        RECT 218.800 53.600 219.600 53.700 ;
        RECT 223.600 53.600 224.400 53.700 ;
        RECT 228.400 53.600 229.200 53.700 ;
        RECT 238.000 53.600 238.800 53.700 ;
        RECT 278.000 54.300 278.800 54.400 ;
        RECT 289.200 54.300 290.000 54.400 ;
        RECT 278.000 53.700 290.000 54.300 ;
        RECT 278.000 53.600 278.800 53.700 ;
        RECT 289.200 53.600 290.000 53.700 ;
        RECT 308.400 54.300 309.200 54.400 ;
        RECT 346.800 54.300 347.600 54.400 ;
        RECT 308.400 53.700 347.600 54.300 ;
        RECT 308.400 53.600 309.200 53.700 ;
        RECT 346.800 53.600 347.600 53.700 ;
        RECT 356.400 54.300 357.200 54.400 ;
        RECT 359.600 54.300 360.400 54.400 ;
        RECT 378.800 54.300 379.600 54.400 ;
        RECT 356.400 53.700 379.600 54.300 ;
        RECT 356.400 53.600 357.200 53.700 ;
        RECT 359.600 53.600 360.400 53.700 ;
        RECT 378.800 53.600 379.600 53.700 ;
        RECT 385.200 54.300 386.000 54.400 ;
        RECT 394.800 54.300 395.600 54.400 ;
        RECT 385.200 53.700 395.600 54.300 ;
        RECT 385.200 53.600 386.000 53.700 ;
        RECT 394.800 53.600 395.600 53.700 ;
        RECT 414.000 54.300 414.800 54.400 ;
        RECT 439.600 54.300 440.400 54.400 ;
        RECT 414.000 53.700 440.400 54.300 ;
        RECT 414.000 53.600 414.800 53.700 ;
        RECT 439.600 53.600 440.400 53.700 ;
        RECT 441.200 54.300 442.000 54.400 ;
        RECT 450.800 54.300 451.600 54.400 ;
        RECT 494.000 54.300 494.800 54.400 ;
        RECT 516.400 54.300 517.200 54.400 ;
        RECT 530.800 54.300 531.600 54.400 ;
        RECT 441.200 53.700 531.600 54.300 ;
        RECT 441.200 53.600 442.000 53.700 ;
        RECT 450.800 53.600 451.600 53.700 ;
        RECT 494.000 53.600 494.800 53.700 ;
        RECT 516.400 53.600 517.200 53.700 ;
        RECT 530.800 53.600 531.600 53.700 ;
        RECT 532.400 54.300 533.200 54.400 ;
        RECT 554.800 54.300 555.600 54.400 ;
        RECT 532.400 53.700 555.600 54.300 ;
        RECT 532.400 53.600 533.200 53.700 ;
        RECT 554.800 53.600 555.600 53.700 ;
        RECT 71.600 52.300 72.400 52.400 ;
        RECT 94.000 52.300 94.800 52.400 ;
        RECT 71.600 51.700 94.800 52.300 ;
        RECT 71.600 51.600 72.400 51.700 ;
        RECT 94.000 51.600 94.800 51.700 ;
        RECT 135.600 52.300 136.400 52.400 ;
        RECT 146.800 52.300 147.600 52.400 ;
        RECT 135.600 51.700 147.600 52.300 ;
        RECT 135.600 51.600 136.400 51.700 ;
        RECT 146.800 51.600 147.600 51.700 ;
        RECT 204.400 52.300 205.200 52.400 ;
        RECT 246.000 52.300 246.800 52.400 ;
        RECT 204.400 51.700 246.800 52.300 ;
        RECT 204.400 51.600 205.200 51.700 ;
        RECT 246.000 51.600 246.800 51.700 ;
        RECT 270.000 52.300 270.800 52.400 ;
        RECT 279.600 52.300 280.400 52.400 ;
        RECT 270.000 51.700 280.400 52.300 ;
        RECT 270.000 51.600 270.800 51.700 ;
        RECT 279.600 51.600 280.400 51.700 ;
        RECT 348.400 52.300 349.200 52.400 ;
        RECT 361.200 52.300 362.000 52.400 ;
        RECT 364.400 52.300 365.200 52.400 ;
        RECT 348.400 51.700 365.200 52.300 ;
        RECT 348.400 51.600 349.200 51.700 ;
        RECT 361.200 51.600 362.000 51.700 ;
        RECT 364.400 51.600 365.200 51.700 ;
        RECT 366.000 52.300 366.800 52.400 ;
        RECT 375.600 52.300 376.400 52.400 ;
        RECT 366.000 51.700 376.400 52.300 ;
        RECT 366.000 51.600 366.800 51.700 ;
        RECT 375.600 51.600 376.400 51.700 ;
        RECT 423.600 52.300 424.400 52.400 ;
        RECT 431.600 52.300 432.400 52.400 ;
        RECT 423.600 51.700 432.400 52.300 ;
        RECT 423.600 51.600 424.400 51.700 ;
        RECT 431.600 51.600 432.400 51.700 ;
        RECT 439.600 52.300 440.400 52.400 ;
        RECT 449.200 52.300 450.000 52.400 ;
        RECT 439.600 51.700 450.000 52.300 ;
        RECT 439.600 51.600 440.400 51.700 ;
        RECT 449.200 51.600 450.000 51.700 ;
        RECT 465.200 52.300 466.000 52.400 ;
        RECT 473.200 52.300 474.000 52.400 ;
        RECT 465.200 51.700 474.000 52.300 ;
        RECT 465.200 51.600 466.000 51.700 ;
        RECT 473.200 51.600 474.000 51.700 ;
        RECT 497.200 52.300 498.000 52.400 ;
        RECT 505.200 52.300 506.000 52.400 ;
        RECT 529.200 52.300 530.000 52.400 ;
        RECT 554.800 52.300 555.600 52.400 ;
        RECT 497.200 51.700 555.600 52.300 ;
        RECT 497.200 51.600 498.000 51.700 ;
        RECT 505.200 51.600 506.000 51.700 ;
        RECT 529.200 51.600 530.000 51.700 ;
        RECT 554.800 51.600 555.600 51.700 ;
        RECT 41.200 50.300 42.000 50.400 ;
        RECT 71.600 50.300 72.400 50.400 ;
        RECT 41.200 49.700 72.400 50.300 ;
        RECT 41.200 49.600 42.000 49.700 ;
        RECT 71.600 49.600 72.400 49.700 ;
        RECT 87.600 50.300 88.400 50.400 ;
        RECT 124.400 50.300 125.200 50.400 ;
        RECT 87.600 49.700 125.200 50.300 ;
        RECT 87.600 49.600 88.400 49.700 ;
        RECT 124.400 49.600 125.200 49.700 ;
        RECT 137.200 50.300 138.000 50.400 ;
        RECT 162.800 50.300 163.600 50.400 ;
        RECT 137.200 49.700 163.600 50.300 ;
        RECT 137.200 49.600 138.000 49.700 ;
        RECT 162.800 49.600 163.600 49.700 ;
        RECT 236.400 50.300 237.200 50.400 ;
        RECT 255.600 50.300 256.400 50.400 ;
        RECT 236.400 49.700 256.400 50.300 ;
        RECT 236.400 49.600 237.200 49.700 ;
        RECT 255.600 49.600 256.400 49.700 ;
        RECT 282.800 50.300 283.600 50.400 ;
        RECT 294.000 50.300 294.800 50.400 ;
        RECT 282.800 49.700 294.800 50.300 ;
        RECT 282.800 49.600 283.600 49.700 ;
        RECT 294.000 49.600 294.800 49.700 ;
        RECT 327.600 50.300 328.400 50.400 ;
        RECT 345.200 50.300 346.000 50.400 ;
        RECT 358.000 50.300 358.800 50.400 ;
        RECT 327.600 49.700 358.800 50.300 ;
        RECT 327.600 49.600 328.400 49.700 ;
        RECT 345.200 49.600 346.000 49.700 ;
        RECT 358.000 49.600 358.800 49.700 ;
        RECT 362.800 50.300 363.600 50.400 ;
        RECT 422.000 50.300 422.800 50.400 ;
        RECT 362.800 49.700 422.800 50.300 ;
        RECT 362.800 49.600 363.600 49.700 ;
        RECT 422.000 49.600 422.800 49.700 ;
        RECT 431.600 50.300 432.400 50.400 ;
        RECT 434.800 50.300 435.600 50.400 ;
        RECT 431.600 49.700 435.600 50.300 ;
        RECT 431.600 49.600 432.400 49.700 ;
        RECT 434.800 49.600 435.600 49.700 ;
        RECT 439.600 50.300 440.400 50.400 ;
        RECT 442.800 50.300 443.600 50.400 ;
        RECT 439.600 49.700 443.600 50.300 ;
        RECT 439.600 49.600 440.400 49.700 ;
        RECT 442.800 49.600 443.600 49.700 ;
        RECT 444.400 50.300 445.200 50.400 ;
        RECT 447.600 50.300 448.400 50.400 ;
        RECT 444.400 49.700 448.400 50.300 ;
        RECT 444.400 49.600 445.200 49.700 ;
        RECT 447.600 49.600 448.400 49.700 ;
        RECT 474.800 50.300 475.600 50.400 ;
        RECT 511.600 50.300 512.400 50.400 ;
        RECT 474.800 49.700 512.400 50.300 ;
        RECT 474.800 49.600 475.600 49.700 ;
        RECT 511.600 49.600 512.400 49.700 ;
        RECT 524.400 50.300 525.200 50.400 ;
        RECT 540.400 50.300 541.200 50.400 ;
        RECT 524.400 49.700 541.200 50.300 ;
        RECT 524.400 49.600 525.200 49.700 ;
        RECT 540.400 49.600 541.200 49.700 ;
        RECT 586.800 50.300 587.600 50.400 ;
        RECT 594.800 50.300 595.600 50.400 ;
        RECT 586.800 49.700 595.600 50.300 ;
        RECT 586.800 49.600 587.600 49.700 ;
        RECT 594.800 49.600 595.600 49.700 ;
        RECT 145.200 48.300 146.000 48.400 ;
        RECT 148.400 48.300 149.200 48.400 ;
        RECT 159.600 48.300 160.400 48.400 ;
        RECT 145.200 47.700 160.400 48.300 ;
        RECT 145.200 47.600 146.000 47.700 ;
        RECT 148.400 47.600 149.200 47.700 ;
        RECT 159.600 47.600 160.400 47.700 ;
        RECT 444.400 48.300 445.200 48.400 ;
        RECT 463.600 48.300 464.400 48.400 ;
        RECT 444.400 47.700 464.400 48.300 ;
        RECT 444.400 47.600 445.200 47.700 ;
        RECT 463.600 47.600 464.400 47.700 ;
        RECT 534.000 48.300 534.800 48.400 ;
        RECT 537.200 48.300 538.000 48.400 ;
        RECT 534.000 47.700 538.000 48.300 ;
        RECT 534.000 47.600 534.800 47.700 ;
        RECT 537.200 47.600 538.000 47.700 ;
        RECT 540.400 48.300 541.200 48.400 ;
        RECT 551.600 48.300 552.400 48.400 ;
        RECT 540.400 47.700 552.400 48.300 ;
        RECT 540.400 47.600 541.200 47.700 ;
        RECT 551.600 47.600 552.400 47.700 ;
        RECT 87.600 46.300 88.400 46.400 ;
        RECT 90.800 46.300 91.600 46.400 ;
        RECT 87.600 45.700 91.600 46.300 ;
        RECT 87.600 45.600 88.400 45.700 ;
        RECT 90.800 45.600 91.600 45.700 ;
        RECT 134.000 46.300 134.800 46.400 ;
        RECT 153.200 46.300 154.000 46.400 ;
        RECT 134.000 45.700 154.000 46.300 ;
        RECT 134.000 45.600 134.800 45.700 ;
        RECT 153.200 45.600 154.000 45.700 ;
        RECT 340.400 46.300 341.200 46.400 ;
        RECT 346.800 46.300 347.600 46.400 ;
        RECT 354.800 46.300 355.600 46.400 ;
        RECT 340.400 45.700 355.600 46.300 ;
        RECT 340.400 45.600 341.200 45.700 ;
        RECT 346.800 45.600 347.600 45.700 ;
        RECT 354.800 45.600 355.600 45.700 ;
        RECT 535.600 46.300 536.400 46.400 ;
        RECT 575.600 46.300 576.400 46.400 ;
        RECT 580.400 46.300 581.200 46.400 ;
        RECT 535.600 45.700 581.200 46.300 ;
        RECT 535.600 45.600 536.400 45.700 ;
        RECT 575.600 45.600 576.400 45.700 ;
        RECT 580.400 45.600 581.200 45.700 ;
        RECT 289.200 44.300 290.000 44.400 ;
        RECT 313.200 44.300 314.000 44.400 ;
        RECT 289.200 43.700 314.000 44.300 ;
        RECT 289.200 43.600 290.000 43.700 ;
        RECT 313.200 43.600 314.000 43.700 ;
        RECT 455.600 44.300 456.400 44.400 ;
        RECT 474.800 44.300 475.600 44.400 ;
        RECT 455.600 43.700 475.600 44.300 ;
        RECT 455.600 43.600 456.400 43.700 ;
        RECT 474.800 43.600 475.600 43.700 ;
        RECT 526.000 44.300 526.800 44.400 ;
        RECT 550.000 44.300 550.800 44.400 ;
        RECT 526.000 43.700 550.800 44.300 ;
        RECT 526.000 43.600 526.800 43.700 ;
        RECT 550.000 43.600 550.800 43.700 ;
        RECT 604.400 42.300 605.200 42.400 ;
        RECT 609.200 42.300 610.000 42.400 ;
        RECT 604.400 41.700 610.000 42.300 ;
        RECT 604.400 41.600 605.200 41.700 ;
        RECT 609.200 41.600 610.000 41.700 ;
        RECT 38.000 40.300 38.800 40.400 ;
        RECT 41.200 40.300 42.000 40.400 ;
        RECT 38.000 39.700 42.000 40.300 ;
        RECT 38.000 39.600 38.800 39.700 ;
        RECT 41.200 39.600 42.000 39.700 ;
        RECT 246.000 40.300 246.800 40.400 ;
        RECT 279.600 40.300 280.400 40.400 ;
        RECT 246.000 39.700 280.400 40.300 ;
        RECT 246.000 39.600 246.800 39.700 ;
        RECT 279.600 39.600 280.400 39.700 ;
        RECT 502.000 40.300 502.800 40.400 ;
        RECT 503.600 40.300 504.400 40.400 ;
        RECT 502.000 39.700 504.400 40.300 ;
        RECT 502.000 39.600 502.800 39.700 ;
        RECT 503.600 39.600 504.400 39.700 ;
        RECT 508.400 40.300 509.200 40.400 ;
        RECT 524.400 40.300 525.200 40.400 ;
        RECT 553.200 40.300 554.000 40.400 ;
        RECT 508.400 39.700 554.000 40.300 ;
        RECT 508.400 39.600 509.200 39.700 ;
        RECT 524.400 39.600 525.200 39.700 ;
        RECT 553.200 39.600 554.000 39.700 ;
        RECT 17.200 38.300 18.000 38.400 ;
        RECT 22.000 38.300 22.800 38.400 ;
        RECT 17.200 37.700 22.800 38.300 ;
        RECT 17.200 37.600 18.000 37.700 ;
        RECT 22.000 37.600 22.800 37.700 ;
        RECT 140.400 38.300 141.200 38.400 ;
        RECT 145.200 38.300 146.000 38.400 ;
        RECT 140.400 37.700 146.000 38.300 ;
        RECT 140.400 37.600 141.200 37.700 ;
        RECT 145.200 37.600 146.000 37.700 ;
        RECT 538.800 38.300 539.600 38.400 ;
        RECT 574.000 38.300 574.800 38.400 ;
        RECT 538.800 37.700 574.800 38.300 ;
        RECT 538.800 37.600 539.600 37.700 ;
        RECT 574.000 37.600 574.800 37.700 ;
        RECT 63.600 36.300 64.400 36.400 ;
        RECT 89.200 36.300 90.000 36.400 ;
        RECT 63.600 35.700 90.000 36.300 ;
        RECT 63.600 35.600 64.400 35.700 ;
        RECT 89.200 35.600 90.000 35.700 ;
        RECT 113.200 36.300 114.000 36.400 ;
        RECT 121.200 36.300 122.000 36.400 ;
        RECT 130.800 36.300 131.600 36.400 ;
        RECT 113.200 35.700 131.600 36.300 ;
        RECT 113.200 35.600 114.000 35.700 ;
        RECT 121.200 35.600 122.000 35.700 ;
        RECT 130.800 35.600 131.600 35.700 ;
        RECT 407.600 36.300 408.400 36.400 ;
        RECT 535.600 36.300 536.400 36.400 ;
        RECT 407.600 35.700 536.400 36.300 ;
        RECT 407.600 35.600 408.400 35.700 ;
        RECT 535.600 35.600 536.400 35.700 ;
        RECT 551.600 36.300 552.400 36.400 ;
        RECT 570.800 36.300 571.600 36.400 ;
        RECT 551.600 35.700 571.600 36.300 ;
        RECT 551.600 35.600 552.400 35.700 ;
        RECT 570.800 35.600 571.600 35.700 ;
        RECT 62.000 34.300 62.800 34.400 ;
        RECT 82.800 34.300 83.600 34.400 ;
        RECT 114.800 34.300 115.600 34.400 ;
        RECT 127.600 34.300 128.400 34.400 ;
        RECT 134.000 34.300 134.800 34.400 ;
        RECT 62.000 33.700 134.800 34.300 ;
        RECT 62.000 33.600 62.800 33.700 ;
        RECT 82.800 33.600 83.600 33.700 ;
        RECT 114.800 33.600 115.600 33.700 ;
        RECT 127.600 33.600 128.400 33.700 ;
        RECT 134.000 33.600 134.800 33.700 ;
        RECT 430.000 34.300 430.800 34.400 ;
        RECT 442.800 34.300 443.600 34.400 ;
        RECT 430.000 33.700 443.600 34.300 ;
        RECT 430.000 33.600 430.800 33.700 ;
        RECT 442.800 33.600 443.600 33.700 ;
        RECT 508.400 34.300 509.200 34.400 ;
        RECT 516.400 34.300 517.200 34.400 ;
        RECT 508.400 33.700 517.200 34.300 ;
        RECT 508.400 33.600 509.200 33.700 ;
        RECT 516.400 33.600 517.200 33.700 ;
        RECT 543.600 34.300 544.400 34.400 ;
        RECT 553.200 34.300 554.000 34.400 ;
        RECT 543.600 33.700 554.000 34.300 ;
        RECT 543.600 33.600 544.400 33.700 ;
        RECT 553.200 33.600 554.000 33.700 ;
        RECT 570.800 33.600 571.600 34.400 ;
        RECT 55.600 32.300 56.400 32.400 ;
        RECT 70.000 32.300 70.800 32.400 ;
        RECT 55.600 31.700 70.800 32.300 ;
        RECT 55.600 31.600 56.400 31.700 ;
        RECT 70.000 31.600 70.800 31.700 ;
        RECT 76.400 32.300 77.200 32.400 ;
        RECT 84.400 32.300 85.200 32.400 ;
        RECT 76.400 31.700 85.200 32.300 ;
        RECT 76.400 31.600 77.200 31.700 ;
        RECT 84.400 31.600 85.200 31.700 ;
        RECT 89.200 32.300 90.000 32.400 ;
        RECT 92.400 32.300 93.200 32.400 ;
        RECT 89.200 31.700 93.200 32.300 ;
        RECT 89.200 31.600 90.000 31.700 ;
        RECT 92.400 31.600 93.200 31.700 ;
        RECT 102.000 32.300 102.800 32.400 ;
        RECT 116.400 32.300 117.200 32.400 ;
        RECT 102.000 31.700 117.200 32.300 ;
        RECT 102.000 31.600 102.800 31.700 ;
        RECT 116.400 31.600 117.200 31.700 ;
        RECT 129.200 32.300 130.000 32.400 ;
        RECT 134.000 32.300 134.800 32.400 ;
        RECT 129.200 31.700 134.800 32.300 ;
        RECT 129.200 31.600 130.000 31.700 ;
        RECT 134.000 31.600 134.800 31.700 ;
        RECT 167.600 32.300 168.400 32.400 ;
        RECT 180.200 32.300 181.000 32.400 ;
        RECT 222.000 32.300 222.800 32.400 ;
        RECT 167.600 31.700 222.800 32.300 ;
        RECT 167.600 31.600 168.400 31.700 ;
        RECT 180.200 31.600 181.000 31.700 ;
        RECT 222.000 31.600 222.800 31.700 ;
        RECT 327.600 32.300 328.400 32.400 ;
        RECT 338.800 32.300 339.600 32.400 ;
        RECT 327.600 31.700 339.600 32.300 ;
        RECT 327.600 31.600 328.400 31.700 ;
        RECT 338.800 31.600 339.600 31.700 ;
        RECT 426.800 32.300 427.600 32.400 ;
        RECT 436.400 32.300 437.200 32.400 ;
        RECT 426.800 31.700 437.200 32.300 ;
        RECT 426.800 31.600 427.600 31.700 ;
        RECT 436.400 31.600 437.200 31.700 ;
        RECT 476.400 32.300 477.200 32.400 ;
        RECT 484.400 32.300 485.200 32.400 ;
        RECT 519.600 32.300 520.400 32.400 ;
        RECT 532.400 32.300 533.200 32.400 ;
        RECT 476.400 31.700 485.200 32.300 ;
        RECT 476.400 31.600 477.200 31.700 ;
        RECT 484.400 31.600 485.200 31.700 ;
        RECT 492.500 31.700 533.200 32.300 ;
        RECT 492.500 30.400 493.100 31.700 ;
        RECT 519.600 31.600 520.400 31.700 ;
        RECT 532.400 31.600 533.200 31.700 ;
        RECT 546.800 32.300 547.600 32.400 ;
        RECT 551.600 32.300 552.400 32.400 ;
        RECT 546.800 31.700 552.400 32.300 ;
        RECT 546.800 31.600 547.600 31.700 ;
        RECT 551.600 31.600 552.400 31.700 ;
        RECT 556.400 32.300 557.200 32.400 ;
        RECT 562.800 32.300 563.600 32.400 ;
        RECT 556.400 31.700 563.600 32.300 ;
        RECT 556.400 31.600 557.200 31.700 ;
        RECT 562.800 31.600 563.600 31.700 ;
        RECT 6.000 30.300 6.800 30.400 ;
        RECT 44.400 30.300 45.200 30.400 ;
        RECT 6.000 29.700 45.200 30.300 ;
        RECT 6.000 29.600 6.800 29.700 ;
        RECT 44.400 29.600 45.200 29.700 ;
        RECT 60.400 30.300 61.200 30.400 ;
        RECT 65.200 30.300 66.000 30.400 ;
        RECT 60.400 29.700 66.000 30.300 ;
        RECT 60.400 29.600 61.200 29.700 ;
        RECT 65.200 29.600 66.000 29.700 ;
        RECT 84.400 30.300 85.200 30.400 ;
        RECT 90.800 30.300 91.600 30.400 ;
        RECT 84.400 29.700 91.600 30.300 ;
        RECT 84.400 29.600 85.200 29.700 ;
        RECT 90.800 29.600 91.600 29.700 ;
        RECT 92.400 30.300 93.200 30.400 ;
        RECT 124.400 30.300 125.200 30.400 ;
        RECT 137.200 30.300 138.000 30.400 ;
        RECT 92.400 29.700 138.000 30.300 ;
        RECT 92.400 29.600 93.200 29.700 ;
        RECT 124.400 29.600 125.200 29.700 ;
        RECT 137.200 29.600 138.000 29.700 ;
        RECT 153.200 30.300 154.000 30.400 ;
        RECT 156.400 30.300 157.200 30.400 ;
        RECT 153.200 29.700 157.200 30.300 ;
        RECT 153.200 29.600 154.000 29.700 ;
        RECT 156.400 29.600 157.200 29.700 ;
        RECT 217.200 30.300 218.000 30.400 ;
        RECT 220.400 30.300 221.200 30.400 ;
        RECT 217.200 29.700 221.200 30.300 ;
        RECT 217.200 29.600 218.000 29.700 ;
        RECT 220.400 29.600 221.200 29.700 ;
        RECT 257.200 30.300 258.000 30.400 ;
        RECT 273.200 30.300 274.000 30.400 ;
        RECT 257.200 29.700 274.000 30.300 ;
        RECT 257.200 29.600 258.000 29.700 ;
        RECT 273.200 29.600 274.000 29.700 ;
        RECT 284.400 30.300 285.200 30.400 ;
        RECT 314.800 30.300 315.600 30.400 ;
        RECT 284.400 29.700 315.600 30.300 ;
        RECT 284.400 29.600 285.200 29.700 ;
        RECT 314.800 29.600 315.600 29.700 ;
        RECT 423.600 30.300 424.400 30.400 ;
        RECT 426.800 30.300 427.600 30.400 ;
        RECT 423.600 29.700 427.600 30.300 ;
        RECT 423.600 29.600 424.400 29.700 ;
        RECT 426.800 29.600 427.600 29.700 ;
        RECT 428.400 30.300 429.200 30.400 ;
        RECT 431.600 30.300 432.400 30.400 ;
        RECT 444.400 30.300 445.200 30.400 ;
        RECT 428.400 29.700 445.200 30.300 ;
        RECT 428.400 29.600 429.200 29.700 ;
        RECT 431.600 29.600 432.400 29.700 ;
        RECT 444.400 29.600 445.200 29.700 ;
        RECT 465.200 30.300 466.000 30.400 ;
        RECT 481.200 30.300 482.000 30.400 ;
        RECT 465.200 29.700 482.000 30.300 ;
        RECT 465.200 29.600 466.000 29.700 ;
        RECT 481.200 29.600 482.000 29.700 ;
        RECT 489.200 30.300 490.000 30.400 ;
        RECT 492.400 30.300 493.200 30.400 ;
        RECT 489.200 29.700 493.200 30.300 ;
        RECT 489.200 29.600 490.000 29.700 ;
        RECT 492.400 29.600 493.200 29.700 ;
        RECT 497.200 30.300 498.000 30.400 ;
        RECT 513.200 30.300 514.000 30.400 ;
        RECT 497.200 29.700 514.000 30.300 ;
        RECT 497.200 29.600 498.000 29.700 ;
        RECT 513.200 29.600 514.000 29.700 ;
        RECT 521.200 30.300 522.000 30.400 ;
        RECT 542.000 30.300 542.800 30.400 ;
        RECT 521.200 29.700 542.800 30.300 ;
        RECT 521.200 29.600 522.000 29.700 ;
        RECT 542.000 29.600 542.800 29.700 ;
        RECT 548.400 30.300 549.200 30.400 ;
        RECT 606.000 30.300 606.800 30.400 ;
        RECT 548.400 29.700 606.800 30.300 ;
        RECT 548.400 29.600 549.200 29.700 ;
        RECT 606.000 29.600 606.800 29.700 ;
        RECT 18.800 28.300 19.600 28.400 ;
        RECT 39.600 28.300 40.400 28.400 ;
        RECT 18.800 27.700 40.400 28.300 ;
        RECT 18.800 27.600 19.600 27.700 ;
        RECT 39.600 27.600 40.400 27.700 ;
        RECT 89.200 28.300 90.000 28.400 ;
        RECT 94.000 28.300 94.800 28.400 ;
        RECT 126.000 28.300 126.800 28.400 ;
        RECT 89.200 27.700 126.800 28.300 ;
        RECT 89.200 27.600 90.000 27.700 ;
        RECT 94.000 27.600 94.800 27.700 ;
        RECT 126.000 27.600 126.800 27.700 ;
        RECT 199.600 28.300 200.400 28.400 ;
        RECT 206.000 28.300 206.800 28.400 ;
        RECT 199.600 27.700 206.800 28.300 ;
        RECT 199.600 27.600 200.400 27.700 ;
        RECT 206.000 27.600 206.800 27.700 ;
        RECT 222.000 28.300 222.800 28.400 ;
        RECT 228.400 28.300 229.200 28.400 ;
        RECT 222.000 27.700 229.200 28.300 ;
        RECT 222.000 27.600 222.800 27.700 ;
        RECT 228.400 27.600 229.200 27.700 ;
        RECT 282.800 28.300 283.600 28.400 ;
        RECT 287.600 28.300 288.400 28.400 ;
        RECT 282.800 27.700 288.400 28.300 ;
        RECT 282.800 27.600 283.600 27.700 ;
        RECT 287.600 27.600 288.400 27.700 ;
        RECT 303.600 28.300 304.400 28.400 ;
        RECT 314.800 28.300 315.600 28.400 ;
        RECT 318.000 28.300 318.800 28.400 ;
        RECT 303.600 27.700 318.800 28.300 ;
        RECT 303.600 27.600 304.400 27.700 ;
        RECT 314.800 27.600 315.600 27.700 ;
        RECT 318.000 27.600 318.800 27.700 ;
        RECT 345.200 28.300 346.000 28.400 ;
        RECT 348.400 28.300 349.200 28.400 ;
        RECT 345.200 27.700 349.200 28.300 ;
        RECT 345.200 27.600 346.000 27.700 ;
        RECT 348.400 27.600 349.200 27.700 ;
        RECT 378.800 28.300 379.600 28.400 ;
        RECT 382.000 28.300 382.800 28.400 ;
        RECT 378.800 27.700 382.800 28.300 ;
        RECT 378.800 27.600 379.600 27.700 ;
        RECT 382.000 27.600 382.800 27.700 ;
        RECT 407.600 27.600 408.400 28.400 ;
        RECT 446.000 28.300 446.800 28.400 ;
        RECT 470.000 28.300 470.800 28.400 ;
        RECT 502.000 28.300 502.800 28.400 ;
        RECT 522.800 28.300 523.600 28.400 ;
        RECT 526.000 28.300 526.800 28.400 ;
        RECT 446.000 27.700 526.800 28.300 ;
        RECT 446.000 27.600 446.800 27.700 ;
        RECT 470.000 27.600 470.800 27.700 ;
        RECT 502.000 27.600 502.800 27.700 ;
        RECT 522.800 27.600 523.600 27.700 ;
        RECT 526.000 27.600 526.800 27.700 ;
        RECT 538.800 28.300 539.600 28.400 ;
        RECT 543.600 28.300 544.400 28.400 ;
        RECT 538.800 27.700 544.400 28.300 ;
        RECT 538.800 27.600 539.600 27.700 ;
        RECT 543.600 27.600 544.400 27.700 ;
        RECT 551.600 28.300 552.400 28.400 ;
        RECT 559.600 28.300 560.400 28.400 ;
        RECT 551.600 27.700 560.400 28.300 ;
        RECT 551.600 27.600 552.400 27.700 ;
        RECT 559.600 27.600 560.400 27.700 ;
        RECT 561.200 28.300 562.000 28.400 ;
        RECT 590.000 28.300 590.800 28.400 ;
        RECT 561.200 27.700 590.800 28.300 ;
        RECT 561.200 27.600 562.000 27.700 ;
        RECT 590.000 27.600 590.800 27.700 ;
        RECT 129.200 26.300 130.000 26.400 ;
        RECT 146.800 26.300 147.600 26.400 ;
        RECT 129.200 25.700 147.600 26.300 ;
        RECT 129.200 25.600 130.000 25.700 ;
        RECT 146.800 25.600 147.600 25.700 ;
        RECT 335.600 26.300 336.400 26.400 ;
        RECT 346.800 26.300 347.600 26.400 ;
        RECT 335.600 25.700 347.600 26.300 ;
        RECT 335.600 25.600 336.400 25.700 ;
        RECT 346.800 25.600 347.600 25.700 ;
        RECT 353.200 26.300 354.000 26.400 ;
        RECT 359.600 26.300 360.400 26.400 ;
        RECT 361.200 26.300 362.000 26.400 ;
        RECT 362.800 26.300 363.600 26.400 ;
        RECT 353.200 25.700 363.600 26.300 ;
        RECT 353.200 25.600 354.000 25.700 ;
        RECT 359.600 25.600 360.400 25.700 ;
        RECT 361.200 25.600 362.000 25.700 ;
        RECT 362.800 25.600 363.600 25.700 ;
        RECT 457.200 26.300 458.000 26.400 ;
        RECT 478.000 26.300 478.800 26.400 ;
        RECT 482.800 26.300 483.600 26.400 ;
        RECT 510.000 26.300 510.800 26.400 ;
        RECT 524.400 26.300 525.200 26.400 ;
        RECT 457.200 25.700 525.200 26.300 ;
        RECT 457.200 25.600 458.000 25.700 ;
        RECT 478.000 25.600 478.800 25.700 ;
        RECT 482.800 25.600 483.600 25.700 ;
        RECT 510.000 25.600 510.800 25.700 ;
        RECT 524.400 25.600 525.200 25.700 ;
        RECT 558.000 26.300 558.800 26.400 ;
        RECT 562.800 26.300 563.600 26.400 ;
        RECT 558.000 25.700 563.600 26.300 ;
        RECT 558.000 25.600 558.800 25.700 ;
        RECT 562.800 25.600 563.600 25.700 ;
        RECT 586.800 26.300 587.600 26.400 ;
        RECT 590.000 26.300 590.800 26.400 ;
        RECT 586.800 25.700 590.800 26.300 ;
        RECT 586.800 25.600 587.600 25.700 ;
        RECT 590.000 25.600 590.800 25.700 ;
        RECT 86.000 24.300 86.800 24.400 ;
        RECT 90.800 24.300 91.600 24.400 ;
        RECT 86.000 23.700 91.600 24.300 ;
        RECT 86.000 23.600 86.800 23.700 ;
        RECT 90.800 23.600 91.600 23.700 ;
        RECT 146.800 24.300 147.600 24.400 ;
        RECT 162.800 24.300 163.600 24.400 ;
        RECT 146.800 23.700 163.600 24.300 ;
        RECT 146.800 23.600 147.600 23.700 ;
        RECT 162.800 23.600 163.600 23.700 ;
        RECT 452.400 24.300 453.200 24.400 ;
        RECT 489.200 24.300 490.000 24.400 ;
        RECT 521.200 24.300 522.000 24.400 ;
        RECT 538.800 24.300 539.600 24.400 ;
        RECT 545.200 24.300 546.000 24.400 ;
        RECT 452.400 23.700 546.000 24.300 ;
        RECT 452.400 23.600 453.200 23.700 ;
        RECT 489.200 23.600 490.000 23.700 ;
        RECT 521.200 23.600 522.000 23.700 ;
        RECT 538.800 23.600 539.600 23.700 ;
        RECT 545.200 23.600 546.000 23.700 ;
        RECT 30.000 22.300 30.800 22.400 ;
        RECT 154.800 22.300 155.600 22.400 ;
        RECT 30.000 21.700 155.600 22.300 ;
        RECT 30.000 21.600 30.800 21.700 ;
        RECT 154.800 21.600 155.600 21.700 ;
        RECT 231.600 22.300 232.400 22.400 ;
        RECT 252.400 22.300 253.200 22.400 ;
        RECT 231.600 21.700 253.200 22.300 ;
        RECT 231.600 21.600 232.400 21.700 ;
        RECT 252.400 21.600 253.200 21.700 ;
        RECT 375.600 22.300 376.400 22.400 ;
        RECT 380.400 22.300 381.200 22.400 ;
        RECT 375.600 21.700 381.200 22.300 ;
        RECT 375.600 21.600 376.400 21.700 ;
        RECT 380.400 21.600 381.200 21.700 ;
        RECT 423.600 22.300 424.400 22.400 ;
        RECT 433.200 22.300 434.000 22.400 ;
        RECT 463.600 22.300 464.400 22.400 ;
        RECT 423.600 21.700 464.400 22.300 ;
        RECT 423.600 21.600 424.400 21.700 ;
        RECT 433.200 21.600 434.000 21.700 ;
        RECT 463.600 21.600 464.400 21.700 ;
        RECT 17.200 20.300 18.000 20.400 ;
        RECT 22.000 20.300 22.800 20.400 ;
        RECT 54.000 20.300 54.800 20.400 ;
        RECT 17.200 19.700 54.800 20.300 ;
        RECT 17.200 19.600 18.000 19.700 ;
        RECT 22.000 19.600 22.800 19.700 ;
        RECT 54.000 19.600 54.800 19.700 ;
        RECT 76.400 20.300 77.200 20.400 ;
        RECT 100.400 20.300 101.200 20.400 ;
        RECT 76.400 19.700 101.200 20.300 ;
        RECT 76.400 19.600 77.200 19.700 ;
        RECT 100.400 19.600 101.200 19.700 ;
        RECT 126.000 20.300 126.800 20.400 ;
        RECT 130.800 20.300 131.600 20.400 ;
        RECT 138.800 20.300 139.600 20.400 ;
        RECT 164.400 20.300 165.200 20.400 ;
        RECT 126.000 19.700 165.200 20.300 ;
        RECT 126.000 19.600 126.800 19.700 ;
        RECT 130.800 19.600 131.600 19.700 ;
        RECT 138.800 19.600 139.600 19.700 ;
        RECT 164.400 19.600 165.200 19.700 ;
        RECT 183.600 20.300 184.400 20.400 ;
        RECT 185.200 20.300 186.000 20.400 ;
        RECT 188.400 20.300 189.200 20.400 ;
        RECT 183.600 19.700 189.200 20.300 ;
        RECT 183.600 19.600 184.400 19.700 ;
        RECT 185.200 19.600 186.000 19.700 ;
        RECT 188.400 19.600 189.200 19.700 ;
        RECT 260.400 20.300 261.200 20.400 ;
        RECT 274.800 20.300 275.600 20.400 ;
        RECT 260.400 19.700 275.600 20.300 ;
        RECT 260.400 19.600 261.200 19.700 ;
        RECT 274.800 19.600 275.600 19.700 ;
        RECT 327.600 20.300 328.400 20.400 ;
        RECT 334.000 20.300 334.800 20.400 ;
        RECT 327.600 19.700 334.800 20.300 ;
        RECT 327.600 19.600 328.400 19.700 ;
        RECT 334.000 19.600 334.800 19.700 ;
        RECT 433.200 20.300 434.000 20.400 ;
        RECT 447.600 20.300 448.400 20.400 ;
        RECT 465.200 20.300 466.000 20.400 ;
        RECT 433.200 19.700 466.000 20.300 ;
        RECT 433.200 19.600 434.000 19.700 ;
        RECT 447.600 19.600 448.400 19.700 ;
        RECT 465.200 19.600 466.000 19.700 ;
        RECT 36.400 18.300 37.200 18.400 ;
        RECT 50.800 18.300 51.600 18.400 ;
        RECT 73.200 18.300 74.000 18.400 ;
        RECT 36.400 17.700 74.000 18.300 ;
        RECT 36.400 17.600 37.200 17.700 ;
        RECT 50.800 17.600 51.600 17.700 ;
        RECT 73.200 17.600 74.000 17.700 ;
        RECT 110.000 18.300 110.800 18.400 ;
        RECT 134.000 18.300 134.800 18.400 ;
        RECT 110.000 17.700 134.800 18.300 ;
        RECT 110.000 17.600 110.800 17.700 ;
        RECT 134.000 17.600 134.800 17.700 ;
        RECT 236.400 18.300 237.200 18.400 ;
        RECT 249.200 18.300 250.000 18.400 ;
        RECT 258.800 18.300 259.600 18.400 ;
        RECT 286.000 18.300 286.800 18.400 ;
        RECT 311.600 18.300 312.400 18.400 ;
        RECT 330.800 18.300 331.600 18.400 ;
        RECT 394.800 18.300 395.600 18.400 ;
        RECT 236.400 17.700 395.600 18.300 ;
        RECT 236.400 17.600 237.200 17.700 ;
        RECT 249.200 17.600 250.000 17.700 ;
        RECT 258.800 17.600 259.600 17.700 ;
        RECT 286.000 17.600 286.800 17.700 ;
        RECT 311.600 17.600 312.400 17.700 ;
        RECT 330.800 17.600 331.600 17.700 ;
        RECT 394.800 17.600 395.600 17.700 ;
        RECT 396.400 18.300 397.200 18.400 ;
        RECT 404.400 18.300 405.200 18.400 ;
        RECT 396.400 17.700 405.200 18.300 ;
        RECT 396.400 17.600 397.200 17.700 ;
        RECT 404.400 17.600 405.200 17.700 ;
        RECT 559.600 18.300 560.400 18.400 ;
        RECT 564.400 18.300 565.200 18.400 ;
        RECT 590.000 18.300 590.800 18.400 ;
        RECT 559.600 17.700 590.800 18.300 ;
        RECT 559.600 17.600 560.400 17.700 ;
        RECT 564.400 17.600 565.200 17.700 ;
        RECT 590.000 17.600 590.800 17.700 ;
        RECT 33.200 16.300 34.000 16.400 ;
        RECT 41.200 16.300 42.000 16.400 ;
        RECT 33.200 15.700 42.000 16.300 ;
        RECT 33.200 15.600 34.000 15.700 ;
        RECT 41.200 15.600 42.000 15.700 ;
        RECT 78.000 16.300 78.800 16.400 ;
        RECT 82.800 16.300 83.600 16.400 ;
        RECT 78.000 15.700 83.600 16.300 ;
        RECT 78.000 15.600 78.800 15.700 ;
        RECT 82.800 15.600 83.600 15.700 ;
        RECT 97.200 16.300 98.000 16.400 ;
        RECT 134.000 16.300 134.800 16.400 ;
        RECT 97.200 15.700 134.800 16.300 ;
        RECT 97.200 15.600 98.000 15.700 ;
        RECT 134.000 15.600 134.800 15.700 ;
        RECT 162.800 16.300 163.600 16.400 ;
        RECT 196.400 16.300 197.200 16.400 ;
        RECT 162.800 15.700 197.200 16.300 ;
        RECT 162.800 15.600 163.600 15.700 ;
        RECT 196.400 15.600 197.200 15.700 ;
        RECT 350.000 16.300 350.800 16.400 ;
        RECT 359.600 16.300 360.400 16.400 ;
        RECT 350.000 15.700 360.400 16.300 ;
        RECT 350.000 15.600 350.800 15.700 ;
        RECT 359.600 15.600 360.400 15.700 ;
        RECT 380.400 16.300 381.200 16.400 ;
        RECT 409.200 16.300 410.000 16.400 ;
        RECT 380.400 15.700 410.000 16.300 ;
        RECT 380.400 15.600 381.200 15.700 ;
        RECT 409.200 15.600 410.000 15.700 ;
        RECT 553.200 16.300 554.000 16.400 ;
        RECT 593.200 16.300 594.000 16.400 ;
        RECT 553.200 15.700 594.000 16.300 ;
        RECT 553.200 15.600 554.000 15.700 ;
        RECT 593.200 15.600 594.000 15.700 ;
        RECT 14.000 14.300 14.800 14.400 ;
        RECT 42.800 14.300 43.600 14.400 ;
        RECT 14.000 13.700 43.600 14.300 ;
        RECT 14.000 13.600 14.800 13.700 ;
        RECT 42.800 13.600 43.600 13.700 ;
        RECT 82.800 14.300 83.600 14.400 ;
        RECT 102.000 14.300 102.800 14.400 ;
        RECT 82.800 13.700 102.800 14.300 ;
        RECT 82.800 13.600 83.600 13.700 ;
        RECT 102.000 13.600 102.800 13.700 ;
        RECT 166.000 14.300 166.800 14.400 ;
        RECT 172.400 14.300 173.200 14.400 ;
        RECT 166.000 13.700 173.200 14.300 ;
        RECT 166.000 13.600 166.800 13.700 ;
        RECT 172.400 13.600 173.200 13.700 ;
        RECT 193.200 14.300 194.000 14.400 ;
        RECT 217.200 14.300 218.000 14.400 ;
        RECT 193.200 13.700 218.000 14.300 ;
        RECT 193.200 13.600 194.000 13.700 ;
        RECT 217.200 13.600 218.000 13.700 ;
        RECT 223.600 14.300 224.400 14.400 ;
        RECT 233.200 14.300 234.000 14.400 ;
        RECT 223.600 13.700 234.000 14.300 ;
        RECT 223.600 13.600 224.400 13.700 ;
        RECT 233.200 13.600 234.000 13.700 ;
        RECT 282.800 13.600 283.600 14.400 ;
        RECT 359.600 14.300 360.400 14.400 ;
        RECT 377.200 14.300 378.000 14.400 ;
        RECT 359.600 13.700 378.000 14.300 ;
        RECT 359.600 13.600 360.400 13.700 ;
        RECT 377.200 13.600 378.000 13.700 ;
        RECT 410.800 14.300 411.600 14.400 ;
        RECT 425.200 14.300 426.000 14.400 ;
        RECT 410.800 13.700 426.000 14.300 ;
        RECT 410.800 13.600 411.600 13.700 ;
        RECT 425.200 13.600 426.000 13.700 ;
        RECT 446.000 14.300 446.800 14.400 ;
        RECT 452.400 14.300 453.200 14.400 ;
        RECT 446.000 13.700 453.200 14.300 ;
        RECT 446.000 13.600 446.800 13.700 ;
        RECT 452.400 13.600 453.200 13.700 ;
        RECT 455.600 14.300 456.400 14.400 ;
        RECT 466.800 14.300 467.600 14.400 ;
        RECT 455.600 13.700 467.600 14.300 ;
        RECT 455.600 13.600 456.400 13.700 ;
        RECT 466.800 13.600 467.600 13.700 ;
        RECT 478.000 14.300 478.800 14.400 ;
        RECT 484.400 14.300 485.200 14.400 ;
        RECT 478.000 13.700 485.200 14.300 ;
        RECT 478.000 13.600 478.800 13.700 ;
        RECT 484.400 13.600 485.200 13.700 ;
        RECT 489.200 14.300 490.000 14.400 ;
        RECT 494.000 14.300 494.800 14.400 ;
        RECT 489.200 13.700 494.800 14.300 ;
        RECT 489.200 13.600 490.000 13.700 ;
        RECT 494.000 13.600 494.800 13.700 ;
        RECT 521.200 14.300 522.000 14.400 ;
        RECT 530.800 14.300 531.600 14.400 ;
        RECT 543.600 14.300 544.400 14.400 ;
        RECT 521.200 13.700 544.400 14.300 ;
        RECT 521.200 13.600 522.000 13.700 ;
        RECT 530.800 13.600 531.600 13.700 ;
        RECT 543.600 13.600 544.400 13.700 ;
        RECT 545.200 14.300 546.000 14.400 ;
        RECT 566.000 14.300 566.800 14.400 ;
        RECT 545.200 13.700 566.800 14.300 ;
        RECT 545.200 13.600 546.000 13.700 ;
        RECT 566.000 13.600 566.800 13.700 ;
        RECT 4.400 12.300 5.200 12.400 ;
        RECT 34.800 12.300 35.600 12.400 ;
        RECT 38.000 12.300 38.800 12.400 ;
        RECT 4.400 11.700 38.800 12.300 ;
        RECT 4.400 11.600 5.200 11.700 ;
        RECT 34.800 11.600 35.600 11.700 ;
        RECT 38.000 11.600 38.800 11.700 ;
        RECT 52.400 12.300 53.200 12.400 ;
        RECT 78.000 12.300 78.800 12.400 ;
        RECT 97.200 12.300 98.000 12.400 ;
        RECT 52.400 11.700 98.000 12.300 ;
        RECT 52.400 11.600 53.200 11.700 ;
        RECT 78.000 11.600 78.800 11.700 ;
        RECT 97.200 11.600 98.000 11.700 ;
        RECT 100.400 12.300 101.200 12.400 ;
        RECT 116.400 12.300 117.200 12.400 ;
        RECT 100.400 11.700 117.200 12.300 ;
        RECT 100.400 11.600 101.200 11.700 ;
        RECT 116.400 11.600 117.200 11.700 ;
        RECT 122.800 12.300 123.600 12.400 ;
        RECT 132.400 12.300 133.200 12.400 ;
        RECT 122.800 11.700 133.200 12.300 ;
        RECT 122.800 11.600 123.600 11.700 ;
        RECT 132.400 11.600 133.200 11.700 ;
        RECT 177.200 12.300 178.000 12.400 ;
        RECT 183.600 12.300 184.400 12.400 ;
        RECT 177.200 11.700 184.400 12.300 ;
        RECT 177.200 11.600 178.000 11.700 ;
        RECT 183.600 11.600 184.400 11.700 ;
        RECT 204.400 12.300 205.200 12.400 ;
        RECT 223.600 12.300 224.400 12.400 ;
        RECT 204.400 11.700 224.400 12.300 ;
        RECT 204.400 11.600 205.200 11.700 ;
        RECT 223.600 11.600 224.400 11.700 ;
        RECT 297.200 12.300 298.000 12.400 ;
        RECT 318.000 12.300 318.800 12.400 ;
        RECT 297.200 11.700 318.800 12.300 ;
        RECT 297.200 11.600 298.000 11.700 ;
        RECT 318.000 11.600 318.800 11.700 ;
        RECT 430.000 12.300 430.800 12.400 ;
        RECT 474.800 12.300 475.600 12.400 ;
        RECT 430.000 11.700 475.600 12.300 ;
        RECT 430.000 11.600 430.800 11.700 ;
        RECT 474.800 11.600 475.600 11.700 ;
        RECT 481.200 12.300 482.000 12.400 ;
        RECT 518.000 12.300 518.800 12.400 ;
        RECT 522.800 12.300 523.600 12.400 ;
        RECT 481.200 11.700 523.600 12.300 ;
        RECT 481.200 11.600 482.000 11.700 ;
        RECT 518.000 11.600 518.800 11.700 ;
        RECT 522.800 11.600 523.600 11.700 ;
        RECT 529.200 12.300 530.000 12.400 ;
        RECT 554.800 12.300 555.600 12.400 ;
        RECT 529.200 11.700 555.600 12.300 ;
        RECT 529.200 11.600 530.000 11.700 ;
        RECT 554.800 11.600 555.600 11.700 ;
        RECT 567.600 12.300 568.400 12.400 ;
        RECT 583.600 12.300 584.400 12.400 ;
        RECT 567.600 11.700 584.400 12.300 ;
        RECT 567.600 11.600 568.400 11.700 ;
        RECT 583.600 11.600 584.400 11.700 ;
        RECT 449.200 10.300 450.000 10.400 ;
        RECT 452.400 10.300 453.200 10.400 ;
        RECT 449.200 9.700 453.200 10.300 ;
        RECT 449.200 9.600 450.000 9.700 ;
        RECT 452.400 9.600 453.200 9.700 ;
        RECT 479.600 10.300 480.400 10.400 ;
        RECT 489.200 10.300 490.000 10.400 ;
        RECT 503.600 10.300 504.400 10.400 ;
        RECT 513.200 10.300 514.000 10.400 ;
        RECT 479.600 9.700 514.000 10.300 ;
        RECT 479.600 9.600 480.400 9.700 ;
        RECT 489.200 9.600 490.000 9.700 ;
        RECT 503.600 9.600 504.400 9.700 ;
        RECT 513.200 9.600 514.000 9.700 ;
        RECT 518.000 10.300 518.800 10.400 ;
        RECT 526.000 10.300 526.800 10.400 ;
        RECT 518.000 9.700 526.800 10.300 ;
        RECT 518.000 9.600 518.800 9.700 ;
        RECT 526.000 9.600 526.800 9.700 ;
        RECT 551.600 10.300 552.400 10.400 ;
        RECT 570.800 10.300 571.600 10.400 ;
        RECT 551.600 9.700 571.600 10.300 ;
        RECT 551.600 9.600 552.400 9.700 ;
        RECT 570.800 9.600 571.600 9.700 ;
        RECT 422.000 8.300 422.800 8.400 ;
        RECT 425.200 8.300 426.000 8.400 ;
        RECT 434.800 8.300 435.600 8.400 ;
        RECT 422.000 7.700 435.600 8.300 ;
        RECT 422.000 7.600 422.800 7.700 ;
        RECT 425.200 7.600 426.000 7.700 ;
        RECT 434.800 7.600 435.600 7.700 ;
        RECT 487.600 8.300 488.400 8.400 ;
        RECT 500.400 8.300 501.200 8.400 ;
        RECT 487.600 7.700 501.200 8.300 ;
        RECT 487.600 7.600 488.400 7.700 ;
        RECT 500.400 7.600 501.200 7.700 ;
      LAYER metal4 ;
        RECT 17.000 435.400 18.200 484.600 ;
        RECT 13.800 319.400 15.000 428.600 ;
        RECT 33.000 411.400 34.200 546.600 ;
        RECT 122.600 541.400 123.800 550.600 ;
        RECT 36.200 427.400 37.400 530.600 ;
        RECT 45.800 513.400 47.000 536.600 ;
        RECT 45.800 457.400 47.000 510.600 ;
        RECT 42.600 387.400 43.800 454.600 ;
        RECT 52.200 453.400 53.400 532.600 ;
        RECT 65.000 489.400 66.200 524.600 ;
        RECT 87.400 441.400 88.600 492.600 ;
        RECT 45.800 383.400 47.000 398.600 ;
        RECT 58.600 389.400 59.800 430.600 ;
        RECT 90.600 373.400 91.800 496.600 ;
        RECT 97.000 493.400 98.200 534.600 ;
        RECT 93.800 467.400 95.000 472.600 ;
        RECT 103.400 451.400 104.600 490.600 ;
        RECT 135.400 469.400 136.600 480.600 ;
        RECT 170.600 467.400 171.800 502.600 ;
        RECT 106.600 375.400 107.800 382.600 ;
        RECT 116.200 351.400 117.400 416.600 ;
        RECT 129.000 377.400 130.200 422.600 ;
        RECT 132.200 375.400 133.400 446.600 ;
        RECT 135.400 423.400 136.600 442.600 ;
        RECT 161.000 411.400 162.200 444.600 ;
        RECT 167.400 409.400 168.600 438.600 ;
        RECT 177.000 411.400 178.200 460.600 ;
        RECT 189.800 449.400 191.000 508.600 ;
        RECT 196.200 429.400 197.400 486.600 ;
        RECT 189.800 375.400 191.000 420.600 ;
        RECT 202.600 401.400 203.800 428.600 ;
        RECT 221.800 361.400 223.000 432.600 ;
        RECT 225.000 391.400 226.200 498.600 ;
        RECT 244.200 495.400 245.400 536.600 ;
        RECT 109.800 273.400 111.000 322.600 ;
        RECT 129.000 317.400 130.200 358.600 ;
        RECT 138.600 267.400 139.800 320.600 ;
        RECT 196.200 275.400 197.400 344.600 ;
        RECT 205.800 283.400 207.000 318.600 ;
        RECT 228.200 281.400 229.400 350.600 ;
        RECT 231.400 341.400 232.600 422.600 ;
        RECT 237.800 315.400 239.000 370.600 ;
        RECT 241.000 359.400 242.200 470.600 ;
        RECT 250.600 441.400 251.800 544.600 ;
        RECT 372.200 513.400 373.400 538.600 ;
        RECT 266.600 389.400 267.800 438.600 ;
        RECT 276.200 373.400 277.400 494.600 ;
        RECT 282.600 381.400 283.800 492.600 ;
        RECT 295.400 489.400 296.600 504.600 ;
        RECT 330.600 471.400 331.800 498.600 ;
        RECT 244.200 283.400 245.400 366.600 ;
        RECT 269.800 307.400 271.000 340.600 ;
        RECT 292.200 339.400 293.400 398.600 ;
        RECT 295.400 327.400 296.600 440.600 ;
        RECT 298.600 329.400 299.800 446.600 ;
        RECT 337.000 347.400 338.200 422.600 ;
        RECT 340.200 397.400 341.400 464.600 ;
        RECT 381.800 409.400 383.000 476.600 ;
        RECT 391.400 475.400 392.600 500.600 ;
        RECT 397.800 479.400 399.000 514.600 ;
        RECT 410.600 485.400 411.800 518.600 ;
        RECT 413.800 463.400 415.000 510.600 ;
        RECT 426.600 467.400 427.800 490.600 ;
        RECT 439.400 485.400 440.600 512.600 ;
        RECT 397.800 427.400 399.000 462.600 ;
        RECT 343.400 339.400 344.600 408.600 ;
        RECT 420.200 371.400 421.400 420.600 ;
        RECT 442.600 375.400 443.800 522.600 ;
        RECT 449.000 475.400 450.200 482.600 ;
        RECT 465.000 481.400 466.200 512.600 ;
        RECT 487.400 503.400 488.600 508.600 ;
        RECT 468.200 453.400 469.400 472.600 ;
        RECT 503.400 471.400 504.600 496.600 ;
        RECT 519.400 483.400 520.600 532.600 ;
        RECT 525.800 507.400 527.000 536.600 ;
        RECT 474.600 405.400 475.800 454.600 ;
        RECT 493.800 431.400 495.000 468.600 ;
        RECT 506.600 437.400 507.800 456.600 ;
        RECT 516.200 451.400 517.400 460.600 ;
        RECT 509.800 411.400 511.000 416.600 ;
        RECT 4.200 69.400 5.400 212.600 ;
        RECT 13.800 129.400 15.000 190.600 ;
        RECT 36.200 183.400 37.400 264.600 ;
        RECT 199.400 259.400 200.600 280.600 ;
        RECT 250.600 277.400 251.800 284.600 ;
        RECT 273.000 279.400 274.200 312.600 ;
        RECT 292.200 283.400 293.400 312.600 ;
        RECT 36.200 95.400 37.400 152.600 ;
        RECT 42.600 123.400 43.800 160.600 ;
        RECT 45.800 63.400 47.000 104.600 ;
        RECT 52.200 11.400 53.400 82.600 ;
        RECT 55.400 55.400 56.600 222.600 ;
        RECT 81.000 93.400 82.200 172.600 ;
        RECT 84.200 91.400 85.400 198.600 ;
        RECT 93.800 111.400 95.000 132.600 ;
        RECT 97.000 93.400 98.200 132.600 ;
        RECT 100.200 91.400 101.400 122.600 ;
        RECT 122.600 111.400 123.800 180.600 ;
        RECT 106.600 85.400 107.800 106.600 ;
        RECT 135.400 87.400 136.600 156.600 ;
        RECT 138.600 107.400 139.800 140.600 ;
        RECT 141.800 121.400 143.000 164.600 ;
        RECT 71.400 67.400 72.600 72.600 ;
        RECT 145.000 55.400 146.200 190.600 ;
        RECT 157.800 129.400 159.000 168.600 ;
        RECT 205.800 163.400 207.000 190.600 ;
        RECT 209.000 175.400 210.200 190.600 ;
        RECT 221.800 177.400 223.000 214.600 ;
        RECT 241.000 175.400 242.200 244.600 ;
        RECT 260.200 215.400 261.400 256.600 ;
        RECT 273.000 231.400 274.200 254.600 ;
        RECT 285.800 249.400 287.000 268.600 ;
        RECT 295.400 253.400 296.600 302.600 ;
        RECT 311.400 297.400 312.600 314.600 ;
        RECT 298.600 231.400 299.800 268.600 ;
        RECT 314.600 265.400 315.800 304.600 ;
        RECT 321.000 251.400 322.200 282.600 ;
        RECT 324.200 281.400 325.400 322.600 ;
        RECT 346.600 317.400 347.800 350.600 ;
        RECT 375.400 309.400 376.600 326.600 ;
        RECT 378.600 325.400 379.800 370.600 ;
        RECT 327.400 267.400 328.600 284.600 ;
        RECT 314.600 231.400 315.800 246.600 ;
        RECT 324.200 243.400 325.400 266.600 ;
        RECT 346.600 237.400 347.800 248.600 ;
        RECT 311.400 201.400 312.600 222.600 ;
        RECT 321.000 203.400 322.200 230.600 ;
        RECT 161.000 79.400 162.200 156.600 ;
        RECT 193.000 73.400 194.200 116.600 ;
        RECT 205.800 27.400 207.000 132.600 ;
        RECT 215.400 53.400 216.600 170.600 ;
        RECT 257.000 29.400 258.200 120.600 ;
        RECT 285.800 113.400 287.000 190.600 ;
        RECT 311.400 149.400 312.600 190.600 ;
        RECT 317.800 175.400 319.000 196.600 ;
        RECT 340.200 169.400 341.400 230.600 ;
        RECT 349.800 223.400 351.000 260.600 ;
        RECT 353.000 241.400 354.200 306.600 ;
        RECT 359.400 229.400 360.600 276.600 ;
        RECT 362.600 259.400 363.800 286.600 ;
        RECT 365.800 271.400 367.000 288.600 ;
        RECT 365.800 225.400 367.000 254.600 ;
        RECT 343.400 181.400 344.600 194.600 ;
        RECT 346.600 189.400 347.800 204.600 ;
        RECT 295.400 93.400 296.600 108.600 ;
        RECT 333.800 97.400 335.000 132.600 ;
        RECT 369.000 113.400 370.200 140.600 ;
        RECT 372.200 127.400 373.400 264.600 ;
        RECT 378.600 263.400 379.800 308.600 ;
        RECT 391.400 293.400 392.600 308.600 ;
        RECT 404.200 303.400 405.400 350.600 ;
        RECT 410.600 311.400 411.800 342.600 ;
        RECT 449.000 307.400 450.200 330.600 ;
        RECT 465.000 313.400 466.200 320.600 ;
        RECT 381.800 275.400 383.000 288.600 ;
        RECT 394.600 267.400 395.800 290.600 ;
        RECT 401.000 277.400 402.200 302.600 ;
        RECT 404.200 235.400 405.400 286.600 ;
        RECT 417.000 241.400 418.200 306.600 ;
        RECT 420.200 249.400 421.400 266.600 ;
        RECT 429.800 255.400 431.000 288.600 ;
        RECT 433.000 261.400 434.200 280.600 ;
        RECT 468.200 263.400 469.400 310.600 ;
        RECT 474.600 263.400 475.800 380.600 ;
        RECT 490.600 353.400 491.800 404.600 ;
        RECT 493.800 305.400 495.000 332.600 ;
        RECT 500.200 301.400 501.400 310.600 ;
        RECT 503.400 307.400 504.600 314.600 ;
        RECT 506.600 297.400 507.800 312.600 ;
        RECT 477.800 259.400 479.000 282.600 ;
        RECT 484.200 249.400 485.400 294.600 ;
        RECT 487.400 253.400 488.600 264.600 ;
        RECT 423.400 239.400 424.600 244.600 ;
        RECT 381.800 221.400 383.000 228.600 ;
        RECT 381.800 105.400 383.000 210.600 ;
        RECT 407.400 183.400 408.600 236.600 ;
        RECT 465.000 223.400 466.200 244.600 ;
        RECT 503.400 243.400 504.600 264.600 ;
        RECT 506.600 263.400 507.800 294.600 ;
        RECT 509.800 293.400 511.000 322.600 ;
        RECT 519.400 321.400 520.600 466.600 ;
        RECT 522.600 311.400 523.800 442.600 ;
        RECT 529.000 331.400 530.200 346.600 ;
        RECT 535.400 321.400 536.600 438.600 ;
        RECT 538.600 333.400 539.800 362.600 ;
        RECT 541.800 357.400 543.000 518.600 ;
        RECT 557.800 493.400 559.000 544.600 ;
        RECT 519.400 269.400 520.600 296.600 ;
        RECT 509.800 251.400 511.000 268.600 ;
        RECT 525.800 253.400 527.000 266.600 ;
        RECT 529.000 255.400 530.200 276.600 ;
        RECT 468.200 227.400 469.400 242.600 ;
        RECT 471.400 231.400 472.600 242.600 ;
        RECT 532.200 231.400 533.400 254.600 ;
        RECT 538.600 243.400 539.800 306.600 ;
        RECT 541.800 267.400 543.000 302.600 ;
        RECT 97.000 11.400 98.200 16.600 ;
        RECT 282.600 13.400 283.800 28.600 ;
        RECT 317.800 27.400 319.000 76.600 ;
        RECT 359.400 53.400 360.600 94.600 ;
        RECT 365.800 51.400 367.000 92.600 ;
        RECT 381.800 27.400 383.000 56.600 ;
        RECT 394.600 53.400 395.800 74.600 ;
        RECT 401.000 61.400 402.200 102.600 ;
        RECT 404.200 17.400 405.400 130.600 ;
        RECT 407.400 27.400 408.600 108.600 ;
        RECT 410.600 107.400 411.800 198.600 ;
        RECT 410.600 69.400 411.800 102.600 ;
        RECT 429.800 91.400 431.000 114.600 ;
        RECT 436.200 77.400 437.400 92.600 ;
        RECT 442.600 91.400 443.800 118.600 ;
        RECT 445.800 71.400 447.000 112.600 ;
        RECT 449.000 91.400 450.200 152.600 ;
        RECT 468.200 125.400 469.400 190.600 ;
        RECT 481.000 149.400 482.200 194.600 ;
        RECT 484.200 97.400 485.400 168.600 ;
        RECT 503.400 135.400 504.600 172.600 ;
        RECT 506.600 135.400 507.800 196.600 ;
        RECT 509.800 123.400 511.000 192.600 ;
        RECT 519.400 127.400 520.600 182.600 ;
        RECT 522.600 143.400 523.800 184.600 ;
        RECT 503.400 113.400 504.600 122.600 ;
        RECT 506.600 97.400 507.800 122.600 ;
        RECT 465.000 55.400 466.200 82.600 ;
        RECT 541.800 73.400 543.000 118.600 ;
        RECT 503.400 9.400 504.600 40.600 ;
        RECT 516.200 33.400 517.400 68.600 ;
        RECT 545.000 13.400 546.200 476.600 ;
        RECT 561.000 423.400 562.200 534.600 ;
        RECT 573.800 387.400 575.000 442.600 ;
        RECT 554.600 291.400 555.800 332.600 ;
        RECT 557.800 273.400 559.000 322.600 ;
        RECT 583.400 313.400 584.600 460.600 ;
        RECT 589.800 451.400 591.000 530.600 ;
        RECT 589.800 371.400 591.000 414.600 ;
        RECT 548.200 231.400 549.400 266.600 ;
        RECT 551.400 9.400 552.600 244.600 ;
        RECT 564.200 167.400 565.400 210.600 ;
        RECT 567.400 107.400 568.600 204.600 ;
        RECT 573.800 185.400 575.000 238.600 ;
        RECT 580.200 181.400 581.400 294.600 ;
        RECT 586.600 237.400 587.800 314.600 ;
        RECT 593.000 293.400 594.200 452.600 ;
        RECT 599.400 399.400 600.600 526.600 ;
        RECT 602.600 267.400 603.800 484.600 ;
        RECT 570.600 109.400 571.800 144.600 ;
        RECT 554.600 51.400 555.800 70.600 ;
        RECT 570.600 33.400 571.800 104.600 ;
        RECT 580.200 45.400 581.400 176.600 ;
        RECT 586.600 147.400 587.800 232.600 ;
        RECT 583.400 11.400 584.600 120.600 ;
        RECT 589.800 117.400 591.000 198.600 ;
        RECT 586.600 67.400 587.800 98.600 ;
        RECT 596.200 97.400 597.400 160.600 ;
        RECT 602.600 133.400 603.800 230.600 ;
        RECT 602.600 97.400 603.800 118.600 ;
        RECT 609.000 41.400 610.200 188.600 ;
  END
END noc_top
END LIBRARY


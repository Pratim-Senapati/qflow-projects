magic
tech scmos
magscale 1 2
timestamp 1740382396
<< metal1 >>
rect 584 2006 590 2014
rect 598 2006 604 2014
rect 612 2006 618 2014
rect 626 2006 632 2014
rect 356 1916 364 1924
rect 381 1904 387 1923
rect 1508 1916 1512 1924
rect 52 1897 67 1903
rect 189 1897 220 1903
rect 61 1877 67 1897
rect 276 1897 355 1903
rect 388 1897 403 1903
rect 1460 1897 1475 1903
rect 157 1877 179 1883
rect 173 1864 179 1877
rect 317 1877 339 1883
rect 317 1863 323 1877
rect 520 1876 524 1884
rect 1469 1877 1475 1897
rect 1693 1897 1708 1903
rect 1725 1877 1763 1883
rect 301 1857 323 1863
rect 1560 1806 1566 1814
rect 1574 1806 1580 1814
rect 1588 1806 1594 1814
rect 1602 1806 1608 1814
rect 1642 1776 1644 1784
rect 1956 1776 1960 1784
rect 605 1757 675 1763
rect 605 1743 611 1757
rect 1869 1757 1891 1763
rect 589 1737 611 1743
rect 1533 1737 1619 1743
rect 580 1717 700 1723
rect 1773 1723 1779 1743
rect 1853 1737 1868 1743
rect 1773 1717 1843 1723
rect 2076 1723 2084 1728
rect 2076 1717 2099 1723
rect 500 1677 515 1683
rect 1476 1676 1480 1684
rect 2173 1677 2188 1683
rect 1716 1636 1720 1644
rect 584 1606 590 1614
rect 598 1606 604 1614
rect 612 1606 618 1614
rect 626 1606 632 1614
rect 1636 1537 1700 1543
rect 1692 1532 1700 1537
rect 157 1517 179 1523
rect 125 1497 140 1503
rect 269 1503 275 1523
rect 349 1503 355 1516
rect 269 1497 307 1503
rect 317 1497 355 1503
rect 2062 1497 2099 1503
rect 216 1477 243 1483
rect 333 1477 348 1483
rect 2173 1477 2188 1483
rect 1706 1436 1708 1444
rect 1560 1406 1566 1414
rect 1574 1406 1580 1414
rect 1588 1406 1594 1414
rect 1602 1406 1608 1414
rect 2004 1376 2008 1384
rect 372 1357 387 1363
rect 1917 1357 1932 1363
rect 388 1337 403 1343
rect 596 1337 674 1343
rect 1188 1337 1203 1343
rect 1213 1337 1228 1343
rect 1693 1337 1747 1343
rect 1693 1323 1699 1337
rect 1684 1317 1699 1323
rect 1837 1323 1843 1336
rect 1837 1317 1859 1323
rect 2116 1317 2131 1323
rect 440 1298 444 1306
rect 2157 1277 2188 1283
rect 1044 1236 1048 1244
rect 1780 1236 1784 1244
rect 584 1206 590 1214
rect 598 1206 604 1214
rect 612 1206 618 1214
rect 626 1206 632 1214
rect 381 1097 396 1103
rect 444 1103 452 1104
rect 444 1097 483 1103
rect 2078 1097 2115 1103
rect 509 1077 588 1083
rect 1325 1077 1340 1083
rect 2141 1077 2188 1083
rect 948 1057 963 1063
rect 328 1036 332 1044
rect 1560 1006 1566 1014
rect 1574 1006 1580 1014
rect 1588 1006 1594 1014
rect 1602 1006 1608 1014
rect 888 976 892 984
rect 2084 976 2088 984
rect 925 937 940 943
rect 989 937 1004 943
rect 1053 937 1084 943
rect 1806 937 1836 943
rect 1933 937 1971 943
rect 1828 917 1875 923
rect 989 897 1004 903
rect 1069 897 1084 903
rect 1021 877 1036 883
rect 584 806 590 814
rect 598 806 604 814
rect 612 806 618 814
rect 626 806 632 814
rect 2052 776 2054 784
rect 308 737 323 743
rect 1060 737 1075 743
rect 413 697 508 703
rect 1108 697 1123 703
rect 2061 697 2083 703
rect 116 677 147 683
rect 285 677 307 683
rect 445 677 530 683
rect 1332 677 1347 683
rect 2141 677 2188 683
rect 141 657 156 663
rect 1524 657 1603 663
rect 2013 657 2028 663
rect 1780 636 1784 644
rect 1560 606 1566 614
rect 1574 606 1580 614
rect 1588 606 1594 614
rect 1602 606 1608 614
rect 824 576 828 584
rect 1604 577 1628 583
rect 372 537 387 543
rect 637 543 643 563
rect 740 557 755 563
rect 941 557 963 563
rect 564 537 643 543
rect 957 543 963 557
rect 1101 557 1116 563
rect 1565 557 1628 563
rect 957 537 979 543
rect 2077 537 2108 543
rect 548 517 675 523
rect 916 517 995 523
rect 1005 517 1036 523
rect 1181 517 1196 523
rect 429 497 451 503
rect 765 497 787 503
rect 2044 484 2052 488
rect 1044 477 1059 483
rect 584 406 590 414
rect 598 406 604 414
rect 612 406 618 414
rect 626 406 632 414
rect 324 376 326 384
rect 141 317 163 323
rect 285 297 300 303
rect 173 277 188 283
rect 173 257 179 277
rect 285 277 291 297
rect 349 303 355 316
rect 308 297 323 303
rect 349 297 387 303
rect 381 283 387 297
rect 680 297 716 303
rect 1469 303 1475 316
rect 1469 297 1491 303
rect 1597 297 1619 303
rect 2116 297 2124 303
rect 381 277 403 283
rect 564 277 627 283
rect 1501 277 1564 283
rect 2109 277 2115 296
rect 2157 277 2188 283
rect 248 236 252 244
rect 557 237 604 243
rect 2052 236 2056 244
rect 1560 206 1566 214
rect 1574 206 1580 214
rect 1588 206 1594 214
rect 1602 206 1608 214
rect 516 157 531 163
rect 1444 157 1475 163
rect 45 117 82 123
rect 445 117 530 123
rect 584 6 590 14
rect 598 6 604 14
rect 612 6 618 14
rect 626 6 632 14
<< m2contact >>
rect 590 2006 598 2014
rect 604 2006 612 2014
rect 618 2006 626 2014
rect 428 1976 436 1984
rect 972 1976 980 1984
rect 1052 1976 1060 1984
rect 1420 1976 1428 1984
rect 1660 1976 1668 1984
rect 1132 1958 1140 1966
rect 1884 1958 1892 1966
rect 508 1936 516 1944
rect 540 1936 548 1944
rect 348 1916 356 1924
rect 476 1916 484 1924
rect 604 1916 612 1924
rect 972 1916 980 1924
rect 1132 1912 1140 1920
rect 1500 1916 1508 1924
rect 1884 1912 1892 1920
rect 44 1896 52 1904
rect 12 1876 20 1884
rect 220 1896 228 1904
rect 268 1896 276 1904
rect 380 1896 388 1904
rect 492 1896 500 1904
rect 682 1896 690 1904
rect 972 1896 980 1904
rect 1020 1896 1028 1904
rect 1100 1896 1108 1904
rect 1390 1896 1398 1904
rect 1452 1896 1460 1904
rect 284 1876 292 1884
rect 172 1856 180 1864
rect 284 1856 292 1864
rect 460 1876 468 1884
rect 524 1876 532 1884
rect 572 1876 580 1884
rect 588 1876 596 1884
rect 876 1876 884 1884
rect 1196 1876 1204 1884
rect 1628 1896 1636 1904
rect 1708 1896 1716 1904
rect 1740 1896 1748 1904
rect 1852 1896 1860 1904
rect 1564 1876 1572 1884
rect 1772 1880 1780 1888
rect 1948 1876 1956 1884
rect 444 1856 452 1864
rect 556 1856 564 1864
rect 844 1856 852 1864
rect 1228 1856 1236 1864
rect 1676 1856 1684 1864
rect 1708 1856 1716 1864
rect 1980 1856 1988 1864
rect 108 1836 116 1844
rect 284 1836 292 1844
rect 1724 1836 1732 1844
rect 1804 1836 1812 1844
rect 2140 1836 2148 1844
rect 1566 1806 1574 1814
rect 1580 1806 1588 1814
rect 1594 1806 1602 1814
rect 28 1776 36 1784
rect 364 1776 372 1784
rect 684 1776 692 1784
rect 908 1776 916 1784
rect 1612 1776 1620 1784
rect 1644 1776 1652 1784
rect 1948 1776 1956 1784
rect 2028 1776 2036 1784
rect 188 1756 196 1764
rect 492 1756 500 1764
rect 524 1756 532 1764
rect 220 1736 228 1744
rect 684 1756 692 1764
rect 1196 1756 1204 1764
rect 1356 1756 1364 1764
rect 1596 1756 1604 1764
rect 1900 1756 1908 1764
rect 684 1736 692 1744
rect 780 1736 788 1744
rect 876 1736 884 1744
rect 1020 1736 1028 1744
rect 1164 1736 1172 1744
rect 1436 1736 1444 1744
rect 1660 1736 1668 1744
rect 1676 1736 1684 1744
rect 108 1716 116 1724
rect 396 1716 404 1724
rect 444 1716 452 1724
rect 476 1716 484 1724
rect 556 1716 564 1724
rect 572 1716 580 1724
rect 700 1716 708 1724
rect 1100 1716 1108 1724
rect 1420 1716 1428 1724
rect 1788 1736 1796 1744
rect 1868 1736 1876 1744
rect 1916 1736 1924 1744
rect 2012 1736 2020 1744
rect 2076 1736 2084 1744
rect 2124 1736 2132 1744
rect 2060 1716 2068 1724
rect 2140 1716 2148 1724
rect 316 1696 324 1704
rect 460 1696 468 1704
rect 540 1696 548 1704
rect 1068 1696 1076 1704
rect 1628 1696 1636 1704
rect 1820 1696 1828 1704
rect 428 1676 436 1684
rect 492 1676 500 1684
rect 1468 1676 1476 1684
rect 2188 1676 2196 1684
rect 108 1654 116 1662
rect 412 1636 420 1644
rect 828 1636 836 1644
rect 1068 1636 1076 1644
rect 1388 1636 1396 1644
rect 1708 1636 1716 1644
rect 590 1606 598 1614
rect 604 1606 612 1614
rect 618 1606 626 1614
rect 716 1576 724 1584
rect 1116 1576 1124 1584
rect 1612 1576 1620 1584
rect 60 1556 68 1564
rect 524 1556 532 1564
rect 924 1556 932 1564
rect 1356 1558 1364 1566
rect 1804 1558 1812 1566
rect 12 1536 20 1544
rect 204 1536 212 1544
rect 1628 1536 1636 1544
rect 2124 1536 2132 1544
rect 44 1496 52 1504
rect 92 1496 100 1504
rect 140 1496 148 1504
rect 188 1496 196 1504
rect 284 1516 292 1524
rect 348 1516 356 1524
rect 460 1512 468 1520
rect 860 1512 868 1520
rect 1356 1512 1364 1520
rect 1692 1516 1700 1524
rect 1804 1512 1812 1520
rect 524 1496 532 1504
rect 924 1496 932 1504
rect 1324 1496 1332 1504
rect 1532 1496 1540 1504
rect 1772 1496 1780 1504
rect 2140 1496 2148 1504
rect 348 1476 356 1484
rect 364 1476 372 1484
rect 380 1476 388 1484
rect 524 1476 532 1484
rect 924 1476 932 1484
rect 1148 1476 1156 1484
rect 1276 1476 1284 1484
rect 1420 1476 1428 1484
rect 1724 1476 1732 1484
rect 1868 1476 1876 1484
rect 2188 1476 2196 1484
rect 108 1456 116 1464
rect 140 1456 148 1464
rect 252 1456 260 1464
rect 556 1456 564 1464
rect 956 1456 964 1464
rect 1452 1456 1460 1464
rect 1900 1456 1908 1464
rect 204 1436 212 1444
rect 1708 1436 1716 1444
rect 2060 1436 2068 1444
rect 1566 1406 1574 1414
rect 1580 1406 1588 1414
rect 1594 1406 1602 1414
rect 28 1376 36 1384
rect 1132 1376 1140 1384
rect 1996 1376 2004 1384
rect 2076 1376 2084 1384
rect 188 1356 196 1364
rect 364 1356 372 1364
rect 828 1356 836 1364
rect 1500 1356 1508 1364
rect 1884 1356 1892 1364
rect 1932 1356 1940 1364
rect 220 1336 228 1344
rect 380 1336 388 1344
rect 492 1336 500 1344
rect 588 1336 596 1344
rect 860 1336 868 1344
rect 1004 1336 1012 1344
rect 1100 1336 1108 1344
rect 1180 1336 1188 1344
rect 1228 1336 1236 1344
rect 1324 1336 1332 1344
rect 1468 1336 1476 1344
rect 1662 1336 1670 1344
rect 316 1316 324 1324
rect 412 1316 420 1324
rect 748 1316 756 1324
rect 1164 1316 1172 1324
rect 1276 1316 1284 1324
rect 1372 1316 1380 1324
rect 1676 1316 1684 1324
rect 1836 1336 1844 1344
rect 1964 1336 1972 1344
rect 2060 1336 2068 1344
rect 2108 1336 2116 1344
rect 1932 1316 1940 1324
rect 2108 1316 2116 1324
rect 316 1296 324 1304
rect 444 1298 452 1306
rect 924 1300 932 1308
rect 1180 1296 1188 1304
rect 1404 1300 1412 1308
rect 1948 1296 1956 1304
rect 2076 1296 2084 1304
rect 540 1276 548 1284
rect 1852 1276 1860 1284
rect 1916 1276 1924 1284
rect 2188 1276 2196 1284
rect 748 1254 756 1262
rect 1404 1254 1412 1262
rect 316 1236 324 1244
rect 1036 1236 1044 1244
rect 1772 1236 1780 1244
rect 590 1206 598 1214
rect 604 1206 612 1214
rect 618 1206 626 1214
rect 60 1176 68 1184
rect 348 1176 356 1184
rect 604 1176 612 1184
rect 892 1176 900 1184
rect 1388 1176 1396 1184
rect 1676 1176 1684 1184
rect 1788 1176 1796 1184
rect 1212 1158 1220 1166
rect 12 1136 20 1144
rect 316 1136 324 1144
rect 236 1116 244 1124
rect 284 1116 292 1124
rect 892 1116 900 1124
rect 1212 1112 1220 1120
rect 1388 1116 1396 1124
rect 1788 1116 1796 1124
rect 44 1096 52 1104
rect 92 1096 100 1104
rect 268 1096 276 1104
rect 300 1096 308 1104
rect 396 1096 404 1104
rect 684 1096 692 1104
rect 908 1096 916 1104
rect 1244 1096 1252 1104
rect 1292 1096 1300 1104
rect 1388 1096 1396 1104
rect 1596 1096 1604 1104
rect 1788 1096 1796 1104
rect 108 1076 116 1084
rect 204 1076 212 1084
rect 460 1076 468 1084
rect 588 1076 596 1084
rect 796 1076 804 1084
rect 1148 1076 1156 1084
rect 1340 1076 1348 1084
rect 1484 1076 1492 1084
rect 1884 1076 1892 1084
rect 2188 1076 2196 1084
rect 220 1056 228 1064
rect 252 1056 260 1064
rect 764 1056 772 1064
rect 940 1056 948 1064
rect 1116 1056 1124 1064
rect 1516 1056 1524 1064
rect 1916 1056 1924 1064
rect 156 1036 164 1044
rect 332 1036 340 1044
rect 444 1036 452 1044
rect 2076 1036 2084 1044
rect 1566 1006 1574 1014
rect 1580 1006 1588 1014
rect 1594 1006 1602 1014
rect 28 976 36 984
rect 380 976 388 984
rect 892 976 900 984
rect 2076 976 2084 984
rect 188 956 196 964
rect 540 956 548 964
rect 1004 956 1012 964
rect 1260 956 1268 964
rect 1644 956 1652 964
rect 220 936 228 944
rect 572 936 580 944
rect 828 936 836 944
rect 940 936 948 944
rect 1004 936 1012 944
rect 1036 936 1044 944
rect 1084 936 1092 944
rect 1292 936 1300 944
rect 1612 936 1620 944
rect 1836 936 1844 944
rect 1980 936 1988 944
rect 2028 936 2036 944
rect 2044 936 2052 944
rect 2140 936 2148 944
rect 108 916 116 924
rect 460 916 468 924
rect 812 916 820 924
rect 956 916 964 924
rect 1388 916 1396 924
rect 1516 916 1524 924
rect 1820 916 1828 924
rect 2156 916 2164 924
rect 316 896 324 904
rect 668 896 676 904
rect 1004 896 1012 904
rect 1084 896 1092 904
rect 1100 896 1108 904
rect 1356 900 1364 908
rect 1516 896 1524 904
rect 1948 896 1956 904
rect 1996 896 2004 904
rect 1036 876 1044 884
rect 2188 876 2196 884
rect 108 854 116 862
rect 460 854 468 862
rect 28 836 36 844
rect 380 836 388 844
rect 780 836 788 844
rect 1356 836 1364 844
rect 1516 836 1524 844
rect 2012 836 2020 844
rect 590 806 598 814
rect 604 806 612 814
rect 618 806 626 814
rect 1084 776 1092 784
rect 1148 776 1156 784
rect 1452 776 1460 784
rect 1916 776 1924 784
rect 2044 776 2052 784
rect 716 756 724 764
rect 12 736 20 744
rect 300 736 308 744
rect 1052 736 1060 744
rect 1724 736 1732 744
rect 284 716 292 724
rect 332 716 340 724
rect 780 712 788 720
rect 1036 716 1044 724
rect 1996 716 2004 724
rect 44 696 52 704
rect 92 696 100 704
rect 156 696 164 704
rect 252 696 260 704
rect 508 696 516 704
rect 716 696 724 704
rect 1052 696 1060 704
rect 1100 696 1108 704
rect 1276 696 1284 704
rect 1516 696 1524 704
rect 1580 696 1588 704
rect 1644 696 1652 704
rect 1676 696 1684 704
rect 1692 696 1700 704
rect 1868 696 1876 704
rect 1900 696 1908 704
rect 1948 696 1956 704
rect 1980 696 1988 704
rect 2108 696 2116 704
rect 60 676 68 684
rect 108 676 116 684
rect 236 676 244 684
rect 348 676 356 684
rect 716 676 724 684
rect 892 676 900 684
rect 1020 676 1028 684
rect 1260 676 1268 684
rect 1324 676 1332 684
rect 1628 676 1636 684
rect 1740 676 1748 684
rect 1836 676 1844 684
rect 1852 676 1860 684
rect 1964 676 1972 684
rect 2188 676 2196 684
rect 156 656 164 664
rect 684 656 692 664
rect 876 656 884 664
rect 1100 656 1108 664
rect 1484 656 1492 664
rect 1516 656 1524 664
rect 1612 656 1620 664
rect 2028 656 2036 664
rect 2092 656 2100 664
rect 140 636 148 644
rect 524 636 532 644
rect 860 636 868 644
rect 1308 636 1316 644
rect 1500 636 1508 644
rect 1772 636 1780 644
rect 2044 636 2052 644
rect 1566 606 1574 614
rect 1580 606 1588 614
rect 1594 606 1602 614
rect 828 576 836 584
rect 924 576 932 584
rect 1596 576 1604 584
rect 1628 576 1636 584
rect 2044 576 2052 584
rect 188 556 196 564
rect 412 556 420 564
rect 220 536 228 544
rect 364 536 372 544
rect 396 536 404 544
rect 556 536 564 544
rect 732 556 740 564
rect 924 556 932 564
rect 652 536 660 544
rect 924 536 932 544
rect 1084 556 1092 564
rect 1116 556 1124 564
rect 1196 556 1204 564
rect 1404 556 1412 564
rect 1628 556 1636 564
rect 1804 556 1812 564
rect 2028 556 2036 564
rect 2124 556 2132 564
rect 2140 556 2148 564
rect 1036 536 1044 544
rect 1132 536 1140 544
rect 1372 536 1380 544
rect 1772 536 1780 544
rect 2012 536 2020 544
rect 2108 536 2116 544
rect 108 516 116 524
rect 460 516 468 524
rect 524 516 532 524
rect 540 516 548 524
rect 796 516 804 524
rect 908 516 916 524
rect 1036 516 1044 524
rect 1116 516 1124 524
rect 1148 516 1156 524
rect 1196 516 1204 524
rect 1228 516 1236 524
rect 1308 516 1316 524
rect 1484 516 1492 524
rect 1676 516 1684 524
rect 1708 516 1716 524
rect 1996 516 2004 524
rect 2092 516 2100 524
rect 2156 516 2164 524
rect 316 496 324 504
rect 364 496 372 504
rect 1020 496 1028 504
rect 1068 496 1076 504
rect 1276 496 1284 504
rect 1676 496 1684 504
rect 476 476 484 484
rect 508 476 516 484
rect 716 476 724 484
rect 812 476 820 484
rect 1036 476 1044 484
rect 1964 476 1972 484
rect 2044 476 2052 484
rect 2188 476 2196 484
rect 108 454 116 462
rect 28 436 36 444
rect 492 436 500 444
rect 1228 436 1236 444
rect 1276 436 1284 444
rect 1676 436 1684 444
rect 590 406 598 414
rect 604 406 612 414
rect 618 406 626 414
rect 124 376 132 384
rect 316 376 324 384
rect 460 376 468 384
rect 492 376 500 384
rect 1052 376 1060 384
rect 1100 376 1108 384
rect 1596 376 1604 384
rect 1980 376 1988 384
rect 796 358 804 366
rect 1180 358 1188 366
rect 1724 358 1732 366
rect 12 336 20 344
rect 108 336 116 344
rect 348 316 356 324
rect 556 316 564 324
rect 44 296 52 304
rect 76 296 84 304
rect 124 296 132 304
rect 60 256 68 264
rect 188 276 196 284
rect 300 296 308 304
rect 796 312 804 320
rect 1356 312 1364 320
rect 1388 316 1396 324
rect 1468 316 1476 324
rect 300 276 308 284
rect 412 296 420 304
rect 716 296 724 304
rect 780 296 788 304
rect 1180 296 1188 304
rect 1724 312 1732 320
rect 1708 296 1716 304
rect 2108 296 2116 304
rect 2124 296 2132 304
rect 524 276 532 284
rect 556 276 564 284
rect 716 276 724 284
rect 860 276 868 284
rect 1292 276 1300 284
rect 1436 276 1444 284
rect 1564 276 1572 284
rect 1788 276 1796 284
rect 2012 276 2020 284
rect 2188 276 2196 284
rect 380 256 388 264
rect 508 256 516 264
rect 892 256 900 264
rect 1260 256 1268 264
rect 1516 256 1524 264
rect 1580 256 1588 264
rect 1644 256 1652 264
rect 1820 256 1828 264
rect 252 236 260 244
rect 604 236 612 244
rect 1100 236 1108 244
rect 1468 236 1476 244
rect 1628 236 1636 244
rect 2044 236 2052 244
rect 1566 206 1574 214
rect 1580 206 1588 214
rect 1594 206 1602 214
rect 76 176 84 184
rect 1068 176 1076 184
rect 2124 176 2132 184
rect 236 156 244 164
rect 508 156 516 164
rect 684 156 692 164
rect 1228 156 1236 164
rect 1436 156 1444 164
rect 1628 156 1636 164
rect 1964 156 1972 164
rect 268 136 276 144
rect 716 136 724 144
rect 1260 136 1268 144
rect 1660 136 1668 144
rect 1932 136 1940 144
rect 332 116 340 124
rect 604 116 612 124
rect 780 116 788 124
rect 892 116 900 124
rect 908 116 916 124
rect 956 116 964 124
rect 1004 116 1012 124
rect 1356 116 1364 124
rect 1740 116 1748 124
rect 1836 116 1844 124
rect 364 96 372 104
rect 812 96 820 104
rect 1356 96 1364 104
rect 1724 100 1732 108
rect 1868 100 1876 108
rect 12 76 20 84
rect 364 36 372 44
rect 412 36 420 44
rect 812 36 820 44
rect 860 36 868 44
rect 940 36 948 44
rect 988 36 996 44
rect 1036 36 1044 44
rect 1356 36 1364 44
rect 1724 36 1732 44
rect 1868 36 1876 44
rect 590 6 598 14
rect 604 6 612 14
rect 618 6 626 14
<< metal2 >>
rect 365 2037 387 2043
rect 413 2037 435 2043
rect 1021 2037 1043 2043
rect 13 1884 19 1896
rect 45 1864 51 1896
rect 45 1803 51 1856
rect 173 1824 179 1856
rect 29 1797 51 1803
rect 29 1784 35 1797
rect 109 1662 115 1716
rect 13 1524 19 1536
rect 189 1523 195 1756
rect 221 1744 227 1836
rect 285 1684 291 1836
rect 365 1784 371 2037
rect 429 1984 435 2037
rect 584 2006 590 2014
rect 598 2006 604 2014
rect 612 2006 618 2014
rect 626 2006 632 2014
rect 973 1924 979 1976
rect 381 1884 387 1896
rect 477 1864 483 1916
rect 493 1884 499 1896
rect 557 1864 563 1896
rect 397 1724 403 1756
rect 493 1704 499 1756
rect 573 1724 579 1876
rect 845 1824 851 1856
rect 909 1784 915 1816
rect 669 1777 684 1783
rect 189 1517 211 1523
rect 45 1464 51 1496
rect 93 1484 99 1496
rect 205 1483 211 1517
rect 189 1477 211 1483
rect 141 1464 147 1476
rect 29 1457 44 1463
rect 29 1384 35 1457
rect 189 1384 195 1477
rect 285 1464 291 1516
rect 253 1444 259 1456
rect 189 1364 195 1376
rect 221 1344 227 1436
rect 317 1324 323 1696
rect 461 1684 467 1696
rect 413 1524 419 1636
rect 381 1484 387 1496
rect 349 1463 355 1476
rect 349 1457 371 1463
rect 365 1364 371 1457
rect 381 1344 387 1456
rect 413 1344 419 1516
rect 413 1324 419 1336
rect 461 1324 467 1512
rect 525 1504 531 1556
rect 557 1504 563 1716
rect 584 1606 590 1614
rect 598 1606 604 1614
rect 612 1606 618 1614
rect 626 1606 632 1614
rect 669 1544 675 1777
rect 877 1744 883 1756
rect 685 1704 691 1736
rect 701 1724 707 1736
rect 717 1584 723 1696
rect 829 1484 835 1636
rect 557 1384 563 1456
rect 829 1364 835 1456
rect 861 1424 867 1512
rect 925 1504 931 1556
rect 957 1464 963 1816
rect 1021 1764 1027 1896
rect 1037 1743 1043 2037
rect 1053 1984 1059 2043
rect 1421 2037 1443 2043
rect 1645 2037 1667 2043
rect 1677 2037 1683 2043
rect 1725 2037 1731 2043
rect 2013 2037 2019 2043
rect 1421 1984 1427 2037
rect 1661 1984 1667 2037
rect 1133 1920 1139 1958
rect 1885 1920 1891 1958
rect 1028 1737 1043 1743
rect 1021 1644 1027 1736
rect 1069 1644 1075 1696
rect 1085 1584 1091 1756
rect 1101 1724 1107 1896
rect 1197 1884 1203 1916
rect 1197 1764 1203 1856
rect 1560 1806 1566 1814
rect 1574 1806 1580 1814
rect 1588 1806 1594 1814
rect 1602 1806 1608 1814
rect 1629 1764 1635 1896
rect 1645 1784 1651 1876
rect 1677 1864 1683 1896
rect 1709 1784 1715 1856
rect 1725 1804 1731 1836
rect 1773 1824 1779 1880
rect 1101 1484 1107 1716
rect 1165 1704 1171 1736
rect 1149 1484 1155 1636
rect 589 1344 595 1356
rect 317 1244 323 1296
rect 349 1184 355 1216
rect 93 1104 99 1176
rect 445 1144 451 1298
rect 461 1104 467 1316
rect 749 1262 755 1316
rect 861 1284 867 1336
rect 925 1308 931 1416
rect 957 1364 963 1456
rect 1133 1384 1139 1476
rect 1149 1424 1155 1476
rect 1197 1464 1203 1756
rect 1661 1744 1667 1756
rect 1677 1744 1683 1756
rect 1789 1744 1795 1796
rect 1629 1704 1635 1736
rect 1469 1684 1475 1696
rect 1389 1604 1395 1636
rect 1357 1520 1363 1558
rect 1629 1544 1635 1696
rect 1677 1584 1683 1736
rect 1325 1484 1331 1496
rect 1277 1464 1283 1476
rect 1453 1404 1459 1456
rect 1560 1406 1566 1414
rect 1574 1406 1580 1414
rect 1588 1406 1594 1414
rect 1602 1406 1608 1414
rect 1501 1364 1507 1396
rect 925 1223 931 1300
rect 909 1217 931 1223
rect 584 1206 590 1214
rect 598 1206 604 1214
rect 612 1206 618 1214
rect 626 1206 632 1214
rect 893 1124 899 1176
rect 909 1104 915 1217
rect 1005 1184 1011 1336
rect 1165 1284 1171 1316
rect 1325 1304 1331 1336
rect 1469 1324 1475 1336
rect 1037 1104 1043 1236
rect 1213 1120 1219 1158
rect 1293 1104 1299 1276
rect 1373 1104 1379 1316
rect 1405 1262 1411 1300
rect 1677 1284 1683 1316
rect 1677 1184 1683 1276
rect 1693 1204 1699 1516
rect 1709 1484 1715 1636
rect 1725 1484 1731 1596
rect 1773 1504 1779 1716
rect 1805 1604 1811 1836
rect 1853 1724 1859 1896
rect 1949 1784 1955 1876
rect 1981 1844 1987 1856
rect 2029 1784 2035 1816
rect 2077 1744 2083 1756
rect 2013 1724 2019 1736
rect 2141 1724 2147 1836
rect 2189 1684 2195 1696
rect 1805 1520 1811 1558
rect 1709 1364 1715 1436
rect 1725 1324 1731 1476
rect 1997 1384 2003 1476
rect 1885 1364 1891 1376
rect 1837 1344 1843 1356
rect 1965 1344 1971 1356
rect 2061 1344 2067 1436
rect 2141 1344 2147 1496
rect 2189 1484 2195 1496
rect 2068 1337 2083 1343
rect 2077 1304 2083 1337
rect 2109 1324 2115 1336
rect 1853 1284 1859 1296
rect 1949 1284 1955 1296
rect 2109 1284 2115 1316
rect 2189 1284 2195 1296
rect 1389 1124 1395 1176
rect 29 1097 44 1103
rect 29 984 35 1097
rect 45 1084 51 1096
rect 205 1024 211 1076
rect 221 1064 227 1076
rect 109 862 115 916
rect 29 684 35 836
rect 45 704 51 716
rect 61 684 67 696
rect 93 564 99 696
rect 109 684 115 716
rect 157 664 163 676
rect 189 664 195 956
rect 221 944 227 1036
rect 253 1024 259 1056
rect 301 744 307 936
rect 141 604 147 636
rect 189 564 195 656
rect 109 462 115 516
rect 29 323 35 436
rect 125 384 131 416
rect 29 317 44 323
rect 45 304 51 316
rect 301 304 307 516
rect 317 504 323 896
rect 333 724 339 1036
rect 381 984 387 1016
rect 397 964 403 1096
rect 589 1084 595 1096
rect 797 1084 803 1096
rect 1245 1084 1251 1096
rect 1341 1084 1347 1096
rect 445 844 451 1036
rect 541 964 547 1056
rect 893 984 899 1076
rect 941 964 947 1056
rect 1117 964 1123 1056
rect 461 862 467 916
rect 381 724 387 836
rect 333 524 339 716
rect 509 684 515 696
rect 324 497 339 503
rect 317 384 323 476
rect 52 297 67 303
rect 61 264 67 297
rect 77 184 83 276
rect 237 164 243 216
rect 253 203 259 236
rect 253 197 275 203
rect 269 144 275 197
rect 333 124 339 497
rect 349 424 355 676
rect 541 664 547 956
rect 941 944 947 956
rect 829 924 835 936
rect 781 844 787 896
rect 813 844 819 916
rect 584 806 590 814
rect 598 806 604 814
rect 612 806 618 814
rect 626 806 632 814
rect 717 704 723 756
rect 781 720 787 836
rect 525 564 531 636
rect 829 584 835 916
rect 893 664 899 676
rect 557 544 563 556
rect 397 524 403 536
rect 365 484 371 496
rect 397 424 403 516
rect 461 404 467 516
rect 509 484 515 536
rect 477 383 483 476
rect 493 424 499 436
rect 493 384 499 396
rect 468 377 483 383
rect 381 264 387 276
rect 509 264 515 476
rect 525 284 531 516
rect 557 424 563 496
rect 557 324 563 416
rect 584 406 590 414
rect 598 406 604 414
rect 612 406 618 414
rect 626 406 632 414
rect 557 284 563 316
rect 733 283 739 556
rect 829 544 835 576
rect 861 524 867 636
rect 877 524 883 656
rect 925 584 931 736
rect 1037 724 1043 876
rect 1085 784 1091 896
rect 1117 824 1123 956
rect 1389 924 1395 1096
rect 1773 1084 1779 1236
rect 1917 1204 1923 1276
rect 1789 1124 1795 1176
rect 2189 1084 2195 1096
rect 1517 1024 1523 1056
rect 1133 664 1139 896
rect 1357 844 1363 900
rect 1149 784 1155 816
rect 1277 704 1283 836
rect 1085 657 1100 663
rect 1085 564 1091 657
rect 925 524 931 536
rect 909 504 915 516
rect 1021 504 1027 516
rect 1037 504 1043 516
rect 797 320 803 358
rect 724 277 739 283
rect 509 164 515 256
rect 605 144 611 236
rect 685 164 691 216
rect 733 204 739 277
rect 781 124 787 296
rect 861 284 867 296
rect 1037 284 1043 476
rect 1053 384 1059 556
rect 893 124 899 196
rect 909 124 915 136
rect 1005 124 1011 176
rect 1085 124 1091 556
rect 1133 544 1139 656
rect 1309 524 1315 636
rect 1405 564 1411 816
rect 1453 784 1459 1016
rect 1517 964 1523 1016
rect 1560 1006 1566 1014
rect 1574 1006 1580 1014
rect 1588 1006 1594 1014
rect 1602 1006 1608 1014
rect 1645 964 1651 1036
rect 1885 1024 1891 1076
rect 1917 1044 1923 1056
rect 2029 944 2035 1036
rect 2077 984 2083 1016
rect 1821 924 1827 936
rect 1837 924 1843 936
rect 1997 904 2003 916
rect 2045 904 2051 936
rect 1517 844 1523 896
rect 1917 784 1923 876
rect 1949 704 1955 716
rect 2013 704 2019 836
rect 2045 784 2051 896
rect 2189 884 2195 896
rect 1517 684 1523 696
rect 1629 684 1635 696
rect 1101 384 1107 516
rect 1101 144 1107 236
rect 1117 184 1123 516
rect 1197 404 1203 516
rect 1277 444 1283 496
rect 1229 424 1235 436
rect 1309 384 1315 516
rect 1181 304 1187 358
rect 1357 320 1363 376
rect 1261 164 1267 256
rect 1389 124 1395 316
rect 1405 264 1411 556
rect 1501 544 1507 636
rect 1560 606 1566 614
rect 1574 606 1580 614
rect 1588 606 1594 614
rect 1602 606 1608 614
rect 1629 584 1635 676
rect 1645 664 1651 696
rect 1677 684 1683 696
rect 1837 684 1843 696
rect 1869 664 1875 696
rect 1901 684 1907 696
rect 2093 664 2099 676
rect 2109 664 2115 696
rect 2189 684 2195 696
rect 1469 324 1475 396
rect 1597 384 1603 576
rect 1645 563 1651 656
rect 1636 557 1651 563
rect 1677 444 1683 496
rect 1709 304 1715 516
rect 1805 383 1811 556
rect 1981 384 1987 656
rect 1997 524 2003 636
rect 2029 623 2035 656
rect 2029 617 2051 623
rect 2045 584 2051 617
rect 2093 524 2099 656
rect 1805 377 1827 383
rect 1725 320 1731 358
rect 1437 264 1443 276
rect 1565 264 1571 276
rect 1437 164 1443 256
rect 1581 244 1587 256
rect 1560 206 1566 214
rect 1574 206 1580 214
rect 1588 206 1594 214
rect 1602 206 1608 214
rect 1629 184 1635 236
rect 1709 204 1715 296
rect 1789 284 1795 376
rect 1821 264 1827 377
rect 2093 364 2099 516
rect 2013 284 2019 356
rect 2109 304 2115 536
rect 2141 484 2147 556
rect 2157 484 2163 516
rect 2189 484 2195 496
rect 1661 144 1667 176
rect 1741 124 1747 196
rect 1821 164 1827 256
rect 1837 124 1843 196
rect 2045 144 2051 236
rect 2125 184 2131 296
rect 2189 284 2195 296
rect 13 84 19 96
rect 365 44 371 96
rect 813 44 819 96
rect 1357 44 1363 96
rect 1725 44 1731 100
rect 1869 44 1875 100
rect 413 -17 419 36
rect 584 6 590 14
rect 598 6 604 14
rect 612 6 618 14
rect 626 6 632 14
rect 861 -17 867 36
rect 941 -17 947 36
rect 989 -17 995 36
rect 1037 -17 1043 36
rect 413 -23 435 -17
rect 477 -23 483 -17
rect 861 -23 883 -17
rect 925 -23 947 -17
rect 973 -23 995 -17
rect 1021 -23 1043 -17
rect 1405 -23 1411 16
rect 1453 -23 1459 -17
<< m3contact >>
rect 348 1916 356 1924
rect 12 1896 20 1904
rect 220 1896 228 1904
rect 268 1896 276 1904
rect 284 1876 292 1884
rect 44 1856 52 1864
rect 284 1856 292 1864
rect 108 1836 116 1844
rect 220 1836 228 1844
rect 172 1816 180 1824
rect 60 1556 68 1564
rect 12 1516 20 1524
rect 590 2006 598 2014
rect 604 2006 612 2014
rect 618 2006 626 2014
rect 508 1936 516 1944
rect 540 1936 548 1944
rect 604 1916 612 1924
rect 380 1896 388 1904
rect 380 1876 388 1884
rect 460 1876 468 1884
rect 556 1896 564 1904
rect 684 1896 690 1904
rect 690 1896 692 1904
rect 972 1896 980 1904
rect 492 1876 500 1884
rect 524 1876 532 1884
rect 572 1876 580 1884
rect 588 1876 596 1884
rect 876 1876 884 1884
rect 444 1856 452 1864
rect 476 1856 484 1864
rect 396 1756 404 1764
rect 492 1756 500 1764
rect 524 1756 532 1764
rect 444 1716 452 1724
rect 476 1716 484 1724
rect 844 1816 852 1824
rect 908 1816 916 1824
rect 956 1816 964 1824
rect 492 1696 500 1704
rect 540 1696 548 1704
rect 284 1676 292 1684
rect 204 1536 212 1544
rect 140 1496 148 1504
rect 188 1496 196 1504
rect 92 1476 100 1484
rect 140 1476 148 1484
rect 44 1456 52 1464
rect 108 1456 116 1464
rect 284 1456 292 1464
rect 204 1436 212 1444
rect 220 1436 228 1444
rect 252 1436 260 1444
rect 188 1376 196 1384
rect 428 1676 436 1684
rect 460 1676 468 1684
rect 492 1676 500 1684
rect 348 1516 356 1524
rect 412 1516 420 1524
rect 380 1496 388 1504
rect 348 1476 356 1484
rect 364 1476 372 1484
rect 380 1456 388 1464
rect 364 1356 372 1364
rect 412 1336 420 1344
rect 590 1606 598 1614
rect 604 1606 612 1614
rect 618 1606 626 1614
rect 684 1756 692 1764
rect 876 1756 884 1764
rect 700 1736 708 1744
rect 780 1736 788 1744
rect 684 1696 692 1704
rect 716 1696 724 1704
rect 668 1536 676 1544
rect 556 1496 564 1504
rect 524 1476 532 1484
rect 828 1476 836 1484
rect 556 1456 564 1464
rect 828 1456 836 1464
rect 556 1376 564 1384
rect 924 1476 932 1484
rect 1020 1756 1028 1764
rect 1196 1916 1204 1924
rect 1500 1916 1508 1924
rect 1100 1896 1108 1904
rect 1084 1756 1092 1764
rect 1020 1636 1028 1644
rect 1388 1896 1390 1904
rect 1390 1896 1396 1904
rect 1452 1896 1460 1904
rect 1676 1896 1684 1904
rect 1708 1896 1716 1904
rect 1740 1896 1748 1904
rect 1564 1876 1572 1884
rect 1196 1856 1204 1864
rect 1228 1856 1236 1864
rect 1566 1806 1574 1814
rect 1580 1806 1588 1814
rect 1594 1806 1602 1814
rect 1612 1776 1620 1784
rect 1644 1876 1652 1884
rect 1772 1816 1780 1824
rect 1724 1796 1732 1804
rect 1788 1796 1796 1804
rect 1708 1776 1716 1784
rect 1356 1756 1364 1764
rect 1596 1756 1604 1764
rect 1628 1756 1636 1764
rect 1660 1756 1668 1764
rect 1676 1756 1684 1764
rect 1084 1576 1092 1584
rect 1164 1696 1172 1704
rect 1148 1636 1156 1644
rect 1116 1576 1124 1584
rect 1100 1476 1108 1484
rect 1132 1476 1140 1484
rect 860 1416 868 1424
rect 924 1416 932 1424
rect 588 1356 596 1364
rect 828 1356 836 1364
rect 492 1336 500 1344
rect 316 1316 324 1324
rect 460 1316 468 1324
rect 348 1216 356 1224
rect 60 1176 68 1184
rect 92 1176 100 1184
rect 12 1136 20 1144
rect 316 1136 324 1144
rect 444 1136 452 1144
rect 236 1116 244 1124
rect 284 1116 292 1124
rect 540 1276 548 1284
rect 1436 1736 1444 1744
rect 1628 1736 1636 1744
rect 1420 1716 1428 1724
rect 1468 1696 1476 1704
rect 1628 1696 1636 1704
rect 1388 1596 1396 1604
rect 1612 1576 1620 1584
rect 1772 1716 1780 1724
rect 1676 1576 1684 1584
rect 1532 1496 1540 1504
rect 1324 1476 1332 1484
rect 1420 1476 1428 1484
rect 1196 1456 1204 1464
rect 1276 1456 1284 1464
rect 1452 1456 1460 1464
rect 1148 1416 1156 1424
rect 1566 1406 1574 1414
rect 1580 1406 1588 1414
rect 1594 1406 1602 1414
rect 1452 1396 1460 1404
rect 1500 1396 1508 1404
rect 956 1356 964 1364
rect 1100 1336 1108 1344
rect 1180 1336 1188 1344
rect 1228 1336 1236 1344
rect 1660 1336 1662 1344
rect 1662 1336 1668 1344
rect 860 1276 868 1284
rect 590 1206 598 1214
rect 604 1206 612 1214
rect 618 1206 626 1214
rect 604 1176 612 1184
rect 1276 1316 1284 1324
rect 1468 1316 1476 1324
rect 1180 1296 1188 1304
rect 1324 1296 1332 1304
rect 1164 1276 1172 1284
rect 1292 1276 1300 1284
rect 1004 1176 1012 1184
rect 1676 1276 1684 1284
rect 1724 1596 1732 1604
rect 1980 1836 1988 1844
rect 2028 1816 2036 1824
rect 1900 1756 1908 1764
rect 2076 1756 2084 1764
rect 1868 1736 1876 1744
rect 1916 1736 1924 1744
rect 2124 1736 2132 1744
rect 1852 1716 1860 1724
rect 2012 1716 2020 1724
rect 2060 1716 2068 1724
rect 2140 1716 2148 1724
rect 1820 1696 1828 1704
rect 2188 1696 2196 1704
rect 1804 1596 1812 1604
rect 2124 1536 2132 1544
rect 1772 1496 1780 1504
rect 2188 1496 2196 1504
rect 1708 1476 1716 1484
rect 1868 1476 1876 1484
rect 1996 1476 2004 1484
rect 1708 1356 1716 1364
rect 1900 1456 1908 1464
rect 1884 1376 1892 1384
rect 1836 1356 1844 1364
rect 1932 1356 1940 1364
rect 1964 1356 1972 1364
rect 2076 1376 2084 1384
rect 1724 1316 1732 1324
rect 1932 1316 1940 1324
rect 2140 1336 2148 1344
rect 1852 1296 1860 1304
rect 2188 1296 2196 1304
rect 1948 1276 1956 1284
rect 2108 1276 2116 1284
rect 1692 1196 1700 1204
rect 268 1096 276 1104
rect 300 1096 308 1104
rect 460 1096 468 1104
rect 588 1096 596 1104
rect 684 1096 692 1104
rect 796 1096 804 1104
rect 1036 1096 1044 1104
rect 1292 1096 1300 1104
rect 1340 1096 1348 1104
rect 1372 1096 1380 1104
rect 1388 1096 1396 1104
rect 1596 1096 1604 1104
rect 44 1076 52 1084
rect 108 1076 116 1084
rect 220 1076 228 1084
rect 156 1036 164 1044
rect 220 1036 228 1044
rect 204 1016 212 1024
rect 12 736 20 744
rect 44 716 52 724
rect 108 716 116 724
rect 60 696 68 704
rect 28 676 36 684
rect 156 696 164 704
rect 156 676 164 684
rect 252 1016 260 1024
rect 300 936 308 944
rect 316 896 324 904
rect 284 716 292 724
rect 252 696 260 704
rect 236 676 244 684
rect 188 656 196 664
rect 140 596 148 604
rect 92 556 100 564
rect 220 536 228 544
rect 300 516 308 524
rect 12 336 20 344
rect 124 416 132 424
rect 108 336 116 344
rect 44 316 52 324
rect 380 1016 388 1024
rect 460 1076 468 1084
rect 892 1076 900 1084
rect 1148 1076 1156 1084
rect 1244 1076 1252 1084
rect 1340 1076 1348 1084
rect 540 1056 548 1064
rect 764 1056 772 1064
rect 396 956 404 964
rect 940 956 948 964
rect 1004 956 1012 964
rect 1116 956 1124 964
rect 1260 956 1268 964
rect 444 836 452 844
rect 380 716 388 724
rect 508 676 516 684
rect 332 516 340 524
rect 316 476 324 484
rect 76 296 84 304
rect 124 296 132 304
rect 300 296 308 304
rect 76 276 84 284
rect 188 276 196 284
rect 300 276 308 284
rect 236 216 244 224
rect 572 936 580 944
rect 1004 936 1012 944
rect 1036 936 1044 944
rect 1084 936 1092 944
rect 828 916 836 924
rect 956 916 964 924
rect 668 896 676 904
rect 780 896 788 904
rect 812 836 820 844
rect 590 806 598 814
rect 604 806 612 814
rect 618 806 626 814
rect 716 676 724 684
rect 540 656 548 664
rect 684 656 692 664
rect 1004 896 1012 904
rect 1100 896 1108 904
rect 924 736 932 744
rect 892 656 900 664
rect 412 556 420 564
rect 524 556 532 564
rect 556 556 564 564
rect 732 556 740 564
rect 364 536 372 544
rect 508 536 516 544
rect 652 536 660 544
rect 396 516 404 524
rect 364 476 372 484
rect 348 416 356 424
rect 396 416 404 424
rect 540 516 548 524
rect 460 396 468 404
rect 492 416 500 424
rect 492 396 500 404
rect 348 316 356 324
rect 412 296 420 304
rect 380 276 388 284
rect 556 496 564 504
rect 716 476 724 484
rect 556 416 564 424
rect 590 406 598 414
rect 604 406 612 414
rect 618 406 626 414
rect 716 296 724 304
rect 828 536 836 544
rect 1292 936 1300 944
rect 1916 1196 1924 1204
rect 1788 1096 1796 1104
rect 2188 1096 2196 1104
rect 1484 1076 1492 1084
rect 1772 1076 1780 1084
rect 1644 1036 1652 1044
rect 1452 1016 1460 1024
rect 1516 1016 1524 1024
rect 1388 916 1396 924
rect 1132 896 1140 904
rect 1116 816 1124 824
rect 1052 736 1060 744
rect 1052 696 1060 704
rect 1100 696 1108 704
rect 1020 676 1028 684
rect 1276 836 1284 844
rect 1148 816 1156 824
rect 1404 816 1412 824
rect 1260 676 1268 684
rect 1324 676 1332 684
rect 1100 656 1108 664
rect 1132 656 1140 664
rect 924 556 932 564
rect 1052 556 1060 564
rect 1116 556 1124 564
rect 1036 536 1044 544
rect 796 516 804 524
rect 860 516 868 524
rect 876 516 884 524
rect 924 516 932 524
rect 1020 516 1028 524
rect 908 496 916 504
rect 1036 496 1044 504
rect 812 476 820 484
rect 860 296 868 304
rect 684 216 692 224
rect 732 196 740 204
rect 604 136 612 144
rect 716 136 724 144
rect 1068 496 1076 504
rect 1036 276 1044 284
rect 892 256 900 264
rect 892 196 900 204
rect 1004 176 1012 184
rect 1068 176 1076 184
rect 908 136 916 144
rect 1196 556 1204 564
rect 1566 1006 1574 1014
rect 1580 1006 1588 1014
rect 1594 1006 1602 1014
rect 1916 1036 1924 1044
rect 2028 1036 2036 1044
rect 2076 1036 2084 1044
rect 1884 1016 1892 1024
rect 1516 956 1524 964
rect 1644 956 1652 964
rect 2076 1016 2084 1024
rect 1612 936 1620 944
rect 1820 936 1828 944
rect 1980 936 1988 944
rect 2028 936 2036 944
rect 2140 936 2148 944
rect 1516 916 1524 924
rect 1836 916 1844 924
rect 1996 916 2004 924
rect 2156 916 2164 924
rect 1948 896 1956 904
rect 2044 896 2052 904
rect 2188 896 2196 904
rect 1916 876 1924 884
rect 1724 736 1732 744
rect 1948 716 1956 724
rect 1996 716 2004 724
rect 1580 696 1588 704
rect 1628 696 1636 704
rect 1644 696 1652 704
rect 1692 696 1700 704
rect 1836 696 1844 704
rect 1868 696 1876 704
rect 1980 696 1988 704
rect 2012 696 2020 704
rect 2188 696 2196 704
rect 1516 676 1524 684
rect 1484 656 1492 664
rect 1516 656 1524 664
rect 1612 656 1620 664
rect 1372 536 1380 544
rect 1100 516 1108 524
rect 1116 516 1124 524
rect 1148 516 1156 524
rect 1196 516 1204 524
rect 1228 516 1236 524
rect 1228 416 1236 424
rect 1196 396 1204 404
rect 1308 376 1316 384
rect 1356 376 1364 384
rect 1292 276 1300 284
rect 1260 256 1268 264
rect 1116 176 1124 184
rect 1228 156 1236 164
rect 1260 156 1268 164
rect 1100 136 1108 144
rect 1260 136 1268 144
rect 1566 606 1574 614
rect 1580 606 1588 614
rect 1594 606 1602 614
rect 1676 676 1684 684
rect 1740 676 1748 684
rect 1852 676 1860 684
rect 1900 676 1908 684
rect 1964 676 1972 684
rect 2092 676 2100 684
rect 1644 656 1652 664
rect 1868 656 1876 664
rect 1980 656 1988 664
rect 2108 656 2116 664
rect 1500 536 1508 544
rect 1484 516 1492 524
rect 1468 396 1476 404
rect 1772 636 1780 644
rect 1804 556 1812 564
rect 1772 536 1780 544
rect 1676 516 1684 524
rect 1788 376 1796 384
rect 1964 476 1972 484
rect 1996 636 2004 644
rect 2044 636 2052 644
rect 2028 556 2036 564
rect 2012 536 2020 544
rect 2124 556 2132 564
rect 2044 476 2052 484
rect 1404 256 1412 264
rect 1436 256 1444 264
rect 1516 256 1524 264
rect 1564 256 1572 264
rect 1644 256 1652 264
rect 1468 236 1476 244
rect 1580 236 1588 244
rect 1566 206 1574 214
rect 1580 206 1588 214
rect 1594 206 1602 214
rect 2012 356 2020 364
rect 2092 356 2100 364
rect 2188 496 2196 504
rect 2140 476 2148 484
rect 2156 476 2164 484
rect 2188 296 2196 304
rect 1708 196 1716 204
rect 1740 196 1748 204
rect 1628 176 1636 184
rect 1660 176 1668 184
rect 1628 156 1636 164
rect 1836 196 1844 204
rect 1820 156 1828 164
rect 1964 156 1972 164
rect 1932 136 1940 144
rect 2044 136 2052 144
rect 332 116 340 124
rect 604 116 612 124
rect 956 116 964 124
rect 1084 116 1092 124
rect 1356 116 1364 124
rect 1388 116 1396 124
rect 12 96 20 104
rect 590 6 598 14
rect 604 6 612 14
rect 618 6 626 14
rect 1404 16 1412 24
<< metal3 >>
rect 584 2014 632 2016
rect 584 2006 588 2014
rect 598 2006 604 2014
rect 612 2006 618 2014
rect 628 2006 632 2014
rect 584 2004 632 2006
rect 516 1937 540 1943
rect 356 1917 604 1923
rect 1204 1917 1500 1923
rect -19 1897 12 1903
rect 228 1897 268 1903
rect 388 1897 556 1903
rect 564 1897 684 1903
rect 980 1897 1100 1903
rect 1396 1897 1452 1903
rect 1460 1897 1676 1903
rect 1716 1897 1740 1903
rect 292 1877 380 1883
rect 468 1877 492 1883
rect 532 1877 572 1883
rect 596 1877 876 1883
rect 1572 1877 1644 1883
rect 52 1857 284 1863
rect 292 1857 444 1863
rect 468 1857 476 1863
rect 1204 1857 1228 1863
rect 116 1837 220 1843
rect 1940 1837 1980 1843
rect 180 1817 460 1823
rect 852 1817 908 1823
rect 916 1817 956 1823
rect 1780 1817 2028 1823
rect 1560 1814 1608 1816
rect 1560 1806 1564 1814
rect 1574 1806 1580 1814
rect 1588 1806 1594 1814
rect 1604 1806 1608 1814
rect 1560 1804 1608 1806
rect 1732 1797 1788 1803
rect 2221 1797 2227 1803
rect 1620 1777 1708 1783
rect 404 1757 492 1763
rect 532 1757 684 1763
rect 692 1757 876 1763
rect 884 1757 1020 1763
rect 1028 1757 1084 1763
rect 1364 1757 1596 1763
rect 1604 1757 1628 1763
rect 1636 1757 1660 1763
rect 1684 1757 1900 1763
rect 1908 1757 2076 1763
rect 708 1737 780 1743
rect 1444 1737 1628 1743
rect 1876 1737 1916 1743
rect 2132 1737 2227 1743
rect 452 1717 476 1723
rect 1780 1717 1852 1723
rect 2020 1717 2060 1723
rect 2068 1717 2140 1723
rect 500 1697 540 1703
rect 548 1697 684 1703
rect 692 1697 716 1703
rect 1172 1697 1468 1703
rect 1636 1697 1820 1703
rect 2196 1697 2227 1703
rect 292 1677 428 1683
rect 468 1677 492 1683
rect 1028 1637 1148 1643
rect 584 1614 632 1616
rect 584 1606 588 1614
rect 598 1606 604 1614
rect 612 1606 618 1614
rect 628 1606 632 1614
rect 584 1604 632 1606
rect 1732 1597 1804 1603
rect 1092 1577 1116 1583
rect 1620 1577 1676 1583
rect -19 1557 60 1563
rect 212 1537 668 1543
rect 2132 1537 2227 1543
rect -19 1517 12 1523
rect 356 1517 412 1523
rect 148 1497 188 1503
rect 388 1497 556 1503
rect 1540 1497 1772 1503
rect 2196 1497 2227 1503
rect -19 1477 -13 1483
rect 100 1477 140 1483
rect 148 1477 348 1483
rect 372 1477 524 1483
rect 836 1477 924 1483
rect 1108 1477 1132 1483
rect 1140 1477 1324 1483
rect 1428 1477 1708 1483
rect 1876 1477 1996 1483
rect 52 1457 108 1463
rect 116 1457 284 1463
rect 292 1457 380 1463
rect 564 1457 828 1463
rect 1204 1457 1276 1463
rect 1284 1457 1452 1463
rect 1460 1457 1900 1463
rect 1908 1457 1932 1463
rect 148 1437 204 1443
rect 228 1437 252 1443
rect -19 1417 -13 1423
rect 868 1417 924 1423
rect 1140 1417 1148 1423
rect 1560 1414 1608 1416
rect 1560 1406 1564 1414
rect 1574 1406 1580 1414
rect 1588 1406 1594 1414
rect 1604 1406 1608 1414
rect 1560 1404 1608 1406
rect 1460 1397 1500 1403
rect 196 1377 556 1383
rect 1892 1377 2076 1383
rect -19 1357 -13 1363
rect 372 1357 588 1363
rect 836 1357 956 1363
rect 1716 1357 1836 1363
rect 1940 1357 1964 1363
rect 420 1337 492 1343
rect 1108 1337 1180 1343
rect 1236 1337 1660 1343
rect 1668 1337 2140 1343
rect 324 1317 460 1323
rect 1284 1317 1468 1323
rect 1732 1317 1932 1323
rect 1188 1297 1324 1303
rect 1332 1297 1852 1303
rect 2196 1297 2227 1303
rect 548 1277 860 1283
rect 1172 1277 1292 1283
rect 1684 1277 1948 1283
rect 1956 1277 2108 1283
rect -19 1257 268 1263
rect -19 1217 348 1223
rect 584 1214 632 1216
rect 584 1206 588 1214
rect 598 1206 604 1214
rect 612 1206 618 1214
rect 628 1206 632 1214
rect 584 1204 632 1206
rect 1700 1197 1900 1203
rect 1908 1197 1916 1203
rect -19 1177 60 1183
rect 100 1177 460 1183
rect 468 1177 604 1183
rect 612 1177 1004 1183
rect 2221 1177 2227 1183
rect -19 1137 12 1143
rect 324 1137 444 1143
rect 244 1117 284 1123
rect -19 1097 -13 1103
rect 276 1097 300 1103
rect 468 1097 588 1103
rect 596 1097 684 1103
rect 804 1097 1036 1103
rect 1348 1097 1372 1103
rect 1380 1097 1388 1103
rect 1604 1097 1788 1103
rect 2196 1097 2227 1103
rect 52 1077 108 1083
rect 116 1077 220 1083
rect 276 1077 460 1083
rect 900 1077 1148 1083
rect 1252 1077 1340 1083
rect 1492 1077 1772 1083
rect 548 1057 764 1063
rect 164 1037 220 1043
rect 1652 1037 1836 1043
rect 1844 1037 1916 1043
rect 2036 1037 2076 1043
rect 148 1017 204 1023
rect 260 1017 380 1023
rect 1460 1017 1516 1023
rect 1892 1017 2076 1023
rect 1560 1014 1608 1016
rect 1560 1006 1564 1014
rect 1574 1006 1580 1014
rect 1588 1006 1594 1014
rect 1604 1006 1608 1014
rect 1560 1004 1608 1006
rect 404 957 940 963
rect 948 957 1004 963
rect 1124 957 1260 963
rect 1524 957 1644 963
rect 2221 957 2227 963
rect 308 937 572 943
rect 1012 937 1036 943
rect 1092 937 1292 943
rect 1620 937 1820 943
rect 1988 937 2028 943
rect 2036 937 2140 943
rect 836 917 956 923
rect 1396 917 1516 923
rect 1844 917 1996 923
rect 2004 917 2156 923
rect 324 897 668 903
rect 676 897 780 903
rect 1012 897 1100 903
rect 1108 897 1132 903
rect 1956 897 2044 903
rect 2196 897 2227 903
rect 1908 877 1916 883
rect 452 837 812 843
rect 820 837 1276 843
rect 1284 837 1292 843
rect 1124 817 1148 823
rect 1156 817 1404 823
rect 584 814 632 816
rect 584 806 588 814
rect 598 806 604 814
rect 612 806 618 814
rect 628 806 632 814
rect 584 804 632 806
rect -19 737 12 743
rect 932 737 1052 743
rect 1732 737 2227 743
rect 52 717 108 723
rect 116 717 284 723
rect 292 717 380 723
rect 1956 717 1996 723
rect -19 697 60 703
rect 148 697 156 703
rect 164 697 252 703
rect 1060 697 1100 703
rect 1588 697 1628 703
rect 1652 697 1692 703
rect 1844 697 1868 703
rect 1988 697 2012 703
rect 2196 697 2227 703
rect 36 677 156 683
rect 164 677 236 683
rect 516 677 716 683
rect 1028 677 1132 683
rect 1140 677 1260 683
rect 1268 677 1324 683
rect 1524 677 1676 683
rect 1684 677 1740 683
rect 1748 677 1852 683
rect 1908 677 1964 683
rect 1972 677 2092 683
rect 196 657 236 663
rect 244 657 540 663
rect 548 657 684 663
rect 692 657 892 663
rect 1108 657 1132 663
rect 1492 657 1516 663
rect 1620 657 1644 663
rect 1876 657 1980 663
rect 1988 657 2108 663
rect 2004 637 2044 643
rect 1560 614 1608 616
rect 1560 606 1564 614
rect 1574 606 1580 614
rect 1588 606 1594 614
rect 1604 606 1608 614
rect 1560 604 1608 606
rect 116 597 140 603
rect 100 557 412 563
rect 420 557 524 563
rect 532 557 556 563
rect 740 557 924 563
rect 932 557 1052 563
rect 1124 557 1196 563
rect 1812 557 1836 563
rect 2036 557 2124 563
rect 228 537 364 543
rect 516 537 652 543
rect 836 537 1036 543
rect 1380 537 1500 543
rect 1780 537 2012 543
rect -19 517 -13 523
rect 308 517 332 523
rect 404 517 540 523
rect 804 517 860 523
rect 884 517 924 523
rect 932 517 1020 523
rect 1028 517 1100 523
rect 1124 517 1148 523
rect 1204 517 1228 523
rect 1492 517 1676 523
rect 564 497 908 503
rect 1044 497 1068 503
rect 2196 497 2227 503
rect 324 477 364 483
rect 724 477 812 483
rect 1972 477 2044 483
rect 2052 477 2140 483
rect 2148 477 2156 483
rect 132 417 348 423
rect 356 417 396 423
rect 500 417 556 423
rect 1236 417 1260 423
rect 584 414 632 416
rect 584 406 588 414
rect 598 406 604 414
rect 612 406 618 414
rect 628 406 632 414
rect 584 404 632 406
rect 468 397 492 403
rect 1204 397 1468 403
rect 1316 377 1356 383
rect 1780 377 1788 383
rect 2020 357 2092 363
rect -19 337 12 343
rect 52 317 348 323
rect -19 297 -13 303
rect 84 297 124 303
rect 308 297 412 303
rect 724 297 860 303
rect 2196 297 2227 303
rect 84 277 188 283
rect 196 277 300 283
rect 308 277 380 283
rect 1044 277 1292 283
rect 900 257 1260 263
rect 1268 257 1404 263
rect 1428 257 1436 263
rect 1444 257 1516 263
rect 1572 257 1644 263
rect 1476 237 1580 243
rect 244 217 684 223
rect 1560 214 1608 216
rect 1560 206 1564 214
rect 1574 206 1580 214
rect 1588 206 1594 214
rect 1604 206 1608 214
rect 1560 204 1608 206
rect 740 197 892 203
rect 1716 197 1740 203
rect 1748 197 1836 203
rect 1012 177 1068 183
rect 1076 177 1116 183
rect 1636 177 1660 183
rect -19 157 -13 163
rect 1236 157 1260 163
rect 1636 157 1820 163
rect 1828 157 1964 163
rect 612 137 716 143
rect 916 137 1100 143
rect 1940 137 2044 143
rect 340 117 604 123
rect 964 117 1084 123
rect 1364 117 1388 123
rect 2221 117 2227 123
rect -19 97 12 103
rect 1396 17 1404 23
rect 584 14 632 16
rect 584 6 588 14
rect 598 6 604 14
rect 612 6 618 14
rect 628 6 632 14
rect 584 4 632 6
<< m4contact >>
rect 588 2006 590 2014
rect 590 2006 596 2014
rect 604 2006 612 2014
rect 620 2006 626 2014
rect 626 2006 628 2014
rect 460 1856 468 1864
rect 1932 1836 1940 1844
rect 460 1816 468 1824
rect 1564 1806 1566 1814
rect 1566 1806 1572 1814
rect 1580 1806 1588 1814
rect 1596 1806 1602 1814
rect 1602 1806 1604 1814
rect 1420 1716 1428 1724
rect 588 1606 590 1614
rect 590 1606 596 1614
rect 604 1606 612 1614
rect 620 1606 626 1614
rect 626 1606 628 1614
rect 1388 1596 1396 1604
rect 1932 1456 1940 1464
rect 140 1436 148 1444
rect 1132 1416 1140 1424
rect 1564 1406 1566 1414
rect 1566 1406 1572 1414
rect 1580 1406 1588 1414
rect 1596 1406 1602 1414
rect 1602 1406 1604 1414
rect 268 1256 276 1264
rect 588 1206 590 1214
rect 590 1206 596 1214
rect 604 1206 612 1214
rect 620 1206 626 1214
rect 626 1206 628 1214
rect 1900 1196 1908 1204
rect 460 1176 468 1184
rect 1292 1096 1300 1104
rect 268 1076 276 1084
rect 1836 1036 1844 1044
rect 140 1016 148 1024
rect 1564 1006 1566 1014
rect 1566 1006 1572 1014
rect 1580 1006 1588 1014
rect 1596 1006 1602 1014
rect 1602 1006 1604 1014
rect 1900 876 1908 884
rect 1292 836 1300 844
rect 588 806 590 814
rect 590 806 596 814
rect 604 806 612 814
rect 620 806 626 814
rect 626 806 628 814
rect 140 696 148 704
rect 1132 676 1140 684
rect 236 656 244 664
rect 1772 636 1780 644
rect 1564 606 1566 614
rect 1566 606 1572 614
rect 1580 606 1588 614
rect 1596 606 1602 614
rect 1602 606 1604 614
rect 108 596 116 604
rect 1836 556 1844 564
rect 1260 416 1268 424
rect 588 406 590 414
rect 590 406 596 414
rect 604 406 612 414
rect 620 406 626 414
rect 626 406 628 414
rect 1772 376 1780 384
rect 108 336 116 344
rect 1420 256 1428 264
rect 236 216 244 224
rect 1564 206 1566 214
rect 1566 206 1572 214
rect 1580 206 1588 214
rect 1596 206 1602 214
rect 1602 206 1604 214
rect 1260 136 1268 144
rect 1388 16 1396 24
rect 588 6 590 14
rect 590 6 596 14
rect 604 6 612 14
rect 620 6 626 14
rect 626 6 628 14
<< metal4 >>
rect 584 2014 632 2040
rect 584 2006 588 2014
rect 596 2006 604 2014
rect 612 2006 620 2014
rect 628 2006 632 2014
rect 458 1864 470 1866
rect 458 1856 460 1864
rect 468 1856 470 1864
rect 458 1824 470 1856
rect 458 1816 460 1824
rect 468 1816 470 1824
rect 138 1444 150 1446
rect 138 1436 140 1444
rect 148 1436 150 1444
rect 138 1024 150 1436
rect 266 1264 278 1266
rect 266 1256 268 1264
rect 276 1256 278 1264
rect 266 1084 278 1256
rect 458 1184 470 1816
rect 458 1176 460 1184
rect 468 1176 470 1184
rect 458 1174 470 1176
rect 584 1614 632 2006
rect 1560 1814 1608 2040
rect 1560 1806 1564 1814
rect 1572 1806 1580 1814
rect 1588 1806 1596 1814
rect 1604 1806 1608 1814
rect 584 1606 588 1614
rect 596 1606 604 1614
rect 612 1606 620 1614
rect 628 1606 632 1614
rect 1418 1724 1430 1726
rect 1418 1716 1420 1724
rect 1428 1716 1430 1724
rect 584 1214 632 1606
rect 1386 1604 1398 1606
rect 1386 1596 1388 1604
rect 1396 1596 1398 1604
rect 584 1206 588 1214
rect 596 1206 604 1214
rect 612 1206 620 1214
rect 628 1206 632 1214
rect 266 1076 268 1084
rect 276 1076 278 1084
rect 266 1074 278 1076
rect 138 1016 140 1024
rect 148 1016 150 1024
rect 138 704 150 1016
rect 138 696 140 704
rect 148 696 150 704
rect 138 694 150 696
rect 584 814 632 1206
rect 584 806 588 814
rect 596 806 604 814
rect 612 806 620 814
rect 628 806 632 814
rect 234 664 246 666
rect 234 656 236 664
rect 244 656 246 664
rect 106 604 118 606
rect 106 596 108 604
rect 116 596 118 604
rect 106 344 118 596
rect 106 336 108 344
rect 116 336 118 344
rect 106 334 118 336
rect 234 224 246 656
rect 234 216 236 224
rect 244 216 246 224
rect 234 214 246 216
rect 584 414 632 806
rect 1130 1424 1142 1426
rect 1130 1416 1132 1424
rect 1140 1416 1142 1424
rect 1130 684 1142 1416
rect 1290 1104 1302 1106
rect 1290 1096 1292 1104
rect 1300 1096 1302 1104
rect 1290 844 1302 1096
rect 1290 836 1292 844
rect 1300 836 1302 844
rect 1290 834 1302 836
rect 1130 676 1132 684
rect 1140 676 1142 684
rect 1130 674 1142 676
rect 584 406 588 414
rect 596 406 604 414
rect 612 406 620 414
rect 628 406 632 414
rect 584 14 632 406
rect 1258 424 1270 426
rect 1258 416 1260 424
rect 1268 416 1270 424
rect 1258 144 1270 416
rect 1258 136 1260 144
rect 1268 136 1270 144
rect 1258 134 1270 136
rect 1386 24 1398 1596
rect 1418 264 1430 1716
rect 1418 256 1420 264
rect 1428 256 1430 264
rect 1418 254 1430 256
rect 1560 1414 1608 1806
rect 1930 1844 1942 1846
rect 1930 1836 1932 1844
rect 1940 1836 1942 1844
rect 1930 1464 1942 1836
rect 1930 1456 1932 1464
rect 1940 1456 1942 1464
rect 1930 1454 1942 1456
rect 1560 1406 1564 1414
rect 1572 1406 1580 1414
rect 1588 1406 1596 1414
rect 1604 1406 1608 1414
rect 1560 1014 1608 1406
rect 1898 1204 1910 1206
rect 1898 1196 1900 1204
rect 1908 1196 1910 1204
rect 1560 1006 1564 1014
rect 1572 1006 1580 1014
rect 1588 1006 1596 1014
rect 1604 1006 1608 1014
rect 1560 614 1608 1006
rect 1834 1044 1846 1046
rect 1834 1036 1836 1044
rect 1844 1036 1846 1044
rect 1560 606 1564 614
rect 1572 606 1580 614
rect 1588 606 1596 614
rect 1604 606 1608 614
rect 1386 16 1388 24
rect 1396 16 1398 24
rect 1386 14 1398 16
rect 1560 214 1608 606
rect 1770 644 1782 646
rect 1770 636 1772 644
rect 1780 636 1782 644
rect 1770 384 1782 636
rect 1834 564 1846 1036
rect 1898 884 1910 1196
rect 1898 876 1900 884
rect 1908 876 1910 884
rect 1898 874 1910 876
rect 1834 556 1836 564
rect 1844 556 1846 564
rect 1834 554 1846 556
rect 1770 376 1772 384
rect 1780 376 1782 384
rect 1770 374 1782 376
rect 1560 206 1564 214
rect 1572 206 1580 214
rect 1588 206 1596 214
rect 1604 206 1608 214
rect 584 6 588 14
rect 596 6 604 14
rect 612 6 620 14
rect 628 6 632 14
rect 584 -40 632 6
rect 1560 -40 1608 206
use DFFSR  DFFSR_31
timestamp 1740382396
transform -1 0 408 0 -1 210
box -16 -6 368 210
use INVX1  INVX1_21
timestamp 1740382396
transform -1 0 184 0 1 210
box -18 -6 52 210
use INVX1  INVX1_20
timestamp 1740382396
transform 1 0 56 0 1 210
box -18 -6 52 210
use BUFX2  BUFX2_31
timestamp 1740382396
transform -1 0 56 0 1 210
box -10 -6 56 210
use BUFX2  BUFX2_30
timestamp 1740382396
transform -1 0 56 0 -1 210
box -10 -6 56 210
use XNOR2X1  XNOR2X1_13
timestamp 1740382396
transform -1 0 296 0 1 210
box -16 -6 128 210
use NAND3X1  NAND3X1_8
timestamp 1740382396
transform -1 0 152 0 1 210
box -16 -6 80 210
use OAI21X1  OAI21X1_7
timestamp 1740382396
transform 1 0 296 0 1 210
box -16 -6 68 210
use NOR3X1  NOR3X1_6
timestamp 1740382396
transform 1 0 360 0 1 210
box -14 -6 136 210
use FILL  FILL_72
timestamp 1740382396
transform 1 0 568 0 1 210
box -16 -6 32 210
use FILL  FILL_73
timestamp 1740382396
transform 1 0 584 0 1 210
box -16 -6 32 210
use FILL  FILL_74
timestamp 1740382396
transform -1 0 472 0 -1 210
box -16 -6 32 210
use FILL  FILL_75
timestamp 1740382396
transform -1 0 488 0 -1 210
box -16 -6 32 210
use FILL  FILL_76
timestamp 1740382396
transform -1 0 504 0 -1 210
box -16 -6 32 210
use INVX1  INVX1_19
timestamp 1740382396
transform -1 0 520 0 1 210
box -18 -6 52 210
use BUFX2  BUFX2_29
timestamp 1740382396
transform -1 0 456 0 -1 210
box -10 -6 56 210
use NAND2X1  NAND2X1_16
timestamp 1740382396
transform 1 0 520 0 1 210
box -16 -6 64 210
use FILL  FILL_71
timestamp 1740382396
transform 1 0 600 0 1 210
box -16 -6 32 210
use XNOR2X1  XNOR2X1_12
timestamp 1740382396
transform 1 0 616 0 1 210
box -16 -6 128 210
use DFFSR  DFFSR_29
timestamp 1740382396
transform -1 0 856 0 -1 210
box -16 -6 368 210
use DFFSR  DFFSR_30
timestamp 1740382396
transform 1 0 728 0 1 210
box -16 -6 368 210
use DFFSR  DFFSR_28
timestamp 1740382396
transform -1 0 1432 0 1 210
box -16 -6 368 210
use DFFSR  DFFSR_27
timestamp 1740382396
transform -1 0 1400 0 -1 210
box -16 -6 368 210
use BUFX2  BUFX2_28
timestamp 1740382396
transform 1 0 1000 0 -1 210
box -10 -6 56 210
use BUFX2  BUFX2_27
timestamp 1740382396
transform 1 0 952 0 -1 210
box -10 -6 56 210
use BUFX2  BUFX2_26
timestamp 1740382396
transform 1 0 904 0 -1 210
box -10 -6 56 210
use BUFX2  BUFX2_25
timestamp 1740382396
transform -1 0 904 0 -1 210
box -10 -6 56 210
use FILL  FILL_70
timestamp 1740382396
transform 1 0 1544 0 1 210
box -16 -6 32 210
use FILL  FILL_69
timestamp 1740382396
transform 1 0 1528 0 1 210
box -16 -6 32 210
use FILL  FILL_68
timestamp 1740382396
transform -1 0 1448 0 -1 210
box -16 -6 32 210
use FILL  FILL_67
timestamp 1740382396
transform -1 0 1432 0 -1 210
box -16 -6 32 210
use FILL  FILL_66
timestamp 1740382396
transform -1 0 1416 0 -1 210
box -16 -6 32 210
use DFFSR  DFFSR_26
timestamp 1740382396
transform -1 0 1800 0 -1 210
box -16 -6 368 210
use NOR2X1  NOR2X1_11
timestamp 1740382396
transform -1 0 1528 0 1 210
box -16 -6 64 210
use NAND2X1  NAND2X1_15
timestamp 1740382396
transform 1 0 1432 0 1 210
box -16 -6 64 210
use FILL  FILL_65
timestamp 1740382396
transform 1 0 1560 0 1 210
box -16 -6 32 210
use DFFSR  DFFSR_25
timestamp 1740382396
transform 1 0 1656 0 1 210
box -16 -6 368 210
use DFFSR  DFFSR_24
timestamp 1740382396
transform 1 0 1800 0 -1 210
box -16 -6 368 210
use NOR2X1  NOR2X1_10
timestamp 1740382396
transform -1 0 1656 0 1 210
box -16 -6 64 210
use INVX1  INVX1_18
timestamp 1740382396
transform 1 0 1576 0 1 210
box -18 -6 52 210
use FILL  FILL_64
timestamp 1740382396
transform 1 0 2184 0 1 210
box -16 -6 32 210
use FILL  FILL_63
timestamp 1740382396
transform -1 0 2200 0 -1 210
box -16 -6 32 210
use FILL  FILL_62
timestamp 1740382396
transform 1 0 2168 0 1 210
box -16 -6 32 210
use FILL  FILL_61
timestamp 1740382396
transform -1 0 2184 0 -1 210
box -16 -6 32 210
use FILL  FILL_60
timestamp 1740382396
transform -1 0 2168 0 -1 210
box -16 -6 32 210
use BUFX2  BUFX2_24
timestamp 1740382396
transform 1 0 2120 0 1 210
box -10 -6 56 210
use XOR2X1  XOR2X1_5
timestamp 1740382396
transform 1 0 2008 0 1 210
box -16 -6 128 210
use DFFSR  DFFSR_23
timestamp 1740382396
transform -1 0 360 0 -1 610
box -16 -6 368 210
use NAND2X1  NAND2X1_14
timestamp 1740382396
transform -1 0 408 0 -1 610
box -16 -6 64 210
use FILL  FILL_59
timestamp 1740382396
transform 1 0 600 0 -1 610
box -16 -6 32 210
use FILL  FILL_58
timestamp 1740382396
transform 1 0 584 0 -1 610
box -16 -6 32 210
use FILL  FILL_57
timestamp 1740382396
transform 1 0 568 0 -1 610
box -16 -6 32 210
use INVX1  INVX1_17
timestamp 1740382396
transform 1 0 744 0 -1 610
box -18 -6 52 210
use INVX1  INVX1_16
timestamp 1740382396
transform 1 0 408 0 -1 610
box -18 -6 52 210
use NAND3X1  NAND3X1_7
timestamp 1740382396
transform 1 0 776 0 -1 610
box -16 -6 80 210
use NAND3X1  NAND3X1_6
timestamp 1740382396
transform 1 0 440 0 -1 610
box -16 -6 80 210
use OAI21X1  OAI21X1_6
timestamp 1740382396
transform -1 0 568 0 -1 610
box -16 -6 68 210
use NOR3X1  NOR3X1_5
timestamp 1740382396
transform 1 0 616 0 -1 610
box -14 -6 136 210
use AND2X2  AND2X2_5
timestamp 1740382396
transform 1 0 1128 0 -1 610
box -16 -6 80 210
use NOR2X1  NOR2X1_9
timestamp 1740382396
transform 1 0 1080 0 -1 610
box -16 -6 64 210
use NAND2X1  NAND2X1_13
timestamp 1740382396
transform 1 0 1032 0 -1 610
box -16 -6 64 210
use OAI21X1  OAI21X1_5
timestamp 1740382396
transform 1 0 968 0 -1 610
box -16 -6 68 210
use NOR3X1  NOR3X1_4
timestamp 1740382396
transform -1 0 968 0 -1 610
box -14 -6 136 210
use DFFSR  DFFSR_22
timestamp 1740382396
transform 1 0 1240 0 -1 610
box -16 -6 368 210
use NOR2X1  NOR2X1_8
timestamp 1740382396
transform 1 0 1192 0 -1 610
box -16 -6 64 210
use FILL  FILL_56
timestamp 1740382396
transform 1 0 1624 0 -1 610
box -16 -6 32 210
use FILL  FILL_55
timestamp 1740382396
transform 1 0 1608 0 -1 610
box -16 -6 32 210
use FILL  FILL_54
timestamp 1740382396
transform 1 0 1592 0 -1 610
box -16 -6 32 210
use DFFSR  DFFSR_21
timestamp 1740382396
transform 1 0 1640 0 -1 610
box -16 -6 368 210
use NOR2X1  NOR2X1_7
timestamp 1740382396
transform -1 0 2040 0 -1 610
box -16 -6 64 210
use BUFX2  BUFX2_23
timestamp 1740382396
transform 1 0 2152 0 -1 610
box -10 -6 56 210
use NAND2X1  NAND2X1_12
timestamp 1740382396
transform -1 0 2088 0 -1 610
box -16 -6 64 210
use AOI21X1  AOI21X1_0
timestamp 1740382396
transform 1 0 2088 0 -1 610
box -14 -6 78 210
use BUFX2  BUFX2_22
timestamp 1740382396
transform -1 0 104 0 1 610
box -10 -6 56 210
use BUFX2  BUFX2_21
timestamp 1740382396
transform -1 0 56 0 1 610
box -10 -6 56 210
use XNOR2X1  XNOR2X1_11
timestamp 1740382396
transform 1 0 344 0 1 610
box -16 -6 128 210
use NAND2X1  NAND2X1_11
timestamp 1740382396
transform 1 0 296 0 1 610
box -16 -6 64 210
use OAI21X1  OAI21X1_4
timestamp 1740382396
transform 1 0 232 0 1 610
box -16 -6 68 210
use NOR3X1  NOR3X1_3
timestamp 1740382396
transform 1 0 104 0 1 610
box -14 -6 136 210
use FILL  FILL_53
timestamp 1740382396
transform -1 0 504 0 1 610
box -16 -6 32 210
use FILL  FILL_52
timestamp 1740382396
transform -1 0 488 0 1 610
box -16 -6 32 210
use FILL  FILL_51
timestamp 1740382396
transform -1 0 472 0 1 610
box -16 -6 32 210
use DFFSR  DFFSR_20
timestamp 1740382396
transform -1 0 856 0 1 610
box -16 -6 368 210
use INVX1  INVX1_15
timestamp 1740382396
transform 1 0 1096 0 1 610
box -18 -6 52 210
use INVX1  INVX1_14
timestamp 1740382396
transform -1 0 888 0 1 610
box -18 -6 52 210
use NAND3X1  NAND3X1_5
timestamp 1740382396
transform 1 0 1032 0 1 610
box -16 -6 80 210
use CLKBUF1  CLKBUF1_4
timestamp 1740382396
transform -1 0 1272 0 1 610
box -16 -6 160 210
use CLKBUF1  CLKBUF1_3
timestamp 1740382396
transform -1 0 1032 0 1 610
box -16 -6 160 210
use FILL  FILL_50
timestamp 1740382396
transform -1 0 1560 0 1 610
box -16 -6 32 210
use FILL  FILL_49
timestamp 1740382396
transform -1 0 1544 0 1 610
box -16 -6 32 210
use NOR2X1  NOR2X1_6
timestamp 1740382396
transform 1 0 1480 0 1 610
box -16 -6 64 210
use CLKBUF1  CLKBUF1_2
timestamp 1740382396
transform 1 0 1336 0 1 610
box -16 -6 160 210
use BUFX4  BUFX4_4
timestamp 1740382396
transform 1 0 1272 0 1 610
box -18 -6 74 210
use FILL  FILL_48
timestamp 1740382396
transform -1 0 1576 0 1 610
box -16 -6 32 210
use AND2X2  AND2X2_4
timestamp 1740382396
transform -1 0 1976 0 1 610
box -16 -6 80 210
use AND2X2  AND2X2_3
timestamp 1740382396
transform 1 0 1848 0 1 610
box -16 -6 80 210
use AND2X2  AND2X2_2
timestamp 1740382396
transform 1 0 1624 0 1 610
box -16 -6 80 210
use NOR2X1  NOR2X1_5
timestamp 1740382396
transform -1 0 1624 0 1 610
box -16 -6 64 210
use BUFX2  BUFX2_20
timestamp 1740382396
transform 1 0 1688 0 1 610
box -10 -6 56 210
use XOR2X1  XOR2X1_4
timestamp 1740382396
transform 1 0 1736 0 1 610
box -16 -6 128 210
use FILL  FILL_47
timestamp 1740382396
transform 1 0 2184 0 1 610
box -16 -6 32 210
use FILL  FILL_46
timestamp 1740382396
transform 1 0 2168 0 1 610
box -16 -6 32 210
use FILL  FILL_45
timestamp 1740382396
transform 1 0 2152 0 1 610
box -16 -6 32 210
use NOR2X1  NOR2X1_4
timestamp 1740382396
transform 1 0 2024 0 1 610
box -16 -6 64 210
use NOR2X1  NOR2X1_3
timestamp 1740382396
transform -1 0 2024 0 1 610
box -16 -6 64 210
use INVX1  INVX1_13
timestamp 1740382396
transform -1 0 2104 0 1 610
box -18 -6 52 210
use BUFX2  BUFX2_19
timestamp 1740382396
transform 1 0 2104 0 1 610
box -10 -6 56 210
use DFFSR  DFFSR_19
timestamp 1740382396
transform -1 0 712 0 -1 1010
box -16 -6 368 210
use DFFSR  DFFSR_18
timestamp 1740382396
transform -1 0 360 0 -1 1010
box -16 -6 368 210
use FILL  FILL_44
timestamp 1740382396
transform -1 0 760 0 -1 1010
box -16 -6 32 210
use FILL  FILL_43
timestamp 1740382396
transform -1 0 744 0 -1 1010
box -16 -6 32 210
use FILL  FILL_42
timestamp 1740382396
transform -1 0 728 0 -1 1010
box -16 -6 32 210
use BUFX4  BUFX4_3
timestamp 1740382396
transform -1 0 824 0 -1 1010
box -18 -6 74 210
use DFFSR  DFFSR_17
timestamp 1740382396
transform -1 0 1432 0 -1 1010
box -16 -6 368 210
use INVX1  INVX1_12
timestamp 1740382396
transform 1 0 1000 0 -1 1010
box -18 -6 52 210
use XNOR2X1  XNOR2X1_10
timestamp 1740382396
transform 1 0 824 0 -1 1010
box -16 -6 128 210
use NAND2X1  NAND2X1_10
timestamp 1740382396
transform 1 0 1032 0 -1 1010
box -16 -6 64 210
use OAI21X1  OAI21X1_3
timestamp 1740382396
transform 1 0 936 0 -1 1010
box -16 -6 68 210
use FILL  FILL_41
timestamp 1740382396
transform 1 0 1464 0 -1 1010
box -16 -6 32 210
use FILL  FILL_40
timestamp 1740382396
transform 1 0 1448 0 -1 1010
box -16 -6 32 210
use FILL  FILL_39
timestamp 1740382396
transform 1 0 1432 0 -1 1010
box -16 -6 32 210
use DFFSR  DFFSR_16
timestamp 1740382396
transform 1 0 1480 0 -1 1010
box -16 -6 368 210
use XNOR2X1  XNOR2X1_9
timestamp 1740382396
transform -1 0 1944 0 -1 1010
box -16 -6 128 210
use BUFX2  BUFX2_18
timestamp 1740382396
transform 1 0 2152 0 -1 1010
box -10 -6 56 210
use NAND2X1  NAND2X1_9
timestamp 1740382396
transform -1 0 2040 0 -1 1010
box -16 -6 64 210
use NAND2X1  NAND2X1_8
timestamp 1740382396
transform -1 0 1992 0 -1 1010
box -16 -6 64 210
use XOR2X1  XOR2X1_3
timestamp 1740382396
transform 1 0 2040 0 -1 1010
box -16 -6 128 210
use INVX1  INVX1_11
timestamp 1740382396
transform 1 0 248 0 1 1010
box -18 -6 52 210
use INVX1  INVX1_10
timestamp 1740382396
transform 1 0 216 0 1 1010
box -18 -6 52 210
use BUFX2  BUFX2_17
timestamp 1740382396
transform -1 0 392 0 1 1010
box -10 -6 56 210
use BUFX2  BUFX2_16
timestamp 1740382396
transform -1 0 104 0 1 1010
box -10 -6 56 210
use BUFX2  BUFX2_15
timestamp 1740382396
transform -1 0 56 0 1 1010
box -10 -6 56 210
use XNOR2X1  XNOR2X1_8
timestamp 1740382396
transform -1 0 216 0 1 1010
box -16 -6 128 210
use NAND3X1  NAND3X1_4
timestamp 1740382396
transform 1 0 280 0 1 1010
box -16 -6 80 210
use FILL  FILL_38
timestamp 1740382396
transform -1 0 584 0 1 1010
box -16 -6 32 210
use FILL  FILL_37
timestamp 1740382396
transform -1 0 568 0 1 1010
box -16 -6 32 210
use FILL  FILL_36
timestamp 1740382396
transform -1 0 552 0 1 1010
box -16 -6 32 210
use DFFSR  DFFSR_15
timestamp 1740382396
transform -1 0 936 0 1 1010
box -16 -6 368 210
use BUFX4  BUFX4_2
timestamp 1740382396
transform 1 0 472 0 1 1010
box -18 -6 74 210
use INVX8  INVX8_0
timestamp 1740382396
transform -1 0 472 0 1 1010
box -18 -6 90 210
use DFFSR  DFFSR_14
timestamp 1740382396
transform -1 0 1288 0 1 1010
box -16 -6 368 210
use DFFSR  DFFSR_13
timestamp 1740382396
transform 1 0 1352 0 1 1010
box -16 -6 368 210
use BUFX4  BUFX4_1
timestamp 1740382396
transform 1 0 1288 0 1 1010
box -18 -6 74 210
use FILL  FILL_35
timestamp 1740382396
transform 1 0 1736 0 1 1010
box -16 -6 32 210
use FILL  FILL_34
timestamp 1740382396
transform 1 0 1720 0 1 1010
box -16 -6 32 210
use FILL  FILL_33
timestamp 1740382396
transform 1 0 1704 0 1 1010
box -16 -6 32 210
use DFFSR  DFFSR_12
timestamp 1740382396
transform 1 0 1752 0 1 1010
box -16 -6 368 210
use FILL  FILL_32
timestamp 1740382396
transform 1 0 2184 0 1 1010
box -16 -6 32 210
use FILL  FILL_31
timestamp 1740382396
transform 1 0 2168 0 1 1010
box -16 -6 32 210
use FILL  FILL_30
timestamp 1740382396
transform 1 0 2152 0 1 1010
box -16 -6 32 210
use BUFX2  BUFX2_14
timestamp 1740382396
transform 1 0 2104 0 1 1010
box -10 -6 56 210
use DFFSR  DFFSR_11
timestamp 1740382396
transform -1 0 360 0 -1 1410
box -16 -6 368 210
use NOR3X1  NOR3X1_2
timestamp 1740382396
transform 1 0 360 0 -1 1410
box -14 -6 136 210
use FILL  FILL_29
timestamp 1740382396
transform -1 0 648 0 -1 1410
box -16 -6 32 210
use FILL  FILL_28
timestamp 1740382396
transform -1 0 632 0 -1 1410
box -16 -6 32 210
use FILL  FILL_27
timestamp 1740382396
transform -1 0 616 0 -1 1410
box -16 -6 32 210
use DFFSR  DFFSR_10
timestamp 1740382396
transform -1 0 1000 0 -1 1410
box -16 -6 368 210
use XNOR2X1  XNOR2X1_7
timestamp 1740382396
transform 1 0 488 0 -1 1410
box -16 -6 128 210
use XNOR2X1  XNOR2X1_6
timestamp 1740382396
transform -1 0 1112 0 -1 1410
box -16 -6 128 210
use BUFX4  BUFX4_0
timestamp 1740382396
transform -1 0 1176 0 -1 1410
box -18 -6 74 210
use DFFSR  DFFSR_9
timestamp 1740382396
transform 1 0 1336 0 -1 1410
box -16 -6 368 210
use NAND2X1  NAND2X1_7
timestamp 1740382396
transform -1 0 1224 0 -1 1410
box -16 -6 64 210
use XOR2X1  XOR2X1_2
timestamp 1740382396
transform -1 0 1336 0 -1 1410
box -16 -6 128 210
use FILL  FILL_26
timestamp 1740382396
transform -1 0 1736 0 -1 1410
box -16 -6 32 210
use FILL  FILL_25
timestamp 1740382396
transform -1 0 1720 0 -1 1410
box -16 -6 32 210
use FILL  FILL_24
timestamp 1740382396
transform -1 0 1704 0 -1 1410
box -16 -6 32 210
use NOR2X1  NOR2X1_2
timestamp 1740382396
transform -1 0 1896 0 -1 1410
box -16 -6 64 210
use XNOR2X1  XNOR2X1_5
timestamp 1740382396
transform -1 0 1848 0 -1 1410
box -16 -6 128 210
use NAND3X1  NAND3X1_3
timestamp 1740382396
transform -1 0 1960 0 -1 1410
box -16 -6 80 210
use FILL  FILL_23
timestamp 1740382396
transform -1 0 2200 0 -1 1410
box -16 -6 32 210
use FILL  FILL_22
timestamp 1740382396
transform -1 0 2184 0 -1 1410
box -16 -6 32 210
use BUFX2  BUFX2_13
timestamp 1740382396
transform 1 0 2120 0 -1 1410
box -10 -6 56 210
use XNOR2X1  XNOR2X1_4
timestamp 1740382396
transform 1 0 1960 0 -1 1410
box -16 -6 128 210
use NAND2X1  NAND2X1_6
timestamp 1740382396
transform -1 0 2120 0 -1 1410
box -16 -6 64 210
use DFFSR  DFFSR_8
timestamp 1740382396
transform 1 0 392 0 1 1410
box -16 -6 368 210
use INVX1  INVX1_9
timestamp 1740382396
transform 1 0 136 0 1 1410
box -18 -6 52 210
use INVX1  INVX1_8
timestamp 1740382396
transform 1 0 104 0 1 1410
box -18 -6 52 210
use BUFX2  BUFX2_12
timestamp 1740382396
transform -1 0 104 0 1 1410
box -10 -6 56 210
use BUFX2  BUFX2_11
timestamp 1740382396
transform -1 0 56 0 1 1410
box -10 -6 56 210
use NAND2X1  NAND2X1_5
timestamp 1740382396
transform -1 0 392 0 1 1410
box -16 -6 64 210
use NAND2X1  NAND2X1_4
timestamp 1740382396
transform 1 0 232 0 1 1410
box -16 -6 64 210
use NAND3X1  NAND3X1_2
timestamp 1740382396
transform 1 0 168 0 1 1410
box -16 -6 80 210
use OAI21X1  OAI21X1_2
timestamp 1740382396
transform -1 0 344 0 1 1410
box -16 -6 68 210
use FILL  FILL_21
timestamp 1740382396
transform 1 0 776 0 1 1410
box -16 -6 32 210
use FILL  FILL_20
timestamp 1740382396
transform 1 0 760 0 1 1410
box -16 -6 32 210
use FILL  FILL_19
timestamp 1740382396
transform 1 0 744 0 1 1410
box -16 -6 32 210
use DFFSR  DFFSR_7
timestamp 1740382396
transform 1 0 792 0 1 1410
box -16 -6 368 210
use CLKBUF1  CLKBUF1_1
timestamp 1740382396
transform 1 0 1144 0 1 1410
box -16 -6 160 210
use DFFSR  DFFSR_6
timestamp 1740382396
transform 1 0 1288 0 1 1410
box -16 -6 368 210
use FILL  FILL_18
timestamp 1740382396
transform -1 0 1688 0 1 1410
box -16 -6 32 210
use FILL  FILL_17
timestamp 1740382396
transform -1 0 1672 0 1 1410
box -16 -6 32 210
use FILL  FILL_16
timestamp 1740382396
transform -1 0 1656 0 1 1410
box -16 -6 32 210
use DFFSR  DFFSR_5
timestamp 1740382396
transform 1 0 1736 0 1 1410
box -16 -6 368 210
use NAND2X1  NAND2X1_3
timestamp 1740382396
transform -1 0 1736 0 1 1410
box -16 -6 64 210
use FILL  FILL_15
timestamp 1740382396
transform 1 0 2184 0 1 1410
box -16 -6 32 210
use BUFX2  BUFX2_10
timestamp 1740382396
transform 1 0 2136 0 1 1410
box -10 -6 56 210
use BUFX2  BUFX2_9
timestamp 1740382396
transform 1 0 2088 0 1 1410
box -10 -6 56 210
use DFFSR  DFFSR_4
timestamp 1740382396
transform -1 0 360 0 -1 1810
box -16 -6 368 210
use BUFX2  BUFX2_8
timestamp 1740382396
transform -1 0 408 0 -1 1810
box -10 -6 56 210
use FILL  FILL_14
timestamp 1740382396
transform 1 0 632 0 -1 1810
box -16 -6 32 210
use FILL  FILL_13
timestamp 1740382396
transform 1 0 616 0 -1 1810
box -16 -6 32 210
use FILL  FILL_12
timestamp 1740382396
transform 1 0 600 0 -1 1810
box -16 -6 32 210
use INVX1  INVX1_7
timestamp 1740382396
transform -1 0 536 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_6
timestamp 1740382396
transform -1 0 504 0 -1 1810
box -18 -6 52 210
use XNOR2X1  XNOR2X1_3
timestamp 1740382396
transform 1 0 776 0 -1 1810
box -16 -6 128 210
use NAND3X1  NAND3X1_1
timestamp 1740382396
transform -1 0 472 0 -1 1810
box -16 -6 80 210
use OAI21X1  OAI21X1_1
timestamp 1740382396
transform -1 0 600 0 -1 1810
box -16 -6 68 210
use NOR3X1  NOR3X1_1
timestamp 1740382396
transform 1 0 648 0 -1 1810
box -14 -6 136 210
use DFFSR  DFFSR_3
timestamp 1740382396
transform 1 0 1032 0 -1 1810
box -16 -6 368 210
use CLKBUF1  CLKBUF1_0
timestamp 1740382396
transform -1 0 1032 0 -1 1810
box -16 -6 160 210
use FILL  FILL_11
timestamp 1740382396
transform 1 0 1544 0 -1 1810
box -16 -6 32 210
use BUFX2  BUFX2_7
timestamp 1740382396
transform -1 0 1432 0 -1 1810
box -10 -6 56 210
use XNOR2X1  XNOR2X1_2
timestamp 1740382396
transform 1 0 1432 0 -1 1810
box -16 -6 128 210
use FILL  FILL_10
timestamp 1740382396
transform 1 0 1576 0 -1 1810
box -16 -6 32 210
use FILL  FILL_9
timestamp 1740382396
transform 1 0 1560 0 -1 1810
box -16 -6 32 210
use NOR2X1  NOR2X1_1
timestamp 1740382396
transform -1 0 1880 0 -1 1810
box -16 -6 64 210
use INVX1  INVX1_5
timestamp 1740382396
transform -1 0 1912 0 -1 1810
box -18 -6 52 210
use INVX1  INVX1_4
timestamp 1740382396
transform 1 0 1592 0 -1 1810
box -18 -6 52 210
use XNOR2X1  XNOR2X1_1
timestamp 1740382396
transform -1 0 1784 0 -1 1810
box -16 -6 128 210
use NAND2X1  NAND2X1_2
timestamp 1740382396
transform 1 0 1784 0 -1 1810
box -16 -6 64 210
use NAND2X1  NAND2X1_1
timestamp 1740382396
transform -1 0 1672 0 -1 1810
box -16 -6 64 210
use XOR2X1  XOR2X1_1
timestamp 1740382396
transform 1 0 1912 0 -1 1810
box -16 -6 128 210
use FILL  FILL_8
timestamp 1740382396
transform -1 0 2200 0 -1 1810
box -16 -6 32 210
use AND2X2  AND2X2_1
timestamp 1740382396
transform -1 0 2088 0 -1 1810
box -16 -6 80 210
use BUFX2  BUFX2_6
timestamp 1740382396
transform 1 0 2136 0 -1 1810
box -10 -6 56 210
use BUFX2  BUFX2_5
timestamp 1740382396
transform 1 0 2088 0 -1 1810
box -10 -6 56 210
use INVX1  INVX1_3
timestamp 1740382396
transform 1 0 168 0 1 1810
box -18 -6 52 210
use BUFX2  BUFX2_4
timestamp 1740382396
transform -1 0 56 0 1 1810
box -10 -6 56 210
use OAI21X1  OAI21X1_0
timestamp 1740382396
transform 1 0 328 0 1 1810
box -16 -6 68 210
use NOR3X1  NOR3X1_0
timestamp 1740382396
transform -1 0 328 0 1 1810
box -14 -6 136 210
use XOR2X1  XOR2X1_0
timestamp 1740382396
transform 1 0 56 0 1 1810
box -16 -6 128 210
use FILL  FILL_7
timestamp 1740382396
transform -1 0 664 0 1 1810
box -16 -6 32 210
use FILL  FILL_6
timestamp 1740382396
transform -1 0 648 0 1 1810
box -16 -6 32 210
use FILL  FILL_5
timestamp 1740382396
transform -1 0 632 0 1 1810
box -16 -6 32 210
use DFFSR  DFFSR_2
timestamp 1740382396
transform -1 0 1016 0 1 1810
box -16 -6 368 210
use INVX1  INVX1_2
timestamp 1740382396
transform -1 0 568 0 1 1810
box -18 -6 52 210
use INVX1  INVX1_1
timestamp 1740382396
transform 1 0 440 0 1 1810
box -18 -6 52 210
use BUFX2  BUFX2_3
timestamp 1740382396
transform 1 0 392 0 1 1810
box -10 -6 56 210
use NAND2X1  NAND2X1_0
timestamp 1740382396
transform 1 0 568 0 1 1810
box -16 -6 64 210
use NAND3X1  NAND3X1_0
timestamp 1740382396
transform 1 0 472 0 1 1810
box -16 -6 80 210
use DFFSR  DFFSR_1
timestamp 1740382396
transform 1 0 1064 0 1 1810
box -16 -6 368 210
use BUFX2  BUFX2_2
timestamp 1740382396
transform 1 0 1016 0 1 1810
box -10 -6 56 210
use BUFX2  BUFX2_1
timestamp 1740382396
transform -1 0 1464 0 1 1810
box -10 -6 56 210
use XNOR2X1  XNOR2X1_0
timestamp 1740382396
transform -1 0 1576 0 1 1810
box -16 -6 128 210
use FILL  FILL_4
timestamp 1740382396
transform 1 0 1608 0 1 1810
box -16 -6 32 210
use FILL  FILL_3
timestamp 1740382396
transform 1 0 1592 0 1 1810
box -16 -6 32 210
use FILL  FILL_2
timestamp 1740382396
transform 1 0 1576 0 1 1810
box -16 -6 32 210
use DFFSR  DFFSR_0
timestamp 1740382396
transform 1 0 1816 0 1 1810
box -16 -6 368 210
use AND2X2  AND2X2_0
timestamp 1740382396
transform 1 0 1752 0 1 1810
box -16 -6 80 210
use NOR2X1  NOR2X1_0
timestamp 1740382396
transform 1 0 1704 0 1 1810
box -16 -6 64 210
use INVX1  INVX1_0
timestamp 1740382396
transform 1 0 1672 0 1 1810
box -18 -6 52 210
use BUFX2  BUFX2_0
timestamp 1740382396
transform 1 0 1624 0 1 1810
box -10 -6 56 210
use FILL  FILL_1
timestamp 1740382396
transform 1 0 2184 0 1 1810
box -16 -6 32 210
use FILL  FILL_0
timestamp 1740382396
transform 1 0 2168 0 1 1810
box -16 -6 32 210
<< labels >>
flabel metal4 608 -28 608 -28 7 FreeSans 30 270 0 0 vdd
flabel metal4 1584 -28 1584 -28 7 FreeSans 30 270 0 0 gnd
flabel metal2 1024 2040 1024 2040 3 FreeSans 30 90 0 0 clk
flabel metal3 -16 1260 -16 1260 7 FreeSans 30 0 0 0 rst
flabel metal3 -16 520 -16 520 7 FreeSans 30 0 0 0 theta[0]
flabel metal3 -16 300 -16 300 7 FreeSans 30 0 0 0 theta[1]
flabel metal3 2224 120 2224 120 3 FreeSans 30 0 0 0 theta[2]
flabel metal3 -16 1420 -16 1420 7 FreeSans 30 0 0 0 theta[3]
flabel metal3 -16 1360 -16 1360 7 FreeSans 30 0 0 0 theta[4]
flabel metal3 2224 1180 2224 1180 3 FreeSans 30 0 0 0 theta[5]
flabel metal2 1728 2040 1728 2040 3 FreeSans 30 90 0 0 theta[6]
flabel metal2 2016 2040 2016 2040 3 FreeSans 30 90 0 0 theta[7]
flabel metal2 480 -20 480 -20 7 FreeSans 30 270 0 0 theta[8]
flabel metal3 -16 160 -16 160 7 FreeSans 30 0 0 0 theta[9]
flabel metal3 -16 1100 -16 1100 7 FreeSans 30 0 0 0 theta[10]
flabel metal2 1456 -20 1456 -20 7 FreeSans 30 270 0 0 theta[11]
flabel metal3 -16 1480 -16 1480 7 FreeSans 30 0 0 0 theta[12]
flabel metal2 1680 2040 1680 2040 3 FreeSans 30 90 0 0 theta[13]
flabel metal3 2224 1800 2224 1800 3 FreeSans 30 0 0 0 theta[14]
flabel metal3 2224 960 2224 960 3 FreeSans 30 0 0 0 theta[15]
flabel metal2 1024 -20 1024 -20 7 FreeSans 30 270 0 0 sine[0]
flabel metal2 1408 -20 1408 -20 7 FreeSans 30 270 0 0 sine[1]
flabel metal3 2224 740 2224 740 3 FreeSans 30 0 0 0 sine[2]
flabel metal3 2224 700 2224 700 3 FreeSans 30 0 0 0 sine[3]
flabel metal3 2224 300 2224 300 3 FreeSans 30 0 0 0 sine[4]
flabel metal3 2224 500 2224 500 3 FreeSans 30 0 0 0 sine[5]
flabel metal3 2224 1100 2224 1100 3 FreeSans 30 0 0 0 sine[6]
flabel metal3 2224 900 2224 900 3 FreeSans 30 0 0 0 sine[7]
flabel metal2 1648 2040 1648 2040 3 FreeSans 30 90 0 0 sine[8]
flabel metal2 1440 2040 1440 2040 3 FreeSans 30 90 0 0 sine[9]
flabel metal3 2224 1740 2224 1740 3 FreeSans 30 0 0 0 sine[10]
flabel metal3 2224 1700 2224 1700 3 FreeSans 30 0 0 0 sine[11]
flabel metal3 2224 1300 2224 1300 3 FreeSans 30 0 0 0 sine[12]
flabel metal3 2224 1540 2224 1540 3 FreeSans 30 0 0 0 sine[13]
flabel metal3 2224 1500 2224 1500 3 FreeSans 30 0 0 0 sine[14]
flabel metal3 -16 1180 -16 1180 7 FreeSans 30 0 0 0 sine[15]
flabel metal3 -16 1900 -16 1900 7 FreeSans 30 0 0 0 cosine[0]
flabel metal2 416 2040 416 2040 3 FreeSans 30 90 0 0 cosine[1]
flabel metal2 1056 2040 1056 2040 3 FreeSans 30 90 0 0 cosine[2]
flabel metal2 384 2040 384 2040 3 FreeSans 30 90 0 0 cosine[3]
flabel metal3 -16 1560 -16 1560 7 FreeSans 30 0 0 0 cosine[4]
flabel metal3 -16 1520 -16 1520 7 FreeSans 30 0 0 0 cosine[5]
flabel metal3 -16 1140 -16 1140 7 FreeSans 30 0 0 0 cosine[6]
flabel metal3 -16 740 -16 740 7 FreeSans 30 0 0 0 cosine[7]
flabel metal3 -16 100 -16 100 7 FreeSans 30 0 0 0 cosine[8]
flabel metal3 -16 340 -16 340 7 FreeSans 30 0 0 0 cosine[9]
flabel metal3 -16 700 -16 700 7 FreeSans 30 0 0 0 cosine[10]
flabel metal2 432 -20 432 -20 7 FreeSans 30 270 0 0 cosine[11]
flabel metal2 880 -20 880 -20 7 FreeSans 30 270 0 0 cosine[12]
flabel metal2 928 -20 928 -20 7 FreeSans 30 270 0 0 cosine[13]
flabel metal3 -16 1220 -16 1220 7 FreeSans 30 0 0 0 cosine[14]
flabel metal2 976 -20 976 -20 7 FreeSans 30 270 0 0 cosine[15]
<< end >>

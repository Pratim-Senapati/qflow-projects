* NGSPICE file created from fft_top.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

.subckt fft_top vdd gnd clk reset start x0[0] x0[1] x0[2] x0[3] x0[4] x0[5] x0[6]
+ x0[7] x1[0] x1[1] x1[2] x1[3] x1[4] x1[5] x1[6] x1[7] x2[0] x2[1] x2[2] x2[3] x2[4]
+ x2[5] x2[6] x2[7] x3[0] x3[1] x3[2] x3[3] x3[4] x3[5] x3[6] x3[7] X0_mag[0] X0_mag[1]
+ X0_mag[2] X0_mag[3] X0_mag[4] X0_mag[5] X0_mag[6] X0_mag[7] X1_mag[0] X1_mag[1]
+ X1_mag[2] X1_mag[3] X1_mag[4] X1_mag[5] X1_mag[6] X1_mag[7] X2_mag[0] X2_mag[1]
+ X2_mag[2] X2_mag[3] X2_mag[4] X2_mag[5] X2_mag[6] X2_mag[7] X3_mag[0] X3_mag[1]
+ X3_mag[2] X3_mag[3] X3_mag[4] X3_mag[5] X3_mag[6] X3_mag[7] done
XFILL_22_0_2 gnd vdd FILL
XFILL_5_1_2 gnd vdd FILL
XAND2X2_5 AND2X2_5/A AND2X2_5/B gnd INVX1_50/A vdd AND2X2
XOAI21X1_360 INVX2_43/A NOR2X1_221/Y AND2X2_45/Y gnd AOI22X1_48/B vdd OAI21X1
XOAI21X1_371 OAI21X1_371/A OAI21X1_371/B NAND2X1_410/Y gnd NAND3X1_335/C vdd OAI21X1
XOAI21X1_382 AOI22X1_51/Y XNOR2X1_49/A AOI21X1_154/Y gnd OAI21X1_382/Y vdd OAI21X1
XFILL_13_0_2 gnd vdd FILL
XINVX1_221 INVX1_221/A gnd INVX1_221/Y vdd INVX1
XINVX1_232 gnd gnd INVX1_232/Y vdd INVX1
XOAI21X1_190 gnd INVX2_12/Y NOR2X1_119/Y gnd AOI22X1_7/D vdd OAI21X1
XINVX1_243 INVX1_243/A gnd INVX1_243/Y vdd INVX1
XINVX1_210 INVX1_210/A gnd INVX1_210/Y vdd INVX1
XNAND2X1_32 x2[0] INVX1_32/Y gnd AOI21X1_6/B vdd NAND2X1
XNAND2X1_21 OAI21X1_34/C NAND2X1_21/B gnd INVX1_40/A vdd NAND2X1
XINVX1_287 INVX1_287/A gnd INVX1_287/Y vdd INVX1
XNAND2X1_43 INVX1_273/A OR2X2_4/B gnd OAI21X1_77/C vdd NAND2X1
XINVX1_276 AND2X2_43/Y gnd INVX1_276/Y vdd INVX1
XNAND2X1_10 OR2X2_3/B BUFX4_12/Y gnd OAI21X1_11/C vdd NAND2X1
XINVX1_298 INVX1_298/A gnd INVX1_298/Y vdd INVX1
XINVX1_254 INVX1_254/A gnd INVX1_254/Y vdd INVX1
XINVX1_265 INVX1_265/A gnd INVX1_265/Y vdd INVX1
XNAND2X1_76 INVX1_116/A INVX1_80/Y gnd AND2X2_12/A vdd NAND2X1
XNAND2X1_65 NAND2X1_65/A NAND2X1_65/B gnd NOR2X1_95/B vdd NAND2X1
XNAND2X1_98 INVX2_23/A BUFX4_12/Y gnd NAND2X1_98/Y vdd NAND2X1
XNAND2X1_54 BUFX4_9/Y INVX1_63/A gnd OAI21X1_91/C vdd NAND2X1
XNAND2X1_87 INVX1_54/A INVX1_83/Y gnd NAND2X1_87/Y vdd NAND2X1
XAOI22X1_30 AOI22X1_30/A INVX1_248/A AOI22X1_31/C AOI22X1_31/D gnd AOI22X1_30/Y vdd
+ AOI22X1
XAOI22X1_41 AOI22X1_37/A AOI22X1_37/B AOI22X1_41/C AOI22X1_41/D gnd AOI22X1_41/Y vdd
+ AOI22X1
XAOI22X1_52 INVX2_36/A INVX1_99/A INVX2_37/A INVX1_98/A gnd AOI22X1_52/Y vdd AOI22X1
XNAND3X1_218 XNOR2X1_40/Y NAND3X1_212/Y NAND3X1_245/C gnd NAND3X1_218/Y vdd NAND3X1
XNAND3X1_229 NAND3X1_232/A NOR2X1_194/Y NAND3X1_232/B gnd NAND3X1_230/B vdd NAND3X1
XNAND3X1_207 INVX1_131/A INVX2_33/A INVX1_242/A gnd INVX1_261/A vdd NAND3X1
XOAI22X1_3 BUFX4_3/Y INVX1_41/Y AND2X2_3/Y OAI22X1_3/D gnd OAI22X1_3/Y vdd OAI22X1
XNAND2X1_409 OR2X2_32/A INVX1_296/A gnd AOI22X1_48/C vdd NAND2X1
XFILL_20_1_0 gnd vdd FILL
XINVX2_34 INVX2_34/A gnd INVX2_34/Y vdd INVX2
XINVX2_23 INVX2_23/A gnd INVX2_23/Y vdd INVX2
XINVX2_12 gnd gnd INVX2_12/Y vdd INVX2
XFILL_3_2_0 gnd vdd FILL
XOAI21X1_19 BUFX4_1/Y INVX2_3/Y OAI21X1_21/C gnd OAI21X1_19/Y vdd OAI21X1
XFILL_11_1_0 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XDFFPOSX1_103 INVX1_29/A CLKBUF1_1/Y OAI21X1_23/Y gnd vdd DFFPOSX1
XFILL_12_3 gnd vdd FILL
XDFFPOSX1_114 BUFX2_10/A DFFSR_1/CLK NOR2X1_132/Y gnd vdd DFFPOSX1
XDFFPOSX1_125 BUFX2_21/A CLKBUF1_6/Y NOR2X1_131/Y gnd vdd DFFPOSX1
XNAND2X1_239 NAND3X1_87/A NAND3X1_87/Y gnd INVX1_217/A vdd NAND2X1
XNAND2X1_217 INVX1_201/Y NOR2X1_148/Y gnd NOR3X1_7/A vdd NAND2X1
XNAND2X1_228 INVX1_219/A NAND3X1_92/B gnd NAND2X1_228/Y vdd NAND2X1
XDFFPOSX1_136 BUFX2_32/A CLKBUF1_6/Y NAND2X1_445/Y gnd vdd DFFPOSX1
XNAND2X1_206 AOI21X1_75/B OR2X2_16/Y gnd NAND2X1_207/B vdd NAND2X1
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XOR2X2_33 OR2X2_33/A OR2X2_33/B gnd OR2X2_33/Y vdd OR2X2
XOR2X2_11 OR2X2_11/A OR2X2_11/B gnd OR2X2_11/Y vdd OR2X2
XOR2X2_22 OR2X2_22/A OR2X2_22/B gnd OR2X2_22/Y vdd OR2X2
XXNOR2X1_6 AOI21X1_4/B AND2X2_2/B gnd XNOR2X1_6/Y vdd XNOR2X1
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 x1[2] gnd INVX1_6/Y vdd INVX1
XFILL_8_1_0 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XOAI21X1_361 INVX2_43/A NOR2X1_221/Y INVX1_296/Y gnd AOI22X1_49/C vdd OAI21X1
XAND2X2_6 OR2X2_4/B XOR2X1_5/A gnd AND2X2_6/Y vdd AND2X2
XOAI21X1_350 INVX2_37/Y INVX1_275/Y NOR2X1_218/Y gnd NAND3X1_278/B vdd OAI21X1
XOAI21X1_372 INVX1_295/A AOI21X1_149/Y NAND3X1_333/B gnd OAI21X1_372/Y vdd OAI21X1
XOAI21X1_383 OAI21X1_383/A NOR2X1_225/Y INVX1_307/Y gnd OAI21X1_383/Y vdd OAI21X1
XINVX1_277 INVX1_277/A gnd INVX1_277/Y vdd INVX1
XAOI22X1_1 BUFX4_14/Y INVX1_52/Y AOI22X1_1/C OR2X2_2/Y gnd AOI22X1_1/Y vdd AOI22X1
XINVX1_266 INVX1_266/A gnd INVX1_266/Y vdd INVX1
XINVX1_222 XOR2X1_16/Y gnd INVX1_222/Y vdd INVX1
XINVX1_244 OR2X2_22/Y gnd INVX1_244/Y vdd INVX1
XINVX1_233 INVX1_233/A gnd INVX1_233/Y vdd INVX1
XOAI21X1_191 INVX1_180/A AND2X2_22/Y INVX1_163/A gnd AOI22X1_8/B vdd OAI21X1
XINVX1_255 INVX1_255/A gnd INVX1_255/Y vdd INVX1
XINVX1_211 INVX1_211/A gnd INVX1_211/Y vdd INVX1
XOAI21X1_180 INVX1_141/Y INVX1_150/Y AND2X2_20/B gnd INVX1_155/A vdd OAI21X1
XINVX1_200 INVX1_200/A gnd INVX1_200/Y vdd INVX1
XNAND2X1_33 AOI21X1_8/Y OAI21X1_48/Y gnd NAND2X1_33/Y vdd NAND2X1
XINVX1_288 INVX1_288/A gnd INVX1_288/Y vdd INVX1
XNAND2X1_11 NOR2X1_5/Y NOR2X1_9/Y gnd NAND2X1_11/Y vdd NAND2X1
XNAND2X1_44 INVX2_2/Y NOR2X1_58/Y gnd NAND2X1_45/B vdd NAND2X1
XINVX1_299 INVX1_99/A gnd INVX1_299/Y vdd INVX1
XNAND2X1_77 INVX1_80/A INVX1_116/Y gnd NAND3X1_9/C vdd NAND2X1
XNAND2X1_22 INVX1_112/A BUFX4_16/Y gnd NAND2X1_22/Y vdd NAND2X1
XNAND2X1_66 INVX1_112/A INVX1_111/Y gnd NAND2X1_68/A vdd NAND2X1
XNAND2X1_55 BUFX4_5/Y INVX1_65/A gnd NAND2X1_55/Y vdd NAND2X1
XNAND2X1_99 INVX1_193/A BUFX4_12/Y gnd NAND2X1_99/Y vdd NAND2X1
XNAND2X1_88 INVX1_152/A BUFX4_10/Y gnd NAND2X1_88/Y vdd NAND2X1
XAOI22X1_53 AND2X2_44/Y AOI22X1_53/B XOR2X1_21/B XOR2X1_21/A gnd AOI22X1_53/Y vdd
+ AOI22X1
XAOI22X1_42 INVX2_36/A NOR2X1_206/Y INVX1_274/A AOI22X1_42/D gnd OR2X2_29/B vdd AOI22X1
XAOI22X1_31 AOI22X1_31/A AOI22X1_31/B AOI22X1_31/C AOI22X1_31/D gnd OR2X2_24/A vdd
+ AOI22X1
XAOI22X1_20 AOI22X1_20/A NAND3X1_86/Y INVX1_218/A AOI22X1_18/A gnd AOI22X1_20/Y vdd
+ AOI22X1
XNAND3X1_219 XNOR2X1_39/Y NAND3X1_214/Y NAND3X1_215/Y gnd NAND3X1_219/Y vdd NAND3X1
XNAND3X1_208 AND2X2_38/Y INVX1_261/A INVX1_260/Y gnd AND2X2_39/B vdd NAND3X1
XOAI22X1_4 BUFX4_3/Y INVX1_47/Y OAI22X1_4/C OAI22X1_4/D gnd OAI22X1_4/Y vdd OAI22X1
XFILL_20_1_1 gnd vdd FILL
XINVX2_35 INVX2_35/A gnd INVX2_35/Y vdd INVX2
XINVX2_24 NOR3X1_7/A gnd INVX2_24/Y vdd INVX2
XINVX2_13 INVX2_13/A gnd INVX2_13/Y vdd INVX2
XFILL_3_2_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_19_2_1 gnd vdd FILL
XDFFPOSX1_104 INVX1_30/A CLKBUF1_4/Y OAI21X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_115 BUFX2_11/A CLKBUF1_10/Y XNOR2X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_126 BUFX2_22/A CLKBUF1_6/Y XNOR2X1_22/Y gnd vdd DFFPOSX1
XNAND2X1_218 INVX2_19/A INVX1_104/A gnd INVX1_205/A vdd NAND2X1
XNAND2X1_229 NAND2X1_229/A OR2X2_20/B gnd INVX1_209/A vdd NAND2X1
XNAND2X1_207 INVX1_196/A NAND2X1_207/B gnd AOI21X1_72/B vdd NAND2X1
XFILL_10_1 gnd vdd FILL
XOR2X2_34 OR2X2_34/A OR2X2_34/B gnd OR2X2_34/Y vdd OR2X2
XOR2X2_23 OR2X2_23/A OR2X2_23/B gnd OR2X2_23/Y vdd OR2X2
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XOR2X2_12 OR2X2_12/A OR2X2_12/B gnd OR2X2_12/Y vdd OR2X2
XXNOR2X1_7 XNOR2X1_7/A AND2X2_2/A gnd XNOR2X1_7/Y vdd XNOR2X1
XFILL_0_0_1 gnd vdd FILL
XINVX1_7 x3[2] gnd INVX1_7/Y vdd INVX1
XFILL_8_1_1 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XAND2X2_7 AND2X2_7/A AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XOAI21X1_351 INVX2_42/Y INVX1_289/Y NAND2X1_391/Y gnd NAND3X1_279/B vdd OAI21X1
XOAI21X1_373 INVX2_43/A NOR2X1_221/Y INVX2_41/A gnd OAI21X1_373/Y vdd OAI21X1
XOAI21X1_362 INVX2_43/A NOR2X1_221/Y OAI21X1_362/C gnd AOI22X1_49/B vdd OAI21X1
XOAI21X1_384 INVX2_43/A OAI21X1_362/C OR2X2_32/Y gnd XOR2X1_25/A vdd OAI21X1
XOAI21X1_340 INVX2_37/A INVX1_275/Y INVX1_278/A gnd NAND3X1_273/A vdd OAI21X1
XNAND2X1_390 INVX2_37/A INVX1_96/A gnd INVX1_290/A vdd NAND2X1
XAOI22X1_2 BUFX4_11/Y AOI22X1_2/B AOI22X1_2/C AOI22X1_2/D gnd AOI22X1_2/Y vdd AOI22X1
XINVX1_289 INVX1_289/A gnd INVX1_289/Y vdd INVX1
XINVX1_278 INVX1_278/A gnd INVX1_278/Y vdd INVX1
XINVX1_212 INVX1_212/A gnd INVX1_212/Y vdd INVX1
XINVX1_245 INVX1_245/A gnd INVX1_245/Y vdd INVX1
XINVX1_267 INVX1_267/A gnd INVX1_267/Y vdd INVX1
XINVX1_256 INVX1_256/A gnd INVX1_256/Y vdd INVX1
XINVX1_223 XOR2X1_14/Y gnd INVX1_223/Y vdd INVX1
XINVX1_234 INVX1_234/A gnd INVX1_234/Y vdd INVX1
XOAI21X1_192 INVX1_180/A AND2X2_22/Y INVX1_164/Y gnd AOI22X1_8/C vdd OAI21X1
XOAI21X1_170 INVX2_8/Y INVX1_142/Y XNOR2X1_19/Y gnd AND2X2_20/A vdd OAI21X1
XINVX1_201 INVX1_201/A gnd INVX1_201/Y vdd INVX1
XOAI21X1_181 INVX2_9/Y INVX2_13/A INVX1_146/A gnd NAND2X1_140/A vdd OAI21X1
XNAND2X1_45 NAND2X1_45/A NAND2X1_45/B gnd NAND2X1_45/Y vdd NAND2X1
XNAND2X1_12 INVX1_79/A NOR2X1_13/B gnd OAI21X1_13/C vdd NAND2X1
XNAND2X1_67 INVX1_111/A INVX1_112/Y gnd NAND2X1_68/B vdd NAND2X1
XNAND2X1_34 INVX1_110/A BUFX4_15/Y gnd NAND2X1_34/Y vdd NAND2X1
XNAND2X1_23 INVX1_114/A BUFX4_16/Y gnd OAI21X1_37/C vdd NAND2X1
XNAND2X1_56 BUFX4_1/Y INVX1_66/A gnd OAI21X1_93/C vdd NAND2X1
XNAND2X1_89 NOR2X1_75/Y NOR2X1_85/Y gnd INVX1_121/A vdd NAND2X1
XNAND2X1_78 INVX2_9/A BUFX4_11/Y gnd NAND2X1_78/Y vdd NAND2X1
XAOI22X1_43 AOI22X1_46/A AOI22X1_46/B AOI22X1_43/C AOI22X1_43/D gnd AOI22X1_43/Y vdd
+ AOI22X1
XAOI22X1_54 NOR2X1_219/A AOI22X1_53/B AOI22X1_54/C OR2X2_34/A gnd AOI22X1_54/Y vdd
+ AOI22X1
XAOI22X1_32 INVX1_248/A AOI22X1_30/A AOI22X1_29/C AOI22X1_32/D gnd AOI22X1_32/Y vdd
+ AOI22X1
XAOI22X1_21 INVX2_21/A INVX1_193/A INVX1_187/A AOI22X1_21/D gnd INVX2_25/A vdd AOI22X1
XAOI22X1_10 INVX2_10/A INVX1_152/A INVX1_139/A INVX1_153/A gnd INVX1_170/A vdd AOI22X1
XNAND3X1_209 NAND3X1_203/Y NAND3X1_206/Y AND2X2_39/Y gnd NAND3X1_245/C vdd NAND3X1
XOAI22X1_5 BUFX4_3/Y INVX1_75/Y OAI22X1_5/C INVX1_76/Y gnd OAI22X1_5/Y vdd OAI22X1
XFILL_20_1_2 gnd vdd FILL
XINVX2_36 INVX2_36/A gnd INVX2_36/Y vdd INVX2
XINVX2_25 INVX2_25/A gnd INVX2_25/Y vdd INVX2
XINVX2_14 INVX2_14/A gnd INVX2_14/Y vdd INVX2
XFILL_3_2_2 gnd vdd FILL
XFILL_11_1_2 gnd vdd FILL
XFILL_19_2_2 gnd vdd FILL
XDFFPOSX1_116 BUFX2_12/A CLKBUF1_10/Y NOR2X1_141/Y gnd vdd DFFPOSX1
XDFFPOSX1_127 BUFX2_23/A CLKBUF1_6/Y XNOR2X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_105 BUFX2_1/A DFFSR_1/CLK NOR2X1_165/Y gnd vdd DFFPOSX1
XNAND2X1_219 NAND3X1_87/A NAND3X1_87/B gnd OAI21X1_235/C vdd NAND2X1
XNAND2X1_208 NAND2X1_207/B INVX1_196/Y gnd NAND3X1_84/C vdd NAND2X1
XINVX8_1 BUFX4_3/Y gnd INVX8_1/Y vdd INVX8
XBUFX4_10 INVX8_1/Y gnd BUFX4_10/Y vdd BUFX4
XFILL_10_2 gnd vdd FILL
XXNOR2X1_8 XNOR2X1_8/A INVX1_60/A gnd XNOR2X1_8/Y vdd XNOR2X1
XOR2X2_24 OR2X2_24/A OR2X2_24/B gnd OR2X2_24/Y vdd OR2X2
XOR2X2_13 OR2X2_13/A OR2X2_13/B gnd OR2X2_13/Y vdd OR2X2
XOR2X2_6 BUFX4_4/Y OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XFILL_0_0_2 gnd vdd FILL
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_8_1_2 gnd vdd FILL
XFILL_16_0_2 gnd vdd FILL
XFILL_9_1 gnd vdd FILL
XOAI21X1_341 INVX2_35/Y INVX1_279/Y NAND2X1_371/Y gnd OAI21X1_341/Y vdd OAI21X1
XOAI21X1_330 AOI22X1_37/Y AOI22X1_38/Y OAI21X1_330/C gnd OAI21X1_330/Y vdd OAI21X1
XOAI21X1_363 NOR3X1_12/Y AOI21X1_142/Y INVX1_297/A gnd OAI21X1_363/Y vdd OAI21X1
XOAI21X1_352 AOI22X1_43/Y AOI22X1_44/Y OAI21X1_355/C gnd INVX1_305/A vdd OAI21X1
XOAI21X1_374 INVX2_39/Y OAI21X1_373/Y OAI21X1_374/C gnd XOR2X1_22/B vdd OAI21X1
XAND2X2_8 AND2X2_8/A AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XOAI21X1_385 AOI21X1_158/Y OAI21X1_385/B XOR2X1_25/Y gnd NAND3X1_356/C vdd OAI21X1
XNAND2X1_380 NAND2X1_380/A INVX1_282/Y gnd NAND2X1_380/Y vdd NAND2X1
XNAND2X1_391 NAND2X1_391/A NAND3X1_278/B gnd NAND2X1_391/Y vdd NAND2X1
XAOI22X1_3 BUFX4_10/Y AOI22X1_3/B AOI22X1_3/C AOI22X1_3/D gnd AOI22X1_3/Y vdd AOI22X1
XOAI21X1_171 INVX2_8/Y INVX1_142/Y NOR2X1_111/Y gnd AND2X2_19/B vdd OAI21X1
XOAI21X1_182 INVX1_139/A INVX1_152/Y OAI21X1_182/C gnd NAND3X1_20/C vdd OAI21X1
XOAI21X1_160 NOR2X1_99/Y AND2X2_17/Y BUFX4_5/Y gnd AND2X2_18/A vdd OAI21X1
XINVX1_279 INVX1_279/A gnd INVX1_279/Y vdd INVX1
XINVX1_224 INVX1_224/A gnd INVX1_224/Y vdd INVX1
XINVX1_235 INVX1_235/A gnd INVX1_235/Y vdd INVX1
XINVX1_246 INVX1_246/A gnd INVX1_246/Y vdd INVX1
XINVX1_257 INVX1_257/A gnd INVX1_257/Y vdd INVX1
XINVX1_268 INVX1_268/A gnd INVX1_268/Y vdd INVX1
XINVX1_213 INVX1_107/A gnd INVX1_213/Y vdd INVX1
XOAI21X1_193 NOR3X1_2/B NOR3X1_2/C NOR3X1_2/A gnd AOI21X1_56/B vdd OAI21X1
XINVX1_202 INVX1_202/A gnd INVX1_202/Y vdd INVX1
XNAND2X1_24 INVX1_60/A INVX1_45/A gnd NAND2X1_24/Y vdd NAND2X1
XNAND2X1_13 BUFX4_8/Y OAI21X1_13/C gnd OAI22X1_2/D vdd NAND2X1
XNAND2X1_46 INVX2_39/A OR2X2_4/B gnd OAI21X1_79/C vdd NAND2X1
XNAND2X1_35 INVX1_111/A BUFX4_15/Y gnd OAI21X1_62/C vdd NAND2X1
XNAND2X1_79 AND2X2_12/A NAND3X1_9/C gnd NOR2X1_66/B vdd NAND2X1
XNAND2X1_68 NAND2X1_68/A NAND2X1_68/B gnd NAND2X1_68/Y vdd NAND2X1
XNAND2X1_57 BUFX4_1/Y INVX1_67/A gnd NAND2X1_57/Y vdd NAND2X1
XAOI22X1_44 AOI22X1_46/D INVX1_304/A AOI22X1_44/C OR2X2_31/Y gnd AOI22X1_44/Y vdd
+ AOI22X1
XNOR3X1_1 INVX1_29/A NOR3X1_1/B NOR3X1_1/C gnd OR2X2_4/A vdd NOR3X1
XAOI22X1_33 gnd gnd gnd gnd gnd NOR3X1_8/A vdd AOI22X1
XAOI22X1_11 AOI22X1_11/A AOI22X1_11/B AOI22X1_11/C AOI22X1_11/D gnd AOI22X1_11/Y vdd
+ AOI22X1
XAOI22X1_22 NAND3X1_99/Y AOI22X1_22/B AOI22X1_22/C AOI22X1_22/D gnd NOR3X1_7/B vdd
+ AOI22X1
XFILL_23_1_0 gnd vdd FILL
XOAI22X1_6 BUFX4_3/Y INVX1_80/Y OAI22X1_6/C OAI22X1_6/D gnd OAI22X1_6/Y vdd OAI22X1
XFILL_6_2_0 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XINVX2_26 INVX2_26/A gnd INVX2_26/Y vdd INVX2
XINVX2_15 INVX2_15/A gnd INVX2_15/Y vdd INVX2
XINVX2_37 INVX2_37/A gnd INVX2_37/Y vdd INVX2
XDFFPOSX1_117 BUFX2_13/A CLKBUF1_4/Y NOR2X1_162/Y gnd vdd DFFPOSX1
XDFFPOSX1_128 BUFX2_24/A CLKBUF1_6/Y NAND2X1_189/Y gnd vdd DFFPOSX1
XDFFPOSX1_106 BUFX2_2/A DFFSR_1/CLK NOR2X1_163/Y gnd vdd DFFPOSX1
XNAND2X1_209 INVX1_196/A XOR2X1_12/Y gnd NAND3X1_84/B vdd NAND2X1
XNOR2X1_220 INVX1_293/Y AOI22X1_46/B gnd INVX1_294/A vdd NOR2X1
XFILL_3_0_0 gnd vdd FILL
XBUFX4_11 INVX8_1/Y gnd BUFX4_11/Y vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XNAND3X1_360 AOI21X1_163/Y NAND3X1_360/B NAND3X1_360/C gnd NAND3X1_360/Y vdd NAND3X1
XOR2X2_14 OR2X2_14/A XOR2X1_9/A gnd OR2X2_14/Y vdd OR2X2
XFILL_10_3 gnd vdd FILL
XXNOR2X1_9 XNOR2X1_9/A INVX1_53/A gnd XNOR2X1_9/Y vdd XNOR2X1
XOR2X2_7 BUFX4_7/Y DFFSR_1/Q gnd OR2X2_7/Y vdd OR2X2
XOR2X2_25 OR2X2_25/A OR2X2_25/B gnd OR2X2_25/Y vdd OR2X2
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XFILL_9_2 gnd vdd FILL
XNAND3X1_190 NAND3X1_194/A NAND3X1_190/B NAND3X1_189/Y gnd NAND2X1_312/A vdd NAND3X1
XOAI21X1_364 NOR3X1_12/B NOR3X1_12/C INVX2_42/A gnd NAND3X1_326/B vdd OAI21X1
XOAI21X1_353 AOI22X1_46/Y AOI22X1_45/Y OAI21X1_353/C gnd NAND3X1_281/C vdd OAI21X1
XOAI21X1_342 INVX2_35/Y INVX1_279/Y NOR2X1_210/Y gnd OAI21X1_342/Y vdd OAI21X1
XOAI21X1_331 AOI22X1_39/Y AOI21X1_133/Y NAND2X1_338/A gnd OAI21X1_332/C vdd OAI21X1
XOAI21X1_320 INVX1_257/A NOR2X1_196/Y OAI21X1_320/C gnd OAI21X1_320/Y vdd OAI21X1
XOAI21X1_386 INVX1_297/Y AOI21X1_142/Y NAND3X1_326/C gnd INVX1_311/A vdd OAI21X1
XAND2X2_9 OR2X2_4/B XOR2X1_5/B gnd AND2X2_9/Y vdd AND2X2
XXOR2X1_20 OR2X2_29/A OR2X2_29/B gnd XOR2X1_20/Y vdd XOR2X1
XOAI21X1_375 OAI21X1_375/A OAI21X1_375/B NAND3X1_302/Y gnd OR2X2_33/A vdd OAI21X1
XNAND2X1_392 NAND3X1_279/B NAND3X1_279/C gnd NAND2X1_395/B vdd NAND2X1
XNAND2X1_381 INVX1_282/A XOR2X1_20/Y gnd NAND3X1_275/B vdd NAND2X1
XNAND2X1_370 INVX2_36/A INVX1_96/A gnd INVX1_278/A vdd NAND2X1
XINVX1_214 INVX1_214/A gnd INVX1_214/Y vdd INVX1
XINVX1_225 INVX1_225/A gnd INVX1_225/Y vdd INVX1
XOAI21X1_172 INVX1_144/Y gnd NOR2X1_110/Y gnd AND2X2_19/A vdd OAI21X1
XINVX1_203 INVX1_203/A gnd INVX1_203/Y vdd INVX1
XAOI22X1_4 BUFX4_11/Y INVX1_131/Y AOI22X1_4/C OR2X2_5/Y gnd AOI22X1_4/Y vdd AOI22X1
XOAI21X1_194 INVX1_154/A NAND2X1_145/Y AND2X2_21/B gnd INVX1_173/A vdd OAI21X1
XOAI21X1_183 INVX2_10/Y INVX1_153/Y OAI21X1_183/C gnd AND2X2_21/A vdd OAI21X1
XOAI21X1_150 BUFX4_13/Y XNOR2X1_15/Y OAI21X1_150/C gnd DFFPOSX1_2/D vdd OAI21X1
XOAI21X1_161 NOR2X1_100/Y AND2X2_17/Y INVX1_128/Y gnd AOI22X1_5/C vdd OAI21X1
XNAND2X1_14 INVX1_90/A BUFX4_14/Y gnd OAI21X1_14/C vdd NAND2X1
XNAND2X1_25 x2[6] INVX1_48/Y gnd AND2X2_5/A vdd NAND2X1
XINVX1_247 INVX1_247/A gnd INVX1_247/Y vdd INVX1
XINVX1_236 INVX1_236/A gnd INVX1_236/Y vdd INVX1
XINVX1_269 INVX1_269/A gnd INVX1_269/Y vdd INVX1
XINVX1_258 OR2X2_6/B gnd INVX1_258/Y vdd INVX1
XNAND2X1_47 INVX2_41/A OR2X2_4/B gnd OAI21X1_81/C vdd NAND2X1
XNAND2X1_36 NOR2X1_5/Y AND2X2_8/Y gnd INVX1_76/A vdd NAND2X1
XNAND2X1_58 BUFX4_1/Y INVX1_68/A gnd OAI21X1_95/C vdd NAND2X1
XNAND2X1_69 INVX1_41/A INVX1_75/Y gnd NAND2X1_69/Y vdd NAND2X1
XAOI22X1_23 AOI22X1_23/A AOI22X1_23/B AOI22X1_23/C AOI22X1_23/D gnd NOR3X1_7/C vdd
+ AOI22X1
XAOI22X1_12 AOI22X1_12/A AOI22X1_12/B AOI22X1_12/C AOI22X1_12/D gnd AOI22X1_12/Y vdd
+ AOI22X1
XAOI22X1_45 AOI22X1_43/D AOI22X1_43/C AOI22X1_44/C OR2X2_31/Y gnd AOI22X1_45/Y vdd
+ AOI22X1
XAOI22X1_34 AND2X2_36/B AND2X2_36/A AOI22X1_34/C AOI22X1_34/D gnd NOR3X1_9/B vdd AOI22X1
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd NOR3X1_3/B vdd NOR3X1
XFILL_23_1_1 gnd vdd FILL
XOAI22X1_7 OAI22X1_7/A OAI22X1_7/B OAI22X1_9/C OAI22X1_9/D gnd OAI22X1_7/Y vdd OAI22X1
XFILL_6_2_1 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XINVX2_38 INVX2_38/A gnd INVX2_38/Y vdd INVX2
XINVX2_27 gnd gnd INVX2_27/Y vdd INVX2
XINVX2_16 INVX2_16/A gnd INVX2_16/Y vdd INVX2
XCLKBUF1_1 clk gnd CLKBUF1_1/Y vdd CLKBUF1
XDFFPOSX1_118 BUFX2_14/A CLKBUF1_2/Y XOR2X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_129 BUFX2_25/A CLKBUF1_6/Y NOR2X1_201/Y gnd vdd DFFPOSX1
XDFFPOSX1_107 BUFX2_3/A CLKBUF1_3/Y XNOR2X1_38/Y gnd vdd DFFPOSX1
XNOR2X1_221 OR2X2_32/A OR2X2_32/B gnd NOR2X1_221/Y vdd NOR2X1
XNOR2X1_210 INVX1_273/A INVX2_39/Y gnd NOR2X1_210/Y vdd NOR2X1
XFILL_3_0_1 gnd vdd FILL
XFILL_19_0_1 gnd vdd FILL
XBUFX4_12 INVX8_1/Y gnd BUFX4_12/Y vdd BUFX4
XNAND3X1_350 OAI22X1_21/Y OAI21X1_377/Y AND2X2_48/Y gnd NAND2X1_435/B vdd NAND3X1
XNAND3X1_361 OAI21X1_390/Y OR2X2_34/Y OAI21X1_392/C gnd NAND3X1_361/Y vdd NAND3X1
XOR2X2_15 OR2X2_15/A OR2X2_15/B gnd OR2X2_15/Y vdd OR2X2
XOR2X2_26 OR2X2_26/A OR2X2_26/B gnd OR2X2_26/Y vdd OR2X2
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XFILL_9_3 gnd vdd FILL
XNAND3X1_191 INVX1_234/Y NAND3X1_191/B INVX1_264/A gnd NAND3X1_194/B vdd NAND3X1
XNAND3X1_180 INVX2_28/A INVX1_131/A NOR2X1_176/Y gnd NAND3X1_180/Y vdd NAND3X1
XOAI21X1_354 AOI22X1_43/Y AOI22X1_44/Y OAI21X1_353/C gnd NAND3X1_282/B vdd OAI21X1
XOAI21X1_343 INVX2_39/Y INVX1_273/A NOR2X1_209/Y gnd NAND2X1_373/B vdd OAI21X1
XOAI21X1_365 INVX1_290/A INVX2_44/A AOI22X1_51/D gnd XNOR2X1_47/A vdd OAI21X1
XOAI21X1_387 NAND2X1_423/Y OAI21X1_371/B NAND3X1_325/B gnd OAI21X1_387/Y vdd OAI21X1
XOAI21X1_376 INVX2_44/A AOI22X1_52/Y NAND3X1_298/C gnd OAI21X1_376/Y vdd OAI21X1
XOAI21X1_321 NAND2X1_333/Y OAI21X1_321/B NAND3X1_203/Y gnd OAI21X1_321/Y vdd OAI21X1
XOAI21X1_310 AOI21X1_109/Y NOR3X1_9/Y INVX1_254/Y gnd OAI21X1_310/Y vdd OAI21X1
XOAI21X1_332 AOI22X1_40/Y AOI22X1_41/Y OAI21X1_332/C gnd NAND2X1_360/B vdd OAI21X1
XXOR2X1_21 XOR2X1_21/A XOR2X1_21/B gnd XOR2X1_21/Y vdd XOR2X1
XXOR2X1_10 XOR2X1_10/A XOR2X1_10/B gnd XOR2X1_10/Y vdd XOR2X1
XNAND2X1_382 INVX1_273/A INVX1_279/A gnd INVX1_286/A vdd NAND2X1
XNAND2X1_393 INVX1_288/A NAND2X1_395/B gnd AOI22X1_43/D vdd NAND2X1
XNAND2X1_371 NAND3X1_273/A NAND2X1_387/A gnd NAND2X1_371/Y vdd NAND2X1
XNAND2X1_360 OAI21X1_330/Y NAND2X1_360/B gnd NAND2X1_360/Y vdd NAND2X1
XOAI21X1_184 NOR3X1_6/B NOR3X1_6/C NOR3X1_6/A gnd AOI21X1_67/B vdd OAI21X1
XOAI21X1_162 INVX2_9/A INVX2_10/Y NOR2X1_105/Y gnd INVX1_135/A vdd OAI21X1
XINVX1_248 INVX1_248/A gnd OR2X2_24/B vdd INVX1
XINVX1_215 INVX1_215/A gnd INVX1_215/Y vdd INVX1
XOAI21X1_173 INVX1_136/A INVX1_143/A OR2X2_10/A gnd OAI21X1_173/Y vdd OAI21X1
XINVX1_259 INVX1_259/A gnd INVX1_259/Y vdd INVX1
XINVX1_237 INVX1_237/A gnd INVX1_237/Y vdd INVX1
XINVX1_226 INVX1_226/A gnd INVX1_226/Y vdd INVX1
XINVX1_204 INVX1_105/A gnd INVX1_204/Y vdd INVX1
XOAI21X1_195 INVX2_9/Y INVX2_16/Y INVX1_153/Y gnd AND2X2_24/B vdd OAI21X1
XOAI21X1_151 NOR2X1_97/A INVX1_130/Y AOI21X1_33/Y gnd XNOR2X1_16/A vdd OAI21X1
XAOI22X1_5 BUFX4_10/Y INVX1_132/Y AOI22X1_5/C AOI22X1_5/D gnd AOI22X1_5/Y vdd AOI22X1
XOAI21X1_140 BUFX4_13/Y INVX2_4/Y NAND2X1_100/Y gnd DFFPOSX1_22/D vdd OAI21X1
XNAND2X1_26 x0[6] INVX1_49/Y gnd AND2X2_5/B vdd NAND2X1
XNAND2X1_15 OAI21X1_27/Y NAND2X1_15/B gnd OAI21X1_29/B vdd NAND2X1
XNAND2X1_48 NOR2X1_60/Y NOR2X1_61/Y gnd INVX1_91/A vdd NAND2X1
XNAND2X1_59 BUFX4_1/Y INVX1_69/A gnd NAND2X1_59/Y vdd NAND2X1
XNAND2X1_37 INVX1_113/A BUFX4_16/Y gnd NAND2X1_37/Y vdd NAND2X1
XNAND2X1_190 INVX1_187/A INVX2_17/Y gnd XNOR2X1_31/B vdd NAND2X1
XAOI22X1_46 AOI22X1_46/A AOI22X1_46/B INVX1_304/A AOI22X1_46/D gnd AOI22X1_46/Y vdd
+ AOI22X1
XAOI22X1_24 INVX2_19/A INVX1_105/A INVX1_104/A INVX1_103/A gnd OAI22X1_18/D vdd AOI22X1
XAOI22X1_35 INVX2_29/A INVX1_242/A INVX1_131/A INVX2_33/A gnd INVX1_255/A vdd AOI22X1
XAOI22X1_13 AOI22X1_13/A AOI22X1_13/B AOI22X1_13/C AOI22X1_13/D gnd NOR3X1_5/C vdd
+ AOI22X1
XNOR3X1_3 INVX2_15/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XFILL_23_1_2 gnd vdd FILL
XOAI22X1_8 INVX2_14/Y OAI22X1_9/B OAI22X1_8/C OAI22X1_8/D gnd OAI22X1_8/Y vdd OAI22X1
XFILL_6_2_2 gnd vdd FILL
XFILL_14_1_2 gnd vdd FILL
XAOI21X1_90 INVX2_25/Y INVX2_23/A NOR2X1_154/Y gnd AOI21X1_90/Y vdd AOI21X1
XFILL_19_1 gnd vdd FILL
XINVX2_39 INVX2_39/A gnd INVX2_39/Y vdd INVX2
XINVX2_28 INVX2_28/A gnd INVX2_28/Y vdd INVX2
XINVX2_17 INVX2_17/A gnd INVX2_17/Y vdd INVX2
XDFFPOSX1_119 BUFX2_15/A CLKBUF1_2/Y XNOR2X1_35/Y gnd vdd DFFPOSX1
XDFFPOSX1_108 BUFX2_4/A DFFSR_1/CLK NOR2X1_175/Y gnd vdd DFFPOSX1
XCLKBUF1_2 clk gnd CLKBUF1_2/Y vdd CLKBUF1
XNOR2X1_222 INVX2_39/A INVX2_41/Y gnd INVX1_296/A vdd NOR2X1
XNOR2X1_211 NOR2X1_211/A INVX1_280/Y gnd INVX1_281/A vdd NOR2X1
XNOR2X1_200 INVX2_35/A INVX2_36/A gnd NOR2X1_201/A vdd NOR2X1
XFILL_3_0_2 gnd vdd FILL
XDFFPOSX1_90 INVX1_4/A CLKBUF1_2/Y OAI21X1_4/Y gnd vdd DFFPOSX1
XFILL_19_0_2 gnd vdd FILL
XBUFX4_13 INVX8_1/Y gnd BUFX4_13/Y vdd BUFX4
XNAND3X1_340 AOI21X1_146/Y NAND3X1_343/B NAND3X1_343/C gnd AOI22X1_54/C vdd NAND3X1
XNAND3X1_362 NAND3X1_362/A OAI22X1_22/Y NAND3X1_361/Y gnd NAND3X1_362/Y vdd NAND3X1
XNAND3X1_351 INVX1_307/A NAND2X1_434/Y NAND3X1_351/C gnd NAND3X1_351/Y vdd NAND3X1
XOR2X2_9 OR2X2_9/A OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XOR2X2_27 OR2X2_27/A OR2X2_27/B gnd OR2X2_27/Y vdd OR2X2
XOR2X2_16 OR2X2_16/A OR2X2_16/B gnd OR2X2_16/Y vdd OR2X2
XFILL_21_2_0 gnd vdd FILL
XFILL_12_2_0 gnd vdd FILL
XNAND3X1_192 INVX1_234/A NAND3X1_189/B NAND3X1_189/C gnd NAND3X1_194/C vdd NAND3X1
XNAND3X1_181 OAI21X1_283/Y XOR2X1_17/A NAND3X1_180/Y gnd NAND2X1_287/A vdd NAND3X1
XNAND3X1_170 OAI21X1_273/Y OR2X2_20/Y NAND3X1_170/C gnd NAND3X1_170/Y vdd NAND3X1
XOAI21X1_355 AOI22X1_46/Y AOI22X1_45/Y OAI21X1_355/C gnd NAND3X1_282/C vdd OAI21X1
XOAI21X1_344 NOR2X1_219/A NOR2X1_219/B AND2X2_44/B gnd OAI21X1_344/Y vdd OAI21X1
XOAI21X1_377 INVX2_41/Y INVX2_43/A OR2X2_32/Y gnd OAI21X1_377/Y vdd OAI21X1
XOAI21X1_333 INVX1_273/Y INVX2_38/Y INVX2_40/Y gnd AND2X2_43/A vdd OAI21X1
XOAI21X1_366 INVX2_36/Y INVX1_299/Y NOR2X1_224/B gnd NAND3X1_298/B vdd OAI21X1
XOAI21X1_388 OAI21X1_389/A INVX1_310/Y NAND2X1_441/Y gnd NAND3X1_358/B vdd OAI21X1
XOAI21X1_300 NOR3X1_8/A NOR3X1_8/C NOR3X1_8/B gnd INVX1_252/A vdd OAI21X1
XOAI21X1_322 NOR3X1_11/B NOR3X1_11/C INVX1_270/A gnd OAI21X1_322/Y vdd OAI21X1
XOAI21X1_311 OAI21X1_312/A OAI21X1_312/B NAND2X1_337/Y gnd NAND3X1_231/C vdd OAI21X1
XNAND2X1_372 NAND2X1_372/A OAI21X1_341/Y gnd OR2X2_29/A vdd NAND2X1
XXOR2X1_22 XOR2X1_22/A XOR2X1_22/B gnd INVX1_309/A vdd XOR2X1
XNAND2X1_361 NAND3X1_184/Y NAND2X1_361/B gnd NOR2X1_197/B vdd NAND2X1
XXOR2X1_11 XOR2X1_11/A XOR2X1_10/B gnd XOR2X1_11/Y vdd XOR2X1
XNAND2X1_350 NAND2X1_343/Y AOI21X1_122/Y gnd NAND2X1_351/A vdd NAND2X1
XNAND2X1_394 OR2X2_31/B OR2X2_31/A gnd AOI22X1_44/C vdd NAND2X1
XNAND2X1_383 INVX2_35/A AOI22X1_47/D gnd INVX1_287/A vdd NAND2X1
XFILL_7_1 gnd vdd FILL
XNAND3X1_1 BUFX4_2/Y NAND3X1_1/B OAI21X1_5/C gnd OAI21X1_4/C vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XOAI21X1_130 BUFX4_10/Y XNOR2X1_14/Y NAND2X1_90/Y gnd OAI21X1_130/Y vdd OAI21X1
XOAI21X1_141 BUFX4_12/Y INVX1_29/Y NAND2X1_101/Y gnd DFFPOSX1_23/D vdd OAI21X1
XAOI22X1_6 AOI22X1_6/A AOI22X1_6/B AOI22X1_6/C AOI22X1_6/D gnd AOI22X1_6/Y vdd AOI22X1
XOAI21X1_185 NOR2X1_112/Y INVX2_11/Y OR2X2_9/Y gnd NAND3X1_33/C vdd OAI21X1
XOAI21X1_174 NOR2X1_112/Y INVX2_11/Y AOI22X1_6/C gnd AOI21X1_43/A vdd OAI21X1
XINVX1_249 NOR3X1_8/Y gnd INVX1_249/Y vdd INVX1
XINVX1_216 INVX1_216/A gnd INVX1_216/Y vdd INVX1
XOAI21X1_163 INVX1_134/Y INVX1_136/A OR2X2_8/B gnd AOI21X1_41/C vdd OAI21X1
XINVX1_205 INVX1_205/A gnd INVX1_205/Y vdd INVX1
XINVX1_238 INVX1_238/A gnd INVX1_238/Y vdd INVX1
XINVX1_227 gnd gnd INVX1_227/Y vdd INVX1
XOAI21X1_152 BUFX4_11/Y XNOR2X1_16/Y OAI21X1_152/C gnd DFFPOSX1_3/D vdd OAI21X1
XOAI21X1_196 INVX2_16/Y XOR2X1_6/B AND2X2_24/B gnd NOR2X1_121/B vdd OAI21X1
XNAND2X1_49 INVX1_279/A BUFX4_14/Y gnd OAI21X1_83/C vdd NAND2X1
XNAND2X1_27 INVX1_50/Y NOR2X1_30/B gnd OR2X2_2/A vdd NAND2X1
XNAND2X1_38 INVX1_79/A NOR2X1_46/Y gnd NAND3X1_6/C vdd NAND2X1
XNAND2X1_16 NOR2X1_64/A BUFX4_16/Y gnd OAI21X1_29/C vdd NAND2X1
XNAND2X1_180 XNOR2X1_28/Y INVX1_177/Y gnd AOI22X1_12/C vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XNAND2X1_191 NAND3X1_77/Y NAND2X1_191/B gnd OR2X2_15/B vdd NAND2X1
XFILL_17_1_0 gnd vdd FILL
XAOI22X1_47 INVX2_39/A INVX1_279/A INVX1_273/A AOI22X1_47/D gnd INVX2_43/A vdd AOI22X1
XAOI22X1_36 OR2X2_26/Y AOI22X1_36/B AOI22X1_36/C AOI22X1_36/D gnd NOR3X1_11/B vdd
+ AOI22X1
XAOI22X1_25 INVX1_205/Y INVX2_26/Y INVX1_212/Y AOI22X1_25/D gnd AOI22X1_25/Y vdd AOI22X1
XAOI22X1_14 AND2X2_25/A AND2X2_25/B NAND3X1_59/A NAND3X1_56/Y gnd AOI22X1_14/Y vdd
+ AOI22X1
XNOR3X1_4 INVX2_15/Y NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_4/Y vdd NOR3X1
XOAI22X1_9 INVX2_14/Y OAI22X1_9/B OAI22X1_9/C OAI22X1_9/D gnd OAI22X1_9/Y vdd OAI22X1
XAOI21X1_91 AOI21X1_91/A AOI21X1_91/B OAI22X1_18/Y gnd AOI21X1_91/Y vdd AOI21X1
XAOI21X1_80 AOI21X1_80/A AOI21X1_80/B INVX1_217/Y gnd AOI21X1_94/C vdd AOI21X1
XFILL_19_2 gnd vdd FILL
XINVX2_29 INVX2_29/A gnd INVX2_29/Y vdd INVX2
XINVX2_18 INVX2_18/A gnd INVX2_18/Y vdd INVX2
XXOR2X1_1 x1[1] x3[1] gnd XOR2X1_1/Y vdd XOR2X1
XFILL_6_0_0 gnd vdd FILL
XDFFPOSX1_109 BUFX2_5/A DFFSR_1/CLK NOR2X1_198/Y gnd vdd DFFPOSX1
XCLKBUF1_3 clk gnd CLKBUF1_3/Y vdd CLKBUF1
XNOR2X1_223 INVX1_304/Y AOI22X1_45/Y gnd NOR2X1_223/Y vdd NOR2X1
XNOR2X1_212 INVX1_286/A INVX1_287/A gnd INVX1_293/A vdd NOR2X1
XNOR2X1_201 NOR2X1_201/A NOR2X1_199/Y gnd NOR2X1_201/Y vdd NOR2X1
XDFFPOSX1_80 XOR2X1_5/B CLKBUF1_7/Y AND2X2_9/Y gnd vdd DFFPOSX1
XBUFX4_14 INVX8_1/Y gnd BUFX4_14/Y vdd BUFX4
XDFFPOSX1_91 INVX1_89/A CLKBUF1_2/Y OAI21X1_6/Y gnd vdd DFFPOSX1
XNAND3X1_341 INVX1_306/A AOI22X1_54/C OR2X2_34/A gnd OAI21X1_391/C vdd NAND3X1
XNAND3X1_330 OAI21X1_358/Y NAND3X1_334/A NAND3X1_334/C gnd NAND3X1_333/B vdd NAND3X1
XNAND3X1_363 OAI21X1_372/Y NAND3X1_360/B NAND3X1_360/C gnd NAND2X1_444/A vdd NAND3X1
XNAND3X1_352 NAND3X1_352/A NAND3X1_351/Y OAI21X1_383/Y gnd NAND2X1_436/B vdd NAND3X1
XOR2X2_28 OR2X2_28/A OR2X2_28/B gnd OR2X2_28/Y vdd OR2X2
XOR2X2_17 OR2X2_17/A OR2X2_17/B gnd OR2X2_17/Y vdd OR2X2
XFILL_21_2_1 gnd vdd FILL
XFILL_12_2_1 gnd vdd FILL
XNAND3X1_193 NAND3X1_194/B NAND3X1_194/C OAI21X1_297/Y gnd NAND2X1_312/B vdd NAND3X1
XNAND3X1_182 INVX1_235/A NAND3X1_182/B NAND3X1_182/C gnd AOI21X1_108/C vdd NAND3X1
XNAND3X1_160 OAI22X1_18/Y AOI21X1_90/Y AND2X2_31/Y gnd AND2X2_32/A vdd NAND3X1
XNAND3X1_171 AOI21X1_84/Y OAI22X1_19/Y NAND3X1_170/Y gnd NAND3X1_171/Y vdd NAND3X1
XOAI21X1_301 NOR3X1_8/Y INVX1_252/Y AND2X2_36/Y gnd NAND3X1_199/C vdd OAI21X1
XOAI21X1_323 OAI21X1_312/B NAND2X1_337/Y NAND3X1_228/A gnd NOR3X1_11/A vdd OAI21X1
XOAI21X1_312 OAI21X1_312/A OAI21X1_312/B OAI21X1_312/C gnd NAND3X1_232/B vdd OAI21X1
XOAI21X1_345 INVX1_282/A NAND2X1_380/A OR2X2_29/Y gnd OAI21X1_355/C vdd OAI21X1
XOAI21X1_356 INVX1_284/A NOR2X1_219/B AOI21X1_141/C gnd NAND3X1_286/A vdd OAI21X1
XOAI21X1_334 INVX1_273/A INVX2_38/A INVX2_40/A gnd AND2X2_43/B vdd OAI21X1
XOAI21X1_378 AOI22X1_51/Y XNOR2X1_49/A OAI21X1_377/Y gnd OAI21X1_378/Y vdd OAI21X1
XOAI21X1_367 INVX1_300/A INVX1_301/Y AND2X2_47/Y gnd NAND2X1_419/B vdd OAI21X1
XOAI21X1_389 OAI21X1_389/A INVX1_310/Y XNOR2X1_52/Y gnd NAND3X1_360/C vdd OAI21X1
XNAND2X1_384 OR2X2_30/B OR2X2_30/A gnd NAND3X1_277/B vdd NAND2X1
XNAND2X1_395 INVX1_288/Y NAND2X1_395/B gnd AOI22X1_46/D vdd NAND2X1
XNAND2X1_373 OAI21X1_342/Y NAND2X1_373/B gnd INVX1_280/A vdd NAND2X1
XNAND2X1_362 INVX1_273/A INVX2_35/Y gnd XNOR2X1_46/B vdd NAND2X1
XXOR2X1_23 XOR2X1_23/A XOR2X1_23/B gnd XOR2X1_23/Y vdd XOR2X1
XNAND2X1_340 OR2X2_26/B OR2X2_26/A gnd AOI22X1_36/B vdd NAND2X1
XNAND2X1_351 NAND2X1_351/A NAND2X1_351/B gnd NAND2X1_351/Y vdd NAND2X1
XXOR2X1_12 OR2X2_16/A OR2X2_16/B gnd XOR2X1_12/Y vdd XOR2X1
XFILL_7_2 gnd vdd FILL
XNAND3X1_2 x0[4] INVX1_44/Y INVX1_60/Y gnd NAND3X1_2/Y vdd NAND3X1
XFILL_1_1_1 gnd vdd FILL
XOAI21X1_120 AND2X2_13/Y OAI21X1_119/Y NAND2X1_84/Y gnd OAI21X1_120/Y vdd OAI21X1
XOAI21X1_164 INVX1_134/Y INVX1_136/A OAI21X1_167/C gnd OAI21X1_165/C vdd OAI21X1
XAOI22X1_7 AOI22X1_7/A AOI22X1_7/B AOI22X1_7/C AOI22X1_7/D gnd NOR3X1_2/C vdd AOI22X1
XOAI21X1_153 NOR2X1_97/B AOI21X1_33/Y AOI21X1_36/Y gnd AOI21X1_37/C vdd OAI21X1
XOAI21X1_131 INVX1_125/A AOI21X1_23/Y INVX1_126/A gnd NOR2X1_94/B vdd OAI21X1
XOAI21X1_142 BUFX4_4/Y INVX1_129/Y OAI21X1_88/C gnd DFFPOSX1_24/D vdd OAI21X1
XINVX1_217 INVX1_217/A gnd INVX1_217/Y vdd INVX1
XOAI21X1_186 NAND3X1_33/Y AOI22X1_6/Y NAND3X1_32/Y gnd AOI21X1_60/B vdd OAI21X1
XINVX1_239 INVX1_239/A gnd INVX1_239/Y vdd INVX1
XINVX1_228 gnd gnd INVX1_228/Y vdd INVX1
XOAI21X1_175 INVX1_158/A NOR2X1_113/Y INVX1_157/A gnd NAND3X1_22/A vdd OAI21X1
XFILL_9_2_1 gnd vdd FILL
XOAI21X1_197 INVX2_13/A INVX1_151/A INVX1_170/Y gnd XOR2X1_7/A vdd OAI21X1
XINVX1_206 OR2X2_16/Y gnd INVX1_206/Y vdd INVX1
XNAND2X1_28 BUFX4_3/Y OR2X2_2/A gnd OAI22X1_4/D vdd NAND2X1
XNAND2X1_39 INVX1_89/Y NOR2X1_55/Y gnd NOR2X1_56/B vdd NAND2X1
XNAND2X1_17 INVX1_109/A BUFX4_15/Y gnd NAND2X1_17/Y vdd NAND2X1
XNAND2X1_181 OR2X2_14/A XOR2X1_9/Y gnd AOI22X1_12/D vdd NAND2X1
XNAND2X1_192 INVX1_188/A AOI22X1_16/D gnd NAND3X1_78/C vdd NAND2X1
XNAND2X1_170 INVX2_10/A INVX2_16/A gnd XNOR2X1_25/A vdd NAND2X1
XFILL_17_1_1 gnd vdd FILL
XAOI22X1_48 AOI22X1_48/A AOI22X1_48/B AOI22X1_48/C AOI22X1_48/D gnd NOR3X1_12/B vdd
+ AOI22X1
XAOI22X1_37 AOI22X1_37/A AOI22X1_37/B AOI22X1_37/C AOI22X1_37/D gnd AOI22X1_37/Y vdd
+ AOI22X1
XAOI22X1_15 NAND3X1_66/Y AOI22X1_15/B NAND3X1_43/Y NAND3X1_71/B gnd AOI22X1_15/Y vdd
+ AOI22X1
XNOR3X1_5 NOR3X1_5/A NOR3X1_5/B NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XAOI22X1_26 AND2X2_27/Y AOI22X1_26/B XOR2X1_13/B XOR2X1_13/A gnd AOI22X1_26/Y vdd
+ AOI22X1
XAOI21X1_70 NAND3X1_80/C INVX1_198/A INVX1_186/Y gnd AOI21X1_70/Y vdd AOI21X1
XAOI21X1_81 AOI21X1_81/A AOI21X1_81/B INVX1_217/A gnd AOI21X1_81/Y vdd AOI21X1
XAOI21X1_92 AOI21X1_92/A AOI21X1_92/B AOI21X1_92/C gnd AOI21X1_92/Y vdd AOI21X1
XINVX2_19 INVX2_19/A gnd INVX2_19/Y vdd INVX2
XXOR2X1_2 XOR2X1_2/A XOR2X1_2/B gnd XOR2X1_2/Y vdd XOR2X1
XFILL_6_0_1 gnd vdd FILL
XCLKBUF1_4 clk gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_24_1 gnd vdd FILL
XNOR2X1_213 INVX1_286/Y INVX1_287/Y gnd NOR2X1_213/Y vdd NOR2X1
XNOR2X1_202 INVX2_36/A INVX2_37/Y gnd INVX2_38/A vdd NOR2X1
XNOR2X1_224 NOR2X1_224/A NOR2X1_224/B gnd NOR2X1_224/Y vdd NOR2X1
XDFFPOSX1_70 INVX1_113/A CLKBUF1_1/Y OAI21X1_65/Y gnd vdd DFFPOSX1
XDFFPOSX1_81 INVX1_63/A CLKBUF1_8/Y OAI21X1_49/Y gnd vdd DFFPOSX1
XBUFX4_15 INVX8_1/Y gnd BUFX4_15/Y vdd BUFX4
XDFFPOSX1_92 NOR2X1_56/A CLKBUF1_2/Y OAI21X1_7/Y gnd vdd DFFPOSX1
XNAND3X1_342 AOI21X1_146/Y NAND3X1_342/B NAND3X1_336/Y gnd NAND3X1_342/Y vdd NAND3X1
XNAND3X1_331 NAND2X1_423/Y NAND3X1_325/B NAND3X1_324/Y gnd NAND3X1_331/Y vdd NAND3X1
XNAND3X1_320 INVX1_302/Y NAND3X1_320/B NAND3X1_320/C gnd NAND3X1_327/C vdd NAND3X1
XNAND3X1_364 AOI21X1_163/Y NAND3X1_358/B NAND3X1_358/C gnd NAND3X1_364/Y vdd NAND3X1
XNAND3X1_353 OR2X2_33/Y NAND3X1_353/B NAND3X1_353/C gnd NAND3X1_353/Y vdd NAND3X1
XOR2X2_29 OR2X2_29/A OR2X2_29/B gnd OR2X2_29/Y vdd OR2X2
XOR2X2_18 OR2X2_18/A OR2X2_18/B gnd OR2X2_18/Y vdd OR2X2
XFILL_21_2_2 gnd vdd FILL
XFILL_12_2_2 gnd vdd FILL
XNAND3X1_150 INVX1_220/A AOI22X1_27/C OR2X2_20/A gnd OAI21X1_274/C vdd NAND3X1
XNAND3X1_194 NAND3X1_194/A NAND3X1_194/B NAND3X1_194/C gnd NAND3X1_196/A vdd NAND3X1
XNAND3X1_183 INVX1_235/Y NAND2X1_294/Y NAND2X1_295/Y gnd NAND2X1_313/B vdd NAND3X1
XNAND3X1_161 NAND3X1_111/Y NAND3X1_127/B NAND3X1_161/C gnd AOI21X1_93/A vdd NAND3X1
XNAND3X1_172 AOI21X1_99/C AOI21X1_99/B AOI21X1_99/A gnd NAND3X1_172/Y vdd NAND3X1
XOAI21X1_346 INVX1_273/A NOR2X1_209/Y INVX2_39/A gnd INVX1_285/A vdd OAI21X1
XOAI21X1_335 INVX1_273/Y INVX2_40/Y INVX1_274/Y gnd OAI21X1_335/Y vdd OAI21X1
XOAI21X1_324 INVX1_254/Y AOI21X1_109/Y NAND3X1_199/Y gnd XNOR2X1_45/B vdd OAI21X1
XOAI21X1_313 INVX1_247/A OAI21X1_313/B NAND3X1_230/C gnd OAI21X1_313/Y vdd OAI21X1
XOAI21X1_302 NOR3X1_8/A NOR3X1_8/C INVX1_253/Y gnd AOI22X1_34/C vdd OAI21X1
XOAI21X1_357 INVX1_286/A INVX1_287/A AOI22X1_46/B gnd NAND2X1_401/A vdd OAI21X1
XOAI21X1_379 NOR2X1_224/B INVX1_300/A INVX1_301/A gnd INVX1_307/A vdd OAI21X1
XOAI21X1_368 INVX1_300/A INVX1_301/Y NOR2X1_224/B gnd NAND2X1_420/B vdd OAI21X1
XNAND2X1_385 NAND3X1_277/B OR2X2_30/Y gnd OR2X2_31/A vdd NAND2X1
XNAND2X1_396 NAND3X1_283/Y NAND3X1_286/Y gnd XOR2X1_21/A vdd NAND2X1
XNAND2X1_374 NOR2X1_211/A INVX1_280/Y gnd NAND2X1_374/Y vdd NAND2X1
XNAND2X1_363 NOR2X1_211/A OAI21X1_335/Y gnd OR2X2_28/B vdd NAND2X1
XXOR2X1_13 XOR2X1_13/A XOR2X1_13/B gnd XOR2X1_13/Y vdd XOR2X1
XXOR2X1_24 XOR2X1_24/A OR2X2_33/B gnd XOR2X1_24/Y vdd XOR2X1
XNAND2X1_352 NAND2X1_351/Y OAI21X1_321/Y gnd NAND2X1_352/Y vdd NAND2X1
XNAND2X1_330 AND2X2_37/Y AND2X2_38/Y gnd OAI21X1_320/C vdd NAND2X1
XNAND2X1_341 INVX2_28/A INVX1_132/A gnd OR2X2_27/B vdd NAND2X1
XFILL_7_3 gnd vdd FILL
XNAND3X1_3 x1[0] x3[0] XOR2X1_1/Y gnd NAND3X1_4/B vdd NAND3X1
XFILL_1_1_2 gnd vdd FILL
XOAI21X1_143 OAI21X1_143/A XNOR2X1_11/Y NAND2X1_103/Y gnd AOI21X1_29/A vdd OAI21X1
XOAI21X1_110 INVX1_114/Y INVX1_113/A NAND2X1_69/Y gnd OAI21X1_111/C vdd OAI21X1
XOAI21X1_165 INVX1_136/A INVX1_143/A OAI21X1_165/C gnd INVX1_138/A vdd OAI21X1
XAOI22X1_8 AOI22X1_8/A AOI22X1_8/B AOI22X1_8/C AOI22X1_8/D gnd NOR3X1_2/B vdd AOI22X1
XOAI21X1_198 INVX1_171/A INVX1_169/Y XOR2X1_7/Y gnd INVX1_178/A vdd OAI21X1
XINVX1_207 INVX1_207/A gnd INVX1_207/Y vdd INVX1
XOAI21X1_154 AND2X2_16/B AND2X2_16/A BUFX4_5/Y gnd OAI21X1_155/B vdd OAI21X1
XOAI21X1_176 gnd NOR2X1_110/Y gnd gnd INVX1_156/A vdd OAI21X1
XOAI21X1_187 INVX1_145/A INVX1_146/A INVX2_14/A gnd NAND2X1_152/A vdd OAI21X1
XOAI21X1_121 NAND2X1_85/Y INVX2_5/A NAND2X1_87/Y gnd AOI21X1_22/A vdd OAI21X1
XOAI21X1_132 INVX2_7/Y AOI21X1_26/Y BUFX4_7/Y gnd OAI21X1_132/Y vdd OAI21X1
XINVX1_229 INVX1_229/A gnd INVX1_229/Y vdd INVX1
XINVX1_218 INVX1_218/A gnd INVX1_218/Y vdd INVX1
XFILL_9_2_2 gnd vdd FILL
XNAND2X1_29 x0[7] x2[7] gnd INVX1_51/A vdd NAND2X1
XNAND2X1_18 AND2X2_2/B AOI21X1_4/B gnd NAND2X1_18/Y vdd NAND2X1
XFILL_17_1_2 gnd vdd FILL
XNAND2X1_193 NAND3X1_78/A NAND3X1_78/C gnd OAI21X1_222/C vdd NAND2X1
XNAND2X1_160 INVX1_164/A NOR2X1_119/Y gnd AOI22X1_8/D vdd NAND2X1
XNAND2X1_182 XOR2X1_9/A OR2X2_14/A gnd NAND3X1_55/A vdd NAND2X1
XNAND2X1_171 INVX2_9/A INVX1_127/A gnd XNOR2X1_25/B vdd NAND2X1
XAOI22X1_49 AOI22X1_49/A AOI22X1_49/B AOI22X1_49/C AOI22X1_49/D gnd NOR3X1_12/C vdd
+ AOI22X1
XAOI22X1_38 AOI22X1_38/A AOI22X1_38/B AOI22X1_41/C AOI22X1_41/D gnd AOI22X1_38/Y vdd
+ AOI22X1
XNOR3X1_6 NOR3X1_6/A NOR3X1_6/B NOR3X1_6/C gnd NOR3X1_6/Y vdd NOR3X1
XAOI22X1_27 AOI21X1_76/C AOI22X1_26/B AOI22X1_27/C OR2X2_20/A gnd AOI22X1_27/Y vdd
+ AOI22X1
XAOI22X1_16 INVX2_18/A NOR2X1_140/B INVX1_188/A AOI22X1_16/D gnd OR2X2_16/B vdd AOI22X1
XAOI21X1_93 AOI21X1_93/A AOI21X1_93/B AOI21X1_93/C gnd AOI21X1_93/Y vdd AOI21X1
XAOI21X1_60 NAND3X1_54/Y AOI21X1_60/B AOI21X1_60/C gnd NAND3X1_73/C vdd AOI21X1
XAOI21X1_82 INVX1_195/A NAND3X1_93/C INVX1_219/Y gnd AOI21X1_82/Y vdd AOI21X1
XAOI21X1_71 NAND3X1_84/C NAND3X1_84/B INVX1_197/Y gnd AOI21X1_76/C vdd AOI21X1
XFILL_6_0_2 gnd vdd FILL
XXOR2X1_3 XOR2X1_3/A NOR2X1_9/Y gnd XOR2X1_3/Y vdd XOR2X1
XCLKBUF1_5 clk gnd CLKBUF1_5/Y vdd CLKBUF1
XFILL_24_2 gnd vdd FILL
XNOR2X1_214 INVX1_293/A NOR2X1_213/Y gnd OR2X2_30/A vdd NOR2X1
XNOR2X1_203 INVX2_35/Y INVX2_39/Y gnd INVX2_40/A vdd NOR2X1
XFILL_17_1 gnd vdd FILL
XNOR2X1_225 NOR2X1_225/A XNOR2X1_51/Y gnd NOR2X1_225/Y vdd NOR2X1
XDFFPOSX1_71 INVX1_78/A CLKBUF1_1/Y OAI21X1_70/Y gnd vdd DFFPOSX1
XDFFPOSX1_93 INVX1_12/A CLKBUF1_1/Y OAI22X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_82 INVX1_65/A CLKBUF1_9/Y OAI21X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_60 INVX1_56/A CLKBUF1_9/Y NOR2X1_36/Y gnd vdd DFFPOSX1
XBUFX4_16 INVX8_1/Y gnd BUFX4_16/Y vdd BUFX4
XNAND3X1_332 NOR2X1_223/Y NAND3X1_331/Y NAND3X1_335/C gnd NAND3X1_333/C vdd NAND3X1
XNAND3X1_321 INVX1_303/A NAND3X1_327/B NAND3X1_327/C gnd NAND3X1_325/B vdd NAND3X1
XFILL_15_2_0 gnd vdd FILL
XNAND3X1_310 OAI22X1_21/Y NAND3X1_304/Y NAND3X1_310/C gnd NAND3X1_315/B vdd NAND3X1
XNAND3X1_343 NAND2X1_400/Y NAND3X1_343/B NAND3X1_343/C gnd NAND3X1_343/Y vdd NAND3X1
XNAND3X1_365 OAI21X1_390/Y OR2X2_34/Y NAND2X1_444/Y gnd NAND3X1_365/Y vdd NAND3X1
XNAND3X1_354 NAND2X1_436/A NAND2X1_436/B XOR2X1_24/Y gnd NAND3X1_354/Y vdd NAND3X1
XOR2X2_19 OR2X2_19/A OR2X2_19/B gnd OR2X2_19/Y vdd OR2X2
XNAND3X1_162 AOI21X1_93/A AOI21X1_93/B AOI21X1_93/C gnd NAND3X1_162/Y vdd NAND3X1
XNAND3X1_184 INVX1_230/A AOI21X1_108/C NAND2X1_313/B gnd NAND3X1_184/Y vdd NAND3X1
XNAND3X1_140 NAND2X1_251/Y NAND3X1_130/Y AOI21X1_94/A gnd AOI21X1_96/B vdd NAND3X1
XNAND3X1_173 AOI21X1_97/Y AOI21X1_98/B AOI21X1_98/A gnd NAND3X1_173/Y vdd NAND3X1
XNAND3X1_151 AOI21X1_82/Y NAND3X1_146/B NAND3X1_146/C gnd AOI21X1_83/B vdd NAND3X1
XNAND3X1_195 NAND3X1_190/B NAND3X1_189/Y OAI21X1_297/Y gnd NAND3X1_195/Y vdd NAND3X1
XOAI21X1_358 OAI21X1_358/A NAND2X1_403/Y INVX1_304/A gnd OAI21X1_358/Y vdd OAI21X1
XOAI21X1_347 INVX2_41/A INVX1_279/A INVX1_273/A gnd OAI21X1_347/Y vdd OAI21X1
XFILL_21_0_0 gnd vdd FILL
XOAI21X1_336 INVX2_37/A INVX1_95/A INVX2_36/A gnd NOR2X1_207/A vdd OAI21X1
XOAI21X1_369 INVX2_36/Y INVX1_299/Y OAI21X1_362/C gnd AND2X2_48/B vdd OAI21X1
XOAI21X1_314 NOR3X1_8/A NOR3X1_8/B OR2X2_25/Y gnd XNOR2X1_42/A vdd OAI21X1
XOAI21X1_303 AOI21X1_109/Y NOR3X1_9/Y INVX1_254/A gnd NAND2X1_326/B vdd OAI21X1
XOAI21X1_325 NOR3X1_10/Y AOI21X1_128/Y XNOR2X1_45/Y gnd NAND3X1_257/B vdd OAI21X1
XXOR2X1_25 XOR2X1_25/A XOR2X1_25/B gnd XOR2X1_25/Y vdd XOR2X1
XBUFX4_1 start gnd BUFX4_1/Y vdd BUFX4
XXOR2X1_14 XOR2X1_14/A XOR2X1_14/B gnd XOR2X1_14/Y vdd XOR2X1
XNAND2X1_320 gnd gnd gnd OR2X2_25/B vdd NAND2X1
XNAND2X1_386 INVX1_285/A OR2X2_31/A gnd AOI22X1_46/A vdd NAND2X1
XNAND2X1_397 NAND3X1_287/B NAND3X1_287/C gnd AOI22X1_53/B vdd NAND2X1
XNAND2X1_375 NAND2X1_374/Y INVX1_281/Y gnd INVX1_282/A vdd NAND2X1
XNAND2X1_364 INVX1_274/A AOI22X1_42/D gnd NAND2X1_364/Y vdd NAND2X1
XNAND2X1_353 NAND2X1_348/Y OAI21X1_321/Y gnd NAND2X1_353/Y vdd NAND2X1
XFILL_4_1_0 gnd vdd FILL
XNAND2X1_331 INVX2_29/A AND2X2_38/B gnd NOR2X1_195/B vdd NAND2X1
XNAND2X1_342 INVX2_29/A OR2X2_6/B gnd OR2X2_27/A vdd NAND2X1
XFILL_12_0_0 gnd vdd FILL
XNAND3X1_4 BUFX4_2/Y NAND3X1_4/B NAND3X1_4/C gnd NAND3X1_4/Y vdd NAND3X1
XOAI21X1_144 NAND2X1_65/A NOR2X1_95/A OAI21X1_144/C gnd AOI21X1_29/C vdd OAI21X1
XOAI21X1_111 INVX1_114/A INVX1_113/Y OAI21X1_111/C gnd OAI21X1_111/Y vdd OAI21X1
XOAI21X1_199 INVX2_9/Y INVX2_16/Y INVX1_163/A gnd NAND2X1_165/A vdd OAI21X1
XAOI22X1_9 INVX1_168/Y INVX1_146/Y AOI22X1_9/C INVX1_167/Y gnd NOR3X1_3/C vdd AOI22X1
XINVX1_208 INVX1_208/A gnd OR2X2_20/B vdd INVX1
XOAI21X1_122 NOR2X1_85/A AND2X2_14/A BUFX4_5/Y gnd OAI21X1_122/Y vdd OAI21X1
XOAI21X1_155 AND2X2_16/Y OAI21X1_155/B NAND2X1_112/Y gnd DFFPOSX1_5/D vdd OAI21X1
XOAI21X1_166 INVX2_10/A INVX1_139/A INVX2_9/A gnd NOR2X1_107/A vdd OAI21X1
XOAI21X1_188 INVX2_12/Y INVX1_145/A NAND3X1_21/C gnd INVX2_15/A vdd OAI21X1
XINVX1_219 INVX1_219/A gnd INVX1_219/Y vdd INVX1
XOAI21X1_100 BUFX4_9/Y INVX1_102/Y NAND2X1_55/Y gnd DFFPOSX1_10/D vdd OAI21X1
XOAI21X1_133 NOR2X1_94/Y OAI21X1_132/Y NAND2X1_91/Y gnd DFFPOSX1_31/D vdd OAI21X1
XOAI21X1_177 gnd gnd gnd gnd INVX1_147/A vdd OAI21X1
XNAND2X1_19 INVX1_38/Y INVX1_39/Y gnd NAND2X1_21/B vdd NAND2X1
XNAND2X1_150 NAND3X1_22/Y NAND3X1_28/Y gnd INVX1_175/A vdd NAND2X1
XNAND2X1_161 INVX2_9/A INVX2_13/Y gnd INVX1_168/A vdd NAND2X1
XNAND2X1_194 NAND3X1_78/Y OAI21X1_222/Y gnd OR2X2_15/A vdd NAND2X1
XNAND2X1_172 gnd gnd gnd XOR2X1_10/B vdd NAND2X1
XNAND2X1_183 NAND3X1_55/A OR2X2_14/Y gnd NAND2X1_183/Y vdd NAND2X1
XAOI22X1_39 NOR2X1_187/Y AOI22X1_39/B XOR2X1_18/B XOR2X1_18/A gnd AOI22X1_39/Y vdd
+ AOI22X1
XAOI22X1_28 INVX2_28/A AOI22X1_28/B INVX1_229/A NOR2X1_172/Y gnd OR2X2_22/B vdd AOI22X1
XAOI22X1_17 AOI22X1_20/A NAND3X1_86/Y AOI22X1_17/C AOI22X1_17/D gnd AOI22X1_17/Y vdd
+ AOI22X1
XNOR3X1_7 NOR3X1_7/A NOR3X1_7/B NOR3X1_7/C gnd NOR3X1_7/Y vdd NOR3X1
XXNOR2X1_50 XNOR2X1_50/A XNOR2X1_50/B gnd XNOR2X1_50/Y vdd XNOR2X1
XFILL_5_1 gnd vdd FILL
XOAI21X1_1 NOR2X1_1/Y NOR2X1_2/Y BUFX4_2/Y gnd OAI21X1_1/Y vdd OAI21X1
XAOI21X1_94 AOI21X1_94/A AOI21X1_94/B AOI21X1_94/C gnd AOI21X1_94/Y vdd AOI21X1
XAOI21X1_50 INVX1_158/Y OR2X2_12/Y INVX1_157/Y gnd NAND3X1_25/A vdd AOI21X1
XAOI21X1_61 NOR2X1_121/B AOI21X1_61/B INVX1_171/A gnd OR2X2_14/A vdd AOI21X1
XAOI21X1_83 AOI21X1_83/A AOI21X1_83/B INVX1_220/Y gnd AOI21X1_84/C vdd AOI21X1
XAOI21X1_72 AOI21X1_72/A AOI21X1_72/B INVX1_197/A gnd AOI21X1_72/Y vdd AOI21X1
XFILL_9_0_0 gnd vdd FILL
XXOR2X1_4 INVX1_47/A INVX1_78/A gnd XOR2X1_4/Y vdd XOR2X1
XCLKBUF1_6 clk gnd CLKBUF1_6/Y vdd CLKBUF1
XNOR2X1_204 INVX2_35/Y INVX2_41/Y gnd INVX1_274/A vdd NOR2X1
XNOR2X1_215 INVX1_278/A NOR2X1_215/B gnd NOR2X1_215/Y vdd NOR2X1
XFILL_24_3 gnd vdd FILL
XFILL_17_2 gnd vdd FILL
XNOR2X1_226 OR2X2_34/B OR2X2_34/A gnd OAI22X1_22/D vdd NOR2X1
XDFFPOSX1_50 NOR2X1_64/A CLKBUF1_2/Y OAI21X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_72 INVX1_80/A CLKBUF1_1/Y OAI22X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_94 OR2X2_3/B CLKBUF1_1/Y OAI21X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_83 INVX1_66/A CLKBUF1_8/Y OAI21X1_51/Y gnd vdd DFFPOSX1
XDFFPOSX1_61 INVX1_57/A CLKBUF1_3/Y NOR2X1_37/Y gnd vdd DFFPOSX1
XBUFX4_17 INVX8_1/Y gnd OR2X2_4/B vdd BUFX4
XNAND3X1_344 INVX1_306/Y NAND3X1_342/Y NAND3X1_343/Y gnd NAND2X1_424/B vdd NAND3X1
XNAND3X1_333 INVX1_295/Y NAND3X1_333/B NAND3X1_333/C gnd NAND3X1_342/B vdd NAND3X1
XNAND3X1_366 NAND3X1_366/A OAI21X1_392/Y NAND3X1_365/Y gnd NAND2X1_445/B vdd NAND3X1
XNAND3X1_322 INVX1_302/Y NAND3X1_317/B NAND3X1_317/C gnd NAND3X1_324/B vdd NAND3X1
XNAND3X1_300 INVX2_37/A INVX1_98/A NOR2X1_224/A gnd NAND3X1_301/C vdd NAND3X1
XNAND3X1_311 AND2X2_47/Y INVX1_301/A INVX1_300/Y gnd NAND2X1_420/A vdd NAND3X1
XFILL_15_2_1 gnd vdd FILL
XNAND3X1_355 INVX1_308/Y NAND3X1_354/Y NAND3X1_353/Y gnd NAND3X1_356/A vdd NAND3X1
XNAND3X1_130 INVX1_217/A AOI21X1_81/A AOI21X1_81/B gnd NAND3X1_130/Y vdd NAND3X1
XNAND3X1_163 AOI21X1_92/A AOI21X1_92/B AOI21X1_92/C gnd NAND3X1_164/B vdd NAND3X1
XNAND3X1_196 NAND3X1_196/A NAND3X1_195/Y XOR2X1_18/B gnd NAND3X1_196/Y vdd NAND3X1
XNAND3X1_185 OAI21X1_290/Y OAI21X1_291/Y NOR2X1_184/Y gnd NAND2X1_307/B vdd NAND3X1
XNAND3X1_141 NOR2X1_156/Y AOI21X1_96/B AOI21X1_96/A gnd AOI21X1_97/B vdd NAND3X1
XNAND3X1_152 NAND2X1_228/Y NAND3X1_149/B NAND3X1_149/C gnd AOI21X1_83/A vdd NAND3X1
XNAND3X1_174 OAI21X1_273/Y OR2X2_20/Y NAND2X1_275/Y gnd NAND3X1_174/Y vdd NAND3X1
XOAI21X1_359 INVX2_41/Y INVX1_286/A NAND3X1_277/B gnd INVX1_297/A vdd OAI21X1
XFILL_21_0_1 gnd vdd FILL
XOAI21X1_348 INVX1_278/A NOR2X1_215/B INVX1_287/A gnd INVX1_289/A vdd OAI21X1
XOAI21X1_337 NOR2X1_207/A NOR2X1_206/Y INVX1_274/Y gnd NAND3X1_269/A vdd OAI21X1
XOAI21X1_315 INVX2_32/Y NOR3X1_8/A OR2X2_25/Y gnd XOR2X1_19/B vdd OAI21X1
XOAI21X1_326 NOR3X1_8/C NOR3X1_8/Y XNOR2X1_45/B gnd OAI21X1_326/Y vdd OAI21X1
XOAI21X1_304 NOR3X1_9/B NOR3X1_9/C INVX2_34/A gnd OAI21X1_304/Y vdd OAI21X1
XBUFX4_2 start gnd BUFX4_2/Y vdd BUFX4
XNAND2X1_321 gnd gnd gnd NOR3X1_8/B vdd NAND2X1
XNAND2X1_354 AOI22X1_36/B OR2X2_26/Y gnd INVX1_271/A vdd NAND2X1
XNAND2X1_310 INVX1_236/A INVX1_239/Y gnd AOI22X1_31/D vdd NAND2X1
XNAND2X1_332 NOR2X1_195/B AND2X2_37/Y gnd NAND2X1_332/Y vdd NAND2X1
XXOR2X1_15 XOR2X1_15/A XOR2X1_15/B gnd XOR2X1_15/Y vdd XOR2X1
XNAND2X1_343 AND2X2_40/B OR2X2_27/Y gnd NAND2X1_343/Y vdd NAND2X1
XNAND2X1_376 XOR2X1_20/Y INVX1_282/Y gnd NAND2X1_376/Y vdd NAND2X1
XNAND2X1_387 NAND2X1_387/A NAND2X1_372/A gnd INVX1_288/A vdd NAND2X1
XNAND2X1_365 NAND3X1_269/A NAND2X1_364/Y gnd NAND2X1_365/Y vdd NAND2X1
XNAND2X1_398 AOI22X1_53/B AND2X2_44/Y gnd NAND2X1_398/Y vdd NAND2X1
XFILL_4_1_1 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XNAND3X1_5 INVX1_8/A XOR2X1_2/B AOI21X1_9/A gnd AND2X2_8/A vdd NAND3X1
XOAI21X1_112 NAND2X1_69/Y NAND3X1_12/B NAND2X1_80/Y gnd AOI21X1_18/A vdd OAI21X1
XOAI21X1_101 BUFX4_4/Y INVX1_103/Y OAI21X1_93/C gnd DFFPOSX1_11/D vdd OAI21X1
XOAI21X1_145 OAI21X1_145/A NAND3X1_8/B NAND2X1_106/Y gnd AOI21X1_31/A vdd OAI21X1
XOAI21X1_134 INVX2_7/Y AOI21X1_26/Y INVX1_124/Y gnd NAND2X1_94/B vdd OAI21X1
XOAI21X1_189 INVX1_180/A AND2X2_22/Y INVX1_163/Y gnd AOI22X1_7/B vdd OAI21X1
XINVX1_209 INVX1_209/A gnd INVX1_209/Y vdd INVX1
XOAI21X1_167 NOR2X1_107/A INVX1_141/A OAI21X1_167/C gnd NAND2X1_122/A vdd OAI21X1
XOAI21X1_123 AND2X2_14/Y OAI21X1_122/Y NAND2X1_86/Y gnd OAI21X1_123/Y vdd OAI21X1
XOAI21X1_156 AND2X2_16/B AND2X2_16/A NOR2X1_98/A gnd XNOR2X1_17/A vdd OAI21X1
XOAI21X1_178 INVX2_12/Y INVX1_145/A INVX1_147/Y gnd INVX1_148/A vdd OAI21X1
XNAND2X1_195 OR2X2_15/B OR2X2_15/A gnd NAND3X1_79/B vdd NAND2X1
XNAND2X1_173 XOR2X1_10/A XOR2X1_8/Y gnd AOI22X1_11/A vdd NAND2X1
XNAND2X1_184 NAND2X1_183/Y INVX1_179/Y gnd NAND3X1_56/C vdd NAND2X1
XNAND2X1_140 NAND2X1_140/A NOR3X1_2/A gnd INVX1_154/A vdd NAND2X1
XNAND2X1_151 NAND3X1_68/A INVX2_14/Y gnd XNOR2X1_30/B vdd NAND2X1
XNAND2X1_162 INVX2_9/A NAND2X1_90/A gnd XOR2X1_7/B vdd NAND2X1
XAOI22X1_29 AOI22X1_31/B AOI22X1_31/A AOI22X1_29/C AOI22X1_32/D gnd AOI22X1_29/Y vdd
+ AOI22X1
XAOI22X1_18 AOI22X1_18/A INVX1_218/A AOI22X1_19/C OR2X2_18/Y gnd AOI22X1_18/Y vdd
+ AOI22X1
XNOR3X1_8 NOR3X1_8/A NOR3X1_8/B NOR3X1_8/C gnd NOR3X1_8/Y vdd NOR3X1
XXNOR2X1_51 XOR2X1_23/A XOR2X1_23/B gnd XNOR2X1_51/Y vdd XNOR2X1
XXNOR2X1_40 XNOR2X1_39/A INVX1_256/A gnd XNOR2X1_40/Y vdd XNOR2X1
XFILL_5_2 gnd vdd FILL
XOAI21X1_2 INVX1_1/Y BUFX4_2/Y OAI21X1_1/Y gnd OAI21X1_2/Y vdd OAI21X1
XAOI21X1_73 AOI21X1_73/A NAND3X1_85/Y INVX1_191/A gnd XOR2X1_13/B vdd AOI21X1
XAOI21X1_95 AOI21X1_95/A AOI21X1_95/B XOR2X1_14/Y gnd AOI21X1_95/Y vdd AOI21X1
XAOI21X1_51 NAND3X1_24/Y NAND3X1_27/Y INVX2_11/A gnd NOR3X1_6/B vdd AOI21X1
XAOI21X1_62 AND2X2_23/Y NAND3X1_36/C INVX1_178/Y gnd AOI21X1_62/Y vdd AOI21X1
XFILL_9_0_1 gnd vdd FILL
XAOI21X1_84 AOI21X1_84/A AOI21X1_84/B AOI21X1_84/C gnd AOI21X1_84/Y vdd AOI21X1
XAOI21X1_40 AOI21X1_40/A XOR2X1_5/Y BUFX4_10/Y gnd AOI22X1_5/D vdd AOI21X1
XXOR2X1_5 XOR2X1_5/A XOR2X1_5/B gnd XOR2X1_5/Y vdd XOR2X1
XCLKBUF1_7 clk gnd CLKBUF1_7/Y vdd CLKBUF1
XNOR2X1_216 INVX1_289/Y INVX2_42/Y gnd NOR2X1_216/Y vdd NOR2X1
XNOR2X1_205 INVX2_38/Y INVX2_40/Y gnd NOR2X1_205/Y vdd NOR2X1
XNOR2X1_227 INVX1_277/Y NOR2X1_227/B gnd NOR2X1_227/Y vdd NOR2X1
XFILL_17_3 gnd vdd FILL
XDFFPOSX1_95 INVX1_20/A CLKBUF1_7/Y OAI22X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_51 INVX1_109/A CLKBUF1_2/Y OAI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_40 INVX1_100/A CLKBUF1_4/Y OAI21X1_98/Y gnd vdd DFFPOSX1
XDFFPOSX1_84 INVX1_67/A CLKBUF1_8/Y OAI21X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_73 INVX1_82/A CLKBUF1_8/Y AOI21X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_62 INVX1_58/A CLKBUF1_3/Y NOR2X1_38/Y gnd vdd DFFPOSX1
XNAND3X1_334 NAND3X1_334/A NOR2X1_223/Y NAND3X1_334/C gnd NAND3X1_334/Y vdd NAND3X1
XNAND3X1_345 OAI22X1_21/Y AOI21X1_154/Y AND2X2_48/Y gnd NAND2X1_431/B vdd NAND3X1
XNAND3X1_323 INVX1_302/A NAND3X1_320/B NAND3X1_320/C gnd NAND3X1_324/C vdd NAND3X1
XNAND3X1_301 INVX2_44/A NAND3X1_301/B NAND3X1_301/C gnd AOI21X1_152/B vdd NAND3X1
XFILL_15_2_2 gnd vdd FILL
XNAND3X1_312 OAI21X1_375/A NAND3X1_315/B NAND3X1_309/Y gnd NAND3X1_318/C vdd NAND3X1
XNAND3X1_356 NAND3X1_356/A INVX1_309/A NAND3X1_356/C gnd INVX1_310/A vdd NAND3X1
XAOI21X1_160 NAND3X1_324/Y NAND2X1_410/Y OAI21X1_371/A gnd XNOR2X1_52/A vdd AOI21X1
XNAND3X1_120 AND2X2_30/Y INVX1_215/A INVX1_214/Y gnd NAND2X1_248/A vdd NAND3X1
XNAND3X1_131 INVX1_216/Y NAND3X1_122/Y AOI21X1_87/A gnd AOI21X1_80/A vdd NAND3X1
XNAND3X1_164 INVX1_222/Y NAND3X1_164/B NAND3X1_162/Y gnd AOI21X1_95/B vdd NAND3X1
XNAND3X1_197 INVX1_251/Y INVX1_250/A OR2X2_25/Y gnd AND2X2_36/A vdd NAND3X1
XNAND3X1_186 INVX1_240/Y NAND2X1_307/A NAND2X1_307/B gnd AOI22X1_31/B vdd NAND3X1
XNAND3X1_142 INVX1_209/Y NAND3X1_142/B AOI21X1_97/B gnd NAND3X1_146/B vdd NAND3X1
XNAND3X1_153 INVX1_220/Y AOI21X1_83/B AOI21X1_83/A gnd AOI21X1_84/A vdd NAND3X1
XNAND3X1_175 NAND3X1_175/A OAI21X1_275/Y NAND3X1_174/Y gnd NAND3X1_175/Y vdd NAND3X1
XFILL_21_0_2 gnd vdd FILL
XOAI21X1_305 INVX1_243/A INVX1_257/A INVX1_255/Y gnd XNOR2X1_39/A vdd OAI21X1
XBUFX4_3 start gnd BUFX4_3/Y vdd BUFX4
XOAI21X1_338 INVX2_38/Y INVX2_40/Y NAND2X1_365/Y gnd OAI21X1_338/Y vdd OAI21X1
XOAI21X1_349 INVX1_290/Y NOR2X1_218/B NOR2X1_206/Y gnd NAND2X1_391/A vdd OAI21X1
XOAI21X1_316 INVX1_262/A OAI21X1_316/B NAND3X1_213/Y gnd OAI21X1_316/Y vdd OAI21X1
XOAI21X1_327 AOI21X1_132/Y NOR3X1_11/Y AND2X2_42/Y gnd NAND3X1_262/C vdd OAI21X1
XNAND2X1_377 OR2X2_29/B OR2X2_29/A gnd AOI21X1_139/B vdd NAND2X1
XNAND2X1_366 OAI21X1_339/C OAI21X1_338/Y gnd OR2X2_28/A vdd NAND2X1
XNAND2X1_355 OAI21X1_326/Y NAND3X1_258/Y gnd NAND2X1_356/B vdd NAND2X1
XNAND2X1_311 INVX1_240/Y NAND2X1_307/Y gnd AOI22X1_30/A vdd NAND2X1
XNAND2X1_300 INVX1_236/Y INVX1_239/Y gnd AOI22X1_32/D vdd NAND2X1
XNAND2X1_322 gnd INVX1_228/Y gnd INVX1_250/A vdd NAND2X1
XNAND2X1_333 AND2X2_39/B AND2X2_39/A gnd NAND2X1_333/Y vdd NAND2X1
XNAND2X1_344 OAI21X1_317/Y AND2X2_40/Y gnd NAND3X1_242/C vdd NAND2X1
XXOR2X1_16 XOR2X1_16/A XOR2X1_16/B gnd XOR2X1_16/Y vdd XOR2X1
XNAND2X1_399 NAND2X1_398/Y NAND3X1_289/Y gnd XNOR2X1_50/B vdd NAND2X1
XNAND2X1_388 INVX2_37/A INVX1_97/A gnd NOR2X1_215/B vdd NAND2X1
XFILL_4_1_2 gnd vdd FILL
XFILL_12_0_2 gnd vdd FILL
XNAND3X1_6 BUFX4_3/Y NAND3X1_6/B NAND3X1_6/C gnd NAND3X1_6/Y vdd NAND3X1
XOAI21X1_113 INVX1_116/Y INVX1_80/A NAND3X1_9/Y gnd INVX1_118/A vdd OAI21X1
XOAI21X1_146 NAND2X1_74/Y AND2X2_12/Y OAI21X1_146/C gnd AOI21X1_31/C vdd OAI21X1
XOAI21X1_135 BUFX4_13/Y INVX1_24/Y NAND2X1_95/Y gnd DFFPOSX1_17/D vdd OAI21X1
XOAI21X1_124 NOR2X1_80/Y NOR2X1_79/Y OR2X2_5/B gnd AOI22X1_2/C vdd OAI21X1
XOAI21X1_102 BUFX4_4/Y INVX1_104/Y NAND2X1_57/Y gnd DFFPOSX1_12/D vdd OAI21X1
XOAI21X1_168 OR2X2_8/B OR2X2_8/A NAND3X1_14/Y gnd OR2X2_11/B vdd OAI21X1
XOAI21X1_157 BUFX4_11/Y XNOR2X1_17/Y NAND2X1_114/Y gnd DFFPOSX1_6/D vdd OAI21X1
XOAI21X1_179 NAND3X1_68/A NOR2X1_115/Y INVX1_148/A gnd NAND3X1_21/B vdd OAI21X1
XNAND2X1_196 NAND3X1_79/B OR2X2_15/Y gnd NAND2X1_197/B vdd NAND2X1
XNAND2X1_185 AND2X2_25/A AND2X2_25/B gnd AOI21X1_63/C vdd NAND2X1
XNAND2X1_174 INVX1_176/Y XNOR2X1_27/Y gnd AOI22X1_11/B vdd NAND2X1
XNAND2X1_163 INVX1_172/A NOR2X1_121/B gnd INVX1_169/A vdd NAND2X1
XNAND2X1_130 NOR2X1_110/Y XOR2X1_6/Y gnd AND2X2_20/B vdd NAND2X1
XNAND2X1_152 NAND2X1_152/A XNOR2X1_30/B gnd INVX1_161/A vdd NAND2X1
XNAND2X1_141 INVX2_10/A INVX1_153/A gnd INVX1_151/A vdd NAND2X1
XNOR3X1_9 INVX2_34/A NOR3X1_9/B NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XAOI22X1_19 AOI22X1_17/D AOI22X1_17/C AOI22X1_19/C OR2X2_18/Y gnd NOR2X1_156/B vdd
+ AOI22X1
XXNOR2X1_30 NAND3X1_48/B XNOR2X1_30/B gnd NAND3X1_71/B vdd XNOR2X1
XXNOR2X1_41 XNOR2X1_41/A XNOR2X1_41/B gnd XNOR2X1_41/Y vdd XNOR2X1
XXNOR2X1_52 XNOR2X1_52/A INVX1_311/A gnd XNOR2X1_52/Y vdd XNOR2X1
XAOI21X1_30 AND2X2_12/A NAND3X1_9/C NAND2X1_75/Y gnd AOI21X1_30/Y vdd AOI21X1
XAOI21X1_41 INVX1_136/A AOI21X1_41/B AOI21X1_41/C gnd INVX1_137/A vdd AOI21X1
XAOI21X1_52 NAND3X1_28/Y NAND3X1_29/Y INVX2_11/Y gnd NOR3X1_6/C vdd AOI21X1
XOAI21X1_3 x1[0] INVX1_2/Y XNOR2X1_1/Y gnd OAI21X1_5/C vdd OAI21X1
XAOI21X1_85 AOI21X1_85/A AOI21X1_85/B AOI21X1_85/C gnd AOI21X1_85/Y vdd AOI21X1
XAOI21X1_63 NAND3X1_60/Y NAND3X1_61/A AOI21X1_63/C gnd AOI21X1_63/Y vdd AOI21X1
XAOI21X1_96 AOI21X1_96/A AOI21X1_96/B NOR2X1_156/Y gnd AOI21X1_96/Y vdd AOI21X1
XFILL_9_0_2 gnd vdd FILL
XAOI21X1_74 INVX1_200/Y INVX2_23/A AOI21X1_74/C gnd OR2X2_17/B vdd AOI21X1
XFILL_2_2_0 gnd vdd FILL
XXOR2X1_6 XOR2X1_6/A XOR2X1_6/B gnd XOR2X1_6/Y vdd XOR2X1
XCLKBUF1_8 clk gnd CLKBUF1_8/Y vdd CLKBUF1
XFILL_10_1_0 gnd vdd FILL
XNOR2X1_206 INVX2_37/Y INVX1_275/Y gnd NOR2X1_206/Y vdd NOR2X1
XNOR2X1_228 XOR2X1_21/B NOR2X1_227/Y gnd NOR2X1_228/Y vdd NOR2X1
XNOR2X1_217 INVX2_36/Y INVX1_291/Y gnd NOR2X1_218/B vdd NOR2X1
XFILL_18_2_0 gnd vdd FILL
XDFFPOSX1_52 INVX1_112/A CLKBUF1_2/Y OAI21X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_41 INVX2_35/A CLKBUF1_4/Y OAI21X1_75/Y gnd vdd DFFPOSX1
XDFFPOSX1_63 INVX1_59/A CLKBUF1_9/Y NOR2X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_30 NAND2X1_90/A CLKBUF1_3/Y OAI21X1_130/Y gnd vdd DFFPOSX1
XDFFPOSX1_96 INVX1_90/A CLKBUF1_7/Y OAI21X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_85 INVX1_68/A CLKBUF1_1/Y OAI21X1_53/Y gnd vdd DFFPOSX1
XDFFPOSX1_74 INVX1_83/A CLKBUF1_5/Y NOR2X1_49/Y gnd vdd DFFPOSX1
XNAND3X1_335 OAI21X1_358/Y NAND3X1_331/Y NAND3X1_335/C gnd NAND3X1_336/C vdd NAND3X1
XNAND3X1_324 INVX1_303/Y NAND3X1_324/B NAND3X1_324/C gnd NAND3X1_324/Y vdd NAND3X1
XNAND3X1_346 INVX1_92/A AND2X2_45/Y AND2X2_46/Y gnd NAND3X1_346/Y vdd NAND3X1
XNAND3X1_313 XNOR2X1_47/Y NAND3X1_318/B NAND3X1_318/C gnd NAND3X1_317/B vdd NAND3X1
XNAND3X1_302 OAI22X1_21/Y AOI21X1_152/B AOI21X1_152/A gnd NAND3X1_302/Y vdd NAND3X1
XNAND3X1_357 INVX1_310/A NAND3X1_357/B XNOR2X1_52/Y gnd NAND3X1_358/C vdd NAND3X1
XFILL_15_1 gnd vdd FILL
XINVX1_190 AND2X2_26/Y gnd INVX1_190/Y vdd INVX1
XAOI21X1_150 AOI21X1_150/A AOI21X1_150/B XNOR2X1_48/Y gnd AOI21X1_150/Y vdd AOI21X1
XAOI21X1_161 NAND3X1_356/C NAND3X1_356/A INVX1_309/A gnd OAI21X1_389/A vdd AOI21X1
XFILL_7_1_0 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XNAND3X1_132 INVX1_216/A NAND3X1_132/B NAND3X1_132/C gnd AOI21X1_80/B vdd NAND3X1
XNAND3X1_121 NAND2X1_248/Y NAND3X1_119/Y NAND3X1_118/Y gnd NAND3X1_127/C vdd NAND3X1
XNAND3X1_110 INVX2_26/A NAND3X1_108/Y NAND3X1_109/Y gnd AOI21X1_91/B vdd NAND3X1
XNAND3X1_198 INVX1_252/A INVX1_249/Y NAND2X1_324/Y gnd NAND3X1_199/B vdd NAND3X1
XNAND3X1_165 AOI21X1_95/B XOR2X1_14/Y AOI21X1_95/A gnd INVX1_224/A vdd NAND3X1
XNAND3X1_187 INVX1_240/A NAND2X1_307/A NAND2X1_307/B gnd INVX1_248/A vdd NAND3X1
XNAND3X1_143 AOI21X1_85/A NOR2X1_156/Y AOI21X1_85/B gnd NAND3X1_145/B vdd NAND3X1
XNAND3X1_176 gnd gnd INVX2_30/Y gnd INVX1_226/A vdd NAND3X1
XNAND3X1_154 INVX1_129/A AND2X2_28/Y AND2X2_29/Y gnd AOI21X1_88/B vdd NAND3X1
XOAI21X1_328 NOR3X1_11/B NOR3X1_11/C NOR3X1_11/A gnd OAI21X1_328/Y vdd OAI21X1
XOAI21X1_317 NOR2X1_195/B INVX1_260/A INVX1_261/A gnd OAI21X1_317/Y vdd OAI21X1
XOAI21X1_306 INVX2_28/Y INVX1_258/Y NOR2X1_195/B gnd OAI21X1_306/Y vdd OAI21X1
XOAI21X1_339 OR2X2_28/B OR2X2_28/A OAI21X1_339/C gnd INVX1_283/A vdd OAI21X1
XBUFX4_4 start gnd BUFX4_4/Y vdd BUFX4
XNAND2X1_389 INVX1_287/Y NOR2X1_215/Y gnd INVX2_42/A vdd NAND2X1
XNAND2X1_378 AOI21X1_139/B OR2X2_29/Y gnd NAND2X1_380/A vdd NAND2X1
XNAND2X1_367 OR2X2_28/B OR2X2_28/A gnd NAND3X1_270/B vdd NAND2X1
XNAND2X1_356 INVX1_267/A NAND2X1_356/B gnd AND2X2_42/A vdd NAND2X1
XNAND2X1_312 NAND2X1_312/A NAND2X1_312/B gnd XOR2X1_18/A vdd NAND2X1
XNAND2X1_301 INVX1_236/A INVX1_239/A gnd AOI22X1_29/C vdd NAND2X1
XXOR2X1_17 XOR2X1_17/A XOR2X1_17/B gnd INVX1_233/A vdd XOR2X1
XNAND2X1_345 AND2X2_41/B AND2X2_41/A gnd NAND2X1_345/Y vdd NAND2X1
XNAND2X1_334 INVX2_28/A OR2X2_6/B gnd NOR2X1_191/B vdd NAND2X1
XNAND2X1_323 OR2X2_25/A INVX1_250/Y gnd AND2X2_36/B vdd NAND2X1
XNAND3X1_7 INVX1_90/Y INVX1_91/Y NAND3X1_7/C gnd NOR3X1_1/C vdd NAND3X1
XOAI21X1_136 BUFX4_12/Y INVX2_2/Y NAND2X1_96/Y gnd DFFPOSX1_18/D vdd OAI21X1
XOAI21X1_147 NAND3X1_12/Y AOI21X1_29/Y AOI21X1_31/Y gnd NOR2X1_96/B vdd OAI21X1
XOAI21X1_114 NAND3X1_8/Y AOI21X1_17/Y AOI21X1_18/Y gnd NOR2X1_70/B vdd OAI21X1
XOAI21X1_169 INVX2_9/Y INVX1_141/Y NAND3X1_13/Y gnd OR2X2_12/B vdd OAI21X1
XOAI21X1_125 NOR2X1_81/Y NOR2X1_82/Y NOR2X1_80/Y gnd OAI21X1_125/Y vdd OAI21X1
XOAI21X1_103 BUFX4_4/Y INVX1_105/Y OAI21X1_95/C gnd DFFPOSX1_13/D vdd OAI21X1
XOAI21X1_158 NOR2X1_90/Y NOR2X1_91/Y INVX1_123/Y gnd OAI21X1_159/A vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd X0_mag[0] vdd BUFX2
XNAND2X1_197 INVX1_190/Y NAND2X1_197/B gnd NAND3X1_80/C vdd NAND2X1
XNAND2X1_120 gnd gnd gnd INVX1_143/A vdd NAND2X1
XNAND2X1_186 NAND3X1_61/Y NAND3X1_59/Y gnd NAND3X1_66/C vdd NAND2X1
XNAND2X1_164 INVX1_163/Y NOR2X1_122/Y gnd XOR2X1_10/A vdd NAND2X1
XNAND2X1_131 AND2X2_20/B AND2X2_20/A gnd XNOR2X1_20/A vdd NAND2X1
XNAND2X1_153 INVX1_162/Y OAI22X1_7/Y gnd INVX1_174/A vdd NAND2X1
XNAND2X1_175 INVX2_10/A NAND2X1_90/A gnd AOI21X1_61/B vdd NAND2X1
XNAND2X1_142 INVX1_139/A INVX1_153/A gnd OAI21X1_182/C vdd NAND2X1
XINVX2_1 x1[6] gnd INVX2_1/Y vdd INVX2
XAOI21X1_1 OAI21X1_5/Y INVX1_8/Y INVX1_9/Y gnd XNOR2X1_3/A vdd AOI21X1
XXNOR2X1_42 XNOR2X1_42/A INVX1_267/A gnd INVX1_270/A vdd XNOR2X1
XXNOR2X1_20 XNOR2X1_20/A OR2X2_12/B gnd XNOR2X1_21/A vdd XNOR2X1
XXNOR2X1_31 INVX2_20/A XNOR2X1_31/B gnd XNOR2X1_31/Y vdd XNOR2X1
XBUFX2_30 BUFX2_30/A gnd X3_mag[5] vdd BUFX2
XAOI21X1_31 AOI21X1_31/A AOI21X1_30/Y AOI21X1_31/C gnd AOI21X1_31/Y vdd AOI21X1
XAOI21X1_42 OR2X2_9/Y NAND3X1_15/B INVX1_135/Y gnd AOI21X1_42/Y vdd AOI21X1
XAOI21X1_86 AOI21X1_86/A AOI21X1_86/B XNOR2X1_33/Y gnd AOI21X1_87/C vdd AOI21X1
XAOI21X1_53 AOI21X1_56/A AOI21X1_56/B INVX2_15/Y gnd OAI22X1_15/C vdd AOI21X1
XAOI21X1_64 NAND3X1_44/B INVX1_183/Y INVX1_184/Y gnd AOI21X1_64/Y vdd AOI21X1
XAOI21X1_20 NOR2X1_70/B NOR2X1_75/Y AOI21X1_22/A gnd AND2X2_14/A vdd AOI21X1
XAOI21X1_75 INVX1_196/Y AOI21X1_75/B INVX1_206/Y gnd AOI21X1_75/Y vdd AOI21X1
XOAI21X1_4 BUFX4_2/Y INVX1_4/Y OAI21X1_4/C gnd OAI21X1_4/Y vdd OAI21X1
XAOI21X1_97 INVX1_209/Y AOI21X1_97/B AOI21X1_96/Y gnd AOI21X1_97/Y vdd AOI21X1
XFILL_3_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XXOR2X1_7 XOR2X1_7/A XOR2X1_7/B gnd XOR2X1_7/Y vdd XOR2X1
XFILL_10_1_1 gnd vdd FILL
XCLKBUF1_9 clk gnd CLKBUF1_9/Y vdd CLKBUF1
XFILL_18_2_1 gnd vdd FILL
XNOR2X1_207 NOR2X1_207/A NOR2X1_206/Y gnd AOI22X1_42/D vdd NOR2X1
XNOR2X1_218 INVX1_290/Y NOR2X1_218/B gnd NOR2X1_218/Y vdd NOR2X1
XDFFPOSX1_64 XOR2X1_5/A CLKBUF1_7/Y AND2X2_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_42 INVX1_273/A CLKBUF1_7/Y OAI21X1_77/Y gnd vdd DFFPOSX1
XDFFPOSX1_86 INVX1_69/A CLKBUF1_1/Y OAI21X1_54/Y gnd vdd DFFPOSX1
XDFFPOSX1_20 INVX2_23/A CLKBUF1_8/Y DFFPOSX1_20/D gnd vdd DFFPOSX1
XDFFPOSX1_53 INVX1_41/A CLKBUF1_10/Y OAI22X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_75 INVX1_84/A CLKBUF1_5/Y NOR2X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_31 INVX2_16/A CLKBUF1_3/Y DFFPOSX1_31/D gnd vdd DFFPOSX1
XDFFPOSX1_97 INVX1_24/A CLKBUF1_7/Y OAI21X1_17/Y gnd vdd DFFPOSX1
XNAND3X1_314 OAI21X1_375/A NAND3X1_302/Y AOI21X1_157/A gnd AOI21X1_150/A vdd NAND3X1
XNAND3X1_303 INVX2_44/A NAND3X1_298/B NAND3X1_298/C gnd NAND3X1_310/C vdd NAND3X1
XNAND3X1_336 INVX1_295/A NAND3X1_334/Y NAND3X1_336/C gnd NAND3X1_336/Y vdd NAND3X1
XNAND3X1_325 NAND2X1_410/Y NAND3X1_325/B NAND3X1_324/Y gnd NAND3X1_334/A vdd NAND3X1
XNAND3X1_358 OAI21X1_372/Y NAND3X1_358/B NAND3X1_358/C gnd NAND3X1_358/Y vdd NAND3X1
XNAND3X1_347 OAI21X1_380/Y NAND3X1_346/Y XOR2X1_23/Y gnd NAND3X1_351/C vdd NAND3X1
XINVX1_191 INVX1_191/A gnd INVX1_191/Y vdd INVX1
XINVX1_180 INVX1_180/A gnd INVX1_180/Y vdd INVX1
XAOI21X1_140 AND2X2_44/B AOI21X1_140/B NOR2X1_219/A gnd NAND3X1_287/A vdd AOI21X1
XAOI21X1_162 NAND3X1_335/C NAND3X1_331/Y NOR2X1_223/Y gnd AOI21X1_162/Y vdd AOI21X1
XAOI21X1_151 NAND3X1_317/C INVX1_302/A AOI21X1_150/Y gnd XOR2X1_22/A vdd AOI21X1
XFILL_7_1_1 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XNAND3X1_133 INVX1_217/Y AOI21X1_80/A AOI21X1_80/B gnd AOI21X1_94/A vdd NAND3X1
XNAND3X1_166 INVX1_224/A NAND3X1_168/B XNOR2X1_37/Y gnd AOI21X1_98/A vdd NAND3X1
XNAND3X1_111 OAI22X1_18/Y AOI21X1_91/B AOI21X1_91/A gnd NAND3X1_111/Y vdd NAND3X1
XNAND3X1_122 XNOR2X1_32/Y NAND3X1_127/B NAND3X1_127/C gnd NAND3X1_122/Y vdd NAND3X1
XNAND3X1_144 AOI21X1_85/C AOI21X1_96/B AOI21X1_96/A gnd NAND3X1_145/C vdd NAND3X1
XNAND3X1_155 AOI21X1_88/A AOI21X1_88/B XOR2X1_15/Y gnd NAND3X1_155/Y vdd NAND3X1
XNAND3X1_100 INVX2_25/Y INVX1_210/A OR2X2_19/Y gnd AOI22X1_23/D vdd NAND3X1
XNAND3X1_188 INVX1_234/A NAND3X1_191/B INVX1_264/A gnd NAND3X1_190/B vdd NAND3X1
XNAND3X1_199 INVX2_34/Y NAND3X1_199/B NAND3X1_199/C gnd NAND3X1_199/Y vdd NAND3X1
XNAND3X1_177 gnd gnd NOR2X1_168/Y gnd NOR2X1_179/A vdd NAND3X1
XOAI21X1_329 INVX1_245/Y AOI22X1_32/D NAND3X1_234/Y gnd AOI22X1_41/D vdd OAI21X1
XOAI21X1_307 INVX2_28/Y INVX1_258/Y AND2X2_38/Y gnd OAI21X1_307/Y vdd OAI21X1
XOAI21X1_318 INVX2_29/Y INVX1_258/Y OR2X2_27/B gnd AND2X2_40/B vdd OAI21X1
XXOR2X1_18 XOR2X1_18/A XOR2X1_18/B gnd XOR2X1_18/Y vdd XOR2X1
XNAND2X1_302 NAND3X1_180/Y NAND2X1_287/A gnd INVX1_240/A vdd NAND2X1
XBUFX4_5 start gnd BUFX4_5/Y vdd BUFX4
XNAND2X1_379 INVX1_282/A NAND2X1_380/A gnd NAND2X1_379/Y vdd NAND2X1
XNAND2X1_368 NAND3X1_270/B OR2X2_28/Y gnd NAND2X1_368/Y vdd NAND2X1
XNAND2X1_335 INVX1_259/A NOR2X1_193/Y gnd XOR2X1_19/A vdd NAND2X1
XNAND2X1_357 AND2X2_42/B AND2X2_42/A gnd NAND3X1_261/B vdd NAND2X1
XNAND2X1_313 AOI21X1_108/C NAND2X1_313/B gnd NOR2X1_187/B vdd NAND2X1
XNAND2X1_324 AND2X2_36/B AND2X2_36/A gnd NAND2X1_324/Y vdd NAND2X1
XNAND2X1_346 AOI21X1_122/Y AND2X2_40/Y gnd NAND2X1_346/Y vdd NAND2X1
XNAND3X1_8 INVX1_115/Y NAND3X1_8/B NOR2X1_66/Y gnd NAND3X1_8/Y vdd NAND3X1
XOAI21X1_115 OAI21X1_111/Y NOR2X1_71/A INVX1_118/Y gnd AOI21X1_19/C vdd OAI21X1
XOAI21X1_126 INVX1_56/Y INVX1_85/A OAI21X1_125/Y gnd AOI21X1_22/C vdd OAI21X1
XOAI21X1_137 BUFX4_13/Y INVX2_3/Y NAND2X1_97/Y gnd DFFPOSX1_19/D vdd OAI21X1
XOAI21X1_104 BUFX4_4/Y INVX1_106/Y NAND2X1_59/Y gnd DFFPOSX1_14/D vdd OAI21X1
XOAI21X1_148 NOR2X1_70/A INVX1_130/Y BUFX4_9/Y gnd OAI21X1_149/B vdd OAI21X1
XOAI21X1_159 OAI21X1_159/A AND2X2_16/A AOI21X1_38/Y gnd AND2X2_17/A vdd OAI21X1
XNAND2X1_132 INVX1_136/Y INVX1_143/Y gnd OR2X2_10/B vdd NAND2X1
XBUFX2_2 BUFX2_2/A gnd X0_mag[1] vdd BUFX2
XNAND2X1_121 gnd gnd gnd OAI21X1_167/C vdd NAND2X1
XNAND2X1_110 INVX2_33/A BUFX4_11/Y gnd OAI21X1_152/C vdd NAND2X1
XNAND2X1_143 INVX2_9/A NAND3X1_20/C gnd OAI21X1_183/C vdd NAND2X1
XNAND2X1_154 gnd gnd gnd AND2X2_22/A vdd NAND2X1
XNAND2X1_176 OR2X2_14/A XNOR2X1_28/Y gnd AOI22X1_11/C vdd NAND2X1
XNAND2X1_165 NAND2X1_165/A XOR2X1_10/A gnd OR2X2_13/A vdd NAND2X1
XNAND2X1_198 INVX2_18/A INVX1_104/A gnd INVX1_192/A vdd NAND2X1
XNAND2X1_187 XNOR2X1_30/B AOI21X1_65/Y gnd NAND3X1_69/A vdd NAND2X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XAOI21X1_2 OAI21X1_5/Y NOR2X1_6/Y AOI21X1_2/C gnd AND2X2_1/A vdd AOI21X1
XXNOR2X1_10 AOI21X1_9/A INVX1_8/A gnd OAI21X1_61/B vdd XNOR2X1
XXNOR2X1_32 XNOR2X1_32/A INVX1_212/Y gnd XNOR2X1_32/Y vdd XNOR2X1
XXNOR2X1_43 NOR2X1_191/Y INVX1_267/Y gnd INVX1_268/A vdd XNOR2X1
XXNOR2X1_21 XNOR2X1_21/A INVX1_158/A gnd OR2X2_11/A vdd XNOR2X1
XBUFX2_31 BUFX2_31/A gnd X3_mag[6] vdd BUFX2
XBUFX2_20 BUFX2_20/A gnd X2_mag[3] vdd BUFX2
XOAI21X1_5 INVX1_5/Y x3[1] OAI21X1_5/C gnd OAI21X1_5/Y vdd OAI21X1
XAOI21X1_10 XOR2X1_2/B NOR2X1_42/Y NOR2X1_43/Y gnd AND2X2_8/B vdd AOI21X1
XAOI21X1_76 INVX1_198/Y NAND3X1_85/C AOI21X1_76/C gnd AOI21X1_76/Y vdd AOI21X1
XAOI21X1_43 AOI21X1_43/A NAND3X1_16/Y INVX1_140/A gnd AOI21X1_67/A vdd AOI21X1
XAOI21X1_87 AOI21X1_87/A INVX1_216/A AOI21X1_87/C gnd XOR2X1_14/A vdd AOI21X1
XAOI21X1_98 AOI21X1_98/A AOI21X1_98/B AOI21X1_97/Y gnd AOI21X1_98/Y vdd AOI21X1
XAOI21X1_54 AOI21X1_57/A NAND3X1_36/Y INVX1_173/A gnd OAI22X1_14/A vdd AOI21X1
XAOI21X1_65 NAND3X1_42/B NAND3X1_42/C INVX1_174/Y gnd AOI21X1_65/Y vdd AOI21X1
XAOI21X1_21 NOR2X1_84/Y INVX1_120/Y BUFX4_11/Y gnd AOI22X1_2/D vdd AOI21X1
XAOI21X1_32 NOR2X1_96/B NOR2X1_69/Y NOR2X1_68/Y gnd XNOR2X1_15/A vdd AOI21X1
XFILL_3_2 gnd vdd FILL
XFILL_2_2_2 gnd vdd FILL
XXOR2X1_8 XOR2X1_9/B XOR2X1_8/B gnd XOR2X1_8/Y vdd XOR2X1
XFILL_10_1_2 gnd vdd FILL
XFILL_18_2_2 gnd vdd FILL
XNOR2X1_219 NOR2X1_219/A NOR2X1_219/B gnd AND2X2_44/A vdd NOR2X1
XNOR2X1_208 NOR2X1_208/A INVX1_277/Y gnd NOR2X1_208/Y vdd NOR2X1
XDFFPOSX1_43 INVX2_39/A CLKBUF1_4/Y OAI21X1_79/Y gnd vdd DFFPOSX1
XDFFPOSX1_98 INVX2_2/A CLKBUF1_4/Y OAI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_65 INVX1_72/A CLKBUF1_2/Y OAI21X1_57/Y gnd vdd DFFPOSX1
XDFFPOSX1_21 INVX1_193/A CLKBUF1_8/Y DFFPOSX1_21/D gnd vdd DFFPOSX1
XDFFPOSX1_87 INVX1_70/A CLKBUF1_8/Y OAI21X1_55/Y gnd vdd DFFPOSX1
XDFFPOSX1_54 INVX1_114/A CLKBUF1_10/Y OAI21X1_37/Y gnd vdd DFFPOSX1
XDFFPOSX1_32 INVX1_127/A CLKBUF1_3/Y AOI22X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_76 INVX1_85/A CLKBUF1_9/Y NOR2X1_51/Y gnd vdd DFFPOSX1
XDFFPOSX1_10 INVX2_19/A CLKBUF1_5/Y DFFPOSX1_10/D gnd vdd DFFPOSX1
XNAND3X1_326 INVX1_297/A NAND3X1_326/B NAND3X1_326/C gnd NAND3X1_326/Y vdd NAND3X1
XNAND3X1_337 NAND2X1_400/Y NAND3X1_342/B NAND3X1_336/Y gnd OR2X2_34/A vdd NAND3X1
XNAND3X1_304 INVX2_44/Y NAND3X1_301/B NAND3X1_301/C gnd NAND3X1_304/Y vdd NAND3X1
XNAND3X1_315 NAND3X1_308/A NAND3X1_315/B NAND3X1_309/Y gnd AOI21X1_150/B vdd NAND3X1
XNAND3X1_348 INVX1_307/Y NAND2X1_434/Y NAND3X1_351/C gnd NAND3X1_349/B vdd NAND3X1
XNAND3X1_359 INVX1_310/A NAND3X1_357/B NAND2X1_441/Y gnd NAND3X1_360/B vdd NAND3X1
XINVX1_170 INVX1_170/A gnd INVX1_170/Y vdd INVX1
XINVX1_181 INVX1_181/A gnd INVX1_181/Y vdd INVX1
XINVX1_192 INVX1_192/A gnd INVX1_192/Y vdd INVX1
XAOI21X1_141 NAND3X1_287/B NAND3X1_287/C AOI21X1_141/C gnd INVX1_306/A vdd AOI21X1
XAOI21X1_163 INVX1_295/Y NAND3X1_333/C AOI21X1_162/Y gnd AOI21X1_163/Y vdd AOI21X1
XAOI21X1_152 AOI21X1_152/A AOI21X1_152/B OAI22X1_21/Y gnd OAI21X1_375/B vdd AOI21X1
XAOI21X1_130 INVX1_247/Y NAND3X1_230/B AOI21X1_130/C gnd AOI21X1_130/Y vdd AOI21X1
XFILL_7_1_2 gnd vdd FILL
XFILL_15_0_2 gnd vdd FILL
XNAND3X1_156 INVX1_221/Y NAND2X1_257/Y NAND3X1_155/Y gnd NAND3X1_157/A vdd NAND3X1
XNAND3X1_189 INVX1_234/Y NAND3X1_189/B NAND3X1_189/C gnd NAND3X1_189/Y vdd NAND3X1
XNAND3X1_123 NAND2X1_248/Y NAND3X1_111/Y NAND3X1_114/Y gnd AOI21X1_86/A vdd NAND3X1
XNAND3X1_134 AOI21X1_94/B NAND3X1_130/Y AOI21X1_94/A gnd AOI21X1_85/A vdd NAND3X1
XNAND3X1_112 INVX2_26/A AOI21X1_89/A NAND2X1_244/Y gnd NAND3X1_112/Y vdd NAND3X1
XNAND3X1_167 AOI21X1_99/C AOI21X1_98/B AOI21X1_98/A gnd NAND3X1_167/Y vdd NAND3X1
XNAND3X1_178 NAND3X1_178/A NOR2X1_170/Y NAND3X1_178/C gnd NAND3X1_178/Y vdd NAND3X1
XNAND3X1_145 INVX1_209/A NAND3X1_145/B NAND3X1_145/C gnd NAND3X1_146/C vdd NAND3X1
XNAND3X1_101 AOI22X1_23/C AOI22X1_23/D NAND3X1_101/C gnd AOI21X1_78/B vdd NAND3X1
XFILL_20_1 gnd vdd FILL
XOAI21X1_319 INVX1_269/A OAI21X1_319/B INVX1_268/Y gnd AND2X2_41/A vdd OAI21X1
XOAI21X1_308 INVX1_260/A INVX1_261/Y NOR2X1_195/B gnd AND2X2_39/A vdd OAI21X1
XBUFX4_6 start gnd BUFX4_6/Y vdd BUFX4
XNAND2X1_314 NAND3X1_194/B NAND3X1_194/C gnd AOI22X1_39/B vdd NAND2X1
XXOR2X1_19 XOR2X1_19/A XOR2X1_19/B gnd OR2X2_26/A vdd XOR2X1
XNAND2X1_336 NAND2X1_336/A XOR2X1_19/A gnd INVX1_262/A vdd NAND2X1
XNAND2X1_325 NOR3X1_8/B INVX1_266/A gnd AOI22X1_34/D vdd NAND2X1
XNAND2X1_303 INVX2_29/A INVX1_242/A gnd NOR2X1_183/B vdd NAND2X1
XNAND2X1_369 INVX1_276/Y NAND2X1_368/Y gnd AOI21X1_134/A vdd NAND2X1
XNAND2X1_358 INVX1_246/A NAND3X1_234/Y gnd AOI22X1_37/C vdd NAND2X1
XNOR3X1_10 INVX1_270/A NOR3X1_11/B NOR3X1_11/C gnd NOR3X1_10/Y vdd NOR3X1
XNAND2X1_347 NAND2X1_343/Y OAI21X1_320/Y gnd NAND2X1_348/B vdd NAND2X1
XNAND3X1_9 INVX1_47/A INVX1_78/Y NAND3X1_9/C gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_138 BUFX4_12/Y INVX1_27/Y NAND2X1_98/Y gnd DFFPOSX1_20/D vdd OAI21X1
XOAI21X1_105 BUFX4_4/Y INVX1_107/Y NAND2X1_60/Y gnd DFFPOSX1_15/D vdd OAI21X1
XOAI21X1_149 NOR2X1_96/Y OAI21X1_149/B NAND2X1_107/Y gnd DFFPOSX1_1/D vdd OAI21X1
XOAI21X1_127 INVX1_121/A AOI21X1_19/Y INVX1_122/A gnd NOR2X1_89/B vdd OAI21X1
XBUFX2_3 BUFX2_3/A gnd X0_mag[2] vdd BUFX2
XOAI21X1_116 NOR2X1_69/Y AOI21X1_19/Y BUFX4_5/Y gnd OAI21X1_116/Y vdd OAI21X1
XNAND2X1_133 OAI21X1_173/Y OR2X2_10/Y gnd INVX1_158/A vdd NAND2X1
XNAND2X1_155 gnd gnd gnd AND2X2_22/B vdd NAND2X1
XNAND2X1_177 XOR2X1_9/Y INVX1_177/Y gnd AOI22X1_11/D vdd NAND2X1
XNAND2X1_166 OR2X2_13/B OR2X2_13/A gnd AND2X2_23/B vdd NAND2X1
XNAND2X1_122 NAND2X1_122/A NAND3X1_13/Y gnd OR2X2_8/A vdd NAND2X1
XNAND2X1_144 INVX1_154/A AND2X2_21/Y gnd AOI21X1_45/A vdd NAND2X1
XNAND2X1_111 NOR2X1_69/Y INVX2_5/A gnd NOR2X1_97/A vdd NAND2X1
XNAND2X1_100 AOI22X1_21/D BUFX4_13/Y gnd NAND2X1_100/Y vdd NAND2X1
XNAND2X1_188 AOI21X1_66/B AOI21X1_66/A gnd NAND3X1_71/C vdd NAND2X1
XNAND2X1_199 NAND3X1_82/A NAND3X1_82/C gnd NAND2X1_199/Y vdd NAND2X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XAOI21X1_3 NOR2X1_9/Y NOR2X1_4/Y NOR2X1_8/Y gnd AOI21X1_3/Y vdd AOI21X1
XINVX1_90 INVX1_90/A gnd INVX1_90/Y vdd INVX1
XXNOR2X1_11 NOR2X1_64/A INVX1_73/A gnd XNOR2X1_11/Y vdd XNOR2X1
XBUFX2_10 BUFX2_10/A gnd X1_mag[1] vdd BUFX2
XXNOR2X1_33 XNOR2X1_32/A INVX1_212/A gnd XNOR2X1_33/Y vdd XNOR2X1
XXNOR2X1_22 XNOR2X1_22/A AOI21X1_67/A gnd XNOR2X1_22/Y vdd XNOR2X1
XXNOR2X1_44 NOR3X1_11/A XNOR2X1_44/B gnd XNOR2X1_44/Y vdd XNOR2X1
XBUFX2_21 BUFX2_21/A gnd X2_mag[4] vdd BUFX2
XBUFX2_32 BUFX2_32/A gnd X3_mag[7] vdd BUFX2
XNOR2X1_1 x1[0] INVX1_2/Y gnd NOR2X1_1/Y vdd NOR2X1
XFILL_22_1_0 gnd vdd FILL
XAOI21X1_11 NAND3X1_6/B INVX1_81/Y INVX1_25/A gnd OAI22X1_6/C vdd AOI21X1
XOAI21X1_6 BUFX4_15/Y OAI21X1_6/B NAND2X1_5/Y gnd OAI21X1_6/Y vdd OAI21X1
XAOI21X1_99 AOI21X1_99/A AOI21X1_99/B AOI21X1_99/C gnd AOI21X1_99/Y vdd AOI21X1
XAOI21X1_88 AOI21X1_88/A AOI21X1_88/B XOR2X1_15/Y gnd AOI21X1_88/Y vdd AOI21X1
XAOI21X1_66 AOI21X1_66/A AOI21X1_66/B NAND3X1_69/Y gnd AOI21X1_66/Y vdd AOI21X1
XAOI21X1_55 AOI21X1_58/A NAND3X1_40/Y INVX1_173/Y gnd OAI22X1_14/B vdd AOI21X1
XAOI21X1_22 AOI21X1_22/A NOR2X1_85/Y AOI21X1_22/C gnd INVX1_122/A vdd AOI21X1
XAOI21X1_44 NAND3X1_21/C NAND3X1_21/B INVX1_156/A gnd OAI22X1_7/B vdd AOI21X1
XAOI21X1_33 INVX2_5/A NOR2X1_68/Y NOR2X1_73/Y gnd AOI21X1_33/Y vdd AOI21X1
XAOI21X1_77 NAND3X1_95/B NAND3X1_95/C NAND3X1_85/B gnd INVX1_220/A vdd AOI21X1
XFILL_5_2_0 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XFILL_3_3 gnd vdd FILL
XXOR2X1_9 XOR2X1_9/A XOR2X1_9/B gnd XOR2X1_9/Y vdd XOR2X1
XNOR2X1_209 INVX2_35/Y INVX1_279/Y gnd NOR2X1_209/Y vdd NOR2X1
XDFFPOSX1_11 INVX1_103/A CLKBUF1_10/Y DFFPOSX1_11/D gnd vdd DFFPOSX1
XDFFPOSX1_44 INVX2_41/A CLKBUF1_7/Y OAI21X1_81/Y gnd vdd DFFPOSX1
XDFFPOSX1_66 INVX1_73/A CLKBUF1_1/Y OAI21X1_59/Y gnd vdd DFFPOSX1
XDFFPOSX1_99 INVX2_3/A CLKBUF1_8/Y OAI21X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_55 INVX1_47/A CLKBUF1_1/Y OAI22X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_33 INVX2_36/A CLKBUF1_4/Y OAI21X1_91/Y gnd vdd DFFPOSX1
XDFFPOSX1_77 INVX1_86/A CLKBUF1_3/Y NOR2X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_88 INVX1_71/A CLKBUF1_5/Y OAI21X1_56/Y gnd vdd DFFPOSX1
XDFFPOSX1_22 AOI22X1_21/D CLKBUF1_5/Y DFFPOSX1_22/D gnd vdd DFFPOSX1
XFILL_2_0_0 gnd vdd FILL
XNAND3X1_338 INVX1_295/A NAND3X1_333/B NAND3X1_333/C gnd NAND3X1_343/B vdd NAND3X1
XNAND3X1_327 INVX1_303/Y NAND3X1_327/B NAND3X1_327/C gnd NAND3X1_327/Y vdd NAND3X1
XNAND3X1_316 XNOR2X1_48/Y AOI21X1_150/A AOI21X1_150/B gnd NAND3X1_317/C vdd NAND3X1
XNAND3X1_305 AOI22X1_51/Y NAND3X1_304/Y NAND3X1_310/C gnd AOI21X1_157/A vdd NAND3X1
XNAND3X1_349 NAND3X1_349/A NAND3X1_349/B OAI21X1_381/Y gnd NAND2X1_436/A vdd NAND3X1
XFILL_18_0_0 gnd vdd FILL
XINVX1_160 NOR3X1_6/A gnd INVX1_160/Y vdd INVX1
XINVX1_182 XOR2X1_11/Y gnd INVX1_182/Y vdd INVX1
XINVX1_171 INVX1_171/A gnd INVX1_171/Y vdd INVX1
XINVX1_193 INVX1_193/A gnd INVX1_193/Y vdd INVX1
XAOI21X1_142 AOI21X1_142/A OAI21X1_374/C INVX2_42/Y gnd AOI21X1_142/Y vdd AOI21X1
XAOI21X1_153 NAND3X1_298/B INVX2_44/Y NOR2X1_224/Y gnd NAND2X1_427/A vdd AOI21X1
XAOI21X1_164 NAND3X1_358/C NAND3X1_358/B AOI21X1_163/Y gnd OAI22X1_22/A vdd AOI21X1
XAOI21X1_131 OAI21X1_312/C NAND3X1_228/B OAI21X1_312/A gnd AOI21X1_131/Y vdd AOI21X1
XAOI21X1_120 OR2X2_27/Y AND2X2_40/B OAI21X1_317/Y gnd INVX1_269/A vdd AOI21X1
XNAND3X1_168 INVX1_224/A NAND3X1_168/B NAND3X1_168/C gnd AOI21X1_99/B vdd NAND3X1
XNAND3X1_124 NAND2X1_247/Y NAND3X1_119/Y NAND3X1_118/Y gnd AOI21X1_86/B vdd NAND3X1
XNAND3X1_113 INVX2_26/Y NAND3X1_108/Y NAND3X1_109/Y gnd NAND3X1_113/Y vdd NAND3X1
XNAND3X1_157 NAND3X1_157/A NAND3X1_157/B NAND3X1_157/C gnd AOI21X1_92/A vdd NAND3X1
XNAND3X1_179 AND2X2_33/Y AOI21X1_101/B OR2X2_21/Y gnd INVX1_230/A vdd NAND3X1
XNAND3X1_135 INVX1_211/A OAI21X1_248/Y NAND3X1_105/Y gnd NAND2X1_251/A vdd NAND3X1
XNAND3X1_102 INVX2_25/Y AND2X2_28/Y OR2X2_19/Y gnd AOI22X1_23/A vdd NAND3X1
XNAND3X1_146 NAND2X1_228/Y NAND3X1_146/B NAND3X1_146/C gnd OR2X2_20/A vdd NAND3X1
XBUFX4_7 start gnd BUFX4_7/Y vdd BUFX4
XOAI21X1_309 NOR2X1_191/Y NOR2X1_192/Y INVX1_259/Y gnd NAND2X1_336/A vdd OAI21X1
XFILL_13_1 gnd vdd FILL
XNAND2X1_337 NAND2X1_337/A OAI21X1_310/Y gnd NAND2X1_337/Y vdd NAND2X1
XNAND2X1_315 NOR2X1_187/Y AOI22X1_39/B gnd NAND2X1_316/A vdd NAND2X1
XNAND2X1_359 NAND3X1_237/B NAND3X1_236/Y gnd NAND2X1_359/Y vdd NAND2X1
XNAND2X1_326 NAND2X1_326/A NAND2X1_326/B gnd OAI21X1_312/C vdd NAND2X1
XNAND2X1_304 INVX1_238/Y NOR2X1_183/Y gnd INVX2_34/A vdd NAND2X1
XNAND2X1_348 NAND2X1_346/Y NAND2X1_348/B gnd NAND2X1_348/Y vdd NAND2X1
XNOR3X1_11 NOR3X1_11/A NOR3X1_11/B NOR3X1_11/C gnd NOR3X1_11/Y vdd NOR3X1
XOAI21X1_106 BUFX4_4/Y INVX1_108/Y OAI21X1_98/C gnd DFFPOSX1_16/D vdd OAI21X1
XOAI21X1_128 INVX1_123/Y AOI21X1_23/Y BUFX4_7/Y gnd OAI21X1_128/Y vdd OAI21X1
XOAI21X1_117 NOR2X1_70/Y OAI21X1_116/Y NAND2X1_78/Y gnd OAI21X1_117/Y vdd OAI21X1
XOAI21X1_139 BUFX4_14/Y INVX1_28/Y NAND2X1_99/Y gnd DFFPOSX1_21/D vdd OAI21X1
XBUFX2_4 BUFX2_4/A gnd X0_mag[3] vdd BUFX2
XNAND2X1_101 AND2X2_28/B BUFX4_13/Y gnd NAND2X1_101/Y vdd NAND2X1
XNAND2X1_123 OR2X2_8/B OR2X2_8/A gnd NAND3X1_14/B vdd NAND2X1
XNAND2X1_134 OR2X2_11/B OR2X2_11/A gnd INVX2_11/A vdd NAND2X1
XNAND2X1_189 NAND3X1_73/Y NAND3X1_75/Y gnd NAND2X1_189/Y vdd NAND2X1
XNAND2X1_167 AND2X2_23/B OR2X2_13/Y gnd NAND3X1_36/A vdd NAND2X1
XNAND2X1_156 gnd gnd gnd INVX1_163/A vdd NAND2X1
XNAND2X1_178 XOR2X1_10/A XNOR2X1_27/Y gnd AOI22X1_12/B vdd NAND2X1
XNAND2X1_112 INVX1_242/A BUFX4_10/Y gnd NAND2X1_112/Y vdd NAND2X1
XNAND2X1_145 AND2X2_21/B AND2X2_21/A gnd NAND2X1_145/Y vdd NAND2X1
XAOI21X1_4 AND2X2_2/Y AOI21X1_4/B AOI21X1_4/C gnd AND2X2_3/A vdd AOI21X1
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XXNOR2X1_12 INVX1_114/A INVX1_113/A gnd NAND3X1_8/B vdd XNOR2X1
XXNOR2X1_23 XOR2X1_7/A XOR2X1_7/B gnd XNOR2X1_23/Y vdd XNOR2X1
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XBUFX2_11 BUFX2_11/A gnd X1_mag[2] vdd BUFX2
XXNOR2X1_34 XNOR2X1_34/A OAI22X1_18/Y gnd INVX1_216/A vdd XNOR2X1
XBUFX2_33 DFFSR_1/Q gnd done vdd BUFX2
XBUFX2_22 BUFX2_22/A gnd X2_mag[5] vdd BUFX2
XXNOR2X1_45 NOR3X1_11/A XNOR2X1_45/B gnd XNOR2X1_45/Y vdd XNOR2X1
XNOR2X1_2 x3[0] INVX1_3/Y gnd NOR2X1_2/Y vdd NOR2X1
XFILL_22_1_1 gnd vdd FILL
XAOI21X1_12 BUFX4_12/Y INVX1_82/Y NOR2X1_48/Y gnd AOI21X1_12/Y vdd AOI21X1
XAOI21X1_34 XNOR2X1_16/A NOR2X1_85/A NOR2X1_77/Y gnd OR2X2_5/A vdd AOI21X1
XAOI21X1_23 NOR2X1_70/B INVX1_121/Y INVX1_122/Y gnd AOI21X1_23/Y vdd AOI21X1
XOAI21X1_7 BUFX4_15/Y OAI21X1_7/B OAI21X1_7/C gnd OAI21X1_7/Y vdd OAI21X1
XAOI21X1_67 AOI21X1_67/A AOI21X1_67/B NOR3X1_6/Y gnd AOI21X1_67/Y vdd AOI21X1
XAOI21X1_89 AOI21X1_89/A INVX2_26/Y AOI21X1_89/C gnd AOI21X1_89/Y vdd AOI21X1
XAOI21X1_78 AOI21X1_78/A AOI21X1_78/B INVX2_24/Y gnd AOI21X1_78/Y vdd AOI21X1
XAOI21X1_56 AOI21X1_56/A AOI21X1_56/B INVX2_15/A gnd OAI22X1_13/C vdd AOI21X1
XAOI21X1_45 AOI21X1_45/A AOI21X1_45/B INVX1_155/A gnd OAI22X1_9/C vdd AOI21X1
XFILL_5_2_1 gnd vdd FILL
XFILL_13_1_1 gnd vdd FILL
XOAI22X1_20 INVX1_243/A INVX1_257/A INVX1_256/A INVX1_255/A gnd INVX1_259/A vdd OAI22X1
XFILL_1_1 gnd vdd FILL
XDFFPOSX1_45 INVX1_279/A CLKBUF1_7/Y OAI21X1_83/Y gnd vdd DFFPOSX1
XDFFPOSX1_23 AND2X2_28/B CLKBUF1_8/Y DFFPOSX1_23/D gnd vdd DFFPOSX1
XDFFPOSX1_12 INVX1_104/A CLKBUF1_5/Y DFFPOSX1_12/D gnd vdd DFFPOSX1
XDFFPOSX1_34 INVX2_37/A CLKBUF1_9/Y OAI21X1_92/Y gnd vdd DFFPOSX1
XDFFPOSX1_56 INVX1_116/A CLKBUF1_1/Y OAI21X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_67 INVX1_110/A CLKBUF1_2/Y OAI21X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_89 INVX1_1/A CLKBUF1_2/Y OAI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_78 INVX1_87/A CLKBUF1_3/Y NOR2X1_53/Y gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XNAND3X1_339 INVX1_295/Y NAND3X1_334/Y NAND3X1_336/C gnd NAND3X1_343/C vdd NAND3X1
XNAND3X1_328 INVX1_303/A NAND3X1_324/B NAND3X1_324/C gnd NAND3X1_329/C vdd NAND3X1
XNAND3X1_306 INVX1_96/A INVX1_95/A INVX1_97/A gnd INVX1_301/A vdd NAND3X1
XNAND3X1_317 INVX1_302/A NAND3X1_317/B NAND3X1_317/C gnd NAND3X1_327/B vdd NAND3X1
XFILL_18_0_1 gnd vdd FILL
XINVX1_183 NOR3X1_5/A gnd INVX1_183/Y vdd INVX1
XINVX1_172 INVX1_172/A gnd OR2X2_13/B vdd INVX1
XINVX1_161 INVX1_161/A gnd INVX1_161/Y vdd INVX1
XINVX1_150 XOR2X1_6/B gnd INVX1_150/Y vdd INVX1
XINVX1_194 INVX1_194/A gnd INVX1_194/Y vdd INVX1
XAOI21X1_110 INVX1_249/Y INVX1_252/A NAND2X1_324/Y gnd NOR3X1_9/C vdd AOI21X1
XAOI21X1_132 NAND3X1_255/C NAND3X1_255/B AOI21X1_131/Y gnd AOI21X1_132/Y vdd AOI21X1
XAOI21X1_121 INVX1_261/A AND2X2_39/B NAND2X1_343/Y gnd OAI21X1_319/B vdd AOI21X1
XAOI21X1_154 INVX2_43/Y INVX2_41/A NOR2X1_221/Y gnd AOI21X1_154/Y vdd AOI21X1
XAOI21X1_143 INVX1_95/A INVX1_97/A INVX1_96/A gnd INVX1_300/A vdd AOI21X1
XAOI21X1_165 NAND3X1_360/C NAND3X1_360/B OAI21X1_372/Y gnd OAI22X1_22/B vdd AOI21X1
XNAND3X1_114 AOI22X1_25/Y NAND3X1_113/Y NAND3X1_112/Y gnd NAND3X1_114/Y vdd NAND3X1
XNAND3X1_103 INVX2_25/Y OR2X2_19/Y INVX1_210/Y gnd AOI22X1_22/D vdd NAND3X1
XNAND3X1_158 INVX1_221/A NAND2X1_257/Y NAND3X1_155/Y gnd NAND3X1_159/A vdd NAND3X1
XNAND3X1_136 INVX1_217/Y AOI21X1_81/A AOI21X1_81/B gnd NAND3X1_136/Y vdd NAND3X1
XNAND3X1_125 XNOR2X1_33/Y AOI21X1_86/A AOI21X1_86/B gnd AOI21X1_87/A vdd NAND3X1
XNAND3X1_169 AOI21X1_97/Y AOI21X1_99/B AOI21X1_99/A gnd NAND3X1_169/Y vdd NAND3X1
XNAND3X1_147 INVX1_209/A NAND3X1_142/B AOI21X1_97/B gnd NAND3X1_149/B vdd NAND3X1
XFILL_13_2 gnd vdd FILL
XBUFX4_8 start gnd BUFX4_8/Y vdd BUFX4
XNAND2X1_316 NAND2X1_316/A NAND3X1_196/Y gnd XNOR2X1_41/B vdd NAND2X1
XNAND2X1_338 NAND2X1_338/A NAND2X1_338/B gnd XNOR2X1_41/A vdd NAND2X1
XNAND2X1_327 OAI21X1_290/Y NAND2X1_307/B gnd INVX1_263/A vdd NAND2X1
XNAND2X1_349 AND2X2_40/Y OAI21X1_320/Y gnd NAND2X1_351/B vdd NAND2X1
XNAND2X1_305 INVX2_29/A INVX1_131/A gnd INVX1_243/A vdd NAND2X1
XNOR3X1_12 INVX2_42/A NOR3X1_12/B NOR3X1_12/C gnd NOR3X1_12/Y vdd NOR3X1
XOAI21X1_107 NOR2X1_63/Y NOR2X1_64/Y NAND2X1_62/Y gnd AOI21X1_17/B vdd OAI21X1
XOAI21X1_118 NOR2X1_69/Y AOI21X1_19/Y NAND2X1_85/Y gnd AND2X2_13/A vdd OAI21X1
XOAI21X1_129 OAI21X1_128/Y NOR2X1_89/Y NAND2X1_88/Y gnd OAI21X1_129/Y vdd OAI21X1
XBUFX2_5 BUFX2_5/A gnd X0_mag[4] vdd BUFX2
XNAND2X1_102 INVX1_31/A INVX1_72/A gnd OAI21X1_143/A vdd NAND2X1
XNAND2X1_124 NAND3X1_14/B OR2X2_8/Y gnd NAND2X1_124/Y vdd NAND2X1
XNAND2X1_168 NAND3X1_51/Y NAND3X1_54/Y gnd XNOR2X1_24/A vdd NAND2X1
XNAND2X1_157 INVX1_163/A NOR2X1_119/Y gnd AOI22X1_7/A vdd NAND2X1
XNAND2X1_179 INVX1_176/Y XOR2X1_8/Y gnd AOI22X1_12/A vdd NAND2X1
XNAND2X1_135 OR2X2_12/B OR2X2_12/A gnd INVX1_157/A vdd NAND2X1
XNAND2X1_146 INVX1_154/Y NAND2X1_145/Y gnd AOI21X1_45/B vdd NAND2X1
XNAND2X1_113 NOR2X1_85/A OR2X2_5/B gnd NOR2X1_97/B vdd NAND2X1
XNOR2X1_190 NOR3X1_8/A NOR3X1_8/C gnd INVX1_266/A vdd NOR2X1
XAOI21X1_5 INVX1_60/A INVX1_46/A AND2X2_4/Y gnd AOI21X1_5/Y vdd AOI21X1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XXNOR2X1_46 INVX2_38/A XNOR2X1_46/B gnd XNOR2X1_46/Y vdd XNOR2X1
XXNOR2X1_13 INVX1_112/A INVX1_111/A gnd NOR2X1_95/A vdd XNOR2X1
XXNOR2X1_24 XNOR2X1_24/A AOI21X1_60/B gnd XNOR2X1_24/Y vdd XNOR2X1
XXNOR2X1_35 XNOR2X1_35/A AOI21X1_84/B gnd XNOR2X1_35/Y vdd XNOR2X1
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XBUFX2_12 BUFX2_12/A gnd X1_mag[3] vdd BUFX2
XBUFX2_23 BUFX2_23/A gnd X2_mag[6] vdd BUFX2
XNOR2X1_3 x1[4] INVX1_13/Y gnd NOR2X1_3/Y vdd NOR2X1
XFILL_22_1_2 gnd vdd FILL
XAOI21X1_13 NAND3X1_7/C INVX1_90/Y INVX1_24/Y gnd OAI21X1_75/A vdd AOI21X1
XAOI21X1_68 INVX1_185/A NAND3X1_50/Y NOR3X1_6/B gnd AOI21X1_68/Y vdd AOI21X1
XAOI21X1_57 AOI21X1_57/A NAND3X1_36/Y INVX1_173/Y gnd NOR3X1_5/A vdd AOI21X1
XAOI21X1_35 OR2X2_5/A OR2X2_5/B BUFX4_11/Y gnd AOI22X1_4/C vdd AOI21X1
XAOI21X1_46 AOI21X1_46/A AOI21X1_46/B INVX1_155/Y gnd OAI22X1_9/D vdd AOI21X1
XAOI21X1_24 NOR2X1_89/B AND2X2_16/B NOR2X1_86/Y gnd XNOR2X1_14/A vdd AOI21X1
XOAI21X1_8 INVX1_9/A INVX1_16/Y OAI21X1_8/C gnd AOI21X1_2/C vdd OAI21X1
XAOI21X1_79 INVX1_103/A INVX1_105/A INVX1_104/A gnd INVX1_214/A vdd AOI21X1
XFILL_5_2_2 gnd vdd FILL
XOAI22X1_21 INVX1_290/A INVX2_44/A INVX1_298/A OAI22X1_21/D gnd OAI22X1_21/Y vdd OAI22X1
XFILL_13_1_2 gnd vdd FILL
XOAI22X1_10 OAI22X1_7/B OAI22X1_7/A OAI22X1_8/C OAI22X1_8/D gnd OAI22X1_10/Y vdd OAI22X1
XINVX1_310 INVX1_310/A gnd INVX1_310/Y vdd INVX1
XOAI21X1_290 INVX1_243/Y NOR2X1_185/Y AOI22X1_28/B gnd OAI21X1_290/Y vdd OAI21X1
XDFFPOSX1_46 AOI22X1_47/D CLKBUF1_7/Y OAI21X1_86/Y gnd vdd DFFPOSX1
XDFFPOSX1_35 INVX1_95/A CLKBUF1_4/Y OAI21X1_93/Y gnd vdd DFFPOSX1
XDFFPOSX1_68 INVX1_111/A CLKBUF1_2/Y OAI21X1_62/Y gnd vdd DFFPOSX1
XDFFPOSX1_57 INVX1_52/A CLKBUF1_8/Y AOI22X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_13 INVX1_105/A CLKBUF1_10/Y DFFPOSX1_13/D gnd vdd DFFPOSX1
XDFFPOSX1_24 INVX1_129/A CLKBUF1_10/Y DFFPOSX1_24/D gnd vdd DFFPOSX1
XDFFPOSX1_79 INVX1_88/A CLKBUF1_4/Y NOR2X1_54/Y gnd vdd DFFPOSX1
XFILL_2_0_2 gnd vdd FILL
XNAND3X1_329 NAND2X1_423/Y NAND3X1_327/Y NAND3X1_329/C gnd NAND3X1_334/C vdd NAND3X1
XNAND3X1_318 XNOR2X1_48/Y NAND3X1_318/B NAND3X1_318/C gnd NAND3X1_320/B vdd NAND3X1
XNAND3X1_307 NOR2X1_224/B INVX1_301/A INVX1_300/Y gnd NAND2X1_419/A vdd NAND3X1
XFILL_18_0_2 gnd vdd FILL
XINVX1_140 INVX1_140/A gnd INVX1_140/Y vdd INVX1
XINVX1_184 NOR3X1_5/B gnd INVX1_184/Y vdd INVX1
XINVX1_173 INVX1_173/A gnd INVX1_173/Y vdd INVX1
XINVX1_162 OAI22X1_8/D gnd INVX1_162/Y vdd INVX1
XINVX1_195 INVX1_195/A gnd INVX1_195/Y vdd INVX1
XINVX1_151 INVX1_151/A gnd INVX1_151/Y vdd INVX1
XFILL_20_2_0 gnd vdd FILL
XAOI21X1_166 AOI21X1_166/A NAND2X1_400/Y INVX1_294/A gnd OAI22X1_22/C vdd AOI21X1
XAOI21X1_144 NAND3X1_324/B NAND3X1_324/C INVX1_303/Y gnd OAI21X1_371/A vdd AOI21X1
XAOI21X1_155 OAI21X1_380/Y NAND3X1_346/Y XOR2X1_23/Y gnd OAI21X1_383/A vdd AOI21X1
XAOI21X1_133 NAND3X1_234/Y NAND3X1_238/C INVX1_265/A gnd AOI21X1_133/Y vdd AOI21X1
XAOI21X1_122 OAI21X1_306/Y INVX1_257/Y NOR2X1_195/Y gnd AOI21X1_122/Y vdd AOI21X1
XAOI21X1_111 INVX2_33/A INVX1_242/A INVX1_131/A gnd INVX1_260/A vdd AOI21X1
XAOI21X1_100 NAND2X1_274/Y NAND2X1_228/Y INVX1_208/A gnd OAI22X1_19/C vdd AOI21X1
XNAND3X1_137 INVX1_217/A AOI21X1_80/A AOI21X1_80/B gnd NAND3X1_137/Y vdd NAND3X1
XNAND3X1_126 INVX1_216/A NAND3X1_122/Y AOI21X1_87/A gnd AOI21X1_81/A vdd NAND3X1
XNAND3X1_115 INVX1_104/A INVX1_103/A INVX1_105/A gnd INVX1_215/A vdd NAND3X1
XNAND3X1_148 INVX1_209/Y NAND3X1_145/B NAND3X1_145/C gnd NAND3X1_149/C vdd NAND3X1
XNAND3X1_104 AOI22X1_22/C AOI22X1_22/D NAND2X1_236/Y gnd AOI21X1_78/A vdd NAND3X1
XNAND3X1_159 NAND3X1_159/A NAND3X1_159/B NAND3X1_159/C gnd AOI21X1_92/B vdd NAND3X1
XFILL_11_2_0 gnd vdd FILL
XBUFX4_9 start gnd BUFX4_9/Y vdd BUFX4
XNAND2X1_339 gnd gnd gnd INVX1_267/A vdd NAND2X1
XNAND2X1_317 INVX1_264/A NAND3X1_190/B gnd NAND2X1_317/Y vdd NAND2X1
XNAND2X1_306 OAI21X1_290/Y OAI21X1_291/Y gnd NAND2X1_306/Y vdd NAND2X1
XNAND2X1_328 INVX2_33/A INVX1_242/A gnd INVX1_257/A vdd NAND2X1
XNOR2X1_90 INVX1_87/A INVX1_58/Y gnd NOR2X1_90/Y vdd NOR2X1
XNAND3X1_90 INVX1_195/A INVX1_219/A NAND3X1_93/C gnd NAND3X1_92/B vdd NAND3X1
XOAI21X1_108 INVX1_112/A INVX1_111/Y NOR2X1_65/Y gnd NAND3X1_11/B vdd OAI21X1
XOAI21X1_119 INVX2_5/Y AND2X2_13/A BUFX4_9/Y gnd OAI21X1_119/Y vdd OAI21X1
XNAND2X1_103 NOR2X1_64/A INVX1_73/A gnd NAND2X1_103/Y vdd NAND2X1
XBUFX2_6 BUFX2_6/A gnd X0_mag[5] vdd BUFX2
XNAND2X1_125 INVX1_138/A NAND2X1_124/Y gnd NAND2X1_126/B vdd NAND2X1
XNAND2X1_114 AND2X2_38/B BUFX4_11/Y gnd NAND2X1_114/Y vdd NAND2X1
XNAND2X1_1 NOR2X1_1/Y XOR2X1_1/Y gnd NAND3X1_1/B vdd NAND2X1
XNAND2X1_158 AND2X2_22/A INVX1_164/A gnd AOI22X1_7/C vdd NAND2X1
XNAND2X1_169 INVX1_178/A AOI21X1_58/A gnd NAND3X1_60/B vdd NAND2X1
XNAND2X1_147 INVX1_154/Y AND2X2_21/Y gnd AOI21X1_46/A vdd NAND2X1
XNAND2X1_136 gnd gnd gnd INVX1_145/A vdd NAND2X1
XNOR2X1_191 NOR3X1_8/B NOR2X1_191/B gnd NOR2X1_191/Y vdd NOR2X1
XFILL_0_1_0 gnd vdd FILL
XNOR2X1_180 INVX1_237/A INVX1_238/A gnd INVX1_245/A vdd NOR2X1
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XAOI21X1_6 AOI21X1_6/A AOI21X1_6/B AOI21X1_6/C gnd AOI21X1_6/Y vdd AOI21X1
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XXNOR2X1_47 XNOR2X1_47/A INVX1_298/Y gnd XNOR2X1_47/Y vdd XNOR2X1
XXNOR2X1_36 XOR2X1_15/A XOR2X1_15/B gnd XNOR2X1_36/Y vdd XNOR2X1
XFILL_8_2_0 gnd vdd FILL
XXNOR2X1_14 XNOR2X1_14/A INVX2_6/Y gnd XNOR2X1_14/Y vdd XNOR2X1
XXNOR2X1_25 XNOR2X1_25/A XNOR2X1_25/B gnd XOR2X1_9/B vdd XNOR2X1
XBUFX2_13 BUFX2_13/A gnd X1_mag[4] vdd BUFX2
XFILL_16_1_0 gnd vdd FILL
XINVX1_93 INVX2_36/A gnd INVX1_93/Y vdd INVX1
XINVX1_82 INVX1_82/A gnd INVX1_82/Y vdd INVX1
XBUFX2_24 BUFX2_24/A gnd X2_mag[7] vdd BUFX2
XDFFPOSX1_1 INVX2_28/A CLKBUF1_5/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XINVX1_71 INVX1_71/A gnd INVX1_71/Y vdd INVX1
XNOR2X1_4 x3[4] NOR2X1_4/B gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_14 AND2X2_10/Y INVX2_3/Y INVX1_27/Y gnd AOI21X1_14/Y vdd AOI21X1
XAOI21X1_69 NOR3X1_6/A NAND3X1_33/C INVX1_140/Y gnd NOR2X1_131/B vdd AOI21X1
XAOI21X1_58 AOI21X1_58/A NAND3X1_40/Y INVX1_173/A gnd AOI21X1_58/Y vdd AOI21X1
XAOI21X1_36 OR2X2_5/B NOR2X1_77/Y NOR2X1_82/Y gnd AOI21X1_36/Y vdd AOI21X1
XAOI21X1_47 NAND3X1_21/C NAND3X1_21/B INVX1_156/Y gnd OAI22X1_9/B vdd AOI21X1
XAOI21X1_25 INVX2_6/A NOR2X1_86/Y NOR2X1_90/Y gnd INVX1_126/A vdd AOI21X1
XOAI21X1_9 INVX1_15/Y AND2X2_1/A BUFX4_2/Y gnd OAI22X1_1/D vdd OAI21X1
XOAI22X1_22 OAI22X1_22/A OAI22X1_22/B OAI22X1_22/C OAI22X1_22/D gnd OAI22X1_22/Y vdd
+ OAI22X1
XOAI22X1_11 INVX2_13/A INVX1_151/A XOR2X1_7/B INVX1_170/A gnd INVX1_172/A vdd OAI22X1
XFILL_5_0_0 gnd vdd FILL
XINVX1_300 INVX1_300/A gnd INVX1_300/Y vdd INVX1
XOAI21X1_291 INVX2_29/Y INVX2_33/Y NOR2X1_186/Y gnd OAI21X1_291/Y vdd OAI21X1
XOAI21X1_280 NOR2X1_172/A AOI22X1_28/B INVX1_229/Y gnd NAND3X1_178/A vdd OAI21X1
XINVX1_311 INVX1_311/A gnd INVX1_311/Y vdd INVX1
XDFFPOSX1_47 AND2X2_45/B CLKBUF1_7/Y OAI21X1_87/Y gnd vdd DFFPOSX1
XDFFPOSX1_69 INVX1_75/A CLKBUF1_1/Y OAI22X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_36 INVX1_96/A CLKBUF1_4/Y OAI21X1_94/Y gnd vdd DFFPOSX1
XDFFPOSX1_14 INVX1_106/A CLKBUF1_10/Y DFFPOSX1_14/D gnd vdd DFFPOSX1
XDFFPOSX1_58 INVX1_54/A CLKBUF1_5/Y NOR2X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_25 INVX2_9/A CLKBUF1_9/Y OAI21X1_117/Y gnd vdd DFFPOSX1
XNAND3X1_319 XNOR2X1_47/Y AOI21X1_150/A AOI21X1_150/B gnd NAND3X1_320/C vdd NAND3X1
XNAND3X1_308 NAND3X1_308/A NAND3X1_302/Y AOI21X1_157/A gnd NAND3X1_318/B vdd NAND3X1
XINVX1_141 INVX1_141/A gnd INVX1_141/Y vdd INVX1
XINVX1_130 NOR2X1_96/B gnd INVX1_130/Y vdd INVX1
XINVX1_152 INVX1_152/A gnd INVX1_152/Y vdd INVX1
XINVX1_185 INVX1_185/A gnd INVX1_185/Y vdd INVX1
XINVX1_163 INVX1_163/A gnd INVX1_163/Y vdd INVX1
XINVX1_174 INVX1_174/A gnd INVX1_174/Y vdd INVX1
XINVX1_196 INVX1_196/A gnd INVX1_196/Y vdd INVX1
XFILL_20_2_1 gnd vdd FILL
XAOI21X1_134 AOI21X1_134/A INVX1_284/A INVX1_272/Y gnd NOR2X1_208/A vdd AOI21X1
XAOI21X1_145 NAND3X1_327/B NAND3X1_327/C INVX1_303/A gnd OAI21X1_371/B vdd AOI21X1
XAOI21X1_156 NAND3X1_310/C NAND3X1_304/Y AOI22X1_51/Y gnd AOI21X1_156/Y vdd AOI21X1
XAOI21X1_123 NAND3X1_202/Y NAND3X1_201/Y INVX1_259/A gnd OAI21X1_321/B vdd AOI21X1
XAOI21X1_112 NAND3X1_224/B NAND3X1_224/C INVX1_263/Y gnd OAI21X1_312/A vdd AOI21X1
XAOI21X1_101 OR2X2_21/Y AOI21X1_101/B AND2X2_33/Y gnd NOR2X1_173/A vdd AOI21X1
XNAND3X1_116 NOR2X1_159/B INVX1_215/A INVX1_214/Y gnd NAND2X1_247/A vdd NAND3X1
XNAND3X1_127 XNOR2X1_33/Y NAND3X1_127/B NAND3X1_127/C gnd NAND3X1_132/B vdd NAND3X1
XNAND3X1_138 NAND2X1_251/Y NAND3X1_136/Y NAND3X1_137/Y gnd AOI21X1_85/B vdd NAND3X1
XNAND3X1_105 INVX2_24/Y AOI21X1_78/B AOI21X1_78/A gnd NAND3X1_105/Y vdd NAND3X1
XNAND3X1_149 AOI21X1_82/Y NAND3X1_149/B NAND3X1_149/C gnd AOI22X1_27/C vdd NAND3X1
XFILL_11_2_1 gnd vdd FILL
XNAND2X1_318 NAND2X1_318/A INVX1_246/Y gnd INVX1_247/A vdd NAND2X1
XNAND2X1_307 NAND2X1_307/A NAND2X1_307/B gnd NAND2X1_307/Y vdd NAND2X1
XNAND2X1_329 INVX2_28/A AND2X2_38/B gnd INVX1_256/A vdd NAND2X1
XNAND3X1_80 INVX1_186/Y INVX1_198/A NAND3X1_80/C gnd INVX1_191/A vdd NAND3X1
XNAND3X1_91 INVX1_195/Y NAND3X1_91/B NAND3X1_91/C gnd NAND3X1_92/C vdd NAND3X1
XNOR2X1_80 INVX1_84/A INVX1_55/Y gnd NOR2X1_80/Y vdd NOR2X1
XNOR2X1_91 INVX1_58/A INVX1_87/Y gnd NOR2X1_91/Y vdd NOR2X1
XOAI21X1_109 INVX1_112/Y INVX1_111/A NAND3X1_11/B gnd AOI21X1_17/C vdd OAI21X1
XBUFX2_7 BUFX2_7/A gnd X0_mag[6] vdd BUFX2
XFILL_11_1 gnd vdd FILL
XNAND2X1_104 INVX1_112/A INVX1_111/A gnd OAI21X1_144/C vdd NAND2X1
XNAND2X1_126 NAND3X1_14/Y NAND2X1_126/B gnd OR2X2_9/A vdd NAND2X1
XNAND2X1_159 INVX1_163/Y NOR2X1_119/Y gnd AOI22X1_8/A vdd NAND2X1
XNAND2X1_148 INVX1_154/A NAND2X1_145/Y gnd AOI21X1_46/B vdd NAND2X1
XNAND2X1_115 INVX1_57/A INVX1_86/A gnd NOR2X1_98/A vdd NAND2X1
XNAND2X1_137 gnd gnd gnd INVX1_146/A vdd NAND2X1
XNAND2X1_2 x3[2] INVX1_6/Y gnd NAND2X1_4/A vdd NAND2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XFILL_0_1_1 gnd vdd FILL
XNOR2X1_192 AND2X2_37/Y INVX1_253/Y gnd NOR2X1_192/Y vdd NOR2X1
XNOR2X1_181 INVX1_237/Y INVX1_238/Y gnd NOR2X1_181/Y vdd NOR2X1
XNOR2X1_170 INVX2_30/Y INVX2_31/Y gnd NOR2X1_170/Y vdd NOR2X1
XAOI21X1_7 INVX1_40/A AOI21X1_7/B NOR2X1_41/Y gnd AOI21X1_7/Y vdd AOI21X1
XINVX1_61 x0[5] gnd INVX1_61/Y vdd INVX1
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XXNOR2X1_48 XNOR2X1_47/A INVX1_298/A gnd XNOR2X1_48/Y vdd XNOR2X1
XXNOR2X1_37 AOI21X1_94/Y INVX1_225/A gnd XNOR2X1_37/Y vdd XNOR2X1
XXNOR2X1_26 INVX2_13/A XOR2X1_10/B gnd XOR2X1_8/B vdd XNOR2X1
XFILL_8_2_1 gnd vdd FILL
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XINVX1_94 INVX2_37/A gnd INVX1_94/Y vdd INVX1
XXNOR2X1_15 XNOR2X1_15/A INVX2_5/Y gnd XNOR2X1_15/Y vdd XNOR2X1
XFILL_16_1_1 gnd vdd FILL
XBUFX2_14 BUFX2_14/A gnd X1_mag[5] vdd BUFX2
XBUFX2_25 BUFX2_25/A gnd X3_mag[0] vdd BUFX2
XDFFPOSX1_2 INVX2_29/A CLKBUF1_5/Y DFFPOSX1_2/D gnd vdd DFFPOSX1
XNOR2X1_5 NOR2X1_3/Y NOR2X1_4/Y gnd NOR2X1_5/Y vdd NOR2X1
XAOI21X1_15 NOR2X1_62/Y INVX2_4/Y INVX1_29/Y gnd OAI21X1_87/A vdd AOI21X1
XAOI21X1_59 NAND3X1_54/B NAND3X1_54/C AOI22X1_6/A gnd AOI21X1_60/C vdd AOI21X1
XAOI21X1_48 AOI21X1_45/A AOI21X1_45/B INVX1_155/Y gnd OAI22X1_8/D vdd AOI21X1
XAOI21X1_37 NOR2X1_96/B NOR2X1_97/Y AOI21X1_37/C gnd AND2X2_16/A vdd AOI21X1
XAOI21X1_26 NOR2X1_89/B INVX1_125/Y INVX1_126/Y gnd AOI21X1_26/Y vdd AOI21X1
XOAI22X1_12 OAI22X1_14/A OAI22X1_14/B OAI22X1_15/C NOR3X1_3/Y gnd NAND3X1_44/B vdd
+ OAI22X1
XFILL_5_0_1 gnd vdd FILL
XINVX1_301 INVX1_301/A gnd INVX1_301/Y vdd INVX1
XOAI21X1_270 NAND2X1_251/Y AOI21X1_81/Y NAND3X1_130/Y gnd NAND2X1_271/B vdd OAI21X1
XOAI21X1_292 INVX2_34/Y INVX1_241/Y NAND2X1_306/Y gnd NAND2X1_307/A vdd OAI21X1
XOAI21X1_281 INVX2_30/Y INVX2_31/Y NAND2X1_281/Y gnd NAND2X1_282/B vdd OAI21X1
XDFFPOSX1_48 INVX1_92/A CLKBUF1_4/Y OAI21X1_90/Y gnd vdd DFFPOSX1
XDFFPOSX1_37 INVX1_97/A CLKBUF1_4/Y OAI21X1_95/Y gnd vdd DFFPOSX1
XDFFPOSX1_26 INVX2_10/A CLKBUF1_9/Y OAI21X1_120/Y gnd vdd DFFPOSX1
XDFFPOSX1_59 INVX1_55/A CLKBUF1_5/Y NOR2X1_35/Y gnd vdd DFFPOSX1
XDFFPOSX1_15 INVX1_107/A CLKBUF1_10/Y DFFPOSX1_15/D gnd vdd DFFPOSX1
XNAND3X1_309 AOI22X1_51/Y AOI21X1_152/B AOI21X1_152/A gnd NAND3X1_309/Y vdd NAND3X1
XINVX1_186 INVX1_186/A gnd INVX1_186/Y vdd INVX1
XINVX1_142 gnd gnd INVX1_142/Y vdd INVX1
XINVX1_164 INVX1_164/A gnd INVX1_164/Y vdd INVX1
XINVX1_175 INVX1_175/A gnd INVX1_175/Y vdd INVX1
XINVX1_131 INVX1_131/A gnd INVX1_131/Y vdd INVX1
XINVX1_120 OR2X2_5/B gnd INVX1_120/Y vdd INVX1
XINVX1_153 INVX1_153/A gnd INVX1_153/Y vdd INVX1
XINVX1_197 INVX1_197/A gnd INVX1_197/Y vdd INVX1
XAOI21X1_146 INVX1_281/A NAND3X1_281/C INVX1_305/Y gnd AOI21X1_146/Y vdd AOI21X1
XAOI21X1_135 NAND2X1_380/Y NAND3X1_275/B INVX1_283/Y gnd NOR2X1_219/A vdd AOI21X1
XFILL_20_2_2 gnd vdd FILL
XAOI21X1_157 AOI21X1_157/A NAND3X1_308/A AOI21X1_156/Y gnd XOR2X1_24/A vdd AOI21X1
XAOI21X1_102 NAND2X1_295/Y NAND2X1_294/Y INVX1_235/Y gnd OAI21X1_285/B vdd AOI21X1
XAOI21X1_124 NAND3X1_215/Y NAND3X1_214/Y XNOR2X1_40/Y gnd AOI21X1_125/C vdd AOI21X1
XAOI21X1_113 NAND3X1_217/Y NAND3X1_221/C INVX1_263/A gnd OAI21X1_312/B vdd AOI21X1
XNAND3X1_128 XNOR2X1_32/Y AOI21X1_86/A AOI21X1_86/B gnd NAND3X1_132/C vdd NAND3X1
XNAND3X1_117 NAND2X1_247/Y NAND3X1_111/Y NAND3X1_114/Y gnd NAND3X1_127/B vdd NAND3X1
XNAND3X1_139 AOI21X1_85/C AOI21X1_85/A AOI21X1_85/B gnd NAND3X1_142/B vdd NAND3X1
XNAND3X1_106 OAI21X1_248/Y INVX1_211/Y NAND3X1_105/Y gnd NAND2X1_238/A vdd NAND3X1
XFILL_11_2_2 gnd vdd FILL
XNAND2X1_308 INVX1_240/A NAND2X1_307/Y gnd AOI22X1_31/A vdd NAND2X1
XNAND2X1_319 gnd gnd gnd OR2X2_25/A vdd NAND2X1
XNAND3X1_92 AOI21X1_76/Y NAND3X1_92/B NAND3X1_92/C gnd NAND3X1_92/Y vdd NAND3X1
XNAND3X1_70 AOI21X1_66/A AOI21X1_66/B NAND3X1_69/Y gnd NAND3X1_70/Y vdd NAND3X1
XNAND3X1_81 INVX2_19/Y INVX1_103/A INVX1_192/Y gnd NAND3X1_82/C vdd NAND3X1
XNOR2X1_81 INVX1_56/A INVX1_85/A gnd NOR2X1_81/Y vdd NOR2X1
XFILL_11_2 gnd vdd FILL
XNOR2X1_70 NOR2X1_70/A NOR2X1_70/B gnd NOR2X1_70/Y vdd NOR2X1
XNOR2X1_92 NOR2X1_90/Y NOR2X1_91/Y gnd INVX2_6/A vdd NOR2X1
XBUFX2_8 BUFX2_8/A gnd X0_mag[7] vdd BUFX2
XNAND2X1_3 x1[2] INVX1_7/Y gnd INVX1_9/A vdd NAND2X1
XNAND2X1_105 INVX1_41/A INVX1_75/A gnd OAI21X1_145/A vdd NAND2X1
XNAND2X1_149 AOI21X1_67/B NAND3X1_32/Y gnd XNOR2X1_22/A vdd NAND2X1
XNAND2X1_127 OR2X2_9/B OR2X2_9/A gnd NAND3X1_15/B vdd NAND2X1
XNAND2X1_116 gnd INVX2_8/Y gnd XNOR2X1_18/B vdd NAND2X1
XNAND2X1_138 INVX1_148/Y NOR2X1_116/Y gnd NAND3X1_21/C vdd NAND2X1
XFILL_0_1_2 gnd vdd FILL
XNOR2X1_160 OR2X2_20/B OR2X2_20/A gnd NOR2X1_160/Y vdd NOR2X1
XAOI21X1_8 INVX1_64/Y x0[7] BUFX4_14/Y gnd AOI21X1_8/Y vdd AOI21X1
XNOR2X1_193 NOR2X1_191/Y NOR2X1_192/Y gnd NOR2X1_193/Y vdd NOR2X1
XINVX2_8 gnd gnd INVX2_8/Y vdd INVX2
XNOR2X1_182 INVX1_245/A NOR2X1_181/Y gnd OR2X2_23/A vdd NOR2X1
XNOR2X1_171 INVX2_29/Y INVX2_33/Y gnd AOI22X1_28/B vdd NOR2X1
XINVX1_62 INVX1_62/A gnd AND2X2_7/B vdd INVX1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XINVX1_40 INVX1_40/A gnd AND2X2_2/A vdd INVX1
XINVX1_73 INVX1_73/A gnd INVX1_73/Y vdd INVX1
XXNOR2X1_49 XNOR2X1_49/A OAI22X1_21/Y gnd INVX1_302/A vdd XNOR2X1
XBUFX2_15 BUFX2_15/A gnd X1_mag[6] vdd BUFX2
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XBUFX2_26 BUFX2_26/A gnd X3_mag[1] vdd BUFX2
XXNOR2X1_38 INVX2_30/A XNOR2X1_38/B gnd XNOR2X1_38/Y vdd XNOR2X1
XXNOR2X1_27 XOR2X1_9/B XOR2X1_8/B gnd XNOR2X1_27/Y vdd XNOR2X1
XFILL_8_2_2 gnd vdd FILL
XXNOR2X1_16 XNOR2X1_16/A NOR2X1_85/A gnd XNOR2X1_16/Y vdd XNOR2X1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XFILL_16_1_2 gnd vdd FILL
XDFFPOSX1_3 INVX2_33/A CLKBUF1_9/Y DFFPOSX1_3/D gnd vdd DFFPOSX1
XNOR2X1_6 INVX1_8/A XOR2X1_2/B gnd NOR2X1_6/Y vdd NOR2X1
XAOI21X1_16 NAND2X1_65/B NAND2X1_65/A NAND2X1_68/Y gnd AOI21X1_17/A vdd AOI21X1
XAOI21X1_49 AOI21X1_46/A AOI21X1_46/B INVX1_155/A gnd OAI22X1_8/C vdd AOI21X1
XAOI21X1_27 NOR2X1_94/B INVX2_7/A INVX1_124/A gnd AOI21X1_27/Y vdd AOI21X1
XAOI21X1_38 INVX1_58/A INVX1_87/A NOR2X1_98/Y gnd AOI21X1_38/Y vdd AOI21X1
XOAI22X1_13 NOR3X1_5/A AOI21X1_58/Y OAI22X1_13/C NOR3X1_4/Y gnd NAND3X1_44/C vdd OAI22X1
XOAI21X1_90 INVX1_30/A OR2X2_4/Y OAI21X1_89/Y gnd OAI21X1_90/Y vdd OAI21X1
XFILL_5_0_2 gnd vdd FILL
XINVX1_302 INVX1_302/A gnd INVX1_302/Y vdd INVX1
XOAI21X1_271 AOI21X1_95/Y INVX1_224/Y NAND3X1_168/C gnd AOI21X1_98/B vdd OAI21X1
XOAI21X1_293 AOI22X1_29/Y AOI22X1_30/Y OAI21X1_286/Y gnd INVX1_264/A vdd OAI21X1
XOAI21X1_282 OR2X2_21/B OR2X2_21/A NAND3X1_178/Y gnd INVX1_235/A vdd OAI21X1
XOAI21X1_260 NAND3X1_99/B NOR2X1_159/A XOR2X1_16/B gnd AOI21X1_88/A vdd OAI21X1
XDFFPOSX1_27 INVX1_139/A CLKBUF1_3/Y OAI21X1_123/Y gnd vdd DFFPOSX1
XDFFPOSX1_16 INVX1_108/A CLKBUF1_10/Y DFFPOSX1_16/D gnd vdd DFFPOSX1
XDFFPOSX1_49 INVX1_31/A CLKBUF1_2/Y OAI21X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_38 INVX1_98/A CLKBUF1_4/Y OAI21X1_96/Y gnd vdd DFFPOSX1
XFILL_23_2_0 gnd vdd FILL
XFILL_14_2_0 gnd vdd FILL
XINVX1_110 INVX1_110/A gnd INVX1_110/Y vdd INVX1
XINVX1_198 INVX1_198/A gnd INVX1_198/Y vdd INVX1
XINVX1_143 INVX1_143/A gnd INVX1_143/Y vdd INVX1
XINVX1_165 NOR3X1_2/A gnd INVX1_165/Y vdd INVX1
XINVX1_176 XOR2X1_10/A gnd INVX1_176/Y vdd INVX1
XINVX1_154 INVX1_154/A gnd INVX1_154/Y vdd INVX1
XINVX1_121 INVX1_121/A gnd INVX1_121/Y vdd INVX1
XINVX1_132 INVX1_132/A gnd INVX1_132/Y vdd INVX1
XINVX1_187 INVX1_187/A gnd INVX1_187/Y vdd INVX1
XAOI21X1_114 INVX1_234/A NAND3X1_191/B INVX1_264/Y gnd AOI21X1_114/Y vdd AOI21X1
XAOI21X1_103 NAND3X1_182/C NAND3X1_182/B INVX1_235/A gnd AOI21X1_103/Y vdd AOI21X1
XAOI21X1_136 NAND2X1_376/Y NAND2X1_379/Y INVX1_283/A gnd NOR2X1_219/B vdd AOI21X1
XAOI21X1_147 NAND3X1_343/Y NAND3X1_342/Y INVX1_306/Y gnd AOI21X1_147/Y vdd AOI21X1
XAOI21X1_158 NAND2X1_436/A NAND2X1_436/B XOR2X1_24/Y gnd AOI21X1_158/Y vdd AOI21X1
XAOI21X1_125 NAND3X1_216/Y INVX1_262/Y AOI21X1_125/C gnd AOI21X1_125/Y vdd AOI21X1
XNAND3X1_118 AOI22X1_25/Y AOI21X1_91/B AOI21X1_91/A gnd NAND3X1_118/Y vdd NAND3X1
XNAND3X1_129 INVX1_216/Y NAND3X1_132/B NAND3X1_132/C gnd AOI21X1_81/B vdd NAND3X1
XNAND3X1_107 INVX2_26/Y AOI21X1_89/A NAND2X1_244/Y gnd AOI21X1_91/A vdd NAND3X1
XNAND2X1_309 INVX1_236/Y INVX1_239/A gnd AOI22X1_31/C vdd NAND2X1
XFILL_20_0_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XNOR2X1_60 INVX1_24/A INVX2_2/A gnd NOR2X1_60/Y vdd NOR2X1
XFILL_19_1_0 gnd vdd FILL
XNOR2X1_71 NOR2X1_71/A NOR2X1_71/B gnd NOR2X1_71/Y vdd NOR2X1
XNAND3X1_60 NAND3X1_55/Y NAND3X1_60/B NAND3X1_56/C gnd NAND3X1_60/Y vdd NAND3X1
XNAND3X1_71 NAND3X1_43/Y NAND3X1_71/B NAND3X1_71/C gnd NAND3X1_71/Y vdd NAND3X1
XNOR2X1_82 INVX1_56/Y INVX1_85/Y gnd NOR2X1_82/Y vdd NOR2X1
XNAND3X1_82 NAND3X1_82/A NOR2X1_142/Y NAND3X1_82/C gnd NAND3X1_82/Y vdd NAND3X1
XNAND3X1_93 INVX1_195/Y INVX1_219/A NAND3X1_93/C gnd NAND3X1_95/B vdd NAND3X1
XNOR2X1_93 INVX1_88/A INVX1_59/Y gnd INVX1_124/A vdd NOR2X1
XFILL_11_3 gnd vdd FILL
XBUFX2_9 BUFX2_9/A gnd X1_mag[0] vdd BUFX2
XNAND2X1_4 NAND2X1_4/A INVX1_9/A gnd INVX1_8/A vdd NAND2X1
XNAND2X1_106 INVX1_114/A INVX1_113/A gnd NAND2X1_106/Y vdd NAND2X1
XNAND2X1_117 gnd gnd gnd INVX1_136/A vdd NAND2X1
XNAND2X1_128 INVX2_9/A INVX1_153/A gnd XOR2X1_6/B vdd NAND2X1
XNAND2X1_139 INVX1_139/A INVX1_152/A gnd INVX2_13/A vdd NAND2X1
XNOR2X1_161 INVX1_191/Y NOR2X1_161/B gnd NOR2X1_161/Y vdd NOR2X1
XNOR2X1_194 OR2X2_24/B OR2X2_24/A gnd NOR2X1_194/Y vdd NOR2X1
XNOR2X1_183 NOR2X1_183/A NOR2X1_183/B gnd NOR2X1_183/Y vdd NOR2X1
XNOR2X1_172 NOR2X1_172/A AOI22X1_28/B gnd NOR2X1_172/Y vdd NOR2X1
XNOR2X1_150 INVX2_18/Y INVX1_204/Y gnd NOR2X1_150/Y vdd NOR2X1
XAOI21X1_9 AOI21X1_9/A INVX1_8/A NOR2X1_42/Y gnd XOR2X1_2/A vdd AOI21X1
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XXNOR2X1_39 XNOR2X1_39/A INVX1_256/Y gnd XNOR2X1_39/Y vdd XNOR2X1
XXNOR2X1_28 XOR2X1_9/A XOR2X1_9/B gnd XNOR2X1_28/Y vdd XNOR2X1
XXNOR2X1_17 XNOR2X1_17/A INVX2_6/Y gnd XNOR2X1_17/Y vdd XNOR2X1
XINVX1_74 x3[1] gnd INVX1_74/Y vdd INVX1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XBUFX2_16 BUFX2_16/A gnd X1_mag[7] vdd BUFX2
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XBUFX2_27 BUFX2_27/A gnd X3_mag[2] vdd BUFX2
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XDFFPOSX1_4 INVX1_131/A CLKBUF1_9/Y AOI22X1_4/Y gnd vdd DFFPOSX1
XNOR2X1_7 x1[5] INVX1_18/Y gnd NOR2X1_9/A vdd NOR2X1
XNAND3X1_290 INVX2_43/Y OAI21X1_362/C OR2X2_32/Y gnd AOI22X1_48/A vdd NAND3X1
XAOI21X1_17 AOI21X1_17/A AOI21X1_17/B AOI21X1_17/C gnd AOI21X1_17/Y vdd AOI21X1
XAOI21X1_39 AND2X2_17/A INVX2_7/Y NOR2X1_100/Y gnd AOI21X1_40/A vdd AOI21X1
XAOI21X1_28 AOI21X1_27/Y INVX1_128/Y BUFX4_10/Y gnd AOI22X1_3/D vdd AOI21X1
XOAI22X1_14 OAI22X1_14/A OAI22X1_14/B OAI22X1_13/C NOR3X1_4/Y gnd NAND3X1_42/B vdd
+ OAI22X1
XFILL_8_0_0 gnd vdd FILL
XOAI21X1_80 INVX1_91/A NOR2X1_58/B BUFX4_6/Y gnd OAI21X1_80/Y vdd OAI21X1
XOAI21X1_91 BUFX4_7/Y INVX1_93/Y OAI21X1_91/C gnd OAI21X1_91/Y vdd OAI21X1
XOAI21X1_250 INVX2_18/Y INVX1_213/Y NOR2X1_159/B gnd AOI21X1_89/A vdd OAI21X1
XINVX1_303 INVX1_303/A gnd INVX1_303/Y vdd INVX1
XOAI21X1_272 AOI21X1_95/Y INVX1_224/Y XNOR2X1_37/Y gnd AOI21X1_99/A vdd OAI21X1
XOAI21X1_294 OR2X2_24/A AOI22X1_32/Y AOI21X1_106/Y gnd NAND3X1_191/B vdd OAI21X1
XOAI21X1_261 AOI21X1_88/Y NOR2X1_157/Y INVX1_221/A gnd NAND3X1_157/C vdd OAI21X1
XOAI21X1_283 INVX2_29/A INVX2_33/Y NOR2X1_183/A gnd OAI21X1_283/Y vdd OAI21X1
XDFFPOSX1_39 INVX1_99/A CLKBUF1_8/Y OAI21X1_97/Y gnd vdd DFFPOSX1
XDFFPOSX1_17 INVX2_17/A CLKBUF1_10/Y DFFPOSX1_17/D gnd vdd DFFPOSX1
XDFFPOSX1_28 INVX1_153/A CLKBUF1_9/Y AOI22X1_2/Y gnd vdd DFFPOSX1
XFILL_23_2_1 gnd vdd FILL
XFILL_14_2_1 gnd vdd FILL
XINVX1_100 INVX1_100/A gnd INVX1_100/Y vdd INVX1
XINVX1_111 INVX1_111/A gnd INVX1_111/Y vdd INVX1
XINVX1_133 reset gnd DFFSR_1/R vdd INVX1
XINVX1_144 gnd gnd INVX1_144/Y vdd INVX1
XINVX1_177 OR2X2_14/A gnd INVX1_177/Y vdd INVX1
XINVX1_166 NOR3X1_2/C gnd AOI22X1_9/C vdd INVX1
XINVX1_155 INVX1_155/A gnd INVX1_155/Y vdd INVX1
XINVX1_199 INVX1_199/A gnd OR2X2_18/B vdd INVX1
XINVX1_122 INVX1_122/A gnd INVX1_122/Y vdd INVX1
XINVX1_188 INVX1_188/A gnd INVX1_188/Y vdd INVX1
XAOI21X1_137 OAI21X1_344/Y NAND3X1_276/Y INVX1_277/A gnd XOR2X1_21/B vdd AOI21X1
XAOI21X1_148 NAND2X1_424/B XNOR2X1_50/B AOI21X1_147/Y gnd NAND3X1_362/A vdd AOI21X1
XAOI21X1_115 NAND3X1_239/Y AOI21X1_115/B INVX1_265/Y gnd AOI21X1_115/Y vdd AOI21X1
XAOI21X1_126 AOI21X1_126/A AOI21X1_126/B INVX1_271/A gnd NOR3X1_11/C vdd AOI21X1
XAOI21X1_104 NAND2X1_361/B NAND3X1_184/Y INVX1_231/A gnd XOR2X1_18/B vdd AOI21X1
XAOI21X1_159 OR2X2_33/Y NAND3X1_353/B NAND3X1_353/C gnd OAI21X1_385/B vdd AOI21X1
XNAND3X1_119 OAI22X1_18/Y NAND3X1_113/Y NAND3X1_112/Y gnd NAND3X1_119/Y vdd NAND3X1
XNAND3X1_108 INVX2_18/A INVX1_107/A NOR2X1_159/B gnd NAND3X1_108/Y vdd NAND3X1
XFILL_20_0_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XNAND3X1_50 INVX1_175/Y NAND3X1_48/Y NAND3X1_49/Y gnd NAND3X1_50/Y vdd NAND3X1
XFILL_19_1_1 gnd vdd FILL
XNOR2X1_61 INVX2_3/A INVX1_27/A gnd NOR2X1_61/Y vdd NOR2X1
XNAND3X1_72 INVX1_185/Y NAND3X1_70/Y NAND3X1_71/Y gnd NAND3X1_72/Y vdd NAND3X1
XNAND3X1_61 NAND3X1_61/A NAND3X1_60/Y AOI21X1_63/C gnd NAND3X1_61/Y vdd NAND3X1
XNOR2X1_83 NOR2X1_81/Y NOR2X1_82/Y gnd OR2X2_5/B vdd NOR2X1
XNOR2X1_50 BUFX4_9/Y INVX1_84/Y gnd NOR2X1_50/Y vdd NOR2X1
XNAND3X1_94 INVX1_195/A NAND3X1_91/B NAND3X1_91/C gnd NAND3X1_95/C vdd NAND3X1
XNOR2X1_72 INVX1_54/A INVX1_83/A gnd NOR2X1_74/A vdd NOR2X1
XNOR2X1_94 INVX2_7/A NOR2X1_94/B gnd NOR2X1_94/Y vdd NOR2X1
XNAND3X1_83 INVX1_197/A AOI21X1_72/B AOI21X1_72/A gnd NAND3X1_85/B vdd NAND3X1
XNAND2X1_107 INVX2_28/A BUFX4_13/Y gnd NAND2X1_107/Y vdd NAND2X1
XNAND2X1_5 INVX1_89/A BUFX4_15/Y gnd NAND2X1_5/Y vdd NAND2X1
XNAND2X1_118 gnd NOR2X1_104/Y gnd AOI21X1_41/B vdd NAND2X1
XNAND2X1_129 INVX1_139/A INVX2_10/Y gnd XOR2X1_6/A vdd NAND2X1
XNOR2X1_162 XOR2X1_13/B NOR2X1_161/Y gnd NOR2X1_162/Y vdd NOR2X1
XNOR2X1_173 NOR2X1_173/A INVX1_230/Y gnd NOR2X1_173/Y vdd NOR2X1
XNOR2X1_195 NOR2X1_191/B NOR2X1_195/B gnd NOR2X1_195/Y vdd NOR2X1
XNOR2X1_184 INVX1_241/Y INVX2_34/Y gnd NOR2X1_184/Y vdd NOR2X1
XNOR2X1_151 INVX1_205/Y NOR2X1_150/Y gnd NOR2X1_151/Y vdd NOR2X1
XNOR2X1_140 NOR2X1_140/A NOR2X1_140/B gnd AOI22X1_16/D vdd NOR2X1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XXNOR2X1_18 NOR2X1_104/Y XNOR2X1_18/B gnd XNOR2X1_18/Y vdd XNOR2X1
XXNOR2X1_29 XOR2X1_10/Y INVX2_13/Y gnd INVX1_179/A vdd XNOR2X1
XINVX1_64 x2[7] gnd INVX1_64/Y vdd INVX1
XINVX1_53 INVX1_53/A gnd OR2X2_2/B vdd INVX1
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XBUFX2_28 BUFX2_28/A gnd X3_mag[3] vdd BUFX2
XBUFX2_17 BUFX2_17/A gnd X2_mag[0] vdd BUFX2
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XDFFPOSX1_5 INVX1_242/A CLKBUF1_9/Y DFFPOSX1_5/D gnd vdd DFFPOSX1
XNOR2X1_8 x3[5] INVX1_19/Y gnd NOR2X1_8/Y vdd NOR2X1
XNAND3X1_280 INVX1_288/A NAND3X1_279/B NAND3X1_279/C gnd INVX1_304/A vdd NAND3X1
XNAND3X1_291 INVX2_43/Y INVX1_296/A OR2X2_32/Y gnd AOI22X1_49/D vdd NAND3X1
XAOI21X1_29 AOI21X1_29/A NOR2X1_95/Y AOI21X1_29/C gnd AOI21X1_29/Y vdd AOI21X1
XAOI21X1_18 AOI21X1_18/A NOR2X1_66/Y INVX1_118/A gnd AOI21X1_18/Y vdd AOI21X1
XOAI22X1_15 NOR3X1_5/A AOI21X1_58/Y OAI22X1_15/C NOR3X1_3/Y gnd NAND3X1_42/C vdd OAI22X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_81 OAI21X1_80/Y AOI21X1_14/Y OAI21X1_81/C gnd OAI21X1_81/Y vdd OAI21X1
XOAI21X1_70 BUFX4_3/Y INVX1_78/Y NAND3X1_6/Y gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_92 BUFX4_5/Y INVX1_94/Y NAND2X1_55/Y gnd OAI21X1_92/Y vdd OAI21X1
XOAI21X1_240 INVX1_198/A AOI21X1_72/Y NAND3X1_85/B gnd NAND3X1_97/A vdd OAI21X1
XOAI21X1_251 INVX1_214/A INVX1_215/Y AND2X2_30/Y gnd NAND2X1_247/B vdd OAI21X1
XOAI21X1_262 INVX2_26/A NOR2X1_158/Y NAND2X1_244/Y gnd NAND2X1_258/B vdd OAI21X1
XOAI21X1_273 INVX1_207/Y NAND3X1_86/Y OR2X2_20/A gnd OAI21X1_273/Y vdd OAI21X1
XINVX1_304 INVX1_304/A gnd INVX1_304/Y vdd INVX1
XOAI21X1_295 AOI22X1_29/Y AOI22X1_30/Y AOI21X1_106/Y gnd NAND3X1_189/B vdd OAI21X1
XOAI21X1_284 INVX2_27/Y INVX1_232/Y NAND2X1_286/Y gnd NAND2X1_287/B vdd OAI21X1
XAND2X2_40 OR2X2_27/Y AND2X2_40/B gnd AND2X2_40/Y vdd AND2X2
XNAND2X1_290 AND2X2_35/Y AND2X2_34/Y gnd NAND3X1_182/C vdd NAND2X1
XDFFPOSX1_18 INVX1_187/A CLKBUF1_8/Y DFFPOSX1_18/D gnd vdd DFFPOSX1
XDFFPOSX1_29 INVX1_152/A CLKBUF1_3/Y OAI21X1_129/Y gnd vdd DFFPOSX1
XFILL_23_2_2 gnd vdd FILL
XFILL_14_2_2 gnd vdd FILL
XINVX1_112 INVX1_112/A gnd INVX1_112/Y vdd INVX1
XINVX1_134 gnd gnd INVX1_134/Y vdd INVX1
XINVX1_123 AND2X2_16/B gnd INVX1_123/Y vdd INVX1
XINVX1_101 INVX2_18/A gnd INVX1_101/Y vdd INVX1
XINVX1_167 NOR3X1_2/B gnd INVX1_167/Y vdd INVX1
XINVX1_178 INVX1_178/A gnd INVX1_178/Y vdd INVX1
XINVX1_189 INVX1_103/A gnd INVX1_189/Y vdd INVX1
XINVX1_145 INVX1_145/A gnd INVX1_145/Y vdd INVX1
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XAOI21X1_138 INVX1_286/Y INVX2_41/A OAI21X1_347/Y gnd OR2X2_30/B vdd AOI21X1
XAOI21X1_149 NAND3X1_334/A NAND3X1_334/C OAI21X1_358/Y gnd AOI21X1_149/Y vdd AOI21X1
XAOI21X1_127 OAI21X1_304/Y INVX1_254/A NOR3X1_9/Y gnd XNOR2X1_44/B vdd AOI21X1
XAOI21X1_116 NAND2X1_338/B XNOR2X1_41/B AOI21X1_115/Y gnd OAI21X1_330/C vdd AOI21X1
XAOI21X1_105 INVX1_237/Y gnd OAI21X1_288/Y gnd OR2X2_23/B vdd AOI21X1
XNAND3X1_109 INVX2_19/A INVX1_106/A NOR2X1_159/A gnd NAND3X1_109/Y vdd NAND3X1
XFILL_20_0_2 gnd vdd FILL
XFILL_3_1_2 gnd vdd FILL
XFILL_11_0_2 gnd vdd FILL
XNAND3X1_51 NOR3X1_6/B INVX1_185/A NAND3X1_50/Y gnd NAND3X1_51/Y vdd NAND3X1
XNAND3X1_73 NAND3X1_72/Y NAND3X1_73/B NAND3X1_73/C gnd NAND3X1_73/Y vdd NAND3X1
XNAND3X1_62 INVX1_183/Y INVX1_184/Y NAND3X1_44/B gnd NAND3X1_62/Y vdd NAND3X1
XNAND3X1_40 NAND3X1_36/A NAND3X1_40/B NAND3X1_37/Y gnd NAND3X1_40/Y vdd NAND3X1
XNAND3X1_84 INVX1_197/Y NAND3X1_84/B NAND3X1_84/C gnd NAND3X1_85/C vdd NAND3X1
XNOR2X1_40 x2[2] INVX1_36/Y gnd AOI21X1_7/B vdd NOR2X1
XNOR2X1_62 INVX1_28/A NOR3X1_1/C gnd NOR2X1_62/Y vdd NOR2X1
XFILL_19_1_2 gnd vdd FILL
XNOR2X1_95 NOR2X1_95/A NOR2X1_95/B gnd NOR2X1_95/Y vdd NOR2X1
XNAND3X1_95 NAND3X1_97/A NAND3X1_95/B NAND3X1_95/C gnd NAND3X1_95/Y vdd NAND3X1
XNOR2X1_84 NOR2X1_80/Y NOR2X1_79/Y gnd NOR2X1_84/Y vdd NOR2X1
XNOR2X1_51 BUFX4_5/Y INVX1_85/Y gnd NOR2X1_51/Y vdd NOR2X1
XNOR2X1_73 INVX1_54/Y INVX1_83/Y gnd NOR2X1_73/Y vdd NOR2X1
XNAND2X1_108 INVX1_116/A INVX1_80/A gnd OAI21X1_146/C vdd NAND2X1
XNAND2X1_119 INVX1_136/Y NOR2X1_104/Y gnd OR2X2_8/B vdd NAND2X1
XNAND2X1_6 x3[3] INVX1_10/Y gnd INVX1_16/A vdd NAND2X1
XNOR2X1_141 AOI21X1_70/Y INVX1_191/Y gnd NOR2X1_141/Y vdd NOR2X1
XNOR2X1_174 INVX1_226/Y NOR2X1_173/Y gnd NOR2X1_175/A vdd NOR2X1
XNOR2X1_130 AOI22X1_14/Y AOI21X1_63/Y gnd NOR2X1_130/Y vdd NOR2X1
XNOR2X1_196 AND2X2_37/Y AND2X2_38/Y gnd NOR2X1_196/Y vdd NOR2X1
XNOR2X1_185 INVX2_28/Y INVX1_242/Y gnd NOR2X1_185/Y vdd NOR2X1
XNOR2X1_163 INVX2_27/Y INVX2_28/Y gnd NOR2X1_163/Y vdd NOR2X1
XNOR2X1_152 AOI21X1_76/C AOI21X1_72/Y gnd AND2X2_27/A vdd NOR2X1
XINVX1_43 x0[4] gnd INVX1_43/Y vdd INVX1
XINVX1_21 x3[6] gnd INVX1_21/Y vdd INVX1
XINVX1_32 x0[0] gnd INVX1_32/Y vdd INVX1
XINVX1_10 x1[3] gnd INVX1_10/Y vdd INVX1
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XXNOR2X1_19 XOR2X1_6/A XOR2X1_6/B gnd XNOR2X1_19/Y vdd XNOR2X1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XBUFX2_29 BUFX2_29/A gnd X3_mag[4] vdd BUFX2
XBUFX2_18 BUFX2_18/A gnd X2_mag[1] vdd BUFX2
XDFFPOSX1_6 AND2X2_38/B CLKBUF1_5/Y DFFPOSX1_6/D gnd vdd DFFPOSX1
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XNOR2X1_9 NOR2X1_9/A NOR2X1_8/Y gnd NOR2X1_9/Y vdd NOR2X1
XNAND3X1_281 INVX1_281/A INVX1_305/A NAND3X1_281/C gnd NAND3X1_281/Y vdd NAND3X1
XNAND3X1_292 AOI22X1_49/C AOI22X1_49/D NAND3X1_292/C gnd OAI21X1_374/C vdd NAND3X1
XNAND3X1_270 AND2X2_43/Y NAND3X1_270/B OR2X2_28/Y gnd INVX1_284/A vdd NAND3X1
XAOI21X1_19 NOR2X1_71/Y AOI21X1_19/B AOI21X1_19/C gnd AOI21X1_19/Y vdd AOI21X1
XOAI22X1_16 NOR3X1_2/C NOR2X1_123/Y OAI22X1_16/C NOR2X1_124/Y gnd NAND3X1_57/B vdd
+ OAI22X1
XFILL_8_0_2 gnd vdd FILL
XFILL_8_1 gnd vdd FILL
XOAI21X1_82 INVX1_28/A NOR3X1_1/C BUFX4_8/Y gnd OAI21X1_82/Y vdd OAI21X1
XOAI21X1_60 INVX1_5/Y INVX1_74/Y NAND3X1_4/B gnd AOI21X1_9/A vdd OAI21X1
XOAI21X1_71 INVX2_1/Y INVX1_21/Y NAND3X1_6/B gnd OAI21X1_72/B vdd OAI21X1
XOAI21X1_93 BUFX4_1/Y INVX1_95/Y OAI21X1_93/C gnd OAI21X1_93/Y vdd OAI21X1
XFILL_1_2_0 gnd vdd FILL
XINVX1_305 INVX1_305/A gnd INVX1_305/Y vdd INVX1
XOAI21X1_296 OR2X2_24/A AOI22X1_32/Y OAI21X1_286/Y gnd NAND3X1_189/C vdd OAI21X1
XOAI21X1_252 INVX1_214/A INVX1_215/Y NOR2X1_159/B gnd NAND2X1_248/B vdd OAI21X1
XOAI21X1_285 AOI21X1_103/Y OAI21X1_285/B INVX1_230/Y gnd NAND2X1_361/B vdd OAI21X1
XOAI21X1_263 AOI21X1_88/Y NOR2X1_157/Y INVX1_221/Y gnd NAND3X1_159/C vdd OAI21X1
XOAI21X1_241 INVX1_200/A INVX1_201/A NAND3X1_86/Y gnd NAND2X1_229/A vdd OAI21X1
XOAI21X1_230 INVX1_187/A NOR2X1_142/Y INVX2_21/A gnd INVX1_199/A vdd OAI21X1
XOAI21X1_274 AOI22X1_26/Y AOI22X1_27/Y OAI21X1_274/C gnd NAND3X1_175/A vdd OAI21X1
XAND2X2_30 INVX2_19/A INVX1_106/A gnd AND2X2_30/Y vdd AND2X2
XAND2X2_41 AND2X2_41/A AND2X2_41/B gnd AND2X2_41/Y vdd AND2X2
XFILL_17_2_0 gnd vdd FILL
XNAND2X1_291 AND2X2_34/B OR2X2_22/Y gnd NAND2X1_293/B vdd NAND2X1
XNAND2X1_280 INVX1_229/A NOR2X1_172/Y gnd NAND3X1_178/C vdd NAND2X1
XDFFPOSX1_19 INVX2_21/A CLKBUF1_5/Y DFFPOSX1_19/D gnd vdd DFFPOSX1
XINVX1_113 INVX1_113/A gnd INVX1_113/Y vdd INVX1
XINVX1_124 INVX1_124/A gnd INVX1_124/Y vdd INVX1
XINVX1_135 INVX1_135/A gnd INVX1_135/Y vdd INVX1
XINVX1_168 INVX1_168/A gnd INVX1_168/Y vdd INVX1
XINVX1_157 INVX1_157/A gnd INVX1_157/Y vdd INVX1
XINVX1_146 INVX1_146/A gnd INVX1_146/Y vdd INVX1
XINVX1_102 INVX2_19/A gnd INVX1_102/Y vdd INVX1
XINVX1_179 INVX1_179/A gnd INVX1_179/Y vdd INVX1
XAOI21X1_139 INVX1_282/Y AOI21X1_139/B INVX1_292/Y gnd OAI21X1_353/C vdd AOI21X1
XAOI21X1_117 NAND3X1_231/C NAND3X1_225/Y OR2X2_24/Y gnd OAI21X1_313/B vdd AOI21X1
XAOI21X1_128 NAND3X1_255/C NAND3X1_255/B INVX1_270/Y gnd AOI21X1_128/Y vdd AOI21X1
XAOI21X1_106 AND2X2_35/Y AND2X2_34/B INVX1_244/Y gnd AOI21X1_106/Y vdd AOI21X1
XFILL_23_0_0 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XNOR2X1_30 INVX1_50/Y NOR2X1_30/B gnd OAI22X1_4/C vdd NOR2X1
XNAND3X1_85 INVX1_198/A NAND3X1_85/B NAND3X1_85/C gnd NAND3X1_85/Y vdd NAND3X1
XNAND3X1_96 AOI21X1_76/Y NAND3X1_95/B NAND3X1_95/C gnd NAND3X1_98/A vdd NAND3X1
XNAND3X1_30 NAND3X1_28/Y NAND3X1_29/Y INVX2_11/Y gnd AOI22X1_6/A vdd NAND3X1
XNAND3X1_74 INVX1_185/A NAND3X1_70/Y NAND3X1_71/Y gnd NAND3X1_74/Y vdd NAND3X1
XNAND3X1_52 INVX1_175/Y NAND3X1_43/Y NAND3X1_52/C gnd NAND3X1_54/B vdd NAND3X1
XNAND3X1_63 INVX2_15/Y AOI21X1_56/B AOI21X1_56/A gnd AOI22X1_13/C vdd NAND3X1
XNAND3X1_41 INVX1_174/A NAND3X1_44/B NAND3X1_44/C gnd NAND3X1_48/B vdd NAND3X1
XNOR2X1_41 x2[3] INVX1_38/Y gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_63 INVX1_31/A INVX1_72/Y gnd NOR2X1_63/Y vdd NOR2X1
XNOR2X1_52 BUFX4_5/Y INVX1_86/Y gnd NOR2X1_52/Y vdd NOR2X1
XNOR2X1_85 NOR2X1_85/A OR2X2_5/B gnd NOR2X1_85/Y vdd NOR2X1
XNOR2X1_96 NOR2X1_69/Y NOR2X1_96/B gnd NOR2X1_96/Y vdd NOR2X1
XNOR2X1_74 NOR2X1_74/A NOR2X1_73/Y gnd INVX2_5/A vdd NOR2X1
XNAND2X1_7 x1[3] INVX1_11/Y gnd OAI21X1_8/C vdd NAND2X1
XNAND2X1_109 INVX2_29/A BUFX4_13/Y gnd OAI21X1_150/C vdd NAND2X1
XNOR2X1_131 AOI21X1_67/A NOR2X1_131/B gnd NOR2X1_131/Y vdd NOR2X1
XNOR2X1_120 gnd INVX2_12/Y gnd INVX1_164/A vdd NOR2X1
XNOR2X1_142 INVX2_17/Y INVX1_193/Y gnd NOR2X1_142/Y vdd NOR2X1
XNOR2X1_175 NOR2X1_175/A INVX1_231/Y gnd NOR2X1_175/Y vdd NOR2X1
XNOR2X1_197 INVX1_231/Y NOR2X1_197/B gnd NOR2X1_197/Y vdd NOR2X1
XNOR2X1_186 INVX1_243/Y NOR2X1_185/Y gnd NOR2X1_186/Y vdd NOR2X1
XNOR2X1_153 INVX1_207/Y NAND3X1_86/Y gnd INVX1_208/A vdd NOR2X1
XNOR2X1_164 gnd INVX2_28/A gnd NOR2X1_164/Y vdd NOR2X1
XINVX1_44 x2[4] gnd INVX1_44/Y vdd INVX1
XINVX1_22 x3[7] gnd INVX1_22/Y vdd INVX1
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XINVX1_33 x2[0] gnd INVX1_33/Y vdd INVX1
XINVX1_11 x3[3] gnd INVX1_11/Y vdd INVX1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XBUFX2_19 BUFX2_19/A gnd X2_mag[2] vdd BUFX2
XDFFPOSX1_7 OR2X2_6/B CLKBUF1_5/Y AND2X2_18/Y gnd vdd DFFPOSX1
XNAND3X1_282 INVX1_281/Y NAND3X1_282/B NAND3X1_282/C gnd NAND3X1_282/Y vdd NAND3X1
XNAND3X1_293 INVX2_43/Y AND2X2_45/Y OR2X2_32/Y gnd AOI22X1_49/A vdd NAND3X1
XNAND3X1_271 INVX1_272/Y INVX1_284/A AOI21X1_134/A gnd INVX1_277/A vdd NAND3X1
XNAND3X1_260 AOI21X1_131/Y NAND3X1_255/B NAND3X1_255/C gnd NAND3X1_261/C vdd NAND3X1
XOAI22X1_17 NOR3X1_2/C NOR2X1_123/Y OAI22X1_17/C NOR2X1_128/Y gnd NAND3X1_58/B vdd
+ OAI22X1
XNAND2X1_440 INVX1_311/A OAI21X1_387/Y gnd NAND2X1_440/Y vdd NAND2X1
XFILL_8_2 gnd vdd FILL
XOAI21X1_83 AND2X2_11/Y OAI21X1_82/Y OAI21X1_83/C gnd OAI21X1_83/Y vdd OAI21X1
XOAI21X1_72 INVX1_25/Y OAI21X1_72/B BUFX4_3/Y gnd OAI22X1_6/D vdd OAI21X1
XOAI21X1_61 BUFX4_15/Y OAI21X1_61/B NAND2X1_34/Y gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_94 BUFX4_1/Y INVX1_96/Y NAND2X1_57/Y gnd OAI21X1_94/Y vdd OAI21X1
XOAI21X1_50 BUFX4_5/Y INVX1_65/Y NAND2X1_33/Y gnd OAI21X1_50/Y vdd OAI21X1
XFILL_1_2_1 gnd vdd FILL
XINVX1_306 INVX1_306/A gnd INVX1_306/Y vdd INVX1
XOAI21X1_297 INVX1_230/A AOI21X1_103/Y AOI21X1_108/C gnd OAI21X1_297/Y vdd OAI21X1
XOAI21X1_286 NAND2X1_293/A NAND2X1_293/B OR2X2_22/Y gnd OAI21X1_286/Y vdd OAI21X1
XAND2X2_31 AND2X2_31/A AND2X2_31/B gnd AND2X2_31/Y vdd AND2X2
XOAI21X1_253 INVX2_18/Y INVX1_213/Y NAND3X1_99/B gnd AND2X2_31/B vdd OAI21X1
XOAI21X1_275 OAI22X1_19/C NOR2X1_160/Y NAND3X1_170/C gnd OAI21X1_275/Y vdd OAI21X1
XOAI21X1_242 OAI21X1_242/A OAI21X1_242/B INVX1_218/A gnd AOI21X1_85/C vdd OAI21X1
XOAI21X1_264 INVX2_23/Y INVX2_25/A OR2X2_19/Y gnd OAI21X1_265/C vdd OAI21X1
XAND2X2_20 AND2X2_20/A AND2X2_20/B gnd OR2X2_12/A vdd AND2X2
XOAI21X1_231 INVX2_23/A INVX1_193/A INVX1_187/A gnd AOI21X1_74/C vdd OAI21X1
XOAI21X1_220 INVX2_19/A INVX1_103/A INVX2_18/A gnd NOR2X1_140/A vdd OAI21X1
XNAND2X1_270 INVX1_225/Y AOI21X1_94/Y gnd NAND2X1_270/Y vdd NAND2X1
XAND2X2_42 AND2X2_42/A AND2X2_42/B gnd AND2X2_42/Y vdd AND2X2
XFILL_17_2_1 gnd vdd FILL
XNAND2X1_292 AND2X2_35/B INVX1_234/Y gnd NAND2X1_293/A vdd NAND2X1
XNAND2X1_281 NAND3X1_178/A NAND3X1_178/C gnd NAND2X1_281/Y vdd NAND2X1
XINVX1_114 INVX1_114/A gnd INVX1_114/Y vdd INVX1
XINVX1_136 INVX1_136/A gnd INVX1_136/Y vdd INVX1
XINVX1_169 INVX1_169/A gnd INVX1_169/Y vdd INVX1
XINVX1_158 INVX1_158/A gnd INVX1_158/Y vdd INVX1
XINVX1_125 INVX1_125/A gnd INVX1_125/Y vdd INVX1
XINVX1_147 INVX1_147/A gnd INVX1_147/Y vdd INVX1
XINVX1_103 INVX1_103/A gnd INVX1_103/Y vdd INVX1
XAOI21X1_118 NOR2X1_168/Y INVX1_266/Y NOR3X1_9/B gnd OR2X2_26/B vdd AOI21X1
XAOI21X1_107 NAND2X1_313/B INVX1_230/Y OAI21X1_285/B gnd NAND3X1_194/A vdd AOI21X1
XAOI21X1_129 NAND3X1_232/B NAND3X1_232/A NOR2X1_194/Y gnd AOI21X1_130/C vdd AOI21X1
XFILL_23_0_1 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XNOR2X1_31 x0[7] x2[7] gnd NOR2X1_31/Y vdd NOR2X1
XNOR2X1_20 x2[1] INVX1_35/Y gnd AOI21X1_6/C vdd NOR2X1
XNOR2X1_42 INVX1_6/Y INVX1_7/Y gnd NOR2X1_42/Y vdd NOR2X1
XNOR2X1_64 NOR2X1_64/A INVX1_73/Y gnd NOR2X1_64/Y vdd NOR2X1
XNAND3X1_97 NAND3X1_97/A NAND3X1_92/B NAND3X1_92/C gnd NAND3X1_97/Y vdd NAND3X1
XNAND3X1_53 INVX1_175/A NAND3X1_48/Y NAND3X1_49/Y gnd NAND3X1_54/C vdd NAND3X1
XNAND3X1_31 INVX2_11/A NAND3X1_24/Y NAND3X1_27/Y gnd AOI22X1_6/B vdd NAND3X1
XNAND3X1_75 NAND3X1_75/A NAND3X1_74/Y NAND3X1_75/C gnd NAND3X1_75/Y vdd NAND3X1
XNAND3X1_64 INVX1_173/Y NAND3X1_40/Y AOI21X1_58/A gnd AOI22X1_13/A vdd NAND3X1
XNAND3X1_42 INVX1_174/Y NAND3X1_42/B NAND3X1_42/C gnd NAND3X1_48/C vdd NAND3X1
XNAND3X1_86 OR2X2_18/B NAND3X1_86/B OR2X2_17/Y gnd NAND3X1_86/Y vdd NAND3X1
XNAND3X1_20 INVX2_9/A INVX1_151/Y NAND3X1_20/C gnd AND2X2_21/B vdd NAND3X1
XNOR2X1_53 BUFX4_7/Y INVX1_87/Y gnd NOR2X1_53/Y vdd NOR2X1
XNOR2X1_97 NOR2X1_97/A NOR2X1_97/B gnd NOR2X1_97/Y vdd NOR2X1
XNOR2X1_75 NOR2X1_69/Y INVX2_5/A gnd NOR2X1_75/Y vdd NOR2X1
XNOR2X1_86 INVX1_86/A INVX1_57/Y gnd NOR2X1_86/Y vdd NOR2X1
XNAND2X1_8 INVX1_16/A OAI21X1_8/C gnd XOR2X1_2/B vdd NAND2X1
XNOR2X1_176 INVX2_29/A INVX2_33/Y gnd NOR2X1_176/Y vdd NOR2X1
XNOR2X1_110 INVX2_8/Y INVX1_142/Y gnd NOR2X1_110/Y vdd NOR2X1
XNOR2X1_154 OR2X2_19/A OR2X2_19/B gnd NOR2X1_154/Y vdd NOR2X1
XNOR2X1_121 INVX1_172/A NOR2X1_121/B gnd INVX1_171/A vdd NOR2X1
XNOR2X1_143 INVX1_187/A INVX2_21/Y gnd NOR2X1_143/Y vdd NOR2X1
XNOR2X1_132 INVX2_17/Y INVX2_18/Y gnd NOR2X1_132/Y vdd NOR2X1
XNOR2X1_165 NOR2X1_164/Y NOR2X1_163/Y gnd NOR2X1_165/Y vdd NOR2X1
XNOR2X1_187 INVX1_230/A NOR2X1_187/B gnd NOR2X1_187/Y vdd NOR2X1
XNOR2X1_198 XOR2X1_18/B NOR2X1_197/Y gnd NOR2X1_198/Y vdd NOR2X1
XINVX1_23 x1[7] gnd INVX1_23/Y vdd INVX1
XINVX1_34 x2[1] gnd INVX1_34/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XDFFPOSX1_8 INVX1_132/A CLKBUF1_9/Y AOI22X1_5/Y gnd vdd DFFPOSX1
XNAND3X1_294 INVX2_43/Y OR2X2_32/Y INVX1_296/Y gnd AOI22X1_48/D vdd NAND3X1
XNAND3X1_272 INVX2_37/Y INVX1_95/A INVX1_278/Y gnd NAND2X1_387/A vdd NAND3X1
XNAND3X1_283 NAND3X1_287/A NAND3X1_281/Y NAND3X1_282/Y gnd NAND3X1_283/Y vdd NAND3X1
XNAND3X1_250 NAND3X1_248/Y AOI21X1_125/Y NAND3X1_249/Y gnd AOI22X1_36/C vdd NAND3X1
XNAND3X1_261 OAI21X1_328/Y NAND3X1_261/B NAND3X1_261/C gnd NAND3X1_262/B vdd NAND3X1
XOAI22X1_18 INVX1_205/A INVX2_26/A INVX1_212/A OAI22X1_18/D gnd OAI22X1_18/Y vdd OAI22X1
XNAND2X1_441 NAND2X1_441/A NAND2X1_440/Y gnd NAND2X1_441/Y vdd NAND2X1
XNAND2X1_430 OR2X2_33/B OR2X2_33/A gnd NAND3X1_353/B vdd NAND2X1
XOAI21X1_84 INVX1_28/A NOR3X1_1/C INVX2_4/A gnd OAI21X1_84/Y vdd OAI21X1
XOAI21X1_73 INVX1_23/Y INVX1_22/Y BUFX4_8/Y gnd NOR2X1_48/A vdd OAI21X1
XOAI21X1_95 BUFX4_6/Y INVX1_97/Y OAI21X1_95/C gnd OAI21X1_95/Y vdd OAI21X1
XOAI21X1_40 BUFX4_12/Y XNOR2X1_9/Y OAI21X1_40/C gnd OAI21X1_40/Y vdd OAI21X1
XOAI21X1_62 BUFX4_15/Y XOR2X1_2/Y OAI21X1_62/C gnd OAI21X1_62/Y vdd OAI21X1
XOAI21X1_51 BUFX4_1/Y INVX1_66/Y NAND2X1_33/Y gnd OAI21X1_51/Y vdd OAI21X1
XFILL_1_2_2 gnd vdd FILL
XOAI21X1_210 NOR3X1_3/B NOR3X1_3/C INVX2_15/A gnd AOI22X1_13/D vdd OAI21X1
XOAI21X1_221 NOR2X1_140/A NOR2X1_140/B INVX1_188/Y gnd NAND3X1_78/A vdd OAI21X1
XAND2X2_43 AND2X2_43/A AND2X2_43/B gnd AND2X2_43/Y vdd AND2X2
XAND2X2_10 NOR2X1_58/Y INVX2_2/Y gnd AND2X2_10/Y vdd AND2X2
XINVX1_307 INVX1_307/A gnd INVX1_307/Y vdd INVX1
XAND2X2_32 AND2X2_32/A AND2X2_32/B gnd AND2X2_32/Y vdd AND2X2
XOAI21X1_265 AOI22X1_25/Y XNOR2X1_34/A OAI21X1_265/C gnd AND2X2_32/B vdd OAI21X1
XOAI21X1_298 INVX1_236/A INVX1_239/A INVX1_245/Y gnd NAND2X1_318/A vdd OAI21X1
XOAI21X1_287 gnd XOR2X1_17/A gnd gnd INVX1_236/A vdd OAI21X1
XOAI21X1_254 NOR3X1_7/Y AOI21X1_78/Y INVX1_211/Y gnd NAND2X1_251/B vdd OAI21X1
XOAI21X1_276 INVX1_227/Y INVX2_30/Y INVX2_31/Y gnd AND2X2_33/A vdd OAI21X1
XOAI21X1_232 INVX1_192/A NOR2X1_148/B INVX1_201/A gnd INVX1_203/A vdd OAI21X1
XOAI21X1_243 INVX2_23/Y INVX1_200/A NAND3X1_86/B gnd INVX1_211/A vdd OAI21X1
XAND2X2_21 AND2X2_21/A AND2X2_21/B gnd AND2X2_21/Y vdd AND2X2
XNAND2X1_271 INVX1_225/A NAND2X1_271/B gnd NAND2X1_272/B vdd NAND2X1
XNAND2X1_293 NAND2X1_293/A NAND2X1_293/B gnd NAND3X1_182/B vdd NAND2X1
XNAND2X1_260 NAND2X1_259/Y NAND2X1_260/B gnd NAND3X1_157/B vdd NAND2X1
XNAND2X1_282 NAND3X1_178/Y NAND2X1_282/B gnd OR2X2_21/A vdd NAND2X1
XFILL_17_2_2 gnd vdd FILL
XINVX1_115 INVX1_115/A gnd INVX1_115/Y vdd INVX1
XINVX1_137 INVX1_137/A gnd OR2X2_9/B vdd INVX1
XINVX1_159 OR2X2_10/Y gnd INVX1_159/Y vdd INVX1
XINVX1_104 INVX1_104/A gnd INVX1_104/Y vdd INVX1
XINVX1_126 INVX1_126/A gnd INVX1_126/Y vdd INVX1
XINVX1_148 INVX1_148/A gnd INVX1_148/Y vdd INVX1
XAOI21X1_119 NAND3X1_245/C NAND3X1_212/Y XNOR2X1_39/Y gnd OAI21X1_316/B vdd AOI21X1
XAOI21X1_108 NAND3X1_194/B NAND3X1_194/C AOI21X1_108/C gnd INVX1_265/A vdd AOI21X1
XFILL_23_0_2 gnd vdd FILL
XFILL_6_1_2 gnd vdd FILL
XFILL_14_0_2 gnd vdd FILL
XFILL_18_1 gnd vdd FILL
XNAND3X1_10 NOR2X1_95/B NOR2X1_95/A AOI21X1_17/B gnd NAND3X1_11/C vdd NAND3X1
XNAND3X1_32 AOI22X1_6/A AOI22X1_6/B INVX1_160/Y gnd NAND3X1_32/Y vdd NAND3X1
XNAND3X1_21 INVX1_156/Y NAND3X1_21/B NAND3X1_21/C gnd INVX2_14/A vdd NAND3X1
XNOR2X1_21 NOR2X1_21/A AOI21X1_6/C gnd AOI21X1_6/A vdd NOR2X1
XNOR2X1_10 x1[6] INVX1_21/Y gnd NOR2X1_10/Y vdd NOR2X1
XNOR2X1_32 NOR2X1_31/Y INVX1_51/Y gnd INVX1_53/A vdd NOR2X1
XNOR2X1_43 INVX1_10/Y INVX1_11/Y gnd NOR2X1_43/Y vdd NOR2X1
XNAND3X1_54 AOI22X1_6/A NAND3X1_54/B NAND3X1_54/C gnd NAND3X1_54/Y vdd NAND3X1
XNOR2X1_65 INVX1_110/A NOR2X1_65/B gnd NOR2X1_65/Y vdd NOR2X1
XNOR2X1_54 BUFX4_7/Y INVX1_88/Y gnd NOR2X1_54/Y vdd NOR2X1
XNAND3X1_76 INVX2_17/A INVX1_187/A INVX2_20/Y gnd INVX1_186/A vdd NAND3X1
XNAND3X1_98 NAND3X1_98/A NAND3X1_97/Y XOR2X1_13/B gnd NAND3X1_98/Y vdd NAND3X1
XNAND3X1_65 INVX1_173/A NAND3X1_36/Y AOI21X1_57/A gnd AOI22X1_13/B vdd NAND3X1
XNAND3X1_87 NAND3X1_87/A NAND3X1_87/B NOR2X1_149/Y gnd NAND3X1_87/Y vdd NAND3X1
XNAND3X1_43 INVX1_161/Y NAND3X1_48/B NAND3X1_48/C gnd NAND3X1_43/Y vdd NAND3X1
XNOR2X1_76 INVX1_55/A INVX1_84/A gnd NOR2X1_78/A vdd NOR2X1
XNOR2X1_87 INVX1_57/A INVX1_86/Y gnd NOR2X1_87/Y vdd NOR2X1
XNOR2X1_98 NOR2X1_98/A INVX2_6/A gnd NOR2X1_98/Y vdd NOR2X1
XNAND2X1_9 NOR2X1_56/A BUFX4_15/Y gnd OAI21X1_7/C vdd NAND2X1
XNOR2X1_199 INVX2_35/Y INVX2_36/Y gnd NOR2X1_199/Y vdd NOR2X1
XNOR2X1_100 INVX1_59/Y INVX1_88/Y gnd NOR2X1_100/Y vdd NOR2X1
XNOR2X1_188 INVX1_245/Y AOI22X1_32/D gnd INVX1_246/A vdd NOR2X1
XNOR2X1_111 gnd INVX1_144/Y gnd NOR2X1_111/Y vdd NOR2X1
XNOR2X1_177 INVX2_27/Y INVX1_232/Y gnd XOR2X1_17/A vdd NOR2X1
XNOR2X1_122 INVX2_9/Y INVX2_16/Y gnd NOR2X1_122/Y vdd NOR2X1
XNOR2X1_166 INVX2_28/A INVX2_29/Y gnd INVX2_30/A vdd NOR2X1
XNOR2X1_155 INVX2_21/A INVX2_23/Y gnd INVX1_210/A vdd NOR2X1
XNOR2X1_144 NAND3X1_77/Y INVX1_194/Y gnd INVX1_195/A vdd NOR2X1
XNOR2X1_133 INVX2_17/A INVX2_18/A gnd NOR2X1_133/Y vdd NOR2X1
XINVX1_13 x3[4] gnd INVX1_13/Y vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XINVX1_35 x0[1] gnd INVX1_35/Y vdd INVX1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XDFFPOSX1_9 INVX2_18/A CLKBUF1_10/Y DFFPOSX1_9/D gnd vdd DFFPOSX1
XNAND3X1_284 INVX1_281/Y INVX1_305/A NAND3X1_281/C gnd NAND3X1_287/B vdd NAND3X1
XNAND3X1_295 AOI22X1_48/C AOI22X1_48/D NAND3X1_295/C gnd AOI21X1_142/A vdd NAND3X1
XNAND3X1_273 NAND3X1_273/A NOR2X1_209/Y NAND2X1_387/A gnd NAND2X1_372/A vdd NAND3X1
XNAND3X1_240 NAND2X1_317/Y NAND3X1_237/B NAND3X1_236/Y gnd AOI21X1_115/B vdd NAND3X1
XNAND3X1_251 NAND3X1_248/Y NAND3X1_249/Y OAI21X1_316/Y gnd AOI21X1_126/A vdd NAND3X1
XNAND3X1_262 AOI21X1_130/Y NAND3X1_262/B NAND3X1_262/C gnd AOI22X1_37/B vdd NAND3X1
XFILL_21_1_0 gnd vdd FILL
XOAI22X1_19 AOI21X1_98/Y AOI21X1_99/Y OAI22X1_19/C NOR2X1_160/Y gnd OAI22X1_19/Y vdd
+ OAI22X1
XNAND2X1_431 OAI21X1_378/Y NAND2X1_431/B gnd NAND3X1_349/A vdd NAND2X1
XNAND2X1_442 NAND3X1_360/Y NAND3X1_358/Y gnd OAI21X1_392/C vdd NAND2X1
XNAND2X1_420 NAND2X1_420/A NAND2X1_420/B gnd OAI21X1_375/A vdd NAND2X1
XFILL_4_2_0 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XOAI21X1_41 OAI21X1_41/A NOR2X1_31/Y INVX1_51/A gnd NOR2X1_33/B vdd OAI21X1
XOAI21X1_30 INVX1_35/Y INVX1_34/Y OAI21X1_27/Y gnd AOI21X1_4/B vdd OAI21X1
XOAI21X1_63 NOR2X1_5/Y AND2X2_8/Y BUFX4_3/Y gnd OAI22X1_5/C vdd OAI21X1
XOAI21X1_52 BUFX4_9/Y INVX1_67/Y NAND2X1_33/Y gnd OAI21X1_52/Y vdd OAI21X1
XOAI21X1_85 NOR3X1_1/C NOR3X1_1/B OAI21X1_84/Y gnd OAI21X1_85/Y vdd OAI21X1
XOAI21X1_74 INVX1_24/A NOR2X1_58/B BUFX4_6/Y gnd OAI21X1_74/Y vdd OAI21X1
XOAI21X1_96 BUFX4_7/Y INVX1_98/Y NAND2X1_59/Y gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_222 INVX2_20/Y INVX2_22/Y OAI21X1_222/C gnd OAI21X1_222/Y vdd OAI21X1
XOAI21X1_255 AOI21X1_94/C AOI21X1_81/Y AOI21X1_94/B gnd AOI21X1_96/A vdd OAI21X1
XOAI21X1_211 NOR3X1_5/A NOR3X1_5/C NOR3X1_5/B gnd NAND3X1_66/B vdd OAI21X1
XOAI21X1_244 INVX2_25/A NOR2X1_154/Y AND2X2_28/Y gnd AOI22X1_22/B vdd OAI21X1
XOAI21X1_200 INVX1_171/A INVX1_169/Y XNOR2X1_23/Y gnd NAND3X1_40/B vdd OAI21X1
XOAI21X1_233 INVX1_205/Y NOR2X1_150/Y NOR2X1_140/B gnd NAND3X1_87/A vdd OAI21X1
XAND2X2_11 NOR3X1_1/C INVX1_28/A gnd AND2X2_11/Y vdd AND2X2
XAND2X2_44 AND2X2_44/A AND2X2_44/B gnd AND2X2_44/Y vdd AND2X2
XINVX1_308 XOR2X1_25/Y gnd INVX1_308/Y vdd INVX1
XOAI21X1_266 NAND2X1_248/Y AOI21X1_91/Y NAND3X1_111/Y gnd OAI21X1_266/Y vdd OAI21X1
XOAI21X1_299 INVX2_32/Y INVX1_237/A NAND2X1_299/A gnd INVX1_254/A vdd OAI21X1
XOAI21X1_288 gnd gnd gnd gnd OAI21X1_288/Y vdd OAI21X1
XOAI21X1_277 gnd INVX2_30/A INVX2_31/A gnd AND2X2_33/B vdd OAI21X1
XAND2X2_33 AND2X2_33/A AND2X2_33/B gnd AND2X2_33/Y vdd AND2X2
XAND2X2_22 AND2X2_22/A AND2X2_22/B gnd AND2X2_22/Y vdd AND2X2
XNAND2X1_272 NAND2X1_270/Y NAND2X1_272/B gnd NAND3X1_168/C vdd NAND2X1
XNAND2X1_294 NAND2X1_293/B AND2X2_35/Y gnd NAND2X1_294/Y vdd NAND2X1
XNAND2X1_283 OR2X2_21/B OR2X2_21/A gnd AOI21X1_101/B vdd NAND2X1
XNAND2X1_250 AND2X2_31/B AND2X2_31/A gnd XNOR2X1_34/A vdd NAND2X1
XNAND2X1_261 AOI21X1_89/Y XOR2X1_15/Y gnd NAND2X1_263/A vdd NAND2X1
XFILL_6_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XINVX1_116 INVX1_116/A gnd INVX1_116/Y vdd INVX1
XINVX1_105 INVX1_105/A gnd INVX1_105/Y vdd INVX1
XINVX1_127 INVX1_127/A gnd AOI22X1_3/B vdd INVX1
XINVX1_138 INVX1_138/A gnd INVX1_138/Y vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XINVX1_149 INVX1_149/A gnd OAI22X1_7/A vdd INVX1
XFILL_17_0_0 gnd vdd FILL
XAOI21X1_109 NAND3X1_199/C NAND3X1_199/B INVX2_34/Y gnd AOI21X1_109/Y vdd AOI21X1
XFILL_18_2 gnd vdd FILL
XNAND3X1_11 NAND2X1_68/A NAND3X1_11/B NAND3X1_11/C gnd AOI21X1_19/B vdd NAND3X1
XNAND3X1_33 NOR3X1_6/A INVX1_140/Y NAND3X1_33/C gnd NAND3X1_33/Y vdd NAND3X1
XNAND3X1_66 NAND3X1_62/Y NAND3X1_66/B NAND3X1_66/C gnd NAND3X1_66/Y vdd NAND3X1
XNAND3X1_55 NAND3X1_55/A OR2X2_14/Y INVX1_179/A gnd NAND3X1_55/Y vdd NAND3X1
XNAND3X1_44 INVX1_174/Y NAND3X1_44/B NAND3X1_44/C gnd NAND3X1_49/B vdd NAND3X1
XNAND3X1_22 NAND3X1_22/A OAI22X1_7/Y OAI22X1_8/Y gnd NAND3X1_22/Y vdd NAND3X1
XNOR2X1_22 x0[2] x2[2] gnd NOR2X1_22/Y vdd NOR2X1
XNOR2X1_11 x3[6] INVX2_1/Y gnd INVX1_26/A vdd NOR2X1
XNOR2X1_33 BUFX4_14/Y NOR2X1_33/B gnd AOI22X1_1/C vdd NOR2X1
XNOR2X1_44 NOR2X1_4/B INVX1_13/Y gnd INVX1_77/A vdd NOR2X1
XNOR2X1_55 INVX1_1/A INVX1_4/A gnd NOR2X1_55/Y vdd NOR2X1
XNOR2X1_66 XOR2X1_4/Y NOR2X1_66/B gnd NOR2X1_66/Y vdd NOR2X1
XNAND3X1_88 INVX1_202/Y NAND3X1_89/B NAND3X1_87/Y gnd AOI22X1_17/C vdd NAND3X1
XNAND3X1_99 INVX2_25/Y NAND3X1_99/B OR2X2_19/Y gnd NAND3X1_99/Y vdd NAND3X1
XNOR2X1_77 INVX1_55/Y INVX1_84/Y gnd NOR2X1_77/Y vdd NOR2X1
XNOR2X1_88 NOR2X1_86/Y NOR2X1_87/Y gnd AND2X2_16/B vdd NOR2X1
XNOR2X1_99 INVX2_7/Y AND2X2_17/A gnd NOR2X1_99/Y vdd NOR2X1
XNAND3X1_77 INVX1_187/A INVX2_23/A INVX2_22/A gnd NAND3X1_77/Y vdd NAND3X1
XNOR2X1_134 NOR2X1_133/Y NOR2X1_132/Y gnd NOR2X1_134/Y vdd NOR2X1
XNOR2X1_101 INVX2_8/Y INVX2_9/Y gnd NOR2X1_101/Y vdd NOR2X1
XNOR2X1_112 OR2X2_11/B OR2X2_11/A gnd NOR2X1_112/Y vdd NOR2X1
XNOR2X1_189 OR2X2_25/A OR2X2_25/B gnd NOR3X1_8/C vdd NOR2X1
XNOR2X1_178 gnd INVX1_228/Y gnd XOR2X1_17/B vdd NOR2X1
XNOR2X1_123 INVX1_144/Y NOR2X1_123/B gnd NOR2X1_123/Y vdd NOR2X1
XNOR2X1_167 INVX2_27/Y INVX1_228/Y gnd INVX2_31/A vdd NOR2X1
XNOR2X1_156 INVX1_218/Y NOR2X1_156/B gnd NOR2X1_156/Y vdd NOR2X1
XNOR2X1_145 INVX1_200/A INVX1_201/A gnd INVX1_207/A vdd NOR2X1
XINVX1_36 x0[2] gnd INVX1_36/Y vdd INVX1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_14 x1[4] gnd NOR2X1_4/B vdd INVX1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XNAND3X1_241 INVX1_265/Y NAND3X1_239/Y AOI21X1_115/B gnd NAND2X1_338/B vdd NAND3X1
XNAND3X1_230 INVX1_247/Y NAND3X1_230/B NAND3X1_230/C gnd NAND3X1_234/B vdd NAND3X1
XNAND3X1_285 INVX1_281/A NAND3X1_282/B NAND3X1_282/C gnd NAND3X1_287/C vdd NAND3X1
XNAND3X1_296 INVX2_42/Y OAI21X1_374/C AOI21X1_142/A gnd NAND3X1_326/C vdd NAND3X1
XNAND3X1_274 INVX1_283/A NAND2X1_379/Y NAND2X1_376/Y gnd AOI21X1_141/C vdd NAND3X1
XNAND3X1_263 NAND2X1_317/Y INVX1_246/Y NAND2X1_359/Y gnd AOI22X1_37/D vdd NAND3X1
XNAND3X1_252 NAND3X1_244/Y AOI21X1_125/Y NAND3X1_246/Y gnd AOI21X1_126/B vdd NAND3X1
XFILL_21_1_1 gnd vdd FILL
XNAND2X1_410 NAND2X1_410/A OAI21X1_363/Y gnd NAND2X1_410/Y vdd NAND2X1
XNAND2X1_432 INVX2_35/A INVX1_92/A gnd XOR2X1_25/B vdd NAND2X1
XNAND2X1_443 NAND3X1_343/B NAND3X1_343/C gnd AOI21X1_166/A vdd NAND2X1
XNAND2X1_421 AND2X2_45/Y AND2X2_46/Y gnd AND2X2_48/A vdd NAND2X1
XFILL_4_2_1 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XOAI21X1_42 NOR2X1_22/Y INVX1_42/A INVX1_40/A gnd OAI21X1_42/Y vdd OAI21X1
XOAI21X1_86 BUFX4_14/Y OAI21X1_85/Y OAI21X1_86/C gnd OAI21X1_86/Y vdd OAI21X1
XOAI21X1_64 NOR2X1_5/Y AND2X2_8/Y INVX1_77/Y gnd XOR2X1_3/A vdd OAI21X1
XOAI21X1_75 OAI21X1_75/A OAI21X1_74/Y OAI21X1_75/C gnd OAI21X1_75/Y vdd OAI21X1
XOAI21X1_53 BUFX4_8/Y INVX1_68/Y NAND2X1_33/Y gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_20 BUFX4_6/Y INVX1_27/Y OAI21X1_21/C gnd OAI21X1_20/Y vdd OAI21X1
XOAI21X1_31 BUFX4_15/Y XNOR2X1_6/Y NAND2X1_17/Y gnd OAI21X1_31/Y vdd OAI21X1
XOAI21X1_97 BUFX4_1/Y INVX1_99/Y NAND2X1_60/Y gnd OAI21X1_97/Y vdd OAI21X1
XOAI21X1_223 OR2X2_15/B OR2X2_15/A NAND3X1_78/Y gnd INVX1_197/A vdd OAI21X1
XOAI21X1_256 INVX1_209/A AOI21X1_85/Y NAND3X1_142/B gnd AOI21X1_99/C vdd OAI21X1
XOAI21X1_278 INVX1_227/Y INVX2_31/Y INVX1_229/Y gnd NAND2X1_279/B vdd OAI21X1
XOAI21X1_212 NOR3X1_5/Y AOI21X1_64/Y NOR2X1_130/Y gnd AOI22X1_15/B vdd OAI21X1
XOAI21X1_289 NOR2X1_183/A NOR2X1_183/B INVX1_238/A gnd INVX1_241/A vdd OAI21X1
XOAI21X1_245 INVX2_25/A NOR2X1_154/Y INVX1_210/Y gnd AOI22X1_23/C vdd OAI21X1
XOAI21X1_267 INVX2_25/A NAND3X1_99/B OR2X2_19/Y gnd XOR2X1_16/A vdd OAI21X1
XOAI21X1_234 INVX2_19/Y INVX1_189/Y NOR2X1_151/Y gnd NAND3X1_87/B vdd OAI21X1
XOAI21X1_201 INVX2_16/Y XOR2X1_6/B AOI21X1_61/B gnd AND2X2_24/A vdd OAI21X1
XAND2X2_45 INVX2_35/A AND2X2_45/B gnd AND2X2_45/Y vdd AND2X2
XAND2X2_12 AND2X2_12/A NAND3X1_9/C gnd AND2X2_12/Y vdd AND2X2
XINVX1_309 INVX1_309/A gnd INVX1_309/Y vdd INVX1
XAND2X2_34 OR2X2_22/Y AND2X2_34/B gnd AND2X2_34/Y vdd AND2X2
XAND2X2_23 OR2X2_13/Y AND2X2_23/B gnd AND2X2_23/Y vdd AND2X2
XNAND2X1_295 NAND2X1_293/A AND2X2_34/Y gnd NAND2X1_295/Y vdd NAND2X1
XNAND2X1_262 XNOR2X1_36/Y NAND2X1_258/B gnd NAND2X1_263/B vdd NAND2X1
XNAND2X1_284 INVX1_226/Y NOR2X1_173/Y gnd INVX1_231/A vdd NAND2X1
XNAND2X1_251 NAND2X1_251/A NAND2X1_251/B gnd NAND2X1_251/Y vdd NAND2X1
XNAND2X1_240 INVX1_103/A INVX1_105/A gnd INVX2_26/A vdd NAND2X1
XNAND2X1_273 NAND3X1_169/Y NAND3X1_167/Y gnd NAND3X1_170/C vdd NAND2X1
XCLKBUF1_10 clk gnd CLKBUF1_10/Y vdd CLKBUF1
XFILL_1_0_1 gnd vdd FILL
XINVX1_139 INVX1_139/A gnd INVX1_139/Y vdd INVX1
XINVX1_106 INVX1_106/A gnd INVX1_106/Y vdd INVX1
XINVX1_117 NOR2X1_69/Y gnd NOR2X1_70/A vdd INVX1
XINVX1_128 XOR2X1_5/Y gnd INVX1_128/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XNOR2X1_12 NOR2X1_10/Y INVX1_26/A gnd INVX1_79/A vdd NOR2X1
XNAND3X1_12 INVX1_115/A NAND3X1_12/B AOI21X1_30/Y gnd NAND3X1_12/Y vdd NAND3X1
XNAND3X1_78 NAND3X1_78/A NAND3X1_78/B NAND3X1_78/C gnd NAND3X1_78/Y vdd NAND3X1
XNAND3X1_67 NAND3X1_62/Y NAND3X1_66/B NOR2X1_130/Y gnd AOI21X1_66/A vdd NAND3X1
XNAND3X1_56 AOI21X1_62/Y NAND3X1_55/Y NAND3X1_56/C gnd NAND3X1_56/Y vdd NAND3X1
XNAND3X1_34 INVX1_165/Y AOI22X1_9/C INVX1_167/Y gnd AOI21X1_56/A vdd NAND3X1
XNAND3X1_45 INVX1_174/A NAND3X1_42/B NAND3X1_42/C gnd NAND3X1_49/C vdd NAND3X1
XNAND3X1_89 INVX1_202/A NAND3X1_89/B NAND3X1_87/Y gnd INVX1_218/A vdd NAND3X1
XNAND3X1_23 NAND3X1_25/A OAI22X1_10/Y OAI22X1_9/Y gnd NAND3X1_23/Y vdd NAND3X1
XNOR2X1_23 INVX1_36/Y INVX1_37/Y gnd INVX1_42/A vdd NOR2X1
XNOR2X1_45 NOR2X1_45/A AND2X2_8/Y gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_56 NOR2X1_56/A NOR2X1_56/B gnd NOR2X1_56/Y vdd NOR2X1
XNOR2X1_67 INVX1_52/A INVX1_82/A gnd NOR2X1_69/A vdd NOR2X1
XNOR2X1_78 NOR2X1_78/A NOR2X1_77/Y gnd NOR2X1_85/A vdd NOR2X1
XNOR2X1_89 AND2X2_16/B NOR2X1_89/B gnd NOR2X1_89/Y vdd NOR2X1
XNOR2X1_34 BUFX4_9/Y INVX1_54/Y gnd NOR2X1_34/Y vdd NOR2X1
XNOR2X1_102 gnd INVX2_9/A gnd NOR2X1_102/Y vdd NOR2X1
XNOR2X1_124 INVX1_181/A OR2X2_13/Y gnd NOR2X1_124/Y vdd NOR2X1
XNOR2X1_113 OR2X2_12/B OR2X2_12/A gnd NOR2X1_113/Y vdd NOR2X1
XFILL_23_1 gnd vdd FILL
XNOR2X1_179 NOR2X1_179/A INVX1_233/Y gnd INVX1_234/A vdd NOR2X1
XNOR2X1_157 NOR2X1_157/A XNOR2X1_36/Y gnd NOR2X1_157/Y vdd NOR2X1
XNOR2X1_168 INVX1_228/Y INVX2_32/Y gnd NOR2X1_168/Y vdd NOR2X1
XNOR2X1_146 INVX1_200/Y INVX1_201/Y gnd NOR2X1_147/B vdd NOR2X1
XNOR2X1_135 INVX2_18/A INVX2_19/Y gnd INVX2_20/A vdd NOR2X1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XINVX1_48 x0[6] gnd INVX1_48/Y vdd INVX1
XINVX1_37 x2[2] gnd INVX1_37/Y vdd INVX1
XINVX1_15 NOR2X1_5/Y gnd INVX1_15/Y vdd INVX1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XNAND3X1_275 INVX1_283/Y NAND3X1_275/B NAND2X1_380/Y gnd AOI21X1_140/B vdd NAND3X1
XNAND3X1_231 NAND3X1_225/Y NOR2X1_194/Y NAND3X1_231/C gnd NAND3X1_233/B vdd NAND3X1
XNAND3X1_253 INVX1_271/A AOI21X1_126/B AOI21X1_126/A gnd NAND3X1_255/B vdd NAND3X1
XNAND3X1_220 INVX1_262/A NAND3X1_218/Y NAND3X1_219/Y gnd NAND3X1_221/C vdd NAND3X1
XNAND3X1_264 OAI21X1_313/Y NAND3X1_262/B NAND3X1_262/C gnd AOI22X1_38/B vdd NAND3X1
XNAND3X1_242 INVX1_268/A INVX1_269/Y NAND3X1_242/C gnd AND2X2_41/B vdd NAND3X1
XNAND3X1_297 NAND3X1_326/B INVX1_297/Y NAND3X1_326/C gnd NAND2X1_410/A vdd NAND3X1
XNAND3X1_286 NAND3X1_286/A NAND3X1_287/B NAND3X1_287/C gnd NAND3X1_286/Y vdd NAND3X1
XFILL_21_1_2 gnd vdd FILL
XNAND2X1_400 INVX1_305/A NAND3X1_281/Y gnd NAND2X1_400/Y vdd NAND2X1
XNAND2X1_411 NAND2X1_391/A NAND3X1_279/C gnd INVX1_303/A vdd NAND2X1
XNAND2X1_422 AND2X2_48/B AND2X2_48/A gnd XNOR2X1_49/A vdd NAND2X1
XNAND2X1_433 OAI21X1_380/Y NAND3X1_346/Y gnd NOR2X1_225/A vdd NAND2X1
XNAND2X1_444 NAND2X1_444/A NAND3X1_364/Y gnd NAND2X1_444/Y vdd NAND2X1
XFILL_4_2_2 gnd vdd FILL
XFILL_12_1_2 gnd vdd FILL
XOAI21X1_43 OAI21X1_42/Y AOI21X1_6/Y AOI21X1_7/Y gnd AND2X2_7/A vdd OAI21X1
XOAI21X1_32 INVX1_36/Y INVX1_37/Y NAND2X1_18/Y gnd XNOR2X1_7/A vdd OAI21X1
XOAI21X1_21 BUFX4_8/Y INVX1_28/Y OAI21X1_21/C gnd OAI21X1_21/Y vdd OAI21X1
XOAI21X1_87 OAI21X1_87/A OR2X2_4/Y OAI21X1_87/C gnd OAI21X1_87/Y vdd OAI21X1
XOAI21X1_76 INVX1_24/A NOR2X1_58/B INVX2_2/A gnd NAND2X1_45/A vdd OAI21X1
XOAI21X1_10 NOR2X1_3/Y AND2X2_1/A INVX1_17/Y gnd XNOR2X1_4/A vdd OAI21X1
XOAI21X1_54 BUFX4_6/Y INVX1_69/Y NAND2X1_33/Y gnd OAI21X1_54/Y vdd OAI21X1
XOAI21X1_65 BUFX4_16/Y XOR2X1_3/Y NAND2X1_37/Y gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_98 BUFX4_7/Y INVX1_100/Y OAI21X1_98/C gnd OAI21X1_98/Y vdd OAI21X1
XAND2X2_13 AND2X2_13/A INVX2_5/Y gnd AND2X2_13/Y vdd AND2X2
XOAI21X1_268 AOI21X1_92/Y AOI21X1_93/Y XOR2X1_16/Y gnd AOI21X1_95/A vdd OAI21X1
XOAI21X1_213 NOR3X1_5/Y AOI21X1_64/Y NAND3X1_66/C gnd AOI21X1_66/B vdd OAI21X1
XOAI21X1_279 INVX2_29/A INVX2_33/A INVX2_28/A gnd NOR2X1_172/A vdd OAI21X1
XOAI21X1_202 AOI22X1_11/Y AOI22X1_12/Y NAND3X1_60/B gnd NAND3X1_59/A vdd OAI21X1
XOAI21X1_235 INVX2_24/Y INVX1_203/Y OAI21X1_235/C gnd NAND3X1_89/B vdd OAI21X1
XOAI21X1_257 INVX2_25/A NOR2X1_154/Y INVX2_23/A gnd OAI21X1_258/B vdd OAI21X1
XOAI21X1_246 INVX2_25/A NOR2X1_154/Y NAND3X1_99/B gnd AOI22X1_23/B vdd OAI21X1
XOAI21X1_224 INVX2_19/A INVX1_189/Y INVX1_192/A gnd NAND3X1_82/A vdd OAI21X1
XAND2X2_46 INVX2_36/A INVX1_99/A gnd AND2X2_46/Y vdd AND2X2
XAND2X2_35 INVX1_234/Y AND2X2_35/B gnd AND2X2_35/Y vdd AND2X2
XNAND2X1_241 INVX1_104/A INVX1_103/A gnd NAND2X1_242/B vdd NAND2X1
XNAND2X1_230 NAND3X1_86/Y AOI22X1_20/A gnd OAI21X1_242/A vdd NAND2X1
XAND2X2_24 AND2X2_24/A AND2X2_24/B gnd XOR2X1_9/A vdd AND2X2
XNAND2X1_252 OAI21X1_274/C AOI21X1_84/A gnd XNOR2X1_35/A vdd NAND2X1
XNAND2X1_263 NAND2X1_263/A NAND2X1_263/B gnd NAND3X1_159/B vdd NAND2X1
XNAND2X1_296 gnd gnd gnd INVX1_237/A vdd NAND2X1
XNAND2X1_285 INVX2_28/A INVX1_131/A gnd NOR2X1_183/A vdd NAND2X1
XNAND2X1_274 NAND3X1_149/B NAND3X1_149/C gnd NAND2X1_274/Y vdd NAND2X1
XCLKBUF1_11 clk gnd DFFSR_1/CLK vdd CLKBUF1
XFILL_1_0_2 gnd vdd FILL
XINVX1_118 INVX1_118/A gnd INVX1_118/Y vdd INVX1
XINVX1_107 INVX1_107/A gnd INVX1_107/Y vdd INVX1
XINVX1_129 INVX1_129/A gnd INVX1_129/Y vdd INVX1
XFILL_9_1_2 gnd vdd FILL
XFILL_17_0_2 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XNOR2X1_24 NOR2X1_22/Y INVX1_42/A gnd AND2X2_2/B vdd NOR2X1
XNOR2X1_46 NOR2X1_46/A NOR2X1_45/Y gnd NOR2X1_46/Y vdd NOR2X1
XNOR2X1_13 INVX1_79/A NOR2X1_13/B gnd NOR2X1_13/Y vdd NOR2X1
XNAND3X1_79 AND2X2_26/Y NAND3X1_79/B OR2X2_15/Y gnd INVX1_198/A vdd NAND3X1
XNAND3X1_46 INVX1_161/A NAND3X1_49/B NAND3X1_49/C gnd NAND3X1_52/C vdd NAND3X1
XNAND3X1_57 INVX1_182/Y NAND3X1_57/B NAND3X1_57/C gnd AND2X2_25/A vdd NAND3X1
XNAND3X1_24 OR2X2_10/Y NAND3X1_22/Y NAND3X1_23/Y gnd NAND3X1_24/Y vdd NAND3X1
XNAND3X1_35 INVX1_169/A INVX1_171/Y XNOR2X1_23/Y gnd NAND3X1_36/C vdd NAND3X1
XNAND3X1_13 gnd gnd NAND3X1_13/C gnd NAND3X1_13/Y vdd NAND3X1
XNAND3X1_68 NAND3X1_68/A INVX2_14/Y NAND3X1_48/B gnd NAND3X1_69/B vdd NAND3X1
XNOR2X1_35 BUFX4_9/Y INVX1_55/Y gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_57 INVX1_20/A OR2X2_3/Y gnd NAND3X1_7/C vdd NOR2X1
XNOR2X1_68 INVX1_52/Y INVX1_82/Y gnd NOR2X1_68/Y vdd NOR2X1
XNOR2X1_79 NOR2X1_85/A AND2X2_14/A gnd NOR2X1_79/Y vdd NOR2X1
XNOR2X1_103 NOR2X1_102/Y NOR2X1_101/Y gnd NOR2X1_103/Y vdd NOR2X1
XNOR2X1_158 AND2X2_29/Y AND2X2_30/Y gnd NOR2X1_158/Y vdd NOR2X1
XNOR2X1_125 OR2X2_13/B OR2X2_13/A gnd NOR2X1_125/Y vdd NOR2X1
XNOR2X1_147 INVX1_207/A NOR2X1_147/B gnd OR2X2_17/A vdd NOR2X1
XNOR2X1_114 INVX1_145/A INVX1_146/A gnd NAND3X1_68/A vdd NOR2X1
XNOR2X1_136 INVX2_17/Y INVX2_21/Y gnd INVX2_22/A vdd NOR2X1
XFILL_23_2 gnd vdd FILL
XFILL_16_1 gnd vdd FILL
XNOR2X1_169 INVX2_27/Y INVX2_32/Y gnd INVX1_229/A vdd NOR2X1
XDFFSR_1 DFFSR_1/Q DFFSR_1/CLK DFFSR_1/R vdd OR2X2_7/Y gnd vdd DFFSR
XINVX1_49 x2[6] gnd INVX1_49/Y vdd INVX1
XINVX1_38 x0[3] gnd INVX1_38/Y vdd INVX1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XINVX1_290 INVX1_290/A gnd INVX1_290/Y vdd INVX1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XNAND2X1_90 NAND2X1_90/A BUFX4_10/Y gnd NAND2X1_90/Y vdd NAND2X1
XFILL_7_2_0 gnd vdd FILL
XNAND3X1_287 NAND3X1_287/A NAND3X1_287/B NAND3X1_287/C gnd NAND3X1_289/A vdd NAND3X1
XNAND3X1_276 INVX1_284/A AOI21X1_141/C AOI21X1_140/B gnd NAND3X1_276/Y vdd NAND3X1
XNAND3X1_298 INVX2_44/Y NAND3X1_298/B NAND3X1_298/C gnd AOI21X1_152/A vdd NAND3X1
XFILL_15_1_0 gnd vdd FILL
XNAND3X1_210 NAND3X1_201/Y NAND3X1_202/Y INVX1_259/Y gnd NAND3X1_215/B vdd NAND3X1
XNAND3X1_243 NAND3X1_203/Y NAND2X1_348/Y NAND3X1_245/C gnd NAND3X1_243/Y vdd NAND3X1
XNAND3X1_232 NAND3X1_232/A NAND3X1_232/B OR2X2_24/Y gnd NAND3X1_232/Y vdd NAND3X1
XNAND3X1_254 AOI22X1_36/D AOI22X1_36/C INVX1_271/Y gnd NAND3X1_255/C vdd NAND3X1
XNAND3X1_265 AOI21X1_130/Y NAND3X1_257/B NAND3X1_257/C gnd AOI22X1_38/A vdd NAND3X1
XNAND3X1_221 INVX1_263/A NAND3X1_217/Y NAND3X1_221/C gnd NAND3X1_228/A vdd NAND3X1
XNAND2X1_423 NAND3X1_326/Y OAI21X1_370/Y gnd NAND2X1_423/Y vdd NAND2X1
XNAND2X1_401 NAND2X1_401/A OR2X2_34/B gnd INVX1_295/A vdd NAND2X1
XNAND2X1_412 INVX1_95/A INVX1_97/A gnd INVX2_44/A vdd NAND2X1
XNAND2X1_445 NAND3X1_362/Y NAND2X1_445/B gnd NAND2X1_445/Y vdd NAND2X1
XNAND2X1_434 NOR2X1_225/A XNOR2X1_51/Y gnd NAND2X1_434/Y vdd NAND2X1
XOAI21X1_11 BUFX4_16/Y XNOR2X1_4/Y OAI21X1_11/C gnd OAI21X1_11/Y vdd OAI21X1
XOAI21X1_44 INVX1_61/Y x2[5] NAND3X1_2/Y gnd OAI21X1_44/Y vdd OAI21X1
XOAI21X1_66 NOR2X1_9/A NOR2X1_8/Y INVX1_77/A gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_77 OR2X2_4/B NAND2X1_45/Y OAI21X1_77/C gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_22 BUFX4_8/Y INVX2_4/Y OAI21X1_21/C gnd OAI21X1_22/Y vdd OAI21X1
XOAI21X1_33 BUFX4_16/Y XNOR2X1_7/Y NAND2X1_22/Y gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_88 BUFX4_6/Y INVX1_92/Y OAI21X1_88/C gnd OAI21X1_89/C vdd OAI21X1
XOAI21X1_55 BUFX4_1/Y INVX1_70/Y NAND2X1_33/Y gnd OAI21X1_55/Y vdd OAI21X1
XOAI21X1_99 BUFX4_4/Y INVX1_101/Y OAI21X1_91/C gnd DFFPOSX1_9/D vdd OAI21X1
XOAI21X1_203 INVX1_180/A AND2X2_22/Y gnd gnd NOR2X1_123/B vdd OAI21X1
XAND2X2_47 INVX2_37/A INVX1_98/A gnd AND2X2_47/Y vdd AND2X2
XAND2X2_36 AND2X2_36/A AND2X2_36/B gnd AND2X2_36/Y vdd AND2X2
XAND2X2_25 AND2X2_25/A AND2X2_25/B gnd AND2X2_25/Y vdd AND2X2
XOAI21X1_269 INVX1_211/Y AOI21X1_78/Y NAND3X1_105/Y gnd INVX1_225/A vdd OAI21X1
XOAI21X1_247 NOR3X1_7/Y AOI21X1_78/Y INVX1_211/A gnd NAND2X1_238/B vdd OAI21X1
XOAI21X1_214 AOI22X1_15/Y AOI21X1_66/Y INVX1_185/A gnd NAND3X1_73/B vdd OAI21X1
XOAI21X1_258 INVX2_21/Y OAI21X1_258/B AOI21X1_78/B gnd XOR2X1_14/B vdd OAI21X1
XAND2X2_14 AND2X2_14/A NOR2X1_85/A gnd AND2X2_14/Y vdd AND2X2
XOAI21X1_236 AOI22X1_17/Y AOI22X1_18/Y OAI21X1_229/Y gnd INVX1_219/A vdd OAI21X1
XOAI21X1_225 INVX2_17/Y INVX1_193/Y NAND2X1_199/Y gnd NAND2X1_200/B vdd OAI21X1
XNAND2X1_264 AOI21X1_92/A AOI21X1_92/B gnd AOI21X1_93/C vdd NAND2X1
XNAND2X1_242 NOR2X1_148/B NAND2X1_242/B gnd AOI22X1_25/D vdd NAND2X1
XNAND2X1_286 OAI21X1_283/Y NAND3X1_180/Y gnd NAND2X1_286/Y vdd NAND2X1
XNAND2X1_275 NAND3X1_172/Y NAND3X1_173/Y gnd NAND2X1_275/Y vdd NAND2X1
XNAND2X1_253 INVX2_19/A INVX1_107/A gnd XOR2X1_15/A vdd NAND2X1
XNAND2X1_231 INVX1_218/A AOI22X1_18/A gnd OAI21X1_242/B vdd NAND2X1
XNAND2X1_220 NAND3X1_89/B NAND3X1_87/Y gnd NAND2X1_221/B vdd NAND2X1
XFILL_4_0_0 gnd vdd FILL
XNAND2X1_297 gnd gnd gnd INVX1_238/A vdd NAND2X1
XINVX1_119 INVX1_153/A gnd AOI22X1_2/B vdd INVX1
XINVX1_108 INVX1_108/A gnd INVX1_108/Y vdd INVX1
XFILL_4_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XNAND3X1_14 INVX1_138/Y NAND3X1_14/B OR2X2_8/Y gnd NAND3X1_14/Y vdd NAND3X1
XNOR2X1_25 x0[4] x2[4] gnd NOR2X1_25/Y vdd NOR2X1
XNOR2X1_14 x1[7] INVX1_22/Y gnd NOR2X1_14/Y vdd NOR2X1
XNOR2X1_47 INVX2_1/Y INVX1_21/Y gnd INVX1_81/A vdd NOR2X1
XNOR2X1_58 INVX1_24/A NOR2X1_58/B gnd NOR2X1_58/Y vdd NOR2X1
XNAND3X1_58 XOR2X1_11/Y NAND3X1_58/B NAND3X1_58/C gnd AND2X2_25/B vdd NAND3X1
XNAND3X1_47 INVX1_175/A NAND3X1_43/Y NAND3X1_52/C gnd INVX1_185/A vdd NAND3X1
XNAND3X1_36 NAND3X1_36/A INVX1_178/A NAND3X1_36/C gnd NAND3X1_36/Y vdd NAND3X1
XNAND3X1_25 NAND3X1_25/A OAI22X1_7/Y OAI22X1_8/Y gnd NAND3X1_25/Y vdd NAND3X1
XNAND3X1_69 NAND3X1_69/A NAND3X1_69/B NAND3X1_43/Y gnd NAND3X1_69/Y vdd NAND3X1
XNOR2X1_36 BUFX4_5/Y INVX1_56/Y gnd NOR2X1_36/Y vdd NOR2X1
XNOR2X1_69 NOR2X1_69/A NOR2X1_68/Y gnd NOR2X1_69/Y vdd NOR2X1
XNOR2X1_104 INVX2_9/A INVX2_10/Y gnd NOR2X1_104/Y vdd NOR2X1
XNOR2X1_159 NOR2X1_159/A NOR2X1_159/B gnd AOI21X1_89/C vdd NOR2X1
XNOR2X1_126 INVX1_181/Y NOR2X1_125/Y gnd OAI22X1_16/C vdd NOR2X1
XNOR2X1_148 INVX1_192/A NOR2X1_148/B gnd NOR2X1_148/Y vdd NOR2X1
XNOR2X1_115 INVX1_145/Y INVX1_146/Y gnd NOR2X1_115/Y vdd NOR2X1
XNOR2X1_137 INVX2_17/Y INVX2_23/Y gnd INVX1_188/A vdd NOR2X1
XFILL_23_3 gnd vdd FILL
XINVX1_280 INVX1_280/A gnd INVX1_280/Y vdd INVX1
XINVX1_291 INVX1_97/A gnd INVX1_291/Y vdd INVX1
XINVX1_39 x2[3] gnd INVX1_39/Y vdd INVX1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XINVX1_17 NOR2X1_4/Y gnd INVX1_17/Y vdd INVX1
XNAND2X1_80 INVX1_114/A INVX1_113/Y gnd NAND2X1_80/Y vdd NAND2X1
XNAND2X1_91 INVX2_16/A BUFX4_10/Y gnd NAND2X1_91/Y vdd NAND2X1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XNAND3X1_277 OR2X2_31/B NAND3X1_277/B OR2X2_30/Y gnd AOI22X1_46/B vdd NAND3X1
XNAND3X1_288 NAND3X1_286/A NAND3X1_281/Y NAND3X1_282/Y gnd NAND3X1_289/B vdd NAND3X1
XNAND3X1_299 INVX2_36/A INVX1_99/A NOR2X1_224/B gnd NAND3X1_301/B vdd NAND3X1
XNAND3X1_200 INVX1_254/Y NAND3X1_199/Y OAI21X1_304/Y gnd NAND2X1_326/A vdd NAND3X1
XNAND3X1_244 NAND3X1_243/Y NAND2X1_345/Y NAND2X1_352/Y gnd NAND3X1_244/Y vdd NAND3X1
XNAND3X1_233 INVX1_247/A NAND3X1_233/B NAND3X1_232/Y gnd NAND3X1_234/C vdd NAND3X1
XNAND3X1_266 NAND2X1_317/Y INVX1_246/A NAND2X1_359/Y gnd AOI22X1_41/C vdd NAND3X1
XNAND3X1_222 INVX1_262/A NAND3X1_213/Y NAND3X1_216/Y gnd NAND3X1_224/B vdd NAND3X1
XNAND3X1_255 INVX1_270/Y NAND3X1_255/B NAND3X1_255/C gnd NAND3X1_255/Y vdd NAND3X1
XNAND3X1_211 INVX1_259/A NAND3X1_204/Y NAND3X1_205/Y gnd NAND3X1_211/Y vdd NAND3X1
XNAND2X1_402 AOI22X1_46/B AOI22X1_46/A gnd OAI21X1_358/A vdd NAND2X1
XNAND2X1_446 NAND3X1_276/Y OAI21X1_344/Y gnd NOR2X1_227/B vdd NAND2X1
XNAND2X1_413 INVX1_96/A INVX1_95/A gnd NAND2X1_413/Y vdd NAND2X1
XNAND2X1_424 OAI21X1_391/C NAND2X1_424/B gnd XNOR2X1_50/A vdd NAND2X1
XNAND2X1_435 OAI21X1_382/Y NAND2X1_435/B gnd NAND3X1_352/A vdd NAND2X1
XOAI21X1_45 NOR2X1_25/Y INVX1_46/A INVX1_60/Y gnd INVX1_62/A vdd OAI21X1
XOAI21X1_34 INVX1_40/A INVX1_42/Y OAI21X1_34/C gnd AOI21X1_4/C vdd OAI21X1
XOAI21X1_23 BUFX4_8/Y INVX1_29/Y OAI21X1_21/C gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_12 NAND2X1_11/Y AND2X2_1/A AOI21X1_3/Y gnd NOR2X1_13/B vdd OAI21X1
XOAI21X1_67 INVX1_19/Y INVX1_18/Y OAI21X1_66/Y gnd NOR2X1_46/A vdd OAI21X1
XOAI21X1_78 INVX2_3/A NAND2X1_45/B BUFX4_6/Y gnd OAI21X1_78/Y vdd OAI21X1
XOAI21X1_89 BUFX4_14/Y OR2X2_4/A OAI21X1_89/C gnd OAI21X1_89/Y vdd OAI21X1
XOAI21X1_56 BUFX4_4/Y INVX1_71/Y NAND2X1_33/Y gnd OAI21X1_56/Y vdd OAI21X1
XOAI21X1_215 AOI21X1_67/Y AOI21X1_68/Y NAND3X1_51/Y gnd NAND3X1_75/C vdd OAI21X1
XOAI21X1_204 INVX2_12/Y AND2X2_22/Y INVX1_180/Y gnd INVX1_181/A vdd OAI21X1
XOAI21X1_237 AOI22X1_20/Y NOR2X1_156/B AOI21X1_75/Y gnd NAND3X1_93/C vdd OAI21X1
XOAI21X1_226 INVX2_17/Y INVX1_193/Y NOR2X1_143/Y gnd NAND2X1_201/A vdd OAI21X1
XAND2X2_48 AND2X2_48/A AND2X2_48/B gnd AND2X2_48/Y vdd AND2X2
XAND2X2_15 INVX1_124/Y AND2X2_15/B gnd INVX2_7/A vdd AND2X2
XOAI21X1_259 NOR2X1_159/B INVX1_214/A INVX1_215/A gnd INVX1_221/A vdd OAI21X1
XOAI21X1_248 NOR3X1_7/B NOR3X1_7/C NOR3X1_7/A gnd OAI21X1_248/Y vdd OAI21X1
XAND2X2_37 INVX2_28/A OR2X2_6/B gnd AND2X2_37/Y vdd AND2X2
XAND2X2_26 AND2X2_26/A AND2X2_26/B gnd AND2X2_26/Y vdd AND2X2
XNAND2X1_265 AND2X2_32/B AND2X2_32/A gnd NAND3X1_161/C vdd NAND2X1
XNAND2X1_298 OR2X2_23/B OR2X2_23/A gnd NAND2X1_299/A vdd NAND2X1
XFILL_4_0_1 gnd vdd FILL
XNAND2X1_243 INVX2_18/A INVX1_106/A gnd INVX1_212/A vdd NAND2X1
XNAND2X1_287 NAND2X1_287/A NAND2X1_287/B gnd OR2X2_22/A vdd NAND2X1
XNAND2X1_221 INVX1_202/A NAND2X1_221/B gnd AOI22X1_17/D vdd NAND2X1
XNAND2X1_232 INVX1_187/A AOI22X1_21/D gnd OR2X2_19/A vdd NAND2X1
XNAND2X1_254 INVX2_18/A INVX1_108/A gnd XOR2X1_15/B vdd NAND2X1
XNAND2X1_276 NAND3X1_171/Y NAND3X1_175/Y gnd NAND2X1_276/Y vdd NAND2X1
XNAND2X1_210 INVX1_187/A INVX1_193/A gnd INVX1_200/A vdd NAND2X1
XINVX1_109 INVX1_109/A gnd NOR2X1_65/B vdd INVX1
XFILL_4_2 gnd vdd FILL
XFILL_10_2_2 gnd vdd FILL
XNAND3X1_48 INVX1_161/A NAND3X1_48/B NAND3X1_48/C gnd NAND3X1_48/Y vdd NAND3X1
XNAND3X1_15 INVX1_135/Y NAND3X1_15/B OR2X2_9/Y gnd INVX1_140/A vdd NAND3X1
XNAND3X1_37 INVX1_169/A INVX1_171/Y XOR2X1_7/Y gnd NAND3X1_37/Y vdd NAND3X1
XNAND3X1_26 NAND3X1_22/A OAI22X1_10/Y OAI22X1_9/Y gnd NAND3X1_26/Y vdd NAND3X1
XNOR2X1_26 INVX1_43/Y INVX1_44/Y gnd INVX1_46/A vdd NOR2X1
XNOR2X1_15 x3[7] INVX1_23/Y gnd NOR2X1_17/A vdd NOR2X1
XNOR2X1_48 NOR2X1_48/A OAI22X1_6/C gnd NOR2X1_48/Y vdd NOR2X1
XNOR2X1_59 INVX2_3/Y AND2X2_10/Y gnd NOR2X1_59/Y vdd NOR2X1
XNAND3X1_59 NAND3X1_59/A NAND3X1_56/Y AND2X2_25/Y gnd NAND3X1_59/Y vdd NAND3X1
XNOR2X1_37 BUFX4_5/Y INVX1_57/Y gnd NOR2X1_37/Y vdd NOR2X1
XNOR2X1_138 INVX2_20/Y INVX2_22/Y gnd NAND3X1_78/B vdd NOR2X1
XNOR2X1_105 INVX2_8/Y INVX1_134/Y gnd NOR2X1_105/Y vdd NOR2X1
XNOR2X1_127 NOR2X1_123/Y NOR3X1_2/C gnd NOR2X1_127/Y vdd NOR2X1
XNOR2X1_149 INVX1_203/Y INVX2_24/Y gnd NOR2X1_149/Y vdd NOR2X1
XNOR2X1_116 NAND3X1_68/A NOR2X1_115/Y gnd NOR2X1_116/Y vdd NOR2X1
XINVX1_18 x3[5] gnd INVX1_18/Y vdd INVX1
XINVX1_281 INVX1_281/A gnd INVX1_281/Y vdd INVX1
XINVX1_292 OR2X2_29/Y gnd INVX1_292/Y vdd INVX1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XINVX1_270 INVX1_270/A gnd INVX1_270/Y vdd INVX1
XNAND2X1_70 INVX1_75/A INVX1_41/Y gnd NAND2X1_71/B vdd NAND2X1
XNAND2X1_81 INVX1_113/A INVX1_114/Y gnd NAND2X1_81/Y vdd NAND2X1
XNAND2X1_92 AND2X2_16/B INVX2_6/A gnd INVX1_125/A vdd NAND2X1
XFILL_7_2_2 gnd vdd FILL
XFILL_15_1_2 gnd vdd FILL
XNAND3X1_223 INVX1_262/Y NAND3X1_218/Y NAND3X1_219/Y gnd NAND3X1_224/C vdd NAND3X1
XNAND3X1_212 NAND2X1_333/Y NAND3X1_211/Y NAND3X1_215/B gnd NAND3X1_212/Y vdd NAND3X1
XNAND3X1_201 INVX1_257/Y OAI21X1_306/Y OAI21X1_320/C gnd NAND3X1_201/Y vdd NAND3X1
XNAND3X1_289 NAND3X1_289/A NAND3X1_289/B XOR2X1_21/B gnd NAND3X1_289/Y vdd NAND3X1
XNAND3X1_278 NAND2X1_391/A NAND3X1_278/B NOR2X1_216/Y gnd NAND3X1_279/C vdd NAND3X1
XNAND3X1_267 INVX2_35/A INVX1_273/A INVX2_38/Y gnd INVX1_272/A vdd NAND3X1
XNAND3X1_234 NAND2X1_317/Y NAND3X1_234/B NAND3X1_234/C gnd NAND3X1_234/Y vdd NAND3X1
XNAND3X1_256 OAI21X1_322/Y NAND3X1_255/Y XNOR2X1_44/Y gnd NAND3X1_257/C vdd NAND3X1
XNAND3X1_245 NAND3X1_203/Y NAND2X1_351/Y NAND3X1_245/C gnd NAND3X1_245/Y vdd NAND3X1
XFILL_21_1 gnd vdd FILL
XNAND2X1_403 INVX1_304/A AOI22X1_46/D gnd NAND2X1_403/Y vdd NAND2X1
XNAND2X1_414 NOR2X1_215/B NAND2X1_413/Y gnd AOI22X1_51/D vdd NAND2X1
XNAND2X1_425 INVX2_37/A INVX1_99/A gnd XOR2X1_23/A vdd NAND2X1
XNAND2X1_436 NAND2X1_436/A NAND2X1_436/B gnd NAND3X1_353/C vdd NAND2X1
XOAI21X1_46 OAI21X1_44/Y AND2X2_7/Y INVX1_50/A gnd OAI21X1_46/Y vdd OAI21X1
XOAI21X1_13 INVX2_1/Y x3[6] OAI21X1_13/C gnd XNOR2X1_5/A vdd OAI21X1
XOAI21X1_68 NOR2X1_9/A NOR2X1_8/Y INVX1_15/Y gnd NOR2X1_45/A vdd OAI21X1
XOAI21X1_35 INVX1_45/Y AND2X2_3/A BUFX4_3/Y gnd OAI22X1_3/D vdd OAI21X1
XOAI21X1_57 BUFX4_2/Y INVX1_72/Y OAI21X1_1/Y gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_24 BUFX4_6/Y INVX1_30/Y OAI21X1_21/C gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_79 OAI21X1_78/Y NOR2X1_59/Y OAI21X1_79/C gnd OAI21X1_79/Y vdd OAI21X1
XOAI21X1_249 INVX1_205/A INVX2_26/A AOI22X1_25/D gnd XNOR2X1_32/A vdd OAI21X1
XOAI21X1_205 NOR2X1_128/Y OAI22X1_17/C NOR2X1_127/Y gnd NAND3X1_57/C vdd OAI21X1
XOAI21X1_216 AOI22X1_15/Y AOI21X1_66/Y INVX1_185/Y gnd NAND3X1_75/A vdd OAI21X1
XOAI21X1_238 AOI22X1_17/Y AOI22X1_18/Y AOI21X1_75/Y gnd NAND3X1_91/B vdd OAI21X1
XOAI21X1_227 INVX2_21/Y INVX1_187/A NOR2X1_142/Y gnd OAI21X1_227/Y vdd OAI21X1
XDFFPOSX1_130 BUFX2_26/A CLKBUF1_6/Y NOR2X1_199/Y gnd vdd DFFPOSX1
XAND2X2_38 INVX2_29/A AND2X2_38/B gnd AND2X2_38/Y vdd AND2X2
XNAND2X1_211 INVX2_17/A AOI22X1_21/D gnd INVX1_201/A vdd NAND2X1
XNAND2X1_200 NAND3X1_82/Y NAND2X1_200/B gnd OR2X2_16/A vdd NAND2X1
XAND2X2_16 AND2X2_16/A AND2X2_16/B gnd AND2X2_16/Y vdd AND2X2
XAND2X2_27 AND2X2_27/A INVX1_198/Y gnd AND2X2_27/Y vdd AND2X2
XNAND2X1_277 NAND3X1_85/Y AOI21X1_73/A gnd NOR2X1_161/B vdd NAND2X1
XNAND2X1_266 OAI21X1_266/Y AND2X2_32/Y gnd AOI21X1_93/B vdd NAND2X1
XNAND2X1_299 NAND2X1_299/A OR2X2_23/Y gnd INVX1_239/A vdd NAND2X1
XNAND2X1_244 AND2X2_29/Y AND2X2_30/Y gnd NAND2X1_244/Y vdd NAND2X1
XFILL_4_0_2 gnd vdd FILL
XNAND2X1_288 OR2X2_22/B OR2X2_22/A gnd AND2X2_34/B vdd NAND2X1
XNAND2X1_255 INVX2_17/A INVX1_129/A gnd XOR2X1_16/B vdd NAND2X1
XNAND2X1_233 INVX2_21/A INVX1_193/A gnd OR2X2_19/B vdd NAND2X1
XNAND2X1_222 OR2X2_18/B OR2X2_18/A gnd AOI22X1_19/C vdd NAND2X1
XFILL_22_2_0 gnd vdd FILL
XFILL_13_2_0 gnd vdd FILL
XNAND3X1_16 OR2X2_9/Y INVX2_11/A OR2X2_11/Y gnd NAND3X1_16/Y vdd NAND3X1
XNAND3X1_27 INVX1_159/Y NAND3X1_26/Y NAND3X1_25/Y gnd NAND3X1_27/Y vdd NAND3X1
XNAND3X1_38 NAND3X1_40/B NAND3X1_37/Y AND2X2_23/Y gnd AOI21X1_57/A vdd NAND3X1
XNAND3X1_49 INVX1_161/Y NAND3X1_49/B NAND3X1_49/C gnd NAND3X1_49/Y vdd NAND3X1
XNOR2X1_16 NOR2X1_14/Y NOR2X1_17/A gnd INVX1_25/A vdd NOR2X1
XNOR2X1_27 NOR2X1_25/Y INVX1_46/A gnd INVX1_45/A vdd NOR2X1
XNOR2X1_38 BUFX4_7/Y INVX1_58/Y gnd NOR2X1_38/Y vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_49 BUFX4_9/Y INVX1_83/Y gnd NOR2X1_49/Y vdd NOR2X1
XFILL_10_0_0 gnd vdd FILL
XFILL_18_1_0 gnd vdd FILL
XNOR2X1_106 INVX2_10/Y INVX1_139/Y gnd INVX1_141/A vdd NOR2X1
XNOR2X1_117 NOR2X1_112/Y INVX2_11/Y gnd AOI22X1_6/D vdd NOR2X1
XNOR2X1_128 INVX1_181/Y OR2X2_13/Y gnd NOR2X1_128/Y vdd NOR2X1
XNOR2X1_139 INVX2_19/Y INVX1_189/Y gnd NOR2X1_140/B vdd NOR2X1
XINVX1_19 x1[5] gnd INVX1_19/Y vdd INVX1
XINVX1_282 INVX1_282/A gnd INVX1_282/Y vdd INVX1
XINVX1_293 INVX1_293/A gnd INVX1_293/Y vdd INVX1
XINVX1_271 INVX1_271/A gnd INVX1_271/Y vdd INVX1
XINVX1_260 INVX1_260/A gnd INVX1_260/Y vdd INVX1
XNAND2X1_71 NAND2X1_69/Y NAND2X1_71/B gnd INVX1_115/A vdd NAND2X1
XNAND2X1_60 BUFX4_1/Y INVX1_70/A gnd NAND2X1_60/Y vdd NAND2X1
XNAND2X1_82 NAND2X1_80/Y NAND2X1_81/Y gnd NAND3X1_12/B vdd NAND2X1
XNAND2X1_93 INVX1_88/A INVX1_59/Y gnd AND2X2_15/B vdd NAND2X1
XNAND3X1_213 XNOR2X1_39/Y NAND3X1_212/Y NAND3X1_245/C gnd NAND3X1_213/Y vdd NAND3X1
XNAND3X1_246 NAND3X1_245/Y NAND2X1_353/Y AND2X2_41/Y gnd NAND3X1_246/Y vdd NAND3X1
XNAND3X1_224 INVX1_263/Y NAND3X1_224/B NAND3X1_224/C gnd NAND3X1_228/B vdd NAND3X1
XNAND3X1_257 OAI21X1_313/Y NAND3X1_257/B NAND3X1_257/C gnd AOI22X1_37/A vdd NAND3X1
XNAND3X1_235 INVX1_247/A NAND3X1_230/B NAND3X1_230/C gnd NAND3X1_237/B vdd NAND3X1
XNAND3X1_202 INVX1_257/A NAND2X1_332/Y OAI21X1_307/Y gnd NAND3X1_202/Y vdd NAND3X1
XNAND3X1_279 INVX1_288/Y NAND3X1_279/B NAND3X1_279/C gnd AOI22X1_43/C vdd NAND3X1
XNAND3X1_268 INVX1_273/A INVX2_41/A INVX2_40/A gnd NOR2X1_211/A vdd NAND3X1
XFILL_14_1 gnd vdd FILL
XNAND2X1_404 INVX1_273/A AOI22X1_47/D gnd OR2X2_32/A vdd NAND2X1
XNAND2X1_415 INVX2_36/A INVX1_98/A gnd INVX1_298/A vdd NAND2X1
XNAND2X1_437 NAND3X1_356/A NAND3X1_356/C gnd NAND2X1_437/Y vdd NAND2X1
XNAND2X1_426 INVX2_36/A INVX1_100/A gnd XOR2X1_23/B vdd NAND2X1
XINVX2_40 INVX2_40/A gnd INVX2_40/Y vdd INVX2
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_14 BUFX4_14/Y XNOR2X1_5/Y OAI21X1_14/C gnd OAI21X1_14/Y vdd OAI21X1
XOAI21X1_47 INVX1_48/Y x2[6] OAI21X1_46/Y gnd OAI21X1_47/Y vdd OAI21X1
XOAI21X1_36 NOR2X1_25/Y AND2X2_3/A INVX1_46/Y gnd XNOR2X1_8/A vdd OAI21X1
XOAI21X1_58 INVX1_3/Y INVX1_2/Y XNOR2X1_1/Y gnd NAND3X1_4/C vdd OAI21X1
XOAI21X1_69 NOR2X1_46/A NOR2X1_45/Y INVX1_79/Y gnd NAND3X1_6/B vdd OAI21X1
XOAI21X1_25 x0[0] x2[0] BUFX4_2/Y gnd OR2X2_1/B vdd OAI21X1
XOAI21X1_206 INVX1_163/A AND2X2_22/Y INVX1_180/Y gnd XOR2X1_11/A vdd OAI21X1
XOAI21X1_239 AOI22X1_20/Y NOR2X1_156/B OAI21X1_229/Y gnd NAND3X1_91/C vdd OAI21X1
XOAI21X1_228 AOI21X1_76/C AOI21X1_72/Y INVX1_198/Y gnd AOI21X1_73/A vdd OAI21X1
XOAI21X1_217 INVX1_187/Y INVX2_20/Y INVX2_22/Y gnd AND2X2_26/A vdd OAI21X1
XDFFPOSX1_120 BUFX2_16/A DFFSR_1/CLK NAND2X1_276/Y gnd vdd DFFPOSX1
XDFFPOSX1_131 BUFX2_27/A DFFSR_1/CLK XNOR2X1_46/Y gnd vdd DFFPOSX1
XAND2X2_39 AND2X2_39/A AND2X2_39/B gnd AND2X2_39/Y vdd AND2X2
XNAND2X1_223 INVX1_202/Y NAND2X1_221/B gnd AOI22X1_18/A vdd NAND2X1
XNAND2X1_234 INVX2_17/A AND2X2_28/B gnd NAND3X1_99/B vdd NAND2X1
XAND2X2_28 INVX2_17/A AND2X2_28/B gnd AND2X2_28/Y vdd AND2X2
XNAND2X1_212 OR2X2_17/B OR2X2_17/A gnd NAND3X1_86/B vdd NAND2X1
XNAND2X1_201 NAND2X1_201/A OAI21X1_227/Y gnd INVX1_194/A vdd NAND2X1
XAND2X2_17 AND2X2_17/A INVX2_7/Y gnd AND2X2_17/Y vdd AND2X2
XNAND2X1_267 AOI21X1_93/A AOI21X1_93/B gnd AOI21X1_92/C vdd NAND2X1
XNAND2X1_289 NOR2X1_179/A INVX1_233/Y gnd AND2X2_35/B vdd NAND2X1
XNAND2X1_256 AOI21X1_88/A AOI21X1_88/B gnd NOR2X1_157/A vdd NAND2X1
XNAND2X1_245 INVX2_19/A INVX1_106/A gnd NOR2X1_159/B vdd NAND2X1
XNAND2X1_278 gnd INVX2_27/Y gnd XNOR2X1_38/B vdd NAND2X1
XFILL_22_2_1 gnd vdd FILL
XXNOR2X1_1 x1[1] x3[1] gnd XNOR2X1_1/Y vdd XNOR2X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XFILL_13_2_1 gnd vdd FILL
XAND2X2_1 AND2X2_1/A INVX1_15/Y gnd AND2X2_1/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XNOR2X1_17 NOR2X1_17/A NOR2X1_17/B gnd NOR2X1_17/Y vdd NOR2X1
XNOR2X1_28 x0[5] x2[5] gnd NOR2X1_29/A vdd NOR2X1
XNAND3X1_17 AOI22X1_6/C INVX2_11/A OR2X2_11/Y gnd NOR3X1_6/A vdd NAND3X1
XNAND3X1_28 INVX1_159/Y NAND3X1_22/Y NAND3X1_23/Y gnd NAND3X1_28/Y vdd NAND3X1
XNAND3X1_39 INVX1_178/A NAND3X1_36/C AND2X2_23/Y gnd AOI21X1_58/A vdd NAND3X1
XNOR2X1_39 BUFX4_7/Y INVX1_59/Y gnd NOR2X1_39/Y vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XFILL_10_0_1 gnd vdd FILL
XFILL_18_1_1 gnd vdd FILL
XNOR2X1_129 INVX1_181/A NOR2X1_125/Y gnd OAI22X1_17/C vdd NOR2X1
XNOR2X1_118 AND2X2_22/A AND2X2_22/B gnd INVX1_180/A vdd NOR2X1
XNOR2X1_107 NOR2X1_107/A INVX1_141/A gnd NAND3X1_13/C vdd NOR2X1
XINVX1_250 INVX1_250/A gnd INVX1_250/Y vdd INVX1
XINVX1_261 INVX1_261/A gnd INVX1_261/Y vdd INVX1
XNAND2X1_50 AOI22X1_47/D BUFX4_14/Y gnd OAI21X1_86/C vdd NAND2X1
XINVX1_283 INVX1_283/A gnd INVX1_283/Y vdd INVX1
XINVX1_272 INVX1_272/A gnd INVX1_272/Y vdd INVX1
XINVX1_294 INVX1_294/A gnd OR2X2_34/B vdd INVX1
XNAND2X1_61 BUFX4_4/Y INVX1_71/A gnd OAI21X1_98/C vdd NAND2X1
XNAND2X1_83 NAND2X1_75/Y AND2X2_12/Y gnd NOR2X1_71/A vdd NAND2X1
XNAND2X1_72 NAND3X1_8/B INVX1_115/Y gnd NOR2X1_71/B vdd NAND2X1
XNAND2X1_94 XOR2X1_5/Y NAND2X1_94/B gnd AOI22X1_3/C vdd NAND2X1
XNAND3X1_269 NAND3X1_269/A NOR2X1_205/Y NAND2X1_364/Y gnd OAI21X1_339/C vdd NAND3X1
XNAND3X1_203 INVX1_259/A NAND3X1_201/Y NAND3X1_202/Y gnd NAND3X1_203/Y vdd NAND3X1
XNAND3X1_258 OR2X2_25/Y INVX1_249/Y XNOR2X1_44/B gnd NAND3X1_258/Y vdd NAND3X1
XNAND3X1_236 INVX1_247/Y NAND3X1_233/B NAND3X1_232/Y gnd NAND3X1_236/Y vdd NAND3X1
XNAND3X1_247 NAND3X1_244/Y NAND3X1_246/Y OAI21X1_316/Y gnd AOI22X1_36/D vdd NAND3X1
XNAND3X1_225 NAND3X1_228/A NAND3X1_228/B OAI21X1_312/C gnd NAND3X1_225/Y vdd NAND3X1
XNAND3X1_214 NAND2X1_333/Y NAND3X1_203/Y NAND3X1_206/Y gnd NAND3X1_214/Y vdd NAND3X1
XFILL_14_2 gnd vdd FILL
XNAND2X1_405 INVX2_39/A INVX1_279/A gnd OR2X2_32/B vdd NAND2X1
XNAND2X1_416 AND2X2_46/Y AND2X2_47/Y gnd NAND3X1_298/C vdd NAND2X1
XNAND2X1_427 NAND2X1_427/A XOR2X1_23/Y gnd NAND2X1_427/Y vdd NAND2X1
XNAND2X1_438 INVX1_309/Y NAND2X1_437/Y gnd NAND3X1_357/B vdd NAND2X1
XINVX2_41 INVX2_41/A gnd INVX2_41/Y vdd INVX2
XINVX2_30 INVX2_30/A gnd INVX2_30/Y vdd INVX2
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_15 NOR2X1_14/Y INVX1_26/Y BUFX4_8/Y gnd NOR2X1_17/B vdd OAI21X1
XOAI21X1_48 NOR2X1_31/Y INVX1_51/Y OAI21X1_47/Y gnd OAI21X1_48/Y vdd OAI21X1
XOAI21X1_59 BUFX4_2/Y INVX1_73/Y NAND3X1_4/Y gnd OAI21X1_59/Y vdd OAI21X1
XOAI21X1_26 BUFX4_2/Y INVX1_31/Y OR2X2_1/Y gnd OAI21X1_26/Y vdd OAI21X1
XOAI21X1_37 BUFX4_16/Y XNOR2X1_8/Y OAI21X1_37/C gnd OAI21X1_37/Y vdd OAI21X1
XDFFPOSX1_121 BUFX2_17/A CLKBUF1_6/Y NOR2X1_103/Y gnd vdd DFFPOSX1
XOAI21X1_207 NOR2X1_124/Y OAI22X1_16/C NOR2X1_127/Y gnd NAND3X1_58/C vdd OAI21X1
XAND2X2_29 INVX2_18/A INVX1_107/A gnd AND2X2_29/Y vdd AND2X2
XAND2X2_18 AND2X2_18/A OR2X2_6/Y gnd AND2X2_18/Y vdd AND2X2
XOAI21X1_229 INVX1_196/A NAND2X1_207/B OR2X2_16/Y gnd OAI21X1_229/Y vdd OAI21X1
XDFFPOSX1_110 BUFX2_6/A CLKBUF1_3/Y XOR2X1_18/Y gnd vdd DFFPOSX1
XOAI21X1_218 INVX1_187/A INVX2_20/A INVX2_22/A gnd AND2X2_26/B vdd OAI21X1
XDFFPOSX1_132 BUFX2_28/A DFFSR_1/CLK NOR2X1_208/Y gnd vdd DFFPOSX1
XNAND2X1_224 NAND3X1_92/Y NAND3X1_95/Y gnd XOR2X1_13/A vdd NAND2X1
XNAND2X1_268 AOI21X1_95/B AOI21X1_95/A gnd NAND2X1_269/B vdd NAND2X1
XNAND2X1_257 NOR2X1_157/A XNOR2X1_36/Y gnd NAND2X1_257/Y vdd NAND2X1
XNAND2X1_235 AOI22X1_22/B NAND3X1_99/Y gnd NAND3X1_101/C vdd NAND2X1
XNAND2X1_246 INVX2_18/A INVX1_107/A gnd NOR2X1_159/A vdd NAND2X1
XNAND2X1_213 NAND3X1_86/B OR2X2_17/Y gnd OR2X2_18/A vdd NAND2X1
XNAND2X1_202 NAND3X1_77/Y INVX1_194/Y gnd NAND2X1_203/A vdd NAND2X1
XNAND2X1_279 NOR2X1_179/A NAND2X1_279/B gnd OR2X2_21/B vdd NAND2X1
XFILL_22_2_2 gnd vdd FILL
XXNOR2X1_2 OAI21X1_5/Y INVX1_8/Y gnd OAI21X1_6/B vdd XNOR2X1
XFILL_13_2_2 gnd vdd FILL
XINVX1_2 x3[0] gnd INVX1_2/Y vdd INVX1
XAND2X2_2 AND2X2_2/A AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XOAI21X1_390 INVX1_293/Y AOI22X1_46/B OR2X2_34/A gnd OAI21X1_390/Y vdd OAI21X1
XNOR2X1_29 NOR2X1_29/A AND2X2_4/Y gnd INVX1_60/A vdd NOR2X1
XNOR2X1_18 INVX1_32/Y INVX1_33/Y gnd OR2X2_1/A vdd NOR2X1
XNAND3X1_29 OR2X2_10/Y NAND3X1_26/Y NAND3X1_25/Y gnd NAND3X1_29/Y vdd NAND3X1
XNAND3X1_18 INVX1_156/A NAND3X1_21/B NAND3X1_21/C gnd INVX1_149/A vdd NAND3X1
XFILL_2_1_2 gnd vdd FILL
XFILL_10_0_2 gnd vdd FILL
XFILL_18_1_2 gnd vdd FILL
XNOR2X1_108 AOI21X1_42/Y INVX1_140/Y gnd NOR2X1_108/Y vdd NOR2X1
XNOR2X1_119 INVX1_180/A AND2X2_22/Y gnd NOR2X1_119/Y vdd NOR2X1
XINVX1_284 INVX1_284/A gnd AND2X2_44/B vdd INVX1
XINVX1_273 INVX1_273/A gnd INVX1_273/Y vdd INVX1
XINVX1_295 INVX1_295/A gnd INVX1_295/Y vdd INVX1
XINVX1_262 INVX1_262/A gnd INVX1_262/Y vdd INVX1
XINVX1_251 NOR3X1_8/A gnd INVX1_251/Y vdd INVX1
XINVX1_240 INVX1_240/A gnd INVX1_240/Y vdd INVX1
XNAND2X1_51 INVX1_28/Y INVX2_4/Y gnd NOR3X1_1/B vdd NAND2X1
XNAND2X1_62 NOR2X1_64/A INVX1_73/Y gnd NAND2X1_62/Y vdd NAND2X1
XNAND2X1_40 INVX1_12/Y NOR2X1_56/Y gnd OR2X2_3/A vdd NAND2X1
XNAND2X1_73 INVX1_47/Y INVX1_78/Y gnd NAND2X1_75/B vdd NAND2X1
XNAND2X1_95 INVX2_17/A BUFX4_13/Y gnd NAND2X1_95/Y vdd NAND2X1
XNAND2X1_84 INVX2_10/A BUFX4_11/Y gnd NAND2X1_84/Y vdd NAND2X1
XNAND3X1_226 INVX1_254/A NAND3X1_199/Y OAI21X1_304/Y gnd NAND2X1_337/A vdd NAND3X1
XNAND3X1_259 INVX1_267/Y OAI21X1_326/Y NAND3X1_258/Y gnd AND2X2_42/B vdd NAND3X1
XNAND3X1_237 AOI21X1_114/Y NAND3X1_237/B NAND3X1_236/Y gnd NAND3X1_238/C vdd NAND3X1
XNAND3X1_248 NAND3X1_245/Y NAND2X1_345/Y NAND2X1_353/Y gnd NAND3X1_248/Y vdd NAND3X1
XNAND3X1_215 NAND3X1_211/Y NAND3X1_215/B AND2X2_39/Y gnd NAND3X1_215/Y vdd NAND3X1
XNAND3X1_204 INVX1_257/A OAI21X1_306/Y OAI21X1_320/C gnd NAND3X1_204/Y vdd NAND3X1
XNAND2X1_406 INVX2_35/A AND2X2_45/B gnd OAI21X1_362/C vdd NAND2X1
XNAND2X1_417 INVX2_37/A INVX1_98/A gnd NOR2X1_224/B vdd NAND2X1
XNAND2X1_439 INVX1_311/Y XNOR2X1_52/A gnd NAND2X1_441/A vdd NAND2X1
XNAND2X1_428 OAI21X1_376/Y XNOR2X1_51/Y gnd NAND2X1_429/A vdd NAND2X1
XINVX2_42 INVX2_42/A gnd INVX2_42/Y vdd INVX2
XINVX2_31 INVX2_31/A gnd INVX2_31/Y vdd INVX2
XFILL_7_0_2 gnd vdd FILL
XINVX2_20 INVX2_20/A gnd INVX2_20/Y vdd INVX2
XOAI21X1_16 INVX1_25/Y OAI21X1_13/C NOR2X1_17/Y gnd OAI21X1_21/C vdd OAI21X1
XOAI21X1_38 NAND2X1_24/Y AND2X2_3/A AOI21X1_5/Y gnd NOR2X1_30/B vdd OAI21X1
XOAI21X1_27 NOR2X1_21/A AOI21X1_6/C OR2X2_1/A gnd OAI21X1_27/Y vdd OAI21X1
XOAI21X1_49 BUFX4_9/Y INVX1_63/Y NAND2X1_33/Y gnd OAI21X1_49/Y vdd OAI21X1
XOAI21X1_208 AOI22X1_11/Y AOI22X1_12/Y AOI21X1_62/Y gnd NAND3X1_61/A vdd OAI21X1
XOAI21X1_219 INVX1_187/Y INVX2_22/Y INVX1_188/Y gnd NAND2X1_191/B vdd OAI21X1
XDFFPOSX1_100 INVX1_27/A CLKBUF1_1/Y OAI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_111 BUFX2_7/A DFFSR_1/CLK XNOR2X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_122 BUFX2_18/A CLKBUF1_6/Y NOR2X1_101/Y gnd vdd DFFPOSX1
XAND2X2_19 AND2X2_19/A AND2X2_19/B gnd OR2X2_10/A vdd AND2X2
XDFFPOSX1_133 BUFX2_29/A CLKBUF1_6/Y NOR2X1_228/Y gnd vdd DFFPOSX1
XNAND2X1_269 INVX1_223/Y NAND2X1_269/B gnd NAND3X1_168/B vdd NAND2X1
XNAND2X1_247 NAND2X1_247/A NAND2X1_247/B gnd NAND2X1_247/Y vdd NAND2X1
XNAND2X1_258 XOR2X1_15/Y NAND2X1_258/B gnd NAND2X1_260/B vdd NAND2X1
XNAND2X1_236 AOI22X1_23/B AOI22X1_23/A gnd NAND2X1_236/Y vdd NAND2X1
XNAND2X1_214 INVX1_199/A OR2X2_18/A gnd AOI22X1_20/A vdd NAND2X1
XNAND2X1_203 NAND2X1_203/A INVX1_195/Y gnd INVX1_196/A vdd NAND2X1
XNAND2X1_225 NAND3X1_95/B NAND3X1_95/C gnd AOI22X1_26/B vdd NAND2X1
XFILL_0_2_0 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XOR2X2_30 OR2X2_30/A OR2X2_30/B gnd OR2X2_30/Y vdd OR2X2
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XXNOR2X1_3 XNOR2X1_3/A XOR2X1_2/B gnd OAI21X1_7/B vdd XNOR2X1
XINVX1_3 x1[0] gnd INVX1_3/Y vdd INVX1
XFILL_22_0_0 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XOAI21X1_391 AOI22X1_53/Y AOI22X1_54/Y OAI21X1_391/C gnd NAND3X1_366/A vdd OAI21X1
XOAI21X1_380 OAI21X1_362/C NOR2X1_224/A XOR2X1_25/B gnd OAI21X1_380/Y vdd OAI21X1
XAND2X2_3 AND2X2_3/A INVX1_45/Y gnd AND2X2_3/Y vdd AND2X2
XNAND3X1_19 INVX2_9/A INVX2_13/Y INVX1_146/Y gnd NOR3X1_2/A vdd NAND3X1
XNOR2X1_19 x0[1] INVX1_34/Y gnd NOR2X1_21/A vdd NOR2X1
XNOR2X1_109 OR2X2_9/B OR2X2_9/A gnd AOI22X1_6/C vdd NOR2X1
XINVX1_285 INVX1_285/A gnd OR2X2_31/B vdd INVX1
XINVX1_296 INVX1_296/A gnd INVX1_296/Y vdd INVX1
XINVX1_274 INVX1_274/A gnd INVX1_274/Y vdd INVX1
XINVX1_252 INVX1_252/A gnd INVX1_252/Y vdd INVX1
XINVX1_263 INVX1_263/A gnd INVX1_263/Y vdd INVX1
XINVX1_230 INVX1_230/A gnd INVX1_230/Y vdd INVX1
XINVX1_241 INVX1_241/A gnd INVX1_241/Y vdd INVX1
XNAND2X1_41 INVX1_90/Y NAND3X1_7/C gnd NOR2X1_58/B vdd NAND2X1
XNAND2X1_52 AND2X2_45/B OR2X2_4/B gnd OAI21X1_87/C vdd NAND2X1
XNAND2X1_30 INVX1_116/A BUFX4_12/Y gnd OAI21X1_40/C vdd NAND2X1
XNAND2X1_74 INVX1_47/A INVX1_78/A gnd NAND2X1_74/Y vdd NAND2X1
XNAND2X1_63 NOR2X1_65/B INVX1_110/Y gnd NAND2X1_65/B vdd NAND2X1
XNAND2X1_96 INVX1_187/A BUFX4_12/Y gnd NAND2X1_96/Y vdd NAND2X1
XNAND2X1_85 INVX1_52/A INVX1_82/Y gnd NAND2X1_85/Y vdd NAND2X1
XAOI22X1_50 INVX2_37/A INVX1_97/A INVX1_96/A INVX1_95/A gnd OAI22X1_21/D vdd AOI22X1
XNAND3X1_205 INVX1_257/Y NAND2X1_332/Y OAI21X1_307/Y gnd NAND3X1_205/Y vdd NAND3X1
XNAND3X1_216 XNOR2X1_40/Y NAND3X1_214/Y NAND3X1_215/Y gnd NAND3X1_216/Y vdd NAND3X1
XNAND3X1_249 NAND3X1_243/Y NAND2X1_352/Y AND2X2_41/Y gnd NAND3X1_249/Y vdd NAND3X1
XNAND3X1_238 INVX1_265/A NAND3X1_234/Y NAND3X1_238/C gnd NAND2X1_338/A vdd NAND3X1
XNAND3X1_227 NAND3X1_225/Y NAND3X1_231/C OR2X2_24/Y gnd NAND3X1_230/C vdd NAND3X1
XOAI22X1_1 BUFX4_2/Y INVX1_12/Y AND2X2_1/Y OAI22X1_1/D gnd OAI22X1_1/Y vdd OAI22X1
XNAND2X1_407 AOI22X1_48/B AOI22X1_48/A gnd NAND3X1_292/C vdd NAND2X1
XNAND2X1_418 INVX2_36/A INVX1_99/A gnd NOR2X1_224/A vdd NAND2X1
XNAND2X1_429 NAND2X1_429/A NAND2X1_427/Y gnd OR2X2_33/B vdd NAND2X1
XINVX2_21 INVX2_21/A gnd INVX2_21/Y vdd INVX2
XINVX2_10 INVX2_10/A gnd INVX2_10/Y vdd INVX2
XINVX2_43 INVX2_43/A gnd INVX2_43/Y vdd INVX2
XINVX2_32 gnd gnd INVX2_32/Y vdd INVX2
XOAI21X1_39 INVX1_48/Y INVX1_49/Y OR2X2_2/A gnd XNOR2X1_9/A vdd OAI21X1
XOAI21X1_17 BUFX4_8/Y INVX1_24/Y OAI21X1_21/C gnd OAI21X1_17/Y vdd OAI21X1
XOAI21X1_28 INVX1_32/Y INVX1_33/Y AOI21X1_6/A gnd NAND2X1_15/B vdd OAI21X1
XOAI21X1_209 INVX2_15/Y NOR3X1_3/C AOI21X1_56/A gnd NOR3X1_5/B vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XDFFPOSX1_134 BUFX2_30/A DFFSR_1/CLK XOR2X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_101 INVX1_28/A CLKBUF1_7/Y OAI21X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_112 BUFX2_8/A CLKBUF1_3/Y NAND2X1_360/Y gnd vdd DFFPOSX1
XDFFPOSX1_123 BUFX2_19/A CLKBUF1_6/Y XNOR2X1_18/Y gnd vdd DFFPOSX1
XNAND2X1_248 NAND2X1_248/A NAND2X1_248/B gnd NAND2X1_248/Y vdd NAND2X1
XNAND2X1_259 AOI21X1_89/Y XNOR2X1_36/Y gnd NAND2X1_259/Y vdd NAND2X1
XNAND2X1_237 OR2X2_19/A INVX1_210/A gnd AOI22X1_22/C vdd NAND2X1
XNAND2X1_215 NAND3X1_82/C NAND3X1_82/Y gnd INVX1_202/A vdd NAND2X1
XNAND2X1_204 XOR2X1_12/Y INVX1_196/Y gnd AOI21X1_72/A vdd NAND2X1
XNAND2X1_226 AOI22X1_26/B AND2X2_27/Y gnd NAND2X1_227/A vdd NAND2X1
XFILL_0_2_1 gnd vdd FILL
XFILL_16_2_1 gnd vdd FILL
XOR2X2_31 OR2X2_31/A OR2X2_31/B gnd OR2X2_31/Y vdd OR2X2
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XXNOR2X1_4 XNOR2X1_4/A NOR2X1_9/Y gnd XNOR2X1_4/Y vdd XNOR2X1
XOR2X2_20 OR2X2_20/A OR2X2_20/B gnd OR2X2_20/Y vdd OR2X2
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_22_0_1 gnd vdd FILL
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XOAI21X1_370 NOR3X1_12/Y AOI21X1_142/Y INVX1_297/Y gnd OAI21X1_370/Y vdd OAI21X1
XAND2X2_4 x0[5] x2[5] gnd AND2X2_4/Y vdd AND2X2
XOAI21X1_392 OAI22X1_22/C OAI22X1_22/D OAI21X1_392/C gnd OAI21X1_392/Y vdd OAI21X1
XOAI21X1_381 OAI21X1_383/A NOR2X1_225/Y INVX1_307/A gnd OAI21X1_381/Y vdd OAI21X1
XINVX1_297 INVX1_297/A gnd INVX1_297/Y vdd INVX1
XINVX1_286 INVX1_286/A gnd INVX1_286/Y vdd INVX1
XINVX1_275 INVX1_95/A gnd INVX1_275/Y vdd INVX1
XINVX1_264 INVX1_264/A gnd INVX1_264/Y vdd INVX1
XINVX1_253 NOR3X1_8/B gnd INVX1_253/Y vdd INVX1
XINVX1_231 INVX1_231/A gnd INVX1_231/Y vdd INVX1
XINVX1_242 INVX1_242/A gnd INVX1_242/Y vdd INVX1
XINVX1_220 INVX1_220/A gnd INVX1_220/Y vdd INVX1
XNAND2X1_31 x0[6] x2[6] gnd OAI21X1_41/A vdd NAND2X1
XNAND2X1_20 x0[3] x2[3] gnd OAI21X1_34/C vdd NAND2X1
XNAND2X1_42 INVX2_35/A OR2X2_4/B gnd OAI21X1_75/C vdd NAND2X1
XNAND2X1_53 BUFX4_6/Y INVX1_30/A gnd OAI21X1_88/C vdd NAND2X1
XNAND2X1_75 NAND2X1_74/Y NAND2X1_75/B gnd NAND2X1_75/Y vdd NAND2X1
XNAND2X1_64 INVX1_109/A INVX1_110/A gnd NAND2X1_65/A vdd NAND2X1
XNAND2X1_97 INVX2_21/A BUFX4_13/Y gnd NAND2X1_97/Y vdd NAND2X1
XNAND2X1_86 INVX1_139/A BUFX4_10/Y gnd NAND2X1_86/Y vdd NAND2X1
XAOI22X1_51 INVX1_290/Y INVX2_44/Y INVX1_298/Y AOI22X1_51/D gnd AOI22X1_51/Y vdd AOI22X1
XAOI22X1_40 AOI22X1_38/A AOI22X1_38/B AOI22X1_37/C AOI22X1_37/D gnd AOI22X1_40/Y vdd
+ AOI22X1
XNAND3X1_239 AOI21X1_114/Y NAND3X1_234/B NAND3X1_234/C gnd NAND3X1_239/Y vdd NAND3X1
XNAND3X1_217 INVX1_262/Y NAND3X1_213/Y NAND3X1_216/Y gnd NAND3X1_217/Y vdd NAND3X1
XNAND3X1_228 NAND3X1_228/A NAND3X1_228/B NAND2X1_337/Y gnd NAND3X1_232/A vdd NAND3X1
XNAND3X1_206 NAND3X1_204/Y NAND3X1_205/Y INVX1_259/Y gnd NAND3X1_206/Y vdd NAND3X1
XOAI22X1_2 BUFX4_8/Y INVX1_20/Y NOR2X1_13/Y OAI22X1_2/D gnd OAI22X1_2/Y vdd OAI22X1
XNAND2X1_408 AOI22X1_49/B AOI22X1_49/A gnd NAND3X1_295/C vdd NAND2X1
XNAND2X1_419 NAND2X1_419/A NAND2X1_419/B gnd NAND3X1_308/A vdd NAND2X1
XINVX2_44 INVX2_44/A gnd INVX2_44/Y vdd INVX2
XINVX2_11 INVX2_11/A gnd INVX2_11/Y vdd INVX2
XINVX2_33 INVX2_33/A gnd INVX2_33/Y vdd INVX2
XINVX2_22 INVX2_22/A gnd INVX2_22/Y vdd INVX2
XOAI21X1_29 BUFX4_16/Y OAI21X1_29/B OAI21X1_29/C gnd OAI21X1_29/Y vdd OAI21X1
XOAI21X1_18 BUFX4_6/Y INVX2_2/Y OAI21X1_21/C gnd OAI21X1_18/Y vdd OAI21X1
XFILL_12_2 gnd vdd FILL
XDFFPOSX1_102 INVX2_4/A CLKBUF1_7/Y OAI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_135 BUFX2_31/A DFFSR_1/CLK XNOR2X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_113 BUFX2_9/A CLKBUF1_3/Y NOR2X1_134/Y gnd vdd DFFPOSX1
XDFFPOSX1_124 BUFX2_20/A CLKBUF1_6/Y NOR2X1_108/Y gnd vdd DFFPOSX1
XNAND2X1_216 INVX2_19/A INVX1_105/A gnd NOR2X1_148/B vdd NAND2X1
XNAND2X1_205 OR2X2_16/B OR2X2_16/A gnd AOI21X1_75/B vdd NAND2X1
XNAND2X1_238 NAND2X1_238/A NAND2X1_238/B gnd AOI21X1_94/B vdd NAND2X1
XNAND2X1_249 AND2X2_28/Y AND2X2_29/Y gnd AND2X2_31/A vdd NAND2X1
XNAND2X1_227 NAND2X1_227/A NAND3X1_98/Y gnd AOI21X1_84/B vdd NAND2X1
XFILL_0_2_2 gnd vdd FILL
XFILL_16_2_2 gnd vdd FILL
XOR2X2_32 OR2X2_32/A OR2X2_32/B gnd OR2X2_32/Y vdd OR2X2
XOR2X2_10 OR2X2_10/A OR2X2_10/B gnd OR2X2_10/Y vdd OR2X2
XOR2X2_21 OR2X2_21/A OR2X2_21/B gnd OR2X2_21/Y vdd OR2X2
XXNOR2X1_5 XNOR2X1_5/A INVX1_25/A gnd XNOR2X1_5/Y vdd XNOR2X1
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XINVX1_5 x1[1] gnd INVX1_5/Y vdd INVX1
.ends


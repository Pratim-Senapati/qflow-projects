VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter
  CLASS BLOCK ;
  FOREIGN counter ;
  ORIGIN 1.900 0.000 ;
  SIZE 88.600 BY 62.000 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 38.600 50.800 39.400 51.000 ;
        RECT 12.400 50.200 39.400 50.800 ;
        RECT 1.200 41.600 2.000 50.200 ;
        RECT 12.400 49.600 13.200 50.200 ;
        RECT 15.800 50.000 16.600 50.200 ;
        RECT 9.200 41.600 10.000 46.200 ;
        RECT 12.400 41.600 13.200 46.200 ;
        RECT 15.600 41.600 16.400 46.200 ;
        RECT 22.000 41.600 22.800 46.200 ;
        RECT 25.200 41.600 26.000 46.200 ;
        RECT 33.200 41.600 34.000 46.200 ;
        RECT 36.400 41.600 37.200 46.200 ;
        RECT 39.600 41.600 40.400 46.200 ;
        RECT 42.800 41.600 43.600 46.200 ;
        RECT 46.000 41.600 46.800 49.000 ;
        RECT 50.800 41.600 51.600 50.200 ;
        RECT 57.200 41.600 58.000 46.200 ;
        RECT 65.200 41.600 66.000 45.800 ;
        RECT 68.400 41.600 69.200 46.200 ;
        RECT 71.600 41.600 72.400 49.000 ;
        RECT 76.400 41.600 77.200 49.000 ;
        RECT 81.200 41.600 82.000 49.000 ;
        RECT 0.400 40.400 84.400 41.600 ;
        RECT 1.200 34.300 2.000 39.800 ;
        RECT 2.800 34.300 3.600 40.400 ;
        RECT 9.200 36.300 10.000 36.400 ;
        RECT 10.800 36.300 11.600 40.400 ;
        RECT 9.200 35.800 11.600 36.300 ;
        RECT 14.000 35.800 14.800 40.400 ;
        RECT 17.200 35.800 18.000 40.400 ;
        RECT 23.600 35.800 24.400 40.400 ;
        RECT 26.800 35.800 27.600 40.400 ;
        RECT 34.800 35.800 35.600 40.400 ;
        RECT 38.000 35.800 38.800 40.400 ;
        RECT 41.200 35.800 42.000 40.400 ;
        RECT 44.400 35.800 45.200 40.400 ;
        RECT 47.800 39.800 48.600 40.400 ;
        RECT 9.200 35.700 11.500 35.800 ;
        RECT 9.200 35.600 10.000 35.700 ;
        RECT 1.200 33.700 3.600 34.300 ;
        RECT 1.200 31.800 2.000 33.700 ;
        RECT 2.800 33.000 3.600 33.700 ;
        RECT 47.600 33.200 48.600 39.800 ;
        RECT 53.800 33.200 54.800 40.400 ;
        RECT 63.800 39.800 64.600 40.400 ;
        RECT 63.600 33.200 64.600 39.800 ;
        RECT 69.800 33.200 70.800 40.400 ;
        RECT 74.800 33.000 75.600 40.400 ;
        RECT 79.600 33.000 80.400 40.400 ;
        RECT 14.000 31.800 14.800 32.400 ;
        RECT 17.400 31.800 18.200 32.000 ;
        RECT 1.200 29.600 1.800 31.800 ;
        RECT 14.000 31.200 41.000 31.800 ;
        RECT 40.200 31.000 41.000 31.200 ;
        RECT 4.400 30.300 5.200 30.400 ;
        RECT 9.200 30.300 10.000 30.400 ;
        RECT 4.400 29.700 10.000 30.300 ;
        RECT 1.200 22.200 2.000 29.600 ;
        RECT 4.400 28.800 5.200 29.700 ;
        RECT 9.200 29.600 10.000 29.700 ;
        RECT 30.600 10.800 31.400 11.000 ;
        RECT 78.600 10.800 79.400 11.000 ;
        RECT 4.400 10.200 31.400 10.800 ;
        RECT 52.400 10.200 79.400 10.800 ;
        RECT 4.400 9.600 5.200 10.200 ;
        RECT 7.800 10.000 8.600 10.200 ;
        RECT 52.400 9.600 53.200 10.200 ;
        RECT 55.800 10.000 56.600 10.200 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 4.400 1.600 5.200 6.200 ;
        RECT 7.600 1.600 8.400 6.200 ;
        RECT 14.000 1.600 14.800 6.200 ;
        RECT 17.200 1.600 18.000 6.200 ;
        RECT 25.200 1.600 26.000 6.200 ;
        RECT 28.400 1.600 29.200 6.200 ;
        RECT 31.600 1.600 32.400 6.200 ;
        RECT 34.800 1.600 35.600 6.200 ;
        RECT 42.800 1.600 43.600 6.200 ;
        RECT 49.200 1.600 50.000 6.200 ;
        RECT 52.400 1.600 53.200 6.200 ;
        RECT 55.600 1.600 56.400 6.200 ;
        RECT 62.000 1.600 62.800 6.200 ;
        RECT 65.200 1.600 66.000 6.200 ;
        RECT 73.200 1.600 74.000 6.200 ;
        RECT 76.400 1.600 77.200 6.200 ;
        RECT 79.600 1.600 80.400 6.200 ;
        RECT 82.800 1.600 83.600 6.200 ;
        RECT 0.400 0.400 84.400 1.600 ;
      LAYER via1 ;
        RECT 12.400 43.600 13.200 44.400 ;
        RECT 15.800 40.600 16.600 41.400 ;
        RECT 17.200 40.600 18.000 41.400 ;
        RECT 18.600 40.600 19.400 41.400 ;
        RECT 14.000 37.600 14.800 38.400 ;
        RECT 14.000 31.600 14.800 32.400 ;
        RECT 4.400 3.600 5.200 4.400 ;
        RECT 52.400 3.600 53.200 4.400 ;
        RECT 15.800 0.600 16.600 1.400 ;
        RECT 17.200 0.600 18.000 1.400 ;
        RECT 18.600 0.600 19.400 1.400 ;
      LAYER metal2 ;
        RECT 12.400 49.600 13.200 50.400 ;
        RECT 12.500 44.400 13.100 49.600 ;
        RECT 12.400 43.600 13.200 44.400 ;
        RECT 15.200 40.600 20.000 41.400 ;
        RECT 14.000 37.600 14.800 38.400 ;
        RECT 9.200 35.600 10.000 36.400 ;
        RECT 9.300 32.400 9.900 35.600 ;
        RECT 14.100 32.400 14.700 37.600 ;
        RECT 9.200 31.600 10.000 32.400 ;
        RECT 14.000 31.600 14.800 32.400 ;
        RECT 9.300 30.400 9.900 31.600 ;
        RECT 9.200 29.600 10.000 30.400 ;
        RECT 4.400 9.600 5.200 10.400 ;
        RECT 52.400 9.600 53.200 10.400 ;
        RECT 4.500 4.400 5.100 9.600 ;
        RECT 52.500 4.400 53.100 9.600 ;
        RECT 4.400 3.600 5.200 4.400 ;
        RECT 52.400 3.600 53.200 4.400 ;
        RECT 15.200 0.600 20.000 1.400 ;
      LAYER via2 ;
        RECT 15.800 40.600 16.600 41.400 ;
        RECT 17.200 40.600 18.000 41.400 ;
        RECT 18.600 40.600 19.400 41.400 ;
        RECT 15.800 0.600 16.600 1.400 ;
        RECT 17.200 0.600 18.000 1.400 ;
        RECT 18.600 0.600 19.400 1.400 ;
      LAYER metal3 ;
        RECT 15.200 40.400 20.000 41.600 ;
        RECT 9.200 32.300 10.000 32.400 ;
        RECT -1.900 31.700 10.000 32.300 ;
        RECT 9.200 31.600 10.000 31.700 ;
        RECT 15.200 0.400 20.000 1.600 ;
      LAYER via3 ;
        RECT 15.600 40.600 16.400 41.400 ;
        RECT 17.200 40.600 18.000 41.400 ;
        RECT 18.800 40.600 19.600 41.400 ;
        RECT 15.600 0.600 16.400 1.400 ;
        RECT 17.200 0.600 18.000 1.400 ;
        RECT 18.800 0.600 19.600 1.400 ;
      LAYER metal4 ;
        RECT 15.200 0.000 20.000 62.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.400 60.400 84.400 61.600 ;
        RECT 1.200 55.800 2.000 60.400 ;
        RECT 12.400 55.800 13.200 60.400 ;
        RECT 22.000 57.800 22.800 60.400 ;
        RECT 25.200 57.800 26.000 60.400 ;
        RECT 36.400 55.800 37.200 60.400 ;
        RECT 42.800 57.800 43.600 60.400 ;
        RECT 45.000 55.800 45.800 60.400 ;
        RECT 49.200 57.800 50.000 60.400 ;
        RECT 50.800 57.800 51.600 60.400 ;
        RECT 54.000 57.800 54.800 60.400 ;
        RECT 57.200 57.800 58.000 60.400 ;
        RECT 68.400 53.800 69.200 60.400 ;
        RECT 71.600 55.800 72.400 60.400 ;
        RECT 76.400 55.800 77.200 60.400 ;
        RECT 81.200 55.800 82.000 60.400 ;
        RECT 81.200 31.800 82.000 39.800 ;
        RECT 78.000 28.800 78.800 30.400 ;
        RECT 81.400 29.600 82.000 31.800 ;
        RECT 81.200 26.300 82.000 29.600 ;
        RECT 79.700 26.200 82.000 26.300 ;
        RECT 2.800 21.600 3.600 26.200 ;
        RECT 14.000 21.600 14.800 26.200 ;
        RECT 23.600 21.600 24.400 24.200 ;
        RECT 26.800 21.600 27.600 24.200 ;
        RECT 38.000 21.600 38.800 26.200 ;
        RECT 44.400 21.600 45.200 24.200 ;
        RECT 47.600 22.200 48.600 25.600 ;
        RECT 47.800 21.600 48.600 22.200 ;
        RECT 53.800 21.600 54.800 25.600 ;
        RECT 63.600 22.200 64.600 25.600 ;
        RECT 63.800 21.600 64.600 22.200 ;
        RECT 69.800 21.600 70.800 25.600 ;
        RECT 74.800 21.600 75.600 26.200 ;
        RECT 79.600 25.700 82.000 26.200 ;
        RECT 79.600 21.600 80.400 25.700 ;
        RECT 81.200 22.200 82.000 25.700 ;
        RECT 0.400 20.400 84.400 21.600 ;
        RECT 4.400 15.800 5.200 20.400 ;
        RECT 14.000 17.800 14.800 20.400 ;
        RECT 17.200 17.800 18.000 20.400 ;
        RECT 28.400 15.800 29.200 20.400 ;
        RECT 34.800 17.800 35.600 20.400 ;
        RECT 42.800 17.800 43.600 20.400 ;
        RECT 52.400 15.800 53.200 20.400 ;
        RECT 62.000 17.800 62.800 20.400 ;
        RECT 65.200 17.800 66.000 20.400 ;
        RECT 76.400 18.300 77.200 20.400 ;
        RECT 78.000 18.300 78.800 18.400 ;
        RECT 76.400 17.700 78.800 18.300 ;
        RECT 82.800 17.800 83.600 20.400 ;
        RECT 76.400 15.800 77.200 17.700 ;
        RECT 78.000 17.600 78.800 17.700 ;
      LAYER via1 ;
        RECT 52.600 60.600 53.400 61.400 ;
        RECT 54.000 60.600 54.800 61.400 ;
        RECT 55.400 60.600 56.200 61.400 ;
        RECT 78.000 29.600 78.800 30.400 ;
        RECT 79.600 25.400 80.400 26.200 ;
        RECT 52.600 20.600 53.400 21.400 ;
        RECT 54.000 20.600 54.800 21.400 ;
        RECT 55.400 20.600 56.200 21.400 ;
      LAYER metal2 ;
        RECT 52.000 60.600 56.800 61.400 ;
        RECT 79.600 31.600 80.400 32.400 ;
        RECT 78.000 29.600 78.800 30.400 ;
        RECT 52.000 20.600 56.800 21.400 ;
        RECT 78.100 18.400 78.700 29.600 ;
        RECT 79.700 26.200 80.300 31.600 ;
        RECT 79.600 25.400 80.400 26.200 ;
        RECT 78.000 17.600 78.800 18.400 ;
      LAYER via2 ;
        RECT 52.600 60.600 53.400 61.400 ;
        RECT 54.000 60.600 54.800 61.400 ;
        RECT 55.400 60.600 56.200 61.400 ;
        RECT 52.600 20.600 53.400 21.400 ;
        RECT 54.000 20.600 54.800 21.400 ;
        RECT 55.400 20.600 56.200 21.400 ;
      LAYER metal3 ;
        RECT 52.000 60.400 56.800 61.600 ;
        RECT 79.600 32.300 80.400 32.400 ;
        RECT 79.600 31.700 86.700 32.300 ;
        RECT 79.600 31.600 80.400 31.700 ;
        RECT 52.000 20.400 56.800 21.600 ;
      LAYER via3 ;
        RECT 52.400 60.600 53.200 61.400 ;
        RECT 54.000 60.600 54.800 61.400 ;
        RECT 55.600 60.600 56.400 61.400 ;
        RECT 52.400 20.600 53.200 21.400 ;
        RECT 54.000 20.600 54.800 21.400 ;
        RECT 55.600 20.600 56.400 21.400 ;
      LAYER metal4 ;
        RECT 52.000 0.000 56.800 62.000 ;
    END
  END gnd
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 25.200 55.600 26.800 56.400 ;
        RECT 26.800 25.600 28.400 26.400 ;
        RECT 17.200 15.600 18.800 16.400 ;
        RECT 65.200 15.600 66.800 16.400 ;
      LAYER metal2 ;
        RECT 25.200 55.600 26.000 56.400 ;
        RECT 25.300 44.300 25.900 55.600 ;
        RECT 25.300 43.700 27.500 44.300 ;
        RECT 17.200 35.600 18.000 36.400 ;
        RECT 17.300 26.400 17.900 35.600 ;
        RECT 26.900 26.400 27.500 43.700 ;
        RECT 17.200 25.600 18.000 26.400 ;
        RECT 26.800 25.600 27.600 26.400 ;
        RECT 17.300 16.400 17.900 25.600 ;
        RECT 26.900 16.400 27.500 25.600 ;
        RECT 17.200 15.600 18.000 16.400 ;
        RECT 26.800 15.600 27.600 16.400 ;
        RECT 65.200 15.600 66.000 16.400 ;
      LAYER metal3 ;
        RECT 17.200 36.300 18.000 36.400 ;
        RECT -1.900 35.700 18.000 36.300 ;
        RECT 17.200 35.600 18.000 35.700 ;
        RECT 17.200 26.300 18.000 26.400 ;
        RECT 26.800 26.300 27.600 26.400 ;
        RECT 17.200 25.700 27.600 26.300 ;
        RECT 17.200 25.600 18.000 25.700 ;
        RECT 26.800 25.600 27.600 25.700 ;
        RECT 26.800 16.300 27.600 16.400 ;
        RECT 65.200 16.300 66.000 16.400 ;
        RECT 26.800 15.700 66.000 16.300 ;
        RECT 26.800 15.600 27.600 15.700 ;
        RECT 65.200 15.600 66.000 15.700 ;
    END
  END clk
  PIN rst
    PORT
      LAYER metal1 ;
        RECT 1.200 53.600 2.000 55.200 ;
      LAYER metal2 ;
        RECT 1.200 53.600 2.000 54.400 ;
        RECT 1.300 50.400 1.900 53.600 ;
        RECT 1.200 49.600 2.000 50.400 ;
      LAYER metal3 ;
        RECT 1.200 50.300 2.000 50.400 ;
        RECT -1.900 49.700 2.000 50.300 ;
        RECT 1.200 49.600 2.000 49.700 ;
    END
  END rst
  PIN count[0]
    PORT
      LAYER metal1 ;
        RECT 73.200 52.400 74.000 59.800 ;
        RECT 73.400 50.200 74.000 52.400 ;
        RECT 73.200 42.200 74.000 50.200 ;
      LAYER via1 ;
        RECT 73.200 57.600 74.000 58.400 ;
      LAYER metal2 ;
        RECT 73.200 57.600 74.000 58.400 ;
      LAYER metal3 ;
        RECT 73.200 58.300 74.000 58.400 ;
        RECT 73.200 57.700 86.700 58.300 ;
        RECT 73.200 57.600 74.000 57.700 ;
    END
  END count[0]
  PIN count[1]
    PORT
      LAYER metal1 ;
        RECT 78.000 52.400 78.800 59.800 ;
        RECT 78.200 50.200 78.800 52.400 ;
        RECT 78.000 42.200 78.800 50.200 ;
      LAYER via1 ;
        RECT 78.000 53.600 78.800 54.400 ;
      LAYER metal2 ;
        RECT 78.000 53.600 78.800 54.400 ;
      LAYER metal3 ;
        RECT 78.000 54.300 78.800 54.400 ;
        RECT 78.000 53.700 86.700 54.300 ;
        RECT 78.000 53.600 78.800 53.700 ;
    END
  END count[1]
  PIN count[2]
    PORT
      LAYER metal1 ;
        RECT 82.800 52.400 83.600 59.800 ;
        RECT 83.000 50.200 83.600 52.400 ;
        RECT 82.800 42.200 83.600 50.200 ;
      LAYER via1 ;
        RECT 82.800 47.600 83.600 48.400 ;
      LAYER metal2 ;
        RECT 82.800 49.600 83.600 50.400 ;
        RECT 82.900 48.400 83.500 49.600 ;
        RECT 82.800 47.600 83.600 48.400 ;
      LAYER metal3 ;
        RECT 82.800 50.300 83.600 50.400 ;
        RECT 82.800 49.700 86.700 50.300 ;
        RECT 82.800 49.600 83.600 49.700 ;
    END
  END count[2]
  PIN count[3]
    PORT
      LAYER metal1 ;
        RECT 76.400 31.800 77.200 39.800 ;
        RECT 76.600 29.600 77.200 31.800 ;
        RECT 76.400 22.200 77.200 29.600 ;
      LAYER via1 ;
        RECT 76.400 27.600 77.200 28.400 ;
      LAYER metal2 ;
        RECT 76.400 29.600 77.200 30.400 ;
        RECT 76.500 28.400 77.100 29.600 ;
        RECT 76.400 27.600 77.200 28.400 ;
      LAYER metal3 ;
        RECT 76.400 30.300 77.200 30.400 ;
        RECT 76.400 29.700 86.700 30.300 ;
        RECT 76.400 29.600 77.200 29.700 ;
    END
  END count[3]
  OBS
      LAYER metal1 ;
        RECT 2.800 52.300 3.600 59.800 ;
        RECT 9.200 53.800 10.000 59.800 ;
        RECT 15.600 56.600 16.400 59.800 ;
        RECT 17.200 57.000 18.000 59.800 ;
        RECT 18.800 57.000 19.600 59.800 ;
        RECT 20.400 57.000 21.200 59.800 ;
        RECT 23.600 57.000 24.400 59.800 ;
        RECT 26.800 57.000 27.600 59.800 ;
        RECT 28.400 57.000 29.200 59.800 ;
        RECT 30.000 57.000 30.800 59.800 ;
        RECT 31.600 57.000 32.400 59.800 ;
        RECT 13.800 55.800 16.400 56.600 ;
        RECT 33.200 56.600 34.000 59.800 ;
        RECT 19.800 55.800 24.400 56.400 ;
        RECT 13.800 55.200 14.600 55.800 ;
        RECT 11.600 54.400 14.600 55.200 ;
        RECT 9.200 53.000 18.000 53.800 ;
        RECT 19.800 53.400 20.600 55.800 ;
        RECT 23.600 55.600 24.400 55.800 ;
        RECT 29.800 55.600 30.800 56.400 ;
        RECT 33.200 55.800 35.600 56.600 ;
        RECT 22.000 53.600 22.800 55.200 ;
        RECT 23.600 54.800 24.400 55.000 ;
        RECT 23.600 54.200 28.000 54.800 ;
        RECT 27.200 54.000 28.000 54.200 ;
        RECT 7.600 52.300 8.400 52.400 ;
        RECT 2.800 51.700 8.400 52.300 ;
        RECT 2.800 42.200 3.600 51.700 ;
        RECT 7.600 51.600 8.400 51.700 ;
        RECT 9.200 47.400 10.000 53.000 ;
        RECT 18.600 52.600 20.600 53.400 ;
        RECT 24.400 52.600 27.600 53.400 ;
        RECT 30.000 52.800 30.800 55.600 ;
        RECT 34.800 55.200 35.600 55.800 ;
        RECT 34.800 54.600 36.600 55.200 ;
        RECT 35.800 53.400 36.600 54.600 ;
        RECT 39.600 54.600 40.400 59.800 ;
        RECT 41.200 56.000 42.000 59.800 ;
        RECT 41.200 55.200 42.200 56.000 ;
        RECT 39.600 54.000 40.800 54.600 ;
        RECT 35.800 52.600 39.600 53.400 ;
        RECT 10.600 52.000 11.400 52.200 ;
        RECT 12.400 52.000 13.200 52.400 ;
        RECT 15.600 52.000 16.400 52.400 ;
        RECT 33.200 52.000 34.000 52.600 ;
        RECT 40.200 52.000 40.800 54.000 ;
        RECT 10.600 51.400 34.000 52.000 ;
        RECT 40.000 51.400 40.800 52.000 ;
        RECT 40.000 49.600 40.600 51.400 ;
        RECT 41.400 50.800 42.200 55.200 ;
        RECT 47.600 55.800 48.400 59.800 ;
        RECT 52.400 57.800 53.200 59.800 ;
        RECT 49.000 56.400 49.800 57.200 ;
        RECT 46.000 52.800 46.800 54.400 ;
        RECT 47.600 54.300 48.200 55.800 ;
        RECT 49.200 55.600 50.000 56.400 ;
        RECT 50.800 55.600 51.600 57.200 ;
        RECT 50.900 54.300 51.500 55.600 ;
        RECT 52.600 54.400 53.200 57.800 ;
        RECT 47.600 53.700 51.500 54.300 ;
        RECT 44.400 52.200 45.200 52.400 ;
        RECT 47.600 52.200 48.200 53.700 ;
        RECT 52.400 53.600 53.200 54.400 ;
        RECT 49.200 52.200 50.000 52.400 ;
        RECT 44.400 51.600 46.000 52.200 ;
        RECT 47.600 51.600 50.000 52.200 ;
        RECT 45.200 51.200 46.000 51.600 ;
        RECT 18.800 49.400 19.600 49.600 ;
        RECT 14.200 49.000 19.600 49.400 ;
        RECT 13.400 48.800 19.600 49.000 ;
        RECT 20.600 49.000 29.200 49.600 ;
        RECT 10.800 48.000 12.400 48.800 ;
        RECT 13.400 48.200 14.800 48.800 ;
        RECT 20.600 48.200 21.200 49.000 ;
        RECT 28.400 48.800 29.200 49.000 ;
        RECT 31.600 49.000 40.600 49.600 ;
        RECT 31.600 48.800 32.400 49.000 ;
        RECT 11.800 47.600 12.400 48.000 ;
        RECT 15.400 47.600 21.200 48.200 ;
        RECT 21.800 47.600 24.400 48.400 ;
        RECT 9.200 46.800 11.200 47.400 ;
        RECT 11.800 46.800 16.000 47.600 ;
        RECT 10.600 46.200 11.200 46.800 ;
        RECT 10.600 45.600 11.600 46.200 ;
        RECT 10.800 42.200 11.600 45.600 ;
        RECT 14.000 42.200 14.800 46.800 ;
        RECT 17.200 42.200 18.000 45.000 ;
        RECT 18.800 42.200 19.600 45.000 ;
        RECT 20.400 42.200 21.200 47.000 ;
        RECT 23.600 42.200 24.400 47.000 ;
        RECT 26.800 42.200 27.600 48.400 ;
        RECT 34.800 47.600 37.400 48.400 ;
        RECT 30.000 46.800 34.200 47.600 ;
        RECT 28.400 42.200 29.200 45.000 ;
        RECT 30.000 42.200 30.800 45.000 ;
        RECT 31.600 42.200 32.400 45.000 ;
        RECT 34.800 42.200 35.600 47.600 ;
        RECT 40.000 47.400 40.600 49.000 ;
        RECT 38.000 46.800 40.600 47.400 ;
        RECT 41.200 50.000 42.200 50.800 ;
        RECT 49.200 50.200 49.800 51.600 ;
        RECT 52.600 50.200 53.200 53.600 ;
        RECT 54.000 52.300 54.800 52.400 ;
        RECT 55.600 52.300 56.400 59.800 ;
        RECT 57.200 56.300 58.000 57.200 ;
        RECT 64.800 56.300 65.600 59.800 ;
        RECT 57.200 55.700 65.600 56.300 ;
        RECT 57.200 55.600 58.000 55.700 ;
        RECT 64.800 54.200 65.600 55.700 ;
        RECT 70.000 55.200 70.800 59.800 ;
        RECT 74.800 55.200 75.600 59.800 ;
        RECT 79.600 55.200 80.400 59.800 ;
        RECT 70.000 54.600 72.200 55.200 ;
        RECT 74.800 54.600 77.000 55.200 ;
        RECT 79.600 54.600 81.800 55.200 ;
        RECT 54.000 51.700 56.400 52.300 ;
        RECT 54.000 50.800 54.800 51.700 ;
        RECT 38.000 42.200 38.800 46.800 ;
        RECT 41.200 42.200 42.000 50.000 ;
        RECT 44.400 49.600 48.400 50.200 ;
        RECT 44.400 42.200 45.200 49.600 ;
        RECT 47.600 42.200 48.400 49.600 ;
        RECT 49.200 42.200 50.000 50.200 ;
        RECT 52.400 49.400 54.200 50.200 ;
        RECT 53.400 42.200 54.200 49.400 ;
        RECT 55.600 42.200 56.400 51.700 ;
        RECT 63.800 53.800 65.600 54.200 ;
        RECT 63.800 53.600 65.400 53.800 ;
        RECT 63.800 50.400 64.400 53.600 ;
        RECT 66.000 51.600 67.600 52.400 ;
        RECT 70.000 52.300 70.800 53.200 ;
        RECT 68.400 51.700 70.800 52.300 ;
        RECT 63.600 49.600 64.400 50.400 ;
        RECT 66.800 50.300 67.600 50.400 ;
        RECT 68.400 50.300 69.200 51.700 ;
        RECT 70.000 51.600 70.800 51.700 ;
        RECT 71.600 51.600 72.200 54.600 ;
        RECT 74.800 51.600 75.600 53.200 ;
        RECT 76.400 51.600 77.000 54.600 ;
        RECT 79.600 51.600 80.400 53.200 ;
        RECT 81.200 51.600 81.800 54.600 ;
        RECT 66.800 49.700 69.200 50.300 ;
        RECT 71.600 50.800 72.800 51.600 ;
        RECT 76.400 50.800 77.600 51.600 ;
        RECT 81.200 50.800 82.400 51.600 ;
        RECT 71.600 50.200 72.200 50.800 ;
        RECT 76.400 50.200 77.000 50.800 ;
        RECT 81.200 50.200 81.800 50.800 ;
        RECT 66.800 49.600 67.600 49.700 ;
        RECT 68.400 49.600 69.200 49.700 ;
        RECT 70.000 49.600 72.200 50.200 ;
        RECT 74.800 49.600 77.000 50.200 ;
        RECT 79.600 49.600 81.800 50.200 ;
        RECT 63.800 47.000 64.400 49.600 ;
        RECT 65.200 47.600 66.000 49.200 ;
        RECT 63.800 46.400 67.400 47.000 ;
        RECT 63.800 46.200 64.400 46.400 ;
        RECT 62.000 44.300 62.800 44.400 ;
        RECT 63.600 44.300 64.400 46.200 ;
        RECT 62.000 43.700 64.400 44.300 ;
        RECT 62.000 43.600 62.800 43.700 ;
        RECT 63.600 42.200 64.400 43.700 ;
        RECT 66.800 46.200 67.400 46.400 ;
        RECT 66.800 42.200 67.600 46.200 ;
        RECT 70.000 42.200 70.800 49.600 ;
        RECT 74.800 42.200 75.600 49.600 ;
        RECT 79.600 42.200 80.400 49.600 ;
        RECT 4.400 32.400 5.200 39.800 ;
        RECT 12.400 36.400 13.200 39.800 ;
        RECT 12.200 35.800 13.200 36.400 ;
        RECT 12.200 35.200 12.800 35.800 ;
        RECT 15.600 35.200 16.400 39.800 ;
        RECT 18.800 37.000 19.600 39.800 ;
        RECT 20.400 37.000 21.200 39.800 ;
        RECT 3.000 31.800 5.200 32.400 ;
        RECT 10.800 34.600 12.800 35.200 ;
        RECT 3.000 31.200 3.600 31.800 ;
        RECT 2.400 30.400 3.600 31.200 ;
        RECT 3.000 27.400 3.600 30.400 ;
        RECT 10.800 29.000 11.600 34.600 ;
        RECT 13.400 34.400 17.600 35.200 ;
        RECT 22.000 35.000 22.800 39.800 ;
        RECT 25.200 35.000 26.000 39.800 ;
        RECT 13.400 34.000 14.000 34.400 ;
        RECT 12.400 33.200 14.000 34.000 ;
        RECT 17.000 33.800 22.800 34.400 ;
        RECT 15.000 33.200 16.400 33.800 ;
        RECT 15.000 33.000 21.200 33.200 ;
        RECT 15.800 32.600 21.200 33.000 ;
        RECT 20.400 32.400 21.200 32.600 ;
        RECT 22.200 33.000 22.800 33.800 ;
        RECT 23.400 33.600 26.000 34.400 ;
        RECT 28.400 33.600 29.200 39.800 ;
        RECT 30.000 37.000 30.800 39.800 ;
        RECT 31.600 37.000 32.400 39.800 ;
        RECT 33.200 37.000 34.000 39.800 ;
        RECT 31.600 34.400 35.800 35.200 ;
        RECT 36.400 34.400 37.200 39.800 ;
        RECT 39.600 35.200 40.400 39.800 ;
        RECT 39.600 34.600 42.200 35.200 ;
        RECT 36.400 33.600 39.000 34.400 ;
        RECT 30.000 33.000 30.800 33.200 ;
        RECT 22.200 32.400 30.800 33.000 ;
        RECT 33.200 33.000 34.000 33.200 ;
        RECT 41.600 33.000 42.200 34.600 ;
        RECT 33.200 32.400 42.200 33.000 ;
        RECT 41.600 30.600 42.200 32.400 ;
        RECT 42.800 32.000 43.600 39.800 ;
        RECT 46.000 32.400 46.800 39.800 ;
        RECT 47.800 32.400 48.600 32.600 ;
        RECT 42.800 31.200 43.800 32.000 ;
        RECT 46.000 31.800 48.600 32.400 ;
        RECT 50.400 31.800 52.000 39.800 ;
        RECT 54.000 32.400 54.800 32.600 ;
        RECT 55.600 32.400 56.400 39.800 ;
        RECT 54.000 31.800 56.400 32.400 ;
        RECT 62.000 32.400 62.800 39.800 ;
        RECT 63.400 32.400 64.200 32.600 ;
        RECT 62.000 31.800 64.200 32.400 ;
        RECT 66.400 32.400 68.000 39.800 ;
        RECT 70.000 32.400 70.800 32.600 ;
        RECT 71.600 32.400 72.400 39.800 ;
        RECT 66.400 31.800 68.400 32.400 ;
        RECT 70.000 31.800 72.400 32.400 ;
        RECT 73.200 32.400 74.000 39.800 ;
        RECT 78.000 32.400 78.800 39.800 ;
        RECT 73.200 31.800 75.400 32.400 ;
        RECT 78.000 31.800 80.200 32.400 ;
        RECT 12.200 30.000 35.600 30.600 ;
        RECT 41.600 30.000 42.400 30.600 ;
        RECT 12.200 29.800 13.000 30.000 ;
        RECT 14.000 29.600 14.800 30.000 ;
        RECT 17.200 29.600 18.000 30.000 ;
        RECT 34.800 29.400 35.600 30.000 ;
        RECT 10.800 28.200 19.600 29.000 ;
        RECT 20.200 28.600 22.200 29.400 ;
        RECT 26.000 28.600 29.200 29.400 ;
        RECT 3.000 26.800 5.200 27.400 ;
        RECT 4.400 22.200 5.200 26.800 ;
        RECT 10.800 22.200 11.600 28.200 ;
        RECT 13.200 26.800 16.200 27.600 ;
        RECT 15.400 26.200 16.200 26.800 ;
        RECT 21.400 26.200 22.200 28.600 ;
        RECT 23.600 26.800 24.400 28.400 ;
        RECT 28.800 27.800 29.600 28.000 ;
        RECT 25.200 27.200 29.600 27.800 ;
        RECT 25.200 27.000 26.000 27.200 ;
        RECT 31.600 26.400 32.400 29.200 ;
        RECT 37.400 28.600 41.200 29.400 ;
        RECT 37.400 27.400 38.200 28.600 ;
        RECT 41.800 28.000 42.400 30.000 ;
        RECT 25.200 26.200 26.000 26.400 ;
        RECT 15.400 25.400 18.000 26.200 ;
        RECT 21.400 25.600 26.000 26.200 ;
        RECT 31.400 25.600 32.400 26.400 ;
        RECT 36.400 26.800 38.200 27.400 ;
        RECT 41.200 27.400 42.400 28.000 ;
        RECT 43.000 30.300 43.800 31.200 ;
        RECT 49.000 30.400 49.800 30.600 ;
        RECT 51.000 30.400 51.600 31.800 ;
        RECT 63.600 31.200 64.200 31.800 ;
        RECT 63.600 30.600 67.000 31.200 ;
        RECT 66.200 30.400 67.000 30.600 ;
        RECT 67.800 30.400 68.400 31.800 ;
        RECT 74.800 31.200 75.400 31.800 ;
        RECT 79.600 31.200 80.200 31.800 ;
        RECT 74.800 30.400 76.000 31.200 ;
        RECT 79.600 30.400 80.800 31.200 ;
        RECT 46.000 30.300 46.800 30.400 ;
        RECT 43.000 29.700 46.800 30.300 ;
        RECT 36.400 26.200 37.200 26.800 ;
        RECT 17.200 22.200 18.000 25.400 ;
        RECT 34.800 25.400 37.200 26.200 ;
        RECT 18.800 22.200 19.600 25.000 ;
        RECT 20.400 22.200 21.200 25.000 ;
        RECT 22.000 22.200 22.800 25.000 ;
        RECT 25.200 22.200 26.000 25.000 ;
        RECT 28.400 22.200 29.200 25.000 ;
        RECT 30.000 22.200 30.800 25.000 ;
        RECT 31.600 22.200 32.400 25.000 ;
        RECT 33.200 22.200 34.000 25.000 ;
        RECT 34.800 22.200 35.600 25.400 ;
        RECT 41.200 22.200 42.000 27.400 ;
        RECT 43.000 26.800 43.800 29.700 ;
        RECT 46.000 29.600 46.800 29.700 ;
        RECT 48.200 29.800 49.800 30.400 ;
        RECT 48.200 29.600 49.000 29.800 ;
        RECT 50.800 29.600 51.600 30.400 ;
        RECT 49.600 28.600 50.400 28.800 ;
        RECT 47.600 28.400 50.400 28.600 ;
        RECT 46.000 28.000 50.400 28.400 ;
        RECT 51.000 28.400 51.600 29.600 ;
        RECT 64.000 29.800 64.800 30.000 ;
        RECT 67.800 29.800 69.200 30.400 ;
        RECT 73.200 30.300 74.000 30.400 ;
        RECT 64.000 29.200 66.600 29.800 ;
        RECT 66.000 28.600 66.600 29.200 ;
        RECT 67.400 29.600 69.200 29.800 ;
        RECT 71.700 29.700 74.000 30.300 ;
        RECT 67.400 29.200 68.400 29.600 ;
        RECT 46.000 27.800 48.200 28.000 ;
        RECT 51.000 27.800 52.000 28.400 ;
        RECT 46.000 27.600 47.600 27.800 ;
        RECT 47.800 26.800 48.600 27.000 ;
        RECT 42.800 26.000 43.800 26.800 ;
        RECT 46.000 26.200 48.600 26.800 ;
        RECT 49.200 26.400 50.800 27.200 ;
        RECT 42.800 22.200 43.600 26.000 ;
        RECT 46.000 22.200 46.800 26.200 ;
        RECT 51.400 25.800 52.000 27.800 ;
        RECT 52.800 27.600 53.600 28.400 ;
        RECT 54.800 27.600 56.400 28.400 ;
        RECT 62.000 28.200 63.600 28.400 ;
        RECT 62.000 27.600 65.400 28.200 ;
        RECT 66.000 27.800 66.800 28.600 ;
        RECT 52.800 27.200 53.400 27.600 ;
        RECT 52.600 26.400 53.400 27.200 ;
        RECT 64.800 27.200 65.400 27.600 ;
        RECT 54.000 26.800 54.800 27.000 ;
        RECT 63.400 26.800 64.200 27.000 ;
        RECT 54.000 26.200 56.400 26.800 ;
        RECT 50.400 22.200 52.000 25.800 ;
        RECT 55.600 22.200 56.400 26.200 ;
        RECT 62.000 26.200 64.200 26.800 ;
        RECT 64.800 26.600 66.800 27.200 ;
        RECT 65.200 26.400 66.800 26.600 ;
        RECT 62.000 22.200 62.800 26.200 ;
        RECT 67.400 25.800 68.000 29.200 ;
        RECT 71.700 28.400 72.300 29.700 ;
        RECT 73.200 28.800 74.000 29.700 ;
        RECT 68.800 27.600 69.600 28.400 ;
        RECT 70.800 27.600 72.400 28.400 ;
        RECT 68.800 27.200 69.400 27.600 ;
        RECT 74.800 27.400 75.400 30.400 ;
        RECT 79.600 27.400 80.200 30.400 ;
        RECT 68.600 26.400 69.400 27.200 ;
        RECT 70.000 26.800 70.800 27.000 ;
        RECT 73.200 26.800 75.400 27.400 ;
        RECT 78.000 26.800 80.200 27.400 ;
        RECT 70.000 26.200 72.400 26.800 ;
        RECT 66.400 24.400 68.000 25.800 ;
        RECT 65.200 23.600 68.000 24.400 ;
        RECT 66.400 22.200 68.000 23.600 ;
        RECT 71.600 22.200 72.400 26.200 ;
        RECT 73.200 22.200 74.000 26.800 ;
        RECT 78.000 22.200 78.800 26.800 ;
        RECT 1.200 13.800 2.000 19.800 ;
        RECT 7.600 16.600 8.400 19.800 ;
        RECT 9.200 17.000 10.000 19.800 ;
        RECT 10.800 17.000 11.600 19.800 ;
        RECT 12.400 17.000 13.200 19.800 ;
        RECT 15.600 17.000 16.400 19.800 ;
        RECT 18.800 17.000 19.600 19.800 ;
        RECT 20.400 17.000 21.200 19.800 ;
        RECT 22.000 17.000 22.800 19.800 ;
        RECT 23.600 17.000 24.400 19.800 ;
        RECT 5.800 15.800 8.400 16.600 ;
        RECT 25.200 16.600 26.000 19.800 ;
        RECT 11.800 15.800 16.400 16.400 ;
        RECT 5.800 15.200 6.600 15.800 ;
        RECT 3.600 14.400 6.600 15.200 ;
        RECT 1.200 13.000 10.000 13.800 ;
        RECT 11.800 13.400 12.600 15.800 ;
        RECT 15.600 15.600 16.400 15.800 ;
        RECT 21.800 15.600 22.800 16.400 ;
        RECT 25.200 15.800 27.600 16.600 ;
        RECT 14.000 13.600 14.800 15.200 ;
        RECT 15.600 14.800 16.400 15.000 ;
        RECT 15.600 14.200 20.000 14.800 ;
        RECT 19.200 14.000 20.000 14.200 ;
        RECT 1.200 7.400 2.000 13.000 ;
        RECT 10.600 12.600 12.600 13.400 ;
        RECT 16.400 12.600 19.600 13.400 ;
        RECT 22.000 12.800 22.800 15.600 ;
        RECT 26.800 15.200 27.600 15.800 ;
        RECT 26.800 14.600 28.600 15.200 ;
        RECT 27.800 13.400 28.600 14.600 ;
        RECT 31.600 14.600 32.400 19.800 ;
        RECT 33.200 16.000 34.000 19.800 ;
        RECT 33.200 15.200 34.200 16.000 ;
        RECT 31.600 14.000 32.800 14.600 ;
        RECT 27.800 12.600 31.600 13.400 ;
        RECT 2.600 12.000 3.400 12.200 ;
        RECT 7.600 12.000 8.400 12.400 ;
        RECT 25.200 12.000 26.000 12.600 ;
        RECT 32.200 12.000 32.800 14.000 ;
        RECT 2.600 11.400 26.000 12.000 ;
        RECT 32.000 11.400 32.800 12.000 ;
        RECT 32.000 9.600 32.600 11.400 ;
        RECT 33.400 10.800 34.200 15.200 ;
        RECT 34.800 14.300 35.600 14.400 ;
        RECT 41.200 14.300 42.000 19.800 ;
        RECT 42.800 16.300 43.600 17.200 ;
        RECT 46.000 16.300 46.800 16.400 ;
        RECT 42.800 15.700 46.800 16.300 ;
        RECT 42.800 15.600 43.600 15.700 ;
        RECT 46.000 15.600 46.800 15.700 ;
        RECT 34.800 13.700 42.000 14.300 ;
        RECT 34.800 13.600 35.600 13.700 ;
        RECT 10.800 9.400 11.600 9.600 ;
        RECT 6.200 9.000 11.600 9.400 ;
        RECT 5.400 8.800 11.600 9.000 ;
        RECT 12.600 9.000 21.200 9.600 ;
        RECT 2.800 8.000 4.400 8.800 ;
        RECT 5.400 8.200 6.800 8.800 ;
        RECT 12.600 8.200 13.200 9.000 ;
        RECT 20.400 8.800 21.200 9.000 ;
        RECT 23.600 9.000 32.600 9.600 ;
        RECT 23.600 8.800 24.400 9.000 ;
        RECT 3.800 7.600 4.400 8.000 ;
        RECT 7.400 7.600 13.200 8.200 ;
        RECT 13.800 7.600 16.400 8.400 ;
        RECT 1.200 6.800 3.200 7.400 ;
        RECT 3.800 6.800 8.000 7.600 ;
        RECT 2.600 6.200 3.200 6.800 ;
        RECT 2.600 5.600 3.600 6.200 ;
        RECT 2.800 2.200 3.600 5.600 ;
        RECT 6.000 2.200 6.800 6.800 ;
        RECT 9.200 2.200 10.000 5.000 ;
        RECT 10.800 2.200 11.600 5.000 ;
        RECT 12.400 2.200 13.200 7.000 ;
        RECT 15.600 2.200 16.400 7.000 ;
        RECT 18.800 2.200 19.600 8.400 ;
        RECT 26.800 7.600 29.400 8.400 ;
        RECT 22.000 6.800 26.200 7.600 ;
        RECT 20.400 2.200 21.200 5.000 ;
        RECT 22.000 2.200 22.800 5.000 ;
        RECT 23.600 2.200 24.400 5.000 ;
        RECT 26.800 2.200 27.600 7.600 ;
        RECT 32.000 7.400 32.600 9.000 ;
        RECT 30.000 6.800 32.600 7.400 ;
        RECT 33.200 10.000 34.200 10.800 ;
        RECT 30.000 2.200 30.800 6.800 ;
        RECT 33.200 2.200 34.000 10.000 ;
        RECT 41.200 2.200 42.000 13.700 ;
        RECT 49.200 13.800 50.000 19.800 ;
        RECT 55.600 16.600 56.400 19.800 ;
        RECT 57.200 17.000 58.000 19.800 ;
        RECT 58.800 17.000 59.600 19.800 ;
        RECT 60.400 17.000 61.200 19.800 ;
        RECT 63.600 17.000 64.400 19.800 ;
        RECT 66.800 17.000 67.600 19.800 ;
        RECT 68.400 17.000 69.200 19.800 ;
        RECT 70.000 17.000 70.800 19.800 ;
        RECT 71.600 17.000 72.400 19.800 ;
        RECT 53.800 15.800 56.400 16.600 ;
        RECT 73.200 16.600 74.000 19.800 ;
        RECT 59.800 15.800 64.400 16.400 ;
        RECT 53.800 15.200 54.600 15.800 ;
        RECT 51.600 14.400 54.600 15.200 ;
        RECT 49.200 13.000 58.000 13.800 ;
        RECT 59.800 13.400 60.600 15.800 ;
        RECT 63.600 15.600 64.400 15.800 ;
        RECT 69.800 15.600 70.800 16.400 ;
        RECT 73.200 15.800 75.600 16.600 ;
        RECT 62.000 13.600 62.800 15.200 ;
        RECT 63.600 14.800 64.400 15.000 ;
        RECT 63.600 14.200 68.000 14.800 ;
        RECT 67.200 14.000 68.000 14.200 ;
        RECT 49.200 7.400 50.000 13.000 ;
        RECT 58.600 12.600 60.600 13.400 ;
        RECT 64.400 12.600 67.600 13.400 ;
        RECT 70.000 12.800 70.800 15.600 ;
        RECT 74.800 15.200 75.600 15.800 ;
        RECT 74.800 14.600 76.600 15.200 ;
        RECT 75.800 13.400 76.600 14.600 ;
        RECT 79.600 14.600 80.400 19.800 ;
        RECT 81.200 16.000 82.000 19.800 ;
        RECT 81.200 15.200 82.200 16.000 ;
        RECT 79.600 14.000 80.800 14.600 ;
        RECT 75.800 12.600 79.600 13.400 ;
        RECT 50.600 12.000 51.400 12.200 ;
        RECT 52.400 12.000 53.200 12.400 ;
        RECT 55.600 12.000 56.400 12.400 ;
        RECT 73.200 12.000 74.000 12.600 ;
        RECT 80.200 12.000 80.800 14.000 ;
        RECT 50.600 11.400 74.000 12.000 ;
        RECT 80.000 11.400 80.800 12.000 ;
        RECT 80.000 9.600 80.600 11.400 ;
        RECT 81.400 10.800 82.200 15.200 ;
        RECT 58.800 9.400 59.600 9.600 ;
        RECT 54.200 9.000 59.600 9.400 ;
        RECT 53.400 8.800 59.600 9.000 ;
        RECT 60.600 9.000 69.200 9.600 ;
        RECT 50.800 8.000 52.400 8.800 ;
        RECT 53.400 8.200 54.800 8.800 ;
        RECT 60.600 8.200 61.200 9.000 ;
        RECT 68.400 8.800 69.200 9.000 ;
        RECT 71.600 9.000 80.600 9.600 ;
        RECT 71.600 8.800 72.400 9.000 ;
        RECT 51.800 7.600 52.400 8.000 ;
        RECT 55.400 7.600 61.200 8.200 ;
        RECT 61.800 7.600 64.400 8.400 ;
        RECT 49.200 6.800 51.200 7.400 ;
        RECT 51.800 6.800 56.000 7.600 ;
        RECT 50.600 6.200 51.200 6.800 ;
        RECT 50.600 5.600 51.600 6.200 ;
        RECT 50.800 2.200 51.600 5.600 ;
        RECT 54.000 2.200 54.800 6.800 ;
        RECT 57.200 2.200 58.000 5.000 ;
        RECT 58.800 2.200 59.600 5.000 ;
        RECT 60.400 2.200 61.200 7.000 ;
        RECT 63.600 2.200 64.400 7.000 ;
        RECT 66.800 2.200 67.600 8.400 ;
        RECT 74.800 7.600 77.400 8.400 ;
        RECT 70.000 6.800 74.200 7.600 ;
        RECT 68.400 2.200 69.200 5.000 ;
        RECT 70.000 2.200 70.800 5.000 ;
        RECT 71.600 2.200 72.400 5.000 ;
        RECT 74.800 2.200 75.600 7.600 ;
        RECT 80.000 7.400 80.600 9.000 ;
        RECT 78.000 6.800 80.600 7.400 ;
        RECT 81.200 10.000 82.200 10.800 ;
        RECT 78.000 2.200 78.800 6.800 ;
        RECT 81.200 2.200 82.000 10.000 ;
      LAYER via1 ;
        RECT 17.200 53.000 18.000 53.800 ;
        RECT 26.800 52.600 27.600 53.400 ;
        RECT 12.400 51.600 13.200 52.400 ;
        RECT 46.000 53.600 46.800 54.400 ;
        RECT 18.800 48.800 19.600 49.600 ;
        RECT 23.600 47.600 24.400 48.400 ;
        RECT 20.400 46.200 21.200 47.000 ;
        RECT 17.200 44.200 18.000 45.000 ;
        RECT 18.800 44.200 19.600 45.000 ;
        RECT 23.600 46.200 24.400 47.000 ;
        RECT 26.800 46.200 27.600 47.000 ;
        RECT 28.400 44.200 29.200 45.000 ;
        RECT 30.000 44.200 30.800 45.000 ;
        RECT 31.600 44.200 32.400 45.000 ;
        RECT 41.200 47.600 42.000 48.400 ;
        RECT 66.800 51.600 67.600 52.400 ;
        RECT 28.400 35.000 29.200 35.800 ;
        RECT 25.200 33.600 26.000 34.400 ;
        RECT 30.000 32.400 30.800 33.200 ;
        RECT 47.800 31.800 48.600 32.600 ;
        RECT 63.400 31.800 64.200 32.600 ;
        RECT 18.800 28.200 19.600 29.000 ;
        RECT 28.400 28.600 29.200 29.400 ;
        RECT 23.600 27.600 24.400 28.400 ;
        RECT 18.800 24.200 19.600 25.000 ;
        RECT 20.400 24.200 21.200 25.000 ;
        RECT 22.000 24.200 22.800 25.000 ;
        RECT 25.200 24.200 26.000 25.000 ;
        RECT 28.400 24.200 29.200 25.000 ;
        RECT 30.000 24.200 30.800 25.000 ;
        RECT 31.600 24.200 32.400 25.000 ;
        RECT 33.200 24.200 34.000 25.000 ;
        RECT 49.000 29.800 49.800 30.600 ;
        RECT 47.800 26.200 48.600 27.000 ;
        RECT 55.600 27.600 56.400 28.400 ;
        RECT 50.800 23.600 51.600 24.400 ;
        RECT 63.400 26.200 64.200 27.000 ;
        RECT 73.200 29.600 74.000 30.400 ;
        RECT 9.200 13.000 10.000 13.800 ;
        RECT 18.800 12.600 19.600 13.400 ;
        RECT 33.200 17.600 34.000 18.400 ;
        RECT 7.600 11.600 8.400 12.400 ;
        RECT 25.200 11.600 26.000 12.400 ;
        RECT 10.800 8.800 11.600 9.600 ;
        RECT 15.600 7.600 16.400 8.400 ;
        RECT 12.400 6.200 13.200 7.000 ;
        RECT 9.200 4.200 10.000 5.000 ;
        RECT 10.800 4.200 11.600 5.000 ;
        RECT 15.600 6.200 16.400 7.000 ;
        RECT 18.800 6.200 19.600 7.000 ;
        RECT 20.400 4.200 21.200 5.000 ;
        RECT 22.000 4.200 22.800 5.000 ;
        RECT 23.600 4.200 24.400 5.000 ;
        RECT 57.200 13.000 58.000 13.800 ;
        RECT 66.800 12.600 67.600 13.400 ;
        RECT 81.200 17.600 82.000 18.400 ;
        RECT 52.400 11.600 53.200 12.400 ;
        RECT 58.800 8.800 59.600 9.600 ;
        RECT 63.600 7.600 64.400 8.400 ;
        RECT 60.400 6.200 61.200 7.000 ;
        RECT 57.200 4.200 58.000 5.000 ;
        RECT 58.800 4.200 59.600 5.000 ;
        RECT 63.600 6.200 64.400 7.000 ;
        RECT 66.800 6.200 67.600 7.000 ;
        RECT 68.400 4.200 69.200 5.000 ;
        RECT 70.000 4.200 70.800 5.000 ;
        RECT 71.600 4.200 72.400 5.000 ;
      LAYER metal2 ;
        RECT 7.600 51.600 8.400 52.400 ;
        RECT 12.400 51.600 13.200 52.400 ;
        RECT 7.700 30.400 8.300 51.600 ;
        RECT 17.200 44.200 18.000 57.800 ;
        RECT 18.800 44.200 19.600 57.800 ;
        RECT 20.400 46.200 21.200 57.800 ;
        RECT 22.000 53.600 22.800 54.400 ;
        RECT 23.600 46.200 24.400 57.800 ;
        RECT 26.800 46.200 27.600 57.800 ;
        RECT 28.400 44.200 29.200 57.800 ;
        RECT 30.000 44.200 30.800 57.800 ;
        RECT 31.600 44.200 32.400 57.800 ;
        RECT 49.200 55.600 50.000 56.400 ;
        RECT 46.000 53.600 46.800 54.400 ;
        RECT 46.100 52.400 46.700 53.600 ;
        RECT 44.400 51.600 45.200 52.400 ;
        RECT 46.000 51.600 46.800 52.400 ;
        RECT 44.500 50.400 45.100 51.600 ;
        RECT 44.400 49.600 45.200 50.400 ;
        RECT 41.200 47.600 42.000 48.400 ;
        RECT 7.600 29.600 8.400 30.400 ;
        RECT 14.000 29.600 14.800 30.400 ;
        RECT 7.700 12.400 8.300 29.600 ;
        RECT 18.800 24.200 19.600 37.800 ;
        RECT 20.400 24.200 21.200 37.800 ;
        RECT 22.000 24.200 22.800 35.800 ;
        RECT 23.600 27.600 24.400 28.400 ;
        RECT 23.700 24.400 24.300 27.600 ;
        RECT 23.600 23.600 24.400 24.400 ;
        RECT 25.200 24.200 26.000 35.800 ;
        RECT 28.400 24.200 29.200 35.800 ;
        RECT 30.000 24.200 30.800 37.800 ;
        RECT 31.600 24.200 32.400 37.800 ;
        RECT 33.200 24.200 34.000 37.800 ;
        RECT 44.500 28.300 45.100 49.600 ;
        RECT 46.100 30.400 46.700 51.600 ;
        RECT 49.300 48.400 49.900 55.600 ;
        RECT 52.400 53.600 53.200 54.400 ;
        RECT 55.600 51.600 56.400 52.400 ;
        RECT 66.800 51.600 67.600 52.400 ;
        RECT 74.800 51.600 75.600 52.400 ;
        RECT 79.600 51.600 80.400 52.400 ;
        RECT 49.200 47.600 50.000 48.400 ;
        RECT 47.800 31.800 48.600 32.600 ;
        RECT 54.000 31.800 54.800 32.600 ;
        RECT 46.000 29.600 46.800 30.400 ;
        RECT 46.000 28.300 46.800 28.400 ;
        RECT 44.500 27.700 46.800 28.300 ;
        RECT 46.000 27.600 46.800 27.700 ;
        RECT 46.100 18.400 46.700 27.600 ;
        RECT 47.800 27.000 48.400 31.800 ;
        RECT 49.000 29.800 49.800 30.600 ;
        RECT 49.200 28.400 49.800 29.800 ;
        RECT 54.200 28.400 54.800 31.800 ;
        RECT 55.700 28.400 56.300 51.600 ;
        RECT 66.800 49.600 67.600 50.400 ;
        RECT 79.700 48.400 80.300 51.600 ;
        RECT 65.200 47.600 66.000 48.400 ;
        RECT 79.600 47.600 80.400 48.400 ;
        RECT 62.000 43.600 62.800 44.400 ;
        RECT 62.100 28.400 62.700 43.600 ;
        RECT 63.400 31.800 64.200 32.600 ;
        RECT 70.000 31.800 70.800 32.600 ;
        RECT 49.200 27.800 54.800 28.400 ;
        RECT 49.200 27.000 50.000 27.200 ;
        RECT 52.600 27.000 53.400 27.200 ;
        RECT 54.200 27.000 54.800 27.800 ;
        RECT 55.600 27.600 56.400 28.400 ;
        RECT 62.000 27.600 62.800 28.400 ;
        RECT 47.800 26.400 53.400 27.000 ;
        RECT 47.800 26.200 48.600 26.400 ;
        RECT 54.000 26.200 54.800 27.000 ;
        RECT 63.400 27.000 64.000 31.800 ;
        RECT 66.000 28.400 66.800 28.600 ;
        RECT 70.200 28.400 70.800 31.800 ;
        RECT 73.200 29.600 74.000 30.400 ;
        RECT 66.000 27.800 70.800 28.400 ;
        RECT 65.200 27.000 66.000 27.200 ;
        RECT 68.600 27.000 69.400 27.200 ;
        RECT 70.200 27.000 70.800 27.800 ;
        RECT 63.400 26.200 64.200 27.000 ;
        RECT 65.200 26.400 69.400 27.000 ;
        RECT 70.000 26.200 70.800 27.000 ;
        RECT 50.800 23.600 51.600 24.400 ;
        RECT 65.200 23.600 66.000 24.400 ;
        RECT 65.300 18.400 65.900 23.600 ;
        RECT 73.300 18.400 73.900 29.600 ;
        RECT 7.600 11.600 8.400 12.400 ;
        RECT 9.200 4.200 10.000 17.800 ;
        RECT 10.800 4.200 11.600 17.800 ;
        RECT 12.400 6.200 13.200 17.800 ;
        RECT 14.000 13.600 14.800 14.400 ;
        RECT 15.600 6.200 16.400 17.800 ;
        RECT 18.800 6.200 19.600 17.800 ;
        RECT 20.400 4.200 21.200 17.800 ;
        RECT 22.000 4.200 22.800 17.800 ;
        RECT 23.600 4.200 24.400 17.800 ;
        RECT 33.200 17.600 34.000 18.400 ;
        RECT 46.000 17.600 46.800 18.400 ;
        RECT 46.100 16.400 46.700 17.600 ;
        RECT 46.000 15.600 46.800 16.400 ;
        RECT 34.800 13.600 35.600 14.400 ;
        RECT 25.200 11.600 26.000 12.400 ;
        RECT 52.400 11.600 53.200 12.400 ;
        RECT 57.200 4.200 58.000 17.800 ;
        RECT 58.800 4.200 59.600 17.800 ;
        RECT 60.400 6.200 61.200 17.800 ;
        RECT 62.000 17.600 62.800 18.400 ;
        RECT 62.100 14.400 62.700 17.600 ;
        RECT 62.000 13.600 62.800 14.400 ;
        RECT 63.600 6.200 64.400 17.800 ;
        RECT 65.200 17.600 66.000 18.400 ;
        RECT 66.800 6.200 67.600 17.800 ;
        RECT 68.400 4.200 69.200 17.800 ;
        RECT 70.000 4.200 70.800 17.800 ;
        RECT 71.600 4.200 72.400 17.800 ;
        RECT 73.200 17.600 74.000 18.400 ;
        RECT 81.200 17.600 82.000 18.400 ;
      LAYER metal3 ;
        RECT 22.000 54.300 22.800 54.400 ;
        RECT 52.400 54.300 53.200 54.400 ;
        RECT 22.000 53.700 53.200 54.300 ;
        RECT 22.000 53.600 22.800 53.700 ;
        RECT 52.400 53.600 53.200 53.700 ;
        RECT 7.600 52.300 8.400 52.400 ;
        RECT 12.400 52.300 13.200 52.400 ;
        RECT 7.600 51.700 13.200 52.300 ;
        RECT 7.600 51.600 8.400 51.700 ;
        RECT 12.400 51.600 13.200 51.700 ;
        RECT 46.000 52.300 46.800 52.400 ;
        RECT 55.600 52.300 56.400 52.400 ;
        RECT 66.800 52.300 67.600 52.400 ;
        RECT 74.800 52.300 75.600 52.400 ;
        RECT 46.000 51.700 75.600 52.300 ;
        RECT 46.000 51.600 46.800 51.700 ;
        RECT 55.600 51.600 56.400 51.700 ;
        RECT 66.800 51.600 67.600 51.700 ;
        RECT 74.800 51.600 75.600 51.700 ;
        RECT 44.400 50.300 45.200 50.400 ;
        RECT 66.800 50.300 67.600 50.400 ;
        RECT 44.400 49.700 67.600 50.300 ;
        RECT 44.400 49.600 45.200 49.700 ;
        RECT 66.800 49.600 67.600 49.700 ;
        RECT 41.200 48.300 42.000 48.400 ;
        RECT 49.200 48.300 50.000 48.400 ;
        RECT 65.200 48.300 66.000 48.400 ;
        RECT 79.600 48.300 80.400 48.400 ;
        RECT 41.200 47.700 80.400 48.300 ;
        RECT 41.200 47.600 42.000 47.700 ;
        RECT 49.200 47.600 50.000 47.700 ;
        RECT 65.200 47.600 66.000 47.700 ;
        RECT 79.600 47.600 80.400 47.700 ;
        RECT 7.600 30.300 8.400 30.400 ;
        RECT 14.000 30.300 14.800 30.400 ;
        RECT 7.600 29.700 14.800 30.300 ;
        RECT 7.600 29.600 8.400 29.700 ;
        RECT 14.000 29.600 14.800 29.700 ;
        RECT 23.600 24.300 24.400 24.400 ;
        RECT 50.800 24.300 51.600 24.400 ;
        RECT 23.600 23.700 51.600 24.300 ;
        RECT 23.600 23.600 24.400 23.700 ;
        RECT 50.800 23.600 51.600 23.700 ;
        RECT 33.200 18.300 34.000 18.400 ;
        RECT 46.000 18.300 46.800 18.400 ;
        RECT 33.200 17.700 46.800 18.300 ;
        RECT 33.200 17.600 34.000 17.700 ;
        RECT 46.000 17.600 46.800 17.700 ;
        RECT 62.000 18.300 62.800 18.400 ;
        RECT 65.200 18.300 66.000 18.400 ;
        RECT 62.000 17.700 66.000 18.300 ;
        RECT 62.000 17.600 62.800 17.700 ;
        RECT 65.200 17.600 66.000 17.700 ;
        RECT 73.200 18.300 74.000 18.400 ;
        RECT 81.200 18.300 82.000 18.400 ;
        RECT 73.200 17.700 82.000 18.300 ;
        RECT 73.200 17.600 74.000 17.700 ;
        RECT 81.200 17.600 82.000 17.700 ;
        RECT 14.000 14.300 14.800 14.400 ;
        RECT 34.800 14.300 35.600 14.400 ;
        RECT 14.000 13.700 35.600 14.300 ;
        RECT 14.000 13.600 14.800 13.700 ;
        RECT 34.800 13.600 35.600 13.700 ;
        RECT 25.200 12.300 26.000 12.400 ;
        RECT 52.400 12.300 53.200 12.400 ;
        RECT 25.200 11.700 53.200 12.300 ;
        RECT 25.200 11.600 26.000 11.700 ;
        RECT 52.400 11.600 53.200 11.700 ;
  END
END counter
END LIBRARY


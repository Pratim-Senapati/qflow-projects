* NGSPICE file created from cordic.ext - technology: scmos

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

.subckt cordic vdd gnd clk rst theta[0] theta[1] theta[2] theta[3] theta[4] theta[5]
+ theta[6] theta[7] theta[8] theta[9] theta[10] theta[11] theta[12] theta[13] theta[14]
+ theta[15] sine[0] sine[1] sine[2] sine[3] sine[4] sine[5] sine[6] sine[7] sine[8]
+ sine[9] sine[10] sine[11] sine[12] sine[13] sine[14] sine[15] cosine[0] cosine[1]
+ cosine[2] cosine[3] cosine[4] cosine[5] cosine[6] cosine[7] cosine[8] cosine[9]
+ cosine[10] cosine[11] cosine[12] cosine[13] cosine[14] cosine[15]
XAND2X2_5 BUFX2_27/A DFFSR_12/Q gnd AND2X2_5/Y vdd AND2X2
XFILL_5_1_2 gnd vdd FILL
XNAND2X1_10 DFFSR_9/Q AND2X2_4/Y gnd XNOR2X1_7/A vdd NAND2X1
XDFFSR_9 DFFSR_9/Q DFFSR_9/CLK DFFSR_9/R vdd DFFSR_9/D gnd vdd DFFSR
XFILL_8_1_0 gnd vdd FILL
XXNOR2X1_6 AND2X2_4/Y INVX1_11/Y gnd DFFSR_9/D vdd XNOR2X1
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XAND2X2_6 AND2X2_6/A AND2X2_5/Y gnd AND2X2_6/Y vdd AND2X2
XNAND2X1_11 AND2X2_6/A AND2X2_4/Y gnd NOR2X1_11/B vdd NAND2X1
XFILL_10_1 gnd vdd FILL
XXNOR2X1_7 XNOR2X1_7/A INVX1_12/A gnd DFFSR_10/D vdd XNOR2X1
XFILL_0_0_1 gnd vdd FILL
XFILL_8_1_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XNAND2X1_12 AND2X2_6/Y AND2X2_4/Y gnd XNOR2X1_9/A vdd NAND2X1
XFILL_10_2 gnd vdd FILL
XFILL_9_1 gnd vdd FILL
XXNOR2X1_8 NOR2X1_11/B BUFX2_27/A gnd DFFSR_11/D vdd XNOR2X1
XFILL_8_1_2 gnd vdd FILL
XINVX8_1 rst gnd BUFX4_1/A vdd INVX8
XFILL_0_0_2 gnd vdd FILL
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XNAND2X1_13 BUFX2_29/A DFFSR_14/Q gnd NOR2X1_12/A vdd NAND2X1
XNOR3X1_1 BUFX2_5/A BUFX2_6/A NOR3X1_1/C gnd NOR3X1_1/Y vdd NOR3X1
XXNOR2X1_9 XNOR2X1_9/A BUFX2_29/A gnd DFFSR_13/D vdd XNOR2X1
XFILL_3_0_0 gnd vdd FILL
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XNAND2X1_14 BUFX2_31/A XOR2X1_5/A gnd XNOR2X1_11/A vdd NAND2X1
XNOR3X1_2 BUFX2_7/A BUFX2_8/A NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XCLKBUF1_1 clk gnd DFFSR_7/CLK vdd CLKBUF1
XFILL_3_0_1 gnd vdd FILL
XNAND2X1_15 NOR3X1_7/C OAI21X1_5/Y gnd DFFSR_18/D vdd NAND2X1
XNOR3X1_3 BUFX2_9/A INVX1_2/A NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XFILL_3_0_2 gnd vdd FILL
XCLKBUF1_2 clk gnd CLKBUF1_2/Y vdd CLKBUF1
XNAND2X1_16 OAI21X1_6/Y NOR3X1_1/C gnd DFFSR_20/D vdd NAND2X1
XFILL_7_1 gnd vdd FILL
XNAND3X1_1 INVX1_21/Y INVX1_22/Y NOR3X1_1/Y gnd NOR3X1_3/C vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XNOR3X1_4 INVX1_3/A INVX1_4/A NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XCLKBUF1_3 clk gnd CLKBUF1_3/Y vdd CLKBUF1
XFILL_6_0_0 gnd vdd FILL
XXOR2X1_1 AND2X2_3/A DFFSR_4/Q gnd DFFSR_4/D vdd XOR2X1
XFILL_7_2 gnd vdd FILL
XNAND3X1_2 INVX1_1/Y INVX1_2/Y NOR3X1_2/Y gnd NOR3X1_4/C vdd NAND3X1
XNAND2X1_17 NOR3X1_2/C OAI21X1_7/Y gnd DFFSR_22/D vdd NAND2X1
XFILL_1_1_1 gnd vdd FILL
XNOR3X1_5 INVX1_5/A INVX1_6/A NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XCLKBUF1_4 clk gnd DFFSR_9/CLK vdd CLKBUF1
XFILL_6_0_1 gnd vdd FILL
XXOR2X1_2 INVX1_10/A DFFSR_5/Q gnd DFFSR_5/D vdd XOR2X1
XNOR3X1_6 BUFX2_1/A BUFX2_2/A INVX1_16/Y gnd NOR3X1_6/Y vdd NOR3X1
XFILL_1_1_2 gnd vdd FILL
XNAND3X1_3 INVX1_3/Y INVX1_4/Y NOR3X1_3/Y gnd NOR3X1_5/C vdd NAND3X1
XFILL_6_0_2 gnd vdd FILL
XXOR2X1_3 NOR2X1_8/B DFFSR_7/Q gnd DFFSR_7/D vdd XOR2X1
XCLKBUF1_5 clk gnd CLKBUF1_5/Y vdd CLKBUF1
XFILL_4_1_0 gnd vdd FILL
XBUFX4_1 BUFX4_1/A gnd DFFSR_3/R vdd BUFX4
XFILL_9_0_0 gnd vdd FILL
XNOR3X1_7 BUFX2_3/A BUFX2_4/A NOR3X1_7/C gnd NOR3X1_7/Y vdd NOR3X1
XOAI21X1_1 BUFX2_9/A NOR3X1_3/C INVX1_2/A gnd OAI21X1_1/Y vdd OAI21X1
XNAND3X1_4 INVX1_5/Y INVX1_6/Y NOR3X1_4/Y gnd OAI21X1_4/B vdd NAND3X1
XXOR2X1_4 XOR2X1_4/A DFFSR_12/Q gnd XOR2X1_4/Y vdd XOR2X1
XFILL_4_1_1 gnd vdd FILL
XBUFX4_2 BUFX4_1/A gnd BUFX4_2/Y vdd BUFX4
XNAND3X1_5 INVX1_7/Y INVX1_8/Y NOR3X1_5/Y gnd NAND3X1_5/Y vdd NAND3X1
XFILL_9_0_1 gnd vdd FILL
XXOR2X1_5 XOR2X1_5/A BUFX2_31/A gnd XOR2X1_5/Y vdd XOR2X1
XOAI21X1_2 INVX1_3/A NOR3X1_4/C INVX1_4/A gnd NAND2X1_3/A vdd OAI21X1
XBUFX4_3 BUFX4_1/A gnd BUFX4_3/Y vdd BUFX4
XFILL_4_1_2 gnd vdd FILL
XNAND3X1_6 BUFX2_29/A AND2X2_6/Y AND2X2_4/Y gnd NAND3X1_6/Y vdd NAND3X1
XFILL_9_0_2 gnd vdd FILL
XXOR2X1_6 BUFX2_1/A INVX1_16/A gnd DFFSR_17/D vdd XOR2X1
XOAI21X1_3 INVX1_5/A NOR3X1_5/C INVX1_6/A gnd OAI21X1_3/Y vdd OAI21X1
XFILL_7_1_0 gnd vdd FILL
XNAND3X1_7 INVX1_16/A INVX1_14/Y INVX1_15/Y gnd NOR3X1_7/C vdd NAND3X1
XBUFX2_1 BUFX2_1/A gnd cosine[0] vdd BUFX2
XBUFX4_4 BUFX4_1/A gnd DFFSR_9/R vdd BUFX4
XBUFX2_30 DFFSR_14/Q gnd sine[13] vdd BUFX2
XOAI21X1_4 INVX1_7/A OAI21X1_4/B INVX1_8/A gnd OAI21X1_4/Y vdd OAI21X1
XAOI21X1_1 INVX1_10/A DFFSR_5/Q DFFSR_6/Q gnd NOR2X1_8/A vdd AOI21X1
XFILL_7_1_1 gnd vdd FILL
XBUFX4_5 BUFX4_1/A gnd DFFSR_7/R vdd BUFX4
XBUFX2_2 BUFX2_2/A gnd cosine[1] vdd BUFX2
XNAND3X1_8 INVX1_17/Y INVX1_18/Y NOR3X1_6/Y gnd NOR3X1_1/C vdd NAND3X1
XBUFX2_31 BUFX2_31/A gnd sine[14] vdd BUFX2
XXNOR2X1_10 NAND3X1_6/Y DFFSR_14/Q gnd DFFSR_14/D vdd XNOR2X1
XBUFX2_20 DFFSR_4/Q gnd sine[3] vdd BUFX2
XOAI21X1_5 BUFX2_1/A INVX1_16/Y BUFX2_2/A gnd OAI21X1_5/Y vdd OAI21X1
XFILL_7_1_2 gnd vdd FILL
XBUFX2_3 BUFX2_3/A gnd cosine[2] vdd BUFX2
XNAND3X1_9 INVX1_19/Y INVX1_20/Y NOR3X1_7/Y gnd NOR3X1_2/C vdd NAND3X1
XOAI21X1_6 BUFX2_3/A NOR3X1_7/C BUFX2_4/A gnd OAI21X1_6/Y vdd OAI21X1
XXNOR2X1_11 XNOR2X1_11/A INVX1_16/A gnd DFFSR_16/D vdd XNOR2X1
XBUFX2_32 INVX1_16/A gnd sine[15] vdd BUFX2
XBUFX2_10 INVX1_2/A gnd cosine[9] vdd BUFX2
XBUFX2_21 DFFSR_5/Q gnd sine[4] vdd BUFX2
XNOR2X1_1 INVX1_8/A DFFSR_1/Q gnd NOR2X1_1/Y vdd NOR2X1
XFILL_2_0_0 gnd vdd FILL
XXNOR2X1_12 NOR3X1_7/C BUFX2_3/A gnd DFFSR_19/D vdd XNOR2X1
XBUFX2_4 BUFX2_4/A gnd cosine[3] vdd BUFX2
XNOR2X1_2 NOR2X1_1/Y NOR2X1_2/B gnd DFFSR_1/D vdd NOR2X1
XBUFX2_22 DFFSR_6/Q gnd sine[5] vdd BUFX2
XBUFX2_11 INVX1_3/A gnd cosine[10] vdd BUFX2
XOAI21X1_7 BUFX2_5/A NOR3X1_1/C BUFX2_6/A gnd OAI21X1_7/Y vdd OAI21X1
XFILL_1_1 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XBUFX2_5 BUFX2_5/A gnd cosine[4] vdd BUFX2
XXNOR2X1_13 NOR3X1_1/C BUFX2_5/A gnd DFFSR_21/D vdd XNOR2X1
XBUFX2_23 DFFSR_7/Q gnd sine[6] vdd BUFX2
XBUFX2_12 INVX1_4/A gnd cosine[11] vdd BUFX2
XNOR2X1_3 DFFSR_2/Q NOR2X1_2/B gnd NOR2X1_3/Y vdd NOR2X1
XOAI21X1_8 BUFX2_7/A NOR3X1_2/C BUFX2_8/A gnd OAI21X1_8/Y vdd OAI21X1
XFILL_1_2 gnd vdd FILL
XFILL_2_0_2 gnd vdd FILL
XBUFX2_6 BUFX2_6/A gnd cosine[5] vdd BUFX2
XXNOR2X1_14 NOR3X1_2/C BUFX2_7/A gnd DFFSR_23/D vdd XNOR2X1
XBUFX2_24 DFFSR_8/Q gnd sine[7] vdd BUFX2
XBUFX2_13 INVX1_5/A gnd cosine[12] vdd BUFX2
XFILL_0_1_0 gnd vdd FILL
XNAND2X1_1 OAI21X1_8/Y NOR3X1_3/C gnd DFFSR_24/D vdd NAND2X1
XNOR2X1_4 NOR2X1_3/Y INVX1_9/Y gnd DFFSR_2/D vdd NOR2X1
XFILL_5_0_0 gnd vdd FILL
XFILL_1_3 gnd vdd FILL
XBUFX2_25 DFFSR_9/Q gnd sine[8] vdd BUFX2
XBUFX2_7 BUFX2_7/A gnd cosine[6] vdd BUFX2
XBUFX2_14 INVX1_6/A gnd cosine[13] vdd BUFX2
XFILL_0_1_1 gnd vdd FILL
XNAND2X1_2 NOR3X1_4/C OAI21X1_1/Y gnd DFFSR_26/D vdd NAND2X1
XNOR2X1_5 DFFSR_3/Q INVX1_9/Y gnd NOR2X1_6/A vdd NOR2X1
XFILL_5_0_1 gnd vdd FILL
XNAND2X1_3 NAND2X1_3/A NOR3X1_5/C gnd DFFSR_28/D vdd NAND2X1
XFILL_0_1_2 gnd vdd FILL
XBUFX2_8 BUFX2_8/A gnd cosine[7] vdd BUFX2
XBUFX2_26 INVX1_12/A gnd sine[9] vdd BUFX2
XBUFX2_15 INVX1_7/A gnd cosine[14] vdd BUFX2
XNOR2X1_6 NOR2X1_6/A AND2X2_3/A gnd DFFSR_3/D vdd NOR2X1
XFILL_5_0_2 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XBUFX2_27 BUFX2_27/A gnd sine[10] vdd BUFX2
XNOR2X1_7 NOR2X1_7/A NOR2X1_7/B gnd NOR2X1_8/B vdd NOR2X1
XBUFX2_9 BUFX2_9/A gnd cosine[8] vdd BUFX2
XBUFX2_16 INVX1_8/A gnd cosine[15] vdd BUFX2
XNAND2X1_4 OAI21X1_4/B OAI21X1_3/Y gnd DFFSR_30/D vdd NAND2X1
XFILL_8_0_0 gnd vdd FILL
XNAND2X1_5 OAI21X1_4/Y NAND3X1_5/Y gnd DFFSR_32/D vdd NAND2X1
XFILL_3_1_1 gnd vdd FILL
XBUFX2_28 DFFSR_12/Q gnd sine[11] vdd BUFX2
XFILL_8_0_1 gnd vdd FILL
XINVX1_20 BUFX2_6/A gnd INVX1_20/Y vdd INVX1
XBUFX2_17 DFFSR_1/Q gnd sine[0] vdd BUFX2
XNOR2X1_8 NOR2X1_8/A NOR2X1_8/B gnd DFFSR_6/D vdd NOR2X1
XBUFX2_18 DFFSR_2/Q gnd sine[1] vdd BUFX2
XBUFX2_29 BUFX2_29/A gnd sine[12] vdd BUFX2
XINVX1_21 BUFX2_7/A gnd INVX1_21/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd NOR2X1_7/B vdd INVX1
XNOR2X1_9 NOR2X1_7/A NOR2X1_9/B gnd AND2X2_4/B vdd NOR2X1
XNAND2X1_6 DFFSR_2/Q NOR2X1_2/B gnd INVX1_9/A vdd NAND2X1
XFILL_3_1_2 gnd vdd FILL
XFILL_8_0_2 gnd vdd FILL
XFILL_8_1 gnd vdd FILL
XDFFSR_30 INVX1_6/A CLKBUF1_5/Y vdd DFFSR_3/R DFFSR_30/D gnd vdd DFFSR
XFILL_6_1_0 gnd vdd FILL
XNAND2X1_7 DFFSR_5/Q DFFSR_6/Q gnd NOR2X1_7/A vdd NAND2X1
XINVX1_11 DFFSR_9/Q gnd INVX1_11/Y vdd INVX1
XINVX1_22 BUFX2_8/A gnd INVX1_22/Y vdd INVX1
XBUFX2_19 DFFSR_3/Q gnd sine[2] vdd BUFX2
XDFFSR_20 BUFX2_4/A CLKBUF1_3/Y vdd BUFX4_3/Y DFFSR_20/D gnd vdd DFFSR
XDFFSR_31 INVX1_7/A CLKBUF1_5/Y DFFSR_7/R vdd DFFSR_31/D gnd vdd DFFSR
XFILL_6_1_1 gnd vdd FILL
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XNAND2X1_8 DFFSR_7/Q NOR2X1_8/B gnd XNOR2X1_5/A vdd NAND2X1
XDFFSR_10 INVX1_12/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_10/D gnd vdd DFFSR
XDFFSR_21 BUFX2_5/A CLKBUF1_3/Y vdd BUFX4_3/Y DFFSR_21/D gnd vdd DFFSR
XDFFSR_32 INVX1_8/A CLKBUF1_5/Y DFFSR_7/R vdd DFFSR_32/D gnd vdd DFFSR
XNOR2X1_10 INVX1_11/Y INVX1_12/Y gnd AND2X2_6/A vdd NOR2X1
XFILL_6_1_2 gnd vdd FILL
XINVX1_13 BUFX2_27/A gnd INVX1_13/Y vdd INVX1
XNAND2X1_9 DFFSR_7/Q DFFSR_8/Q gnd NOR2X1_9/B vdd NAND2X1
XFILL_6_1 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XDFFSR_11 BUFX2_27/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_11/D gnd vdd DFFSR
XDFFSR_22 BUFX2_6/A CLKBUF1_3/Y BUFX4_3/Y vdd DFFSR_22/D gnd vdd DFFSR
XFILL_1_0_0 gnd vdd FILL
XINVX1_14 BUFX2_1/A gnd INVX1_14/Y vdd INVX1
XNOR2X1_11 INVX1_13/Y NOR2X1_11/B gnd XOR2X1_4/A vdd NOR2X1
XDFFSR_12 DFFSR_12/Q DFFSR_9/CLK DFFSR_9/R vdd XOR2X1_4/Y gnd vdd DFFSR
XFILL_9_1_1 gnd vdd FILL
XFILL_6_2 gnd vdd FILL
XDFFSR_23 BUFX2_7/A CLKBUF1_2/Y vdd BUFX4_2/Y DFFSR_23/D gnd vdd DFFSR
XFILL_1_0_1 gnd vdd FILL
XNOR2X1_12 NOR2X1_12/A XNOR2X1_9/A gnd XOR2X1_5/A vdd NOR2X1
XINVX1_15 BUFX2_2/A gnd INVX1_15/Y vdd INVX1
XFILL_6_3 gnd vdd FILL
XFILL_9_1_2 gnd vdd FILL
XDFFSR_13 BUFX2_29/A DFFSR_7/CLK DFFSR_7/R vdd DFFSR_13/D gnd vdd DFFSR
XDFFSR_24 BUFX2_8/A CLKBUF1_2/Y vdd BUFX4_2/Y DFFSR_24/D gnd vdd DFFSR
XFILL_1_0_2 gnd vdd FILL
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XDFFSR_1 DFFSR_1/Q CLKBUF1_5/Y DFFSR_3/R vdd DFFSR_1/D gnd vdd DFFSR
XDFFSR_14 DFFSR_14/Q DFFSR_9/CLK DFFSR_9/R vdd DFFSR_14/D gnd vdd DFFSR
XFILL_4_0_0 gnd vdd FILL
XDFFSR_25 BUFX2_9/A CLKBUF1_2/Y BUFX4_2/Y vdd DFFSR_25/D gnd vdd DFFSR
XFILL_4_1 gnd vdd FILL
XINVX1_17 BUFX2_3/A gnd INVX1_17/Y vdd INVX1
XDFFSR_2 DFFSR_2/Q DFFSR_7/CLK DFFSR_3/R vdd DFFSR_2/D gnd vdd DFFSR
XFILL_4_0_1 gnd vdd FILL
XDFFSR_15 BUFX2_31/A DFFSR_9/CLK DFFSR_7/R vdd XOR2X1_5/Y gnd vdd DFFSR
XFILL_4_2 gnd vdd FILL
XDFFSR_26 INVX1_2/A CLKBUF1_2/Y vdd BUFX4_2/Y DFFSR_26/D gnd vdd DFFSR
XDFFSR_3 DFFSR_3/Q CLKBUF1_5/Y DFFSR_3/R vdd DFFSR_3/D gnd vdd DFFSR
XINVX1_18 BUFX2_4/A gnd INVX1_18/Y vdd INVX1
XDFFSR_16 INVX1_16/A CLKBUF1_2/Y BUFX4_3/Y vdd DFFSR_16/D gnd vdd DFFSR
XFILL_4_0_2 gnd vdd FILL
XDFFSR_27 INVX1_3/A CLKBUF1_2/Y vdd BUFX4_2/Y DFFSR_27/D gnd vdd DFFSR
XFILL_4_3 gnd vdd FILL
XINVX1_19 BUFX2_5/A gnd INVX1_19/Y vdd INVX1
XDFFSR_4 DFFSR_4/Q DFFSR_7/CLK DFFSR_3/R vdd DFFSR_4/D gnd vdd DFFSR
XFILL_2_1_0 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XDFFSR_17 BUFX2_1/A CLKBUF1_3/Y vdd BUFX4_3/Y DFFSR_17/D gnd vdd DFFSR
XINVX1_1 BUFX2_9/A gnd INVX1_1/Y vdd INVX1
XXNOR2X1_1 NOR3X1_3/C BUFX2_9/A gnd DFFSR_25/D vdd XNOR2X1
XDFFSR_28 INVX1_4/A CLKBUF1_2/Y BUFX4_2/Y vdd DFFSR_28/D gnd vdd DFFSR
XFILL_2_1 gnd vdd FILL
XAND2X2_1 INVX1_8/A DFFSR_1/Q gnd NOR2X1_2/B vdd AND2X2
XFILL_2_1_1 gnd vdd FILL
XDFFSR_5 DFFSR_5/Q DFFSR_7/CLK DFFSR_3/R vdd DFFSR_5/D gnd vdd DFFSR
XDFFSR_18 BUFX2_2/A CLKBUF1_3/Y DFFSR_9/R vdd DFFSR_18/D gnd vdd DFFSR
XFILL_7_0_1 gnd vdd FILL
XDFFSR_29 INVX1_5/A CLKBUF1_5/Y BUFX4_2/Y vdd DFFSR_29/D gnd vdd DFFSR
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XXNOR2X1_2 NOR3X1_4/C INVX1_3/A gnd DFFSR_27/D vdd XNOR2X1
XAND2X2_2 INVX1_9/Y DFFSR_3/Q gnd AND2X2_3/A vdd AND2X2
XFILL_2_2 gnd vdd FILL
XFILL_2_1_2 gnd vdd FILL
XDFFSR_6 DFFSR_6/Q DFFSR_7/CLK DFFSR_3/R vdd DFFSR_6/D gnd vdd DFFSR
XFILL_7_0_2 gnd vdd FILL
XDFFSR_19 BUFX2_3/A CLKBUF1_3/Y vdd BUFX4_3/Y DFFSR_19/D gnd vdd DFFSR
XXNOR2X1_3 NOR3X1_5/C INVX1_5/A gnd DFFSR_29/D vdd XNOR2X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_5_1_0 gnd vdd FILL
XAND2X2_3 AND2X2_3/A DFFSR_4/Q gnd INVX1_10/A vdd AND2X2
XDFFSR_7 DFFSR_7/Q DFFSR_7/CLK DFFSR_7/R vdd DFFSR_7/D gnd vdd DFFSR
XFILL_5_1_1 gnd vdd FILL
XXNOR2X1_4 OAI21X1_4/B INVX1_7/A gnd DFFSR_31/D vdd XNOR2X1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XDFFSR_8 DFFSR_8/Q DFFSR_7/CLK DFFSR_7/R vdd DFFSR_8/D gnd vdd DFFSR
XAND2X2_4 INVX1_10/A AND2X2_4/B gnd AND2X2_4/Y vdd AND2X2
XXNOR2X1_5 XNOR2X1_5/A DFFSR_8/Q gnd DFFSR_8/D vdd XNOR2X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
.ends

